

module b15_C_gen_AntiSAT_k_128_6 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, 
        U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, 
        U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, 
        U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, 
        U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, 
        U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, 
        U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, 
        U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, 
        U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, 
        U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, 
        U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, 
        U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, 
        U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, 
        U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, 
        U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, 
        U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, 
        U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, 
        U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, 
        U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, 
        U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, 
        U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, 
        U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, 
        U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, 
        U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, 
        U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, 
        U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, 
        U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, 
        U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, 
        U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, 
        U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, 
        U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, 
        U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, 
        U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, 
        U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, 
        U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, 
        U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, 
        U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, 
        U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, 
        U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, 
        U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, 
        U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, 
        U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, 
        U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, 
        U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, 
        U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, 
        U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780;

  INV_X1 U3429 ( .A(n5945), .ZN(n5963) );
  INV_X1 U3430 ( .A(n6159), .ZN(n6134) );
  BUF_X2 U3431 ( .A(n3555), .Z(n2990) );
  XNOR2_X1 U3432 ( .A(n3271), .B(n3270), .ZN(n3359) );
  CLKBUF_X2 U3433 ( .A(n3213), .Z(n4176) );
  CLKBUF_X2 U3434 ( .A(n3176), .Z(n4178) );
  CLKBUF_X2 U3435 ( .A(n3205), .Z(n4167) );
  CLKBUF_X2 U3436 ( .A(n3182), .Z(n4170) );
  CLKBUF_X2 U3437 ( .A(n3254), .Z(n3195) );
  CLKBUF_X2 U3438 ( .A(n3203), .Z(n4133) );
  CLKBUF_X2 U3439 ( .A(n3223), .Z(n2983) );
  CLKBUF_X2 U3440 ( .A(n3194), .Z(n4169) );
  CLKBUF_X2 U3441 ( .A(n3212), .Z(n4177) );
  NOR2_X1 U3444 ( .A1(n3636), .A2(n3134), .ZN(n3126) );
  AND4_X1 U34450 ( .A1(n3093), .A2(n3092), .A3(n3091), .A4(n3090), .ZN(n3104)
         );
  AND2_X2 U34460 ( .A1(n4317), .A2(n3011), .ZN(n3254) );
  INV_X1 U34470 ( .A(n3555), .ZN(n4349) );
  AND4_X1 U34480 ( .A1(n3020), .A2(n3019), .A3(n3018), .A4(n3017), .ZN(n3021)
         );
  AND4_X1 U3449 ( .A1(n3101), .A2(n3100), .A3(n3099), .A4(n3098), .ZN(n3102)
         );
  CLKBUF_X2 U3450 ( .A(n3119), .Z(n3540) );
  AND2_X1 U34510 ( .A1(n3123), .A2(n3147), .ZN(n3526) );
  OR2_X1 U34520 ( .A1(n3083), .A2(n3082), .ZN(n3133) );
  AND2_X1 U34530 ( .A1(n5482), .A2(n5483), .ZN(n5480) );
  OAI21_X1 U3454 ( .B1(n5229), .B2(n5210), .A(n5209), .ZN(n5211) );
  INV_X1 U34550 ( .A(n3636), .ZN(n4497) );
  AND2_X1 U34560 ( .A1(n5022), .A2(n5059), .ZN(n5107) );
  XNOR2_X1 U3457 ( .A(n5239), .B(n5238), .ZN(n5352) );
  XNOR2_X1 U3458 ( .A(n3372), .B(n3335), .ZN(n4395) );
  NAND2_X1 U34590 ( .A1(n5834), .A2(n4900), .ZN(n5916) );
  AND2_X1 U34600 ( .A1(n3360), .A2(n3359), .ZN(n2981) );
  CLKBUF_X3 U34610 ( .A(n5385), .Z(n2989) );
  AND2_X1 U34620 ( .A1(n2981), .A2(n3293), .ZN(n2982) );
  NOR2_X2 U34630 ( .A1(n3456), .A2(n5480), .ZN(n5454) );
  AND2_X4 U34640 ( .A1(n3016), .A2(n4327), .ZN(n3221) );
  AOI21_X1 U34650 ( .B1(n5313), .B2(n6128), .A(n5307), .ZN(n5308) );
  OAI21_X1 U3466 ( .B1(n5749), .B2(n4200), .A(n5596), .ZN(n4203) );
  CLKBUF_X1 U3467 ( .A(n3451), .Z(n5752) );
  OAI21_X1 U34680 ( .B1(n4247), .B2(n4215), .A(n5259), .ZN(n5293) );
  NAND2_X1 U34690 ( .A1(n4214), .A2(n4215), .ZN(n5259) );
  NAND2_X1 U34700 ( .A1(n5358), .A2(n2992), .ZN(n5359) );
  NOR2_X1 U34710 ( .A1(n5233), .A2(n3695), .ZN(n3696) );
  AND2_X1 U34720 ( .A1(n5125), .A2(n2996), .ZN(n3445) );
  AND2_X1 U34730 ( .A1(n5153), .A2(n3444), .ZN(n5125) );
  INV_X8 U34740 ( .A(n5596), .ZN(n3447) );
  INV_X1 U3475 ( .A(n3440), .ZN(n5596) );
  NAND2_X1 U3476 ( .A1(n3327), .A2(n3326), .ZN(n3385) );
  NAND2_X2 U3477 ( .A1(n3425), .A2(n3424), .ZN(n3440) );
  NAND2_X1 U3478 ( .A1(n5414), .A2(n3599), .ZN(n5417) );
  NAND2_X1 U3479 ( .A1(n3362), .A2(n3361), .ZN(n3363) );
  CLKBUF_X1 U3480 ( .A(n4467), .Z(n5063) );
  CLKBUF_X1 U3481 ( .A(n4406), .Z(n6218) );
  NAND2_X1 U3482 ( .A1(n3268), .A2(n3267), .ZN(n3271) );
  CLKBUF_X1 U3483 ( .A(n5984), .Z(n5719) );
  NAND2_X1 U3484 ( .A1(n3157), .A2(n3244), .ZN(n3246) );
  OR2_X1 U3485 ( .A1(n3641), .A2(n3175), .ZN(n3191) );
  NAND2_X1 U3486 ( .A1(n3526), .A2(n4475), .ZN(n4289) );
  CLKBUF_X1 U3487 ( .A(n3531), .Z(n4313) );
  AND2_X1 U3488 ( .A1(n3140), .A2(n3139), .ZN(n3525) );
  CLKBUF_X1 U3489 ( .A(n3565), .Z(n4223) );
  NAND2_X1 U3490 ( .A1(n4349), .A2(n2989), .ZN(n3673) );
  INV_X1 U3491 ( .A(n5287), .ZN(n3635) );
  INV_X1 U3492 ( .A(n3145), .ZN(n3121) );
  CLKBUF_X2 U3493 ( .A(n3142), .Z(n3164) );
  INV_X1 U3494 ( .A(n3134), .ZN(n5289) );
  OR2_X1 U3495 ( .A1(n3211), .A2(n3210), .ZN(n3426) );
  CLKBUF_X2 U3496 ( .A(n3118), .Z(n3698) );
  CLKBUF_X2 U3497 ( .A(n3134), .Z(n3510) );
  INV_X1 U3498 ( .A(n3545), .ZN(n3135) );
  NAND2_X1 U3499 ( .A1(n3006), .A2(n3021), .ZN(n3118) );
  NAND4_X1 U3500 ( .A1(n3062), .A2(n3061), .A3(n3060), .A4(n3059), .ZN(n3119)
         );
  OR2_X2 U3501 ( .A1(n3117), .A2(n3116), .ZN(n3545) );
  AND4_X1 U3502 ( .A1(n3046), .A2(n3045), .A3(n3044), .A4(n3043), .ZN(n3062)
         );
  AND4_X1 U3503 ( .A1(n3058), .A2(n3057), .A3(n3056), .A4(n3055), .ZN(n3059)
         );
  AND4_X1 U3504 ( .A1(n3050), .A2(n3049), .A3(n3048), .A4(n3047), .ZN(n3061)
         );
  AND4_X1 U3505 ( .A1(n3089), .A2(n3088), .A3(n3087), .A4(n3086), .ZN(n3105)
         );
  BUF_X2 U3506 ( .A(n3220), .Z(n4168) );
  NAND2_X2 U3507 ( .A1(n4216), .A2(n6310), .ZN(n6142) );
  BUF_X2 U3508 ( .A(n3196), .Z(n4175) );
  AND2_X2 U3509 ( .A1(n6476), .A2(n4434), .ZN(n6031) );
  OR2_X2 U3510 ( .A1(n3624), .A2(n3625), .ZN(n5565) );
  INV_X1 U3511 ( .A(n5208), .ZN(n2984) );
  NAND2_X1 U3512 ( .A1(n2981), .A2(n3293), .ZN(n2985) );
  NAND2_X1 U3513 ( .A1(n3360), .A2(n3359), .ZN(n2986) );
  NAND2_X1 U3514 ( .A1(n5450), .A2(n5451), .ZN(n2987) );
  CLKBUF_X1 U3515 ( .A(n4882), .Z(n2988) );
  INV_X1 U3516 ( .A(n5208), .ZN(n5442) );
  NAND2_X1 U3517 ( .A1(n2981), .A2(n3293), .ZN(n3376) );
  NAND2_X1 U3518 ( .A1(n5450), .A2(n5451), .ZN(n5449) );
  OAI22_X2 U3519 ( .A1(n4225), .A2(n5396), .B1(n4227), .B2(n4224), .ZN(n5232)
         );
  XNOR2_X2 U3521 ( .A(n4222), .B(n5210), .ZN(n5265) );
  OR2_X2 U3522 ( .A1(n5442), .A2(n4221), .ZN(n2991) );
  NOR2_X2 U3524 ( .A1(n4453), .A2(n4452), .ZN(n4567) );
  NAND2_X1 U3525 ( .A1(n3545), .A2(n3133), .ZN(n5385) );
  NAND2_X1 U3526 ( .A1(n3545), .A2(n3138), .ZN(n3555) );
  NOR2_X1 U3528 ( .A1(n5359), .A2(n4246), .ZN(n4214) );
  AND2_X1 U3529 ( .A1(n5343), .A2(n5365), .ZN(n5358) );
  XNOR2_X1 U3530 ( .A(n3425), .B(n3412), .ZN(n3757) );
  NAND2_X1 U3531 ( .A1(n6466), .A2(n6723), .ZN(n4164) );
  OR2_X1 U3532 ( .A1(n3280), .A2(n6476), .ZN(n3485) );
  NAND2_X1 U3534 ( .A1(n3536), .A2(n3535), .ZN(n3647) );
  AND3_X1 U3535 ( .A1(n4305), .A2(n4304), .A3(n4303), .ZN(n6435) );
  AND2_X1 U3536 ( .A1(n6011), .A2(n5290), .ZN(n6004) );
  INV_X1 U3537 ( .A(n6011), .ZN(n6003) );
  NAND2_X1 U3538 ( .A1(n3146), .A2(n3636), .ZN(n3148) );
  NAND2_X1 U3539 ( .A1(n3318), .A2(n3317), .ZN(n3403) );
  INV_X1 U3540 ( .A(n3319), .ZN(n3317) );
  NAND2_X1 U3541 ( .A1(n5834), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4954) );
  AND2_X1 U3542 ( .A1(n4045), .A2(n5253), .ZN(n5254) );
  OR2_X1 U3543 ( .A1(n5267), .A2(n6476), .ZN(n4161) );
  INV_X1 U3544 ( .A(n4800), .ZN(n3747) );
  AND2_X1 U3545 ( .A1(n4347), .A2(n4348), .ZN(n3720) );
  OR2_X1 U3546 ( .A1(n5524), .A2(n3441), .ZN(n5513) );
  OAI21_X2 U3547 ( .B1(n3246), .B2(n3245), .A(n3244), .ZN(n3272) );
  CLKBUF_X1 U3548 ( .A(n3724), .Z(n4608) );
  NAND2_X1 U3549 ( .A1(n4406), .A2(n6476), .ZN(n3292) );
  OAI21_X1 U3550 ( .B1(n6582), .B2(n4434), .A(n6565), .ZN(n4473) );
  AND2_X1 U3551 ( .A1(n3280), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3507) );
  NOR2_X1 U3552 ( .A1(n3485), .A2(n3484), .ZN(n3504) );
  INV_X1 U3553 ( .A(n5863), .ZN(n5924) );
  NOR2_X2 U3554 ( .A1(n5417), .A2(n5130), .ZN(n5407) );
  AND2_X1 U3555 ( .A1(n3572), .A2(n3002), .ZN(n4566) );
  OR2_X1 U3556 ( .A1(n4144), .A2(n4213), .ZN(n4145) );
  OR2_X1 U3557 ( .A1(n4145), .A2(n5335), .ZN(n4898) );
  NOR2_X2 U3558 ( .A1(n5259), .A2(n5260), .ZN(n5298) );
  AND2_X1 U3559 ( .A1(n5411), .A2(n5410), .ZN(n5760) );
  OR2_X1 U3560 ( .A1(n5434), .A2(n5435), .ZN(n5432) );
  AOI21_X1 U3561 ( .B1(n3757), .B2(n4020), .A(n3756), .ZN(n4924) );
  INV_X1 U3562 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3749) );
  AND2_X1 U3563 ( .A1(n4322), .A2(n6473), .ZN(n6035) );
  NAND2_X1 U3564 ( .A1(n3447), .A2(n5548), .ZN(n4204) );
  AND2_X1 U3565 ( .A1(n3598), .A2(n3597), .ZN(n5415) );
  NOR2_X2 U3566 ( .A1(n4891), .A2(n4890), .ZN(n4936) );
  NAND2_X1 U3567 ( .A1(n6476), .A2(n4473), .ZN(n4974) );
  AND2_X1 U3568 ( .A1(n4432), .A2(n4431), .ZN(n6458) );
  AND2_X1 U3569 ( .A1(n5834), .A2(n4901), .ZN(n5945) );
  AND2_X2 U3570 ( .A1(n3701), .A2(n6473), .ZN(n5988) );
  NAND2_X1 U3571 ( .A1(n5988), .A2(n5310), .ZN(n5983) );
  NAND2_X1 U3572 ( .A1(n6118), .A2(n4375), .ZN(n6011) );
  OR2_X1 U3573 ( .A1(n4248), .A2(n4247), .ZN(n5728) );
  INV_X1 U3574 ( .A(n6135), .ZN(n6129) );
  NAND2_X1 U3575 ( .A1(n6035), .A2(n6453), .ZN(n6135) );
  INV_X1 U3576 ( .A(n5769), .ZN(n6139) );
  NOR2_X1 U3577 ( .A1(n3697), .A2(n3696), .ZN(n5333) );
  INV_X1 U3578 ( .A(n3694), .ZN(n3695) );
  OR2_X1 U3579 ( .A1(n5206), .A2(n4232), .ZN(n5241) );
  AND2_X1 U3580 ( .A1(n3647), .A2(n3629), .ZN(n6161) );
  AND2_X2 U3581 ( .A1(n3717), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3011)
         );
  NAND2_X1 U3582 ( .A1(n2993), .A2(n3005), .ZN(n3167) );
  AOI22_X1 U3583 ( .A1(n3196), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3014) );
  NAND2_X1 U3584 ( .A1(n3134), .A2(n3702), .ZN(n3142) );
  CLKBUF_X1 U3585 ( .A(n3222), .Z(n3202) );
  AND2_X1 U3586 ( .A1(n3316), .A2(n3315), .ZN(n3319) );
  OR2_X1 U3587 ( .A1(n3397), .A2(n3396), .ZN(n3414) );
  OR2_X1 U3588 ( .A1(n3303), .A2(n3302), .ZN(n3377) );
  OR2_X1 U3589 ( .A1(n3265), .A2(n3264), .ZN(n3322) );
  AOI22_X1 U3590 ( .A1(n3127), .A2(n5289), .B1(n5288), .B2(n3636), .ZN(n3122)
         );
  AND2_X1 U3591 ( .A1(n3126), .A2(n3133), .ZN(n3084) );
  INV_X1 U3592 ( .A(n3485), .ZN(n3478) );
  AND2_X2 U3593 ( .A1(n4327), .A2(n4409), .ZN(n3212) );
  NAND2_X1 U3594 ( .A1(n4037), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4010)
         );
  OR2_X1 U3595 ( .A1(n3236), .A2(n6476), .ZN(n3423) );
  INV_X1 U3596 ( .A(n3402), .ZN(n3400) );
  INV_X1 U3597 ( .A(n3565), .ZN(n3670) );
  INV_X1 U3598 ( .A(n3191), .ZN(n3192) );
  NAND2_X1 U3599 ( .A1(n3708), .A2(n6476), .ZN(n3346) );
  NAND2_X1 U3600 ( .A1(n3274), .A2(n3273), .ZN(n4307) );
  AND2_X1 U3601 ( .A1(n3130), .A2(n3250), .ZN(n4843) );
  INV_X1 U3602 ( .A(n3529), .ZN(n3276) );
  NOR2_X1 U3603 ( .A1(n4608), .A2(n6179), .ZN(n5064) );
  AND2_X1 U3604 ( .A1(n6218), .A2(n6314), .ZN(n4812) );
  INV_X1 U3605 ( .A(n3760), .ZN(n3775) );
  NAND2_X1 U3606 ( .A1(n5567), .A2(n5345), .ZN(n5370) );
  AND2_X1 U3607 ( .A1(n4084), .A2(n4083), .ZN(n5365) );
  AND2_X1 U3608 ( .A1(n6035), .A2(n4265), .ZN(n6013) );
  AND2_X1 U3609 ( .A1(n6035), .A2(n4278), .ZN(n6036) );
  INV_X1 U3610 ( .A(n3842), .ZN(n5299) );
  AND2_X1 U3611 ( .A1(n5326), .A2(n4191), .ZN(n4192) );
  OR2_X1 U3612 ( .A1(n5648), .A2(n4164), .ZN(n4125) );
  BUF_X1 U3613 ( .A(n5358), .Z(n5364) );
  NOR2_X1 U3614 ( .A1(n4081), .A2(n5447), .ZN(n4120) );
  CLKBUF_X1 U3615 ( .A(n5343), .Z(n5366) );
  NOR2_X1 U3616 ( .A1(n3922), .A2(n5249), .ZN(n3887) );
  AND2_X1 U3617 ( .A1(n4046), .A2(n5254), .ZN(n4047) );
  AND2_X1 U3618 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n3886), .ZN(n3923)
         );
  NAND2_X1 U3619 ( .A1(n3923), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3922)
         );
  NOR2_X1 U3620 ( .A1(n3992), .A2(n5499), .ZN(n3957) );
  AND2_X1 U3621 ( .A1(n3996), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3993)
         );
  NOR2_X1 U3622 ( .A1(n4010), .A2(n4011), .ZN(n3996) );
  NOR2_X1 U3624 ( .A1(n3822), .A2(n5119), .ZN(n3841) );
  INV_X1 U3625 ( .A(n3857), .ZN(n5167) );
  NAND2_X1 U3626 ( .A1(n3806), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3822)
         );
  NOR2_X1 U3627 ( .A1(n3791), .A2(n5034), .ZN(n3806) );
  NAND2_X1 U3628 ( .A1(n3775), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3791)
         );
  INV_X1 U3630 ( .A(n4924), .ZN(n3758) );
  AOI21_X1 U3631 ( .B1(n3746), .B2(n4020), .A(n3745), .ZN(n4800) );
  CLKBUF_X1 U3632 ( .A(n4797), .Z(n4923) );
  NAND2_X1 U3633 ( .A1(n3739), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3750)
         );
  NOR2_X1 U3634 ( .A1(n3734), .A2(n5943), .ZN(n3739) );
  NAND2_X1 U3635 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3725) );
  NAND2_X1 U3636 ( .A1(n3716), .A2(n4346), .ZN(n4445) );
  AND2_X1 U3637 ( .A1(n3539), .A2(n3538), .ZN(n6453) );
  OR2_X1 U3638 ( .A1(n4354), .A2(n3714), .ZN(n4355) );
  INV_X1 U3639 ( .A(n5233), .ZN(n5234) );
  INV_X1 U3640 ( .A(n4225), .ZN(n3692) );
  INV_X1 U3641 ( .A(n5470), .ZN(n5456) );
  CLKBUF_X1 U3642 ( .A(n5492), .Z(n5493) );
  AND2_X1 U3643 ( .A1(n5151), .A2(n2998), .ZN(n3438) );
  OR2_X1 U3644 ( .A1(n3440), .A2(n5613), .ZN(n5127) );
  INV_X1 U3645 ( .A(n5415), .ZN(n3599) );
  OR2_X1 U3646 ( .A1(n5525), .A2(n5513), .ZN(n5529) );
  AND2_X1 U3647 ( .A1(n3590), .A2(n3589), .ZN(n5112) );
  CLKBUF_X1 U3648 ( .A(n5141), .Z(n5152) );
  INV_X1 U3649 ( .A(n4738), .ZN(n3576) );
  INV_X1 U3650 ( .A(n4739), .ZN(n3577) );
  AND2_X1 U3651 ( .A1(n3571), .A2(n3570), .ZN(n4452) );
  NAND2_X1 U3652 ( .A1(n3564), .A2(n3563), .ZN(n4453) );
  INV_X1 U3653 ( .A(n4400), .ZN(n3563) );
  INV_X1 U3654 ( .A(n4443), .ZN(n3564) );
  NAND2_X1 U3655 ( .A1(n3561), .A2(n3560), .ZN(n4443) );
  INV_X1 U3656 ( .A(n4441), .ZN(n3561) );
  INV_X1 U3657 ( .A(n4440), .ZN(n3560) );
  AND2_X1 U3658 ( .A1(n3647), .A2(n5266), .ZN(n5625) );
  NAND2_X1 U3659 ( .A1(n3683), .A2(n2989), .ZN(n5236) );
  NOR2_X1 U3660 ( .A1(n4268), .A2(n4475), .ZN(n3125) );
  NAND2_X1 U3662 ( .A1(n3233), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3350) );
  INV_X1 U3663 ( .A(n3232), .ZN(n3233) );
  XNOR2_X1 U3664 ( .A(n3272), .B(n3273), .ZN(n4328) );
  NAND2_X1 U3665 ( .A1(n3376), .A2(n3329), .ZN(n3724) );
  XNOR2_X1 U3666 ( .A(n4307), .B(n6375), .ZN(n4406) );
  INV_X1 U3668 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4332) );
  OR2_X1 U3669 ( .A1(n3521), .A2(n3636), .ZN(n5267) );
  AND2_X2 U3670 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4409) );
  CLKBUF_X1 U3671 ( .A(n4289), .Z(n4290) );
  INV_X1 U3672 ( .A(n4974), .ZN(n4763) );
  AND2_X1 U3673 ( .A1(n5064), .A2(n4965), .ZN(n4817) );
  AND2_X1 U3674 ( .A1(n5067), .A2(n6218), .ZN(n6315) );
  OR2_X1 U3675 ( .A1(n4707), .A2(n5065), .ZN(n6372) );
  INV_X1 U3676 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6446) );
  NAND2_X1 U3677 ( .A1(n4474), .A2(n4473), .ZN(n4507) );
  AND2_X1 U3678 ( .A1(n3509), .A2(n3508), .ZN(n4322) );
  INV_X2 U3679 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U3680 ( .A1(n4279), .A2(n5639), .ZN(n6578) );
  INV_X1 U3681 ( .A(n6036), .ZN(n4279) );
  INV_X1 U3682 ( .A(n5916), .ZN(n5881) );
  INV_X1 U3683 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5119) );
  NAND2_X1 U3684 ( .A1(n4951), .A2(n4903), .ZN(n5863) );
  NAND2_X1 U3685 ( .A1(n4913), .A2(n4912), .ZN(n5969) );
  NOR2_X1 U3686 ( .A1(n6013), .A2(n6031), .ZN(n6024) );
  BUF_X1 U3687 ( .A(n6024), .Z(n6030) );
  CLKBUF_X1 U3688 ( .A(n6059), .Z(n6098) );
  NAND2_X1 U3689 ( .A1(n6036), .A2(n4370), .ZN(n6118) );
  NOR2_X1 U3690 ( .A1(n4898), .A2(n5222), .ZN(n4899) );
  INV_X1 U3691 ( .A(n5732), .ZN(n5661) );
  AND2_X1 U3692 ( .A1(n5762), .A2(n5761), .ZN(n5996) );
  OR2_X1 U3693 ( .A1(n5760), .A2(n5759), .ZN(n5761) );
  AND2_X1 U3694 ( .A1(n5432), .A2(n5409), .ZN(n5412) );
  INV_X1 U3696 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5943) );
  AND2_X1 U3697 ( .A1(n2984), .A2(n4205), .ZN(n4207) );
  INV_X1 U3698 ( .A(n5162), .ZN(n6162) );
  INV_X1 U3699 ( .A(n5636), .ZN(n6166) );
  NOR2_X1 U3700 ( .A1(n4884), .A2(n4365), .ZN(n6169) );
  INV_X1 U3701 ( .A(n6161), .ZN(n5631) );
  INV_X1 U3702 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6369) );
  INV_X1 U3703 ( .A(n6310), .ZN(n6374) );
  CLKBUF_X1 U3704 ( .A(n4311), .Z(n4312) );
  CLKBUF_X1 U3705 ( .A(n4328), .Z(n4329) );
  INV_X1 U3706 ( .A(n4607), .ZN(n6179) );
  OAI21_X1 U3707 ( .B1(n4433), .B2(n6559), .A(n4974), .ZN(n6174) );
  INV_X1 U3708 ( .A(n6469), .ZN(n6565) );
  INV_X1 U3709 ( .A(n6191), .ZN(n6386) );
  INV_X1 U3710 ( .A(n6194), .ZN(n6392) );
  INV_X1 U3711 ( .A(n6200), .ZN(n6404) );
  INV_X1 U3712 ( .A(n6203), .ZN(n6410) );
  AND2_X1 U3713 ( .A1(n4477), .A2(n6304), .ZN(n4792) );
  INV_X1 U3714 ( .A(n4645), .ZN(n4511) );
  INV_X1 U3715 ( .A(n6213), .ZN(n6424) );
  INV_X1 U3716 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6476) );
  AND2_X1 U3717 ( .A1(n4322), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6469) );
  INV_X1 U3718 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U3719 ( .A1(n5325), .A2(n4196), .ZN(n4198) );
  INV_X1 U3720 ( .A(n5325), .ZN(n5296) );
  INV_X1 U3721 ( .A(n4251), .ZN(n4252) );
  OAI21_X1 U3722 ( .B1(n5728), .B2(n6142), .A(n4250), .ZN(n4251) );
  OR2_X1 U3723 ( .A1(n5245), .A2(n5244), .ZN(n5246) );
  INV_X1 U3724 ( .A(n5300), .ZN(n3824) );
  NOR2_X4 U3725 ( .A1(n5288), .A2(n6466), .ZN(n5300) );
  AND2_X1 U3726 ( .A1(n5048), .A2(n5112), .ZN(n5113) );
  INV_X1 U3727 ( .A(n6541), .ZN(n6778) );
  INV_X1 U3728 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6500) );
  AND2_X1 U3729 ( .A1(n4102), .A2(n4101), .ZN(n2992) );
  AND2_X1 U3730 ( .A1(n3141), .A2(n5288), .ZN(n2993) );
  AND2_X1 U3731 ( .A1(n3338), .A2(n3337), .ZN(n2994) );
  INV_X1 U3732 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4411) );
  NOR2_X2 U3733 ( .A1(n4707), .A2(n6304), .ZN(n2995) );
  NAND2_X1 U3734 ( .A1(n3447), .A2(n5613), .ZN(n2996) );
  NOR2_X1 U3735 ( .A1(n3447), .A2(n5515), .ZN(n2997) );
  NOR2_X1 U3736 ( .A1(n5513), .A2(n2997), .ZN(n2998) );
  OR2_X2 U3737 ( .A1(n5370), .A2(n5369), .ZN(n2999) );
  OR2_X1 U3738 ( .A1(n5236), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3000)
         );
  OR2_X1 U3739 ( .A1(n5236), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3001)
         );
  OR2_X1 U3740 ( .A1(n5236), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3002)
         );
  INV_X1 U3741 ( .A(n3169), .ZN(n3170) );
  NAND2_X1 U3742 ( .A1(n3447), .A2(n3650), .ZN(n3003) );
  NAND2_X1 U3743 ( .A1(n3440), .A2(n5052), .ZN(n3004) );
  OR2_X1 U3744 ( .A1(n3142), .A2(n3540), .ZN(n3005) );
  AND2_X1 U3745 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3007) );
  INV_X1 U3746 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3717) );
  OR2_X1 U3747 ( .A1(n3350), .A2(n3349), .ZN(n3008) );
  AND3_X1 U3748 ( .A1(n5450), .A2(n5596), .A3(n5539), .ZN(n3009) );
  INV_X1 U3749 ( .A(n4600), .ZN(n3293) );
  AND2_X1 U3750 ( .A1(n3634), .A2(n3144), .ZN(n3150) );
  AOI21_X1 U3751 ( .B1(n4278), .B2(n3512), .A(n3541), .ZN(n3128) );
  OAI21_X1 U3752 ( .B1(n5385), .B2(n3137), .A(n3136), .ZN(n3163) );
  AND2_X1 U3754 ( .A1(n3537), .A2(n3473), .ZN(n3497) );
  AOI22_X1 U3755 ( .A1(n3218), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3012) );
  OR2_X1 U3756 ( .A1(n3482), .A2(n3480), .ZN(n3463) );
  OR2_X1 U3757 ( .A1(n3314), .A2(n3313), .ZN(n3324) );
  OR2_X1 U3758 ( .A1(n3188), .A2(n3187), .ZN(n3341) );
  OR2_X1 U3759 ( .A1(n3472), .A2(n3471), .ZN(n3513) );
  OR2_X1 U3760 ( .A1(n3230), .A2(n3229), .ZN(n3353) );
  AND2_X1 U3761 ( .A1(n3469), .A2(n3470), .ZN(n3467) );
  INV_X1 U3762 ( .A(n3403), .ZN(n3401) );
  NAND2_X1 U3763 ( .A1(n3121), .A2(n3540), .ZN(n3169) );
  NAND2_X1 U3764 ( .A1(n3106), .A2(n3540), .ZN(n3280) );
  OR2_X1 U3765 ( .A1(n3290), .A2(n3289), .ZN(n3332) );
  AOI22_X1 U3766 ( .A1(n3203), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3028) );
  AOI21_X1 U3767 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6446), .A(n3467), 
        .ZN(n3503) );
  NOR2_X1 U3768 ( .A1(n3555), .A2(n5385), .ZN(n3565) );
  AND2_X2 U3769 ( .A1(n3011), .A2(n4316), .ZN(n3218) );
  NAND2_X1 U3770 ( .A1(n5167), .A2(n3858), .ZN(n3859) );
  INV_X1 U3771 ( .A(n5168), .ZN(n3839) );
  NOR2_X1 U3772 ( .A1(n3750), .A2(n3749), .ZN(n3751) );
  AND2_X1 U3773 ( .A1(n3399), .A2(n3398), .ZN(n3402) );
  INV_X1 U3774 ( .A(n3721), .ZN(n3716) );
  NAND2_X1 U3775 ( .A1(n3401), .A2(n3400), .ZN(n3425) );
  MUX2_X1 U3776 ( .A(n3670), .B(n3683), .S(EBX_REG_2__SCAN_IN), .Z(n3559) );
  OR2_X1 U3777 ( .A1(n6304), .A2(n3484), .ZN(n3356) );
  AND4_X1 U3778 ( .A1(n3168), .A2(n3120), .A3(n3141), .A4(n3145), .ZN(n3123)
         );
  NAND2_X1 U3779 ( .A1(n3253), .A2(n3252), .ZN(n3273) );
  INV_X1 U3780 ( .A(n3348), .ZN(n3349) );
  AND4_X1 U3781 ( .A1(n3054), .A2(n3053), .A3(n3052), .A4(n3051), .ZN(n3060)
         );
  NAND2_X1 U3782 ( .A1(n3135), .A2(n4506), .ZN(n3537) );
  AOI22_X1 U3783 ( .A1(n3254), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3196), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3033) );
  AND2_X1 U3784 ( .A1(n3698), .A2(n5288), .ZN(n3127) );
  AND4_X1 U3785 ( .A1(n3097), .A2(n3096), .A3(n3095), .A4(n3094), .ZN(n3103)
         );
  OR2_X1 U3786 ( .A1(n4080), .A2(n5462), .ZN(n4081) );
  NOR2_X1 U3787 ( .A1(n3885), .A2(n5865), .ZN(n4037) );
  NAND2_X1 U3788 ( .A1(n3841), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3885)
         );
  NAND2_X1 U3789 ( .A1(n3751), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3760)
         );
  INV_X1 U3790 ( .A(n3725), .ZN(n3726) );
  INV_X1 U3791 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5210) );
  AND2_X1 U3792 ( .A1(n3559), .A2(n3558), .ZN(n4440) );
  XNOR2_X1 U3793 ( .A(n3246), .B(n3245), .ZN(n4311) );
  AND2_X2 U3794 ( .A1(n3709), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4316)
         );
  XNOR2_X1 U3795 ( .A(n3193), .B(n3192), .ZN(n3708) );
  AND2_X1 U3796 ( .A1(n3292), .A2(n3291), .ZN(n4600) );
  NAND2_X1 U3797 ( .A1(n3279), .A2(n3278), .ZN(n6375) );
  INV_X1 U3798 ( .A(n4271), .ZN(n4266) );
  OR2_X1 U3799 ( .A1(n5643), .A2(n5314), .ZN(n5338) );
  AND2_X1 U3800 ( .A1(n4120), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4121)
         );
  INV_X1 U3801 ( .A(n3956), .ZN(n3886) );
  INV_X1 U3802 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5865) );
  INV_X1 U3803 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5034) );
  AND2_X1 U3804 ( .A1(n5306), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4901) );
  INV_X1 U3805 ( .A(n4954), .ZN(n4951) );
  NAND2_X1 U3806 ( .A1(n5184), .A2(n4226), .ZN(n4225) );
  NAND2_X1 U3807 ( .A1(n5407), .A2(n5406), .ZN(n5405) );
  AND2_X1 U3808 ( .A1(n3575), .A2(n3574), .ZN(n4738) );
  INV_X1 U3809 ( .A(n4164), .ZN(n4191) );
  XNOR2_X1 U3810 ( .A(n4899), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5306)
         );
  INV_X1 U3811 ( .A(n5297), .ZN(n4195) );
  AND2_X1 U3812 ( .A1(n5377), .A2(n5376), .ZN(n5253) );
  INV_X1 U3813 ( .A(n4041), .ZN(n4020) );
  AND2_X1 U3814 ( .A1(n5025), .A2(n5024), .ZN(n5022) );
  NAND2_X1 U3815 ( .A1(n3726), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3734)
         );
  INV_X1 U3816 ( .A(n5237), .ZN(n5238) );
  NAND2_X1 U3817 ( .A1(n2984), .A2(n4220), .ZN(n5229) );
  NAND2_X1 U3818 ( .A1(n5456), .A2(n5569), .ZN(n5457) );
  AND2_X1 U3819 ( .A1(n4258), .A2(n5624), .ZN(n4884) );
  OAI21_X1 U3820 ( .B1(n3340), .B2(n3337), .A(n3339), .ZN(n4467) );
  AND2_X1 U3821 ( .A1(n4516), .A2(n4608), .ZN(n4837) );
  OR2_X1 U3822 ( .A1(n4966), .A2(n4521), .ZN(n4660) );
  NAND2_X1 U3823 ( .A1(n6179), .A2(n4600), .ZN(n4966) );
  INV_X1 U3824 ( .A(n5063), .ZN(n4965) );
  INV_X1 U3825 ( .A(n6218), .ZN(n6367) );
  AND2_X1 U3826 ( .A1(n6477), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3529) );
  NAND2_X1 U3827 ( .A1(n4121), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4144)
         );
  NAND2_X1 U3828 ( .A1(n3887), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4080)
         );
  NAND2_X1 U3829 ( .A1(n3993), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3992)
         );
  AND2_X1 U3830 ( .A1(n5834), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5913) );
  INV_X1 U3831 ( .A(n5941), .ZN(n5921) );
  OR2_X1 U3832 ( .A1(n6578), .A2(n4897), .ZN(n5834) );
  AND2_X1 U3833 ( .A1(n4911), .A2(n4907), .ZN(n5926) );
  INV_X1 U3834 ( .A(n5719), .ZN(n4196) );
  NAND2_X1 U3835 ( .A1(n3577), .A2(n3576), .ZN(n4891) );
  INV_X1 U3836 ( .A(n5983), .ZN(n5977) );
  AND2_X1 U3837 ( .A1(n6011), .A2(n5287), .ZN(n5994) );
  CLKBUF_X1 U3838 ( .A(n4403), .Z(n4447) );
  XNOR2_X1 U3839 ( .A(n5298), .B(n4195), .ZN(n5325) );
  NOR2_X1 U3840 ( .A1(n5712), .A2(n5711), .ZN(n5755) );
  NAND2_X1 U3841 ( .A1(n3957), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3956)
         );
  AND2_X1 U3842 ( .A1(n5434), .A2(n5420), .ZN(n5859) );
  INV_X1 U3843 ( .A(n6133), .ZN(n5763) );
  NAND2_X1 U3844 ( .A1(n3663), .A2(n3662), .ZN(n3664) );
  AND2_X1 U3845 ( .A1(n5611), .A2(n3658), .ZN(n5776) );
  NOR2_X1 U3846 ( .A1(n5137), .A2(n5791), .ZN(n5611) );
  AND2_X1 U3847 ( .A1(n5154), .A2(n5153), .ZN(n5525) );
  NOR2_X1 U3848 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6564) );
  AND2_X1 U3849 ( .A1(n4837), .A2(n6304), .ZN(n6208) );
  AND2_X1 U3850 ( .A1(n4837), .A2(n5065), .ZN(n6209) );
  NOR2_X1 U3851 ( .A1(n4966), .A2(n4965), .ZN(n6215) );
  OR2_X1 U3852 ( .A1(n4976), .A2(n4975), .ZN(n6300) );
  AND2_X1 U3853 ( .A1(n4817), .A2(n6304), .ZN(n6299) );
  INV_X1 U3854 ( .A(n6357), .ZN(n5101) );
  INV_X1 U3855 ( .A(n6304), .ZN(n5065) );
  OR2_X1 U3856 ( .A1(n6380), .A2(n6379), .ZN(n6427) );
  INV_X1 U3857 ( .A(n6372), .ZN(n6425) );
  INV_X1 U3858 ( .A(n6188), .ZN(n6371) );
  INV_X1 U3859 ( .A(n6197), .ZN(n6398) );
  INV_X1 U3860 ( .A(n6206), .ZN(n6416) );
  AND2_X1 U3861 ( .A1(n3529), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6473) );
  AND2_X1 U3862 ( .A1(n6462), .A2(n6461), .ZN(n6467) );
  INV_X1 U3863 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6723) );
  INV_X1 U3864 ( .A(n5913), .ZN(n5959) );
  INV_X1 U3865 ( .A(n5926), .ZN(n5962) );
  INV_X1 U3866 ( .A(n5969), .ZN(n5909) );
  AND2_X1 U3867 ( .A1(n4952), .A2(n5916), .ZN(n5965) );
  OR2_X1 U3868 ( .A1(n5391), .A2(n5390), .ZN(n5743) );
  NAND2_X1 U3869 ( .A1(n5988), .A2(n5288), .ZN(n5984) );
  NAND2_X1 U3870 ( .A1(n6011), .A2(n4377), .ZN(n6010) );
  INV_X1 U3871 ( .A(n6013), .ZN(n6033) );
  AOI211_X1 U3872 ( .C1(n5763), .C2(n5280), .A(n4218), .B(n4217), .ZN(n4219)
         );
  NAND2_X1 U3873 ( .A1(n6135), .A2(n4210), .ZN(n5769) );
  OR2_X1 U3874 ( .A1(n5412), .A2(n5760), .ZN(n6001) );
  NAND2_X1 U3875 ( .A1(n5769), .A2(n6138), .ZN(n6133) );
  OR2_X1 U3876 ( .A1(n5581), .A2(n4233), .ZN(n5574) );
  INV_X1 U3877 ( .A(n6146), .ZN(n5791) );
  NAND2_X1 U3878 ( .A1(n3647), .A2(n3544), .ZN(n5636) );
  INV_X1 U3879 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6439) );
  AOI21_X1 U3880 ( .B1(n4613), .B2(n4671), .A(n4612), .ZN(n4649) );
  NAND2_X1 U3881 ( .A1(n4670), .A2(n5065), .ZN(n4878) );
  AOI21_X1 U3882 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6178), .A(n6177), .ZN(
        n6214) );
  NOR2_X1 U3883 ( .A1(n4520), .A2(n4519), .ZN(n4557) );
  NAND2_X1 U3884 ( .A1(n6215), .A2(n6304), .ZN(n6287) );
  NAND2_X1 U3885 ( .A1(n6215), .A2(n5065), .ZN(n6303) );
  INV_X1 U3886 ( .A(n6300), .ZN(n5001) );
  NAND2_X1 U3887 ( .A1(n4817), .A2(n5065), .ZN(n5099) );
  AOI22_X1 U3888 ( .A1(n5072), .A2(n6315), .B1(n5069), .B2(n5068), .ZN(n5103)
         );
  OR2_X1 U3889 ( .A1(n6305), .A2(n5065), .ZN(n6357) );
  OR2_X1 U3890 ( .A1(n6305), .A2(n6304), .ZN(n6430) );
  AND3_X1 U3891 ( .A1(n4765), .A2(n4764), .A3(n6225), .ZN(n4796) );
  INV_X1 U3892 ( .A(n6558), .ZN(n6489) );
  INV_X1 U3893 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6496) );
  INV_X1 U3894 ( .A(n6551), .ZN(n6549) );
  INV_X1 U3895 ( .A(n6778), .ZN(n6777) );
  OAI211_X1 U3896 ( .C1(n5333), .C2(n5983), .A(n4198), .B(n4197), .ZN(U2829)
         );
  OAI21_X1 U3897 ( .B1(n5265), .B2(n5636), .A(n4241), .ZN(U2989) );
  OR2_X1 U3898 ( .A1(n3667), .A2(n3666), .ZN(U2996) );
  INV_X1 U3899 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3010) );
  AND2_X2 U3900 ( .A1(n3010), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4317)
         );
  NOR2_X4 U3901 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4428) );
  AND2_X2 U3902 ( .A1(n3011), .A2(n4428), .ZN(n3194) );
  AOI22_X1 U3903 ( .A1(n3254), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3015) );
  AND2_X4 U3904 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4327) );
  INV_X1 U3905 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3709) );
  AND2_X4 U3906 ( .A1(n4316), .A2(n4409), .ZN(n3213) );
  AND2_X2 U3907 ( .A1(n4411), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3016)
         );
  AND2_X2 U3908 ( .A1(n4316), .A2(n3016), .ZN(n3220) );
  AOI22_X1 U3909 ( .A1(n3220), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3013) );
  AND2_X2 U3910 ( .A1(n4428), .A2(n4409), .ZN(n3182) );
  NOR2_X4 U3911 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4408) );
  AND2_X2 U3912 ( .A1(n4316), .A2(n4408), .ZN(n3176) );
  AND2_X2 U3913 ( .A1(n4317), .A2(n4408), .ZN(n3222) );
  AOI22_X1 U3914 ( .A1(n3176), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3020) );
  AND2_X2 U3915 ( .A1(n3016), .A2(n4428), .ZN(n3203) );
  AND2_X4 U3916 ( .A1(n4317), .A2(n4409), .ZN(n3204) );
  AOI22_X1 U3917 ( .A1(n3203), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3019) );
  AND2_X2 U3918 ( .A1(n4408), .A2(n4327), .ZN(n3223) );
  AOI22_X1 U3919 ( .A1(n3223), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3018) );
  AND2_X2 U3920 ( .A1(n4317), .A2(n3016), .ZN(n3205) );
  AND2_X4 U3921 ( .A1(n4428), .A2(n4408), .ZN(n4179) );
  AOI22_X1 U3922 ( .A1(n3205), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4179), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3017) );
  AOI22_X1 U3923 ( .A1(n3254), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3025) );
  AOI22_X1 U3924 ( .A1(n3196), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3024) );
  AOI22_X1 U3925 ( .A1(n3220), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3023) );
  AOI22_X1 U3926 ( .A1(n3218), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3022) );
  NAND4_X1 U3927 ( .A1(n3025), .A2(n3024), .A3(n3023), .A4(n3022), .ZN(n3031)
         );
  AOI22_X1 U3928 ( .A1(n3176), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3029) );
  AOI22_X1 U3929 ( .A1(n3223), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3027) );
  AOI22_X1 U3930 ( .A1(n3205), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        INSTQUEUE_REG_0__5__SCAN_IN), .B2(n4179), .ZN(n3026) );
  NAND4_X1 U3931 ( .A1(n3029), .A2(n3028), .A3(n3027), .A4(n3026), .ZN(n3030)
         );
  OR2_X2 U3932 ( .A1(n3031), .A2(n3030), .ZN(n3134) );
  INV_X1 U3933 ( .A(n3134), .ZN(n3032) );
  NAND2_X1 U3934 ( .A1(n3698), .A2(n3032), .ZN(n3141) );
  AOI22_X1 U3935 ( .A1(n3220), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3036) );
  AOI22_X1 U3936 ( .A1(n3205), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3035) );
  AOI22_X1 U3937 ( .A1(n3203), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3034) );
  AND4_X2 U3938 ( .A1(n3036), .A2(n3035), .A3(n3034), .A4(n3033), .ZN(n3042)
         );
  AOI22_X1 U3939 ( .A1(n3176), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3040) );
  AOI22_X1 U3940 ( .A1(n4179), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3223), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3039) );
  AOI22_X1 U3941 ( .A1(n3204), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3038) );
  AOI22_X1 U3942 ( .A1(n3218), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3037) );
  AND4_X2 U3943 ( .A1(n3040), .A2(n3039), .A3(n3038), .A4(n3037), .ZN(n3041)
         );
  NAND2_X4 U3944 ( .A1(n3042), .A2(n3041), .ZN(n5288) );
  NAND2_X1 U3945 ( .A1(n3254), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3046) );
  NAND2_X1 U3946 ( .A1(n3194), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3045) );
  NAND2_X1 U3947 ( .A1(n3213), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3044)
         );
  NAND2_X1 U3948 ( .A1(n3196), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3043)
         );
  NAND2_X1 U3949 ( .A1(n3205), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3050) );
  NAND2_X1 U3950 ( .A1(n3204), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3049)
         );
  NAND2_X1 U3951 ( .A1(n3203), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3048) );
  NAND2_X1 U3952 ( .A1(n4179), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3047) );
  NAND2_X1 U3953 ( .A1(n3218), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3054)
         );
  NAND2_X1 U3954 ( .A1(n3220), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3053) );
  NAND2_X1 U3955 ( .A1(n3221), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3052) );
  NAND2_X1 U3956 ( .A1(n3182), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3051)
         );
  NAND2_X1 U3957 ( .A1(n3176), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3058) );
  NAND2_X1 U3958 ( .A1(n3222), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3057) );
  NAND2_X1 U3959 ( .A1(n3223), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3056) );
  NAND2_X1 U3960 ( .A1(n3212), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3055)
         );
  INV_X2 U3961 ( .A(n3119), .ZN(n4493) );
  AND2_X1 U3962 ( .A1(n5288), .A2(n4493), .ZN(n3063) );
  NAND2_X1 U3963 ( .A1(n3141), .A2(n3063), .ZN(n3139) );
  INV_X1 U3964 ( .A(n3139), .ZN(n3085) );
  AOI22_X1 U3965 ( .A1(n3205), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3203), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3067) );
  AOI22_X1 U3966 ( .A1(n3254), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3066) );
  AOI22_X1 U3967 ( .A1(n3220), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3196), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3065) );
  AOI22_X1 U3968 ( .A1(n3222), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3223), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3064) );
  NAND4_X1 U3969 ( .A1(n3067), .A2(n3066), .A3(n3065), .A4(n3064), .ZN(n3073)
         );
  AOI22_X1 U3970 ( .A1(n3218), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3071) );
  AOI22_X1 U3971 ( .A1(n3204), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4179), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3070) );
  AOI22_X1 U3972 ( .A1(n3213), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3069) );
  AOI22_X1 U3973 ( .A1(n3176), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3068) );
  NAND4_X1 U3974 ( .A1(n3071), .A2(n3070), .A3(n3069), .A4(n3068), .ZN(n3072)
         );
  OR2_X2 U3975 ( .A1(n3073), .A2(n3072), .ZN(n3636) );
  AOI22_X1 U3976 ( .A1(n3254), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3077) );
  AOI22_X1 U3977 ( .A1(n3196), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3076) );
  AOI22_X1 U3978 ( .A1(n3220), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3075) );
  AOI22_X1 U3979 ( .A1(n3218), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3074) );
  NAND4_X1 U3980 ( .A1(n3077), .A2(n3076), .A3(n3075), .A4(n3074), .ZN(n3083)
         );
  AOI22_X1 U3981 ( .A1(n3176), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3081) );
  AOI22_X1 U3982 ( .A1(n3203), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3080) );
  AOI22_X1 U3983 ( .A1(n3223), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3079) );
  AOI22_X1 U3984 ( .A1(n3205), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4179), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3078) );
  NAND4_X1 U3985 ( .A1(n3081), .A2(n3080), .A3(n3079), .A4(n3078), .ZN(n3082)
         );
  NAND2_X1 U3986 ( .A1(n3085), .A2(n3084), .ZN(n3531) );
  INV_X1 U3987 ( .A(n3531), .ZN(n3107) );
  NAND2_X1 U3988 ( .A1(n3196), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3089)
         );
  NAND2_X1 U3989 ( .A1(n3205), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3088) );
  NAND2_X1 U3990 ( .A1(n3221), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3087) );
  NAND2_X1 U3991 ( .A1(n3213), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3086)
         );
  NAND2_X1 U3992 ( .A1(n3254), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3093) );
  NAND2_X1 U3993 ( .A1(n3220), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3092) );
  NAND2_X1 U3994 ( .A1(n3218), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3091)
         );
  NAND2_X1 U3995 ( .A1(n3182), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3090)
         );
  NAND2_X1 U3996 ( .A1(n3203), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3097) );
  NAND2_X1 U3997 ( .A1(n3194), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3096) );
  NAND2_X1 U3998 ( .A1(n3204), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3095)
         );
  NAND2_X1 U3999 ( .A1(n4179), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3094) );
  NAND2_X1 U4000 ( .A1(n3176), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3101) );
  NAND2_X1 U4001 ( .A1(n3222), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3100) );
  NAND2_X1 U4002 ( .A1(n3223), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3099) );
  NAND2_X1 U4003 ( .A1(n3212), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3098)
         );
  NAND4_X4 U4004 ( .A1(n3105), .A2(n3104), .A3(n3103), .A4(n3102), .ZN(n3138)
         );
  INV_X4 U4005 ( .A(n3138), .ZN(n4506) );
  INV_X2 U4006 ( .A(n4506), .ZN(n3106) );
  NAND2_X1 U4007 ( .A1(n3107), .A2(n3106), .ZN(n4268) );
  AOI22_X1 U4008 ( .A1(n3205), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3176), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3111) );
  AOI22_X1 U4009 ( .A1(n3196), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3110) );
  AOI22_X1 U4010 ( .A1(n3221), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3109) );
  AOI22_X1 U4011 ( .A1(n3203), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4179), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3108) );
  NAND4_X1 U4012 ( .A1(n3111), .A2(n3110), .A3(n3109), .A4(n3108), .ZN(n3117)
         );
  AOI22_X1 U4013 ( .A1(n3220), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3115) );
  AOI22_X1 U4014 ( .A1(n3222), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3114) );
  AOI22_X1 U4015 ( .A1(n3194), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3223), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3113) );
  AOI22_X1 U4016 ( .A1(n3254), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3112) );
  NAND4_X1 U4017 ( .A1(n3115), .A2(n3114), .A3(n3113), .A4(n3112), .ZN(n3116)
         );
  INV_X2 U4018 ( .A(n3545), .ZN(n4475) );
  INV_X2 U4019 ( .A(n3118), .ZN(n3702) );
  NAND2_X1 U4020 ( .A1(n3142), .A2(n3133), .ZN(n3168) );
  NOR2_X1 U4021 ( .A1(n3138), .A2(n3540), .ZN(n3120) );
  NAND2_X2 U4022 ( .A1(n3702), .A2(n5288), .ZN(n3145) );
  NAND2_X1 U4023 ( .A1(n3122), .A2(n3169), .ZN(n3147) );
  INV_X1 U4024 ( .A(n4289), .ZN(n3124) );
  NOR2_X2 U4025 ( .A1(n3125), .A2(n3124), .ZN(n3543) );
  INV_X1 U4026 ( .A(n4268), .ZN(n4278) );
  XNOR2_X1 U4027 ( .A(n6496), .B(STATE_REG_2__SCAN_IN), .ZN(n3512) );
  INV_X2 U4028 ( .A(n3133), .ZN(n4501) );
  NAND2_X1 U4029 ( .A1(n3126), .A2(n4501), .ZN(n3699) );
  NOR2_X2 U4031 ( .A1(n4372), .A2(n3635), .ZN(n3541) );
  NAND2_X1 U4032 ( .A1(n3543), .A2(n3128), .ZN(n3129) );
  NAND2_X2 U4033 ( .A1(n3129), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3155) );
  NAND2_X1 U4034 ( .A1(n6564), .A2(n6476), .ZN(n4209) );
  INV_X1 U4035 ( .A(n4209), .ZN(n3277) );
  NAND2_X1 U4036 ( .A1(n6369), .A2(n6439), .ZN(n3130) );
  NAND2_X1 U4037 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3250) );
  AOI22_X1 U4038 ( .A1(n3277), .A2(n4843), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n3276), .ZN(n3153) );
  INV_X1 U4039 ( .A(n3153), .ZN(n3131) );
  NOR2_X1 U4040 ( .A1(n3131), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3132)
         );
  OR2_X2 U4041 ( .A1(n3155), .A2(n3132), .ZN(n3157) );
  AND2_X2 U4042 ( .A1(n4493), .A2(n3510), .ZN(n3538) );
  INV_X1 U4043 ( .A(n3538), .ZN(n3137) );
  AND2_X4 U4044 ( .A1(n3135), .A2(n3138), .ZN(n6037) );
  NAND2_X1 U4045 ( .A1(n3139), .A2(n6037), .ZN(n3136) );
  AND2_X1 U4046 ( .A1(n3164), .A2(n3138), .ZN(n3140) );
  NOR2_X1 U4047 ( .A1(n3163), .A2(n3525), .ZN(n3151) );
  NAND2_X1 U4048 ( .A1(n4497), .A2(n3133), .ZN(n3143) );
  NOR2_X2 U4049 ( .A1(n3167), .A2(n3143), .ZN(n3634) );
  OAI21_X1 U4050 ( .B1(n3512), .B2(n3545), .A(n5289), .ZN(n3144) );
  NAND2_X1 U4051 ( .A1(n3538), .A2(n3145), .ZN(n3146) );
  NAND4_X1 U4052 ( .A1(n3148), .A2(n3147), .A3(n3168), .A4(n4475), .ZN(n3149)
         );
  NAND2_X1 U4053 ( .A1(n3149), .A2(n4506), .ZN(n3162) );
  NAND3_X1 U4054 ( .A1(n3151), .A2(n3150), .A3(n3162), .ZN(n3152) );
  NAND2_X1 U4055 ( .A1(n3152), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3158) );
  INV_X1 U4056 ( .A(n3158), .ZN(n3154) );
  AOI21_X2 U4057 ( .B1(n3154), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3131), 
        .ZN(n3156) );
  NAND2_X2 U4058 ( .A1(n3156), .A2(n3155), .ZN(n3244) );
  INV_X1 U4059 ( .A(n3158), .ZN(n3247) );
  NAND2_X1 U4060 ( .A1(n3247), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3160) );
  MUX2_X1 U4061 ( .A(n3529), .B(n4209), .S(n6369), .Z(n3159) );
  NAND2_X1 U4062 ( .A1(n3160), .A2(n3159), .ZN(n3193) );
  NAND2_X1 U4063 ( .A1(n3510), .A2(n3545), .ZN(n3484) );
  NOR2_X1 U4064 ( .A1(n3484), .A2(n3540), .ZN(n3161) );
  OAI22_X1 U4065 ( .A1(n3162), .A2(n3161), .B1(n4506), .B2(n4497), .ZN(n3641)
         );
  INV_X1 U4066 ( .A(n3163), .ZN(n3174) );
  NAND2_X1 U4067 ( .A1(n3164), .A2(n3540), .ZN(n3165) );
  NAND2_X1 U4068 ( .A1(n3165), .A2(n3133), .ZN(n3166) );
  OAI21_X1 U4069 ( .B1(n3167), .B2(n3166), .A(n3545), .ZN(n3173) );
  NAND2_X1 U4070 ( .A1(n6564), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6480) );
  AOI21_X1 U4071 ( .B1(n3168), .B2(n6037), .A(n6480), .ZN(n3172) );
  NAND2_X1 U4072 ( .A1(n3170), .A2(n4501), .ZN(n3171) );
  NAND4_X1 U4073 ( .A1(n3174), .A2(n3173), .A3(n3172), .A4(n3171), .ZN(n3175)
         );
  AND2_X2 U4074 ( .A1(n3193), .A2(n3191), .ZN(n3245) );
  NAND2_X1 U4075 ( .A1(n4311), .A2(n6476), .ZN(n3190) );
  NOR2_X1 U4076 ( .A1(n3540), .A2(n6476), .ZN(n3266) );
  AOI22_X1 U4077 ( .A1(n4167), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3180) );
  AOI22_X1 U4078 ( .A1(n3224), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4133), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3179) );
  AOI22_X1 U4079 ( .A1(n4175), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3178) );
  AOI22_X1 U4080 ( .A1(n4178), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3177) );
  NAND4_X1 U4081 ( .A1(n3180), .A2(n3179), .A3(n3178), .A4(n3177), .ZN(n3188)
         );
  AOI22_X1 U4082 ( .A1(n4413), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3186) );
  AOI22_X1 U4083 ( .A1(n3219), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3185) );
  INV_X1 U4084 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U4085 ( .A1(n4168), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3184) );
  AOI22_X1 U4086 ( .A1(n4169), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3183) );
  NAND4_X1 U4087 ( .A1(n3186), .A2(n3185), .A3(n3184), .A4(n3183), .ZN(n3187)
         );
  NAND2_X1 U4088 ( .A1(n3266), .A2(n3341), .ZN(n3189) );
  NAND2_X1 U4089 ( .A1(n3190), .A2(n3189), .ZN(n3242) );
  AOI22_X1 U4090 ( .A1(n3195), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3201) );
  AOI22_X1 U4091 ( .A1(n3196), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3200) );
  AOI22_X1 U4092 ( .A1(n3220), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3199) );
  CLKBUF_X1 U4093 ( .A(n3218), .Z(n3197) );
  AOI22_X1 U4094 ( .A1(n3197), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3198) );
  NAND4_X1 U4095 ( .A1(n3201), .A2(n3200), .A3(n3199), .A4(n3198), .ZN(n3211)
         );
  AOI22_X1 U4096 ( .A1(n3176), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3209) );
  AOI22_X1 U4097 ( .A1(n4133), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3208) );
  AOI22_X1 U4098 ( .A1(n2983), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3207) );
  AOI22_X1 U4099 ( .A1(n3205), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3206) );
  NAND4_X1 U4100 ( .A1(n3209), .A2(n3208), .A3(n3207), .A4(n3206), .ZN(n3210)
         );
  NAND2_X1 U4101 ( .A1(n4493), .A2(n3426), .ZN(n3236) );
  INV_X1 U4102 ( .A(n3426), .ZN(n3238) );
  NAND2_X1 U4103 ( .A1(n3238), .A2(n4493), .ZN(n3231) );
  AOI22_X1 U4104 ( .A1(n3205), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4133), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3217) );
  AOI22_X1 U4105 ( .A1(n3195), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3196), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3216) );
  AOI22_X1 U4106 ( .A1(n3176), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3215) );
  AOI22_X1 U4107 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n3213), .B1(n3182), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3214) );
  NAND4_X1 U4108 ( .A1(n3217), .A2(n3216), .A3(n3215), .A4(n3214), .ZN(n3230)
         );
  CLKBUF_X1 U4109 ( .A(n3218), .Z(n3219) );
  AOI22_X1 U4110 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3219), .B1(n4169), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3228) );
  AOI22_X1 U4111 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n3220), .B1(n4413), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3227) );
  BUF_X1 U4112 ( .A(n3222), .Z(n3224) );
  AOI22_X1 U4113 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n3224), .B1(n2983), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3226) );
  AOI22_X1 U4114 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n3259), .B1(n4103), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3225) );
  NAND4_X1 U4115 ( .A1(n3228), .A2(n3227), .A3(n3226), .A4(n3225), .ZN(n3229)
         );
  MUX2_X1 U4116 ( .A(n3236), .B(n3231), .S(n3353), .Z(n3232) );
  NAND2_X1 U4117 ( .A1(n3346), .A2(n3350), .ZN(n3235) );
  INV_X1 U4118 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4621) );
  AOI21_X1 U4119 ( .B1(n4506), .B2(n3353), .A(n6476), .ZN(n3234) );
  OAI211_X1 U4120 ( .C1(n3485), .C2(n4621), .A(n3234), .B(n3236), .ZN(n3348)
         );
  NAND2_X1 U4121 ( .A1(n3235), .A2(n3348), .ZN(n3237) );
  NAND2_X1 U4122 ( .A1(n3237), .A2(n3423), .ZN(n3241) );
  OR2_X2 U4123 ( .A1(n3242), .A2(n3241), .ZN(n3340) );
  NOR2_X1 U4124 ( .A1(n3106), .A2(n6476), .ZN(n3269) );
  NAND2_X1 U4125 ( .A1(n3269), .A2(n3341), .ZN(n3240) );
  NAND2_X1 U4126 ( .A1(n3266), .A2(n3238), .ZN(n3239) );
  OAI211_X1 U4127 ( .C1(n3485), .C2(n3181), .A(n3240), .B(n3239), .ZN(n3336)
         );
  NAND2_X1 U4128 ( .A1(n3340), .A2(n3336), .ZN(n3243) );
  NAND2_X1 U4129 ( .A1(n3242), .A2(n3241), .ZN(n3338) );
  NAND2_X1 U4130 ( .A1(n3243), .A2(n3338), .ZN(n3360) );
  NAND2_X1 U4131 ( .A1(n3247), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3253) );
  INV_X1 U4132 ( .A(n3250), .ZN(n3249) );
  INV_X1 U4133 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3248) );
  NAND2_X1 U4134 ( .A1(n3249), .A2(n3248), .ZN(n6306) );
  NAND2_X1 U4135 ( .A1(n3250), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3251) );
  NAND2_X1 U4136 ( .A1(n6306), .A2(n3251), .ZN(n4522) );
  AOI22_X1 U4137 ( .A1(n3277), .A2(n4522), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3276), .ZN(n3252) );
  NAND2_X1 U4138 ( .A1(n4328), .A2(n6476), .ZN(n3268) );
  AOI22_X1 U4139 ( .A1(n3195), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3258) );
  AOI22_X1 U4140 ( .A1(n4175), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4141 ( .A1(n4168), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3256) );
  AOI22_X1 U4142 ( .A1(n3219), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3255) );
  NAND4_X1 U4143 ( .A1(n3258), .A2(n3257), .A3(n3256), .A4(n3255), .ZN(n3265)
         );
  AOI22_X1 U4144 ( .A1(n4178), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U4145 ( .A1(n4133), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3262) );
  AOI22_X1 U4146 ( .A1(n2983), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3261) );
  AOI22_X1 U4147 ( .A1(n4167), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3260) );
  NAND4_X1 U4148 ( .A1(n3263), .A2(n3262), .A3(n3261), .A4(n3260), .ZN(n3264)
         );
  NAND2_X1 U4149 ( .A1(n3266), .A2(n3322), .ZN(n3267) );
  AOI22_X1 U4150 ( .A1(n3478), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3269), 
        .B2(n3322), .ZN(n3270) );
  INV_X1 U4151 ( .A(n3272), .ZN(n3274) );
  NAND2_X1 U4152 ( .A1(n3154), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3279) );
  NAND3_X1 U4153 ( .A1(n6446), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6263) );
  INV_X1 U4154 ( .A(n6263), .ZN(n6262) );
  NAND2_X1 U4155 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6262), .ZN(n6286) );
  NAND2_X1 U4156 ( .A1(n6446), .A2(n6286), .ZN(n3275) );
  NOR3_X1 U4157 ( .A1(n6446), .A2(n3248), .A3(n6439), .ZN(n4762) );
  NAND2_X1 U4158 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4762), .ZN(n4466) );
  AND2_X1 U4159 ( .A1(n3275), .A2(n4466), .ZN(n4972) );
  AOI22_X1 U4160 ( .A1(n3277), .A2(n4972), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3276), .ZN(n3278) );
  AOI22_X1 U4161 ( .A1(n3195), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4162 ( .A1(n4175), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3283) );
  AOI22_X1 U4163 ( .A1(n4168), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3282) );
  AOI22_X1 U4164 ( .A1(n3219), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3281) );
  NAND4_X1 U4165 ( .A1(n3284), .A2(n3283), .A3(n3282), .A4(n3281), .ZN(n3290)
         );
  AOI22_X1 U4166 ( .A1(n4178), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3288) );
  AOI22_X1 U4167 ( .A1(n4133), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4168 ( .A1(n2983), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4169 ( .A1(n4167), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3285) );
  NAND4_X1 U4170 ( .A1(n3288), .A2(n3287), .A3(n3286), .A4(n3285), .ZN(n3289)
         );
  AOI22_X1 U4171 ( .A1(n3478), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3507), 
        .B2(n3332), .ZN(n3291) );
  INV_X1 U4172 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4641) );
  AOI22_X1 U4173 ( .A1(n3195), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4174 ( .A1(n4175), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4175 ( .A1(n4168), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3295) );
  AOI22_X1 U4176 ( .A1(n3219), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3294) );
  NAND4_X1 U4177 ( .A1(n3297), .A2(n3296), .A3(n3295), .A4(n3294), .ZN(n3303)
         );
  AOI22_X1 U4178 ( .A1(n4178), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4179 ( .A1(n4133), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4180 ( .A1(n2983), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4181 ( .A1(n4167), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3298) );
  NAND4_X1 U4182 ( .A1(n3301), .A2(n3300), .A3(n3299), .A4(n3298), .ZN(n3302)
         );
  NAND2_X1 U4183 ( .A1(n3507), .A2(n3377), .ZN(n3304) );
  OAI21_X1 U4184 ( .B1(n3485), .B2(n4641), .A(n3304), .ZN(n3375) );
  NAND2_X1 U4185 ( .A1(n2982), .A2(n3375), .ZN(n3320) );
  INV_X1 U4186 ( .A(n3320), .ZN(n3318) );
  NAND2_X1 U4187 ( .A1(n3478), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4188 ( .A1(n4178), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4189 ( .A1(n4167), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U4190 ( .A1(n4413), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4191 ( .A1(n2983), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3305) );
  NAND4_X1 U4192 ( .A1(n3308), .A2(n3307), .A3(n3306), .A4(n3305), .ZN(n3314)
         );
  AOI22_X1 U4193 ( .A1(n4168), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U4194 ( .A1(n3195), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4195 ( .A1(n4133), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4196 ( .A1(n4176), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3309) );
  NAND4_X1 U4197 ( .A1(n3312), .A2(n3311), .A3(n3310), .A4(n3309), .ZN(n3313)
         );
  NAND2_X1 U4198 ( .A1(n3507), .A2(n3324), .ZN(n3315) );
  NAND2_X1 U4199 ( .A1(n3320), .A2(n3319), .ZN(n3321) );
  NAND2_X1 U4200 ( .A1(n3403), .A2(n3321), .ZN(n3742) );
  OR2_X1 U4201 ( .A1(n3742), .A2(n3484), .ZN(n3327) );
  NAND2_X1 U4202 ( .A1(n3353), .A2(n3341), .ZN(n3365) );
  INV_X1 U4203 ( .A(n3322), .ZN(n3366) );
  NAND2_X1 U4204 ( .A1(n3365), .A2(n3366), .ZN(n3364) );
  NAND2_X1 U4205 ( .A1(n3364), .A2(n3332), .ZN(n3378) );
  INV_X1 U4206 ( .A(n3377), .ZN(n3323) );
  NOR2_X1 U4207 ( .A1(n3378), .A2(n3323), .ZN(n3325) );
  NAND2_X1 U4208 ( .A1(n3325), .A2(n3324), .ZN(n3413) );
  OAI211_X1 U4209 ( .C1(n3325), .C2(n3324), .A(n3413), .B(n6037), .ZN(n3326)
         );
  INV_X1 U4210 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3328) );
  XNOR2_X1 U4211 ( .A(n3385), .B(n3328), .ZN(n4747) );
  NAND2_X1 U4212 ( .A1(n2986), .A2(n4600), .ZN(n3329) );
  INV_X1 U4213 ( .A(n3724), .ZN(n3331) );
  INV_X1 U4214 ( .A(n3484), .ZN(n3330) );
  NAND2_X1 U4215 ( .A1(n3331), .A2(n3330), .ZN(n3334) );
  OAI211_X1 U4216 ( .C1(n3332), .C2(n3364), .A(n3378), .B(n6037), .ZN(n3333)
         );
  NAND2_X1 U4217 ( .A1(n3334), .A2(n3333), .ZN(n3372) );
  INV_X1 U4218 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3335) );
  INV_X1 U4219 ( .A(n3336), .ZN(n3337) );
  NAND2_X1 U4220 ( .A1(n3340), .A2(n2994), .ZN(n3339) );
  NAND2_X1 U4221 ( .A1(n4467), .A2(n3330), .ZN(n3345) );
  OAI21_X1 U4222 ( .B1(n3341), .B2(n3353), .A(n3365), .ZN(n3342) );
  INV_X1 U4223 ( .A(n6037), .ZN(n6581) );
  OAI211_X1 U4224 ( .C1(n3342), .C2(n6581), .A(n4497), .B(n3510), .ZN(n3343)
         );
  INV_X1 U4225 ( .A(n3343), .ZN(n3344) );
  NAND2_X1 U4226 ( .A1(n3345), .A2(n3344), .ZN(n4359) );
  NAND2_X1 U4227 ( .A1(n3346), .A2(n3348), .ZN(n3347) );
  NAND2_X1 U4228 ( .A1(n3347), .A2(n3350), .ZN(n3351) );
  NAND2_X2 U4229 ( .A1(n3351), .A2(n3008), .ZN(n6304) );
  AND2_X1 U4230 ( .A1(n4506), .A2(n3133), .ZN(n3367) );
  INV_X1 U4231 ( .A(n3367), .ZN(n3352) );
  OAI21_X1 U4232 ( .B1(n6581), .B2(n3353), .A(n3352), .ZN(n3354) );
  INV_X1 U4233 ( .A(n3354), .ZN(n3355) );
  NAND2_X1 U4234 ( .A1(n3356), .A2(n3355), .ZN(n4255) );
  NAND2_X1 U4235 ( .A1(n4255), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4257)
         );
  XNOR2_X1 U4236 ( .A(n4257), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4358)
         );
  NAND2_X1 U4237 ( .A1(n4359), .A2(n4358), .ZN(n4361) );
  INV_X1 U4238 ( .A(n4257), .ZN(n3357) );
  NAND2_X1 U4239 ( .A1(n3357), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3358)
         );
  AND2_X1 U4240 ( .A1(n4361), .A2(n3358), .ZN(n6126) );
  INV_X1 U4241 ( .A(n3359), .ZN(n3362) );
  INV_X1 U4242 ( .A(n3360), .ZN(n3361) );
  NAND2_X2 U4243 ( .A1(n2986), .A2(n3363), .ZN(n4607) );
  OAI21_X1 U4244 ( .B1(n3366), .B2(n3365), .A(n3364), .ZN(n3368) );
  AOI21_X1 U4245 ( .B1(n3368), .B2(n6037), .A(n3367), .ZN(n3369) );
  OAI21_X1 U4246 ( .B1(n4607), .B2(n3484), .A(n3369), .ZN(n3370) );
  NAND2_X1 U4247 ( .A1(n3370), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6123)
         );
  NAND2_X1 U4248 ( .A1(n6126), .A2(n6123), .ZN(n3371) );
  OR2_X1 U4249 ( .A1(n3370), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6124)
         );
  AND2_X1 U4250 ( .A1(n3371), .A2(n6124), .ZN(n4396) );
  NAND2_X1 U4251 ( .A1(n4395), .A2(n4396), .ZN(n3374) );
  NAND2_X1 U4252 ( .A1(n3372), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3373)
         );
  NAND2_X1 U4253 ( .A1(n3374), .A2(n3373), .ZN(n4458) );
  XNOR2_X1 U4254 ( .A(n2985), .B(n3375), .ZN(n3738) );
  NAND2_X1 U4255 ( .A1(n3738), .A2(n3330), .ZN(n3381) );
  XNOR2_X1 U4256 ( .A(n3378), .B(n3377), .ZN(n3379) );
  NAND2_X1 U4257 ( .A1(n3379), .A2(n6037), .ZN(n3380) );
  NAND2_X1 U4258 ( .A1(n3381), .A2(n3380), .ZN(n3382) );
  INV_X1 U4259 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3566) );
  XNOR2_X1 U4260 ( .A(n3382), .B(n3566), .ZN(n4459) );
  NAND2_X1 U4261 ( .A1(n4458), .A2(n4459), .ZN(n3384) );
  NAND2_X1 U4262 ( .A1(n3382), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3383)
         );
  NAND2_X1 U4263 ( .A1(n3384), .A2(n3383), .ZN(n4748) );
  NAND2_X1 U4264 ( .A1(n4747), .A2(n4748), .ZN(n3387) );
  NAND2_X1 U4265 ( .A1(n3385), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3386)
         );
  NAND2_X1 U4266 ( .A1(n3387), .A2(n3386), .ZN(n4735) );
  NAND2_X1 U4267 ( .A1(n3478), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4268 ( .A1(n3195), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3391) );
  AOI22_X1 U4269 ( .A1(n4175), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4270 ( .A1(n4168), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4271 ( .A1(n3197), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3388) );
  NAND4_X1 U4272 ( .A1(n3391), .A2(n3390), .A3(n3389), .A4(n3388), .ZN(n3397)
         );
  AOI22_X1 U4273 ( .A1(n4178), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3395) );
  AOI22_X1 U4274 ( .A1(n4133), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4275 ( .A1(n2983), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4276 ( .A1(n4167), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3392) );
  NAND4_X1 U4277 ( .A1(n3395), .A2(n3394), .A3(n3393), .A4(n3392), .ZN(n3396)
         );
  NAND2_X1 U4278 ( .A1(n3507), .A2(n3414), .ZN(n3398) );
  NAND2_X1 U4279 ( .A1(n3403), .A2(n3402), .ZN(n3746) );
  NAND3_X1 U4280 ( .A1(n3425), .A2(n3330), .A3(n3746), .ZN(n3406) );
  XNOR2_X1 U4281 ( .A(n3413), .B(n3414), .ZN(n3404) );
  NAND2_X1 U4282 ( .A1(n3404), .A2(n6037), .ZN(n3405) );
  NAND2_X1 U4283 ( .A1(n3406), .A2(n3405), .ZN(n3408) );
  INV_X1 U4284 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3407) );
  XNOR2_X1 U4285 ( .A(n3408), .B(n3407), .ZN(n4736) );
  NAND2_X1 U4286 ( .A1(n4735), .A2(n4736), .ZN(n3410) );
  NAND2_X1 U4287 ( .A1(n3408), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3409)
         );
  NAND2_X1 U4288 ( .A1(n3410), .A2(n3409), .ZN(n4882) );
  INV_X1 U4289 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4633) );
  NAND2_X1 U4290 ( .A1(n3507), .A2(n3426), .ZN(n3411) );
  OAI21_X1 U4291 ( .B1(n4633), .B2(n3485), .A(n3411), .ZN(n3412) );
  NAND2_X1 U4292 ( .A1(n3757), .A2(n3330), .ZN(n3418) );
  INV_X1 U4293 ( .A(n3413), .ZN(n3415) );
  NAND2_X1 U4294 ( .A1(n3415), .A2(n3414), .ZN(n3428) );
  XNOR2_X1 U4295 ( .A(n3428), .B(n3426), .ZN(n3416) );
  NAND2_X1 U4296 ( .A1(n3416), .A2(n6037), .ZN(n3417) );
  NAND2_X1 U4297 ( .A1(n3418), .A2(n3417), .ZN(n3420) );
  INV_X1 U4298 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3419) );
  XNOR2_X1 U4299 ( .A(n3420), .B(n3419), .ZN(n4883) );
  NAND2_X1 U4300 ( .A1(n4882), .A2(n4883), .ZN(n3422) );
  NAND2_X1 U4301 ( .A1(n3420), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3421)
         );
  NAND2_X1 U4302 ( .A1(n3422), .A2(n3421), .ZN(n4932) );
  NOR2_X1 U4303 ( .A1(n3423), .A2(n3484), .ZN(n3424) );
  NAND2_X1 U4304 ( .A1(n6037), .A2(n3426), .ZN(n3427) );
  OR2_X1 U4305 ( .A1(n3428), .A2(n3427), .ZN(n3429) );
  NAND2_X1 U4306 ( .A1(n3440), .A2(n3429), .ZN(n3430) );
  INV_X1 U4307 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3579) );
  XNOR2_X1 U4308 ( .A(n3430), .B(n3579), .ZN(n4933) );
  NAND2_X1 U4309 ( .A1(n4932), .A2(n4933), .ZN(n3432) );
  NAND2_X1 U4310 ( .A1(n3430), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3431)
         );
  NAND2_X1 U4311 ( .A1(n3432), .A2(n3431), .ZN(n5039) );
  INV_X1 U4312 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5053) );
  NOR2_X1 U4313 ( .A1(n3447), .A2(n5053), .ZN(n3433) );
  NOR2_X1 U4314 ( .A1(n5039), .A2(n3433), .ZN(n3434) );
  INV_X1 U4315 ( .A(n3434), .ZN(n3436) );
  NAND2_X1 U4316 ( .A1(n3447), .A2(n5053), .ZN(n3435) );
  NAND2_X1 U4317 ( .A1(n3436), .A2(n3435), .ZN(n5045) );
  INV_X1 U4318 ( .A(n5045), .ZN(n3437) );
  INV_X1 U4319 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5052) );
  NAND2_X1 U4320 ( .A1(n3437), .A2(n3004), .ZN(n5141) );
  OR2_X1 U4321 ( .A1(n3447), .A2(n5052), .ZN(n5142) );
  INV_X1 U4322 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6151) );
  OR2_X1 U4323 ( .A1(n3440), .A2(n6151), .ZN(n5143) );
  AND2_X1 U4324 ( .A1(n5142), .A2(n5143), .ZN(n5151) );
  INV_X1 U4325 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3439) );
  NOR2_X1 U4326 ( .A1(n3440), .A2(n3439), .ZN(n5524) );
  XNOR2_X1 U4327 ( .A(n3440), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5531)
         );
  INV_X1 U4328 ( .A(n5531), .ZN(n3441) );
  INV_X1 U4329 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5515) );
  NAND2_X1 U4330 ( .A1(n5141), .A2(n3438), .ZN(n5126) );
  NAND2_X1 U4331 ( .A1(n3447), .A2(n6151), .ZN(n5153) );
  INV_X1 U4332 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U4333 ( .A1(n3447), .A2(n5622), .ZN(n3442) );
  NAND2_X1 U4334 ( .A1(n3440), .A2(n3439), .ZN(n5526) );
  OR2_X1 U4335 ( .A1(n3441), .A2(n5526), .ZN(n5528) );
  AND2_X1 U4336 ( .A1(n3442), .A2(n5528), .ZN(n5514) );
  NAND2_X1 U4337 ( .A1(n3447), .A2(n5515), .ZN(n3443) );
  AND2_X1 U4338 ( .A1(n5514), .A2(n3443), .ZN(n3444) );
  INV_X1 U4339 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U4340 ( .A1(n5126), .A2(n3445), .ZN(n3446) );
  NAND2_X1 U4341 ( .A1(n3446), .A2(n5127), .ZN(n5492) );
  INV_X1 U4342 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U4343 ( .A1(n3447), .A2(n5620), .ZN(n3448) );
  NAND2_X1 U4344 ( .A1(n5492), .A2(n3448), .ZN(n5495) );
  INV_X1 U4345 ( .A(n5495), .ZN(n3449) );
  NAND2_X1 U4346 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3650) );
  NAND2_X1 U4347 ( .A1(n3449), .A2(n3003), .ZN(n3451) );
  INV_X1 U4348 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U4349 ( .A1(n5603), .A2(n5620), .ZN(n5494) );
  OAI21_X1 U4350 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5494), .A(n5596), 
        .ZN(n3450) );
  AND2_X2 U4351 ( .A1(n3451), .A2(n3450), .ZN(n5751) );
  INV_X1 U4352 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5750) );
  NAND2_X2 U4353 ( .A1(n5751), .A2(n5750), .ZN(n5749) );
  NAND2_X1 U4354 ( .A1(n5749), .A2(n5596), .ZN(n3453) );
  INV_X1 U4355 ( .A(n5752), .ZN(n5468) );
  NAND2_X1 U4356 ( .A1(n5468), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3452) );
  NAND2_X1 U4357 ( .A1(n3453), .A2(n3452), .ZN(n5487) );
  XNOR2_X1 U4358 ( .A(n3447), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5488)
         );
  INV_X1 U4359 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5587) );
  NOR2_X1 U4360 ( .A1(n3440), .A2(n5587), .ZN(n3454) );
  AOI21_X1 U4361 ( .B1(n5487), .B2(n5488), .A(n3454), .ZN(n5482) );
  XNOR2_X1 U4362 ( .A(n3440), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5483)
         );
  NOR2_X1 U4363 ( .A1(n3447), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5455)
         );
  AOI21_X1 U4364 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n3447), .A(n5455), 
        .ZN(n3458) );
  INV_X1 U4365 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3660) );
  AND2_X1 U4366 ( .A1(n3447), .A2(n3660), .ZN(n3456) );
  OR2_X1 U4367 ( .A1(n3458), .A2(n3456), .ZN(n3455) );
  OR2_X1 U4368 ( .A1(n5480), .A2(n3455), .ZN(n3460) );
  INV_X1 U4369 ( .A(n5454), .ZN(n3457) );
  NAND2_X1 U4370 ( .A1(n3458), .A2(n3457), .ZN(n3459) );
  NAND2_X1 U4371 ( .A1(n3460), .A2(n3459), .ZN(n5248) );
  INV_X1 U4372 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3502) );
  NAND2_X1 U4373 ( .A1(n6439), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3462) );
  NAND2_X1 U4374 ( .A1(n4332), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3461) );
  NAND2_X1 U4375 ( .A1(n3462), .A2(n3461), .ZN(n3482) );
  NAND2_X1 U4376 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6369), .ZN(n3480) );
  NAND2_X1 U4377 ( .A1(n3463), .A2(n3462), .ZN(n3476) );
  MUX2_X1 U4378 ( .A(n3248), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n3474) );
  NAND2_X1 U4379 ( .A1(n3476), .A2(n3474), .ZN(n3465) );
  NAND2_X1 U4380 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n3248), .ZN(n3464) );
  NAND2_X1 U4381 ( .A1(n3465), .A2(n3464), .ZN(n3469) );
  XNOR2_X1 U4382 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3470) );
  NAND2_X1 U4383 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3503), .ZN(n3466) );
  NOR2_X1 U4384 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n3466), .ZN(n3472)
         );
  INV_X1 U4385 ( .A(n3467), .ZN(n3468) );
  OAI21_X1 U4386 ( .B1(n3470), .B2(n3469), .A(n3468), .ZN(n3471) );
  NAND2_X1 U4387 ( .A1(n3513), .A2(n3485), .ZN(n3499) );
  NAND2_X1 U4388 ( .A1(n4475), .A2(n3510), .ZN(n3473) );
  INV_X1 U4389 ( .A(n3474), .ZN(n3475) );
  XNOR2_X1 U4390 ( .A(n3476), .B(n3475), .ZN(n3517) );
  NAND2_X1 U4391 ( .A1(n3517), .A2(n3507), .ZN(n3496) );
  INV_X1 U4392 ( .A(n3517), .ZN(n3477) );
  NAND2_X1 U4393 ( .A1(n3478), .A2(n3477), .ZN(n3479) );
  AND3_X1 U4394 ( .A1(n3497), .A2(n3479), .A3(n3496), .ZN(n3495) );
  OAI21_X1 U4395 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6369), .A(n3480), 
        .ZN(n3487) );
  OAI21_X1 U4396 ( .B1(n3538), .B2(n3487), .A(n3106), .ZN(n3483) );
  AOI21_X1 U4397 ( .B1(n3507), .B2(n3545), .A(n5289), .ZN(n3490) );
  INV_X1 U4398 ( .A(n3480), .ZN(n3481) );
  XNOR2_X1 U4399 ( .A(n3482), .B(n3481), .ZN(n3515) );
  NAND2_X1 U4400 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n3515), .ZN(n3489) );
  AOI22_X1 U4401 ( .A1(n3497), .A2(n3483), .B1(n3490), .B2(n3489), .ZN(n3493)
         );
  INV_X1 U4402 ( .A(n3507), .ZN(n3486) );
  INV_X1 U4403 ( .A(n3504), .ZN(n3488) );
  OAI21_X1 U4404 ( .B1(n3487), .B2(n3486), .A(n3488), .ZN(n3492) );
  OAI22_X1 U4405 ( .A1(n3490), .A2(n3489), .B1(n3488), .B2(n3515), .ZN(n3491)
         );
  AOI21_X1 U4406 ( .B1(n3493), .B2(n3492), .A(n3491), .ZN(n3494) );
  OAI22_X1 U4407 ( .A1(n3497), .A2(n3496), .B1(n3495), .B2(n3494), .ZN(n3498)
         );
  NAND2_X1 U4408 ( .A1(n3499), .A2(n3498), .ZN(n3501) );
  NAND2_X1 U4409 ( .A1(n3513), .A2(n3504), .ZN(n3500) );
  OAI211_X1 U4410 ( .C1(STATE2_REG_0__SCAN_IN), .C2(n3502), .A(n3501), .B(
        n3500), .ZN(n3506) );
  OAI222_X1 U4411 ( .A1(n3502), .A2(n3503), .B1(n3502), .B2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C1(n3503), .C2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3519) );
  NAND2_X1 U4412 ( .A1(n3519), .A2(n3504), .ZN(n3505) );
  NAND2_X1 U4413 ( .A1(n3506), .A2(n3505), .ZN(n3509) );
  NAND2_X1 U4414 ( .A1(n3519), .A2(n3507), .ZN(n3508) );
  INV_X1 U4415 ( .A(n4322), .ZN(n4275) );
  NAND2_X1 U4416 ( .A1(n3170), .A2(n3510), .ZN(n3521) );
  OR2_X1 U4417 ( .A1(n5267), .A2(n4475), .ZN(n3630) );
  INV_X1 U4418 ( .A(n3630), .ZN(n3511) );
  NAND2_X1 U4419 ( .A1(n4275), .A2(n3511), .ZN(n4303) );
  NAND2_X1 U4420 ( .A1(n3512), .A2(n6500), .ZN(n6495) );
  NAND2_X1 U4421 ( .A1(n3545), .A2(n6495), .ZN(n3520) );
  INV_X1 U4422 ( .A(n3513), .ZN(n3514) );
  AND2_X1 U4423 ( .A1(n3515), .A2(n3514), .ZN(n3516) );
  AND2_X1 U4424 ( .A1(n3517), .A2(n3516), .ZN(n3518) );
  OR2_X1 U4425 ( .A1(n3519), .A2(n3518), .ZN(n4272) );
  NOR2_X1 U4426 ( .A1(READY_N), .A2(n4272), .ZN(n4291) );
  NAND3_X1 U4427 ( .A1(n3520), .A2(n4291), .A3(n3636), .ZN(n3528) );
  NAND2_X1 U4428 ( .A1(n3521), .A2(n4506), .ZN(n3522) );
  AND2_X1 U4429 ( .A1(n3634), .A2(n3522), .ZN(n3539) );
  INV_X1 U4430 ( .A(n3164), .ZN(n3523) );
  AND2_X1 U4431 ( .A1(n3523), .A2(n6037), .ZN(n3524) );
  NOR2_X1 U4432 ( .A1(n3525), .A2(n3524), .ZN(n3639) );
  NAND2_X1 U4433 ( .A1(n3539), .A2(n3639), .ZN(n3527) );
  NAND2_X1 U4434 ( .A1(n3527), .A2(n4266), .ZN(n4300) );
  NAND3_X1 U4435 ( .A1(n4303), .A2(n3528), .A3(n4300), .ZN(n3530) );
  NAND2_X1 U4436 ( .A1(n3530), .A2(n6473), .ZN(n3536) );
  INV_X1 U4437 ( .A(READY_N), .ZN(n6761) );
  AND2_X1 U4438 ( .A1(n3545), .A2(n6761), .ZN(n4370) );
  INV_X1 U4439 ( .A(n4370), .ZN(n3533) );
  INV_X1 U4440 ( .A(n6495), .ZN(n3532) );
  NAND2_X1 U4441 ( .A1(n3532), .A2(n6761), .ZN(n4908) );
  NAND2_X1 U4442 ( .A1(n3533), .A2(n4908), .ZN(n4902) );
  INV_X1 U4443 ( .A(n4902), .ZN(n4296) );
  OAI211_X1 U4444 ( .C1(n4313), .C2(n4296), .A(n3106), .B(n3635), .ZN(n3534)
         );
  NAND3_X1 U4445 ( .A1(n6035), .A2(n4497), .A3(n3534), .ZN(n3535) );
  INV_X1 U4446 ( .A(n3537), .ZN(n4950) );
  AND2_X1 U4447 ( .A1(n3539), .A2(n4950), .ZN(n4288) );
  INV_X1 U4448 ( .A(n4288), .ZN(n4330) );
  INV_X1 U4449 ( .A(n6453), .ZN(n4269) );
  NAND2_X1 U4450 ( .A1(n3541), .A2(n3540), .ZN(n3542) );
  NAND4_X1 U4451 ( .A1(n3543), .A2(n4330), .A3(n4269), .A4(n3542), .ZN(n3544)
         );
  NOR2_X1 U4452 ( .A1(n5248), .A2(n5636), .ZN(n3667) );
  INV_X1 U4453 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3547) );
  NAND2_X1 U4454 ( .A1(n3565), .A2(n3547), .ZN(n3551) );
  NAND2_X4 U4455 ( .A1(n4501), .A2(n3106), .ZN(n3683) );
  INV_X1 U4456 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3546) );
  NAND2_X1 U4457 ( .A1(n3683), .A2(n3546), .ZN(n3549) );
  NAND2_X1 U4458 ( .A1(n4349), .A2(n3547), .ZN(n3548) );
  NAND3_X1 U4459 ( .A1(n3549), .A2(n2989), .A3(n3548), .ZN(n3550) );
  NAND2_X1 U4460 ( .A1(n3551), .A2(n3550), .ZN(n3554) );
  NAND2_X1 U4461 ( .A1(n3683), .A2(EBX_REG_0__SCAN_IN), .ZN(n3553) );
  INV_X1 U4462 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5015) );
  NAND2_X1 U4463 ( .A1(n2989), .A2(n5015), .ZN(n3552) );
  NAND2_X1 U4464 ( .A1(n3553), .A2(n3552), .ZN(n4260) );
  XNOR2_X1 U4465 ( .A(n3554), .B(n4260), .ZN(n4350) );
  NAND2_X1 U4466 ( .A1(n4350), .A2(n4349), .ZN(n4352) );
  NAND2_X1 U4467 ( .A1(n4352), .A2(n3554), .ZN(n4441) );
  INV_X1 U4468 ( .A(n3683), .ZN(n3556) );
  NAND2_X1 U4469 ( .A1(n3556), .A2(n2990), .ZN(n3621) );
  NAND2_X1 U4470 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n2990), .ZN(n3557)
         );
  AND2_X1 U4471 ( .A1(n3621), .A2(n3557), .ZN(n3558) );
  MUX2_X1 U4472 ( .A(n3673), .B(n2989), .S(EBX_REG_3__SCAN_IN), .Z(n3562) );
  OAI21_X1 U4473 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n5236), .A(n3562), 
        .ZN(n4400) );
  INV_X1 U4474 ( .A(EBX_REG_4__SCAN_IN), .ZN(n3567) );
  NAND2_X1 U4475 ( .A1(n4223), .A2(n3567), .ZN(n3571) );
  NAND2_X1 U4476 ( .A1(n3683), .A2(n3566), .ZN(n3569) );
  NAND2_X1 U4477 ( .A1(n4349), .A2(n3567), .ZN(n3568) );
  NAND3_X1 U4478 ( .A1(n3569), .A2(n2989), .A3(n3568), .ZN(n3570) );
  MUX2_X1 U4479 ( .A(n3673), .B(n2989), .S(EBX_REG_5__SCAN_IN), .Z(n3572) );
  NAND2_X1 U4480 ( .A1(n4567), .A2(n4566), .ZN(n4739) );
  MUX2_X1 U4481 ( .A(n3670), .B(n3683), .S(EBX_REG_6__SCAN_IN), .Z(n3575) );
  NAND2_X1 U4482 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n2990), .ZN(n3573)
         );
  AND2_X1 U4483 ( .A1(n3621), .A2(n3573), .ZN(n3574) );
  MUX2_X1 U4484 ( .A(n3673), .B(n2989), .S(EBX_REG_7__SCAN_IN), .Z(n3578) );
  NAND2_X1 U4485 ( .A1(n3001), .A2(n3578), .ZN(n4890) );
  INV_X1 U4486 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U4487 ( .A1(n4223), .A2(n5908), .ZN(n3583) );
  NAND2_X1 U4488 ( .A1(n3683), .A2(n3579), .ZN(n3581) );
  NAND2_X1 U4489 ( .A1(n4349), .A2(n5908), .ZN(n3580) );
  NAND3_X1 U4490 ( .A1(n3581), .A2(n2989), .A3(n3580), .ZN(n3582) );
  NAND2_X1 U4491 ( .A1(n3583), .A2(n3582), .ZN(n4935) );
  NAND2_X1 U4492 ( .A1(n4936), .A2(n4935), .ZN(n5027) );
  MUX2_X1 U4493 ( .A(n3673), .B(n2989), .S(EBX_REG_9__SCAN_IN), .Z(n3584) );
  NAND2_X1 U4494 ( .A1(n3000), .A2(n3584), .ZN(n5028) );
  NOR2_X2 U4495 ( .A1(n5027), .A2(n5028), .ZN(n5026) );
  MUX2_X1 U4496 ( .A(n3670), .B(n3683), .S(EBX_REG_10__SCAN_IN), .Z(n3587) );
  NAND2_X1 U4497 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n2990), .ZN(n3585) );
  AND2_X1 U4498 ( .A1(n3621), .A2(n3585), .ZN(n3586) );
  NAND2_X1 U4499 ( .A1(n3587), .A2(n3586), .ZN(n5049) );
  AND2_X2 U4500 ( .A1(n5026), .A2(n5049), .ZN(n5048) );
  INV_X1 U4501 ( .A(n3673), .ZN(n3679) );
  INV_X1 U4502 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5111) );
  NAND2_X1 U4503 ( .A1(n3679), .A2(n5111), .ZN(n3590) );
  NAND2_X1 U4504 ( .A1(n2989), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3588) );
  OAI211_X1 U4505 ( .C1(n2990), .C2(EBX_REG_11__SCAN_IN), .A(n3683), .B(n3588), 
        .ZN(n3589) );
  MUX2_X1 U4506 ( .A(n3670), .B(n3683), .S(EBX_REG_12__SCAN_IN), .Z(n3593) );
  NAND2_X1 U4507 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n2990), .ZN(n3591) );
  AND2_X1 U4508 ( .A1(n3621), .A2(n3591), .ZN(n3592) );
  NAND2_X1 U4509 ( .A1(n3593), .A2(n3592), .ZN(n5158) );
  NAND2_X1 U4510 ( .A1(n5113), .A2(n5158), .ZN(n5157) );
  NAND2_X1 U4511 ( .A1(n2989), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3594) );
  OAI211_X1 U4512 ( .C1(n2990), .C2(EBX_REG_13__SCAN_IN), .A(n3683), .B(n3594), 
        .ZN(n3595) );
  OAI21_X1 U4513 ( .B1(n3673), .B2(EBX_REG_13__SCAN_IN), .A(n3595), .ZN(n5782)
         );
  NOR2_X2 U4514 ( .A1(n5157), .A2(n5782), .ZN(n5414) );
  MUX2_X1 U4515 ( .A(n3670), .B(n3683), .S(EBX_REG_14__SCAN_IN), .Z(n3598) );
  NAND2_X1 U4516 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n2990), .ZN(n3596) );
  AND2_X1 U4517 ( .A1(n3621), .A2(n3596), .ZN(n3597) );
  NAND2_X1 U4518 ( .A1(n2989), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3600) );
  OAI211_X1 U4519 ( .C1(n2990), .C2(EBX_REG_15__SCAN_IN), .A(n3683), .B(n3600), 
        .ZN(n3601) );
  OAI21_X1 U4520 ( .B1(n3673), .B2(EBX_REG_15__SCAN_IN), .A(n3601), .ZN(n5130)
         );
  MUX2_X1 U4521 ( .A(n3670), .B(n3683), .S(EBX_REG_16__SCAN_IN), .Z(n3604) );
  NAND2_X1 U4522 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n2990), .ZN(n3602) );
  AND2_X1 U4523 ( .A1(n3621), .A2(n3602), .ZN(n3603) );
  NAND2_X1 U4524 ( .A1(n3604), .A2(n3603), .ZN(n5406) );
  NAND2_X1 U4525 ( .A1(n2989), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3605) );
  OAI211_X1 U4526 ( .C1(n2990), .C2(EBX_REG_17__SCAN_IN), .A(n3683), .B(n3605), 
        .ZN(n3606) );
  OAI21_X1 U4527 ( .B1(n3673), .B2(EBX_REG_17__SCAN_IN), .A(n3606), .ZN(n5600)
         );
  OR2_X2 U4528 ( .A1(n5405), .A2(n5600), .ZN(n5602) );
  INV_X1 U4529 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5727) );
  NAND2_X1 U4530 ( .A1(n4223), .A2(n5727), .ZN(n3610) );
  NAND2_X1 U4531 ( .A1(n3683), .A2(n5750), .ZN(n3608) );
  NAND2_X1 U4532 ( .A1(n4349), .A2(n5727), .ZN(n3607) );
  NAND3_X1 U4533 ( .A1(n3608), .A2(n2989), .A3(n3607), .ZN(n3609) );
  AND2_X1 U4534 ( .A1(n3610), .A2(n3609), .ZN(n5713) );
  NOR2_X2 U4535 ( .A1(n5602), .A2(n5713), .ZN(n5384) );
  INV_X1 U4536 ( .A(n5236), .ZN(n3633) );
  NOR2_X1 U4537 ( .A1(n2990), .A2(EBX_REG_20__SCAN_IN), .ZN(n3611) );
  AOI21_X1 U4538 ( .B1(n3633), .B2(n5587), .A(n3611), .ZN(n5386) );
  OR2_X1 U4539 ( .A1(n5236), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3612)
         );
  INV_X1 U4540 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U4541 ( .A1(n4349), .A2(n5404), .ZN(n5397) );
  NAND2_X1 U4542 ( .A1(n3612), .A2(n5397), .ZN(n5398) );
  INV_X1 U4543 ( .A(EBX_REG_20__SCAN_IN), .ZN(n3613) );
  NOR2_X1 U4544 ( .A1(n2989), .A2(n3613), .ZN(n3614) );
  AOI21_X1 U4545 ( .B1(n5398), .B2(n2989), .A(n3614), .ZN(n3615) );
  OAI21_X1 U4546 ( .B1(n5386), .B2(n5398), .A(n3615), .ZN(n3616) );
  INV_X1 U4547 ( .A(n3616), .ZN(n3617) );
  AND2_X2 U4548 ( .A1(n5384), .A2(n3617), .ZN(n5381) );
  MUX2_X1 U4549 ( .A(n3673), .B(n2989), .S(EBX_REG_21__SCAN_IN), .Z(n3618) );
  OAI21_X1 U4550 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5236), .A(n3618), 
        .ZN(n3619) );
  INV_X1 U4551 ( .A(n3619), .ZN(n5380) );
  NAND2_X1 U4552 ( .A1(n5381), .A2(n5380), .ZN(n3624) );
  MUX2_X1 U4553 ( .A(n3670), .B(n3683), .S(EBX_REG_22__SCAN_IN), .Z(n3623) );
  NAND2_X1 U4554 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n2990), .ZN(n3620) );
  AND2_X1 U4555 ( .A1(n3621), .A2(n3620), .ZN(n3622) );
  AND2_X1 U4556 ( .A1(n3623), .A2(n3622), .ZN(n3625) );
  NAND2_X1 U4557 ( .A1(n3624), .A2(n3625), .ZN(n3626) );
  NAND2_X1 U4558 ( .A1(n5565), .A2(n3626), .ZN(n5685) );
  OR2_X1 U4559 ( .A1(n4313), .A2(n6581), .ZN(n6034) );
  INV_X1 U4560 ( .A(n4372), .ZN(n3627) );
  NAND3_X1 U4561 ( .A1(n3627), .A2(n4493), .A3(n5287), .ZN(n3628) );
  NAND2_X1 U4562 ( .A1(n6034), .A2(n3628), .ZN(n3629) );
  NAND2_X1 U4563 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4934) );
  INV_X1 U4564 ( .A(n4934), .ZN(n5051) );
  NAND3_X1 U4565 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n5051), .ZN(n5135) );
  AOI21_X1 U4566 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n4398) );
  NAND2_X1 U4567 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4460) );
  NOR2_X1 U4568 ( .A1(n4398), .A2(n4460), .ZN(n4746) );
  NAND3_X1 U4569 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n4746), .ZN(n4888) );
  NOR2_X1 U4570 ( .A1(n5135), .A2(n4888), .ZN(n3657) );
  NAND3_X1 U4571 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5630) );
  OR2_X1 U4572 ( .A1(n5515), .A2(n5630), .ZN(n5137) );
  NAND2_X1 U4573 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5617) );
  NOR2_X1 U4574 ( .A1(n5137), .A2(n5617), .ZN(n3645) );
  NAND2_X1 U4575 ( .A1(n3657), .A2(n3645), .ZN(n5582) );
  INV_X1 U4576 ( .A(n5582), .ZN(n3653) );
  NOR2_X1 U4577 ( .A1(n3630), .A2(n4506), .ZN(n3631) );
  NAND2_X1 U4578 ( .A1(n4300), .A2(n3631), .ZN(n4331) );
  INV_X1 U4579 ( .A(n4331), .ZN(n3632) );
  NAND2_X1 U4580 ( .A1(n3647), .A2(n3632), .ZN(n5162) );
  AND2_X1 U4581 ( .A1(n4271), .A2(n3545), .ZN(n5266) );
  INV_X1 U4582 ( .A(n5625), .ZN(n4258) );
  OR2_X1 U4583 ( .A1(n3634), .A2(n3633), .ZN(n3638) );
  NAND2_X1 U4584 ( .A1(n3635), .A2(n3636), .ZN(n3637) );
  NAND2_X1 U4585 ( .A1(n4506), .A2(n3545), .ZN(n4953) );
  OR2_X1 U4586 ( .A1(n4953), .A2(n3636), .ZN(n4299) );
  NAND4_X1 U4587 ( .A1(n3639), .A2(n3638), .A3(n3637), .A4(n4299), .ZN(n3640)
         );
  NOR2_X1 U4588 ( .A1(n3641), .A2(n3640), .ZN(n4315) );
  NAND2_X1 U4589 ( .A1(n4501), .A2(n4506), .ZN(n3642) );
  OR2_X1 U4590 ( .A1(n5267), .A2(n3642), .ZN(n4418) );
  OAI211_X1 U4591 ( .C1(n4372), .C2(n3145), .A(n4315), .B(n4418), .ZN(n3643)
         );
  NAND2_X1 U4592 ( .A1(n3647), .A2(n3643), .ZN(n5624) );
  INV_X1 U4593 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6168) );
  NOR2_X1 U4594 ( .A1(n6168), .A2(n3546), .ZN(n4397) );
  INV_X1 U4595 ( .A(n4397), .ZN(n3644) );
  NOR2_X1 U4596 ( .A1(n3644), .A2(n4460), .ZN(n4750) );
  NAND3_X1 U4597 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n4750), .ZN(n4885) );
  NOR2_X1 U4598 ( .A1(n4885), .A2(n5135), .ZN(n3656) );
  AND2_X1 U4599 ( .A1(n3656), .A2(n3645), .ZN(n3646) );
  OR2_X1 U4600 ( .A1(n4884), .A2(n3646), .ZN(n3649) );
  NOR2_X1 U4601 ( .A1(n5624), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3648)
         );
  NOR2_X1 U4602 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6488) );
  AND2_X2 U4603 ( .A1(n6564), .A2(n6488), .ZN(n6159) );
  NOR2_X1 U4604 ( .A1(n3647), .A2(n6159), .ZN(n4363) );
  NOR2_X1 U4605 ( .A1(n3648), .A2(n4363), .ZN(n5585) );
  AND2_X1 U4606 ( .A1(n3649), .A2(n5585), .ZN(n5605) );
  NAND2_X1 U4607 ( .A1(n4884), .A2(n5162), .ZN(n5214) );
  INV_X1 U4608 ( .A(n3650), .ZN(n5589) );
  AND2_X1 U4609 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5467) );
  AND2_X1 U4610 ( .A1(n5589), .A2(n5467), .ZN(n3659) );
  INV_X1 U4611 ( .A(n3659), .ZN(n3651) );
  NAND2_X1 U4612 ( .A1(n5214), .A2(n3651), .ZN(n3652) );
  OAI211_X1 U4613 ( .C1(n3653), .C2(n5162), .A(n5605), .B(n3652), .ZN(n5578)
         );
  AND2_X1 U4614 ( .A1(n6159), .A2(REIP_REG_22__SCAN_IN), .ZN(n5251) );
  AOI21_X1 U4615 ( .B1(n5578), .B2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5251), 
        .ZN(n3654) );
  OAI21_X1 U4616 ( .B1(n5685), .B2(n5631), .A(n3654), .ZN(n3655) );
  INV_X1 U4617 ( .A(n3655), .ZN(n3665) );
  NOR2_X1 U4618 ( .A1(n5625), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4365)
         );
  NAND2_X1 U4619 ( .A1(n6169), .A2(n3656), .ZN(n5163) );
  NAND2_X1 U4620 ( .A1(n6162), .A2(n3657), .ZN(n5623) );
  NAND2_X1 U4621 ( .A1(n5163), .A2(n5623), .ZN(n6146) );
  INV_X1 U4622 ( .A(n5617), .ZN(n3658) );
  NAND2_X1 U4623 ( .A1(n5776), .A2(n3659), .ZN(n5581) );
  INV_X1 U4624 ( .A(n5581), .ZN(n3663) );
  NOR2_X1 U4625 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4199) );
  INV_X1 U4626 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3661) );
  NOR2_X1 U4627 ( .A1(n3661), .A2(n3660), .ZN(n5466) );
  NOR2_X1 U4628 ( .A1(n4199), .A2(n5466), .ZN(n3662) );
  NAND2_X1 U4629 ( .A1(n3665), .A2(n3664), .ZN(n3666) );
  INV_X1 U4630 ( .A(n5385), .ZN(n5396) );
  NAND2_X1 U4631 ( .A1(n2989), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3668) );
  OAI211_X1 U4632 ( .C1(n2990), .C2(EBX_REG_23__SCAN_IN), .A(n3683), .B(n3668), 
        .ZN(n3669) );
  OAI21_X1 U4633 ( .B1(n3673), .B2(EBX_REG_23__SCAN_IN), .A(n3669), .ZN(n5564)
         );
  NOR2_X4 U4634 ( .A1(n5565), .A2(n5564), .ZN(n5567) );
  MUX2_X1 U4635 ( .A(n3670), .B(n3683), .S(EBX_REG_24__SCAN_IN), .Z(n3672) );
  NAND2_X1 U4636 ( .A1(n2990), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3671) );
  NAND2_X1 U4637 ( .A1(n3672), .A2(n3671), .ZN(n5345) );
  MUX2_X1 U4638 ( .A(n3673), .B(n2989), .S(EBX_REG_25__SCAN_IN), .Z(n3674) );
  OAI21_X1 U4639 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5236), .A(n3674), 
        .ZN(n5369) );
  INV_X1 U4640 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U4641 ( .A1(n4223), .A2(n5658), .ZN(n3678) );
  INV_X1 U4642 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U4643 ( .A1(n3683), .A2(n5537), .ZN(n3676) );
  NAND2_X1 U4644 ( .A1(n4349), .A2(n5658), .ZN(n3675) );
  NAND3_X1 U4645 ( .A1(n3676), .A2(n2989), .A3(n3675), .ZN(n3677) );
  AND2_X1 U4646 ( .A1(n3678), .A2(n3677), .ZN(n5360) );
  NOR2_X2 U4647 ( .A1(n2999), .A2(n5360), .ZN(n5197) );
  INV_X1 U4648 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5722) );
  NAND2_X1 U4649 ( .A1(n3679), .A2(n5722), .ZN(n3682) );
  NAND2_X1 U4650 ( .A1(n2989), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3680) );
  OAI211_X1 U4651 ( .C1(n2990), .C2(EBX_REG_27__SCAN_IN), .A(n3683), .B(n3680), 
        .ZN(n3681) );
  AND2_X1 U4652 ( .A1(n3682), .A2(n3681), .ZN(n5198) );
  AND2_X2 U4653 ( .A1(n5197), .A2(n5198), .ZN(n5200) );
  INV_X1 U4654 ( .A(EBX_REG_28__SCAN_IN), .ZN(n3684) );
  NAND2_X1 U4655 ( .A1(n4223), .A2(n3684), .ZN(n3688) );
  INV_X1 U4656 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U4657 ( .A1(n3683), .A2(n5190), .ZN(n3686) );
  NAND2_X1 U4658 ( .A1(n4349), .A2(n3684), .ZN(n3685) );
  NAND3_X1 U4659 ( .A1(n3686), .A2(n2989), .A3(n3685), .ZN(n3687) );
  NAND2_X1 U4660 ( .A1(n3688), .A2(n3687), .ZN(n5183) );
  AND2_X4 U4661 ( .A1(n5200), .A2(n5183), .ZN(n5184) );
  INV_X1 U4662 ( .A(n5184), .ZN(n4224) );
  AND2_X1 U4663 ( .A1(n2990), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3689)
         );
  AOI21_X1 U4664 ( .B1(n5236), .B2(EBX_REG_30__SCAN_IN), .A(n3689), .ZN(n5231)
         );
  OR2_X1 U4665 ( .A1(n5236), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3691)
         );
  INV_X1 U4666 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5357) );
  NAND2_X1 U4667 ( .A1(n4349), .A2(n5357), .ZN(n3690) );
  AND2_X1 U4668 ( .A1(n3691), .A2(n3690), .ZN(n4226) );
  AOI211_X1 U4669 ( .C1(n5396), .C2(n4224), .A(n5231), .B(n3692), .ZN(n3697)
         );
  NOR2_X1 U4670 ( .A1(n3692), .A2(n5396), .ZN(n5233) );
  INV_X1 U4671 ( .A(n5231), .ZN(n3693) );
  AOI21_X1 U4672 ( .B1(n4225), .B2(n5184), .A(n3693), .ZN(n3694) );
  INV_X1 U4673 ( .A(n5288), .ZN(n5310) );
  NAND3_X1 U4674 ( .A1(n5310), .A2(n4493), .A3(n3698), .ZN(n4371) );
  OR3_X1 U4675 ( .A1(n4371), .A2(n3699), .A3(n2990), .ZN(n3700) );
  OAI21_X1 U4676 ( .B1(n4331), .B2(n4322), .A(n3700), .ZN(n3701) );
  NAND2_X1 U4677 ( .A1(n3702), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4041) );
  NAND2_X1 U4678 ( .A1(n6466), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3842) );
  OAI21_X2 U4679 ( .B1(n4607), .B2(n4041), .A(n3842), .ZN(n3721) );
  NAND2_X1 U4680 ( .A1(n4467), .A2(n4020), .ZN(n3706) );
  AOI22_X1 U4681 ( .A1(n5300), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6466), .ZN(n3704) );
  AND2_X1 U4682 ( .A1(n5287), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3732) );
  NAND2_X1 U4683 ( .A1(n3732), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3703) );
  AND2_X1 U4684 ( .A1(n3704), .A2(n3703), .ZN(n3705) );
  NAND2_X1 U4685 ( .A1(n3706), .A2(n3705), .ZN(n4347) );
  NAND2_X1 U4686 ( .A1(n6304), .A2(n3121), .ZN(n3707) );
  NAND2_X1 U4687 ( .A1(n3707), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4354) );
  INV_X1 U4688 ( .A(n3732), .ZN(n3729) );
  CLKBUF_X1 U4689 ( .A(n3709), .Z(n3710) );
  NAND2_X1 U4690 ( .A1(n5300), .A2(EAX_REG_0__SCAN_IN), .ZN(n3712) );
  NAND2_X1 U4691 ( .A1(n6466), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3711)
         );
  OAI211_X1 U4692 ( .C1(n3729), .C2(n3710), .A(n3712), .B(n3711), .ZN(n3713)
         );
  AOI21_X1 U4693 ( .B1(n6314), .B2(n4020), .A(n3713), .ZN(n3714) );
  INV_X1 U4694 ( .A(n3714), .ZN(n4356) );
  OR2_X1 U4695 ( .A1(n4356), .A2(n4164), .ZN(n3715) );
  NAND2_X1 U4696 ( .A1(n4355), .A2(n3715), .ZN(n4348) );
  INV_X1 U4697 ( .A(n3720), .ZN(n4346) );
  OAI21_X1 U4698 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3725), .ZN(n6132) );
  AOI22_X1 U4699 ( .A1(n5299), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n4191), 
        .B2(n6132), .ZN(n3719) );
  NAND2_X1 U4700 ( .A1(n5300), .A2(EAX_REG_2__SCAN_IN), .ZN(n3718) );
  OAI211_X1 U4701 ( .C1(n3729), .C2(n3717), .A(n3719), .B(n3718), .ZN(n4444)
         );
  NAND2_X1 U4702 ( .A1(n4445), .A2(n4444), .ZN(n3723) );
  NAND2_X1 U4703 ( .A1(n3721), .A2(n3720), .ZN(n3722) );
  NAND2_X1 U4704 ( .A1(n3723), .A2(n3722), .ZN(n4403) );
  OAI21_X1 U4705 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3726), .A(n3734), 
        .ZN(n5964) );
  AOI22_X1 U4706 ( .A1(n4191), .A2(n5964), .B1(n5299), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3728) );
  NAND2_X1 U4707 ( .A1(n5300), .A2(EAX_REG_3__SCAN_IN), .ZN(n3727) );
  OAI211_X1 U4708 ( .C1(n3729), .C2(n4411), .A(n3728), .B(n3727), .ZN(n3730)
         );
  INV_X1 U4709 ( .A(n3730), .ZN(n3731) );
  OAI21_X1 U4710 ( .B1(n4608), .B2(n4041), .A(n3731), .ZN(n4404) );
  NAND2_X1 U4711 ( .A1(n4403), .A2(n4404), .ZN(n4450) );
  NAND2_X1 U4712 ( .A1(n3732), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3736) );
  AOI21_X1 U4713 ( .B1(n5943), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3733) );
  AOI21_X1 U4714 ( .B1(n5300), .B2(EAX_REG_4__SCAN_IN), .A(n3733), .ZN(n3735)
         );
  AOI21_X1 U4715 ( .B1(n5943), .B2(n3734), .A(n3739), .ZN(n5946) );
  AOI22_X1 U4716 ( .A1(n3736), .A2(n3735), .B1(n4191), .B2(n5946), .ZN(n3737)
         );
  AOI21_X1 U4717 ( .B1(n3738), .B2(n4020), .A(n3737), .ZN(n4449) );
  NOR2_X2 U4718 ( .A1(n4450), .A2(n4449), .ZN(n4565) );
  OAI21_X1 U4719 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3739), .A(n3750), 
        .ZN(n5935) );
  AOI22_X1 U4720 ( .A1(n4191), .A2(n5935), .B1(n5299), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3741) );
  NAND2_X1 U4721 ( .A1(n5300), .A2(EAX_REG_5__SCAN_IN), .ZN(n3740) );
  OAI211_X1 U4722 ( .C1(n3742), .C2(n4041), .A(n3741), .B(n3740), .ZN(n4564)
         );
  NAND2_X1 U4723 ( .A1(n4565), .A2(n4564), .ZN(n4799) );
  INV_X1 U4724 ( .A(n4799), .ZN(n3748) );
  NAND2_X1 U4725 ( .A1(n5300), .A2(EAX_REG_6__SCAN_IN), .ZN(n3744) );
  OAI21_X1 U4726 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6723), .A(n6466), 
        .ZN(n3743) );
  XOR2_X1 U4727 ( .A(n3749), .B(n3750), .Z(n4919) );
  AOI22_X1 U4728 ( .A1(n3744), .A2(n3743), .B1(n4191), .B2(n4919), .ZN(n3745)
         );
  NAND2_X1 U4729 ( .A1(n3748), .A2(n3747), .ZN(n4797) );
  INV_X1 U4730 ( .A(n4797), .ZN(n3759) );
  INV_X1 U4731 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3755) );
  OR2_X1 U4732 ( .A1(n3751), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3752) );
  NAND2_X1 U4733 ( .A1(n3752), .A2(n3760), .ZN(n5915) );
  NAND2_X1 U4734 ( .A1(n5915), .A2(n4191), .ZN(n3754) );
  NAND2_X1 U4735 ( .A1(n5299), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3753)
         );
  OAI211_X1 U4736 ( .C1(n3824), .C2(n3755), .A(n3754), .B(n3753), .ZN(n3756)
         );
  NAND2_X1 U4737 ( .A1(n3759), .A2(n3758), .ZN(n4941) );
  XOR2_X1 U4738 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3775), .Z(n5903) );
  INV_X1 U4739 ( .A(n5903), .ZN(n4946) );
  AOI22_X1 U4740 ( .A1(n4175), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4133), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4741 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n3197), .B1(n4176), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4742 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n4168), .B1(n4413), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4743 ( .A1(n4167), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3761) );
  NAND4_X1 U4744 ( .A1(n3764), .A2(n3763), .A3(n3762), .A4(n3761), .ZN(n3770)
         );
  AOI22_X1 U4745 ( .A1(n4178), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4746 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n3259), .B1(n4169), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4747 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n4103), .B1(n2983), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4748 ( .A1(n3195), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3765) );
  NAND4_X1 U4749 ( .A1(n3768), .A2(n3767), .A3(n3766), .A4(n3765), .ZN(n3769)
         );
  OAI21_X1 U4750 ( .B1(n3770), .B2(n3769), .A(n4020), .ZN(n3773) );
  NAND2_X1 U4751 ( .A1(n5300), .A2(EAX_REG_8__SCAN_IN), .ZN(n3772) );
  NAND2_X1 U4752 ( .A1(n5299), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3771)
         );
  NAND3_X1 U4753 ( .A1(n3773), .A2(n3772), .A3(n3771), .ZN(n3774) );
  AOI21_X1 U4754 ( .B1(n4946), .B2(n4191), .A(n3774), .ZN(n4942) );
  NOR2_X2 U4755 ( .A1(n4941), .A2(n4942), .ZN(n5025) );
  XNOR2_X1 U4756 ( .A(n3791), .B(n5034), .ZN(n5041) );
  NAND2_X1 U4757 ( .A1(n5041), .A2(n4191), .ZN(n3790) );
  AOI22_X1 U4758 ( .A1(n4167), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4133), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4759 ( .A1(n3195), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4760 ( .A1(n4168), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4761 ( .A1(n3202), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3776) );
  NAND4_X1 U4762 ( .A1(n3779), .A2(n3778), .A3(n3777), .A4(n3776), .ZN(n3785)
         );
  AOI22_X1 U4763 ( .A1(n4175), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4764 ( .A1(n3259), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4765 ( .A1(n3219), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4766 ( .A1(n4178), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3780) );
  NAND4_X1 U4767 ( .A1(n3783), .A2(n3782), .A3(n3781), .A4(n3780), .ZN(n3784)
         );
  OAI21_X1 U4768 ( .B1(n3785), .B2(n3784), .A(n4020), .ZN(n3787) );
  NAND2_X1 U4769 ( .A1(n5300), .A2(EAX_REG_9__SCAN_IN), .ZN(n3786) );
  OAI211_X1 U4770 ( .C1(n3842), .C2(n5034), .A(n3787), .B(n3786), .ZN(n3788)
         );
  INV_X1 U4771 ( .A(n3788), .ZN(n3789) );
  NAND2_X1 U4772 ( .A1(n3790), .A2(n3789), .ZN(n5024) );
  XOR2_X1 U4773 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3806), .Z(n5892) );
  AOI22_X1 U4774 ( .A1(n4167), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4178), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4775 ( .A1(n3197), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4776 ( .A1(n4133), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4777 ( .A1(n4176), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3792) );
  NAND4_X1 U4778 ( .A1(n3795), .A2(n3794), .A3(n3793), .A4(n3792), .ZN(n3801)
         );
  AOI22_X1 U4779 ( .A1(n3195), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4780 ( .A1(n4168), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4781 ( .A1(n3202), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4782 ( .A1(n3259), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3796) );
  NAND4_X1 U4783 ( .A1(n3799), .A2(n3798), .A3(n3797), .A4(n3796), .ZN(n3800)
         );
  OAI21_X1 U4784 ( .B1(n3801), .B2(n3800), .A(n4020), .ZN(n3804) );
  NAND2_X1 U4785 ( .A1(n5300), .A2(EAX_REG_10__SCAN_IN), .ZN(n3803) );
  NAND2_X1 U4786 ( .A1(n5299), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3802)
         );
  AND3_X1 U4787 ( .A1(n3804), .A2(n3803), .A3(n3802), .ZN(n3805) );
  OAI21_X1 U4788 ( .B1(n5892), .B2(n4164), .A(n3805), .ZN(n5059) );
  XNOR2_X1 U4789 ( .A(n3822), .B(n5119), .ZN(n5146) );
  NAND2_X1 U4790 ( .A1(n5146), .A2(n4191), .ZN(n3821) );
  AOI22_X1 U4791 ( .A1(n4167), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4133), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4792 ( .A1(n3195), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4793 ( .A1(n3202), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4794 ( .A1(n4175), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3807) );
  NAND4_X1 U4795 ( .A1(n3810), .A2(n3809), .A3(n3808), .A4(n3807), .ZN(n3816)
         );
  AOI22_X1 U4796 ( .A1(n3197), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4797 ( .A1(n4168), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4798 ( .A1(n4178), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4799 ( .A1(n4169), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3811) );
  NAND4_X1 U4800 ( .A1(n3814), .A2(n3813), .A3(n3812), .A4(n3811), .ZN(n3815)
         );
  OAI21_X1 U4801 ( .B1(n3816), .B2(n3815), .A(n4020), .ZN(n3818) );
  NAND2_X1 U4802 ( .A1(n5300), .A2(EAX_REG_11__SCAN_IN), .ZN(n3817) );
  OAI211_X1 U4803 ( .C1(n3842), .C2(n5119), .A(n3818), .B(n3817), .ZN(n3819)
         );
  INV_X1 U4804 ( .A(n3819), .ZN(n3820) );
  NAND2_X1 U4805 ( .A1(n3821), .A2(n3820), .ZN(n5106) );
  NAND2_X1 U4806 ( .A1(n5107), .A2(n5106), .ZN(n5105) );
  INV_X1 U4807 ( .A(n5105), .ZN(n3840) );
  XOR2_X1 U4808 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3841), .Z(n5880) );
  NAND2_X1 U4809 ( .A1(n5880), .A2(n4191), .ZN(n3838) );
  INV_X1 U4810 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5169) );
  OAI21_X1 U4811 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6723), .A(n6466), 
        .ZN(n3823) );
  OAI21_X1 U4812 ( .B1(n3824), .B2(n5169), .A(n3823), .ZN(n3837) );
  AOI22_X1 U4813 ( .A1(n4167), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4133), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4814 ( .A1(n4169), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4815 ( .A1(n4175), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4816 ( .A1(n3197), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3825) );
  NAND4_X1 U4817 ( .A1(n3828), .A2(n3827), .A3(n3826), .A4(n3825), .ZN(n3834)
         );
  AOI22_X1 U4818 ( .A1(n4178), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4819 ( .A1(n4168), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4820 ( .A1(n2983), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4821 ( .A1(n3195), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3829) );
  NAND4_X1 U4822 ( .A1(n3832), .A2(n3831), .A3(n3830), .A4(n3829), .ZN(n3833)
         );
  NOR2_X1 U4823 ( .A1(n3834), .A2(n3833), .ZN(n3835) );
  NOR2_X1 U4824 ( .A1(n4041), .A2(n3835), .ZN(n3836) );
  AOI21_X1 U4825 ( .B1(n3838), .B2(n3837), .A(n3836), .ZN(n5168) );
  NAND2_X1 U4826 ( .A1(n3840), .A2(n3839), .ZN(n3857) );
  XNOR2_X1 U4827 ( .A(n3885), .B(n5865), .ZN(n5868) );
  NAND2_X1 U4828 ( .A1(n5868), .A2(n4191), .ZN(n3845) );
  NOR2_X1 U4829 ( .A1(n3842), .A2(n5865), .ZN(n3843) );
  AOI21_X1 U4830 ( .B1(n5300), .B2(EAX_REG_13__SCAN_IN), .A(n3843), .ZN(n3844)
         );
  NAND2_X1 U4831 ( .A1(n3845), .A2(n3844), .ZN(n3858) );
  XNOR2_X1 U4832 ( .A(n3857), .B(n3858), .ZN(n5521) );
  AOI22_X1 U4833 ( .A1(n3195), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4834 ( .A1(n4175), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4835 ( .A1(n4168), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4836 ( .A1(n3197), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3846) );
  NAND4_X1 U4837 ( .A1(n3849), .A2(n3848), .A3(n3847), .A4(n3846), .ZN(n3855)
         );
  AOI22_X1 U4838 ( .A1(n4178), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4839 ( .A1(n4133), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4840 ( .A1(n2983), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4841 ( .A1(n4167), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4179), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3850) );
  NAND4_X1 U4842 ( .A1(n3853), .A2(n3852), .A3(n3851), .A4(n3850), .ZN(n3854)
         );
  OR2_X1 U4843 ( .A1(n3855), .A2(n3854), .ZN(n3856) );
  AND2_X1 U4844 ( .A1(n4020), .A2(n3856), .ZN(n5522) );
  NAND2_X1 U4845 ( .A1(n5521), .A2(n5522), .ZN(n3860) );
  NAND2_X1 U4846 ( .A1(n3860), .A2(n3859), .ZN(n5252) );
  AOI22_X1 U4847 ( .A1(n4178), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4848 ( .A1(n3195), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4849 ( .A1(n4169), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4850 ( .A1(n4167), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3861) );
  NAND4_X1 U4851 ( .A1(n3864), .A2(n3863), .A3(n3862), .A4(n3861), .ZN(n3870)
         );
  AOI22_X1 U4852 ( .A1(n4175), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4133), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4853 ( .A1(n4168), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4854 ( .A1(n2983), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4855 ( .A1(n4176), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3865) );
  NAND4_X1 U4856 ( .A1(n3868), .A2(n3867), .A3(n3866), .A4(n3865), .ZN(n3869)
         );
  NOR2_X1 U4857 ( .A1(n3870), .A2(n3869), .ZN(n4048) );
  AOI22_X1 U4858 ( .A1(n4178), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4859 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n3195), .B1(n4169), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4860 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n3197), .B1(n4176), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4861 ( .A1(n4167), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3871) );
  NAND4_X1 U4862 ( .A1(n3874), .A2(n3873), .A3(n3872), .A4(n3871), .ZN(n3880)
         );
  AOI22_X1 U4863 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n3259), .B1(n4133), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4864 ( .A1(n4168), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4865 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n4179), .B1(n2983), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4866 ( .A1(n4175), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3875) );
  NAND4_X1 U4867 ( .A1(n3878), .A2(n3877), .A3(n3876), .A4(n3875), .ZN(n3879)
         );
  NOR2_X1 U4868 ( .A1(n3880), .A2(n3879), .ZN(n4049) );
  XNOR2_X1 U4869 ( .A(n4048), .B(n4049), .ZN(n3884) );
  NAND2_X1 U4870 ( .A1(n6466), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3881)
         );
  NAND2_X1 U4871 ( .A1(n4164), .A2(n3881), .ZN(n3882) );
  AOI21_X1 U4872 ( .B1(n5300), .B2(EAX_REG_23__SCAN_IN), .A(n3882), .ZN(n3883)
         );
  OAI21_X1 U4873 ( .B1(n4161), .B2(n3884), .A(n3883), .ZN(n3890) );
  INV_X1 U4874 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4011) );
  INV_X1 U4875 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5499) );
  INV_X1 U4876 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5249) );
  OR2_X1 U4877 ( .A1(n3887), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3888)
         );
  NAND2_X1 U4878 ( .A1(n4080), .A2(n3888), .ZN(n5675) );
  OR2_X1 U4879 ( .A1(n5675), .A2(n4164), .ZN(n3889) );
  NAND2_X1 U4880 ( .A1(n3890), .A2(n3889), .ZN(n5475) );
  INV_X1 U4881 ( .A(n5475), .ZN(n4046) );
  AOI22_X1 U4882 ( .A1(n4167), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4883 ( .A1(n4168), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4133), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4884 ( .A1(n4178), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4885 ( .A1(n4179), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3891) );
  NAND4_X1 U4886 ( .A1(n3894), .A2(n3893), .A3(n3892), .A4(n3891), .ZN(n3902)
         );
  AOI22_X1 U4887 ( .A1(n3202), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4888 ( .A1(n4176), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3899) );
  AOI21_X1 U4889 ( .B1(n2983), .B2(INSTQUEUE_REG_6__6__SCAN_IN), .A(n4191), 
        .ZN(n3896) );
  NAND2_X1 U4890 ( .A1(n3219), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3895)
         );
  AND2_X1 U4891 ( .A1(n3896), .A2(n3895), .ZN(n3898) );
  AOI22_X1 U4892 ( .A1(n3195), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3897) );
  NAND4_X1 U4893 ( .A1(n3900), .A2(n3899), .A3(n3898), .A4(n3897), .ZN(n3901)
         );
  NAND2_X1 U4894 ( .A1(n4161), .A2(n4164), .ZN(n3970) );
  OAI21_X1 U4895 ( .B1(n3902), .B2(n3901), .A(n3970), .ZN(n3905) );
  NOR2_X1 U4896 ( .A1(n5249), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3903) );
  AOI21_X1 U4897 ( .B1(n5300), .B2(EAX_REG_22__SCAN_IN), .A(n3903), .ZN(n3904)
         );
  NAND2_X1 U4898 ( .A1(n3905), .A2(n3904), .ZN(n3907) );
  XNOR2_X1 U4899 ( .A(n3922), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5683)
         );
  NAND2_X1 U4900 ( .A1(n5683), .A2(n4191), .ZN(n3906) );
  NAND2_X1 U4901 ( .A1(n3907), .A2(n3906), .ZN(n5256) );
  INV_X1 U4902 ( .A(n5256), .ZN(n4045) );
  AOI22_X1 U4903 ( .A1(n4133), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4904 ( .A1(n3195), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4905 ( .A1(n3197), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4906 ( .A1(n4179), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3908) );
  NAND4_X1 U4907 ( .A1(n3911), .A2(n3910), .A3(n3909), .A4(n3908), .ZN(n3917)
         );
  AOI22_X1 U4908 ( .A1(n4178), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4909 ( .A1(n4175), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4910 ( .A1(n4167), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4911 ( .A1(n4168), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3912) );
  NAND4_X1 U4912 ( .A1(n3915), .A2(n3914), .A3(n3913), .A4(n3912), .ZN(n3916)
         );
  NOR2_X1 U4913 ( .A1(n3917), .A2(n3916), .ZN(n3921) );
  OAI21_X1 U4914 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6723), .A(n6466), 
        .ZN(n3918) );
  INV_X1 U4915 ( .A(n3918), .ZN(n3919) );
  AOI21_X1 U4916 ( .B1(n5300), .B2(EAX_REG_21__SCAN_IN), .A(n3919), .ZN(n3920)
         );
  OAI21_X1 U4917 ( .B1(n4161), .B2(n3921), .A(n3920), .ZN(n3925) );
  OAI21_X1 U4918 ( .B1(n3923), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n3922), 
        .ZN(n5693) );
  OR2_X1 U4919 ( .A1(n5693), .A2(n4164), .ZN(n3924) );
  AND2_X1 U4920 ( .A1(n3925), .A2(n3924), .ZN(n5377) );
  AOI22_X1 U4921 ( .A1(n3202), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4133), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3931) );
  NAND2_X1 U4922 ( .A1(n4167), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3927) );
  NAND2_X1 U4923 ( .A1(n4413), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3926)
         );
  AND3_X1 U4924 ( .A1(n3927), .A2(n3926), .A3(n4164), .ZN(n3930) );
  AOI22_X1 U4925 ( .A1(n4175), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4926 ( .A1(n3259), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3928) );
  NAND4_X1 U4927 ( .A1(n3931), .A2(n3930), .A3(n3929), .A4(n3928), .ZN(n3937)
         );
  AOI22_X1 U4928 ( .A1(n3195), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4168), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4929 ( .A1(n3197), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4178), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4930 ( .A1(n4169), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4931 ( .A1(n4176), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4179), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3932) );
  NAND4_X1 U4932 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n3936)
         );
  OR2_X1 U4933 ( .A1(n3937), .A2(n3936), .ZN(n3938) );
  NAND2_X1 U4934 ( .A1(n3970), .A2(n3938), .ZN(n3941) );
  AOI22_X1 U4935 ( .A1(n5300), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6466), .ZN(n3940) );
  XNOR2_X1 U4936 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n3956), .ZN(n5699)
         );
  AND2_X1 U4937 ( .A1(n5699), .A2(n4191), .ZN(n3939) );
  AOI21_X1 U4938 ( .B1(n3941), .B2(n3940), .A(n3939), .ZN(n5389) );
  AOI22_X1 U4939 ( .A1(n4167), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4940 ( .A1(n4176), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4941 ( .A1(n3219), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4942 ( .A1(n4133), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3942) );
  NAND4_X1 U4943 ( .A1(n3945), .A2(n3944), .A3(n3943), .A4(n3942), .ZN(n3951)
         );
  AOI22_X1 U4944 ( .A1(n3195), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4945 ( .A1(n3259), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4946 ( .A1(n4168), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4947 ( .A1(n4178), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3946) );
  NAND4_X1 U4948 ( .A1(n3949), .A2(n3948), .A3(n3947), .A4(n3946), .ZN(n3950)
         );
  NOR2_X1 U4949 ( .A1(n3951), .A2(n3950), .ZN(n3955) );
  NAND2_X1 U4950 ( .A1(n6466), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3952)
         );
  NAND2_X1 U4951 ( .A1(n4164), .A2(n3952), .ZN(n3953) );
  AOI21_X1 U4952 ( .B1(n5300), .B2(EAX_REG_19__SCAN_IN), .A(n3953), .ZN(n3954)
         );
  OAI21_X1 U4953 ( .B1(n4161), .B2(n3955), .A(n3954), .ZN(n3959) );
  OAI21_X1 U4954 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n3957), .A(n3956), 
        .ZN(n5758) );
  OR2_X1 U4955 ( .A1(n4164), .A2(n5758), .ZN(n3958) );
  NAND2_X1 U4956 ( .A1(n3959), .A2(n3958), .ZN(n5709) );
  INV_X1 U4957 ( .A(n5709), .ZN(n4044) );
  AOI22_X1 U4958 ( .A1(n4167), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4959 ( .A1(n4176), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4133), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4960 ( .A1(n3202), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4961 ( .A1(n4169), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3960) );
  NAND4_X1 U4962 ( .A1(n3963), .A2(n3962), .A3(n3961), .A4(n3960), .ZN(n3972)
         );
  AOI22_X1 U4963 ( .A1(n4175), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3969) );
  NAND2_X1 U4964 ( .A1(n4168), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3965) );
  NAND2_X1 U4965 ( .A1(n4178), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3964) );
  AND3_X1 U4966 ( .A1(n3965), .A2(n3964), .A3(n4164), .ZN(n3968) );
  AOI22_X1 U4967 ( .A1(n3195), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4968 ( .A1(n3259), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3966) );
  NAND4_X1 U4969 ( .A1(n3969), .A2(n3968), .A3(n3967), .A4(n3966), .ZN(n3971)
         );
  OAI21_X1 U4970 ( .B1(n3972), .B2(n3971), .A(n3970), .ZN(n3975) );
  NOR2_X1 U4971 ( .A1(n5499), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3973) );
  AOI21_X1 U4972 ( .B1(n5300), .B2(EAX_REG_18__SCAN_IN), .A(n3973), .ZN(n3974)
         );
  NAND2_X1 U4973 ( .A1(n3975), .A2(n3974), .ZN(n3977) );
  XNOR2_X1 U4974 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3992), .ZN(n5815)
         );
  NAND2_X1 U4975 ( .A1(n4191), .A2(n5815), .ZN(n3976) );
  NAND2_X1 U4976 ( .A1(n3977), .A2(n3976), .ZN(n5394) );
  INV_X1 U4977 ( .A(n5394), .ZN(n4043) );
  AOI22_X1 U4978 ( .A1(n3195), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4979 ( .A1(n3197), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4980 ( .A1(n4168), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4981 ( .A1(n4103), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3978) );
  NAND4_X1 U4982 ( .A1(n3981), .A2(n3980), .A3(n3979), .A4(n3978), .ZN(n3987)
         );
  AOI22_X1 U4983 ( .A1(n4178), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4984 ( .A1(n4133), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4985 ( .A1(n4167), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4986 ( .A1(n4175), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3982) );
  NAND4_X1 U4987 ( .A1(n3985), .A2(n3984), .A3(n3983), .A4(n3982), .ZN(n3986)
         );
  NOR2_X1 U4988 ( .A1(n3987), .A2(n3986), .ZN(n3991) );
  NAND2_X1 U4989 ( .A1(n6466), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3988)
         );
  NAND2_X1 U4990 ( .A1(n4164), .A2(n3988), .ZN(n3989) );
  AOI21_X1 U4991 ( .B1(n5300), .B2(EAX_REG_17__SCAN_IN), .A(n3989), .ZN(n3990)
         );
  OAI21_X1 U4992 ( .B1(n4161), .B2(n3991), .A(n3990), .ZN(n3995) );
  OAI21_X1 U4993 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3993), .A(n3992), 
        .ZN(n5832) );
  OR2_X1 U4994 ( .A1(n4164), .A2(n5832), .ZN(n3994) );
  AND2_X1 U4995 ( .A1(n3995), .A2(n3994), .ZN(n5759) );
  XNOR2_X1 U4996 ( .A(n3996), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5840)
         );
  AOI22_X1 U4997 ( .A1(n4178), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4998 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n4169), .B1(n3259), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4999 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n3197), .B1(n4176), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U5000 ( .A1(n4167), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3997) );
  NAND4_X1 U5001 ( .A1(n4000), .A2(n3999), .A3(n3998), .A4(n3997), .ZN(n4006)
         );
  AOI22_X1 U5002 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n3195), .B1(n4133), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U5003 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4168), .B1(n4413), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U5004 ( .A1(n4103), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U5005 ( .A1(n4175), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4001) );
  NAND4_X1 U5006 ( .A1(n4004), .A2(n4003), .A3(n4002), .A4(n4001), .ZN(n4005)
         );
  NOR2_X1 U5007 ( .A1(n4006), .A2(n4005), .ZN(n4008) );
  AOI22_X1 U5008 ( .A1(n5300), .A2(EAX_REG_16__SCAN_IN), .B1(n5299), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4007) );
  OAI21_X1 U5009 ( .B1(n4161), .B2(n4008), .A(n4007), .ZN(n4009) );
  AOI21_X1 U5010 ( .B1(n5840), .B2(n4191), .A(n4009), .ZN(n5409) );
  XOR2_X1 U5011 ( .A(n4011), .B(n4010), .Z(n5847) );
  INV_X1 U5012 ( .A(n5847), .ZN(n5509) );
  AOI22_X1 U5013 ( .A1(n4167), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U5014 ( .A1(n4175), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U5015 ( .A1(n3219), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U5016 ( .A1(n3224), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4012) );
  NAND4_X1 U5017 ( .A1(n4015), .A2(n4014), .A3(n4013), .A4(n4012), .ZN(n4022)
         );
  AOI22_X1 U5018 ( .A1(n4178), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4133), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U5019 ( .A1(n4169), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U5020 ( .A1(n3195), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U5021 ( .A1(n4168), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4016) );
  NAND4_X1 U5022 ( .A1(n4019), .A2(n4018), .A3(n4017), .A4(n4016), .ZN(n4021)
         );
  OAI21_X1 U5023 ( .B1(n4022), .B2(n4021), .A(n4020), .ZN(n4025) );
  NAND2_X1 U5024 ( .A1(n5300), .A2(EAX_REG_15__SCAN_IN), .ZN(n4024) );
  NAND2_X1 U5025 ( .A1(n5299), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4023)
         );
  NAND3_X1 U5026 ( .A1(n4025), .A2(n4024), .A3(n4023), .ZN(n4026) );
  AOI21_X1 U5027 ( .B1(n5509), .B2(n4191), .A(n4026), .ZN(n5435) );
  NOR2_X1 U5028 ( .A1(n5409), .A2(n5435), .ZN(n5410) );
  AND2_X1 U5029 ( .A1(n5759), .A2(n5410), .ZN(n4042) );
  AOI22_X1 U5030 ( .A1(n4178), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U5031 ( .A1(n4133), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U5032 ( .A1(n4168), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U5033 ( .A1(n4103), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4027) );
  NAND4_X1 U5034 ( .A1(n4030), .A2(n4029), .A3(n4028), .A4(n4027), .ZN(n4036)
         );
  AOI22_X1 U5035 ( .A1(n3195), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U5036 ( .A1(n3219), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U5037 ( .A1(n4167), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U5038 ( .A1(n4176), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4031) );
  NAND4_X1 U5039 ( .A1(n4034), .A2(n4033), .A3(n4032), .A4(n4031), .ZN(n4035)
         );
  NOR2_X1 U5040 ( .A1(n4036), .A2(n4035), .ZN(n4040) );
  XNOR2_X1 U5041 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4037), .ZN(n5857)
         );
  AOI22_X1 U5042 ( .A1(n4191), .A2(n5857), .B1(n5299), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4039) );
  NAND2_X1 U5043 ( .A1(n5300), .A2(EAX_REG_14__SCAN_IN), .ZN(n4038) );
  OAI211_X1 U5044 ( .C1(n4041), .C2(n4040), .A(n4039), .B(n4038), .ZN(n5418)
         );
  AND2_X1 U5045 ( .A1(n4042), .A2(n5418), .ZN(n5393) );
  AND2_X1 U5046 ( .A1(n4043), .A2(n5393), .ZN(n5392) );
  AND2_X1 U5047 ( .A1(n4044), .A2(n5392), .ZN(n5388) );
  AND2_X1 U5048 ( .A1(n5389), .A2(n5388), .ZN(n5376) );
  NAND2_X1 U5049 ( .A1(n5252), .A2(n4047), .ZN(n5472) );
  INV_X1 U5050 ( .A(n4161), .ZN(n4188) );
  NOR2_X1 U5051 ( .A1(n4049), .A2(n4048), .ZN(n4066) );
  AOI22_X1 U5052 ( .A1(n3195), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U5053 ( .A1(n4175), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U5054 ( .A1(n4168), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U5055 ( .A1(n3197), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4050) );
  NAND4_X1 U5056 ( .A1(n4053), .A2(n4052), .A3(n4051), .A4(n4050), .ZN(n4059)
         );
  AOI22_X1 U5057 ( .A1(n4178), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U5058 ( .A1(n4133), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U5059 ( .A1(n2983), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U5060 ( .A1(n4167), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4054) );
  NAND4_X1 U5061 ( .A1(n4057), .A2(n4056), .A3(n4055), .A4(n4054), .ZN(n4058)
         );
  OR2_X1 U5062 ( .A1(n4059), .A2(n4058), .ZN(n4065) );
  INV_X1 U5063 ( .A(n4065), .ZN(n4060) );
  XNOR2_X1 U5064 ( .A(n4066), .B(n4060), .ZN(n4064) );
  XNOR2_X1 U5065 ( .A(n4080), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5460)
         );
  NAND2_X1 U5066 ( .A1(n5300), .A2(EAX_REG_24__SCAN_IN), .ZN(n4062) );
  NAND2_X1 U5067 ( .A1(n5299), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4061)
         );
  OAI211_X1 U5068 ( .C1(n5460), .C2(n4164), .A(n4062), .B(n4061), .ZN(n4063)
         );
  AOI21_X1 U5069 ( .B1(n4188), .B2(n4064), .A(n4063), .ZN(n5344) );
  NOR2_X1 U5070 ( .A1(n5472), .A2(n5344), .ZN(n5343) );
  NAND2_X1 U5071 ( .A1(n4066), .A2(n4065), .ZN(n4085) );
  AOI22_X1 U5072 ( .A1(n4168), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U5073 ( .A1(n4176), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U5074 ( .A1(n4167), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U5075 ( .A1(n4133), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4067) );
  NAND4_X1 U5076 ( .A1(n4070), .A2(n4069), .A3(n4068), .A4(n4067), .ZN(n4076)
         );
  AOI22_X1 U5077 ( .A1(n4178), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4074) );
  AOI22_X1 U5078 ( .A1(n3195), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U5079 ( .A1(n4169), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U5080 ( .A1(n4413), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4071) );
  NAND4_X1 U5081 ( .A1(n4074), .A2(n4073), .A3(n4072), .A4(n4071), .ZN(n4075)
         );
  NOR2_X1 U5082 ( .A1(n4076), .A2(n4075), .ZN(n4086) );
  XNOR2_X1 U5083 ( .A(n4085), .B(n4086), .ZN(n4079) );
  INV_X1 U5084 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5447) );
  OAI21_X1 U5085 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5447), .A(n4164), .ZN(
        n4077) );
  AOI21_X1 U5086 ( .B1(n5300), .B2(EAX_REG_25__SCAN_IN), .A(n4077), .ZN(n4078)
         );
  OAI21_X1 U5087 ( .B1(n4161), .B2(n4079), .A(n4078), .ZN(n4084) );
  INV_X1 U5088 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5462) );
  AND2_X1 U5089 ( .A1(n4081), .A2(n5447), .ZN(n4082) );
  NOR2_X1 U5090 ( .A1(n4082), .A2(n4120), .ZN(n5664) );
  NAND2_X1 U5091 ( .A1(n5664), .A2(n4191), .ZN(n4083) );
  NOR2_X1 U5092 ( .A1(n4086), .A2(n4085), .ZN(n4115) );
  AOI22_X1 U5093 ( .A1(n3195), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U5094 ( .A1(n4175), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U5095 ( .A1(n4168), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U5096 ( .A1(n3197), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4087) );
  NAND4_X1 U5097 ( .A1(n4090), .A2(n4089), .A3(n4088), .A4(n4087), .ZN(n4096)
         );
  AOI22_X1 U5098 ( .A1(n4178), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4094) );
  AOI22_X1 U5099 ( .A1(n4133), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4093) );
  AOI22_X1 U5100 ( .A1(n2983), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4092) );
  AOI22_X1 U5101 ( .A1(n4167), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4091) );
  NAND4_X1 U5102 ( .A1(n4094), .A2(n4093), .A3(n4092), .A4(n4091), .ZN(n4095)
         );
  OR2_X1 U5103 ( .A1(n4096), .A2(n4095), .ZN(n4114) );
  XNOR2_X1 U5104 ( .A(n4115), .B(n4114), .ZN(n4100) );
  NAND2_X1 U5105 ( .A1(n6466), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4097)
         );
  NAND2_X1 U5106 ( .A1(n4164), .A2(n4097), .ZN(n4098) );
  AOI21_X1 U5107 ( .B1(n5300), .B2(EAX_REG_26__SCAN_IN), .A(n4098), .ZN(n4099)
         );
  OAI21_X1 U5108 ( .B1(n4100), .B2(n4161), .A(n4099), .ZN(n4102) );
  INV_X1 U5109 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5443) );
  XNOR2_X1 U5110 ( .A(n4120), .B(n5443), .ZN(n5649) );
  NAND2_X1 U5111 ( .A1(n5649), .A2(n4191), .ZN(n4101) );
  AOI22_X1 U5112 ( .A1(n4169), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U5113 ( .A1(n3195), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U5114 ( .A1(n4178), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U5115 ( .A1(n4133), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4104) );
  NAND4_X1 U5116 ( .A1(n4107), .A2(n4106), .A3(n4105), .A4(n4104), .ZN(n4113)
         );
  AOI22_X1 U5117 ( .A1(n4168), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4111) );
  AOI22_X1 U5118 ( .A1(n4167), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4110) );
  AOI22_X1 U5119 ( .A1(n3202), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5120 ( .A1(n4176), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4108) );
  NAND4_X1 U5121 ( .A1(n4111), .A2(n4110), .A3(n4109), .A4(n4108), .ZN(n4112)
         );
  NOR2_X1 U5122 ( .A1(n4113), .A2(n4112), .ZN(n4128) );
  NAND2_X1 U5123 ( .A1(n4115), .A2(n4114), .ZN(n4127) );
  XNOR2_X1 U5124 ( .A(n4128), .B(n4127), .ZN(n4119) );
  NAND2_X1 U5125 ( .A1(n6466), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4116)
         );
  NAND2_X1 U5126 ( .A1(n4164), .A2(n4116), .ZN(n4117) );
  AOI21_X1 U5127 ( .B1(n5300), .B2(EAX_REG_27__SCAN_IN), .A(n4117), .ZN(n4118)
         );
  OAI21_X1 U5128 ( .B1(n4119), .B2(n4161), .A(n4118), .ZN(n4126) );
  INV_X1 U5129 ( .A(n4121), .ZN(n4123) );
  INV_X1 U5130 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4122) );
  NAND2_X1 U5131 ( .A1(n4123), .A2(n4122), .ZN(n4124) );
  NAND2_X1 U5132 ( .A1(n4144), .A2(n4124), .ZN(n5648) );
  NAND2_X1 U5133 ( .A1(n4126), .A2(n4125), .ZN(n4246) );
  XNOR2_X1 U5134 ( .A(n4144), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5280)
         );
  INV_X1 U5135 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4213) );
  OAI21_X1 U5136 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4213), .A(n4164), .ZN(
        n4142) );
  NOR2_X1 U5137 ( .A1(n4128), .A2(n4127), .ZN(n4158) );
  AOI22_X1 U5138 ( .A1(n3195), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U5139 ( .A1(n4175), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U5140 ( .A1(n4168), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U5141 ( .A1(n3219), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4129) );
  NAND4_X1 U5142 ( .A1(n4132), .A2(n4131), .A3(n4130), .A4(n4129), .ZN(n4139)
         );
  AOI22_X1 U5143 ( .A1(n4178), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4137) );
  AOI22_X1 U5144 ( .A1(n4133), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U5145 ( .A1(n2983), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U5146 ( .A1(n4167), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4179), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4134) );
  NAND4_X1 U5147 ( .A1(n4137), .A2(n4136), .A3(n4135), .A4(n4134), .ZN(n4138)
         );
  OR2_X1 U5148 ( .A1(n4139), .A2(n4138), .ZN(n4157) );
  XNOR2_X1 U5149 ( .A(n4158), .B(n4157), .ZN(n4140) );
  NOR2_X1 U5150 ( .A1(n4140), .A2(n4161), .ZN(n4141) );
  AOI211_X1 U5151 ( .C1(n5300), .C2(EAX_REG_28__SCAN_IN), .A(n4142), .B(n4141), 
        .ZN(n4143) );
  AOI21_X1 U5152 ( .B1(n4191), .B2(n5280), .A(n4143), .ZN(n4215) );
  INV_X1 U5153 ( .A(n4145), .ZN(n4146) );
  INV_X1 U5154 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5335) );
  OAI21_X1 U5155 ( .B1(n4146), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n4898), 
        .ZN(n5334) );
  AOI22_X1 U5156 ( .A1(n4133), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U5157 ( .A1(n4168), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U5158 ( .A1(n3202), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U5159 ( .A1(n4167), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4147) );
  NAND4_X1 U5160 ( .A1(n4150), .A2(n4149), .A3(n4148), .A4(n4147), .ZN(n4156)
         );
  AOI22_X1 U5161 ( .A1(n3195), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5162 ( .A1(n3197), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4413), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U5163 ( .A1(n4178), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4179), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4152) );
  AOI22_X1 U5164 ( .A1(n4176), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4151) );
  NAND4_X1 U5165 ( .A1(n4154), .A2(n4153), .A3(n4152), .A4(n4151), .ZN(n4155)
         );
  NOR2_X1 U5166 ( .A1(n4156), .A2(n4155), .ZN(n4166) );
  NAND2_X1 U5167 ( .A1(n4158), .A2(n4157), .ZN(n4165) );
  XNOR2_X1 U5168 ( .A(n4166), .B(n4165), .ZN(n4162) );
  AOI21_X1 U5169 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6466), .A(n4191), 
        .ZN(n4160) );
  NAND2_X1 U5170 ( .A1(n5300), .A2(EAX_REG_29__SCAN_IN), .ZN(n4159) );
  OAI211_X1 U5171 ( .C1(n4162), .C2(n4161), .A(n4160), .B(n4159), .ZN(n4163)
         );
  OAI21_X1 U5172 ( .B1(n4164), .B2(n5334), .A(n4163), .ZN(n5260) );
  NOR2_X1 U5173 ( .A1(n4166), .A2(n4165), .ZN(n4187) );
  AOI22_X1 U5174 ( .A1(n4167), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U5175 ( .A1(n4168), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4173) );
  AOI22_X1 U5176 ( .A1(n4133), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4172) );
  AOI22_X1 U5177 ( .A1(n3195), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4170), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4171) );
  NAND4_X1 U5178 ( .A1(n4174), .A2(n4173), .A3(n4172), .A4(n4171), .ZN(n4185)
         );
  AOI22_X1 U5179 ( .A1(n4175), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4183) );
  AOI22_X1 U5180 ( .A1(n4413), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4176), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4182) );
  AOI22_X1 U5181 ( .A1(n4178), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4181) );
  AOI22_X1 U5182 ( .A1(n4179), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4180) );
  NAND4_X1 U5183 ( .A1(n4183), .A2(n4182), .A3(n4181), .A4(n4180), .ZN(n4184)
         );
  NOR2_X1 U5184 ( .A1(n4185), .A2(n4184), .ZN(n4186) );
  XNOR2_X1 U5185 ( .A(n4187), .B(n4186), .ZN(n4189) );
  NAND2_X1 U5186 ( .A1(n4189), .A2(n4188), .ZN(n4194) );
  INV_X1 U5187 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5222) );
  AOI21_X1 U5188 ( .B1(n5222), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4190) );
  AOI21_X1 U5189 ( .B1(n5300), .B2(EAX_REG_30__SCAN_IN), .A(n4190), .ZN(n4193)
         );
  XNOR2_X1 U5190 ( .A(n4898), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5326)
         );
  AOI21_X1 U5191 ( .B1(n4194), .B2(n4193), .A(n4192), .ZN(n5297) );
  INV_X1 U5192 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5328) );
  OR2_X1 U5193 ( .A1(n5988), .A2(n5328), .ZN(n4197) );
  INV_X1 U5194 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5569) );
  INV_X1 U5195 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5555) );
  NAND4_X1 U5196 ( .A1(n4199), .A2(n5587), .A3(n5569), .A4(n5555), .ZN(n4200)
         );
  INV_X1 U5197 ( .A(n5751), .ZN(n4201) );
  AND2_X1 U5198 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4236) );
  NAND4_X1 U5199 ( .A1(n4201), .A2(n5467), .A3(n4236), .A4(n5466), .ZN(n4202)
         );
  AND2_X2 U5200 ( .A1(n4203), .A2(n4202), .ZN(n5450) );
  XNOR2_X1 U5201 ( .A(n3447), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5451)
         );
  INV_X1 U5202 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5548) );
  NAND2_X2 U5203 ( .A1(n5449), .A2(n4204), .ZN(n5208) );
  INV_X1 U5204 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4206) );
  AND2_X1 U5205 ( .A1(n3440), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4205)
         );
  NOR2_X1 U5206 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5539) );
  OAI22_X1 U5207 ( .A1(n4207), .A2(n3009), .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n4206), .ZN(n4208) );
  XNOR2_X1 U5208 ( .A(n4208), .B(n5190), .ZN(n5194) );
  NOR2_X2 U5209 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6310) );
  NAND2_X1 U5210 ( .A1(n6374), .A2(n4209), .ZN(n6579) );
  NAND2_X1 U5211 ( .A1(n6579), .A2(n6476), .ZN(n4210) );
  NAND2_X1 U5212 ( .A1(n6476), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4212) );
  NAND2_X1 U5213 ( .A1(n6723), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4211) );
  NAND2_X1 U5214 ( .A1(n4212), .A2(n4211), .ZN(n6138) );
  NAND2_X1 U5215 ( .A1(n6159), .A2(REIP_REG_28__SCAN_IN), .ZN(n5189) );
  OAI21_X1 U5216 ( .B1(n5769), .B2(n4213), .A(n5189), .ZN(n4218) );
  NAND3_X1 U5217 ( .A1(n6476), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6486) );
  INV_X1 U5218 ( .A(n6486), .ZN(n4216) );
  NOR2_X1 U5219 ( .A1(n5293), .A2(n6142), .ZN(n4217) );
  OAI21_X1 U5220 ( .B1(n5194), .B2(n6135), .A(n4219), .ZN(U2958) );
  AND2_X1 U5221 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5187) );
  AND2_X1 U5222 ( .A1(n3440), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4242)
         );
  AND2_X1 U5223 ( .A1(n5187), .A2(n4242), .ZN(n4220) );
  NOR2_X1 U5224 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5188) );
  NAND2_X1 U5225 ( .A1(n5596), .A2(n5188), .ZN(n5207) );
  OR2_X1 U5226 ( .A1(n5207), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4221)
         );
  AND2_X2 U5227 ( .A1(n5229), .A2(n2991), .ZN(n4222) );
  NAND2_X1 U5228 ( .A1(n4223), .A2(n5357), .ZN(n4227) );
  NAND2_X1 U5229 ( .A1(n4226), .A2(n2989), .ZN(n4228) );
  NAND2_X1 U5230 ( .A1(n4228), .A2(n4227), .ZN(n4229) );
  NOR2_X1 U5231 ( .A1(n5184), .A2(n4229), .ZN(n4230) );
  OR2_X1 U5232 ( .A1(n5232), .A2(n4230), .ZN(n5356) );
  INV_X1 U5233 ( .A(n5356), .ZN(n4240) );
  INV_X1 U5234 ( .A(n5466), .ZN(n4233) );
  INV_X1 U5235 ( .A(n4236), .ZN(n4231) );
  NOR2_X1 U5236 ( .A1(n5574), .A2(n4231), .ZN(n5538) );
  AND2_X1 U5237 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U5238 ( .A1(n5538), .A2(n5540), .ZN(n5206) );
  INV_X1 U5239 ( .A(n5187), .ZN(n4232) );
  INV_X1 U5240 ( .A(n5214), .ZN(n5584) );
  INV_X1 U5241 ( .A(n5540), .ZN(n4237) );
  NOR2_X1 U5242 ( .A1(n6169), .A2(n6162), .ZN(n4235) );
  AND2_X1 U5243 ( .A1(n5214), .A2(n4233), .ZN(n4234) );
  NOR2_X1 U5244 ( .A1(n5578), .A2(n4234), .ZN(n5570) );
  OAI21_X1 U5245 ( .B1(n4236), .B2(n4235), .A(n5570), .ZN(n5560) );
  AOI21_X1 U5246 ( .B1(n4237), .B2(n5214), .A(n5560), .ZN(n5196) );
  OAI21_X1 U5247 ( .B1(n5187), .B2(n5584), .A(n5196), .ZN(n5213) );
  INV_X1 U5248 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6629) );
  NOR2_X1 U5249 ( .A1(n6134), .A2(n6629), .ZN(n5261) );
  AOI21_X1 U5250 ( .B1(n5213), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5261), 
        .ZN(n4238) );
  OAI21_X1 U5251 ( .B1(n5241), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n4238), 
        .ZN(n4239) );
  AOI21_X1 U5252 ( .B1(n4240), .B2(n6161), .A(n4239), .ZN(n4241) );
  INV_X1 U5253 ( .A(n4242), .ZN(n4243) );
  NOR2_X1 U5254 ( .A1(n5208), .A2(n4243), .ZN(n4244) );
  NOR2_X1 U5255 ( .A1(n4244), .A2(n3009), .ZN(n4245) );
  XNOR2_X1 U5256 ( .A(n4245), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5195)
         );
  NAND2_X1 U5257 ( .A1(n5195), .A2(n6129), .ZN(n4253) );
  AND2_X1 U5258 ( .A1(n5359), .A2(n4246), .ZN(n4248) );
  INV_X1 U5259 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6649) );
  NOR2_X1 U5260 ( .A1(n6134), .A2(n6649), .ZN(n5202) );
  NOR2_X1 U5261 ( .A1(n6133), .A2(n5648), .ZN(n4249) );
  AOI211_X1 U5262 ( .C1(n6139), .C2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5202), 
        .B(n4249), .ZN(n4250) );
  NAND2_X1 U5263 ( .A1(n4253), .A2(n4252), .ZN(U2959) );
  INV_X1 U5264 ( .A(n5624), .ZN(n4254) );
  NOR2_X1 U5265 ( .A1(n4254), .A2(n6162), .ZN(n5627) );
  NOR2_X1 U5266 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5627), .ZN(n4362)
         );
  OR2_X1 U5267 ( .A1(n4255), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4256)
         );
  NAND2_X1 U5268 ( .A1(n4257), .A2(n4256), .ZN(n6136) );
  NOR2_X1 U5269 ( .A1(n6136), .A2(n5636), .ZN(n4264) );
  INV_X1 U5270 ( .A(n4363), .ZN(n4259) );
  INV_X1 U5271 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4340) );
  AOI21_X1 U5272 ( .B1(n4259), .B2(n4258), .A(n4340), .ZN(n4263) );
  OR2_X1 U5273 ( .A1(n5236), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4261)
         );
  NAND2_X1 U5274 ( .A1(n4261), .A2(n4260), .ZN(n5013) );
  INV_X1 U5275 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6576) );
  OAI22_X1 U5276 ( .A1(n5631), .A2(n5013), .B1(n6576), .B2(n6134), .ZN(n4262)
         );
  OR4_X1 U5277 ( .A1(n4362), .A2(n4264), .A3(n4263), .A4(n4262), .ZN(U3018) );
  INV_X1 U5278 ( .A(n5266), .ZN(n6434) );
  AOI21_X1 U5279 ( .B1(n6434), .B2(n6034), .A(n6495), .ZN(n4265) );
  NOR2_X1 U5280 ( .A1(n6477), .A2(n6466), .ZN(n4434) );
  AND2_X1 U5281 ( .A1(n6030), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  NOR2_X1 U5282 ( .A1(n4272), .A2(n4266), .ZN(n4277) );
  OAI22_X1 U5283 ( .A1(n4322), .A2(n4950), .B1(n4277), .B2(n4278), .ZN(n5793)
         );
  INV_X1 U5284 ( .A(n4953), .ZN(n4267) );
  OR2_X1 U5285 ( .A1(n6037), .A2(n4267), .ZN(n4283) );
  AOI21_X1 U5286 ( .B1(n4283), .B2(n6495), .A(READY_N), .ZN(n6580) );
  NOR2_X1 U5287 ( .A1(n5793), .A2(n6580), .ZN(n6455) );
  INV_X1 U5288 ( .A(n6473), .ZN(n6481) );
  NOR2_X1 U5289 ( .A1(n6455), .A2(n6481), .ZN(n5799) );
  INV_X1 U5290 ( .A(MORE_REG_SCAN_IN), .ZN(n6763) );
  CLKBUF_X1 U5291 ( .A(n4268), .Z(n4297) );
  NAND3_X1 U5292 ( .A1(n4330), .A2(n4269), .A3(n4297), .ZN(n4270) );
  NAND2_X1 U5293 ( .A1(n4270), .A2(n4275), .ZN(n4274) );
  NAND2_X1 U5294 ( .A1(n4272), .A2(n4271), .ZN(n4273) );
  OAI211_X1 U5295 ( .C1(n4275), .C2(n4331), .A(n4274), .B(n4273), .ZN(n6454)
         );
  NAND2_X1 U5296 ( .A1(n5799), .A2(n6454), .ZN(n4276) );
  OAI21_X1 U5297 ( .B1(n5799), .B2(n6763), .A(n4276), .ZN(U3471) );
  NAND2_X1 U5298 ( .A1(n4277), .A2(n6473), .ZN(n5639) );
  INV_X1 U5299 ( .A(n6578), .ZN(n4281) );
  INV_X1 U5300 ( .A(n4283), .ZN(n4280) );
  AND2_X1 U5301 ( .A1(n6310), .A2(n6477), .ZN(n4914) );
  OR2_X1 U5302 ( .A1(n6036), .A2(n4914), .ZN(n5638) );
  OAI22_X1 U5303 ( .A1(n4281), .A2(n4280), .B1(READREQUEST_REG_SCAN_IN), .B2(
        n5638), .ZN(n4282) );
  OAI21_X1 U5304 ( .B1(n4283), .B2(n5639), .A(n4282), .ZN(U3474) );
  INV_X1 U5305 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U5306 ( .A1(n6013), .A2(n3106), .ZN(n4394) );
  AOI22_X1 U5307 ( .A1(n6031), .A2(UWORD_REG_10__SCAN_IN), .B1(n6024), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4284) );
  OAI21_X1 U5308 ( .B1(n6062), .B2(n4394), .A(n4284), .ZN(U2897) );
  INV_X1 U5309 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6070) );
  AOI22_X1 U5310 ( .A1(n6031), .A2(UWORD_REG_13__SCAN_IN), .B1(n6024), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4285) );
  OAI21_X1 U5311 ( .B1(n6070), .B2(n4394), .A(n4285), .ZN(U2894) );
  INV_X1 U5312 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6068) );
  AOI22_X1 U5313 ( .A1(n6031), .A2(UWORD_REG_12__SCAN_IN), .B1(n6024), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4286) );
  OAI21_X1 U5314 ( .B1(n6068), .B2(n4394), .A(n4286), .ZN(U2895) );
  INV_X1 U5315 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6056) );
  AOI22_X1 U5316 ( .A1(n6031), .A2(UWORD_REG_8__SCAN_IN), .B1(n6024), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4287) );
  OAI21_X1 U5317 ( .B1(n6056), .B2(n4394), .A(n4287), .ZN(U2899) );
  NAND2_X1 U5318 ( .A1(n6476), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6560) );
  INV_X1 U5319 ( .A(n6560), .ZN(n4474) );
  NAND2_X1 U5320 ( .A1(n4322), .A2(n4288), .ZN(n4294) );
  INV_X1 U5321 ( .A(n4290), .ZN(n4292) );
  NAND2_X1 U5322 ( .A1(n4292), .A2(n4291), .ZN(n4293) );
  NAND2_X1 U5323 ( .A1(n4294), .A2(n4293), .ZN(n4374) );
  INV_X1 U5324 ( .A(n4374), .ZN(n4305) );
  INV_X1 U5325 ( .A(n4908), .ZN(n4295) );
  NAND2_X1 U5326 ( .A1(n5266), .A2(n4295), .ZN(n4298) );
  AOI21_X1 U5327 ( .B1(n4298), .B2(n4297), .A(n4296), .ZN(n4302) );
  NAND2_X1 U5328 ( .A1(n4300), .A2(n4299), .ZN(n4301) );
  AOI21_X1 U5329 ( .B1(n4322), .B2(n4302), .A(n4301), .ZN(n4304) );
  INV_X1 U5330 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6660) );
  NAND2_X1 U5331 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4434), .ZN(n6559) );
  OAI22_X1 U5332 ( .A1(n6435), .A2(n6481), .B1(n6660), .B2(n6559), .ZN(n4306)
         );
  NOR2_X1 U5333 ( .A1(n4474), .A2(n4306), .ZN(n5272) );
  INV_X1 U5334 ( .A(n5272), .ZN(n6569) );
  INV_X1 U5335 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6562) );
  NAND2_X1 U5336 ( .A1(n6562), .A2(n4306), .ZN(n4310) );
  INV_X1 U5337 ( .A(n6375), .ZN(n4517) );
  NOR2_X1 U5338 ( .A1(n4307), .A2(n4517), .ZN(n4308) );
  XNOR2_X1 U5339 ( .A(n4308), .B(n3502), .ZN(n5940) );
  NOR2_X1 U5340 ( .A1(n4290), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4309) );
  NAND2_X1 U5341 ( .A1(n5940), .A2(n4309), .ZN(n4432) );
  OAI22_X1 U5342 ( .A1(n6569), .A2(n3502), .B1(n4310), .B2(n4432), .ZN(U3455)
         );
  INV_X1 U5343 ( .A(n4312), .ZN(n4960) );
  AND3_X1 U5344 ( .A1(n4290), .A2(n4313), .A3(n4372), .ZN(n4314) );
  NAND2_X1 U5345 ( .A1(n4315), .A2(n4314), .ZN(n4407) );
  INV_X1 U5346 ( .A(n4407), .ZN(n5268) );
  INV_X1 U5347 ( .A(n5267), .ZN(n4320) );
  INV_X1 U5348 ( .A(n4316), .ZN(n4319) );
  INV_X1 U5349 ( .A(n4317), .ZN(n4318) );
  NAND2_X1 U5350 ( .A1(n4319), .A2(n4318), .ZN(n4323) );
  AOI22_X1 U5351 ( .A1(n5266), .A2(n4332), .B1(n4320), .B2(n4323), .ZN(n4321)
         );
  OAI21_X1 U5352 ( .B1(n4960), .B2(n5268), .A(n4321), .ZN(n6437) );
  INV_X1 U5353 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5242) );
  AOI22_X1 U5354 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5242), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n3546), .ZN(n4339) );
  NOR2_X1 U5355 ( .A1(n6477), .A2(n4340), .ZN(n4324) );
  AOI222_X1 U5356 ( .A1(n6437), .A2(n6564), .B1(n4339), .B2(n4324), .C1(n4323), 
        .C2(n6469), .ZN(n4326) );
  NAND2_X1 U5357 ( .A1(n5272), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4325) );
  OAI21_X1 U5358 ( .B1(n5272), .B2(n4326), .A(n4325), .ZN(U3460) );
  INV_X1 U5359 ( .A(n4327), .ZN(n4341) );
  AOI21_X1 U5360 ( .B1(n6469), .B2(n4341), .A(n5272), .ZN(n4345) );
  NAND2_X1 U5361 ( .A1(n4329), .A2(n4407), .ZN(n4338) );
  NAND2_X1 U5362 ( .A1(n4331), .A2(n4330), .ZN(n4421) );
  XNOR2_X1 U5363 ( .A(n4327), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4336)
         );
  XNOR2_X1 U5364 ( .A(n4332), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4333)
         );
  NAND2_X1 U5365 ( .A1(n5266), .A2(n4333), .ZN(n4334) );
  OAI21_X1 U5366 ( .B1(n4336), .B2(n4418), .A(n4334), .ZN(n4335) );
  AOI21_X1 U5367 ( .B1(n4421), .B2(n4336), .A(n4335), .ZN(n4337) );
  NAND2_X1 U5368 ( .A1(n4338), .A2(n4337), .ZN(n4424) );
  NOR3_X1 U5369 ( .A1(n6477), .A2(n4340), .A3(n4339), .ZN(n4343) );
  NOR3_X1 U5370 ( .A1(n6565), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n4341), 
        .ZN(n4342) );
  AOI211_X1 U5371 ( .C1(n4424), .C2(n6564), .A(n4343), .B(n4342), .ZN(n4344)
         );
  OAI22_X1 U5372 ( .A1(n4345), .A2(n3717), .B1(n5272), .B2(n4344), .ZN(U3459)
         );
  OAI21_X1 U5373 ( .B1(n4348), .B2(n4347), .A(n4346), .ZN(n4963) );
  OR2_X1 U5374 ( .A1(n4350), .A2(n4349), .ZN(n4351) );
  AND2_X1 U5375 ( .A1(n4352), .A2(n4351), .ZN(n4955) );
  INV_X1 U5376 ( .A(n4955), .ZN(n4368) );
  INV_X1 U5377 ( .A(n5988), .ZN(n5362) );
  AOI22_X1 U5378 ( .A1(n5977), .A2(n4368), .B1(EBX_REG_1__SCAN_IN), .B2(n5362), 
        .ZN(n4353) );
  OAI21_X1 U5379 ( .B1(n4963), .B2(n5984), .A(n4353), .ZN(U2858) );
  INV_X1 U5380 ( .A(n4354), .ZN(n4357) );
  OAI21_X1 U5381 ( .B1(n4357), .B2(n4356), .A(n4355), .ZN(n6143) );
  OAI222_X1 U5382 ( .A1(n6143), .A2(n5719), .B1(n5015), .B2(n5988), .C1(n5013), 
        .C2(n5983), .ZN(U2859) );
  OR2_X1 U5383 ( .A1(n4359), .A2(n4358), .ZN(n4360) );
  NAND2_X1 U5384 ( .A1(n4361), .A2(n4360), .ZN(n4382) );
  NOR2_X1 U5385 ( .A1(n4363), .A2(n4362), .ZN(n4364) );
  NAND2_X1 U5386 ( .A1(n6159), .A2(REIP_REG_1__SCAN_IN), .ZN(n4378) );
  OAI21_X1 U5387 ( .B1(n4364), .B2(n3546), .A(n4378), .ZN(n4367) );
  NOR3_X1 U5388 ( .A1(n5584), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4365), 
        .ZN(n4366) );
  AOI211_X1 U5389 ( .C1(n6161), .C2(n4368), .A(n4367), .B(n4366), .ZN(n4369)
         );
  OAI21_X1 U5390 ( .B1(n5636), .B2(n4382), .A(n4369), .ZN(U3017) );
  NOR2_X1 U5391 ( .A1(n4372), .A2(n4371), .ZN(n4373) );
  OAI21_X1 U5392 ( .B1(n4374), .B2(n4373), .A(n6473), .ZN(n4375) );
  NAND2_X1 U5393 ( .A1(n3164), .A2(n5288), .ZN(n4376) );
  NAND2_X2 U5394 ( .A1(n6011), .A2(n4376), .ZN(n6012) );
  INV_X1 U5395 ( .A(n4376), .ZN(n4377) );
  INV_X1 U5396 ( .A(DATAI_1_), .ZN(n6714) );
  INV_X1 U5397 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6079) );
  OAI222_X1 U5398 ( .A1(n4963), .A2(n6012), .B1(n6010), .B2(n6714), .C1(n6011), 
        .C2(n6079), .ZN(U2890) );
  INV_X1 U5399 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4958) );
  OAI21_X1 U5400 ( .B1(n5769), .B2(n4958), .A(n4378), .ZN(n4380) );
  NOR2_X1 U5401 ( .A1(n4963), .A2(n6142), .ZN(n4379) );
  AOI211_X1 U5402 ( .C1(n5763), .C2(n4958), .A(n4380), .B(n4379), .ZN(n4381)
         );
  OAI21_X1 U5403 ( .B1(n6135), .B2(n4382), .A(n4381), .ZN(U2985) );
  INV_X1 U5404 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6073) );
  AOI22_X1 U5405 ( .A1(n6031), .A2(UWORD_REG_14__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4383) );
  OAI21_X1 U5406 ( .B1(n6073), .B2(n4394), .A(n4383), .ZN(U2893) );
  INV_X1 U5407 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6058) );
  AOI22_X1 U5408 ( .A1(n6031), .A2(UWORD_REG_9__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4384) );
  OAI21_X1 U5409 ( .B1(n6058), .B2(n4394), .A(n4384), .ZN(U2898) );
  INV_X1 U5410 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6065) );
  AOI22_X1 U5411 ( .A1(n6031), .A2(UWORD_REG_11__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4385) );
  OAI21_X1 U5412 ( .B1(n6065), .B2(n4394), .A(n4385), .ZN(U2896) );
  INV_X1 U5413 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6050) );
  AOI22_X1 U5414 ( .A1(n6031), .A2(UWORD_REG_5__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4386) );
  OAI21_X1 U5415 ( .B1(n6050), .B2(n4394), .A(n4386), .ZN(U2902) );
  INV_X1 U5416 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6052) );
  AOI22_X1 U5417 ( .A1(n6031), .A2(UWORD_REG_6__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4387) );
  OAI21_X1 U5418 ( .B1(n6052), .B2(n4394), .A(n4387), .ZN(U2901) );
  INV_X1 U5419 ( .A(EAX_REG_20__SCAN_IN), .ZN(n6047) );
  AOI22_X1 U5420 ( .A1(n6031), .A2(UWORD_REG_4__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4388) );
  OAI21_X1 U5421 ( .B1(n6047), .B2(n4394), .A(n4388), .ZN(U2903) );
  INV_X1 U5422 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6054) );
  AOI22_X1 U5423 ( .A1(n6031), .A2(UWORD_REG_7__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4389) );
  OAI21_X1 U5424 ( .B1(n6054), .B2(n4394), .A(n4389), .ZN(U2900) );
  INV_X1 U5425 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6043) );
  AOI22_X1 U5426 ( .A1(n6031), .A2(UWORD_REG_2__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4390) );
  OAI21_X1 U5427 ( .B1(n6043), .B2(n4394), .A(n4390), .ZN(U2905) );
  INV_X1 U5428 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6045) );
  AOI22_X1 U5429 ( .A1(n6031), .A2(UWORD_REG_3__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4391) );
  OAI21_X1 U5430 ( .B1(n6045), .B2(n4394), .A(n4391), .ZN(U2904) );
  INV_X1 U5431 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6039) );
  AOI22_X1 U5432 ( .A1(n6031), .A2(UWORD_REG_0__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4392) );
  OAI21_X1 U5433 ( .B1(n6039), .B2(n4394), .A(n4392), .ZN(U2907) );
  INV_X1 U5434 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6041) );
  AOI22_X1 U5435 ( .A1(n6031), .A2(UWORD_REG_1__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4393) );
  OAI21_X1 U5436 ( .B1(n6041), .B2(n4394), .A(n4393), .ZN(U2906) );
  XNOR2_X1 U5437 ( .A(n4396), .B(n4395), .ZN(n4563) );
  OAI21_X1 U5438 ( .B1(n4884), .B2(n4397), .A(n5585), .ZN(n4737) );
  INV_X1 U5439 ( .A(n4737), .ZN(n6164) );
  NAND2_X1 U5440 ( .A1(n6162), .A2(n4398), .ZN(n6171) );
  NAND2_X1 U5441 ( .A1(n6164), .A2(n6171), .ZN(n4463) );
  AOI21_X1 U5442 ( .B1(n4397), .B2(n6169), .A(n6162), .ZN(n4889) );
  NOR2_X1 U5443 ( .A1(n4398), .A2(n4889), .ZN(n4461) );
  AOI22_X1 U5444 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4463), .B1(n4461), 
        .B2(n3335), .ZN(n4402) );
  INV_X1 U5445 ( .A(n4453), .ZN(n4399) );
  AOI21_X1 U5446 ( .B1(n4443), .B2(n4400), .A(n4399), .ZN(n5957) );
  INV_X1 U5447 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6510) );
  NOR2_X1 U5448 ( .A1(n6134), .A2(n6510), .ZN(n4558) );
  AOI21_X1 U5449 ( .B1(n6161), .B2(n5957), .A(n4558), .ZN(n4401) );
  OAI211_X1 U5450 ( .C1(n4563), .C2(n5636), .A(n4402), .B(n4401), .ZN(U3015)
         );
  OAI21_X1 U5451 ( .B1(n4447), .B2(n4404), .A(n4450), .ZN(n5966) );
  AOI22_X1 U5452 ( .A1(n5977), .A2(n5957), .B1(EBX_REG_3__SCAN_IN), .B2(n5362), 
        .ZN(n4405) );
  OAI21_X1 U5453 ( .B1(n5966), .B2(n5984), .A(n4405), .ZN(U2856) );
  NAND2_X1 U5454 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6660), .ZN(n4427) );
  INV_X1 U5455 ( .A(n4409), .ZN(n4426) );
  NAND2_X1 U5456 ( .A1(n6218), .A2(n4407), .ZN(n4423) );
  MUX2_X1 U5457 ( .A(n4408), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4327), 
        .Z(n4410) );
  NOR2_X1 U5458 ( .A1(n4410), .A2(n4409), .ZN(n4420) );
  AOI21_X1 U5459 ( .B1(n4327), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n4411), 
        .ZN(n4412) );
  NOR2_X1 U5460 ( .A1(n4413), .A2(n4412), .ZN(n6566) );
  AND2_X1 U5461 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4415) );
  INV_X1 U5462 ( .A(n4415), .ZN(n4414) );
  MUX2_X1 U5463 ( .A(n4415), .B(n4414), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4416) );
  NAND2_X1 U5464 ( .A1(n5266), .A2(n4416), .ZN(n4417) );
  OAI21_X1 U5465 ( .B1(n6566), .B2(n4418), .A(n4417), .ZN(n4419) );
  AOI21_X1 U5466 ( .B1(n4421), .B2(n4420), .A(n4419), .ZN(n4422) );
  NAND2_X1 U5467 ( .A1(n4423), .A2(n4422), .ZN(n6563) );
  MUX2_X1 U5468 ( .A(n6563), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6435), 
        .Z(n6445) );
  MUX2_X1 U5469 ( .A(n4424), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(n6435), 
        .Z(n6444) );
  NAND3_X1 U5470 ( .A1(n6445), .A2(n6444), .A3(n6477), .ZN(n4425) );
  OAI21_X1 U5471 ( .B1(n4427), .B2(n4426), .A(n4425), .ZN(n6460) );
  INV_X1 U5472 ( .A(n4428), .ZN(n4429) );
  NAND2_X1 U5473 ( .A1(n6460), .A2(n4429), .ZN(n4435) );
  MUX2_X1 U5474 ( .A(n6435), .B(n6660), .S(STATE2_REG_1__SCAN_IN), .Z(n4430)
         );
  NAND2_X1 U5475 ( .A1(n4430), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4431) );
  AND3_X1 U5476 ( .A1(n4435), .A2(n6660), .A3(n6458), .ZN(n4433) );
  NOR2_X1 U5477 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6582) );
  NAND3_X1 U5478 ( .A1(n4435), .A2(n6458), .A3(n4434), .ZN(n6475) );
  INV_X1 U5479 ( .A(n6475), .ZN(n4438) );
  INV_X1 U5480 ( .A(n6314), .ZN(n5269) );
  NAND2_X1 U5481 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6562), .ZN(n4667) );
  INV_X1 U5482 ( .A(n4667), .ZN(n4436) );
  OAI22_X1 U5483 ( .A1(n6304), .A2(n6374), .B1(n5269), .B2(n4436), .ZN(n4437)
         );
  OAI21_X1 U5484 ( .B1(n4438), .B2(n4437), .A(n6174), .ZN(n4439) );
  OAI21_X1 U5485 ( .B1(n6174), .B2(n6369), .A(n4439), .ZN(U3465) );
  NAND2_X1 U5486 ( .A1(n4441), .A2(n4440), .ZN(n4442) );
  AND2_X1 U5487 ( .A1(n4443), .A2(n4442), .ZN(n6160) );
  INV_X1 U5488 ( .A(n6160), .ZN(n4448) );
  INV_X1 U5489 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5008) );
  NOR2_X1 U5490 ( .A1(n4445), .A2(n4444), .ZN(n4446) );
  NOR2_X1 U5491 ( .A1(n4447), .A2(n4446), .ZN(n6127) );
  INV_X1 U5492 ( .A(n6127), .ZN(n5012) );
  OAI222_X1 U5493 ( .A1(n4448), .A2(n5983), .B1(n5988), .B2(n5008), .C1(n5012), 
        .C2(n5984), .ZN(U2857) );
  AND2_X1 U5494 ( .A1(n4450), .A2(n4449), .ZN(n4451) );
  OR2_X1 U5495 ( .A1(n4451), .A2(n4565), .ZN(n5944) );
  INV_X1 U5496 ( .A(n4567), .ZN(n4455) );
  NAND2_X1 U5497 ( .A1(n4453), .A2(n4452), .ZN(n4454) );
  NAND2_X1 U5498 ( .A1(n4455), .A2(n4454), .ZN(n5950) );
  INV_X1 U5499 ( .A(n5950), .ZN(n4456) );
  AOI22_X1 U5500 ( .A1(n4456), .A2(n5977), .B1(EBX_REG_4__SCAN_IN), .B2(n5362), 
        .ZN(n4457) );
  OAI21_X1 U5501 ( .B1(n5944), .B2(n5719), .A(n4457), .ZN(U2855) );
  INV_X1 U5502 ( .A(DATAI_2_), .ZN(n6618) );
  INV_X1 U5503 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6082) );
  OAI222_X1 U5504 ( .A1(n5012), .A2(n6012), .B1(n6010), .B2(n6618), .C1(n6011), 
        .C2(n6082), .ZN(U2889) );
  INV_X1 U5505 ( .A(DATAI_3_), .ZN(n6754) );
  INV_X1 U5506 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6085) );
  OAI222_X1 U5507 ( .A1(n5966), .A2(n6012), .B1(n6010), .B2(n6754), .C1(n6011), 
        .C2(n6085), .ZN(U2888) );
  XNOR2_X1 U5508 ( .A(n4458), .B(n4459), .ZN(n4809) );
  OAI211_X1 U5509 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4461), .B(n4460), .ZN(n4465) );
  INV_X1 U5510 ( .A(REIP_REG_4__SCAN_IN), .ZN(n5954) );
  OAI22_X1 U5511 ( .A1(n5631), .A2(n5950), .B1(n5954), .B2(n6134), .ZN(n4462)
         );
  AOI21_X1 U5512 ( .B1(n4463), .B2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4462), 
        .ZN(n4464) );
  OAI211_X1 U5513 ( .C1(n4809), .C2(n5636), .A(n4465), .B(n4464), .ZN(U3014)
         );
  NAND2_X1 U5514 ( .A1(n4329), .A2(n4312), .ZN(n6221) );
  INV_X1 U5515 ( .A(n6221), .ZN(n4766) );
  INV_X1 U5516 ( .A(n4466), .ZN(n4508) );
  AOI21_X1 U5517 ( .B1(n4812), .B2(n4766), .A(n4508), .ZN(n4472) );
  NAND2_X1 U5518 ( .A1(n3293), .A2(n5063), .ZN(n4468) );
  NOR2_X1 U5519 ( .A1(n4607), .A2(n4468), .ZN(n4477) );
  NAND2_X1 U5520 ( .A1(n6310), .A2(n6723), .ZN(n4969) );
  OAI21_X1 U5521 ( .B1(n4477), .B2(n6142), .A(n4969), .ZN(n4470) );
  AOI21_X1 U5522 ( .B1(n6369), .B2(STATE2_REG_3__SCAN_IN), .A(n4974), .ZN(
        n6261) );
  OAI21_X1 U5523 ( .B1(n4762), .B2(n6310), .A(n6261), .ZN(n4469) );
  AOI21_X1 U5524 ( .B1(n4472), .B2(n4470), .A(n4469), .ZN(n4515) );
  INV_X1 U5525 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4480) );
  NAND2_X1 U5526 ( .A1(DATAI_1_), .A2(n4763), .ZN(n6191) );
  INV_X1 U5527 ( .A(n4762), .ZN(n4471) );
  OAI22_X1 U5528 ( .A1(n4472), .A2(n6374), .B1(n4471), .B2(n6466), .ZN(n4509)
         );
  NOR2_X2 U5529 ( .A1(n4507), .A2(n4475), .ZN(n6385) );
  AOI22_X1 U5530 ( .A1(n6386), .A2(n4509), .B1(n4508), .B2(n6385), .ZN(n4479)
         );
  NAND2_X1 U5531 ( .A1(n4477), .A2(n5065), .ZN(n4645) );
  INV_X1 U5532 ( .A(DATAI_17_), .ZN(n4476) );
  OR2_X1 U5533 ( .A1(n6142), .A2(n4476), .ZN(n6329) );
  INV_X1 U5534 ( .A(n6329), .ZN(n6387) );
  INV_X1 U5535 ( .A(DATAI_25_), .ZN(n6748) );
  OR2_X1 U5536 ( .A1(n6142), .A2(n6748), .ZN(n6390) );
  INV_X1 U5537 ( .A(n6390), .ZN(n6230) );
  AOI22_X1 U5538 ( .A1(n4511), .A2(n6387), .B1(n4792), .B2(n6230), .ZN(n4478)
         );
  OAI211_X1 U5539 ( .C1(n4515), .C2(n4480), .A(n4479), .B(n4478), .ZN(U3141)
         );
  INV_X1 U5540 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4484) );
  NAND2_X1 U5541 ( .A1(DATAI_5_), .A2(n4763), .ZN(n6203) );
  NOR2_X2 U5542 ( .A1(n4507), .A2(n5289), .ZN(n6409) );
  AOI22_X1 U5543 ( .A1(n6410), .A2(n4509), .B1(n4508), .B2(n6409), .ZN(n4483)
         );
  INV_X1 U5544 ( .A(DATAI_21_), .ZN(n5738) );
  OR2_X1 U5545 ( .A1(n6142), .A2(n5738), .ZN(n6346) );
  INV_X1 U5546 ( .A(n6346), .ZN(n6411) );
  INV_X1 U5547 ( .A(DATAI_29_), .ZN(n4481) );
  OR2_X1 U5548 ( .A1(n6142), .A2(n4481), .ZN(n6414) );
  INV_X1 U5549 ( .A(n6414), .ZN(n6242) );
  AOI22_X1 U5550 ( .A1(n4511), .A2(n6411), .B1(n4792), .B2(n6242), .ZN(n4482)
         );
  OAI211_X1 U5551 ( .C1(n4515), .C2(n4484), .A(n4483), .B(n4482), .ZN(U3145)
         );
  INV_X1 U5552 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4488) );
  NAND2_X1 U5553 ( .A1(DATAI_6_), .A2(n4763), .ZN(n6206) );
  NOR2_X2 U5554 ( .A1(n4507), .A2(n3702), .ZN(n6415) );
  AOI22_X1 U5555 ( .A1(n6416), .A2(n4509), .B1(n4508), .B2(n6415), .ZN(n4487)
         );
  INV_X1 U5556 ( .A(DATAI_22_), .ZN(n4485) );
  OR2_X1 U5557 ( .A1(n6142), .A2(n4485), .ZN(n6351) );
  INV_X1 U5558 ( .A(n6351), .ZN(n6417) );
  INV_X1 U5559 ( .A(DATAI_30_), .ZN(n6755) );
  OR2_X1 U5560 ( .A1(n6142), .A2(n6755), .ZN(n6420) );
  INV_X1 U5561 ( .A(n6420), .ZN(n6245) );
  AOI22_X1 U5562 ( .A1(n4511), .A2(n6417), .B1(n4792), .B2(n6245), .ZN(n4486)
         );
  OAI211_X1 U5563 ( .C1(n4515), .C2(n4488), .A(n4487), .B(n4486), .ZN(U3146)
         );
  INV_X1 U5564 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4492) );
  NAND2_X1 U5565 ( .A1(DATAI_7_), .A2(n4763), .ZN(n6213) );
  NOR2_X2 U5566 ( .A1(n4507), .A2(n5310), .ZN(n6422) );
  AOI22_X1 U5567 ( .A1(n6424), .A2(n4509), .B1(n4508), .B2(n6422), .ZN(n4491)
         );
  INV_X1 U5568 ( .A(DATAI_23_), .ZN(n4489) );
  OR2_X1 U5569 ( .A1(n6142), .A2(n4489), .ZN(n6363) );
  INV_X1 U5570 ( .A(n6363), .ZN(n6426) );
  INV_X1 U5571 ( .A(DATAI_31_), .ZN(n6731) );
  OR2_X1 U5572 ( .A1(n6142), .A2(n6731), .ZN(n6431) );
  INV_X1 U5573 ( .A(n6431), .ZN(n6250) );
  AOI22_X1 U5574 ( .A1(n4511), .A2(n6426), .B1(n4792), .B2(n6250), .ZN(n4490)
         );
  OAI211_X1 U5575 ( .C1(n4515), .C2(n4492), .A(n4491), .B(n4490), .ZN(U3147)
         );
  INV_X1 U5576 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4496) );
  NAND2_X1 U5577 ( .A1(DATAI_4_), .A2(n4763), .ZN(n6200) );
  NOR2_X2 U5578 ( .A1(n4507), .A2(n4493), .ZN(n6403) );
  AOI22_X1 U5579 ( .A1(n6404), .A2(n4509), .B1(n4508), .B2(n6403), .ZN(n4495)
         );
  OR2_X1 U5580 ( .A1(n6142), .A2(n6747), .ZN(n6344) );
  INV_X1 U5581 ( .A(n6344), .ZN(n6405) );
  INV_X1 U5582 ( .A(DATAI_28_), .ZN(n6760) );
  OR2_X1 U5583 ( .A1(n6142), .A2(n6760), .ZN(n6408) );
  INV_X1 U5584 ( .A(n6408), .ZN(n6239) );
  AOI22_X1 U5585 ( .A1(n4511), .A2(n6405), .B1(n4792), .B2(n6239), .ZN(n4494)
         );
  OAI211_X1 U5586 ( .C1(n4515), .C2(n4496), .A(n4495), .B(n4494), .ZN(U3144)
         );
  INV_X1 U5587 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4500) );
  NAND2_X1 U5588 ( .A1(DATAI_2_), .A2(n4763), .ZN(n6194) );
  NOR2_X2 U5589 ( .A1(n4507), .A2(n4497), .ZN(n6391) );
  AOI22_X1 U5590 ( .A1(n6392), .A2(n4509), .B1(n4508), .B2(n6391), .ZN(n4499)
         );
  INV_X1 U5591 ( .A(DATAI_18_), .ZN(n5989) );
  OR2_X1 U5592 ( .A1(n6142), .A2(n5989), .ZN(n6334) );
  INV_X1 U5593 ( .A(n6334), .ZN(n6393) );
  INV_X1 U5594 ( .A(DATAI_26_), .ZN(n6742) );
  OR2_X1 U5595 ( .A1(n6142), .A2(n6742), .ZN(n6396) );
  INV_X1 U5596 ( .A(n6396), .ZN(n6233) );
  AOI22_X1 U5597 ( .A1(n4511), .A2(n6393), .B1(n4792), .B2(n6233), .ZN(n4498)
         );
  OAI211_X1 U5598 ( .C1(n4515), .C2(n4500), .A(n4499), .B(n4498), .ZN(U3142)
         );
  INV_X1 U5599 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4505) );
  NAND2_X1 U5600 ( .A1(DATAI_3_), .A2(n4763), .ZN(n6197) );
  NOR2_X2 U5601 ( .A1(n4507), .A2(n4501), .ZN(n6397) );
  AOI22_X1 U5602 ( .A1(n6398), .A2(n4509), .B1(n4508), .B2(n6397), .ZN(n4504)
         );
  INV_X1 U5603 ( .A(DATAI_19_), .ZN(n4502) );
  OR2_X1 U5604 ( .A1(n6142), .A2(n4502), .ZN(n6336) );
  INV_X1 U5605 ( .A(n6336), .ZN(n6399) );
  INV_X1 U5606 ( .A(DATAI_27_), .ZN(n6657) );
  OR2_X1 U5607 ( .A1(n6142), .A2(n6657), .ZN(n6402) );
  INV_X1 U5608 ( .A(n6402), .ZN(n6236) );
  AOI22_X1 U5609 ( .A1(n4511), .A2(n6399), .B1(n4792), .B2(n6236), .ZN(n4503)
         );
  OAI211_X1 U5610 ( .C1(n4515), .C2(n4505), .A(n4504), .B(n4503), .ZN(U3143)
         );
  INV_X1 U5611 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4514) );
  NAND2_X1 U5612 ( .A1(DATAI_0_), .A2(n4763), .ZN(n6188) );
  NOR2_X2 U5613 ( .A1(n4507), .A2(n4506), .ZN(n6370) );
  AOI22_X1 U5614 ( .A1(n6371), .A2(n4509), .B1(n4508), .B2(n6370), .ZN(n4513)
         );
  INV_X1 U5615 ( .A(DATAI_16_), .ZN(n5999) );
  OR2_X1 U5616 ( .A1(n6142), .A2(n5999), .ZN(n6324) );
  INV_X1 U5617 ( .A(n6324), .ZN(n6381) );
  INV_X1 U5618 ( .A(DATAI_24_), .ZN(n4510) );
  OR2_X1 U5619 ( .A1(n6142), .A2(n4510), .ZN(n6384) );
  INV_X1 U5620 ( .A(n6384), .ZN(n6227) );
  AOI22_X1 U5621 ( .A1(n4511), .A2(n6381), .B1(n4792), .B2(n6227), .ZN(n4512)
         );
  OAI211_X1 U5622 ( .C1(n4515), .C2(n4514), .A(n4513), .B(n4512), .ZN(U3140)
         );
  INV_X1 U5623 ( .A(DATAI_4_), .ZN(n6740) );
  INV_X1 U5624 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6088) );
  OAI222_X1 U5625 ( .A1(n5944), .A2(n6012), .B1(n6010), .B2(n6740), .C1(n6011), 
        .C2(n6088), .ZN(U2887) );
  AND2_X1 U5626 ( .A1(n4607), .A2(n5063), .ZN(n4516) );
  AND2_X1 U5627 ( .A1(n4329), .A2(n4960), .ZN(n6376) );
  AND2_X1 U5628 ( .A1(n6376), .A2(n4517), .ZN(n4569) );
  NAND2_X1 U5629 ( .A1(n4965), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4518) );
  OAI21_X1 U5630 ( .B1(n4966), .B2(n4518), .A(n6310), .ZN(n4575) );
  AOI211_X1 U5631 ( .C1(n6209), .C2(n4969), .A(n4569), .B(n4575), .ZN(n4520)
         );
  NAND2_X1 U5632 ( .A1(n6439), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4704) );
  OR2_X1 U5633 ( .A1(n4704), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4573)
         );
  NOR2_X1 U5634 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4573), .ZN(n4551)
         );
  NOR2_X1 U5635 ( .A1(n4522), .A2(n6466), .ZN(n5069) );
  INV_X1 U5636 ( .A(n5069), .ZN(n6378) );
  OR2_X1 U5637 ( .A1(n4972), .A2(n4843), .ZN(n4614) );
  AOI21_X1 U5638 ( .B1(n4614), .B2(STATE2_REG_2__SCAN_IN), .A(n4974), .ZN(
        n4611) );
  OAI211_X1 U5639 ( .C1(n6562), .C2(n4551), .A(n6378), .B(n4611), .ZN(n4519)
         );
  INV_X1 U5640 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4526) );
  NAND2_X1 U5641 ( .A1(n4965), .A2(n6304), .ZN(n4521) );
  NAND2_X1 U5642 ( .A1(n6376), .A2(n6310), .ZN(n6366) );
  AND2_X1 U5643 ( .A1(n4522), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4841) );
  INV_X1 U5644 ( .A(n4841), .ZN(n6365) );
  OAI22_X1 U5645 ( .A1(n6366), .A2(n6218), .B1(n4614), .B2(n6365), .ZN(n4552)
         );
  AOI22_X1 U5646 ( .A1(n6416), .A2(n4552), .B1(n6415), .B2(n4551), .ZN(n4523)
         );
  OAI21_X1 U5647 ( .B1(n6351), .B2(n4660), .A(n4523), .ZN(n4524) );
  AOI21_X1 U5648 ( .B1(n6245), .B2(n6209), .A(n4524), .ZN(n4525) );
  OAI21_X1 U5649 ( .B1(n4557), .B2(n4526), .A(n4525), .ZN(U3058) );
  INV_X1 U5650 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4530) );
  AOI22_X1 U5651 ( .A1(n6386), .A2(n4552), .B1(n6385), .B2(n4551), .ZN(n4527)
         );
  OAI21_X1 U5652 ( .B1(n6329), .B2(n4660), .A(n4527), .ZN(n4528) );
  AOI21_X1 U5653 ( .B1(n6230), .B2(n6209), .A(n4528), .ZN(n4529) );
  OAI21_X1 U5654 ( .B1(n4557), .B2(n4530), .A(n4529), .ZN(U3053) );
  INV_X1 U5655 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4534) );
  AOI22_X1 U5656 ( .A1(n6398), .A2(n4552), .B1(n6397), .B2(n4551), .ZN(n4531)
         );
  OAI21_X1 U5657 ( .B1(n6336), .B2(n4660), .A(n4531), .ZN(n4532) );
  AOI21_X1 U5658 ( .B1(n6236), .B2(n6209), .A(n4532), .ZN(n4533) );
  OAI21_X1 U5659 ( .B1(n4557), .B2(n4534), .A(n4533), .ZN(U3055) );
  INV_X1 U5660 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4538) );
  AOI22_X1 U5661 ( .A1(n6410), .A2(n4552), .B1(n6409), .B2(n4551), .ZN(n4535)
         );
  OAI21_X1 U5662 ( .B1(n6346), .B2(n4660), .A(n4535), .ZN(n4536) );
  AOI21_X1 U5663 ( .B1(n6242), .B2(n6209), .A(n4536), .ZN(n4537) );
  OAI21_X1 U5664 ( .B1(n4557), .B2(n4538), .A(n4537), .ZN(U3057) );
  INV_X1 U5665 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4542) );
  AOI22_X1 U5666 ( .A1(n6371), .A2(n4552), .B1(n6370), .B2(n4551), .ZN(n4539)
         );
  OAI21_X1 U5667 ( .B1(n6324), .B2(n4660), .A(n4539), .ZN(n4540) );
  AOI21_X1 U5668 ( .B1(n6227), .B2(n6209), .A(n4540), .ZN(n4541) );
  OAI21_X1 U5669 ( .B1(n4557), .B2(n4542), .A(n4541), .ZN(U3052) );
  INV_X1 U5670 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4546) );
  AOI22_X1 U5671 ( .A1(n6404), .A2(n4552), .B1(n6403), .B2(n4551), .ZN(n4543)
         );
  OAI21_X1 U5672 ( .B1(n6344), .B2(n4660), .A(n4543), .ZN(n4544) );
  AOI21_X1 U5673 ( .B1(n6239), .B2(n6209), .A(n4544), .ZN(n4545) );
  OAI21_X1 U5674 ( .B1(n4557), .B2(n4546), .A(n4545), .ZN(U3056) );
  INV_X1 U5675 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4550) );
  AOI22_X1 U5676 ( .A1(n6392), .A2(n4552), .B1(n6391), .B2(n4551), .ZN(n4547)
         );
  OAI21_X1 U5677 ( .B1(n6334), .B2(n4660), .A(n4547), .ZN(n4548) );
  AOI21_X1 U5678 ( .B1(n6233), .B2(n6209), .A(n4548), .ZN(n4549) );
  OAI21_X1 U5679 ( .B1(n4557), .B2(n4550), .A(n4549), .ZN(U3054) );
  INV_X1 U5680 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4556) );
  AOI22_X1 U5681 ( .A1(n6424), .A2(n4552), .B1(n6422), .B2(n4551), .ZN(n4553)
         );
  OAI21_X1 U5682 ( .B1(n6363), .B2(n4660), .A(n4553), .ZN(n4554) );
  AOI21_X1 U5683 ( .B1(n6250), .B2(n6209), .A(n4554), .ZN(n4555) );
  OAI21_X1 U5684 ( .B1(n4557), .B2(n4556), .A(n4555), .ZN(U3059) );
  INV_X1 U5685 ( .A(n5966), .ZN(n4561) );
  INV_X1 U5686 ( .A(n6142), .ZN(n6128) );
  AOI21_X1 U5687 ( .B1(n6139), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4558), 
        .ZN(n4559) );
  OAI21_X1 U5688 ( .B1(n5964), .B2(n6133), .A(n4559), .ZN(n4560) );
  AOI21_X1 U5689 ( .B1(n4561), .B2(n6128), .A(n4560), .ZN(n4562) );
  OAI21_X1 U5690 ( .B1(n4563), .B2(n6135), .A(n4562), .ZN(U2983) );
  OAI21_X1 U5691 ( .B1(n4565), .B2(n4564), .A(n4799), .ZN(n5929) );
  INV_X1 U5692 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6091) );
  OAI222_X1 U5693 ( .A1(n5929), .A2(n6012), .B1(n6010), .B2(n6048), .C1(n6011), 
        .C2(n6091), .ZN(U2886) );
  INV_X1 U5694 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4568) );
  OAI21_X1 U5695 ( .B1(n4567), .B2(n4566), .A(n4739), .ZN(n4749) );
  OAI222_X1 U5696 ( .A1(n5929), .A2(n5984), .B1(n4568), .B2(n5988), .C1(n5983), 
        .C2(n4749), .ZN(U2854) );
  INV_X1 U5697 ( .A(n4575), .ZN(n4572) );
  NOR2_X1 U5698 ( .A1(n6369), .A2(n4573), .ZN(n4658) );
  AOI21_X1 U5699 ( .B1(n4569), .B2(n6314), .A(n4658), .ZN(n4574) );
  INV_X1 U5700 ( .A(n6261), .ZN(n6316) );
  INV_X1 U5701 ( .A(n4573), .ZN(n4570) );
  NOR2_X1 U5702 ( .A1(n6310), .A2(n4570), .ZN(n4571) );
  AOI211_X2 U5703 ( .C1(n4572), .C2(n4574), .A(n6316), .B(n4571), .ZN(n4665)
         );
  INV_X1 U5704 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4579) );
  OAI22_X1 U5705 ( .A1(n4575), .A2(n4574), .B1(n4573), .B2(n6466), .ZN(n4662)
         );
  NOR3_X4 U5706 ( .A1(n4966), .A2(n5063), .A3(n6304), .ZN(n6251) );
  AOI22_X1 U5707 ( .A1(n6251), .A2(n6387), .B1(n6385), .B2(n4658), .ZN(n4576)
         );
  OAI21_X1 U5708 ( .B1(n6390), .B2(n4660), .A(n4576), .ZN(n4577) );
  AOI21_X1 U5709 ( .B1(n6386), .B2(n4662), .A(n4577), .ZN(n4578) );
  OAI21_X1 U5710 ( .B1(n4665), .B2(n4579), .A(n4578), .ZN(U3061) );
  INV_X1 U5711 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4583) );
  AOI22_X1 U5712 ( .A1(n6251), .A2(n6399), .B1(n6397), .B2(n4658), .ZN(n4580)
         );
  OAI21_X1 U5713 ( .B1(n6402), .B2(n4660), .A(n4580), .ZN(n4581) );
  AOI21_X1 U5714 ( .B1(n6398), .B2(n4662), .A(n4581), .ZN(n4582) );
  OAI21_X1 U5715 ( .B1(n4665), .B2(n4583), .A(n4582), .ZN(U3063) );
  INV_X1 U5716 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4587) );
  AOI22_X1 U5717 ( .A1(n6251), .A2(n6426), .B1(n6422), .B2(n4658), .ZN(n4584)
         );
  OAI21_X1 U5718 ( .B1(n6431), .B2(n4660), .A(n4584), .ZN(n4585) );
  AOI21_X1 U5719 ( .B1(n6424), .B2(n4662), .A(n4585), .ZN(n4586) );
  OAI21_X1 U5720 ( .B1(n4665), .B2(n4587), .A(n4586), .ZN(U3067) );
  INV_X1 U5721 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4591) );
  AOI22_X1 U5722 ( .A1(n6251), .A2(n6381), .B1(n6370), .B2(n4658), .ZN(n4588)
         );
  OAI21_X1 U5723 ( .B1(n6384), .B2(n4660), .A(n4588), .ZN(n4589) );
  AOI21_X1 U5724 ( .B1(n6371), .B2(n4662), .A(n4589), .ZN(n4590) );
  OAI21_X1 U5725 ( .B1(n4665), .B2(n4591), .A(n4590), .ZN(U3060) );
  INV_X1 U5726 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4595) );
  AOI22_X1 U5727 ( .A1(n6251), .A2(n6393), .B1(n6391), .B2(n4658), .ZN(n4592)
         );
  OAI21_X1 U5728 ( .B1(n6396), .B2(n4660), .A(n4592), .ZN(n4593) );
  AOI21_X1 U5729 ( .B1(n6392), .B2(n4662), .A(n4593), .ZN(n4594) );
  OAI21_X1 U5730 ( .B1(n4665), .B2(n4595), .A(n4594), .ZN(U3062) );
  INV_X1 U5731 ( .A(n6174), .ZN(n4606) );
  NOR2_X1 U5732 ( .A1(n4606), .A2(n6374), .ZN(n4666) );
  NAND2_X1 U5733 ( .A1(n5063), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6311) );
  XNOR2_X1 U5734 ( .A(n6179), .B(n6311), .ZN(n4596) );
  NAND2_X1 U5735 ( .A1(n4666), .A2(n4596), .ZN(n4598) );
  NAND3_X1 U5736 ( .A1(n6174), .A2(n4667), .A3(n4329), .ZN(n4597) );
  OAI211_X1 U5737 ( .C1(n3248), .C2(n6174), .A(n4598), .B(n4597), .ZN(U3463)
         );
  NOR2_X1 U5738 ( .A1(n4966), .A2(n6311), .ZN(n6256) );
  INV_X1 U5739 ( .A(n4969), .ZN(n4599) );
  AOI222_X1 U5740 ( .A1(n6218), .A2(n4667), .B1(n6310), .B2(n6256), .C1(n4599), 
        .C2(n3331), .ZN(n4605) );
  INV_X1 U5741 ( .A(n5064), .ZN(n6312) );
  NOR2_X1 U5742 ( .A1(n5063), .A2(n4600), .ZN(n4601) );
  NAND2_X1 U5743 ( .A1(n6179), .A2(n4601), .ZN(n4707) );
  INV_X1 U5744 ( .A(n4707), .ZN(n4602) );
  NAND2_X1 U5745 ( .A1(n4602), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4700) );
  NAND2_X1 U5746 ( .A1(n6312), .A2(n4700), .ZN(n6180) );
  NAND2_X1 U5747 ( .A1(n4666), .A2(n6180), .ZN(n4604) );
  NAND2_X1 U5748 ( .A1(n4606), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4603) );
  OAI211_X1 U5749 ( .C1(n4606), .C2(n4605), .A(n4604), .B(n4603), .ZN(U3462)
         );
  AND2_X1 U5750 ( .A1(n4607), .A2(n4965), .ZN(n4609) );
  NAND2_X1 U5751 ( .A1(n4609), .A2(n4608), .ZN(n4673) );
  NOR2_X2 U5752 ( .A1(n4673), .A2(n5065), .ZN(n4697) );
  NAND2_X1 U5753 ( .A1(n4645), .A2(n6310), .ZN(n4610) );
  OAI21_X1 U5754 ( .B1(n4697), .B2(n4610), .A(n4969), .ZN(n4613) );
  NOR2_X1 U5755 ( .A1(n4329), .A2(n4312), .ZN(n4968) );
  NAND2_X1 U5756 ( .A1(n6367), .A2(n4968), .ZN(n4671) );
  NAND3_X1 U5757 ( .A1(n6446), .A2(n3248), .A3(n6439), .ZN(n4677) );
  NOR2_X1 U5758 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4677), .ZN(n4642)
         );
  OAI211_X1 U5759 ( .C1(n6562), .C2(n4642), .A(n6365), .B(n4611), .ZN(n4612)
         );
  OAI22_X1 U5760 ( .A1(n4671), .A2(n6374), .B1(n6378), .B2(n4614), .ZN(n4643)
         );
  AOI22_X1 U5761 ( .A1(n6386), .A2(n4643), .B1(n6385), .B2(n4642), .ZN(n4615)
         );
  OAI21_X1 U5762 ( .B1(n6390), .B2(n4645), .A(n4615), .ZN(n4616) );
  AOI21_X1 U5763 ( .B1(n6387), .B2(n4697), .A(n4616), .ZN(n4617) );
  OAI21_X1 U5764 ( .B1(n4649), .B2(n3181), .A(n4617), .ZN(U3021) );
  AOI22_X1 U5765 ( .A1(n6371), .A2(n4643), .B1(n6370), .B2(n4642), .ZN(n4618)
         );
  OAI21_X1 U5766 ( .B1(n6384), .B2(n4645), .A(n4618), .ZN(n4619) );
  AOI21_X1 U5767 ( .B1(n6381), .B2(n4697), .A(n4619), .ZN(n4620) );
  OAI21_X1 U5768 ( .B1(n4649), .B2(n4621), .A(n4620), .ZN(U3020) );
  INV_X1 U5769 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4625) );
  AOI22_X1 U5770 ( .A1(n6416), .A2(n4643), .B1(n6415), .B2(n4642), .ZN(n4622)
         );
  OAI21_X1 U5771 ( .B1(n6420), .B2(n4645), .A(n4622), .ZN(n4623) );
  AOI21_X1 U5772 ( .B1(n6417), .B2(n4697), .A(n4623), .ZN(n4624) );
  OAI21_X1 U5773 ( .B1(n4649), .B2(n4625), .A(n4624), .ZN(U3026) );
  INV_X1 U5774 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4629) );
  AOI22_X1 U5775 ( .A1(n6398), .A2(n4643), .B1(n6397), .B2(n4642), .ZN(n4626)
         );
  OAI21_X1 U5776 ( .B1(n6402), .B2(n4645), .A(n4626), .ZN(n4627) );
  AOI21_X1 U5777 ( .B1(n6399), .B2(n4697), .A(n4627), .ZN(n4628) );
  OAI21_X1 U5778 ( .B1(n4649), .B2(n4629), .A(n4628), .ZN(U3023) );
  AOI22_X1 U5779 ( .A1(n6424), .A2(n4643), .B1(n6422), .B2(n4642), .ZN(n4630)
         );
  OAI21_X1 U5780 ( .B1(n6431), .B2(n4645), .A(n4630), .ZN(n4631) );
  AOI21_X1 U5781 ( .B1(n6426), .B2(n4697), .A(n4631), .ZN(n4632) );
  OAI21_X1 U5782 ( .B1(n4649), .B2(n4633), .A(n4632), .ZN(U3027) );
  INV_X1 U5783 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4637) );
  AOI22_X1 U5784 ( .A1(n6410), .A2(n4643), .B1(n6409), .B2(n4642), .ZN(n4634)
         );
  OAI21_X1 U5785 ( .B1(n6414), .B2(n4645), .A(n4634), .ZN(n4635) );
  AOI21_X1 U5786 ( .B1(n6411), .B2(n4697), .A(n4635), .ZN(n4636) );
  OAI21_X1 U5787 ( .B1(n4649), .B2(n4637), .A(n4636), .ZN(U3025) );
  AOI22_X1 U5788 ( .A1(n6404), .A2(n4643), .B1(n6403), .B2(n4642), .ZN(n4638)
         );
  OAI21_X1 U5789 ( .B1(n6408), .B2(n4645), .A(n4638), .ZN(n4639) );
  AOI21_X1 U5790 ( .B1(n6405), .B2(n4697), .A(n4639), .ZN(n4640) );
  OAI21_X1 U5791 ( .B1(n4649), .B2(n4641), .A(n4640), .ZN(U3024) );
  INV_X1 U5792 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4648) );
  AOI22_X1 U5793 ( .A1(n6392), .A2(n4643), .B1(n6391), .B2(n4642), .ZN(n4644)
         );
  OAI21_X1 U5794 ( .B1(n6396), .B2(n4645), .A(n4644), .ZN(n4646) );
  AOI21_X1 U5795 ( .B1(n6393), .B2(n4697), .A(n4646), .ZN(n4647) );
  OAI21_X1 U5796 ( .B1(n4649), .B2(n4648), .A(n4647), .ZN(U3022) );
  INV_X1 U5797 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4653) );
  AOI22_X1 U5798 ( .A1(n6251), .A2(n6405), .B1(n6403), .B2(n4658), .ZN(n4650)
         );
  OAI21_X1 U5799 ( .B1(n6408), .B2(n4660), .A(n4650), .ZN(n4651) );
  AOI21_X1 U5800 ( .B1(n6404), .B2(n4662), .A(n4651), .ZN(n4652) );
  OAI21_X1 U5801 ( .B1(n4665), .B2(n4653), .A(n4652), .ZN(U3064) );
  INV_X1 U5802 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4657) );
  AOI22_X1 U5803 ( .A1(n6251), .A2(n6417), .B1(n6415), .B2(n4658), .ZN(n4654)
         );
  OAI21_X1 U5804 ( .B1(n6420), .B2(n4660), .A(n4654), .ZN(n4655) );
  AOI21_X1 U5805 ( .B1(n6416), .B2(n4662), .A(n4655), .ZN(n4656) );
  OAI21_X1 U5806 ( .B1(n4665), .B2(n4657), .A(n4656), .ZN(U3066) );
  INV_X1 U5807 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4664) );
  AOI22_X1 U5808 ( .A1(n6251), .A2(n6411), .B1(n6409), .B2(n4658), .ZN(n4659)
         );
  OAI21_X1 U5809 ( .B1(n6414), .B2(n4660), .A(n4659), .ZN(n4661) );
  AOI21_X1 U5810 ( .B1(n6410), .B2(n4662), .A(n4661), .ZN(n4663) );
  OAI21_X1 U5811 ( .B1(n4665), .B2(n4664), .A(n4663), .ZN(U3065) );
  OAI211_X1 U5812 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n5063), .A(n4666), .B(
        n6311), .ZN(n4669) );
  NAND3_X1 U5813 ( .A1(n6174), .A2(n4312), .A3(n4667), .ZN(n4668) );
  OAI211_X1 U5814 ( .C1(n6174), .C2(n6439), .A(n4669), .B(n4668), .ZN(U3464)
         );
  INV_X1 U5815 ( .A(n4673), .ZN(n4670) );
  INV_X1 U5816 ( .A(n4671), .ZN(n4672) );
  NOR2_X1 U5817 ( .A1(n6369), .A2(n4677), .ZN(n4696) );
  AOI21_X1 U5818 ( .B1(n4672), .B2(n6314), .A(n4696), .ZN(n4679) );
  OR2_X1 U5819 ( .A1(n4673), .A2(n6723), .ZN(n4674) );
  NAND2_X1 U5820 ( .A1(n4674), .A2(n6310), .ZN(n4678) );
  INV_X1 U5821 ( .A(n4678), .ZN(n4675) );
  AOI22_X1 U5822 ( .A1(n4679), .A2(n4675), .B1(n6374), .B2(n4677), .ZN(n4676)
         );
  NAND2_X1 U5823 ( .A1(n6261), .A2(n4676), .ZN(n4695) );
  OAI22_X1 U5824 ( .A1(n4679), .A2(n4678), .B1(n6466), .B2(n4677), .ZN(n4694)
         );
  AOI22_X1 U5825 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4695), .B1(n6371), 
        .B2(n4694), .ZN(n4681) );
  AOI22_X1 U5826 ( .A1(n4697), .A2(n6227), .B1(n6370), .B2(n4696), .ZN(n4680)
         );
  OAI211_X1 U5827 ( .C1(n6324), .C2(n4878), .A(n4681), .B(n4680), .ZN(U3028)
         );
  AOI22_X1 U5828 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4695), .B1(n6410), 
        .B2(n4694), .ZN(n4683) );
  AOI22_X1 U5829 ( .A1(n4697), .A2(n6242), .B1(n6409), .B2(n4696), .ZN(n4682)
         );
  OAI211_X1 U5830 ( .C1(n6346), .C2(n4878), .A(n4683), .B(n4682), .ZN(U3033)
         );
  AOI22_X1 U5831 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4695), .B1(n6404), 
        .B2(n4694), .ZN(n4685) );
  AOI22_X1 U5832 ( .A1(n4697), .A2(n6239), .B1(n6403), .B2(n4696), .ZN(n4684)
         );
  OAI211_X1 U5833 ( .C1(n6344), .C2(n4878), .A(n4685), .B(n4684), .ZN(U3032)
         );
  AOI22_X1 U5834 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4695), .B1(n6416), 
        .B2(n4694), .ZN(n4687) );
  AOI22_X1 U5835 ( .A1(n4697), .A2(n6245), .B1(n6415), .B2(n4696), .ZN(n4686)
         );
  OAI211_X1 U5836 ( .C1(n6351), .C2(n4878), .A(n4687), .B(n4686), .ZN(U3034)
         );
  AOI22_X1 U5837 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4695), .B1(n6392), 
        .B2(n4694), .ZN(n4689) );
  AOI22_X1 U5838 ( .A1(n4697), .A2(n6233), .B1(n6391), .B2(n4696), .ZN(n4688)
         );
  OAI211_X1 U5839 ( .C1(n6334), .C2(n4878), .A(n4689), .B(n4688), .ZN(U3030)
         );
  AOI22_X1 U5840 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4695), .B1(n6386), 
        .B2(n4694), .ZN(n4691) );
  AOI22_X1 U5841 ( .A1(n4697), .A2(n6230), .B1(n6385), .B2(n4696), .ZN(n4690)
         );
  OAI211_X1 U5842 ( .C1(n6329), .C2(n4878), .A(n4691), .B(n4690), .ZN(U3029)
         );
  AOI22_X1 U5843 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4695), .B1(n6398), 
        .B2(n4694), .ZN(n4693) );
  AOI22_X1 U5844 ( .A1(n4697), .A2(n6236), .B1(n6397), .B2(n4696), .ZN(n4692)
         );
  OAI211_X1 U5845 ( .C1(n6336), .C2(n4878), .A(n4693), .B(n4692), .ZN(U3031)
         );
  AOI22_X1 U5846 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4695), .B1(n6424), 
        .B2(n4694), .ZN(n4699) );
  AOI22_X1 U5847 ( .A1(n4697), .A2(n6250), .B1(n6422), .B2(n4696), .ZN(n4698)
         );
  OAI211_X1 U5848 ( .C1(n6363), .C2(n4878), .A(n4699), .B(n4698), .ZN(U3035)
         );
  NOR2_X1 U5849 ( .A1(n6446), .A2(n4704), .ZN(n6368) );
  INV_X1 U5850 ( .A(n6368), .ZN(n4703) );
  AND2_X1 U5851 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6368), .ZN(n4729)
         );
  AOI21_X1 U5852 ( .B1(n4812), .B2(n6376), .A(n4729), .ZN(n4706) );
  NAND2_X1 U5853 ( .A1(n4706), .A2(n4700), .ZN(n4701) );
  NOR2_X1 U5854 ( .A1(n6374), .A2(n4701), .ZN(n4702) );
  AOI211_X2 U5855 ( .C1(n6374), .C2(n4703), .A(n4702), .B(n6316), .ZN(n4734)
         );
  INV_X1 U5856 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U5857 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4705) );
  OAI22_X1 U5858 ( .A1(n4706), .A2(n6374), .B1(n4705), .B2(n4704), .ZN(n4730)
         );
  AOI22_X1 U5859 ( .A1(n6424), .A2(n4730), .B1(n6422), .B2(n4729), .ZN(n4709)
         );
  AOI22_X1 U5860 ( .A1(n6250), .A2(n6425), .B1(n2995), .B2(n6426), .ZN(n4708)
         );
  OAI211_X1 U5861 ( .C1(n4734), .C2(n4710), .A(n4709), .B(n4708), .ZN(U3131)
         );
  INV_X1 U5862 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4713) );
  AOI22_X1 U5863 ( .A1(n6416), .A2(n4730), .B1(n6415), .B2(n4729), .ZN(n4712)
         );
  AOI22_X1 U5864 ( .A1(n6245), .A2(n6425), .B1(n2995), .B2(n6417), .ZN(n4711)
         );
  OAI211_X1 U5865 ( .C1(n4734), .C2(n4713), .A(n4712), .B(n4711), .ZN(U3130)
         );
  INV_X1 U5866 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4716) );
  AOI22_X1 U5867 ( .A1(n6404), .A2(n4730), .B1(n6403), .B2(n4729), .ZN(n4715)
         );
  AOI22_X1 U5868 ( .A1(n6239), .A2(n6425), .B1(n2995), .B2(n6405), .ZN(n4714)
         );
  OAI211_X1 U5869 ( .C1(n4734), .C2(n4716), .A(n4715), .B(n4714), .ZN(U3128)
         );
  INV_X1 U5870 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4719) );
  AOI22_X1 U5871 ( .A1(n6398), .A2(n4730), .B1(n6397), .B2(n4729), .ZN(n4718)
         );
  AOI22_X1 U5872 ( .A1(n6236), .A2(n6425), .B1(n2995), .B2(n6399), .ZN(n4717)
         );
  OAI211_X1 U5873 ( .C1(n4734), .C2(n4719), .A(n4718), .B(n4717), .ZN(U3127)
         );
  INV_X1 U5874 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4722) );
  AOI22_X1 U5875 ( .A1(n6392), .A2(n4730), .B1(n6391), .B2(n4729), .ZN(n4721)
         );
  AOI22_X1 U5876 ( .A1(n6233), .A2(n6425), .B1(n2995), .B2(n6393), .ZN(n4720)
         );
  OAI211_X1 U5877 ( .C1(n4734), .C2(n4722), .A(n4721), .B(n4720), .ZN(U3126)
         );
  INV_X1 U5878 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4725) );
  AOI22_X1 U5879 ( .A1(n6386), .A2(n4730), .B1(n6385), .B2(n4729), .ZN(n4724)
         );
  AOI22_X1 U5880 ( .A1(n6230), .A2(n6425), .B1(n2995), .B2(n6387), .ZN(n4723)
         );
  OAI211_X1 U5881 ( .C1(n4734), .C2(n4725), .A(n4724), .B(n4723), .ZN(U3125)
         );
  INV_X1 U5882 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4728) );
  AOI22_X1 U5883 ( .A1(n6371), .A2(n4730), .B1(n6370), .B2(n4729), .ZN(n4727)
         );
  AOI22_X1 U5884 ( .A1(n6227), .A2(n6425), .B1(n2995), .B2(n6381), .ZN(n4726)
         );
  OAI211_X1 U5885 ( .C1(n4734), .C2(n4728), .A(n4727), .B(n4726), .ZN(U3124)
         );
  INV_X1 U5886 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4733) );
  AOI22_X1 U5887 ( .A1(n6410), .A2(n4730), .B1(n6409), .B2(n4729), .ZN(n4732)
         );
  AOI22_X1 U5888 ( .A1(n6242), .A2(n6425), .B1(n2995), .B2(n6411), .ZN(n4731)
         );
  OAI211_X1 U5889 ( .C1(n4734), .C2(n4733), .A(n4732), .B(n4731), .ZN(U3129)
         );
  XNOR2_X1 U5890 ( .A(n4735), .B(n4736), .ZN(n4805) );
  NAND2_X1 U5891 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4746), .ZN(n4741)
         );
  AOI21_X1 U5892 ( .B1(n5214), .B2(n4741), .A(n4737), .ZN(n4755) );
  INV_X1 U5893 ( .A(n4755), .ZN(n4744) );
  NAND2_X1 U5894 ( .A1(n4739), .A2(n4738), .ZN(n4740) );
  NAND2_X1 U5895 ( .A1(n4891), .A2(n4740), .ZN(n4916) );
  INV_X1 U5896 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6515) );
  OAI22_X1 U5897 ( .A1(n5631), .A2(n4916), .B1(n6515), .B2(n6134), .ZN(n4743)
         );
  NOR3_X1 U5898 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4889), .A3(n4741), 
        .ZN(n4742) );
  AOI211_X1 U5899 ( .C1(INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n4744), .A(n4743), 
        .B(n4742), .ZN(n4745) );
  OAI21_X1 U5900 ( .B1(n5636), .B2(n4805), .A(n4745), .ZN(U3012) );
  AOI21_X1 U5901 ( .B1(n6162), .B2(n4746), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n4754) );
  XOR2_X1 U5902 ( .A(n4748), .B(n4747), .Z(n4756) );
  NAND2_X1 U5903 ( .A1(n4756), .A2(n6166), .ZN(n4753) );
  INV_X1 U5904 ( .A(n4749), .ZN(n5925) );
  AND2_X1 U5905 ( .A1(n6159), .A2(REIP_REG_5__SCAN_IN), .ZN(n4758) );
  AND3_X1 U5906 ( .A1(n6169), .A2(n3328), .A3(n4750), .ZN(n4751) );
  AOI211_X1 U5907 ( .C1(n6161), .C2(n5925), .A(n4758), .B(n4751), .ZN(n4752)
         );
  OAI211_X1 U5908 ( .C1(n4755), .C2(n4754), .A(n4753), .B(n4752), .ZN(U3013)
         );
  NAND2_X1 U5909 ( .A1(n4756), .A2(n6129), .ZN(n4760) );
  NOR2_X1 U5910 ( .A1(n6133), .A2(n5935), .ZN(n4757) );
  AOI211_X1 U5911 ( .C1(n6139), .C2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4758), 
        .B(n4757), .ZN(n4759) );
  OAI211_X1 U5912 ( .C1(n6142), .C2(n5929), .A(n4760), .B(n4759), .ZN(U2981)
         );
  OAI21_X1 U5913 ( .B1(n2995), .B2(n4792), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4761) );
  NAND3_X1 U5914 ( .A1(n6221), .A2(n6310), .A3(n4761), .ZN(n4765) );
  NAND2_X1 U5915 ( .A1(n6369), .A2(n4762), .ZN(n4768) );
  AOI21_X1 U5916 ( .B1(n4768), .B2(STATE2_REG_3__SCAN_IN), .A(n6446), .ZN(
        n4764) );
  OAI21_X1 U5917 ( .B1(n4843), .B2(n6466), .A(n4763), .ZN(n4840) );
  NOR2_X1 U5918 ( .A1(n5069), .A2(n4840), .ZN(n6225) );
  INV_X1 U5919 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4771) );
  NAND2_X1 U5920 ( .A1(n4766), .A2(n6310), .ZN(n6219) );
  INV_X1 U5921 ( .A(n4843), .ZN(n4973) );
  NOR2_X1 U5922 ( .A1(n4973), .A2(n6446), .ZN(n5068) );
  INV_X1 U5923 ( .A(n5068), .ZN(n4767) );
  OAI22_X1 U5924 ( .A1(n6367), .A2(n6219), .B1(n6365), .B2(n4767), .ZN(n4791)
         );
  INV_X1 U5925 ( .A(n4768), .ZN(n4790) );
  AOI22_X1 U5926 ( .A1(n6371), .A2(n4791), .B1(n6370), .B2(n4790), .ZN(n4770)
         );
  AOI22_X1 U5927 ( .A1(n2995), .A2(n6227), .B1(n4792), .B2(n6381), .ZN(n4769)
         );
  OAI211_X1 U5928 ( .C1(n4796), .C2(n4771), .A(n4770), .B(n4769), .ZN(U3132)
         );
  INV_X1 U5929 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4774) );
  AOI22_X1 U5930 ( .A1(n6392), .A2(n4791), .B1(n6391), .B2(n4790), .ZN(n4773)
         );
  AOI22_X1 U5931 ( .A1(n2995), .A2(n6233), .B1(n4792), .B2(n6393), .ZN(n4772)
         );
  OAI211_X1 U5932 ( .C1(n4796), .C2(n4774), .A(n4773), .B(n4772), .ZN(U3134)
         );
  INV_X1 U5933 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4777) );
  AOI22_X1 U5934 ( .A1(n6398), .A2(n4791), .B1(n6397), .B2(n4790), .ZN(n4776)
         );
  AOI22_X1 U5935 ( .A1(n2995), .A2(n6236), .B1(n4792), .B2(n6399), .ZN(n4775)
         );
  OAI211_X1 U5936 ( .C1(n4796), .C2(n4777), .A(n4776), .B(n4775), .ZN(U3135)
         );
  INV_X1 U5937 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4780) );
  AOI22_X1 U5938 ( .A1(n6386), .A2(n4791), .B1(n6385), .B2(n4790), .ZN(n4779)
         );
  AOI22_X1 U5939 ( .A1(n2995), .A2(n6230), .B1(n4792), .B2(n6387), .ZN(n4778)
         );
  OAI211_X1 U5940 ( .C1(n4796), .C2(n4780), .A(n4779), .B(n4778), .ZN(U3133)
         );
  INV_X1 U5941 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4783) );
  AOI22_X1 U5942 ( .A1(n6410), .A2(n4791), .B1(n6409), .B2(n4790), .ZN(n4782)
         );
  AOI22_X1 U5943 ( .A1(n2995), .A2(n6242), .B1(n4792), .B2(n6411), .ZN(n4781)
         );
  OAI211_X1 U5944 ( .C1(n4796), .C2(n4783), .A(n4782), .B(n4781), .ZN(U3137)
         );
  INV_X1 U5945 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4786) );
  AOI22_X1 U5946 ( .A1(n6416), .A2(n4791), .B1(n6415), .B2(n4790), .ZN(n4785)
         );
  AOI22_X1 U5947 ( .A1(n2995), .A2(n6245), .B1(n4792), .B2(n6417), .ZN(n4784)
         );
  OAI211_X1 U5948 ( .C1(n4796), .C2(n4786), .A(n4785), .B(n4784), .ZN(U3138)
         );
  INV_X1 U5949 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4789) );
  AOI22_X1 U5950 ( .A1(n6424), .A2(n4791), .B1(n6422), .B2(n4790), .ZN(n4788)
         );
  AOI22_X1 U5951 ( .A1(n2995), .A2(n6250), .B1(n4792), .B2(n6426), .ZN(n4787)
         );
  OAI211_X1 U5952 ( .C1(n4796), .C2(n4789), .A(n4788), .B(n4787), .ZN(U3139)
         );
  INV_X1 U5953 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4795) );
  AOI22_X1 U5954 ( .A1(n6404), .A2(n4791), .B1(n6403), .B2(n4790), .ZN(n4794)
         );
  AOI22_X1 U5955 ( .A1(n2995), .A2(n6239), .B1(n4792), .B2(n6405), .ZN(n4793)
         );
  OAI211_X1 U5956 ( .C1(n4796), .C2(n4795), .A(n4794), .B(n4793), .ZN(U3136)
         );
  INV_X1 U5957 ( .A(n4923), .ZN(n4798) );
  AOI21_X1 U5958 ( .B1(n4800), .B2(n4799), .A(n4798), .ZN(n4810) );
  INV_X1 U5959 ( .A(n4919), .ZN(n4802) );
  AOI22_X1 U5960 ( .A1(n6139), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .B1(n6159), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n4801) );
  OAI21_X1 U5961 ( .B1(n4802), .B2(n6133), .A(n4801), .ZN(n4803) );
  AOI21_X1 U5962 ( .B1(n4810), .B2(n6128), .A(n4803), .ZN(n4804) );
  OAI21_X1 U5963 ( .B1(n6135), .B2(n4805), .A(n4804), .ZN(U2980) );
  OAI22_X1 U5964 ( .A1(n5769), .A2(n5943), .B1(n6134), .B2(n5954), .ZN(n4807)
         );
  NOR2_X1 U5965 ( .A1(n5944), .A2(n6142), .ZN(n4806) );
  AOI211_X1 U5966 ( .C1(n5763), .C2(n5946), .A(n4807), .B(n4806), .ZN(n4808)
         );
  OAI21_X1 U5967 ( .B1(n6135), .B2(n4809), .A(n4808), .ZN(U2982) );
  INV_X1 U5968 ( .A(n4810), .ZN(n4921) );
  INV_X1 U5969 ( .A(DATAI_6_), .ZN(n6663) );
  INV_X1 U5970 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6094) );
  OAI222_X1 U5971 ( .A1(n4921), .A2(n6012), .B1(n6010), .B2(n6663), .C1(n6011), 
        .C2(n6094), .ZN(U2885) );
  INV_X1 U5972 ( .A(n4817), .ZN(n4811) );
  OAI21_X1 U5973 ( .B1(n4811), .B2(n6723), .A(n6310), .ZN(n4815) );
  NAND3_X1 U5974 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n3248), .A3(n6439), .ZN(n4971) );
  NOR2_X1 U5975 ( .A1(n6369), .A2(n4971), .ZN(n4834) );
  AOI21_X1 U5976 ( .B1(n4812), .B2(n4968), .A(n4834), .ZN(n4816) );
  INV_X1 U5977 ( .A(n4816), .ZN(n4814) );
  AOI21_X1 U5978 ( .B1(n6374), .B2(n4971), .A(n6316), .ZN(n4813) );
  OAI21_X1 U5979 ( .B1(n4815), .B2(n4814), .A(n4813), .ZN(n4833) );
  OAI22_X1 U5980 ( .A1(n4816), .A2(n4815), .B1(n6466), .B2(n4971), .ZN(n4832)
         );
  AOI22_X1 U5981 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4833), .B1(n6392), 
        .B2(n4832), .ZN(n4819) );
  AOI22_X1 U5982 ( .A1(n6299), .A2(n6233), .B1(n4834), .B2(n6391), .ZN(n4818)
         );
  OAI211_X1 U5983 ( .C1(n5099), .C2(n6334), .A(n4819), .B(n4818), .ZN(U3094)
         );
  AOI22_X1 U5984 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4833), .B1(n6371), 
        .B2(n4832), .ZN(n4821) );
  AOI22_X1 U5985 ( .A1(n6299), .A2(n6227), .B1(n6370), .B2(n4834), .ZN(n4820)
         );
  OAI211_X1 U5986 ( .C1(n6324), .C2(n5099), .A(n4821), .B(n4820), .ZN(U3092)
         );
  AOI22_X1 U5987 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4833), .B1(n6386), 
        .B2(n4832), .ZN(n4823) );
  AOI22_X1 U5988 ( .A1(n6299), .A2(n6230), .B1(n4834), .B2(n6385), .ZN(n4822)
         );
  OAI211_X1 U5989 ( .C1(n5099), .C2(n6329), .A(n4823), .B(n4822), .ZN(U3093)
         );
  AOI22_X1 U5990 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4833), .B1(n6424), 
        .B2(n4832), .ZN(n4825) );
  AOI22_X1 U5991 ( .A1(n6299), .A2(n6250), .B1(n4834), .B2(n6422), .ZN(n4824)
         );
  OAI211_X1 U5992 ( .C1(n5099), .C2(n6363), .A(n4825), .B(n4824), .ZN(U3099)
         );
  AOI22_X1 U5993 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4833), .B1(n6416), 
        .B2(n4832), .ZN(n4827) );
  AOI22_X1 U5994 ( .A1(n6299), .A2(n6245), .B1(n4834), .B2(n6415), .ZN(n4826)
         );
  OAI211_X1 U5995 ( .C1(n5099), .C2(n6351), .A(n4827), .B(n4826), .ZN(U3098)
         );
  AOI22_X1 U5996 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4833), .B1(n6398), 
        .B2(n4832), .ZN(n4829) );
  AOI22_X1 U5997 ( .A1(n6299), .A2(n6236), .B1(n4834), .B2(n6397), .ZN(n4828)
         );
  OAI211_X1 U5998 ( .C1(n5099), .C2(n6336), .A(n4829), .B(n4828), .ZN(U3095)
         );
  AOI22_X1 U5999 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4833), .B1(n6404), 
        .B2(n4832), .ZN(n4831) );
  AOI22_X1 U6000 ( .A1(n6299), .A2(n6239), .B1(n4834), .B2(n6403), .ZN(n4830)
         );
  OAI211_X1 U6001 ( .C1(n5099), .C2(n6344), .A(n4831), .B(n4830), .ZN(U3096)
         );
  AOI22_X1 U6002 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4833), .B1(n6410), 
        .B2(n4832), .ZN(n4836) );
  AOI22_X1 U6003 ( .A1(n6299), .A2(n6242), .B1(n4834), .B2(n6409), .ZN(n4835)
         );
  OAI211_X1 U6004 ( .C1(n5099), .C2(n6346), .A(n4836), .B(n4835), .ZN(U3097)
         );
  INV_X1 U6005 ( .A(n4878), .ZN(n4838) );
  OAI21_X1 U6006 ( .B1(n4838), .B2(n6208), .A(n4969), .ZN(n4839) );
  NOR2_X1 U6007 ( .A1(n4329), .A2(n4960), .ZN(n5067) );
  NAND2_X1 U6008 ( .A1(n6367), .A2(n5067), .ZN(n6175) );
  AOI21_X1 U6009 ( .B1(n4839), .B2(n6175), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4842) );
  NOR3_X1 U6010 ( .A1(n6439), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6178) );
  INV_X1 U6011 ( .A(n6178), .ZN(n6182) );
  NOR2_X1 U6012 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6182), .ZN(n4874)
         );
  NOR2_X1 U6013 ( .A1(n4841), .A2(n4840), .ZN(n5074) );
  OAI21_X1 U6014 ( .B1(n4842), .B2(n4874), .A(n5074), .ZN(n4880) );
  OR2_X1 U6015 ( .A1(n6175), .A2(n6374), .ZN(n4845) );
  AND2_X1 U6016 ( .A1(n4843), .A2(n6446), .ZN(n6216) );
  NAND2_X1 U6017 ( .A1(n5069), .A2(n6216), .ZN(n4844) );
  NAND2_X1 U6018 ( .A1(n4845), .A2(n4844), .ZN(n4875) );
  AOI22_X1 U6019 ( .A1(n6416), .A2(n4875), .B1(n6415), .B2(n4874), .ZN(n4847)
         );
  NAND2_X1 U6020 ( .A1(n6208), .A2(n6417), .ZN(n4846) );
  OAI211_X1 U6021 ( .C1(n4878), .C2(n6420), .A(n4847), .B(n4846), .ZN(n4848)
         );
  AOI21_X1 U6022 ( .B1(n4880), .B2(INSTQUEUE_REG_2__6__SCAN_IN), .A(n4848), 
        .ZN(n4849) );
  INV_X1 U6023 ( .A(n4849), .ZN(U3042) );
  AOI22_X1 U6024 ( .A1(n6404), .A2(n4875), .B1(n6403), .B2(n4874), .ZN(n4851)
         );
  NAND2_X1 U6025 ( .A1(n6208), .A2(n6405), .ZN(n4850) );
  OAI211_X1 U6026 ( .C1(n4878), .C2(n6408), .A(n4851), .B(n4850), .ZN(n4852)
         );
  AOI21_X1 U6027 ( .B1(n4880), .B2(INSTQUEUE_REG_2__4__SCAN_IN), .A(n4852), 
        .ZN(n4853) );
  INV_X1 U6028 ( .A(n4853), .ZN(U3040) );
  AOI22_X1 U6029 ( .A1(n6398), .A2(n4875), .B1(n6397), .B2(n4874), .ZN(n4855)
         );
  NAND2_X1 U6030 ( .A1(n6208), .A2(n6399), .ZN(n4854) );
  OAI211_X1 U6031 ( .C1(n4878), .C2(n6402), .A(n4855), .B(n4854), .ZN(n4856)
         );
  AOI21_X1 U6032 ( .B1(n4880), .B2(INSTQUEUE_REG_2__3__SCAN_IN), .A(n4856), 
        .ZN(n4857) );
  INV_X1 U6033 ( .A(n4857), .ZN(U3039) );
  AOI22_X1 U6034 ( .A1(n6424), .A2(n4875), .B1(n6422), .B2(n4874), .ZN(n4859)
         );
  NAND2_X1 U6035 ( .A1(n6208), .A2(n6426), .ZN(n4858) );
  OAI211_X1 U6036 ( .C1(n4878), .C2(n6431), .A(n4859), .B(n4858), .ZN(n4860)
         );
  AOI21_X1 U6037 ( .B1(n4880), .B2(INSTQUEUE_REG_2__7__SCAN_IN), .A(n4860), 
        .ZN(n4861) );
  INV_X1 U6038 ( .A(n4861), .ZN(U3043) );
  AOI22_X1 U6039 ( .A1(n6410), .A2(n4875), .B1(n6409), .B2(n4874), .ZN(n4863)
         );
  NAND2_X1 U6040 ( .A1(n6208), .A2(n6411), .ZN(n4862) );
  OAI211_X1 U6041 ( .C1(n4878), .C2(n6414), .A(n4863), .B(n4862), .ZN(n4864)
         );
  AOI21_X1 U6042 ( .B1(n4880), .B2(INSTQUEUE_REG_2__5__SCAN_IN), .A(n4864), 
        .ZN(n4865) );
  INV_X1 U6043 ( .A(n4865), .ZN(U3041) );
  AOI22_X1 U6044 ( .A1(n6386), .A2(n4875), .B1(n6385), .B2(n4874), .ZN(n4867)
         );
  NAND2_X1 U6045 ( .A1(n6208), .A2(n6387), .ZN(n4866) );
  OAI211_X1 U6046 ( .C1(n4878), .C2(n6390), .A(n4867), .B(n4866), .ZN(n4868)
         );
  AOI21_X1 U6047 ( .B1(n4880), .B2(INSTQUEUE_REG_2__1__SCAN_IN), .A(n4868), 
        .ZN(n4869) );
  INV_X1 U6048 ( .A(n4869), .ZN(U3037) );
  AOI22_X1 U6049 ( .A1(n6392), .A2(n4875), .B1(n6391), .B2(n4874), .ZN(n4871)
         );
  NAND2_X1 U6050 ( .A1(n6208), .A2(n6393), .ZN(n4870) );
  OAI211_X1 U6051 ( .C1(n4878), .C2(n6396), .A(n4871), .B(n4870), .ZN(n4872)
         );
  AOI21_X1 U6052 ( .B1(n4880), .B2(INSTQUEUE_REG_2__2__SCAN_IN), .A(n4872), 
        .ZN(n4873) );
  INV_X1 U6053 ( .A(n4873), .ZN(U3038) );
  AOI22_X1 U6054 ( .A1(n6371), .A2(n4875), .B1(n6370), .B2(n4874), .ZN(n4877)
         );
  NAND2_X1 U6055 ( .A1(n6208), .A2(n6381), .ZN(n4876) );
  OAI211_X1 U6056 ( .C1(n4878), .C2(n6384), .A(n4877), .B(n4876), .ZN(n4879)
         );
  AOI21_X1 U6057 ( .B1(n4880), .B2(INSTQUEUE_REG_2__0__SCAN_IN), .A(n4879), 
        .ZN(n4881) );
  INV_X1 U6058 ( .A(n4881), .ZN(U3036) );
  XNOR2_X1 U6059 ( .A(n2988), .B(n4883), .ZN(n4931) );
  INV_X1 U6060 ( .A(n4884), .ZN(n4886) );
  AOI22_X1 U6061 ( .A1(n6162), .A2(n4888), .B1(n4886), .B2(n4885), .ZN(n4887)
         );
  NAND2_X1 U6062 ( .A1(n5585), .A2(n4887), .ZN(n5134) );
  NOR2_X1 U6063 ( .A1(n4889), .A2(n4888), .ZN(n5050) );
  AOI22_X1 U6064 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n5134), .B1(n5050), 
        .B2(n3419), .ZN(n4894) );
  AND2_X1 U6065 ( .A1(n4891), .A2(n4890), .ZN(n4892) );
  NOR2_X1 U6066 ( .A1(n4936), .A2(n4892), .ZN(n5910) );
  INV_X1 U6067 ( .A(REIP_REG_7__SCAN_IN), .ZN(n5912) );
  NOR2_X1 U6068 ( .A1(n6134), .A2(n5912), .ZN(n4926) );
  AOI21_X1 U6069 ( .B1(n5910), .B2(n6161), .A(n4926), .ZN(n4893) );
  OAI211_X1 U6070 ( .C1(n4931), .C2(n5636), .A(n4894), .B(n4893), .ZN(U3011)
         );
  INV_X1 U6071 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4895) );
  OAI222_X1 U6072 ( .A1(n4916), .A2(n5983), .B1(n5988), .B2(n4895), .C1(n4921), 
        .C2(n5984), .ZN(U2853) );
  INV_X1 U6073 ( .A(n6582), .ZN(n6485) );
  NOR3_X1 U6074 ( .A1(n6476), .A2(n6562), .A3(n6485), .ZN(n6471) );
  INV_X1 U6075 ( .A(n6488), .ZN(n4896) );
  NOR3_X1 U6076 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n4896), .A3(n6477), .ZN(
        n6484) );
  OR3_X1 U6077 ( .A1(n6471), .A2(n6484), .A3(n6159), .ZN(n4897) );
  NOR2_X1 U6078 ( .A1(n5306), .A2(n6477), .ZN(n4900) );
  AND3_X1 U6079 ( .A1(n4902), .A2(n3106), .A3(n6723), .ZN(n4903) );
  INV_X1 U6080 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6513) );
  NAND3_X1 U6081 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5937) );
  NOR3_X1 U6082 ( .A1(n6513), .A2(n5954), .A3(n5937), .ZN(n5030) );
  OR2_X1 U6083 ( .A1(n5863), .A2(n5030), .ZN(n4904) );
  NAND2_X1 U6084 ( .A1(n4904), .A2(n5834), .ZN(n5933) );
  INV_X1 U6085 ( .A(n5933), .ZN(n4905) );
  NAND2_X1 U6086 ( .A1(n5924), .A2(n5030), .ZN(n5911) );
  AOI22_X1 U6087 ( .A1(REIP_REG_6__SCAN_IN), .A2(n4905), .B1(n5911), .B2(n6515), .ZN(n4918) );
  NOR2_X1 U6088 ( .A1(STATEBS16_REG_SCAN_IN), .A2(READY_N), .ZN(n4906) );
  NOR2_X1 U6089 ( .A1(n4954), .A2(n4906), .ZN(n4911) );
  INV_X1 U6090 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5353) );
  NOR2_X1 U6091 ( .A1(n2990), .A2(n5353), .ZN(n4907) );
  NOR2_X1 U6092 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n4908), .ZN(n6464) );
  INV_X1 U6093 ( .A(n6464), .ZN(n4909) );
  NAND2_X1 U6094 ( .A1(n6037), .A2(n4909), .ZN(n4910) );
  NOR2_X1 U6095 ( .A1(n4954), .A2(n4910), .ZN(n5317) );
  INV_X1 U6096 ( .A(n5317), .ZN(n4913) );
  NAND3_X1 U6097 ( .A1(n4911), .A2(n3106), .A3(n5353), .ZN(n4912) );
  AOI22_X1 U6098 ( .A1(EBX_REG_6__SCAN_IN), .A2(n5969), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n5913), .ZN(n4915) );
  NAND2_X1 U6099 ( .A1(n5834), .A2(n4914), .ZN(n5941) );
  OAI211_X1 U6100 ( .C1(n5962), .C2(n4916), .A(n4915), .B(n5941), .ZN(n4917)
         );
  AOI211_X1 U6101 ( .C1(n5945), .C2(n4919), .A(n4918), .B(n4917), .ZN(n4920)
         );
  OAI21_X1 U6102 ( .B1(n5916), .B2(n4921), .A(n4920), .ZN(U2821) );
  INV_X1 U6103 ( .A(n4941), .ZN(n4922) );
  AOI21_X1 U6104 ( .B1(n4924), .B2(n4923), .A(n4922), .ZN(n4929) );
  INV_X1 U6105 ( .A(n4929), .ZN(n5917) );
  AOI22_X1 U6106 ( .A1(n5910), .A2(n5977), .B1(EBX_REG_7__SCAN_IN), .B2(n5362), 
        .ZN(n4925) );
  OAI21_X1 U6107 ( .B1(n5917), .B2(n5984), .A(n4925), .ZN(U2852) );
  AOI21_X1 U6108 ( .B1(n6139), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n4926), 
        .ZN(n4927) );
  OAI21_X1 U6109 ( .B1(n5915), .B2(n6133), .A(n4927), .ZN(n4928) );
  AOI21_X1 U6110 ( .B1(n4929), .B2(n6128), .A(n4928), .ZN(n4930) );
  OAI21_X1 U6111 ( .B1(n6135), .B2(n4931), .A(n4930), .ZN(U2979) );
  INV_X1 U6112 ( .A(DATAI_7_), .ZN(n6719) );
  OAI222_X1 U6113 ( .A1(n5917), .A2(n6012), .B1(n6010), .B2(n6719), .C1(n6011), 
        .C2(n3755), .ZN(U2884) );
  XNOR2_X1 U6114 ( .A(n4932), .B(n4933), .ZN(n4949) );
  OAI211_X1 U6115 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n5050), .B(n4934), .ZN(n4940) );
  OR2_X1 U6116 ( .A1(n4936), .A2(n4935), .ZN(n4937) );
  NAND2_X1 U6117 ( .A1(n5027), .A2(n4937), .ZN(n5898) );
  INV_X1 U6118 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6518) );
  OAI22_X1 U6119 ( .A1(n5898), .A2(n5631), .B1(n6518), .B2(n6134), .ZN(n4938)
         );
  AOI21_X1 U6120 ( .B1(n5134), .B2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n4938), 
        .ZN(n4939) );
  OAI211_X1 U6121 ( .C1(n4949), .C2(n5636), .A(n4940), .B(n4939), .ZN(U3010)
         );
  AOI21_X1 U6122 ( .B1(n4942), .B2(n4941), .A(n5025), .ZN(n4964) );
  OAI22_X1 U6123 ( .A1(n5898), .A2(n5983), .B1(n5908), .B2(n5988), .ZN(n4943)
         );
  AOI21_X1 U6124 ( .B1(n4964), .B2(n4196), .A(n4943), .ZN(n4944) );
  INV_X1 U6125 ( .A(n4944), .ZN(U2851) );
  AOI22_X1 U6126 ( .A1(n6139), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6159), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n4945) );
  OAI21_X1 U6127 ( .B1(n4946), .B2(n6133), .A(n4945), .ZN(n4947) );
  AOI21_X1 U6128 ( .B1(n4964), .B2(n6128), .A(n4947), .ZN(n4948) );
  OAI21_X1 U6129 ( .B1(n6135), .B2(n4949), .A(n4948), .ZN(U2978) );
  NAND2_X1 U6130 ( .A1(n4951), .A2(n4950), .ZN(n4952) );
  NOR2_X1 U6131 ( .A1(n4954), .A2(n4953), .ZN(n5939) );
  INV_X1 U6132 ( .A(n5939), .ZN(n5960) );
  INV_X1 U6133 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6571) );
  OAI22_X1 U6134 ( .A1(n4955), .A2(n5962), .B1(n5834), .B2(n6571), .ZN(n4957)
         );
  NOR2_X1 U6135 ( .A1(n5959), .A2(n4958), .ZN(n4956) );
  AOI211_X1 U6136 ( .C1(n4958), .C2(n5945), .A(n4957), .B(n4956), .ZN(n4959)
         );
  OR2_X1 U6137 ( .A1(n5863), .A2(REIP_REG_1__SCAN_IN), .ZN(n5006) );
  OAI211_X1 U6138 ( .C1(n5960), .C2(n4960), .A(n4959), .B(n5006), .ZN(n4961)
         );
  AOI21_X1 U6139 ( .B1(EBX_REG_1__SCAN_IN), .B2(n5969), .A(n4961), .ZN(n4962)
         );
  OAI21_X1 U6140 ( .B1(n4963), .B2(n5965), .A(n4962), .ZN(U2826) );
  INV_X1 U6141 ( .A(n4964), .ZN(n5901) );
  INV_X1 U6142 ( .A(DATAI_8_), .ZN(n6757) );
  INV_X1 U6143 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6100) );
  OAI222_X1 U6144 ( .A1(n5901), .A2(n6012), .B1(n6010), .B2(n6757), .C1(n6011), 
        .C2(n6100), .ZN(U2883) );
  INV_X1 U6145 ( .A(n6299), .ZN(n4967) );
  NAND3_X1 U6146 ( .A1(n4967), .A2(n6310), .A3(n6303), .ZN(n4970) );
  AND2_X1 U6147 ( .A1(n4968), .A2(n6218), .ZN(n4977) );
  AOI21_X1 U6148 ( .B1(n4970), .B2(n4969), .A(n4977), .ZN(n4976) );
  NOR2_X1 U6149 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4971), .ZN(n6297)
         );
  NAND2_X1 U6150 ( .A1(n4973), .A2(n4972), .ZN(n6364) );
  AOI21_X1 U6151 ( .B1(n6364), .B2(STATE2_REG_2__SCAN_IN), .A(n4974), .ZN(
        n6377) );
  OAI211_X1 U6152 ( .C1(n6562), .C2(n6297), .A(n6365), .B(n6377), .ZN(n4975)
         );
  INV_X1 U6153 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4984) );
  NAND2_X1 U6154 ( .A1(n4977), .A2(n6310), .ZN(n4980) );
  INV_X1 U6155 ( .A(n6364), .ZN(n4978) );
  NAND2_X1 U6156 ( .A1(n4978), .A2(n5069), .ZN(n4979) );
  NAND2_X1 U6157 ( .A1(n4980), .A2(n4979), .ZN(n6298) );
  AOI22_X1 U6158 ( .A1(n6410), .A2(n6298), .B1(n6409), .B2(n6297), .ZN(n4981)
         );
  OAI21_X1 U6159 ( .B1(n6303), .B2(n6414), .A(n4981), .ZN(n4982) );
  AOI21_X1 U6160 ( .B1(n6299), .B2(n6411), .A(n4982), .ZN(n4983) );
  OAI21_X1 U6161 ( .B1(n5001), .B2(n4984), .A(n4983), .ZN(U3089) );
  INV_X1 U6162 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4988) );
  AOI22_X1 U6163 ( .A1(n6424), .A2(n6298), .B1(n6422), .B2(n6297), .ZN(n4985)
         );
  OAI21_X1 U6164 ( .B1(n6303), .B2(n6431), .A(n4985), .ZN(n4986) );
  AOI21_X1 U6165 ( .B1(n6299), .B2(n6426), .A(n4986), .ZN(n4987) );
  OAI21_X1 U6166 ( .B1(n5001), .B2(n4988), .A(n4987), .ZN(U3091) );
  INV_X1 U6167 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4992) );
  AOI22_X1 U6168 ( .A1(n6398), .A2(n6298), .B1(n6397), .B2(n6297), .ZN(n4989)
         );
  OAI21_X1 U6169 ( .B1(n6303), .B2(n6402), .A(n4989), .ZN(n4990) );
  AOI21_X1 U6170 ( .B1(n6299), .B2(n6399), .A(n4990), .ZN(n4991) );
  OAI21_X1 U6171 ( .B1(n5001), .B2(n4992), .A(n4991), .ZN(U3087) );
  INV_X1 U6172 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4996) );
  AOI22_X1 U6173 ( .A1(n6416), .A2(n6298), .B1(n6415), .B2(n6297), .ZN(n4993)
         );
  OAI21_X1 U6174 ( .B1(n6303), .B2(n6420), .A(n4993), .ZN(n4994) );
  AOI21_X1 U6175 ( .B1(n6299), .B2(n6417), .A(n4994), .ZN(n4995) );
  OAI21_X1 U6176 ( .B1(n5001), .B2(n4996), .A(n4995), .ZN(U3090) );
  INV_X1 U6177 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5000) );
  AOI22_X1 U6178 ( .A1(n6371), .A2(n6298), .B1(n6370), .B2(n6297), .ZN(n4997)
         );
  OAI21_X1 U6179 ( .B1(n6303), .B2(n6384), .A(n4997), .ZN(n4998) );
  AOI21_X1 U6180 ( .B1(n6381), .B2(n6299), .A(n4998), .ZN(n4999) );
  OAI21_X1 U6181 ( .B1(n5001), .B2(n5000), .A(n4999), .ZN(U3084) );
  INV_X1 U6182 ( .A(REIP_REG_2__SCAN_IN), .ZN(n5007) );
  NAND2_X1 U6183 ( .A1(n5007), .A2(REIP_REG_1__SCAN_IN), .ZN(n5005) );
  INV_X1 U6184 ( .A(n6132), .ZN(n5002) );
  AOI22_X1 U6185 ( .A1(n5913), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n5945), 
        .B2(n5002), .ZN(n5004) );
  NAND2_X1 U6186 ( .A1(n5939), .A2(n4329), .ZN(n5003) );
  OAI211_X1 U6187 ( .C1(n5863), .C2(n5005), .A(n5004), .B(n5003), .ZN(n5010)
         );
  AND2_X1 U6188 ( .A1(n5006), .A2(n5834), .ZN(n5956) );
  OAI22_X1 U6189 ( .A1(n5909), .A2(n5008), .B1(n5956), .B2(n5007), .ZN(n5009)
         );
  AOI211_X1 U6190 ( .C1(n5926), .C2(n6160), .A(n5010), .B(n5009), .ZN(n5011)
         );
  OAI21_X1 U6191 ( .B1(n5012), .B2(n5965), .A(n5011), .ZN(U2825) );
  INV_X1 U6192 ( .A(n5013), .ZN(n5014) );
  NAND2_X1 U6193 ( .A1(n5926), .A2(n5014), .ZN(n5019) );
  NAND2_X1 U6194 ( .A1(n5959), .A2(n5963), .ZN(n5017) );
  AND2_X1 U6195 ( .A1(n5863), .A2(n5834), .ZN(n5278) );
  OAI22_X1 U6196 ( .A1(n5278), .A2(n6576), .B1(n5909), .B2(n5015), .ZN(n5016)
         );
  AOI21_X1 U6197 ( .B1(n5017), .B2(PHYADDRPOINTER_REG_0__SCAN_IN), .A(n5016), 
        .ZN(n5018) );
  OAI211_X1 U6198 ( .C1(n5960), .C2(n5269), .A(n5019), .B(n5018), .ZN(n5020)
         );
  INV_X1 U6199 ( .A(n5020), .ZN(n5021) );
  OAI21_X1 U6200 ( .B1(n6143), .B2(n5965), .A(n5021), .ZN(U2827) );
  INV_X1 U6201 ( .A(n5060), .ZN(n5023) );
  OAI21_X1 U6202 ( .B1(n5025), .B2(n5024), .A(n5023), .ZN(n5058) );
  AOI21_X1 U6203 ( .B1(n5028), .B2(n5027), .A(n5026), .ZN(n6153) );
  AOI22_X1 U6204 ( .A1(n6153), .A2(n5977), .B1(EBX_REG_9__SCAN_IN), .B2(n5362), 
        .ZN(n5029) );
  OAI21_X1 U6205 ( .B1(n5058), .B2(n5719), .A(n5029), .ZN(U2850) );
  INV_X1 U6206 ( .A(n5041), .ZN(n5037) );
  NAND3_X1 U6207 ( .A1(n5030), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .ZN(n5032) );
  NOR2_X1 U6208 ( .A1(n6518), .A2(n5032), .ZN(n5109) );
  OR2_X1 U6209 ( .A1(n5863), .A2(n5109), .ZN(n5031) );
  AND2_X1 U6210 ( .A1(n5031), .A2(n5834), .ZN(n5887) );
  NOR2_X1 U6211 ( .A1(n5863), .A2(n5032), .ZN(n5905) );
  NAND2_X1 U6212 ( .A1(REIP_REG_8__SCAN_IN), .A2(n5905), .ZN(n5885) );
  INV_X1 U6213 ( .A(REIP_REG_9__SCAN_IN), .ZN(n5886) );
  AOI22_X1 U6214 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5887), .B1(n5885), .B2(n5886), .ZN(n5036) );
  AOI22_X1 U6215 ( .A1(EBX_REG_9__SCAN_IN), .A2(n5969), .B1(n5926), .B2(n6153), 
        .ZN(n5033) );
  OAI211_X1 U6216 ( .C1(n5959), .C2(n5034), .A(n5033), .B(n5941), .ZN(n5035)
         );
  AOI211_X1 U6217 ( .C1(n5945), .C2(n5037), .A(n5036), .B(n5035), .ZN(n5038)
         );
  OAI21_X1 U6218 ( .B1(n5058), .B2(n5916), .A(n5038), .ZN(U2818) );
  XNOR2_X1 U6219 ( .A(n3440), .B(n5053), .ZN(n5040) );
  XNOR2_X1 U6220 ( .A(n5039), .B(n5040), .ZN(n6155) );
  NAND2_X1 U6221 ( .A1(n6155), .A2(n6129), .ZN(n5044) );
  AND2_X1 U6222 ( .A1(n6159), .A2(REIP_REG_9__SCAN_IN), .ZN(n6152) );
  NOR2_X1 U6223 ( .A1(n6133), .A2(n5041), .ZN(n5042) );
  AOI211_X1 U6224 ( .C1(n6139), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6152), 
        .B(n5042), .ZN(n5043) );
  OAI211_X1 U6225 ( .C1(n6142), .C2(n5058), .A(n5044), .B(n5043), .ZN(U2977)
         );
  NAND2_X1 U6226 ( .A1(n3004), .A2(n5142), .ZN(n5046) );
  XNOR2_X1 U6227 ( .A(n5045), .B(n5046), .ZN(n5182) );
  INV_X1 U6228 ( .A(n5134), .ZN(n5047) );
  OAI21_X1 U6229 ( .B1(n5584), .B2(n5051), .A(n5047), .ZN(n6154) );
  INV_X1 U6230 ( .A(n5048), .ZN(n5114) );
  OAI21_X1 U6231 ( .B1(n5026), .B2(n5049), .A(n5114), .ZN(n5889) );
  OAI22_X1 U6232 ( .A1(n5889), .A2(n5631), .B1(n5177), .B2(n6134), .ZN(n5055)
         );
  NAND2_X1 U6233 ( .A1(n5051), .A2(n5050), .ZN(n6158) );
  AOI221_X1 U6234 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n5053), .C2(n5052), .A(n6158), 
        .ZN(n5054) );
  AOI211_X1 U6235 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n6154), .A(n5055), .B(n5054), .ZN(n5056) );
  OAI21_X1 U6236 ( .B1(n5182), .B2(n5636), .A(n5056), .ZN(U3008) );
  INV_X1 U6237 ( .A(DATAI_9_), .ZN(n5057) );
  INV_X1 U6238 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6103) );
  OAI222_X1 U6239 ( .A1(n5058), .A2(n6012), .B1(n6010), .B2(n5057), .C1(n6011), 
        .C2(n6103), .ZN(U2882) );
  NOR2_X1 U6240 ( .A1(n5060), .A2(n5059), .ZN(n5061) );
  OR2_X1 U6241 ( .A1(n5107), .A2(n5061), .ZN(n5894) );
  INV_X1 U6242 ( .A(n6010), .ZN(n5438) );
  AOI22_X1 U6243 ( .A1(n5438), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n6003), .ZN(n5062) );
  OAI21_X1 U6244 ( .B1(n5894), .B2(n6012), .A(n5062), .ZN(U2881) );
  NAND2_X1 U6245 ( .A1(n5064), .A2(n5063), .ZN(n6305) );
  NAND2_X1 U6246 ( .A1(n5099), .A2(n6357), .ZN(n5066) );
  AOI21_X1 U6247 ( .B1(n5066), .B2(STATEBS16_REG_SCAN_IN), .A(n6374), .ZN(
        n5072) );
  NAND3_X1 U6248 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n3248), .ZN(n6319) );
  NOR2_X1 U6249 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6319), .ZN(n5097)
         );
  INV_X1 U6250 ( .A(n6315), .ZN(n5071) );
  INV_X1 U6251 ( .A(n5097), .ZN(n5070) );
  AOI22_X1 U6252 ( .A1(n5072), .A2(n5071), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5070), .ZN(n5073) );
  OAI211_X1 U6253 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6466), .A(n5074), .B(n5073), .ZN(n5096) );
  AOI22_X1 U6254 ( .A1(n6415), .A2(n5097), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5096), .ZN(n5075) );
  OAI21_X1 U6255 ( .B1(n5099), .B2(n6420), .A(n5075), .ZN(n5076) );
  AOI21_X1 U6256 ( .B1(n6417), .B2(n5101), .A(n5076), .ZN(n5077) );
  OAI21_X1 U6257 ( .B1(n5103), .B2(n6206), .A(n5077), .ZN(U3106) );
  AOI22_X1 U6258 ( .A1(n6422), .A2(n5097), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5096), .ZN(n5078) );
  OAI21_X1 U6259 ( .B1(n5099), .B2(n6431), .A(n5078), .ZN(n5079) );
  AOI21_X1 U6260 ( .B1(n6426), .B2(n5101), .A(n5079), .ZN(n5080) );
  OAI21_X1 U6261 ( .B1(n5103), .B2(n6213), .A(n5080), .ZN(U3107) );
  AOI22_X1 U6262 ( .A1(n6397), .A2(n5097), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5096), .ZN(n5081) );
  OAI21_X1 U6263 ( .B1(n5099), .B2(n6402), .A(n5081), .ZN(n5082) );
  AOI21_X1 U6264 ( .B1(n6399), .B2(n5101), .A(n5082), .ZN(n5083) );
  OAI21_X1 U6265 ( .B1(n5103), .B2(n6197), .A(n5083), .ZN(U3103) );
  AOI22_X1 U6266 ( .A1(n6409), .A2(n5097), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5096), .ZN(n5084) );
  OAI21_X1 U6267 ( .B1(n5099), .B2(n6414), .A(n5084), .ZN(n5085) );
  AOI21_X1 U6268 ( .B1(n6411), .B2(n5101), .A(n5085), .ZN(n5086) );
  OAI21_X1 U6269 ( .B1(n5103), .B2(n6203), .A(n5086), .ZN(U3105) );
  AOI22_X1 U6270 ( .A1(n6370), .A2(n5097), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5096), .ZN(n5087) );
  OAI21_X1 U6271 ( .B1(n5099), .B2(n6384), .A(n5087), .ZN(n5088) );
  AOI21_X1 U6272 ( .B1(n6381), .B2(n5101), .A(n5088), .ZN(n5089) );
  OAI21_X1 U6273 ( .B1(n5103), .B2(n6188), .A(n5089), .ZN(U3100) );
  AOI22_X1 U6274 ( .A1(n6391), .A2(n5097), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5096), .ZN(n5090) );
  OAI21_X1 U6275 ( .B1(n5099), .B2(n6396), .A(n5090), .ZN(n5091) );
  AOI21_X1 U6276 ( .B1(n6393), .B2(n5101), .A(n5091), .ZN(n5092) );
  OAI21_X1 U6277 ( .B1(n5103), .B2(n6194), .A(n5092), .ZN(U3102) );
  AOI22_X1 U6278 ( .A1(n6385), .A2(n5097), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5096), .ZN(n5093) );
  OAI21_X1 U6279 ( .B1(n5099), .B2(n6390), .A(n5093), .ZN(n5094) );
  AOI21_X1 U6280 ( .B1(n6387), .B2(n5101), .A(n5094), .ZN(n5095) );
  OAI21_X1 U6281 ( .B1(n5103), .B2(n6191), .A(n5095), .ZN(U3101) );
  AOI22_X1 U6282 ( .A1(n6403), .A2(n5097), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5096), .ZN(n5098) );
  OAI21_X1 U6283 ( .B1(n5099), .B2(n6408), .A(n5098), .ZN(n5100) );
  AOI21_X1 U6284 ( .B1(n6405), .B2(n5101), .A(n5100), .ZN(n5102) );
  OAI21_X1 U6285 ( .B1(n5103), .B2(n6200), .A(n5102), .ZN(U3104) );
  INV_X1 U6286 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5104) );
  OAI222_X1 U6287 ( .A1(n5894), .A2(n5719), .B1(n5104), .B2(n5988), .C1(n5983), 
        .C2(n5889), .ZN(U2849) );
  OAI21_X1 U6288 ( .B1(n5107), .B2(n5106), .A(n5105), .ZN(n5150) );
  AOI22_X1 U6289 ( .A1(n5438), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n6003), .ZN(n5108) );
  OAI21_X1 U6290 ( .B1(n5150), .B2(n6012), .A(n5108), .ZN(U2880) );
  INV_X1 U6291 ( .A(n5146), .ZN(n5122) );
  INV_X1 U6292 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6522) );
  INV_X1 U6293 ( .A(n5834), .ZN(n5938) );
  NAND3_X1 U6294 ( .A1(n5109), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .ZN(n5116) );
  NOR2_X1 U6295 ( .A1(n6522), .A2(n5116), .ZN(n5875) );
  INV_X1 U6296 ( .A(n5875), .ZN(n5110) );
  INV_X1 U6297 ( .A(n5278), .ZN(n5936) );
  OAI21_X1 U6298 ( .B1(n5938), .B2(n5110), .A(n5936), .ZN(n5873) );
  OAI22_X1 U6299 ( .A1(n5909), .A2(n5111), .B1(n6522), .B2(n5873), .ZN(n5121)
         );
  INV_X1 U6300 ( .A(n5112), .ZN(n5115) );
  AOI21_X1 U6301 ( .B1(n5115), .B2(n5114), .A(n5113), .ZN(n6145) );
  NOR3_X1 U6302 ( .A1(n5863), .A2(REIP_REG_11__SCAN_IN), .A3(n5116), .ZN(n5117) );
  AOI211_X1 U6303 ( .C1(n5926), .C2(n6145), .A(n5921), .B(n5117), .ZN(n5118)
         );
  OAI21_X1 U6304 ( .B1(n5119), .B2(n5959), .A(n5118), .ZN(n5120) );
  AOI211_X1 U6305 ( .C1(n5945), .C2(n5122), .A(n5121), .B(n5120), .ZN(n5123)
         );
  OAI21_X1 U6306 ( .B1(n5150), .B2(n5916), .A(n5123), .ZN(U2816) );
  AOI22_X1 U6307 ( .A1(n6145), .A2(n5977), .B1(EBX_REG_11__SCAN_IN), .B2(n5362), .ZN(n5124) );
  OAI21_X1 U6308 ( .B1(n5150), .B2(n5984), .A(n5124), .ZN(U2848) );
  NAND2_X1 U6309 ( .A1(n5126), .A2(n5125), .ZN(n5129) );
  NAND2_X1 U6310 ( .A1(n2996), .A2(n5127), .ZN(n5128) );
  XNOR2_X1 U6311 ( .A(n5129), .B(n5128), .ZN(n5512) );
  AND2_X1 U6312 ( .A1(n5417), .A2(n5130), .ZN(n5131) );
  NOR2_X1 U6313 ( .A1(n5407), .A2(n5131), .ZN(n5976) );
  INV_X1 U6314 ( .A(n5976), .ZN(n5132) );
  NAND2_X1 U6315 ( .A1(n6159), .A2(REIP_REG_15__SCAN_IN), .ZN(n5508) );
  OAI21_X1 U6316 ( .B1(n5132), .B2(n5631), .A(n5508), .ZN(n5139) );
  NAND2_X1 U6317 ( .A1(n5585), .A2(n5584), .ZN(n5133) );
  OAI21_X1 U6318 ( .B1(n5135), .B2(n5134), .A(n5133), .ZN(n6150) );
  INV_X1 U6319 ( .A(n6150), .ZN(n5136) );
  AOI21_X1 U6320 ( .B1(n5214), .B2(n5137), .A(n5136), .ZN(n5621) );
  NOR2_X1 U6321 ( .A1(n5621), .A2(n5613), .ZN(n5138) );
  AOI211_X1 U6322 ( .C1(n5611), .C2(n5613), .A(n5139), .B(n5138), .ZN(n5140)
         );
  OAI21_X1 U6323 ( .B1(n5512), .B2(n5636), .A(n5140), .ZN(U3003) );
  NAND2_X1 U6324 ( .A1(n5152), .A2(n5142), .ZN(n5145) );
  NAND2_X1 U6325 ( .A1(n5143), .A2(n5153), .ZN(n5144) );
  XNOR2_X1 U6326 ( .A(n5145), .B(n5144), .ZN(n6147) );
  NAND2_X1 U6327 ( .A1(n6147), .A2(n6129), .ZN(n5149) );
  AND2_X1 U6328 ( .A1(n6159), .A2(REIP_REG_11__SCAN_IN), .ZN(n6144) );
  NOR2_X1 U6329 ( .A1(n6133), .A2(n5146), .ZN(n5147) );
  AOI211_X1 U6330 ( .C1(n6139), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6144), 
        .B(n5147), .ZN(n5148) );
  OAI211_X1 U6331 ( .C1(n6142), .C2(n5150), .A(n5149), .B(n5148), .ZN(U2975)
         );
  NAND2_X1 U6332 ( .A1(n5152), .A2(n5151), .ZN(n5154) );
  INV_X1 U6333 ( .A(n5526), .ZN(n5155) );
  NOR2_X1 U6334 ( .A1(n5524), .A2(n5155), .ZN(n5156) );
  XNOR2_X1 U6335 ( .A(n5525), .B(n5156), .ZN(n5176) );
  NOR2_X1 U6336 ( .A1(n5791), .A2(n6151), .ZN(n5161) );
  OR2_X1 U6337 ( .A1(n5113), .A2(n5158), .ZN(n5159) );
  NAND2_X1 U6338 ( .A1(n5157), .A2(n5159), .ZN(n5874) );
  INV_X1 U6339 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6524) );
  OAI22_X1 U6340 ( .A1(n5874), .A2(n5631), .B1(n6524), .B2(n6134), .ZN(n5160)
         );
  AOI21_X1 U6341 ( .B1(n5161), .B2(n3439), .A(n5160), .ZN(n5166) );
  OAI221_X1 U6342 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n5163), .C1(
        INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n5162), .A(n6150), .ZN(n5164) );
  NAND2_X1 U6343 ( .A1(n5164), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5165) );
  OAI211_X1 U6344 ( .C1(n5176), .C2(n5636), .A(n5166), .B(n5165), .ZN(U3006)
         );
  AOI21_X1 U6345 ( .B1(n5168), .B2(n5105), .A(n5167), .ZN(n5882) );
  INV_X1 U6346 ( .A(n5882), .ZN(n5171) );
  INV_X1 U6347 ( .A(DATAI_12_), .ZN(n6066) );
  OAI222_X1 U6348 ( .A1(n5171), .A2(n6012), .B1(n6011), .B2(n5169), .C1(n6066), 
        .C2(n6010), .ZN(U2879) );
  INV_X1 U6349 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5170) );
  OAI222_X1 U6350 ( .A1(n5171), .A2(n5984), .B1(n5170), .B2(n5988), .C1(n5983), 
        .C2(n5874), .ZN(U2847) );
  INV_X1 U6351 ( .A(n5880), .ZN(n5173) );
  AOI22_X1 U6352 ( .A1(n6139), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n6159), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n5172) );
  OAI21_X1 U6353 ( .B1(n5173), .B2(n6133), .A(n5172), .ZN(n5174) );
  AOI21_X1 U6354 ( .B1(n5882), .B2(n6128), .A(n5174), .ZN(n5175) );
  OAI21_X1 U6355 ( .B1(n5176), .B2(n6135), .A(n5175), .ZN(U2974) );
  INV_X1 U6356 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5178) );
  INV_X1 U6357 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5177) );
  OAI22_X1 U6358 ( .A1(n5769), .A2(n5178), .B1(n6134), .B2(n5177), .ZN(n5180)
         );
  NOR2_X1 U6359 ( .A1(n5894), .A2(n6142), .ZN(n5179) );
  AOI211_X1 U6360 ( .C1(n5763), .C2(n5892), .A(n5180), .B(n5179), .ZN(n5181)
         );
  OAI21_X1 U6361 ( .B1(n6135), .B2(n5182), .A(n5181), .ZN(U2976) );
  INV_X1 U6362 ( .A(n5183), .ZN(n5186) );
  INV_X1 U6363 ( .A(n5200), .ZN(n5185) );
  AOI21_X1 U6364 ( .B1(n5186), .B2(n5185), .A(n5184), .ZN(n5285) );
  NOR3_X1 U6365 ( .A1(n5206), .A2(n5188), .A3(n5187), .ZN(n5192) );
  OAI21_X1 U6366 ( .B1(n5196), .B2(n5190), .A(n5189), .ZN(n5191) );
  AOI211_X1 U6367 ( .C1(n5285), .C2(n6161), .A(n5192), .B(n5191), .ZN(n5193)
         );
  OAI21_X1 U6368 ( .B1(n5194), .B2(n5636), .A(n5193), .ZN(U2990) );
  NAND2_X1 U6369 ( .A1(n5195), .A2(n6166), .ZN(n5205) );
  INV_X1 U6370 ( .A(n5196), .ZN(n5203) );
  NOR2_X1 U6371 ( .A1(n5197), .A2(n5198), .ZN(n5199) );
  OR2_X1 U6372 ( .A1(n5200), .A2(n5199), .ZN(n5718) );
  NOR2_X1 U6373 ( .A1(n5718), .A2(n5631), .ZN(n5201) );
  AOI211_X1 U6374 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5203), .A(n5202), .B(n5201), .ZN(n5204) );
  OAI211_X1 U6375 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5206), .A(n5205), .B(n5204), .ZN(U2991) );
  NOR3_X1 U6376 ( .A1(n5207), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6377 ( .A1(n5208), .A2(n5227), .ZN(n5209) );
  INV_X1 U6378 ( .A(n5211), .ZN(n5212) );
  INV_X1 U6379 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5226) );
  XNOR2_X1 U6380 ( .A(n5212), .B(n5226), .ZN(n5225) );
  INV_X1 U6381 ( .A(n5333), .ZN(n5218) );
  NAND2_X1 U6382 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5240) );
  AOI21_X1 U6383 ( .B1(n5240), .B2(n5214), .A(n5213), .ZN(n5243) );
  INV_X1 U6384 ( .A(n5241), .ZN(n5215) );
  NAND3_X1 U6385 ( .A1(n5215), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5226), .ZN(n5216) );
  NAND2_X1 U6386 ( .A1(n6159), .A2(REIP_REG_30__SCAN_IN), .ZN(n5220) );
  OAI211_X1 U6387 ( .C1(n5243), .C2(n5226), .A(n5216), .B(n5220), .ZN(n5217)
         );
  AOI21_X1 U6388 ( .B1(n5218), .B2(n6161), .A(n5217), .ZN(n5219) );
  OAI21_X1 U6389 ( .B1(n5225), .B2(n5636), .A(n5219), .ZN(U2988) );
  NAND2_X1 U6390 ( .A1(n5763), .A2(n5326), .ZN(n5221) );
  OAI211_X1 U6391 ( .C1(n5769), .C2(n5222), .A(n5221), .B(n5220), .ZN(n5223)
         );
  AOI21_X1 U6392 ( .B1(n5325), .B2(n6128), .A(n5223), .ZN(n5224) );
  OAI21_X1 U6393 ( .B1(n5225), .B2(n6135), .A(n5224), .ZN(U2956) );
  NAND2_X1 U6394 ( .A1(n5227), .A2(n5226), .ZN(n5228) );
  OAI22_X1 U6395 ( .A1(n5229), .A2(n5240), .B1(n2987), .B2(n5228), .ZN(n5230)
         );
  XNOR2_X1 U6396 ( .A(n5230), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5309)
         );
  NAND2_X1 U6397 ( .A1(n5232), .A2(n5231), .ZN(n5235) );
  NAND2_X1 U6398 ( .A1(n5235), .A2(n5234), .ZN(n5239) );
  OAI22_X1 U6399 ( .A1(n5236), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n2990), .ZN(n5237) );
  NOR3_X1 U6400 ( .A1(n5241), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5240), 
        .ZN(n5245) );
  NAND2_X1 U6401 ( .A1(n6159), .A2(REIP_REG_31__SCAN_IN), .ZN(n5305) );
  OAI21_X1 U6402 ( .B1(n5243), .B2(n5242), .A(n5305), .ZN(n5244) );
  AOI21_X1 U6403 ( .B1(n5352), .B2(n6161), .A(n5246), .ZN(n5247) );
  OAI21_X1 U6404 ( .B1(n5309), .B2(n5636), .A(n5247), .ZN(U2987) );
  NOR2_X1 U6405 ( .A1(n5769), .A2(n5249), .ZN(n5250) );
  AOI211_X1 U6406 ( .C1(n5763), .C2(n5683), .A(n5251), .B(n5250), .ZN(n5258)
         );
  NAND2_X1 U6407 ( .A1(n5419), .A2(n5253), .ZN(n5379) );
  NAND2_X1 U6408 ( .A1(n5419), .A2(n5254), .ZN(n5474) );
  INV_X1 U6409 ( .A(n5474), .ZN(n5255) );
  AOI21_X1 U6410 ( .B1(n5256), .B2(n5379), .A(n5255), .ZN(n5374) );
  NAND2_X1 U6411 ( .A1(n5374), .A2(n6128), .ZN(n5257) );
  OAI211_X1 U6412 ( .C1(n5248), .C2(n6135), .A(n5258), .B(n5257), .ZN(U2964)
         );
  AOI21_X1 U6413 ( .B1(n5260), .B2(n5259), .A(n5298), .ZN(n5355) );
  AOI21_X1 U6414 ( .B1(n6139), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5261), 
        .ZN(n5262) );
  OAI21_X1 U6415 ( .B1(n5334), .B2(n6133), .A(n5262), .ZN(n5263) );
  AOI21_X1 U6416 ( .B1(n5355), .B2(n6128), .A(n5263), .ZN(n5264) );
  OAI21_X1 U6417 ( .B1(n5265), .B2(n6135), .A(n5264), .ZN(U2957) );
  AOI21_X1 U6418 ( .B1(n5266), .B2(n6564), .A(n5272), .ZN(n5273) );
  OAI22_X1 U6419 ( .A1(n5269), .A2(n5268), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5267), .ZN(n6432) );
  OAI22_X1 U6420 ( .A1(n6565), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n6477), .ZN(n5270) );
  AOI21_X1 U6421 ( .B1(n6432), .B2(n6564), .A(n5270), .ZN(n5271) );
  OAI22_X1 U6422 ( .A1(n5273), .A2(n3710), .B1(n5272), .B2(n5271), .ZN(U3461)
         );
  AOI22_X1 U6423 ( .A1(n5285), .A2(n5977), .B1(EBX_REG_28__SCAN_IN), .B2(n5362), .ZN(n5274) );
  OAI21_X1 U6424 ( .B1(n5293), .B2(n5984), .A(n5274), .ZN(U2831) );
  INV_X1 U6425 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6666) );
  INV_X1 U6426 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6538) );
  INV_X1 U6427 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6536) );
  INV_X1 U6428 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6533) );
  INV_X1 U6429 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6527) );
  NAND3_X1 U6430 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .A3(
        n5875), .ZN(n5855) );
  NOR2_X1 U6431 ( .A1(n6527), .A2(n5855), .ZN(n5823) );
  NAND4_X1 U6432 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .A4(n5823), .ZN(n5704) );
  NOR2_X1 U6433 ( .A1(n6533), .A2(n5704), .ZN(n5705) );
  NAND2_X1 U6434 ( .A1(REIP_REG_19__SCAN_IN), .A2(n5705), .ZN(n5694) );
  NOR2_X1 U6435 ( .A1(n6536), .A2(n5694), .ZN(n5275) );
  NAND2_X1 U6436 ( .A1(n5924), .A2(n5275), .ZN(n5676) );
  NOR2_X1 U6437 ( .A1(n6538), .A2(n5676), .ZN(n5678) );
  NAND2_X1 U6438 ( .A1(REIP_REG_22__SCAN_IN), .A2(n5678), .ZN(n5669) );
  NOR2_X1 U6439 ( .A1(n6666), .A2(n5669), .ZN(n5650) );
  AND3_X1 U6440 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5279) );
  NAND2_X1 U6441 ( .A1(n5650), .A2(n5279), .ZN(n5643) );
  NOR3_X1 U6442 ( .A1(n5643), .A2(REIP_REG_28__SCAN_IN), .A3(n6649), .ZN(n5284) );
  NAND2_X1 U6443 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5314) );
  NAND3_X1 U6444 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5277) );
  OR2_X1 U6445 ( .A1(n5863), .A2(n5275), .ZN(n5276) );
  NAND2_X1 U6446 ( .A1(n5276), .A2(n5834), .ZN(n5696) );
  AOI21_X1 U6447 ( .B1(n5936), .B2(n5277), .A(n5696), .ZN(n5668) );
  OAI21_X1 U6448 ( .B1(n5279), .B2(n5278), .A(n5668), .ZN(n5655) );
  AOI21_X1 U6449 ( .B1(n5924), .B2(n5314), .A(n5655), .ZN(n5315) );
  INV_X1 U6450 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6632) );
  AOI22_X1 U6451 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n5913), .B1(n5945), 
        .B2(n5280), .ZN(n5282) );
  NAND2_X1 U6452 ( .A1(n5969), .A2(EBX_REG_28__SCAN_IN), .ZN(n5281) );
  OAI211_X1 U6453 ( .C1(n5315), .C2(n6632), .A(n5282), .B(n5281), .ZN(n5283)
         );
  AOI211_X1 U6454 ( .C1(n5285), .C2(n5926), .A(n5284), .B(n5283), .ZN(n5286)
         );
  OAI21_X1 U6455 ( .B1(n5293), .B2(n5916), .A(n5286), .ZN(U2799) );
  AOI22_X1 U6456 ( .A1(n5994), .A2(DATAI_28_), .B1(n6003), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5292) );
  AND2_X1 U6457 ( .A1(n5289), .A2(n5288), .ZN(n5290) );
  NAND2_X1 U6458 ( .A1(n6004), .A2(DATAI_12_), .ZN(n5291) );
  OAI211_X1 U6459 ( .C1(n5293), .C2(n6012), .A(n5292), .B(n5291), .ZN(U2863)
         );
  AOI22_X1 U6460 ( .A1(n5994), .A2(DATAI_30_), .B1(n6003), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5295) );
  NAND2_X1 U6461 ( .A1(n6004), .A2(DATAI_14_), .ZN(n5294) );
  OAI211_X1 U6462 ( .C1(n5296), .C2(n6012), .A(n5295), .B(n5294), .ZN(U2861)
         );
  NAND2_X1 U6463 ( .A1(n5298), .A2(n5297), .ZN(n5303) );
  AOI22_X1 U6464 ( .A1(n5300), .A2(EAX_REG_31__SCAN_IN), .B1(n5299), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5301) );
  INV_X1 U6465 ( .A(n5301), .ZN(n5302) );
  NAND2_X1 U6467 ( .A1(n6139), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5304)
         );
  OAI211_X1 U6468 ( .C1(n6133), .C2(n5306), .A(n5305), .B(n5304), .ZN(n5307)
         );
  OAI21_X1 U6469 ( .B1(n5309), .B2(n6135), .A(n5308), .ZN(U2955) );
  NAND3_X1 U6470 ( .A1(n5313), .A2(n5310), .A3(n6011), .ZN(n5312) );
  AOI22_X1 U6471 ( .A1(n5994), .A2(DATAI_31_), .B1(n6003), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U6472 ( .A1(n5312), .A2(n5311), .ZN(U2860) );
  INV_X1 U6473 ( .A(n5313), .ZN(n5324) );
  OAI21_X1 U6474 ( .B1(n5338), .B2(REIP_REG_29__SCAN_IN), .A(n5315), .ZN(n5336) );
  INV_X1 U6475 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6764) );
  NAND2_X1 U6476 ( .A1(n6764), .A2(REIP_REG_29__SCAN_IN), .ZN(n5316) );
  NOR2_X1 U6477 ( .A1(n5338), .A2(n5316), .ZN(n5329) );
  OAI21_X1 U6478 ( .B1(n5336), .B2(n5329), .A(REIP_REG_31__SCAN_IN), .ZN(n5321) );
  AOI22_X1 U6479 ( .A1(n5317), .A2(EBX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n5913), .ZN(n5320) );
  INV_X1 U6480 ( .A(n5338), .ZN(n5318) );
  INV_X1 U6481 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6554) );
  NAND4_X1 U6482 ( .A1(n5318), .A2(REIP_REG_30__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .A4(n6554), .ZN(n5319) );
  NAND3_X1 U6483 ( .A1(n5321), .A2(n5320), .A3(n5319), .ZN(n5322) );
  AOI21_X1 U6484 ( .B1(n5352), .B2(n5926), .A(n5322), .ZN(n5323) );
  OAI21_X1 U6485 ( .B1(n5324), .B2(n5916), .A(n5323), .ZN(U2796) );
  NAND2_X1 U6486 ( .A1(n5325), .A2(n5881), .ZN(n5332) );
  AOI22_X1 U6487 ( .A1(n5326), .A2(n5945), .B1(n5913), .B2(
        PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5327) );
  OAI21_X1 U6488 ( .B1(n5909), .B2(n5328), .A(n5327), .ZN(n5330) );
  AOI211_X1 U6489 ( .C1(REIP_REG_30__SCAN_IN), .C2(n5336), .A(n5330), .B(n5329), .ZN(n5331) );
  OAI211_X1 U6490 ( .C1(n5333), .C2(n5962), .A(n5332), .B(n5331), .ZN(U2797)
         );
  NAND2_X1 U6491 ( .A1(n5355), .A2(n5881), .ZN(n5342) );
  OAI22_X1 U6492 ( .A1(n5335), .A2(n5959), .B1(n5963), .B2(n5334), .ZN(n5340)
         );
  INV_X1 U6493 ( .A(n5336), .ZN(n5337) );
  AOI21_X1 U6494 ( .B1(n6629), .B2(n5338), .A(n5337), .ZN(n5339) );
  AOI211_X1 U6495 ( .C1(EBX_REG_29__SCAN_IN), .C2(n5969), .A(n5340), .B(n5339), 
        .ZN(n5341) );
  OAI211_X1 U6496 ( .C1(n5962), .C2(n5356), .A(n5342), .B(n5341), .ZN(U2798)
         );
  AOI21_X1 U6497 ( .B1(n5344), .B2(n5472), .A(n5366), .ZN(n5464) );
  INV_X1 U6498 ( .A(n5464), .ZN(n5429) );
  XNOR2_X1 U6499 ( .A(n5567), .B(n5345), .ZN(n5557) );
  INV_X1 U6500 ( .A(n5557), .ZN(n5350) );
  INV_X1 U6501 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6720) );
  NAND2_X1 U6502 ( .A1(n5650), .A2(n6720), .ZN(n5659) );
  INV_X1 U6503 ( .A(n5659), .ZN(n5349) );
  INV_X1 U6504 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5373) );
  OAI22_X1 U6505 ( .A1(n5668), .A2(n6720), .B1(n5462), .B2(n5959), .ZN(n5346)
         );
  AOI21_X1 U6506 ( .B1(n5945), .B2(n5460), .A(n5346), .ZN(n5347) );
  OAI21_X1 U6507 ( .B1(n5909), .B2(n5373), .A(n5347), .ZN(n5348) );
  AOI211_X1 U6508 ( .C1(n5350), .C2(n5926), .A(n5349), .B(n5348), .ZN(n5351)
         );
  OAI21_X1 U6509 ( .B1(n5429), .B2(n5916), .A(n5351), .ZN(U2803) );
  INV_X1 U6510 ( .A(n5352), .ZN(n5354) );
  OAI22_X1 U6511 ( .A1(n5354), .A2(n5983), .B1(n5988), .B2(n5353), .ZN(U2828)
         );
  INV_X1 U6512 ( .A(n5355), .ZN(n5424) );
  OAI222_X1 U6513 ( .A1(n5719), .A2(n5424), .B1(n5357), .B2(n5988), .C1(n5356), 
        .C2(n5983), .ZN(U2830) );
  OAI21_X1 U6514 ( .B1(n5364), .B2(n2992), .A(n5359), .ZN(n5652) );
  AND2_X1 U6515 ( .A1(n2999), .A2(n5360), .ZN(n5361) );
  OR2_X1 U6516 ( .A1(n5361), .A2(n5197), .ZN(n5651) );
  INV_X1 U6517 ( .A(n5651), .ZN(n5543) );
  AOI22_X1 U6518 ( .A1(n5543), .A2(n5977), .B1(EBX_REG_26__SCAN_IN), .B2(n5362), .ZN(n5363) );
  OAI21_X1 U6519 ( .B1(n5652), .B2(n5984), .A(n5363), .ZN(U2833) );
  INV_X1 U6520 ( .A(n5364), .ZN(n5368) );
  OR2_X1 U6521 ( .A1(n5366), .A2(n5365), .ZN(n5367) );
  AND2_X1 U6522 ( .A1(n5368), .A2(n5367), .ZN(n5732) );
  INV_X1 U6523 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5372) );
  NAND2_X1 U6524 ( .A1(n5370), .A2(n5369), .ZN(n5371) );
  NAND2_X1 U6525 ( .A1(n2999), .A2(n5371), .ZN(n5660) );
  OAI222_X1 U6526 ( .A1(n5661), .A2(n5984), .B1(n5988), .B2(n5372), .C1(n5660), 
        .C2(n5983), .ZN(U2834) );
  OAI222_X1 U6527 ( .A1(n5429), .A2(n5984), .B1(n5373), .B2(n5988), .C1(n5983), 
        .C2(n5557), .ZN(U2835) );
  INV_X1 U6528 ( .A(n5374), .ZN(n5681) );
  INV_X1 U6529 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5375) );
  OAI222_X1 U6530 ( .A1(n5984), .A2(n5681), .B1(n5988), .B2(n5375), .C1(n5685), 
        .C2(n5983), .ZN(U2837) );
  AND2_X1 U6531 ( .A1(n5419), .A2(n5376), .ZN(n5391) );
  OR2_X1 U6532 ( .A1(n5391), .A2(n5377), .ZN(n5378) );
  NAND2_X1 U6533 ( .A1(n5379), .A2(n5378), .ZN(n5739) );
  INV_X1 U6534 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5383) );
  OR2_X1 U6535 ( .A1(n5381), .A2(n5380), .ZN(n5382) );
  NAND2_X1 U6536 ( .A1(n3624), .A2(n5382), .ZN(n5689) );
  OAI222_X1 U6537 ( .A1(n5739), .A2(n5719), .B1(n5383), .B2(n5988), .C1(n5983), 
        .C2(n5689), .ZN(U2838) );
  MUX2_X1 U6538 ( .A(n5385), .B(n5398), .S(n5384), .Z(n5387) );
  XNOR2_X1 U6539 ( .A(n5387), .B(n5386), .ZN(n5593) );
  INV_X1 U6540 ( .A(n5593), .ZN(n5697) );
  AND2_X1 U6541 ( .A1(n5419), .A2(n5388), .ZN(n5711) );
  NOR2_X1 U6542 ( .A1(n5711), .A2(n5389), .ZN(n5390) );
  OAI222_X1 U6543 ( .A1(n5697), .A2(n5983), .B1(n5988), .B2(n3613), .C1(n5743), 
        .C2(n5984), .ZN(U2839) );
  NAND2_X1 U6544 ( .A1(n5419), .A2(n5392), .ZN(n5710) );
  NAND2_X1 U6545 ( .A1(n5419), .A2(n5393), .ZN(n5762) );
  NAND2_X1 U6546 ( .A1(n5762), .A2(n5394), .ZN(n5395) );
  NAND2_X1 U6547 ( .A1(n5710), .A2(n5395), .ZN(n5990) );
  MUX2_X1 U6548 ( .A(n5398), .B(n5397), .S(n5396), .Z(n5402) );
  INV_X1 U6549 ( .A(n5602), .ZN(n5400) );
  INV_X1 U6550 ( .A(n5402), .ZN(n5399) );
  NAND2_X1 U6551 ( .A1(n5400), .A2(n5399), .ZN(n5715) );
  INV_X1 U6552 ( .A(n5715), .ZN(n5401) );
  AOI21_X1 U6553 ( .B1(n5602), .B2(n5402), .A(n5401), .ZN(n5818) );
  INV_X1 U6554 ( .A(n5818), .ZN(n5403) );
  OAI222_X1 U6555 ( .A1(n5990), .A2(n5984), .B1(n5404), .B2(n5988), .C1(n5983), 
        .C2(n5403), .ZN(U2841) );
  OR2_X1 U6556 ( .A1(n5407), .A2(n5406), .ZN(n5408) );
  NAND2_X1 U6557 ( .A1(n5405), .A2(n5408), .ZN(n5844) );
  INV_X1 U6558 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U6559 ( .A1(n5419), .A2(n5418), .ZN(n5434) );
  AND2_X1 U6560 ( .A1(n5419), .A2(n5418), .ZN(n5411) );
  OAI222_X1 U6561 ( .A1(n5844), .A2(n5983), .B1(n5988), .B2(n5413), .C1(n6001), 
        .C2(n5719), .ZN(U2843) );
  INV_X1 U6562 ( .A(n5414), .ZN(n5784) );
  NAND2_X1 U6563 ( .A1(n5784), .A2(n5415), .ZN(n5416) );
  NAND2_X1 U6564 ( .A1(n5417), .A2(n5416), .ZN(n5862) );
  INV_X1 U6565 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5421) );
  OR2_X1 U6566 ( .A1(n5419), .A2(n5418), .ZN(n5420) );
  INV_X1 U6567 ( .A(n5859), .ZN(n5440) );
  OAI222_X1 U6568 ( .A1(n5862), .A2(n5983), .B1(n5988), .B2(n5421), .C1(n5440), 
        .C2(n5984), .ZN(U2845) );
  AOI22_X1 U6569 ( .A1(n5994), .A2(DATAI_29_), .B1(n6003), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U6570 ( .A1(n6004), .A2(DATAI_13_), .ZN(n5422) );
  OAI211_X1 U6571 ( .C1(n5424), .C2(n6012), .A(n5423), .B(n5422), .ZN(U2862)
         );
  AOI22_X1 U6572 ( .A1(n6004), .A2(DATAI_10_), .B1(n6003), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U6573 ( .A1(n5994), .A2(DATAI_26_), .ZN(n5425) );
  OAI211_X1 U6574 ( .C1(n5652), .C2(n6012), .A(n5426), .B(n5425), .ZN(U2865)
         );
  AOI22_X1 U6575 ( .A1(n5994), .A2(DATAI_24_), .B1(n6003), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U6576 ( .A1(n6004), .A2(DATAI_8_), .ZN(n5427) );
  OAI211_X1 U6577 ( .C1(n5429), .C2(n6012), .A(n5428), .B(n5427), .ZN(U2867)
         );
  AOI22_X1 U6578 ( .A1(n6004), .A2(DATAI_6_), .B1(n6003), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6579 ( .A1(n5994), .A2(DATAI_22_), .ZN(n5430) );
  OAI211_X1 U6580 ( .C1(n5681), .C2(n6012), .A(n5431), .B(n5430), .ZN(U2869)
         );
  INV_X1 U6581 ( .A(n5432), .ZN(n5433) );
  AOI21_X1 U6582 ( .B1(n5435), .B2(n5434), .A(n5433), .ZN(n5978) );
  INV_X1 U6583 ( .A(n5978), .ZN(n5437) );
  AOI22_X1 U6584 ( .A1(n5438), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6003), .ZN(n5436) );
  OAI21_X1 U6585 ( .B1(n5437), .B2(n6012), .A(n5436), .ZN(U2876) );
  AOI22_X1 U6586 ( .A1(n5438), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n6003), .ZN(n5439) );
  OAI21_X1 U6587 ( .B1(n5440), .B2(n6012), .A(n5439), .ZN(U2877) );
  XNOR2_X1 U6588 ( .A(n3440), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5441)
         );
  XNOR2_X1 U6589 ( .A(n5442), .B(n5441), .ZN(n5545) );
  NAND2_X1 U6590 ( .A1(n6159), .A2(REIP_REG_26__SCAN_IN), .ZN(n5536) );
  OAI21_X1 U6591 ( .B1(n5769), .B2(n5443), .A(n5536), .ZN(n5445) );
  NOR2_X1 U6592 ( .A1(n5652), .A2(n6142), .ZN(n5444) );
  AOI211_X1 U6593 ( .C1(n5763), .C2(n5649), .A(n5445), .B(n5444), .ZN(n5446)
         );
  OAI21_X1 U6594 ( .B1(n6135), .B2(n5545), .A(n5446), .ZN(U2960) );
  NAND2_X1 U6595 ( .A1(n6159), .A2(REIP_REG_25__SCAN_IN), .ZN(n5547) );
  OAI21_X1 U6596 ( .B1(n5769), .B2(n5447), .A(n5547), .ZN(n5448) );
  AOI21_X1 U6597 ( .B1(n5763), .B2(n5664), .A(n5448), .ZN(n5453) );
  OAI21_X1 U6598 ( .B1(n5451), .B2(n5450), .A(n2987), .ZN(n5546) );
  NAND2_X1 U6599 ( .A1(n5546), .A2(n6129), .ZN(n5452) );
  OAI211_X1 U6600 ( .C1(n5661), .C2(n6142), .A(n5453), .B(n5452), .ZN(U2961)
         );
  NAND3_X1 U6601 ( .A1(n5454), .A2(n3440), .A3(n3007), .ZN(n5458) );
  NAND2_X1 U6602 ( .A1(n5480), .A2(n5455), .ZN(n5470) );
  NAND2_X1 U6603 ( .A1(n5458), .A2(n5457), .ZN(n5459) );
  XNOR2_X1 U6604 ( .A(n5459), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5562)
         );
  NAND2_X1 U6605 ( .A1(n5763), .A2(n5460), .ZN(n5461) );
  NAND2_X1 U6606 ( .A1(n6159), .A2(REIP_REG_24__SCAN_IN), .ZN(n5556) );
  OAI211_X1 U6607 ( .C1(n5769), .C2(n5462), .A(n5461), .B(n5556), .ZN(n5463)
         );
  AOI21_X1 U6608 ( .B1(n5464), .B2(n6128), .A(n5463), .ZN(n5465) );
  OAI21_X1 U6609 ( .B1(n5562), .B2(n6135), .A(n5465), .ZN(U2962) );
  NAND4_X1 U6610 ( .A1(n5468), .A2(n5467), .A3(n5466), .A4(n3440), .ZN(n5469)
         );
  NAND2_X1 U6611 ( .A1(n5470), .A2(n5469), .ZN(n5471) );
  XNOR2_X1 U6612 ( .A(n5471), .B(n5569), .ZN(n5563) );
  INV_X1 U6613 ( .A(n5563), .ZN(n5479) );
  INV_X1 U6614 ( .A(n5472), .ZN(n5473) );
  AOI21_X1 U6615 ( .B1(n5475), .B2(n5474), .A(n5473), .ZN(n5735) );
  NAND2_X1 U6616 ( .A1(n6159), .A2(REIP_REG_23__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U6617 ( .A1(n6139), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5476)
         );
  OAI211_X1 U6618 ( .C1(n6133), .C2(n5675), .A(n5568), .B(n5476), .ZN(n5477)
         );
  AOI21_X1 U6619 ( .B1(n5735), .B2(n6128), .A(n5477), .ZN(n5478) );
  OAI21_X1 U6620 ( .B1(n5479), .B2(n6135), .A(n5478), .ZN(U2963) );
  INV_X1 U6621 ( .A(n5480), .ZN(n5481) );
  OAI21_X1 U6622 ( .B1(n5483), .B2(n5482), .A(n5481), .ZN(n5575) );
  NAND2_X1 U6623 ( .A1(n5575), .A2(n6129), .ZN(n5486) );
  NOR2_X1 U6624 ( .A1(n6134), .A2(n6538), .ZN(n5577) );
  NOR2_X1 U6625 ( .A1(n6133), .A2(n5693), .ZN(n5484) );
  AOI211_X1 U6626 ( .C1(n6139), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5577), 
        .B(n5484), .ZN(n5485) );
  OAI211_X1 U6627 ( .C1(n6142), .C2(n5739), .A(n5486), .B(n5485), .ZN(U2965)
         );
  XNOR2_X1 U6628 ( .A(n5487), .B(n5488), .ZN(n5595) );
  INV_X1 U6629 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U6630 ( .A1(n6159), .A2(REIP_REG_20__SCAN_IN), .ZN(n5586) );
  OAI21_X1 U6631 ( .B1(n5769), .B2(n5702), .A(n5586), .ZN(n5490) );
  NOR2_X1 U6632 ( .A1(n5743), .A2(n6142), .ZN(n5489) );
  AOI211_X1 U6633 ( .C1(n5763), .C2(n5699), .A(n5490), .B(n5489), .ZN(n5491)
         );
  OAI21_X1 U6634 ( .B1(n5595), .B2(n6135), .A(n5491), .ZN(U2966) );
  NOR2_X1 U6635 ( .A1(n5493), .A2(n5494), .ZN(n5497) );
  NOR2_X1 U6636 ( .A1(n5495), .A2(n5603), .ZN(n5496) );
  MUX2_X1 U6637 ( .A(n5497), .B(n5496), .S(n3440), .Z(n5498) );
  XOR2_X1 U6638 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(n5498), .Z(n5777) );
  NAND2_X1 U6639 ( .A1(n5777), .A2(n6129), .ZN(n5502) );
  OAI22_X1 U6640 ( .A1(n5769), .A2(n5499), .B1(n6134), .B2(n6533), .ZN(n5500)
         );
  AOI21_X1 U6641 ( .B1(n5763), .B2(n5815), .A(n5500), .ZN(n5501) );
  OAI211_X1 U6642 ( .C1(n6142), .C2(n5990), .A(n5502), .B(n5501), .ZN(U2968)
         );
  XNOR2_X1 U6643 ( .A(n3440), .B(n5620), .ZN(n5503) );
  XNOR2_X1 U6644 ( .A(n5493), .B(n5503), .ZN(n5610) );
  NAND2_X1 U6645 ( .A1(n5610), .A2(n6129), .ZN(n5506) );
  NOR2_X1 U6646 ( .A1(n6134), .A2(n6530), .ZN(n5615) );
  NOR2_X1 U6647 ( .A1(n6133), .A2(n5840), .ZN(n5504) );
  AOI211_X1 U6648 ( .C1(n6139), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5615), 
        .B(n5504), .ZN(n5505) );
  OAI211_X1 U6649 ( .C1(n6142), .C2(n6001), .A(n5506), .B(n5505), .ZN(U2970)
         );
  NAND2_X1 U6650 ( .A1(n6139), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5507)
         );
  OAI211_X1 U6651 ( .C1(n6133), .C2(n5509), .A(n5508), .B(n5507), .ZN(n5510)
         );
  AOI21_X1 U6652 ( .B1(n5978), .B2(n6128), .A(n5510), .ZN(n5511) );
  OAI21_X1 U6653 ( .B1(n6135), .B2(n5512), .A(n5511), .ZN(U2971) );
  NAND2_X1 U6654 ( .A1(n5529), .A2(n5514), .ZN(n5517) );
  XNOR2_X1 U6655 ( .A(n3440), .B(n5515), .ZN(n5516) );
  XNOR2_X1 U6656 ( .A(n5517), .B(n5516), .ZN(n5637) );
  AOI22_X1 U6657 ( .A1(n6139), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6159), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5518) );
  OAI21_X1 U6658 ( .B1(n5857), .B2(n6133), .A(n5518), .ZN(n5519) );
  AOI21_X1 U6659 ( .B1(n5859), .B2(n6128), .A(n5519), .ZN(n5520) );
  OAI21_X1 U6660 ( .B1(n5637), .B2(n6135), .A(n5520), .ZN(U2972) );
  XNOR2_X1 U6661 ( .A(n5523), .B(n5522), .ZN(n6007) );
  OR2_X1 U6662 ( .A1(n5525), .A2(n5524), .ZN(n5527) );
  NAND2_X1 U6663 ( .A1(n5527), .A2(n5526), .ZN(n5532) );
  AND2_X1 U6664 ( .A1(n5529), .A2(n5528), .ZN(n5530) );
  OAI21_X1 U6665 ( .B1(n5532), .B2(n5531), .A(n5530), .ZN(n5787) );
  NAND2_X1 U6666 ( .A1(n5787), .A2(n6129), .ZN(n5535) );
  AND2_X1 U6667 ( .A1(n6159), .A2(REIP_REG_13__SCAN_IN), .ZN(n5785) );
  NOR2_X1 U6668 ( .A1(n6133), .A2(n5868), .ZN(n5533) );
  AOI211_X1 U6669 ( .C1(n6139), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5785), 
        .B(n5533), .ZN(n5534) );
  OAI211_X1 U6670 ( .C1(n6007), .C2(n6142), .A(n5535), .B(n5534), .ZN(U2973)
         );
  INV_X1 U6671 ( .A(n5560), .ZN(n5549) );
  OAI21_X1 U6672 ( .B1(n5549), .B2(n5537), .A(n5536), .ZN(n5542) );
  INV_X1 U6673 ( .A(n5538), .ZN(n5554) );
  NOR3_X1 U6674 ( .A1(n5554), .A2(n5540), .A3(n5539), .ZN(n5541) );
  AOI211_X1 U6675 ( .C1(n5543), .C2(n6161), .A(n5542), .B(n5541), .ZN(n5544)
         );
  OAI21_X1 U6676 ( .B1(n5545), .B2(n5636), .A(n5544), .ZN(U2992) );
  NAND2_X1 U6677 ( .A1(n5546), .A2(n6166), .ZN(n5553) );
  INV_X1 U6678 ( .A(n5660), .ZN(n5551) );
  OAI21_X1 U6679 ( .B1(n5549), .B2(n5548), .A(n5547), .ZN(n5550) );
  AOI21_X1 U6680 ( .B1(n5551), .B2(n6161), .A(n5550), .ZN(n5552) );
  OAI211_X1 U6681 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5554), .A(n5553), .B(n5552), .ZN(U2993) );
  OAI21_X1 U6682 ( .B1(n5574), .B2(n5569), .A(n5555), .ZN(n5559) );
  OAI21_X1 U6683 ( .B1(n5557), .B2(n5631), .A(n5556), .ZN(n5558) );
  AOI21_X1 U6684 ( .B1(n5560), .B2(n5559), .A(n5558), .ZN(n5561) );
  OAI21_X1 U6685 ( .B1(n5562), .B2(n5636), .A(n5561), .ZN(U2994) );
  NAND2_X1 U6686 ( .A1(n5563), .A2(n6166), .ZN(n5573) );
  AND2_X1 U6687 ( .A1(n5565), .A2(n5564), .ZN(n5566) );
  NOR2_X1 U6688 ( .A1(n5567), .A2(n5566), .ZN(n5723) );
  OAI21_X1 U6689 ( .B1(n5570), .B2(n5569), .A(n5568), .ZN(n5571) );
  AOI21_X1 U6690 ( .B1(n5723), .B2(n6161), .A(n5571), .ZN(n5572) );
  OAI211_X1 U6691 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5574), .A(n5573), .B(n5572), .ZN(U2995) );
  NAND2_X1 U6692 ( .A1(n5575), .A2(n6166), .ZN(n5580) );
  NOR2_X1 U6693 ( .A1(n5689), .A2(n5631), .ZN(n5576) );
  AOI211_X1 U6694 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5578), .A(n5577), .B(n5576), .ZN(n5579) );
  OAI211_X1 U6695 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5581), .A(n5580), .B(n5579), .ZN(U2997) );
  OAI21_X1 U6696 ( .B1(n5603), .B2(n5582), .A(n6162), .ZN(n5604) );
  NAND3_X1 U6697 ( .A1(n5605), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n5604), .ZN(n5583) );
  AOI21_X1 U6698 ( .B1(n6169), .B2(n5603), .A(n5583), .ZN(n5781) );
  AOI21_X1 U6699 ( .B1(n5585), .B2(n5584), .A(n5781), .ZN(n5770) );
  INV_X1 U6700 ( .A(n5770), .ZN(n5588) );
  OAI21_X1 U6701 ( .B1(n5588), .B2(n5587), .A(n5586), .ZN(n5592) );
  NAND2_X1 U6702 ( .A1(n5776), .A2(n5589), .ZN(n5775) );
  XNOR2_X1 U6703 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .B(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5590) );
  NOR2_X1 U6704 ( .A1(n5775), .A2(n5590), .ZN(n5591) );
  AOI211_X1 U6705 ( .C1(n6161), .C2(n5593), .A(n5592), .B(n5591), .ZN(n5594)
         );
  OAI21_X1 U6706 ( .B1(n5595), .B2(n5636), .A(n5594), .ZN(U2998) );
  INV_X1 U6707 ( .A(n5776), .ZN(n5609) );
  NAND2_X1 U6708 ( .A1(n5596), .A2(n5620), .ZN(n5598) );
  NAND3_X1 U6709 ( .A1(n5493), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n3447), .ZN(n5597) );
  OAI21_X1 U6710 ( .B1(n5493), .B2(n5598), .A(n5597), .ZN(n5599) );
  XNOR2_X1 U6711 ( .A(n5599), .B(n5603), .ZN(n5765) );
  NAND2_X1 U6712 ( .A1(n5765), .A2(n6166), .ZN(n5608) );
  NAND2_X1 U6713 ( .A1(n5405), .A2(n5600), .ZN(n5601) );
  AND2_X1 U6714 ( .A1(n5602), .A2(n5601), .ZN(n5973) );
  INV_X1 U6715 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5825) );
  NOR2_X1 U6716 ( .A1(n6134), .A2(n5825), .ZN(n5766) );
  AOI21_X1 U6717 ( .B1(n5605), .B2(n5604), .A(n5603), .ZN(n5606) );
  AOI211_X1 U6718 ( .C1(n5973), .C2(n6161), .A(n5766), .B(n5606), .ZN(n5607)
         );
  OAI211_X1 U6719 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5609), .A(n5608), .B(n5607), .ZN(U3001) );
  NAND2_X1 U6720 ( .A1(n5610), .A2(n6166), .ZN(n5619) );
  INV_X1 U6721 ( .A(n5611), .ZN(n5612) );
  AOI21_X1 U6722 ( .B1(n5613), .B2(n5620), .A(n5612), .ZN(n5616) );
  NOR2_X1 U6723 ( .A1(n5844), .A2(n5631), .ZN(n5614) );
  AOI211_X1 U6724 ( .C1(n5617), .C2(n5616), .A(n5615), .B(n5614), .ZN(n5618)
         );
  OAI211_X1 U6725 ( .C1(n5621), .C2(n5620), .A(n5619), .B(n5618), .ZN(U3002)
         );
  NAND3_X1 U6726 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n5622), .ZN(n5790) );
  AOI21_X1 U6727 ( .B1(n5624), .B2(n5623), .A(n5790), .ZN(n5629) );
  NOR2_X1 U6728 ( .A1(n6151), .A2(n3439), .ZN(n5628) );
  NAND2_X1 U6729 ( .A1(n5625), .A2(n5630), .ZN(n5626) );
  OAI211_X1 U6730 ( .C1(n5628), .C2(n5627), .A(n5626), .B(n6150), .ZN(n5786)
         );
  OAI21_X1 U6731 ( .B1(n5629), .B2(n5786), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5635) );
  NOR3_X1 U6732 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5791), .A3(n5630), 
        .ZN(n5633) );
  OAI22_X1 U6733 ( .A1(n5862), .A2(n5631), .B1(n6527), .B2(n6134), .ZN(n5632)
         );
  NOR2_X1 U6734 ( .A1(n5633), .A2(n5632), .ZN(n5634) );
  OAI211_X1 U6735 ( .C1(n5637), .C2(n5636), .A(n5635), .B(n5634), .ZN(U3004)
         );
  AOI21_X1 U6736 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n5639), .A(n5638), .ZN(
        n5640) );
  INV_X1 U6737 ( .A(n5640), .ZN(U2788) );
  INV_X1 U6738 ( .A(n5655), .ZN(n5642) );
  AOI22_X1 U6739 ( .A1(n5969), .A2(EBX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n5913), .ZN(n5641) );
  OAI221_X1 U6740 ( .B1(n5643), .B2(REIP_REG_27__SCAN_IN), .C1(n5642), .C2(
        n6649), .A(n5641), .ZN(n5644) );
  INV_X1 U6741 ( .A(n5644), .ZN(n5647) );
  OAI22_X1 U6742 ( .A1(n5728), .A2(n5916), .B1(n5718), .B2(n5962), .ZN(n5645)
         );
  INV_X1 U6743 ( .A(n5645), .ZN(n5646) );
  OAI211_X1 U6744 ( .C1(n5648), .C2(n5963), .A(n5647), .B(n5646), .ZN(U2800)
         );
  AOI22_X1 U6745 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n5913), .B1(n5649), 
        .B2(n5945), .ZN(n5657) );
  INV_X1 U6746 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6544) );
  NAND2_X1 U6747 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5650), .ZN(n5667) );
  INV_X1 U6748 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6722) );
  OAI21_X1 U6749 ( .B1(n6544), .B2(n5667), .A(n6722), .ZN(n5654) );
  OAI22_X1 U6750 ( .A1(n5652), .A2(n5916), .B1(n5651), .B2(n5962), .ZN(n5653)
         );
  AOI21_X1 U6751 ( .B1(n5655), .B2(n5654), .A(n5653), .ZN(n5656) );
  OAI211_X1 U6752 ( .C1(n5909), .C2(n5658), .A(n5657), .B(n5656), .ZN(U2801)
         );
  AOI22_X1 U6753 ( .A1(EBX_REG_25__SCAN_IN), .A2(n5969), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5913), .ZN(n5666) );
  AOI21_X1 U6754 ( .B1(n5668), .B2(n5659), .A(n6544), .ZN(n5663) );
  OAI22_X1 U6755 ( .A1(n5661), .A2(n5916), .B1(n5962), .B2(n5660), .ZN(n5662)
         );
  AOI211_X1 U6756 ( .C1(n5945), .C2(n5664), .A(n5663), .B(n5662), .ZN(n5665)
         );
  OAI211_X1 U6757 ( .C1(REIP_REG_25__SCAN_IN), .C2(n5667), .A(n5666), .B(n5665), .ZN(U2802) );
  AOI21_X1 U6758 ( .B1(n5669), .B2(n6666), .A(n5668), .ZN(n5672) );
  AOI22_X1 U6759 ( .A1(n5969), .A2(EBX_REG_23__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n5913), .ZN(n5670) );
  INV_X1 U6760 ( .A(n5670), .ZN(n5671) );
  NOR2_X1 U6761 ( .A1(n5672), .A2(n5671), .ZN(n5674) );
  AOI22_X1 U6762 ( .A1(n5735), .A2(n5881), .B1(n5723), .B2(n5926), .ZN(n5673)
         );
  OAI211_X1 U6763 ( .C1(n5675), .C2(n5963), .A(n5674), .B(n5673), .ZN(U2804)
         );
  AOI22_X1 U6764 ( .A1(n5969), .A2(EBX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n5913), .ZN(n5680) );
  NOR2_X1 U6765 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5676), .ZN(n5688) );
  INV_X1 U6766 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6634) );
  OR3_X1 U6767 ( .A1(n5696), .A2(n5688), .A3(n6634), .ZN(n5677) );
  OAI21_X1 U6768 ( .B1(n5678), .B2(REIP_REG_22__SCAN_IN), .A(n5677), .ZN(n5679) );
  OAI211_X1 U6769 ( .C1(n5681), .C2(n5916), .A(n5680), .B(n5679), .ZN(n5682)
         );
  AOI21_X1 U6770 ( .B1(n5683), .B2(n5945), .A(n5682), .ZN(n5684) );
  OAI21_X1 U6771 ( .B1(n5685), .B2(n5962), .A(n5684), .ZN(U2805) );
  AOI22_X1 U6772 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n5913), .B1(
        REIP_REG_21__SCAN_IN), .B2(n5696), .ZN(n5686) );
  INV_X1 U6773 ( .A(n5686), .ZN(n5687) );
  AOI211_X1 U6774 ( .C1(EBX_REG_21__SCAN_IN), .C2(n5969), .A(n5688), .B(n5687), 
        .ZN(n5692) );
  OAI22_X1 U6775 ( .A1(n5739), .A2(n5916), .B1(n5962), .B2(n5689), .ZN(n5690)
         );
  INV_X1 U6776 ( .A(n5690), .ZN(n5691) );
  OAI211_X1 U6777 ( .C1(n5693), .C2(n5963), .A(n5692), .B(n5691), .ZN(U2806)
         );
  OAI21_X1 U6778 ( .B1(n5863), .B2(n5694), .A(n6536), .ZN(n5695) );
  AOI22_X1 U6779 ( .A1(EBX_REG_20__SCAN_IN), .A2(n5969), .B1(n5696), .B2(n5695), .ZN(n5701) );
  OAI22_X1 U6780 ( .A1(n5743), .A2(n5916), .B1(n5962), .B2(n5697), .ZN(n5698)
         );
  AOI21_X1 U6781 ( .B1(n5699), .B2(n5945), .A(n5698), .ZN(n5700) );
  OAI211_X1 U6782 ( .C1(n5702), .C2(n5959), .A(n5701), .B(n5700), .ZN(U2807)
         );
  INV_X1 U6783 ( .A(n5704), .ZN(n5703) );
  OAI21_X1 U6784 ( .B1(n5863), .B2(n5703), .A(n5834), .ZN(n5829) );
  NOR3_X1 U6785 ( .A1(n5863), .A2(REIP_REG_18__SCAN_IN), .A3(n5704), .ZN(n5814) );
  OAI21_X1 U6786 ( .B1(n5829), .B2(n5814), .A(REIP_REG_19__SCAN_IN), .ZN(n5707) );
  INV_X1 U6787 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6734) );
  NAND3_X1 U6788 ( .A1(n5924), .A2(n6734), .A3(n5705), .ZN(n5706) );
  OAI211_X1 U6789 ( .C1(n5909), .C2(n5727), .A(n5707), .B(n5706), .ZN(n5708)
         );
  AOI211_X1 U6790 ( .C1(n5913), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5921), 
        .B(n5708), .ZN(n5717) );
  AND2_X1 U6791 ( .A1(n5710), .A2(n5709), .ZN(n5712) );
  INV_X1 U6792 ( .A(n5713), .ZN(n5714) );
  XNOR2_X1 U6793 ( .A(n5715), .B(n5714), .ZN(n5771) );
  AOI22_X1 U6794 ( .A1(n5755), .A2(n5881), .B1(n5926), .B2(n5771), .ZN(n5716)
         );
  OAI211_X1 U6795 ( .C1(n5758), .C2(n5963), .A(n5717), .B(n5716), .ZN(U2808)
         );
  OAI22_X1 U6796 ( .A1(n5728), .A2(n5719), .B1(n5718), .B2(n5983), .ZN(n5720)
         );
  INV_X1 U6797 ( .A(n5720), .ZN(n5721) );
  OAI21_X1 U6798 ( .B1(n5988), .B2(n5722), .A(n5721), .ZN(U2832) );
  INV_X1 U6799 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5725) );
  AOI22_X1 U6800 ( .A1(n5735), .A2(n4196), .B1(n5723), .B2(n5977), .ZN(n5724)
         );
  OAI21_X1 U6801 ( .B1(n5988), .B2(n5725), .A(n5724), .ZN(U2836) );
  AOI22_X1 U6802 ( .A1(n5755), .A2(n4196), .B1(n5977), .B2(n5771), .ZN(n5726)
         );
  OAI21_X1 U6803 ( .B1(n5988), .B2(n5727), .A(n5726), .ZN(U2840) );
  INV_X1 U6804 ( .A(n5994), .ZN(n6000) );
  OAI22_X1 U6805 ( .A1(n5728), .A2(n6012), .B1(n6000), .B2(n6657), .ZN(n5729)
         );
  INV_X1 U6806 ( .A(n5729), .ZN(n5731) );
  AOI22_X1 U6807 ( .A1(n6004), .A2(DATAI_11_), .B1(n6003), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U6808 ( .A1(n5731), .A2(n5730), .ZN(U2864) );
  INV_X1 U6809 ( .A(n6012), .ZN(n5995) );
  AOI22_X1 U6810 ( .A1(n5732), .A2(n5995), .B1(n5994), .B2(DATAI_25_), .ZN(
        n5734) );
  AOI22_X1 U6811 ( .A1(n6004), .A2(DATAI_9_), .B1(n6003), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U6812 ( .A1(n5734), .A2(n5733), .ZN(U2866) );
  AOI22_X1 U6813 ( .A1(n5735), .A2(n5995), .B1(n5994), .B2(DATAI_23_), .ZN(
        n5737) );
  AOI22_X1 U6814 ( .A1(n6004), .A2(DATAI_7_), .B1(n6003), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U6815 ( .A1(n5737), .A2(n5736), .ZN(U2868) );
  OAI22_X1 U6816 ( .A1(n5739), .A2(n6012), .B1(n6000), .B2(n5738), .ZN(n5740)
         );
  INV_X1 U6817 ( .A(n5740), .ZN(n5742) );
  AOI22_X1 U6818 ( .A1(n6004), .A2(DATAI_5_), .B1(n6003), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5741) );
  NAND2_X1 U6819 ( .A1(n5742), .A2(n5741), .ZN(U2870) );
  INV_X1 U6820 ( .A(n5743), .ZN(n5744) );
  AOI22_X1 U6821 ( .A1(n5744), .A2(n5995), .B1(n5994), .B2(DATAI_20_), .ZN(
        n5746) );
  AOI22_X1 U6822 ( .A1(n6004), .A2(DATAI_4_), .B1(n6003), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5745) );
  NAND2_X1 U6823 ( .A1(n5746), .A2(n5745), .ZN(U2871) );
  AOI22_X1 U6824 ( .A1(n5755), .A2(n5995), .B1(n5994), .B2(DATAI_19_), .ZN(
        n5748) );
  AOI22_X1 U6825 ( .A1(n6004), .A2(DATAI_3_), .B1(n6003), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5747) );
  NAND2_X1 U6826 ( .A1(n5748), .A2(n5747), .ZN(U2872) );
  AOI22_X1 U6827 ( .A1(n6159), .A2(REIP_REG_19__SCAN_IN), .B1(n6139), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5757) );
  OAI21_X1 U6828 ( .B1(n5751), .B2(n5750), .A(n5749), .ZN(n5754) );
  XNOR2_X1 U6829 ( .A(n5752), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5753)
         );
  MUX2_X1 U6830 ( .A(n5754), .B(n5753), .S(n3440), .Z(n5772) );
  AOI22_X1 U6831 ( .A1(n5772), .A2(n6129), .B1(n6128), .B2(n5755), .ZN(n5756)
         );
  OAI211_X1 U6832 ( .C1(n6133), .C2(n5758), .A(n5757), .B(n5756), .ZN(U2967)
         );
  INV_X1 U6833 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5826) );
  INV_X1 U6834 ( .A(n5832), .ZN(n5764) );
  AOI222_X1 U6835 ( .A1(n5765), .A2(n6129), .B1(n5764), .B2(n5763), .C1(n6128), 
        .C2(n5996), .ZN(n5768) );
  INV_X1 U6836 ( .A(n5766), .ZN(n5767) );
  OAI211_X1 U6837 ( .C1(n5826), .C2(n5769), .A(n5768), .B(n5767), .ZN(U2969)
         );
  AOI22_X1 U6838 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n5770), .B1(n6159), .B2(REIP_REG_19__SCAN_IN), .ZN(n5774) );
  AOI22_X1 U6839 ( .A1(n5772), .A2(n6166), .B1(n6161), .B2(n5771), .ZN(n5773)
         );
  OAI211_X1 U6840 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5775), .A(n5774), .B(n5773), .ZN(U2999) );
  AOI21_X1 U6841 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5776), .A(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5780) );
  AOI22_X1 U6842 ( .A1(n5777), .A2(n6166), .B1(n6161), .B2(n5818), .ZN(n5779)
         );
  NAND2_X1 U6843 ( .A1(n6159), .A2(REIP_REG_18__SCAN_IN), .ZN(n5778) );
  OAI211_X1 U6844 ( .C1(n5781), .C2(n5780), .A(n5779), .B(n5778), .ZN(U3000)
         );
  NAND2_X1 U6845 ( .A1(n5157), .A2(n5782), .ZN(n5783) );
  AND2_X1 U6846 ( .A1(n5784), .A2(n5783), .ZN(n5981) );
  AOI21_X1 U6847 ( .B1(n5981), .B2(n6161), .A(n5785), .ZN(n5789) );
  AOI22_X1 U6848 ( .A1(n5787), .A2(n6166), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5786), .ZN(n5788) );
  OAI211_X1 U6849 ( .C1(n5791), .C2(n5790), .A(n5789), .B(n5788), .ZN(U3005)
         );
  INV_X1 U6850 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6506) );
  AOI21_X1 U6851 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6506), .A(n6500), .ZN(n5797) );
  INV_X1 U6852 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5792) );
  NAND2_X1 U6853 ( .A1(n6500), .A2(STATE_REG_1__SCAN_IN), .ZN(n6541) );
  AOI21_X1 U6854 ( .B1(n5797), .B2(n5792), .A(n6778), .ZN(U2789) );
  NAND2_X1 U6855 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6582), .ZN(n5795) );
  OAI21_X1 U6856 ( .B1(n5793), .B2(n6481), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5794) );
  OAI21_X1 U6857 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5795), .A(n5794), .ZN(
        U2790) );
  INV_X1 U6858 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6651) );
  NOR2_X1 U6859 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5798) );
  NOR2_X1 U6860 ( .A1(n6778), .A2(n5798), .ZN(n5796) );
  AOI22_X1 U6861 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n6778), .B1(n6651), .B2(
        n5796), .ZN(U2791) );
  NOR2_X1 U6862 ( .A1(n6778), .A2(n5797), .ZN(n6558) );
  OAI21_X1 U6863 ( .B1(BS16_N), .B2(n5798), .A(n6558), .ZN(n6556) );
  OAI21_X1 U6864 ( .B1(n6558), .B2(n6723), .A(n6556), .ZN(U2792) );
  OAI21_X1 U6865 ( .B1(n5799), .B2(n6660), .A(n6135), .ZN(U2793) );
  NOR4_X1 U6866 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5803) );
  NOR4_X1 U6867 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n5802) );
  NOR4_X1 U6868 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5801) );
  NOR4_X1 U6869 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5800) );
  NAND4_X1 U6870 ( .A1(n5803), .A2(n5802), .A3(n5801), .A4(n5800), .ZN(n5809)
         );
  NOR4_X1 U6871 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n5807) );
  AOI211_X1 U6872 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_2__SCAN_IN), .B(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n5806) );
  NOR4_X1 U6873 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n5805) );
  NOR4_X1 U6874 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n5804) );
  NAND4_X1 U6875 ( .A1(n5807), .A2(n5806), .A3(n5805), .A4(n5804), .ZN(n5808)
         );
  NOR2_X1 U6876 ( .A1(n5809), .A2(n5808), .ZN(n6574) );
  INV_X1 U6877 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6662) );
  NOR3_X1 U6878 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5811) );
  OAI21_X1 U6879 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5811), .A(n6574), .ZN(n5810)
         );
  OAI21_X1 U6880 ( .B1(n6574), .B2(n6662), .A(n5810), .ZN(U2794) );
  INV_X1 U6881 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6557) );
  AOI21_X1 U6882 ( .B1(n6571), .B2(n6557), .A(n5811), .ZN(n5813) );
  INV_X1 U6883 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5812) );
  INV_X1 U6884 ( .A(n6574), .ZN(n6577) );
  AOI22_X1 U6885 ( .A1(n6574), .A2(n5813), .B1(n5812), .B2(n6577), .ZN(U2795)
         );
  AOI22_X1 U6886 ( .A1(EBX_REG_18__SCAN_IN), .A2(n5969), .B1(
        REIP_REG_18__SCAN_IN), .B2(n5829), .ZN(n5822) );
  AOI211_X1 U6887 ( .C1(n5913), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5814), 
        .B(n5921), .ZN(n5821) );
  INV_X1 U6888 ( .A(n5815), .ZN(n5816) );
  OAI22_X1 U6889 ( .A1(n5990), .A2(n5916), .B1(n5816), .B2(n5963), .ZN(n5817)
         );
  INV_X1 U6890 ( .A(n5817), .ZN(n5820) );
  NAND2_X1 U6891 ( .A1(n5926), .A2(n5818), .ZN(n5819) );
  NAND4_X1 U6892 ( .A1(n5822), .A2(n5821), .A3(n5820), .A4(n5819), .ZN(U2809)
         );
  INV_X1 U6893 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6530) );
  INV_X1 U6894 ( .A(n5823), .ZN(n5833) );
  OR2_X1 U6895 ( .A1(n5863), .A2(n5833), .ZN(n5845) );
  INV_X1 U6896 ( .A(n5845), .ZN(n5824) );
  NAND2_X1 U6897 ( .A1(n5824), .A2(REIP_REG_15__SCAN_IN), .ZN(n5838) );
  OAI21_X1 U6898 ( .B1(n6530), .B2(n5838), .A(n5825), .ZN(n5828) );
  INV_X1 U6899 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5975) );
  OAI22_X1 U6900 ( .A1(n5909), .A2(n5975), .B1(n5826), .B2(n5959), .ZN(n5827)
         );
  AOI211_X1 U6901 ( .C1(n5829), .C2(n5828), .A(n5921), .B(n5827), .ZN(n5831)
         );
  AOI22_X1 U6902 ( .A1(n5996), .A2(n5881), .B1(n5926), .B2(n5973), .ZN(n5830)
         );
  OAI211_X1 U6903 ( .C1(n5832), .C2(n5963), .A(n5831), .B(n5830), .ZN(U2810)
         );
  NAND2_X1 U6904 ( .A1(n5924), .A2(n5833), .ZN(n5854) );
  NAND2_X1 U6905 ( .A1(n5854), .A2(n5834), .ZN(n5852) );
  INV_X1 U6906 ( .A(n5852), .ZN(n5835) );
  OAI21_X1 U6907 ( .B1(REIP_REG_15__SCAN_IN), .B2(n5863), .A(n5835), .ZN(n5836) );
  AOI22_X1 U6908 ( .A1(EBX_REG_16__SCAN_IN), .A2(n5969), .B1(
        REIP_REG_16__SCAN_IN), .B2(n5836), .ZN(n5837) );
  OAI21_X1 U6909 ( .B1(REIP_REG_16__SCAN_IN), .B2(n5838), .A(n5837), .ZN(n5839) );
  AOI211_X1 U6910 ( .C1(n5913), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5921), 
        .B(n5839), .ZN(n5843) );
  OAI22_X1 U6911 ( .A1(n6001), .A2(n5916), .B1(n5840), .B2(n5963), .ZN(n5841)
         );
  INV_X1 U6912 ( .A(n5841), .ZN(n5842) );
  OAI211_X1 U6913 ( .C1(n5962), .C2(n5844), .A(n5843), .B(n5842), .ZN(U2811)
         );
  AOI22_X1 U6914 ( .A1(EBX_REG_15__SCAN_IN), .A2(n5969), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5852), .ZN(n5851) );
  NOR2_X1 U6915 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5845), .ZN(n5846) );
  AOI211_X1 U6916 ( .C1(n5913), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5921), 
        .B(n5846), .ZN(n5850) );
  AOI22_X1 U6917 ( .A1(n5978), .A2(n5881), .B1(n5945), .B2(n5847), .ZN(n5849)
         );
  NAND2_X1 U6918 ( .A1(n5926), .A2(n5976), .ZN(n5848) );
  NAND4_X1 U6919 ( .A1(n5851), .A2(n5850), .A3(n5849), .A4(n5848), .ZN(U2812)
         );
  AOI22_X1 U6920 ( .A1(EBX_REG_14__SCAN_IN), .A2(n5969), .B1(
        REIP_REG_14__SCAN_IN), .B2(n5852), .ZN(n5853) );
  OAI21_X1 U6921 ( .B1(n5855), .B2(n5854), .A(n5853), .ZN(n5856) );
  AOI211_X1 U6922 ( .C1(n5913), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5921), 
        .B(n5856), .ZN(n5861) );
  INV_X1 U6923 ( .A(n5857), .ZN(n5858) );
  AOI22_X1 U6924 ( .A1(n5859), .A2(n5881), .B1(n5858), .B2(n5945), .ZN(n5860)
         );
  OAI211_X1 U6925 ( .C1(n5962), .C2(n5862), .A(n5861), .B(n5860), .ZN(U2813)
         );
  OAI21_X1 U6926 ( .B1(REIP_REG_12__SCAN_IN), .B2(n5863), .A(n5873), .ZN(n5864) );
  AOI22_X1 U6927 ( .A1(n5926), .A2(n5981), .B1(REIP_REG_13__SCAN_IN), .B2(
        n5864), .ZN(n5872) );
  NAND3_X1 U6928 ( .A1(n5924), .A2(REIP_REG_12__SCAN_IN), .A3(n5875), .ZN(
        n5866) );
  OAI22_X1 U6929 ( .A1(REIP_REG_13__SCAN_IN), .A2(n5866), .B1(n5865), .B2(
        n5959), .ZN(n5867) );
  AOI211_X1 U6930 ( .C1(EBX_REG_13__SCAN_IN), .C2(n5969), .A(n5921), .B(n5867), 
        .ZN(n5871) );
  OAI22_X1 U6931 ( .A1(n6007), .A2(n5916), .B1(n5868), .B2(n5963), .ZN(n5869)
         );
  INV_X1 U6932 ( .A(n5869), .ZN(n5870) );
  NAND3_X1 U6933 ( .A1(n5872), .A2(n5871), .A3(n5870), .ZN(U2814) );
  OAI22_X1 U6934 ( .A1(n5962), .A2(n5874), .B1(n6524), .B2(n5873), .ZN(n5879)
         );
  INV_X1 U6935 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5877) );
  NAND3_X1 U6936 ( .A1(n5924), .A2(n6524), .A3(n5875), .ZN(n5876) );
  OAI211_X1 U6937 ( .C1(n5959), .C2(n5877), .A(n5941), .B(n5876), .ZN(n5878)
         );
  AOI211_X1 U6938 ( .C1(EBX_REG_12__SCAN_IN), .C2(n5969), .A(n5879), .B(n5878), 
        .ZN(n5884) );
  AOI22_X1 U6939 ( .A1(n5882), .A2(n5881), .B1(n5880), .B2(n5945), .ZN(n5883)
         );
  NAND2_X1 U6940 ( .A1(n5884), .A2(n5883), .ZN(U2815) );
  AOI221_X1 U6941 ( .B1(REIP_REG_10__SCAN_IN), .B2(REIP_REG_9__SCAN_IN), .C1(
        n5177), .C2(n5886), .A(n5885), .ZN(n5891) );
  INV_X1 U6942 ( .A(n5887), .ZN(n5904) );
  AOI22_X1 U6943 ( .A1(PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n5913), .B1(
        REIP_REG_10__SCAN_IN), .B2(n5904), .ZN(n5888) );
  OAI211_X1 U6944 ( .C1(n5962), .C2(n5889), .A(n5888), .B(n5941), .ZN(n5890)
         );
  AOI211_X1 U6945 ( .C1(EBX_REG_10__SCAN_IN), .C2(n5969), .A(n5891), .B(n5890), 
        .ZN(n5897) );
  INV_X1 U6946 ( .A(n5892), .ZN(n5893) );
  OAI22_X1 U6947 ( .A1(n5894), .A2(n5916), .B1(n5963), .B2(n5893), .ZN(n5895)
         );
  INV_X1 U6948 ( .A(n5895), .ZN(n5896) );
  NAND2_X1 U6949 ( .A1(n5897), .A2(n5896), .ZN(U2817) );
  NOR2_X1 U6950 ( .A1(n5962), .A2(n5898), .ZN(n5899) );
  AOI211_X1 U6951 ( .C1(n5913), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n5921), 
        .B(n5899), .ZN(n5900) );
  OAI21_X1 U6952 ( .B1(n5901), .B2(n5916), .A(n5900), .ZN(n5902) );
  AOI21_X1 U6953 ( .B1(n5903), .B2(n5945), .A(n5902), .ZN(n5907) );
  OAI21_X1 U6954 ( .B1(REIP_REG_8__SCAN_IN), .B2(n5905), .A(n5904), .ZN(n5906)
         );
  OAI211_X1 U6955 ( .C1(n5909), .C2(n5908), .A(n5907), .B(n5906), .ZN(U2819)
         );
  AOI22_X1 U6956 ( .A1(EBX_REG_7__SCAN_IN), .A2(n5969), .B1(n5926), .B2(n5910), 
        .ZN(n5923) );
  AOI221_X1 U6957 ( .B1(REIP_REG_7__SCAN_IN), .B2(REIP_REG_6__SCAN_IN), .C1(
        n5912), .C2(n6515), .A(n5911), .ZN(n5920) );
  AOI22_X1 U6958 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n5913), .B1(
        REIP_REG_7__SCAN_IN), .B2(n5933), .ZN(n5914) );
  INV_X1 U6959 ( .A(n5914), .ZN(n5919) );
  OAI22_X1 U6960 ( .A1(n5917), .A2(n5916), .B1(n5915), .B2(n5963), .ZN(n5918)
         );
  NOR4_X1 U6961 ( .A1(n5921), .A2(n5920), .A3(n5919), .A4(n5918), .ZN(n5922)
         );
  NAND2_X1 U6962 ( .A1(n5923), .A2(n5922), .ZN(U2820) );
  NAND4_X1 U6963 ( .A1(n5924), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .A4(REIP_REG_1__SCAN_IN), .ZN(n5955) );
  OAI21_X1 U6964 ( .B1(n5955), .B2(n5954), .A(n6513), .ZN(n5932) );
  INV_X1 U6965 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5928) );
  AOI22_X1 U6966 ( .A1(EBX_REG_5__SCAN_IN), .A2(n5969), .B1(n5926), .B2(n5925), 
        .ZN(n5927) );
  OAI211_X1 U6967 ( .C1(n5959), .C2(n5928), .A(n5927), .B(n5941), .ZN(n5931)
         );
  NOR2_X1 U6968 ( .A1(n5929), .A2(n5965), .ZN(n5930) );
  AOI211_X1 U6969 ( .C1(n5933), .C2(n5932), .A(n5931), .B(n5930), .ZN(n5934)
         );
  OAI21_X1 U6970 ( .B1(n5935), .B2(n5963), .A(n5934), .ZN(U2822) );
  OAI21_X1 U6971 ( .B1(n5938), .B2(n5937), .A(n5936), .ZN(n5972) );
  AOI22_X1 U6972 ( .A1(EBX_REG_4__SCAN_IN), .A2(n5969), .B1(n5940), .B2(n5939), 
        .ZN(n5942) );
  OAI211_X1 U6973 ( .C1(n5959), .C2(n5943), .A(n5942), .B(n5941), .ZN(n5952)
         );
  INV_X1 U6974 ( .A(n5944), .ZN(n5948) );
  INV_X1 U6975 ( .A(n5965), .ZN(n5947) );
  AOI22_X1 U6976 ( .A1(n5948), .A2(n5947), .B1(n5946), .B2(n5945), .ZN(n5949)
         );
  OAI21_X1 U6977 ( .B1(n5962), .B2(n5950), .A(n5949), .ZN(n5951) );
  NOR2_X1 U6978 ( .A1(n5952), .A2(n5951), .ZN(n5953) );
  OAI221_X1 U6979 ( .B1(REIP_REG_4__SCAN_IN), .B2(n5955), .C1(n5954), .C2(
        n5972), .A(n5953), .ZN(U2823) );
  NAND2_X1 U6980 ( .A1(n5956), .A2(REIP_REG_2__SCAN_IN), .ZN(n5971) );
  INV_X1 U6981 ( .A(n5957), .ZN(n5961) );
  INV_X1 U6982 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5958) );
  OAI222_X1 U6983 ( .A1(n5962), .A2(n5961), .B1(n5960), .B2(n6367), .C1(n5959), 
        .C2(n5958), .ZN(n5968) );
  OAI22_X1 U6984 ( .A1(n5966), .A2(n5965), .B1(n5964), .B2(n5963), .ZN(n5967)
         );
  AOI211_X1 U6985 ( .C1(EBX_REG_3__SCAN_IN), .C2(n5969), .A(n5968), .B(n5967), 
        .ZN(n5970) );
  OAI221_X1 U6986 ( .B1(n5972), .B2(n6510), .C1(n5972), .C2(n5971), .A(n5970), 
        .ZN(U2824) );
  AOI22_X1 U6987 ( .A1(n5996), .A2(n4196), .B1(n5977), .B2(n5973), .ZN(n5974)
         );
  OAI21_X1 U6988 ( .B1(n5988), .B2(n5975), .A(n5974), .ZN(U2842) );
  INV_X1 U6989 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5980) );
  AOI22_X1 U6990 ( .A1(n5978), .A2(n4196), .B1(n5977), .B2(n5976), .ZN(n5979)
         );
  OAI21_X1 U6991 ( .B1(n5988), .B2(n5980), .A(n5979), .ZN(U2844) );
  INV_X1 U6992 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5987) );
  INV_X1 U6993 ( .A(n5981), .ZN(n5982) );
  OAI22_X1 U6994 ( .A1(n6007), .A2(n5984), .B1(n5983), .B2(n5982), .ZN(n5985)
         );
  INV_X1 U6995 ( .A(n5985), .ZN(n5986) );
  OAI21_X1 U6996 ( .B1(n5988), .B2(n5987), .A(n5986), .ZN(U2846) );
  OAI22_X1 U6997 ( .A1(n5990), .A2(n6012), .B1(n6000), .B2(n5989), .ZN(n5991)
         );
  INV_X1 U6998 ( .A(n5991), .ZN(n5993) );
  AOI22_X1 U6999 ( .A1(n6004), .A2(DATAI_2_), .B1(n6003), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7000 ( .A1(n5993), .A2(n5992), .ZN(U2873) );
  AOI22_X1 U7001 ( .A1(n5996), .A2(n5995), .B1(n5994), .B2(DATAI_17_), .ZN(
        n5998) );
  AOI22_X1 U7002 ( .A1(n6004), .A2(DATAI_1_), .B1(n6003), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U7003 ( .A1(n5998), .A2(n5997), .ZN(U2874) );
  OAI22_X1 U7004 ( .A1(n6001), .A2(n6012), .B1(n6000), .B2(n5999), .ZN(n6002)
         );
  INV_X1 U7005 ( .A(n6002), .ZN(n6006) );
  AOI22_X1 U7006 ( .A1(n6004), .A2(DATAI_0_), .B1(n6003), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U7007 ( .A1(n6006), .A2(n6005), .ZN(U2875) );
  INV_X1 U7008 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6114) );
  OAI22_X1 U7009 ( .A1(n6007), .A2(n6012), .B1(n6758), .B2(n6010), .ZN(n6008)
         );
  INV_X1 U7010 ( .A(n6008), .ZN(n6009) );
  OAI21_X1 U7011 ( .B1(n6114), .B2(n6011), .A(n6009), .ZN(U2878) );
  INV_X1 U7012 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6076) );
  INV_X1 U7013 ( .A(DATAI_0_), .ZN(n6656) );
  OAI222_X1 U7014 ( .A1(n6143), .A2(n6012), .B1(n6011), .B2(n6076), .C1(n6010), 
        .C2(n6656), .ZN(U2891) );
  INV_X1 U7015 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6122) );
  AOI22_X1 U7016 ( .A1(n6031), .A2(LWORD_REG_15__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6014) );
  OAI21_X1 U7017 ( .B1(n6122), .B2(n6033), .A(n6014), .ZN(U2908) );
  INV_X1 U7018 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6117) );
  AOI22_X1 U7019 ( .A1(n6031), .A2(LWORD_REG_14__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6015) );
  OAI21_X1 U7020 ( .B1(n6117), .B2(n6033), .A(n6015), .ZN(U2909) );
  AOI22_X1 U7021 ( .A1(n6031), .A2(LWORD_REG_13__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6016) );
  OAI21_X1 U7022 ( .B1(n6114), .B2(n6033), .A(n6016), .ZN(U2910) );
  AOI22_X1 U7023 ( .A1(n6031), .A2(LWORD_REG_12__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6017) );
  OAI21_X1 U7024 ( .B1(n5169), .B2(n6033), .A(n6017), .ZN(U2911) );
  INV_X1 U7025 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6109) );
  AOI22_X1 U7026 ( .A1(n6031), .A2(LWORD_REG_11__SCAN_IN), .B1(n6024), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6018) );
  OAI21_X1 U7027 ( .B1(n6109), .B2(n6033), .A(n6018), .ZN(U2912) );
  INV_X1 U7028 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6106) );
  AOI22_X1 U7029 ( .A1(n6031), .A2(LWORD_REG_10__SCAN_IN), .B1(n6024), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6019) );
  OAI21_X1 U7030 ( .B1(n6106), .B2(n6033), .A(n6019), .ZN(U2913) );
  AOI22_X1 U7031 ( .A1(n6031), .A2(LWORD_REG_9__SCAN_IN), .B1(n6024), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6020) );
  OAI21_X1 U7032 ( .B1(n6103), .B2(n6033), .A(n6020), .ZN(U2914) );
  AOI22_X1 U7033 ( .A1(n6031), .A2(LWORD_REG_8__SCAN_IN), .B1(n6024), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6021) );
  OAI21_X1 U7034 ( .B1(n6100), .B2(n6033), .A(n6021), .ZN(U2915) );
  AOI22_X1 U7035 ( .A1(n6031), .A2(LWORD_REG_7__SCAN_IN), .B1(n6024), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6022) );
  OAI21_X1 U7036 ( .B1(n3755), .B2(n6033), .A(n6022), .ZN(U2916) );
  AOI22_X1 U7037 ( .A1(n6031), .A2(LWORD_REG_6__SCAN_IN), .B1(n6024), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6023) );
  OAI21_X1 U7038 ( .B1(n6094), .B2(n6033), .A(n6023), .ZN(U2917) );
  AOI22_X1 U7039 ( .A1(n6031), .A2(LWORD_REG_5__SCAN_IN), .B1(n6024), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6025) );
  OAI21_X1 U7040 ( .B1(n6091), .B2(n6033), .A(n6025), .ZN(U2918) );
  AOI22_X1 U7041 ( .A1(n6031), .A2(LWORD_REG_4__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6026) );
  OAI21_X1 U7042 ( .B1(n6088), .B2(n6033), .A(n6026), .ZN(U2919) );
  AOI22_X1 U7043 ( .A1(n6031), .A2(LWORD_REG_3__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6027) );
  OAI21_X1 U7044 ( .B1(n6085), .B2(n6033), .A(n6027), .ZN(U2920) );
  AOI22_X1 U7045 ( .A1(n6031), .A2(LWORD_REG_2__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6028) );
  OAI21_X1 U7046 ( .B1(n6082), .B2(n6033), .A(n6028), .ZN(U2921) );
  AOI22_X1 U7047 ( .A1(n6031), .A2(LWORD_REG_1__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6029) );
  OAI21_X1 U7048 ( .B1(n6079), .B2(n6033), .A(n6029), .ZN(U2922) );
  AOI22_X1 U7049 ( .A1(n6031), .A2(LWORD_REG_0__SCAN_IN), .B1(n6030), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6032) );
  OAI21_X1 U7050 ( .B1(n6076), .B2(n6033), .A(n6032), .ZN(U2923) );
  INV_X1 U7051 ( .A(n6034), .ZN(n6465) );
  NAND2_X2 U7052 ( .A1(n6035), .A2(n6465), .ZN(n6121) );
  OAI21_X1 U7053 ( .B1(n6037), .B2(n6761), .A(n6036), .ZN(n6059) );
  NOR2_X1 U7054 ( .A1(n6118), .A2(n6656), .ZN(n6074) );
  AOI21_X1 U7055 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n6059), .A(n6074), .ZN(n6038) );
  OAI21_X1 U7056 ( .B1(n6039), .B2(n6121), .A(n6038), .ZN(U2924) );
  NOR2_X1 U7057 ( .A1(n6118), .A2(n6714), .ZN(n6077) );
  AOI21_X1 U7058 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n6059), .A(n6077), .ZN(n6040) );
  OAI21_X1 U7059 ( .B1(n6041), .B2(n6121), .A(n6040), .ZN(U2925) );
  NOR2_X1 U7060 ( .A1(n6118), .A2(n6618), .ZN(n6080) );
  AOI21_X1 U7061 ( .B1(UWORD_REG_2__SCAN_IN), .B2(n6059), .A(n6080), .ZN(n6042) );
  OAI21_X1 U7062 ( .B1(n6043), .B2(n6121), .A(n6042), .ZN(U2926) );
  NOR2_X1 U7063 ( .A1(n6118), .A2(n6754), .ZN(n6083) );
  AOI21_X1 U7064 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n6059), .A(n6083), .ZN(n6044) );
  OAI21_X1 U7065 ( .B1(n6045), .B2(n6121), .A(n6044), .ZN(U2927) );
  NOR2_X1 U7066 ( .A1(n6118), .A2(n6740), .ZN(n6086) );
  AOI21_X1 U7067 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n6059), .A(n6086), .ZN(n6046) );
  OAI21_X1 U7068 ( .B1(n6047), .B2(n6121), .A(n6046), .ZN(U2928) );
  INV_X1 U7069 ( .A(DATAI_5_), .ZN(n6048) );
  NOR2_X1 U7070 ( .A1(n6118), .A2(n6048), .ZN(n6089) );
  AOI21_X1 U7071 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n6059), .A(n6089), .ZN(n6049) );
  OAI21_X1 U7072 ( .B1(n6050), .B2(n6121), .A(n6049), .ZN(U2929) );
  NOR2_X1 U7073 ( .A1(n6118), .A2(n6663), .ZN(n6092) );
  AOI21_X1 U7074 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n6059), .A(n6092), .ZN(n6051) );
  OAI21_X1 U7075 ( .B1(n6052), .B2(n6121), .A(n6051), .ZN(U2930) );
  NOR2_X1 U7076 ( .A1(n6118), .A2(n6719), .ZN(n6095) );
  AOI21_X1 U7077 ( .B1(UWORD_REG_7__SCAN_IN), .B2(n6059), .A(n6095), .ZN(n6053) );
  OAI21_X1 U7078 ( .B1(n6054), .B2(n6121), .A(n6053), .ZN(U2931) );
  NOR2_X1 U7079 ( .A1(n6118), .A2(n6757), .ZN(n6097) );
  AOI21_X1 U7080 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6059), .A(n6097), .ZN(n6055) );
  OAI21_X1 U7081 ( .B1(n6056), .B2(n6121), .A(n6055), .ZN(U2932) );
  NOR2_X1 U7082 ( .A1(n6118), .A2(n5057), .ZN(n6101) );
  AOI21_X1 U7083 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6098), .A(n6101), .ZN(n6057) );
  OAI21_X1 U7084 ( .B1(n6058), .B2(n6121), .A(n6057), .ZN(U2933) );
  INV_X1 U7085 ( .A(DATAI_10_), .ZN(n6060) );
  NOR2_X1 U7086 ( .A1(n6118), .A2(n6060), .ZN(n6104) );
  AOI21_X1 U7087 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6098), .A(n6104), .ZN(
        n6061) );
  OAI21_X1 U7088 ( .B1(n6062), .B2(n6121), .A(n6061), .ZN(U2934) );
  INV_X1 U7089 ( .A(DATAI_11_), .ZN(n6063) );
  NOR2_X1 U7090 ( .A1(n6118), .A2(n6063), .ZN(n6107) );
  AOI21_X1 U7091 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6098), .A(n6107), .ZN(
        n6064) );
  OAI21_X1 U7092 ( .B1(n6065), .B2(n6121), .A(n6064), .ZN(U2935) );
  NOR2_X1 U7093 ( .A1(n6118), .A2(n6066), .ZN(n6110) );
  AOI21_X1 U7094 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6098), .A(n6110), .ZN(
        n6067) );
  OAI21_X1 U7095 ( .B1(n6068), .B2(n6121), .A(n6067), .ZN(U2936) );
  NOR2_X1 U7096 ( .A1(n6118), .A2(n6758), .ZN(n6112) );
  AOI21_X1 U7097 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6098), .A(n6112), .ZN(
        n6069) );
  OAI21_X1 U7098 ( .B1(n6070), .B2(n6121), .A(n6069), .ZN(U2937) );
  INV_X1 U7099 ( .A(DATAI_14_), .ZN(n6071) );
  NOR2_X1 U7100 ( .A1(n6118), .A2(n6071), .ZN(n6115) );
  AOI21_X1 U7101 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6098), .A(n6115), .ZN(
        n6072) );
  OAI21_X1 U7102 ( .B1(n6073), .B2(n6121), .A(n6072), .ZN(U2938) );
  AOI21_X1 U7103 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n6098), .A(n6074), .ZN(n6075) );
  OAI21_X1 U7104 ( .B1(n6076), .B2(n6121), .A(n6075), .ZN(U2939) );
  AOI21_X1 U7105 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n6098), .A(n6077), .ZN(n6078) );
  OAI21_X1 U7106 ( .B1(n6079), .B2(n6121), .A(n6078), .ZN(U2940) );
  AOI21_X1 U7107 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n6098), .A(n6080), .ZN(n6081) );
  OAI21_X1 U7108 ( .B1(n6082), .B2(n6121), .A(n6081), .ZN(U2941) );
  AOI21_X1 U7109 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n6098), .A(n6083), .ZN(n6084) );
  OAI21_X1 U7110 ( .B1(n6085), .B2(n6121), .A(n6084), .ZN(U2942) );
  AOI21_X1 U7111 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n6098), .A(n6086), .ZN(n6087) );
  OAI21_X1 U7112 ( .B1(n6088), .B2(n6121), .A(n6087), .ZN(U2943) );
  AOI21_X1 U7113 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n6098), .A(n6089), .ZN(n6090) );
  OAI21_X1 U7114 ( .B1(n6091), .B2(n6121), .A(n6090), .ZN(U2944) );
  AOI21_X1 U7115 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n6098), .A(n6092), .ZN(n6093) );
  OAI21_X1 U7116 ( .B1(n6094), .B2(n6121), .A(n6093), .ZN(U2945) );
  AOI21_X1 U7117 ( .B1(LWORD_REG_7__SCAN_IN), .B2(n6098), .A(n6095), .ZN(n6096) );
  OAI21_X1 U7118 ( .B1(n3755), .B2(n6121), .A(n6096), .ZN(U2946) );
  AOI21_X1 U7119 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6098), .A(n6097), .ZN(n6099) );
  OAI21_X1 U7120 ( .B1(n6100), .B2(n6121), .A(n6099), .ZN(U2947) );
  AOI21_X1 U7121 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6098), .A(n6101), .ZN(n6102) );
  OAI21_X1 U7122 ( .B1(n6103), .B2(n6121), .A(n6102), .ZN(U2948) );
  AOI21_X1 U7123 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6098), .A(n6104), .ZN(
        n6105) );
  OAI21_X1 U7124 ( .B1(n6106), .B2(n6121), .A(n6105), .ZN(U2949) );
  AOI21_X1 U7125 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6098), .A(n6107), .ZN(
        n6108) );
  OAI21_X1 U7126 ( .B1(n6109), .B2(n6121), .A(n6108), .ZN(U2950) );
  AOI21_X1 U7127 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6098), .A(n6110), .ZN(
        n6111) );
  OAI21_X1 U7128 ( .B1(n5169), .B2(n6121), .A(n6111), .ZN(U2951) );
  AOI21_X1 U7129 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n6098), .A(n6112), .ZN(
        n6113) );
  OAI21_X1 U7130 ( .B1(n6114), .B2(n6121), .A(n6113), .ZN(U2952) );
  AOI21_X1 U7131 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6059), .A(n6115), .ZN(
        n6116) );
  OAI21_X1 U7132 ( .B1(n6117), .B2(n6121), .A(n6116), .ZN(U2953) );
  INV_X1 U7133 ( .A(n6118), .ZN(n6119) );
  AOI22_X1 U7134 ( .A1(n6119), .A2(DATAI_15_), .B1(n6059), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n6120) );
  OAI21_X1 U7135 ( .B1(n6122), .B2(n6121), .A(n6120), .ZN(U2954) );
  AOI22_X1 U7136 ( .A1(n6159), .A2(REIP_REG_2__SCAN_IN), .B1(n6139), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7137 ( .A1(n6124), .A2(n6123), .ZN(n6125) );
  XOR2_X1 U7138 ( .A(n6126), .B(n6125), .Z(n6165) );
  AOI22_X1 U7139 ( .A1(n6165), .A2(n6129), .B1(n6128), .B2(n6127), .ZN(n6130)
         );
  OAI211_X1 U7140 ( .C1(n6133), .C2(n6132), .A(n6131), .B(n6130), .ZN(U2984)
         );
  OAI22_X1 U7141 ( .A1(n6136), .A2(n6135), .B1(n6134), .B2(n6576), .ZN(n6137)
         );
  INV_X1 U7142 ( .A(n6137), .ZN(n6141) );
  OAI21_X1 U7143 ( .B1(n6139), .B2(n6138), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6140) );
  OAI211_X1 U7144 ( .C1(n6143), .C2(n6142), .A(n6141), .B(n6140), .ZN(U2986)
         );
  AOI21_X1 U7145 ( .B1(n6145), .B2(n6161), .A(n6144), .ZN(n6149) );
  AOI22_X1 U7146 ( .A1(n6147), .A2(n6166), .B1(n6146), .B2(n6151), .ZN(n6148)
         );
  OAI211_X1 U7147 ( .C1(n6151), .C2(n6150), .A(n6149), .B(n6148), .ZN(U3007)
         );
  AOI21_X1 U7148 ( .B1(n6153), .B2(n6161), .A(n6152), .ZN(n6157) );
  AOI22_X1 U7149 ( .A1(n6155), .A2(n6166), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6154), .ZN(n6156) );
  OAI211_X1 U7150 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6158), .A(n6157), 
        .B(n6156), .ZN(U3009) );
  AOI22_X1 U7151 ( .A1(n6161), .A2(n6160), .B1(n6159), .B2(REIP_REG_2__SCAN_IN), .ZN(n6173) );
  NAND3_X1 U7152 ( .A1(n6162), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7153 ( .A1(n6164), .A2(n6163), .ZN(n6167) );
  AOI22_X1 U7154 ( .A1(n6167), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6166), 
        .B2(n6165), .ZN(n6172) );
  NAND3_X1 U7155 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6169), .A3(n6168), 
        .ZN(n6170) );
  NAND4_X1 U7156 ( .A1(n6173), .A2(n6172), .A3(n6171), .A4(n6170), .ZN(U3016)
         );
  INV_X1 U7157 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6451) );
  NOR2_X1 U7158 ( .A1(n6451), .A2(n6174), .ZN(U3019) );
  INV_X1 U7159 ( .A(n6175), .ZN(n6176) );
  NOR2_X1 U7160 ( .A1(n6306), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6207)
         );
  AOI21_X1 U7161 ( .B1(n6176), .B2(n6314), .A(n6207), .ZN(n6181) );
  NOR2_X1 U7162 ( .A1(n6181), .A2(n6374), .ZN(n6177) );
  AOI22_X1 U7163 ( .A1(n6208), .A2(n6227), .B1(n6370), .B2(n6207), .ZN(n6187)
         );
  NOR3_X1 U7164 ( .A1(n6180), .A2(n6179), .A3(n6311), .ZN(n6185) );
  NAND2_X1 U7165 ( .A1(n6181), .A2(n6310), .ZN(n6184) );
  AOI21_X1 U7166 ( .B1(n6374), .B2(n6182), .A(n6316), .ZN(n6183) );
  OAI21_X1 U7167 ( .B1(n6185), .B2(n6184), .A(n6183), .ZN(n6210) );
  AOI22_X1 U7168 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6210), .B1(n6381), 
        .B2(n6209), .ZN(n6186) );
  OAI211_X1 U7169 ( .C1(n6214), .C2(n6188), .A(n6187), .B(n6186), .ZN(U3044)
         );
  AOI22_X1 U7170 ( .A1(n6208), .A2(n6230), .B1(n6385), .B2(n6207), .ZN(n6190)
         );
  AOI22_X1 U7171 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6210), .B1(n6387), 
        .B2(n6209), .ZN(n6189) );
  OAI211_X1 U7172 ( .C1(n6214), .C2(n6191), .A(n6190), .B(n6189), .ZN(U3045)
         );
  AOI22_X1 U7173 ( .A1(n6208), .A2(n6233), .B1(n6391), .B2(n6207), .ZN(n6193)
         );
  AOI22_X1 U7174 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6210), .B1(n6393), 
        .B2(n6209), .ZN(n6192) );
  OAI211_X1 U7175 ( .C1(n6214), .C2(n6194), .A(n6193), .B(n6192), .ZN(U3046)
         );
  AOI22_X1 U7176 ( .A1(n6208), .A2(n6236), .B1(n6397), .B2(n6207), .ZN(n6196)
         );
  AOI22_X1 U7177 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6210), .B1(n6399), 
        .B2(n6209), .ZN(n6195) );
  OAI211_X1 U7178 ( .C1(n6214), .C2(n6197), .A(n6196), .B(n6195), .ZN(U3047)
         );
  AOI22_X1 U7179 ( .A1(n6208), .A2(n6239), .B1(n6403), .B2(n6207), .ZN(n6199)
         );
  AOI22_X1 U7180 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6210), .B1(n6405), 
        .B2(n6209), .ZN(n6198) );
  OAI211_X1 U7181 ( .C1(n6214), .C2(n6200), .A(n6199), .B(n6198), .ZN(U3048)
         );
  AOI22_X1 U7182 ( .A1(n6208), .A2(n6242), .B1(n6409), .B2(n6207), .ZN(n6202)
         );
  AOI22_X1 U7183 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6210), .B1(n6411), 
        .B2(n6209), .ZN(n6201) );
  OAI211_X1 U7184 ( .C1(n6214), .C2(n6203), .A(n6202), .B(n6201), .ZN(U3049)
         );
  AOI22_X1 U7185 ( .A1(n6208), .A2(n6245), .B1(n6415), .B2(n6207), .ZN(n6205)
         );
  AOI22_X1 U7186 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6210), .B1(n6417), 
        .B2(n6209), .ZN(n6204) );
  OAI211_X1 U7187 ( .C1(n6214), .C2(n6206), .A(n6205), .B(n6204), .ZN(U3050)
         );
  AOI22_X1 U7188 ( .A1(n6208), .A2(n6250), .B1(n6422), .B2(n6207), .ZN(n6212)
         );
  AOI22_X1 U7189 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6210), .B1(n6426), 
        .B2(n6209), .ZN(n6211) );
  OAI211_X1 U7190 ( .C1(n6214), .C2(n6213), .A(n6212), .B(n6211), .ZN(U3051)
         );
  INV_X1 U7191 ( .A(n6216), .ZN(n6217) );
  OAI22_X1 U7192 ( .A1(n6219), .A2(n6218), .B1(n6217), .B2(n6365), .ZN(n6249)
         );
  NAND2_X1 U7193 ( .A1(n6369), .A2(n6262), .ZN(n6224) );
  INV_X1 U7194 ( .A(n6224), .ZN(n6248) );
  AOI22_X1 U7195 ( .A1(n6371), .A2(n6249), .B1(n6370), .B2(n6248), .ZN(n6229)
         );
  INV_X1 U7196 ( .A(n6251), .ZN(n6220) );
  AOI21_X1 U7197 ( .B1(n6220), .B2(n6287), .A(n6723), .ZN(n6222) );
  NOR2_X1 U7198 ( .A1(n6221), .A2(n6375), .ZN(n6258) );
  NOR2_X1 U7199 ( .A1(n6222), .A2(n6258), .ZN(n6223) );
  AOI22_X1 U7200 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6224), .B1(n6310), .B2(
        n6223), .ZN(n6226) );
  NAND3_X1 U7201 ( .A1(n6446), .A2(n6226), .A3(n6225), .ZN(n6252) );
  AOI22_X1 U7202 ( .A1(n6252), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6227), 
        .B2(n6251), .ZN(n6228) );
  OAI211_X1 U7203 ( .C1(n6324), .C2(n6287), .A(n6229), .B(n6228), .ZN(U3068)
         );
  AOI22_X1 U7204 ( .A1(n6386), .A2(n6249), .B1(n6385), .B2(n6248), .ZN(n6232)
         );
  AOI22_X1 U7205 ( .A1(n6252), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6251), 
        .B2(n6230), .ZN(n6231) );
  OAI211_X1 U7206 ( .C1(n6329), .C2(n6287), .A(n6232), .B(n6231), .ZN(U3069)
         );
  AOI22_X1 U7207 ( .A1(n6392), .A2(n6249), .B1(n6391), .B2(n6248), .ZN(n6235)
         );
  AOI22_X1 U7208 ( .A1(n6252), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6251), 
        .B2(n6233), .ZN(n6234) );
  OAI211_X1 U7209 ( .C1(n6334), .C2(n6287), .A(n6235), .B(n6234), .ZN(U3070)
         );
  AOI22_X1 U7210 ( .A1(n6398), .A2(n6249), .B1(n6397), .B2(n6248), .ZN(n6238)
         );
  AOI22_X1 U7211 ( .A1(n6252), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6251), 
        .B2(n6236), .ZN(n6237) );
  OAI211_X1 U7212 ( .C1(n6336), .C2(n6287), .A(n6238), .B(n6237), .ZN(U3071)
         );
  AOI22_X1 U7213 ( .A1(n6404), .A2(n6249), .B1(n6403), .B2(n6248), .ZN(n6241)
         );
  AOI22_X1 U7214 ( .A1(n6252), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6251), 
        .B2(n6239), .ZN(n6240) );
  OAI211_X1 U7215 ( .C1(n6344), .C2(n6287), .A(n6241), .B(n6240), .ZN(U3072)
         );
  AOI22_X1 U7216 ( .A1(n6410), .A2(n6249), .B1(n6409), .B2(n6248), .ZN(n6244)
         );
  AOI22_X1 U7217 ( .A1(n6252), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6251), 
        .B2(n6242), .ZN(n6243) );
  OAI211_X1 U7218 ( .C1(n6346), .C2(n6287), .A(n6244), .B(n6243), .ZN(U3073)
         );
  AOI22_X1 U7219 ( .A1(n6416), .A2(n6249), .B1(n6415), .B2(n6248), .ZN(n6247)
         );
  AOI22_X1 U7220 ( .A1(n6252), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6251), 
        .B2(n6245), .ZN(n6246) );
  OAI211_X1 U7221 ( .C1(n6351), .C2(n6287), .A(n6247), .B(n6246), .ZN(U3074)
         );
  AOI22_X1 U7222 ( .A1(n6424), .A2(n6249), .B1(n6422), .B2(n6248), .ZN(n6254)
         );
  AOI22_X1 U7223 ( .A1(n6252), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6251), 
        .B2(n6250), .ZN(n6253) );
  OAI211_X1 U7224 ( .C1(n6363), .C2(n6287), .A(n6254), .B(n6253), .ZN(U3075)
         );
  INV_X1 U7225 ( .A(n6370), .ZN(n6308) );
  OAI22_X1 U7226 ( .A1(n6303), .A2(n6324), .B1(n6286), .B2(n6308), .ZN(n6255)
         );
  INV_X1 U7227 ( .A(n6255), .ZN(n6267) );
  OR2_X1 U7228 ( .A1(n6256), .A2(n6374), .ZN(n6265) );
  INV_X1 U7229 ( .A(n6265), .ZN(n6259) );
  INV_X1 U7230 ( .A(n6286), .ZN(n6257) );
  AOI21_X1 U7231 ( .B1(n6258), .B2(n6314), .A(n6257), .ZN(n6264) );
  NAND2_X1 U7232 ( .A1(n6259), .A2(n6264), .ZN(n6260) );
  OAI211_X1 U7233 ( .C1(n6262), .C2(n6310), .A(n6261), .B(n6260), .ZN(n6290)
         );
  OAI22_X1 U7234 ( .A1(n6265), .A2(n6264), .B1(n6263), .B2(n6466), .ZN(n6289)
         );
  AOI22_X1 U7235 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6290), .B1(n6371), 
        .B2(n6289), .ZN(n6266) );
  OAI211_X1 U7236 ( .C1(n6384), .C2(n6287), .A(n6267), .B(n6266), .ZN(U3076)
         );
  INV_X1 U7237 ( .A(n6385), .ZN(n6325) );
  OAI22_X1 U7238 ( .A1(n6287), .A2(n6390), .B1(n6286), .B2(n6325), .ZN(n6268)
         );
  INV_X1 U7239 ( .A(n6268), .ZN(n6270) );
  AOI22_X1 U7240 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6290), .B1(n6386), 
        .B2(n6289), .ZN(n6269) );
  OAI211_X1 U7241 ( .C1(n6329), .C2(n6303), .A(n6270), .B(n6269), .ZN(U3077)
         );
  INV_X1 U7242 ( .A(n6391), .ZN(n6330) );
  OAI22_X1 U7243 ( .A1(n6303), .A2(n6334), .B1(n6286), .B2(n6330), .ZN(n6271)
         );
  INV_X1 U7244 ( .A(n6271), .ZN(n6273) );
  AOI22_X1 U7245 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6290), .B1(n6392), 
        .B2(n6289), .ZN(n6272) );
  OAI211_X1 U7246 ( .C1(n6396), .C2(n6287), .A(n6273), .B(n6272), .ZN(U3078)
         );
  INV_X1 U7247 ( .A(n6397), .ZN(n6335) );
  OAI22_X1 U7248 ( .A1(n6287), .A2(n6402), .B1(n6286), .B2(n6335), .ZN(n6274)
         );
  INV_X1 U7249 ( .A(n6274), .ZN(n6276) );
  AOI22_X1 U7250 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6290), .B1(n6398), 
        .B2(n6289), .ZN(n6275) );
  OAI211_X1 U7251 ( .C1(n6336), .C2(n6303), .A(n6276), .B(n6275), .ZN(U3079)
         );
  INV_X1 U7252 ( .A(n6403), .ZN(n6340) );
  OAI22_X1 U7253 ( .A1(n6303), .A2(n6344), .B1(n6286), .B2(n6340), .ZN(n6277)
         );
  INV_X1 U7254 ( .A(n6277), .ZN(n6279) );
  AOI22_X1 U7255 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6290), .B1(n6404), 
        .B2(n6289), .ZN(n6278) );
  OAI211_X1 U7256 ( .C1(n6408), .C2(n6287), .A(n6279), .B(n6278), .ZN(U3080)
         );
  INV_X1 U7257 ( .A(n6409), .ZN(n6345) );
  OAI22_X1 U7258 ( .A1(n6287), .A2(n6414), .B1(n6286), .B2(n6345), .ZN(n6280)
         );
  INV_X1 U7259 ( .A(n6280), .ZN(n6282) );
  AOI22_X1 U7260 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6290), .B1(n6410), 
        .B2(n6289), .ZN(n6281) );
  OAI211_X1 U7261 ( .C1(n6346), .C2(n6303), .A(n6282), .B(n6281), .ZN(U3081)
         );
  INV_X1 U7262 ( .A(n6415), .ZN(n6350) );
  OAI22_X1 U7263 ( .A1(n6287), .A2(n6420), .B1(n6286), .B2(n6350), .ZN(n6283)
         );
  INV_X1 U7264 ( .A(n6283), .ZN(n6285) );
  AOI22_X1 U7265 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6290), .B1(n6416), 
        .B2(n6289), .ZN(n6284) );
  OAI211_X1 U7266 ( .C1(n6351), .C2(n6303), .A(n6285), .B(n6284), .ZN(U3082)
         );
  INV_X1 U7267 ( .A(n6422), .ZN(n6356) );
  OAI22_X1 U7268 ( .A1(n6287), .A2(n6431), .B1(n6286), .B2(n6356), .ZN(n6288)
         );
  INV_X1 U7269 ( .A(n6288), .ZN(n6292) );
  AOI22_X1 U7270 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6290), .B1(n6424), 
        .B2(n6289), .ZN(n6291) );
  OAI211_X1 U7271 ( .C1(n6363), .C2(n6303), .A(n6292), .B(n6291), .ZN(U3083)
         );
  AOI22_X1 U7272 ( .A1(n6386), .A2(n6298), .B1(n6385), .B2(n6297), .ZN(n6294)
         );
  AOI22_X1 U7273 ( .A1(n6300), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6299), 
        .B2(n6387), .ZN(n6293) );
  OAI211_X1 U7274 ( .C1(n6390), .C2(n6303), .A(n6294), .B(n6293), .ZN(U3085)
         );
  AOI22_X1 U7275 ( .A1(n6392), .A2(n6298), .B1(n6391), .B2(n6297), .ZN(n6296)
         );
  AOI22_X1 U7276 ( .A1(n6300), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6299), 
        .B2(n6393), .ZN(n6295) );
  OAI211_X1 U7277 ( .C1(n6396), .C2(n6303), .A(n6296), .B(n6295), .ZN(U3086)
         );
  AOI22_X1 U7278 ( .A1(n6404), .A2(n6298), .B1(n6403), .B2(n6297), .ZN(n6302)
         );
  AOI22_X1 U7279 ( .A1(n6300), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6299), 
        .B2(n6405), .ZN(n6301) );
  OAI211_X1 U7280 ( .C1(n6408), .C2(n6303), .A(n6302), .B(n6301), .ZN(U3088)
         );
  INV_X1 U7281 ( .A(n6306), .ZN(n6307) );
  NAND2_X1 U7282 ( .A1(n6307), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6355) );
  OAI22_X1 U7283 ( .A1(n6357), .A2(n6384), .B1(n6308), .B2(n6355), .ZN(n6309)
         );
  INV_X1 U7284 ( .A(n6309), .ZN(n6323) );
  OAI21_X1 U7285 ( .B1(n6312), .B2(n6311), .A(n6310), .ZN(n6321) );
  INV_X1 U7286 ( .A(n6355), .ZN(n6313) );
  AOI21_X1 U7287 ( .B1(n6315), .B2(n6314), .A(n6313), .ZN(n6320) );
  INV_X1 U7288 ( .A(n6320), .ZN(n6318) );
  AOI21_X1 U7289 ( .B1(n6374), .B2(n6319), .A(n6316), .ZN(n6317) );
  OAI21_X1 U7290 ( .B1(n6321), .B2(n6318), .A(n6317), .ZN(n6360) );
  OAI22_X1 U7291 ( .A1(n6321), .A2(n6320), .B1(n6319), .B2(n6466), .ZN(n6359)
         );
  AOI22_X1 U7292 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6360), .B1(n6371), 
        .B2(n6359), .ZN(n6322) );
  OAI211_X1 U7293 ( .C1(n6324), .C2(n6430), .A(n6323), .B(n6322), .ZN(U3108)
         );
  OAI22_X1 U7294 ( .A1(n6357), .A2(n6390), .B1(n6325), .B2(n6355), .ZN(n6326)
         );
  INV_X1 U7295 ( .A(n6326), .ZN(n6328) );
  AOI22_X1 U7296 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6360), .B1(n6386), 
        .B2(n6359), .ZN(n6327) );
  OAI211_X1 U7297 ( .C1(n6329), .C2(n6430), .A(n6328), .B(n6327), .ZN(U3109)
         );
  OAI22_X1 U7298 ( .A1(n6357), .A2(n6396), .B1(n6330), .B2(n6355), .ZN(n6331)
         );
  INV_X1 U7299 ( .A(n6331), .ZN(n6333) );
  AOI22_X1 U7300 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6360), .B1(n6392), 
        .B2(n6359), .ZN(n6332) );
  OAI211_X1 U7301 ( .C1(n6334), .C2(n6430), .A(n6333), .B(n6332), .ZN(U3110)
         );
  OAI22_X1 U7302 ( .A1(n6430), .A2(n6336), .B1(n6335), .B2(n6355), .ZN(n6337)
         );
  INV_X1 U7303 ( .A(n6337), .ZN(n6339) );
  AOI22_X1 U7304 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6360), .B1(n6398), 
        .B2(n6359), .ZN(n6338) );
  OAI211_X1 U7305 ( .C1(n6402), .C2(n6357), .A(n6339), .B(n6338), .ZN(U3111)
         );
  OAI22_X1 U7306 ( .A1(n6357), .A2(n6408), .B1(n6340), .B2(n6355), .ZN(n6341)
         );
  INV_X1 U7307 ( .A(n6341), .ZN(n6343) );
  AOI22_X1 U7308 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6360), .B1(n6404), 
        .B2(n6359), .ZN(n6342) );
  OAI211_X1 U7309 ( .C1(n6344), .C2(n6430), .A(n6343), .B(n6342), .ZN(U3112)
         );
  OAI22_X1 U7310 ( .A1(n6430), .A2(n6346), .B1(n6345), .B2(n6355), .ZN(n6347)
         );
  INV_X1 U7311 ( .A(n6347), .ZN(n6349) );
  AOI22_X1 U7312 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6360), .B1(n6410), 
        .B2(n6359), .ZN(n6348) );
  OAI211_X1 U7313 ( .C1(n6414), .C2(n6357), .A(n6349), .B(n6348), .ZN(U3113)
         );
  OAI22_X1 U7314 ( .A1(n6430), .A2(n6351), .B1(n6350), .B2(n6355), .ZN(n6352)
         );
  INV_X1 U7315 ( .A(n6352), .ZN(n6354) );
  AOI22_X1 U7316 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6360), .B1(n6416), 
        .B2(n6359), .ZN(n6353) );
  OAI211_X1 U7317 ( .C1(n6420), .C2(n6357), .A(n6354), .B(n6353), .ZN(U3114)
         );
  OAI22_X1 U7318 ( .A1(n6357), .A2(n6431), .B1(n6356), .B2(n6355), .ZN(n6358)
         );
  INV_X1 U7319 ( .A(n6358), .ZN(n6362) );
  AOI22_X1 U7320 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6360), .B1(n6424), 
        .B2(n6359), .ZN(n6361) );
  OAI211_X1 U7321 ( .C1(n6363), .C2(n6430), .A(n6362), .B(n6361), .ZN(U3115)
         );
  OAI22_X1 U7322 ( .A1(n6367), .A2(n6366), .B1(n6365), .B2(n6364), .ZN(n6423)
         );
  AND2_X1 U7323 ( .A1(n6369), .A2(n6368), .ZN(n6421) );
  AOI22_X1 U7324 ( .A1(n6371), .A2(n6423), .B1(n6370), .B2(n6421), .ZN(n6383)
         );
  AOI21_X1 U7325 ( .B1(n6430), .B2(n6372), .A(n6723), .ZN(n6373) );
  AOI211_X1 U7326 ( .C1(n6376), .C2(n6375), .A(n6374), .B(n6373), .ZN(n6380)
         );
  OAI211_X1 U7327 ( .C1(n6562), .C2(n6421), .A(n6378), .B(n6377), .ZN(n6379)
         );
  AOI22_X1 U7328 ( .A1(n6427), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n6381), 
        .B2(n6425), .ZN(n6382) );
  OAI211_X1 U7329 ( .C1(n6384), .C2(n6430), .A(n6383), .B(n6382), .ZN(U3116)
         );
  AOI22_X1 U7330 ( .A1(n6386), .A2(n6423), .B1(n6385), .B2(n6421), .ZN(n6389)
         );
  AOI22_X1 U7331 ( .A1(n6427), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n6387), 
        .B2(n6425), .ZN(n6388) );
  OAI211_X1 U7332 ( .C1(n6390), .C2(n6430), .A(n6389), .B(n6388), .ZN(U3117)
         );
  AOI22_X1 U7333 ( .A1(n6392), .A2(n6423), .B1(n6391), .B2(n6421), .ZN(n6395)
         );
  AOI22_X1 U7334 ( .A1(n6427), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n6393), 
        .B2(n6425), .ZN(n6394) );
  OAI211_X1 U7335 ( .C1(n6396), .C2(n6430), .A(n6395), .B(n6394), .ZN(U3118)
         );
  AOI22_X1 U7336 ( .A1(n6398), .A2(n6423), .B1(n6397), .B2(n6421), .ZN(n6401)
         );
  AOI22_X1 U7337 ( .A1(n6427), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n6399), 
        .B2(n6425), .ZN(n6400) );
  OAI211_X1 U7338 ( .C1(n6402), .C2(n6430), .A(n6401), .B(n6400), .ZN(U3119)
         );
  AOI22_X1 U7339 ( .A1(n6404), .A2(n6423), .B1(n6403), .B2(n6421), .ZN(n6407)
         );
  AOI22_X1 U7340 ( .A1(n6427), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n6405), 
        .B2(n6425), .ZN(n6406) );
  OAI211_X1 U7341 ( .C1(n6408), .C2(n6430), .A(n6407), .B(n6406), .ZN(U3120)
         );
  AOI22_X1 U7342 ( .A1(n6410), .A2(n6423), .B1(n6409), .B2(n6421), .ZN(n6413)
         );
  AOI22_X1 U7343 ( .A1(n6427), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n6411), 
        .B2(n6425), .ZN(n6412) );
  OAI211_X1 U7344 ( .C1(n6414), .C2(n6430), .A(n6413), .B(n6412), .ZN(U3121)
         );
  AOI22_X1 U7345 ( .A1(n6416), .A2(n6423), .B1(n6415), .B2(n6421), .ZN(n6419)
         );
  AOI22_X1 U7346 ( .A1(n6427), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6417), 
        .B2(n6425), .ZN(n6418) );
  OAI211_X1 U7347 ( .C1(n6420), .C2(n6430), .A(n6419), .B(n6418), .ZN(U3122)
         );
  AOI22_X1 U7348 ( .A1(n6424), .A2(n6423), .B1(n6422), .B2(n6421), .ZN(n6429)
         );
  AOI22_X1 U7349 ( .A1(n6427), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6426), 
        .B2(n6425), .ZN(n6428) );
  OAI211_X1 U7350 ( .C1(n6431), .C2(n6430), .A(n6429), .B(n6428), .ZN(U3123)
         );
  INV_X1 U7351 ( .A(n6432), .ZN(n6433) );
  OAI211_X1 U7352 ( .C1(n3710), .C2(n6434), .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n6433), .ZN(n6438) );
  INV_X1 U7353 ( .A(n6435), .ZN(n6436) );
  OAI211_X1 U7354 ( .C1(n6439), .C2(n6438), .A(n6437), .B(n6436), .ZN(n6441)
         );
  NAND2_X1 U7355 ( .A1(n6439), .A2(n6438), .ZN(n6440) );
  NAND2_X1 U7356 ( .A1(n6441), .A2(n6440), .ZN(n6442) );
  AND2_X1 U7357 ( .A1(n3248), .A2(n6442), .ZN(n6443) );
  OAI22_X1 U7358 ( .A1(n6444), .A2(n6443), .B1(n3248), .B2(n6442), .ZN(n6450)
         );
  INV_X1 U7359 ( .A(n6445), .ZN(n6449) );
  NAND2_X1 U7360 ( .A1(n6449), .A2(n6450), .ZN(n6447) );
  NAND2_X1 U7361 ( .A1(n6447), .A2(n6446), .ZN(n6448) );
  OAI21_X1 U7362 ( .B1(n6450), .B2(n6449), .A(n6448), .ZN(n6452) );
  NAND2_X1 U7363 ( .A1(n6452), .A2(n6451), .ZN(n6462) );
  NOR2_X1 U7364 ( .A1(n6454), .A2(n6453), .ZN(n6457) );
  OAI21_X1 U7365 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6455), 
        .ZN(n6456) );
  NAND3_X1 U7366 ( .A1(n6458), .A2(n6457), .A3(n6456), .ZN(n6459) );
  NOR2_X1 U7367 ( .A1(n6460), .A2(n6459), .ZN(n6461) );
  AOI21_X1 U7368 ( .B1(STATE2_REG_1__SCAN_IN), .B2(READY_N), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n6463) );
  AOI211_X1 U7369 ( .C1(n6465), .C2(n6464), .A(n6463), .B(n6466), .ZN(n6468)
         );
  OAI221_X1 U7370 ( .B1(n6477), .B2(n6476), .C1(n6467), .C2(n6476), .A(n6468), 
        .ZN(n6561) );
  INV_X1 U7371 ( .A(n6561), .ZN(n6479) );
  AOI21_X1 U7372 ( .B1(READY_N), .B2(n6466), .A(n6479), .ZN(n6478) );
  INV_X1 U7373 ( .A(n6467), .ZN(n6472) );
  AOI211_X1 U7374 ( .C1(n6582), .C2(n6469), .A(STATE2_REG_0__SCAN_IN), .B(
        n6468), .ZN(n6470) );
  AOI211_X1 U7375 ( .C1(n6473), .C2(n6472), .A(n6471), .B(n6470), .ZN(n6474)
         );
  OAI221_X1 U7376 ( .B1(n6476), .B2(n6478), .C1(n6476), .C2(n6475), .A(n6474), 
        .ZN(U3148) );
  NOR3_X1 U7377 ( .A1(n6488), .A2(n6478), .A3(n6477), .ZN(n6483) );
  AOI221_X1 U7378 ( .B1(READY_N), .B2(n6481), .C1(n6480), .C2(n6481), .A(n6479), .ZN(n6482) );
  OR3_X1 U7379 ( .A1(n6484), .A2(n6483), .A3(n6482), .ZN(U3149) );
  OAI211_X1 U7380 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6761), .A(n6559), .B(
        n6485), .ZN(n6487) );
  OAI21_X1 U7381 ( .B1(n6488), .B2(n6487), .A(n6486), .ZN(U3150) );
  AND2_X1 U7382 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6489), .ZN(U3151) );
  AND2_X1 U7383 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6489), .ZN(U3152) );
  AND2_X1 U7384 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6489), .ZN(U3153) );
  AND2_X1 U7385 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6489), .ZN(U3154) );
  AND2_X1 U7386 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6489), .ZN(U3155) );
  AND2_X1 U7387 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6489), .ZN(U3156) );
  AND2_X1 U7388 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6489), .ZN(U3157) );
  AND2_X1 U7389 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6489), .ZN(U3158) );
  AND2_X1 U7390 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6489), .ZN(U3159) );
  AND2_X1 U7391 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6489), .ZN(U3160) );
  AND2_X1 U7392 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6489), .ZN(U3161) );
  AND2_X1 U7393 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6489), .ZN(U3162) );
  AND2_X1 U7394 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6489), .ZN(U3163) );
  AND2_X1 U7395 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6489), .ZN(U3164) );
  AND2_X1 U7396 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6489), .ZN(U3165) );
  AND2_X1 U7397 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6489), .ZN(U3166) );
  AND2_X1 U7398 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6489), .ZN(U3167) );
  AND2_X1 U7399 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6489), .ZN(U3168) );
  AND2_X1 U7400 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6489), .ZN(U3169) );
  AND2_X1 U7401 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6489), .ZN(U3170) );
  AND2_X1 U7402 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6489), .ZN(U3171) );
  AND2_X1 U7403 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6489), .ZN(U3172) );
  AND2_X1 U7404 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6489), .ZN(U3173) );
  AND2_X1 U7405 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6489), .ZN(U3174) );
  AND2_X1 U7406 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6489), .ZN(U3175) );
  AND2_X1 U7407 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6489), .ZN(U3176) );
  AND2_X1 U7408 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6489), .ZN(U3177) );
  AND2_X1 U7409 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6489), .ZN(U3178) );
  AND2_X1 U7410 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6489), .ZN(U3179) );
  AND2_X1 U7411 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6489), .ZN(U3180) );
  NOR2_X1 U7412 ( .A1(n6506), .A2(n6496), .ZN(n6497) );
  AOI22_X1 U7413 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6505) );
  AND2_X1 U7414 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6493) );
  INV_X1 U7415 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6491) );
  INV_X1 U7416 ( .A(NA_N), .ZN(n6498) );
  AOI221_X1 U7417 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6498), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6502) );
  AOI221_X1 U7418 ( .B1(n6493), .B2(n6777), .C1(n6491), .C2(n6777), .A(n6502), 
        .ZN(n6490) );
  OAI21_X1 U7419 ( .B1(n6497), .B2(n6505), .A(n6490), .ZN(U3181) );
  NOR2_X1 U7420 ( .A1(n6500), .A2(n6491), .ZN(n6499) );
  NAND2_X1 U7421 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6492) );
  OAI21_X1 U7422 ( .B1(n6499), .B2(n6493), .A(n6492), .ZN(n6494) );
  OAI211_X1 U7423 ( .C1(n6496), .C2(n6761), .A(n6495), .B(n6494), .ZN(U3182)
         );
  AOI21_X1 U7424 ( .B1(n6499), .B2(n6498), .A(n6497), .ZN(n6504) );
  AOI221_X1 U7425 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6761), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6501) );
  AOI221_X1 U7426 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6501), .C2(HOLD), .A(n6500), .ZN(n6503) );
  OAI22_X1 U7427 ( .A1(n6505), .A2(n6504), .B1(n6503), .B2(n6502), .ZN(U3183)
         );
  NOR2_X2 U7428 ( .A1(n6506), .A2(n6777), .ZN(n6551) );
  NAND2_X1 U7429 ( .A1(n6506), .A2(n6778), .ZN(n6553) );
  INV_X1 U7430 ( .A(n6553), .ZN(n6547) );
  AOI22_X1 U7431 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6541), .ZN(n6507) );
  OAI21_X1 U7432 ( .B1(n6571), .B2(n6549), .A(n6507), .ZN(U3184) );
  AOI22_X1 U7433 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6551), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6541), .ZN(n6508) );
  OAI21_X1 U7434 ( .B1(n6510), .B2(n6553), .A(n6508), .ZN(U3185) );
  AOI22_X1 U7435 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6541), .ZN(n6509) );
  OAI21_X1 U7436 ( .B1(n6510), .B2(n6549), .A(n6509), .ZN(U3186) );
  AOI22_X1 U7437 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6551), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6541), .ZN(n6511) );
  OAI21_X1 U7438 ( .B1(n6513), .B2(n6553), .A(n6511), .ZN(U3187) );
  AOI22_X1 U7439 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6541), .ZN(n6512) );
  OAI21_X1 U7440 ( .B1(n6513), .B2(n6549), .A(n6512), .ZN(U3188) );
  AOI22_X1 U7441 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6541), .ZN(n6514) );
  OAI21_X1 U7442 ( .B1(n6515), .B2(n6549), .A(n6514), .ZN(U3189) );
  AOI22_X1 U7443 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6551), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6541), .ZN(n6516) );
  OAI21_X1 U7444 ( .B1(n6518), .B2(n6553), .A(n6516), .ZN(U3190) );
  AOI22_X1 U7445 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6541), .ZN(n6517) );
  OAI21_X1 U7446 ( .B1(n6518), .B2(n6549), .A(n6517), .ZN(U3191) );
  AOI22_X1 U7447 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6551), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6541), .ZN(n6519) );
  OAI21_X1 U7448 ( .B1(n5177), .B2(n6553), .A(n6519), .ZN(U3192) );
  AOI22_X1 U7449 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6551), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6541), .ZN(n6520) );
  OAI21_X1 U7450 ( .B1(n6522), .B2(n6553), .A(n6520), .ZN(U3193) );
  AOI22_X1 U7451 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6777), .ZN(n6521) );
  OAI21_X1 U7452 ( .B1(n6522), .B2(n6549), .A(n6521), .ZN(U3194) );
  AOI22_X1 U7453 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6541), .ZN(n6523) );
  OAI21_X1 U7454 ( .B1(n6524), .B2(n6549), .A(n6523), .ZN(U3195) );
  AOI22_X1 U7455 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6551), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6541), .ZN(n6525) );
  OAI21_X1 U7456 ( .B1(n6527), .B2(n6553), .A(n6525), .ZN(U3196) );
  AOI22_X1 U7457 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6541), .ZN(n6526) );
  OAI21_X1 U7458 ( .B1(n6527), .B2(n6549), .A(n6526), .ZN(U3197) );
  AOI22_X1 U7459 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6551), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6541), .ZN(n6528) );
  OAI21_X1 U7460 ( .B1(n6530), .B2(n6553), .A(n6528), .ZN(U3198) );
  AOI22_X1 U7461 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6541), .ZN(n6529) );
  OAI21_X1 U7462 ( .B1(n6530), .B2(n6549), .A(n6529), .ZN(U3199) );
  AOI22_X1 U7463 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6551), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6541), .ZN(n6531) );
  OAI21_X1 U7464 ( .B1(n6533), .B2(n6553), .A(n6531), .ZN(U3200) );
  AOI22_X1 U7465 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6541), .ZN(n6532) );
  OAI21_X1 U7466 ( .B1(n6533), .B2(n6549), .A(n6532), .ZN(U3201) );
  AOI22_X1 U7467 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6551), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6541), .ZN(n6534) );
  OAI21_X1 U7468 ( .B1(n6536), .B2(n6553), .A(n6534), .ZN(U3202) );
  AOI22_X1 U7469 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6541), .ZN(n6535) );
  OAI21_X1 U7470 ( .B1(n6536), .B2(n6549), .A(n6535), .ZN(U3203) );
  AOI22_X1 U7471 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6541), .ZN(n6537) );
  OAI21_X1 U7472 ( .B1(n6538), .B2(n6549), .A(n6537), .ZN(U3204) );
  AOI22_X1 U7473 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6541), .ZN(n6539) );
  OAI21_X1 U7474 ( .B1(n6634), .B2(n6549), .A(n6539), .ZN(U3205) );
  AOI22_X1 U7475 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6541), .ZN(n6540) );
  OAI21_X1 U7476 ( .B1(n6666), .B2(n6549), .A(n6540), .ZN(U3206) );
  AOI22_X1 U7477 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6541), .ZN(n6542) );
  OAI21_X1 U7478 ( .B1(n6720), .B2(n6549), .A(n6542), .ZN(U3207) );
  AOI22_X1 U7479 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6777), .ZN(n6543) );
  OAI21_X1 U7480 ( .B1(n6544), .B2(n6549), .A(n6543), .ZN(U3208) );
  AOI22_X1 U7481 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6551), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6777), .ZN(n6545) );
  OAI21_X1 U7482 ( .B1(n6649), .B2(n6553), .A(n6545), .ZN(U3209) );
  AOI22_X1 U7483 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6551), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6777), .ZN(n6546) );
  OAI21_X1 U7484 ( .B1(n6632), .B2(n6553), .A(n6546), .ZN(U3210) );
  AOI22_X1 U7485 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6777), .ZN(n6548) );
  OAI21_X1 U7486 ( .B1(n6632), .B2(n6549), .A(n6548), .ZN(U3211) );
  AOI22_X1 U7487 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6551), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6777), .ZN(n6550) );
  OAI21_X1 U7488 ( .B1(n6764), .B2(n6553), .A(n6550), .ZN(U3212) );
  AOI22_X1 U7489 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6551), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6777), .ZN(n6552) );
  OAI21_X1 U7490 ( .B1(n6554), .B2(n6553), .A(n6552), .ZN(U3213) );
  MUX2_X1 U7491 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6777), .Z(U3446) );
  MUX2_X1 U7492 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6777), .Z(U3447) );
  MUX2_X1 U7493 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6777), .Z(U3448) );
  OAI21_X1 U7494 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6558), .A(n6556), .ZN(
        n6555) );
  INV_X1 U7495 ( .A(n6555), .ZN(U3451) );
  OAI21_X1 U7496 ( .B1(n6558), .B2(n6557), .A(n6556), .ZN(U3452) );
  OAI211_X1 U7497 ( .C1(n6562), .C2(n6561), .A(n6560), .B(n6559), .ZN(U3453)
         );
  INV_X1 U7498 ( .A(n6563), .ZN(n6568) );
  INV_X1 U7499 ( .A(n6564), .ZN(n6567) );
  OAI22_X1 U7500 ( .A1(n6568), .A2(n6567), .B1(n6566), .B2(n6565), .ZN(n6570)
         );
  MUX2_X1 U7501 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6570), .S(n6569), 
        .Z(U3456) );
  AOI21_X1 U7502 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6572) );
  AOI22_X1 U7503 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6572), .B2(n6571), .ZN(n6573) );
  INV_X1 U7504 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6659) );
  AOI22_X1 U7505 ( .A1(n6574), .A2(n6573), .B1(n6659), .B2(n6577), .ZN(U3468)
         );
  INV_X1 U7506 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6665) );
  NOR2_X1 U7507 ( .A1(n6577), .A2(REIP_REG_1__SCAN_IN), .ZN(n6575) );
  AOI22_X1 U7508 ( .A1(n6665), .A2(n6577), .B1(n6576), .B2(n6575), .ZN(U3469)
         );
  INV_X1 U7509 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6745) );
  AOI22_X1 U7510 ( .A1(n6778), .A2(READREQUEST_REG_SCAN_IN), .B1(n6745), .B2(
        n6777), .ZN(U3470) );
  AOI211_X1 U7511 ( .C1(n6031), .C2(n6761), .A(n6579), .B(n6578), .ZN(n6586)
         );
  OAI211_X1 U7512 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6581), .A(n6580), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6583) );
  AOI21_X1 U7513 ( .B1(n6583), .B2(STATE2_REG_0__SCAN_IN), .A(n6582), .ZN(
        n6585) );
  NAND2_X1 U7514 ( .A1(n6586), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6584) );
  OAI21_X1 U7515 ( .B1(n6586), .B2(n6585), .A(n6584), .ZN(U3472) );
  INV_X1 U7516 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6732) );
  INV_X1 U7517 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6717) );
  AOI22_X1 U7518 ( .A1(n6778), .A2(n6732), .B1(n6717), .B2(n6777), .ZN(U3473)
         );
  AOI22_X1 U7519 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(REIP_REG_21__SCAN_IN), 
        .B2(keyinput_f61), .ZN(n6587) );
  OAI221_X1 U7520 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(REIP_REG_21__SCAN_IN), .C2(keyinput_f61), .A(n6587), .ZN(n6646) );
  AOI22_X1 U7521 ( .A1(keyinput_f36), .A2(HOLD), .B1(
        REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_f42), .ZN(n6588) );
  OAI221_X1 U7522 ( .B1(keyinput_f36), .B2(HOLD), .C1(
        REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_f42), .A(n6588), .ZN(n6645)
         );
  INV_X1 U7523 ( .A(DATAI_20_), .ZN(n6747) );
  AOI22_X1 U7524 ( .A1(DATAI_9_), .A2(keyinput_f22), .B1(n6747), .B2(
        keyinput_f11), .ZN(n6589) );
  OAI221_X1 U7525 ( .B1(DATAI_9_), .B2(keyinput_f22), .C1(n6747), .C2(
        keyinput_f11), .A(n6589), .ZN(n6599) );
  OAI22_X1 U7526 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput_f51), .B1(
        REIP_REG_25__SCAN_IN), .B2(keyinput_f57), .ZN(n6590) );
  AOI221_X1 U7527 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_f51), .C1(
        keyinput_f57), .C2(REIP_REG_25__SCAN_IN), .A(n6590), .ZN(n6597) );
  OAI22_X1 U7528 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(W_R_N_REG_SCAN_IN), 
        .B2(keyinput_f46), .ZN(n6591) );
  AOI221_X1 U7529 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(keyinput_f46), .C2(
        W_R_N_REG_SCAN_IN), .A(n6591), .ZN(n6596) );
  OAI22_X1 U7530 ( .A1(DATAI_14_), .A2(keyinput_f17), .B1(DATAI_15_), .B2(
        keyinput_f16), .ZN(n6592) );
  AOI221_X1 U7531 ( .B1(DATAI_14_), .B2(keyinput_f17), .C1(keyinput_f16), .C2(
        DATAI_15_), .A(n6592), .ZN(n6595) );
  OAI22_X1 U7532 ( .A1(DATAI_13_), .A2(keyinput_f18), .B1(keyinput_f38), .B2(
        ADS_N_REG_SCAN_IN), .ZN(n6593) );
  AOI221_X1 U7533 ( .B1(DATAI_13_), .B2(keyinput_f18), .C1(ADS_N_REG_SCAN_IN), 
        .C2(keyinput_f38), .A(n6593), .ZN(n6594) );
  NAND4_X1 U7534 ( .A1(n6597), .A2(n6596), .A3(n6595), .A4(n6594), .ZN(n6598)
         );
  AOI211_X1 U7535 ( .C1(keyinput_f0), .C2(DATAI_31_), .A(n6599), .B(n6598), 
        .ZN(n6600) );
  OAI21_X1 U7536 ( .B1(keyinput_f0), .B2(DATAI_31_), .A(n6600), .ZN(n6644) );
  AOI22_X1 U7537 ( .A1(keyinput_f40), .A2(M_IO_N_REG_SCAN_IN), .B1(
        MORE_REG_SCAN_IN), .B2(keyinput_f44), .ZN(n6601) );
  OAI221_X1 U7538 ( .B1(keyinput_f40), .B2(M_IO_N_REG_SCAN_IN), .C1(
        MORE_REG_SCAN_IN), .C2(keyinput_f44), .A(n6601), .ZN(n6608) );
  AOI22_X1 U7539 ( .A1(DATAI_23_), .A2(keyinput_f8), .B1(REIP_REG_19__SCAN_IN), 
        .B2(keyinput_f63), .ZN(n6602) );
  OAI221_X1 U7540 ( .B1(DATAI_23_), .B2(keyinput_f8), .C1(REIP_REG_19__SCAN_IN), .C2(keyinput_f63), .A(n6602), .ZN(n6607) );
  INV_X1 U7541 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6744) );
  AOI22_X1 U7542 ( .A1(DATAI_8_), .A2(keyinput_f23), .B1(n6744), .B2(
        keyinput_f39), .ZN(n6603) );
  OAI221_X1 U7543 ( .B1(DATAI_8_), .B2(keyinput_f23), .C1(n6744), .C2(
        keyinput_f39), .A(n6603), .ZN(n6606) );
  AOI22_X1 U7544 ( .A1(DATAI_22_), .A2(keyinput_f9), .B1(REIP_REG_26__SCAN_IN), 
        .B2(keyinput_f56), .ZN(n6604) );
  OAI221_X1 U7545 ( .B1(DATAI_22_), .B2(keyinput_f9), .C1(REIP_REG_26__SCAN_IN), .C2(keyinput_f56), .A(n6604), .ZN(n6605) );
  NOR4_X1 U7546 ( .A1(n6608), .A2(n6607), .A3(n6606), .A4(n6605), .ZN(n6642)
         );
  AOI22_X1 U7547 ( .A1(DATAI_7_), .A2(keyinput_f24), .B1(DATAI_29_), .B2(
        keyinput_f2), .ZN(n6609) );
  OAI221_X1 U7548 ( .B1(DATAI_7_), .B2(keyinput_f24), .C1(DATAI_29_), .C2(
        keyinput_f2), .A(n6609), .ZN(n6616) );
  AOI22_X1 U7549 ( .A1(keyinput_f33), .A2(NA_N), .B1(DATAI_4_), .B2(
        keyinput_f27), .ZN(n6610) );
  OAI221_X1 U7550 ( .B1(keyinput_f33), .B2(NA_N), .C1(DATAI_4_), .C2(
        keyinput_f27), .A(n6610), .ZN(n6615) );
  AOI22_X1 U7551 ( .A1(DATAI_12_), .A2(keyinput_f19), .B1(REIP_REG_20__SCAN_IN), .B2(keyinput_f62), .ZN(n6611) );
  OAI221_X1 U7552 ( .B1(DATAI_12_), .B2(keyinput_f19), .C1(
        REIP_REG_20__SCAN_IN), .C2(keyinput_f62), .A(n6611), .ZN(n6614) );
  AOI22_X1 U7553 ( .A1(DATAI_3_), .A2(keyinput_f28), .B1(DATAI_25_), .B2(
        keyinput_f6), .ZN(n6612) );
  OAI221_X1 U7554 ( .B1(DATAI_3_), .B2(keyinput_f28), .C1(DATAI_25_), .C2(
        keyinput_f6), .A(n6612), .ZN(n6613) );
  NOR4_X1 U7555 ( .A1(n6616), .A2(n6615), .A3(n6614), .A4(n6613), .ZN(n6641)
         );
  AOI22_X1 U7556 ( .A1(n6618), .A2(keyinput_f29), .B1(n6761), .B2(keyinput_f35), .ZN(n6617) );
  OAI221_X1 U7557 ( .B1(n6618), .B2(keyinput_f29), .C1(n6761), .C2(
        keyinput_f35), .A(n6617), .ZN(n6627) );
  AOI22_X1 U7558 ( .A1(n4502), .A2(keyinput_f12), .B1(keyinput_f15), .B2(n5999), .ZN(n6619) );
  OAI221_X1 U7559 ( .B1(n4502), .B2(keyinput_f12), .C1(n5999), .C2(
        keyinput_f15), .A(n6619), .ZN(n6626) );
  INV_X1 U7560 ( .A(keyinput_f50), .ZN(n6621) );
  AOI22_X1 U7561 ( .A1(n6764), .A2(keyinput_f52), .B1(
        BYTEENABLE_REG_3__SCAN_IN), .B2(n6621), .ZN(n6620) );
  OAI221_X1 U7562 ( .B1(n6764), .B2(keyinput_f52), .C1(n6621), .C2(
        BYTEENABLE_REG_3__SCAN_IN), .A(n6620), .ZN(n6625) );
  INV_X1 U7563 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6623) );
  AOI22_X1 U7564 ( .A1(n6623), .A2(keyinput_f37), .B1(n6723), .B2(keyinput_f43), .ZN(n6622) );
  OAI221_X1 U7565 ( .B1(n6623), .B2(keyinput_f37), .C1(n6723), .C2(
        keyinput_f43), .A(n6622), .ZN(n6624) );
  NOR4_X1 U7566 ( .A1(n6627), .A2(n6626), .A3(n6625), .A4(n6624), .ZN(n6640)
         );
  AOI22_X1 U7567 ( .A1(n5989), .A2(keyinput_f13), .B1(n6629), .B2(keyinput_f53), .ZN(n6628) );
  OAI221_X1 U7568 ( .B1(n5989), .B2(keyinput_f13), .C1(n6629), .C2(
        keyinput_f53), .A(n6628), .ZN(n6638) );
  AOI22_X1 U7569 ( .A1(n6720), .A2(keyinput_f58), .B1(keyinput_f14), .B2(n4476), .ZN(n6630) );
  OAI221_X1 U7570 ( .B1(n6720), .B2(keyinput_f58), .C1(n4476), .C2(
        keyinput_f14), .A(n6630), .ZN(n6637) );
  AOI22_X1 U7571 ( .A1(n6742), .A2(keyinput_f5), .B1(n6632), .B2(keyinput_f54), 
        .ZN(n6631) );
  OAI221_X1 U7572 ( .B1(n6742), .B2(keyinput_f5), .C1(n6632), .C2(keyinput_f54), .A(n6631), .ZN(n6636) );
  AOI22_X1 U7573 ( .A1(n6760), .A2(keyinput_f3), .B1(n6634), .B2(keyinput_f60), 
        .ZN(n6633) );
  OAI221_X1 U7574 ( .B1(n6760), .B2(keyinput_f3), .C1(n6634), .C2(keyinput_f60), .A(n6633), .ZN(n6635) );
  NOR4_X1 U7575 ( .A1(n6638), .A2(n6637), .A3(n6636), .A4(n6635), .ZN(n6639)
         );
  NAND4_X1 U7576 ( .A1(n6642), .A2(n6641), .A3(n6640), .A4(n6639), .ZN(n6643)
         );
  NOR4_X1 U7577 ( .A1(n6646), .A2(n6645), .A3(n6644), .A4(n6643), .ZN(n6677)
         );
  AOI22_X1 U7578 ( .A1(n6714), .A2(keyinput_f30), .B1(n6063), .B2(keyinput_f20), .ZN(n6647) );
  OAI221_X1 U7579 ( .B1(n6714), .B2(keyinput_f30), .C1(n6063), .C2(
        keyinput_f20), .A(n6647), .ZN(n6674) );
  AOI22_X1 U7580 ( .A1(n6048), .A2(keyinput_f26), .B1(n6649), .B2(keyinput_f55), .ZN(n6648) );
  OAI221_X1 U7581 ( .B1(n6048), .B2(keyinput_f26), .C1(n6649), .C2(
        keyinput_f55), .A(n6648), .ZN(n6673) );
  XOR2_X1 U7582 ( .A(keyinput_f34), .B(BS16_N), .Z(n6653) );
  AOI22_X1 U7583 ( .A1(n5738), .A2(keyinput_f10), .B1(keyinput_f41), .B2(n6651), .ZN(n6650) );
  OAI221_X1 U7584 ( .B1(n5738), .B2(keyinput_f10), .C1(n6651), .C2(
        keyinput_f41), .A(n6650), .ZN(n6652) );
  AOI211_X1 U7585 ( .C1(n6732), .C2(keyinput_f32), .A(n6653), .B(n6652), .ZN(
        n6654) );
  OAI21_X1 U7586 ( .B1(n6732), .B2(keyinput_f32), .A(n6654), .ZN(n6672) );
  OAI22_X1 U7587 ( .A1(n6657), .A2(keyinput_f4), .B1(n6656), .B2(keyinput_f31), 
        .ZN(n6655) );
  AOI221_X1 U7588 ( .B1(n6657), .B2(keyinput_f4), .C1(keyinput_f31), .C2(n6656), .A(n6655), .ZN(n6670) );
  OAI22_X1 U7589 ( .A1(n6660), .A2(keyinput_f45), .B1(n6659), .B2(keyinput_f49), .ZN(n6658) );
  AOI221_X1 U7590 ( .B1(n6660), .B2(keyinput_f45), .C1(keyinput_f49), .C2(
        n6659), .A(n6658), .ZN(n6669) );
  OAI22_X1 U7591 ( .A1(n6663), .A2(keyinput_f25), .B1(n6662), .B2(keyinput_f48), .ZN(n6661) );
  AOI221_X1 U7592 ( .B1(n6663), .B2(keyinput_f25), .C1(keyinput_f48), .C2(
        n6662), .A(n6661), .ZN(n6668) );
  OAI22_X1 U7593 ( .A1(n6666), .A2(keyinput_f59), .B1(n6665), .B2(keyinput_f47), .ZN(n6664) );
  AOI221_X1 U7594 ( .B1(n6666), .B2(keyinput_f59), .C1(keyinput_f47), .C2(
        n6665), .A(n6664), .ZN(n6667) );
  NAND4_X1 U7595 ( .A1(n6670), .A2(n6669), .A3(n6668), .A4(n6667), .ZN(n6671)
         );
  NOR4_X1 U7596 ( .A1(n6674), .A2(n6673), .A3(n6672), .A4(n6671), .ZN(n6676)
         );
  NOR2_X1 U7597 ( .A1(DATAI_10_), .A2(keyinput_f21), .ZN(n6675) );
  AOI221_X1 U7598 ( .B1(n6677), .B2(n6676), .C1(keyinput_f21), .C2(DATAI_10_), 
        .A(n6675), .ZN(n6776) );
  AOI22_X1 U7599 ( .A1(DATAI_24_), .A2(keyinput_g7), .B1(DATAI_29_), .B2(
        keyinput_g2), .ZN(n6678) );
  OAI221_X1 U7600 ( .B1(DATAI_24_), .B2(keyinput_g7), .C1(DATAI_29_), .C2(
        keyinput_g2), .A(n6678), .ZN(n6685) );
  AOI22_X1 U7601 ( .A1(DATAI_22_), .A2(keyinput_g9), .B1(DATAI_9_), .B2(
        keyinput_g22), .ZN(n6679) );
  OAI221_X1 U7602 ( .B1(DATAI_22_), .B2(keyinput_g9), .C1(DATAI_9_), .C2(
        keyinput_g22), .A(n6679), .ZN(n6684) );
  AOI22_X1 U7603 ( .A1(ADS_N_REG_SCAN_IN), .A2(keyinput_g38), .B1(DATAI_11_), 
        .B2(keyinput_g20), .ZN(n6680) );
  OAI221_X1 U7604 ( .B1(ADS_N_REG_SCAN_IN), .B2(keyinput_g38), .C1(DATAI_11_), 
        .C2(keyinput_g20), .A(n6680), .ZN(n6683) );
  AOI22_X1 U7605 ( .A1(DATAI_21_), .A2(keyinput_g10), .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_g60), .ZN(n6681) );
  OAI221_X1 U7606 ( .B1(DATAI_21_), .B2(keyinput_g10), .C1(
        REIP_REG_22__SCAN_IN), .C2(keyinput_g60), .A(n6681), .ZN(n6682) );
  NOR4_X1 U7607 ( .A1(n6685), .A2(n6684), .A3(n6683), .A4(n6682), .ZN(n6712)
         );
  XOR2_X1 U7608 ( .A(HOLD), .B(keyinput_g36), .Z(n6692) );
  AOI22_X1 U7609 ( .A1(DATAI_18_), .A2(keyinput_g13), .B1(REIP_REG_27__SCAN_IN), .B2(keyinput_g55), .ZN(n6686) );
  OAI221_X1 U7610 ( .B1(DATAI_18_), .B2(keyinput_g13), .C1(
        REIP_REG_27__SCAN_IN), .C2(keyinput_g55), .A(n6686), .ZN(n6691) );
  AOI22_X1 U7611 ( .A1(DATAI_5_), .A2(keyinput_g26), .B1(DATAI_12_), .B2(
        keyinput_g19), .ZN(n6687) );
  OAI221_X1 U7612 ( .B1(DATAI_5_), .B2(keyinput_g26), .C1(DATAI_12_), .C2(
        keyinput_g19), .A(n6687), .ZN(n6690) );
  AOI22_X1 U7613 ( .A1(REIP_REG_25__SCAN_IN), .A2(keyinput_g57), .B1(
        REIP_REG_28__SCAN_IN), .B2(keyinput_g54), .ZN(n6688) );
  OAI221_X1 U7614 ( .B1(REIP_REG_25__SCAN_IN), .B2(keyinput_g57), .C1(
        REIP_REG_28__SCAN_IN), .C2(keyinput_g54), .A(n6688), .ZN(n6689) );
  NOR4_X1 U7615 ( .A1(n6692), .A2(n6691), .A3(n6690), .A4(n6689), .ZN(n6711)
         );
  AOI22_X1 U7616 ( .A1(DATAI_2_), .A2(keyinput_g29), .B1(DATAI_6_), .B2(
        keyinput_g25), .ZN(n6693) );
  OAI221_X1 U7617 ( .B1(DATAI_2_), .B2(keyinput_g29), .C1(DATAI_6_), .C2(
        keyinput_g25), .A(n6693), .ZN(n6700) );
  AOI22_X1 U7618 ( .A1(NA_N), .A2(keyinput_g33), .B1(REIP_REG_20__SCAN_IN), 
        .B2(keyinput_g62), .ZN(n6694) );
  OAI221_X1 U7619 ( .B1(NA_N), .B2(keyinput_g33), .C1(REIP_REG_20__SCAN_IN), 
        .C2(keyinput_g62), .A(n6694), .ZN(n6699) );
  AOI22_X1 U7620 ( .A1(DATAI_16_), .A2(keyinput_g15), .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_g51), .ZN(n6695) );
  OAI221_X1 U7621 ( .B1(DATAI_16_), .B2(keyinput_g15), .C1(
        REIP_REG_31__SCAN_IN), .C2(keyinput_g51), .A(n6695), .ZN(n6698) );
  AOI22_X1 U7622 ( .A1(BS16_N), .A2(keyinput_g34), .B1(FLUSH_REG_SCAN_IN), 
        .B2(keyinput_g45), .ZN(n6696) );
  OAI221_X1 U7623 ( .B1(BS16_N), .B2(keyinput_g34), .C1(FLUSH_REG_SCAN_IN), 
        .C2(keyinput_g45), .A(n6696), .ZN(n6697) );
  NOR4_X1 U7624 ( .A1(n6700), .A2(n6699), .A3(n6698), .A4(n6697), .ZN(n6710)
         );
  AOI22_X1 U7625 ( .A1(D_C_N_REG_SCAN_IN), .A2(keyinput_g41), .B1(
        REIP_REG_21__SCAN_IN), .B2(keyinput_g61), .ZN(n6701) );
  OAI221_X1 U7626 ( .B1(D_C_N_REG_SCAN_IN), .B2(keyinput_g41), .C1(
        REIP_REG_21__SCAN_IN), .C2(keyinput_g61), .A(n6701), .ZN(n6708) );
  AOI22_X1 U7627 ( .A1(BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_g48), .B1(
        BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_g47), .ZN(n6702) );
  OAI221_X1 U7628 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_g48), .C1(
        BYTEENABLE_REG_0__SCAN_IN), .C2(keyinput_g47), .A(n6702), .ZN(n6707)
         );
  AOI22_X1 U7629 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_g50), .B1(
        REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_g42), .ZN(n6703) );
  OAI221_X1 U7630 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_g50), .C1(
        REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_g42), .A(n6703), .ZN(n6706)
         );
  AOI22_X1 U7631 ( .A1(DATAI_27_), .A2(keyinput_g4), .B1(REIP_REG_29__SCAN_IN), 
        .B2(keyinput_g53), .ZN(n6704) );
  OAI221_X1 U7632 ( .B1(DATAI_27_), .B2(keyinput_g4), .C1(REIP_REG_29__SCAN_IN), .C2(keyinput_g53), .A(n6704), .ZN(n6705) );
  NOR4_X1 U7633 ( .A1(n6708), .A2(n6707), .A3(n6706), .A4(n6705), .ZN(n6709)
         );
  NAND4_X1 U7634 ( .A1(n6712), .A2(n6711), .A3(n6710), .A4(n6709), .ZN(n6774)
         );
  INV_X1 U7635 ( .A(DATAI_15_), .ZN(n6715) );
  AOI22_X1 U7636 ( .A1(n6715), .A2(keyinput_g16), .B1(n6714), .B2(keyinput_g30), .ZN(n6713) );
  OAI221_X1 U7637 ( .B1(n6715), .B2(keyinput_g16), .C1(n6714), .C2(
        keyinput_g30), .A(n6713), .ZN(n6727) );
  AOI22_X1 U7638 ( .A1(n6717), .A2(keyinput_g40), .B1(n4502), .B2(keyinput_g12), .ZN(n6716) );
  OAI221_X1 U7639 ( .B1(n6717), .B2(keyinput_g40), .C1(n4502), .C2(
        keyinput_g12), .A(n6716), .ZN(n6726) );
  AOI22_X1 U7640 ( .A1(n6720), .A2(keyinput_g58), .B1(keyinput_g24), .B2(n6719), .ZN(n6718) );
  OAI221_X1 U7641 ( .B1(n6720), .B2(keyinput_g58), .C1(n6719), .C2(
        keyinput_g24), .A(n6718), .ZN(n6725) );
  AOI22_X1 U7642 ( .A1(n6723), .A2(keyinput_g43), .B1(keyinput_g56), .B2(n6722), .ZN(n6721) );
  OAI221_X1 U7643 ( .B1(n6723), .B2(keyinput_g43), .C1(n6722), .C2(
        keyinput_g56), .A(n6721), .ZN(n6724) );
  NOR4_X1 U7644 ( .A1(n6727), .A2(n6726), .A3(n6725), .A4(n6724), .ZN(n6772)
         );
  AOI22_X1 U7645 ( .A1(DATAI_0_), .A2(keyinput_g31), .B1(DATAI_23_), .B2(
        keyinput_g8), .ZN(n6728) );
  OAI221_X1 U7646 ( .B1(DATAI_0_), .B2(keyinput_g31), .C1(DATAI_23_), .C2(
        keyinput_g8), .A(n6728), .ZN(n6738) );
  AOI22_X1 U7647 ( .A1(BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput_g49), .B1(
        READREQUEST_REG_SCAN_IN), .B2(keyinput_g37), .ZN(n6729) );
  OAI221_X1 U7648 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_g49), .C1(
        READREQUEST_REG_SCAN_IN), .C2(keyinput_g37), .A(n6729), .ZN(n6737) );
  AOI22_X1 U7649 ( .A1(n6732), .A2(keyinput_g32), .B1(n6731), .B2(keyinput_g0), 
        .ZN(n6730) );
  OAI221_X1 U7650 ( .B1(n6732), .B2(keyinput_g32), .C1(n6731), .C2(keyinput_g0), .A(n6730), .ZN(n6736) );
  AOI22_X1 U7651 ( .A1(REIP_REG_23__SCAN_IN), .A2(keyinput_g59), .B1(n6734), 
        .B2(keyinput_g63), .ZN(n6733) );
  OAI221_X1 U7652 ( .B1(REIP_REG_23__SCAN_IN), .B2(keyinput_g59), .C1(n6734), 
        .C2(keyinput_g63), .A(n6733), .ZN(n6735) );
  NOR4_X1 U7653 ( .A1(n6738), .A2(n6737), .A3(n6736), .A4(n6735), .ZN(n6771)
         );
  AOI22_X1 U7654 ( .A1(n6740), .A2(keyinput_g27), .B1(keyinput_g14), .B2(n4476), .ZN(n6739) );
  OAI221_X1 U7655 ( .B1(n6740), .B2(keyinput_g27), .C1(n4476), .C2(
        keyinput_g14), .A(n6739), .ZN(n6752) );
  AOI22_X1 U7656 ( .A1(n6071), .A2(keyinput_g17), .B1(keyinput_g5), .B2(n6742), 
        .ZN(n6741) );
  OAI221_X1 U7657 ( .B1(n6071), .B2(keyinput_g17), .C1(n6742), .C2(keyinput_g5), .A(n6741), .ZN(n6751) );
  AOI22_X1 U7658 ( .A1(n6745), .A2(keyinput_g46), .B1(n6744), .B2(keyinput_g39), .ZN(n6743) );
  OAI221_X1 U7659 ( .B1(n6745), .B2(keyinput_g46), .C1(n6744), .C2(
        keyinput_g39), .A(n6743), .ZN(n6750) );
  AOI22_X1 U7660 ( .A1(n6748), .A2(keyinput_g6), .B1(keyinput_g11), .B2(n6747), 
        .ZN(n6746) );
  OAI221_X1 U7661 ( .B1(n6748), .B2(keyinput_g6), .C1(n6747), .C2(keyinput_g11), .A(n6746), .ZN(n6749) );
  NOR4_X1 U7662 ( .A1(n6752), .A2(n6751), .A3(n6750), .A4(n6749), .ZN(n6770)
         );
  AOI22_X1 U7663 ( .A1(n6755), .A2(keyinput_g1), .B1(keyinput_g28), .B2(n6754), 
        .ZN(n6753) );
  OAI221_X1 U7664 ( .B1(n6755), .B2(keyinput_g1), .C1(n6754), .C2(keyinput_g28), .A(n6753), .ZN(n6768) );
  INV_X1 U7665 ( .A(DATAI_13_), .ZN(n6758) );
  AOI22_X1 U7666 ( .A1(n6758), .A2(keyinput_g18), .B1(keyinput_g23), .B2(n6757), .ZN(n6756) );
  OAI221_X1 U7667 ( .B1(n6758), .B2(keyinput_g18), .C1(n6757), .C2(
        keyinput_g23), .A(n6756), .ZN(n6767) );
  AOI22_X1 U7668 ( .A1(n6761), .A2(keyinput_g35), .B1(keyinput_g3), .B2(n6760), 
        .ZN(n6759) );
  OAI221_X1 U7669 ( .B1(n6761), .B2(keyinput_g35), .C1(n6760), .C2(keyinput_g3), .A(n6759), .ZN(n6766) );
  AOI22_X1 U7670 ( .A1(n6764), .A2(keyinput_g52), .B1(keyinput_g44), .B2(n6763), .ZN(n6762) );
  OAI221_X1 U7671 ( .B1(n6764), .B2(keyinput_g52), .C1(n6763), .C2(
        keyinput_g44), .A(n6762), .ZN(n6765) );
  NOR4_X1 U7672 ( .A1(n6768), .A2(n6767), .A3(n6766), .A4(n6765), .ZN(n6769)
         );
  NAND4_X1 U7673 ( .A1(n6772), .A2(n6771), .A3(n6770), .A4(n6769), .ZN(n6773)
         );
  OAI22_X1 U7674 ( .A1(DATAI_10_), .A2(keyinput_g21), .B1(n6774), .B2(n6773), 
        .ZN(n6775) );
  AOI211_X1 U7675 ( .C1(DATAI_10_), .C2(keyinput_g21), .A(n6776), .B(n6775), 
        .ZN(n6780) );
  AOI22_X1 U7676 ( .A1(n6778), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6777), .ZN(n6779) );
  XNOR2_X1 U7677 ( .A(n6780), .B(n6779), .ZN(U3445) );
  AND2_X2 U3523 ( .A1(n3011), .A2(n4327), .ZN(n3196) );
  CLKBUF_X2 U3443 ( .A(n3204), .Z(n3259) );
  CLKBUF_X2 U3442 ( .A(n3221), .Z(n4413) );
  XNOR2_X1 U6466 ( .A(n5303), .B(n5302), .ZN(n5313) );
  CLKBUF_X1 U3520 ( .A(n4179), .Z(n4103) );
  AND4_X1 U3527 ( .A1(n3015), .A2(n3014), .A3(n3013), .A4(n3012), .ZN(n3006)
         );
  OR2_X1 U3533 ( .A1(n3699), .A2(n3537), .ZN(n4372) );
  CLKBUF_X1 U3623 ( .A(n3127), .Z(n5287) );
  CLKBUF_X1 U3629 ( .A(n5252), .Z(n5419) );
  CLKBUF_X1 U3661 ( .A(n5022), .Z(n5060) );
  CLKBUF_X1 U3667 ( .A(n3526), .Z(n4271) );
  CLKBUF_X1 U3695 ( .A(n3708), .Z(n6314) );
  CLKBUF_X1 U3753 ( .A(n4214), .Z(n4247) );
  CLKBUF_X1 U4030 ( .A(n5521), .Z(n5523) );
endmodule

