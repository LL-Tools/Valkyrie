

module b15_C_gen_AntiSAT_k_128_7 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, 
        U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, 
        U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, 
        U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, 
        U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, 
        U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, 
        U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, 
        U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, 
        U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, 
        U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, 
        U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, 
        U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, 
        U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, 
        U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, 
        U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, 
        U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, 
        U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, 
        U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, 
        U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, 
        U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, 
        U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, 
        U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, 
        U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, 
        U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, 
        U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, 
        U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, 
        U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, 
        U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, 
        U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, 
        U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, 
        U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, 
        U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, 
        U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, 
        U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, 
        U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, 
        U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, 
        U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, 
        U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, 
        U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, 
        U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, 
        U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, 
        U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, 
        U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, 
        U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, 
        U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, 
        U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741;

  AOI21_X1 U3430 ( .B1(n5609), .B2(n2983), .A(n5608), .ZN(n5610) );
  AOI21_X1 U3431 ( .B1(n5422), .B2(n5421), .A(n5420), .ZN(n5602) );
  OR2_X1 U3432 ( .A1(n5307), .A2(n5308), .ZN(n5421) );
  OR2_X1 U3433 ( .A1(n5307), .A2(n5407), .ZN(n5419) );
  OR2_X1 U3434 ( .A1(n5538), .A2(n5539), .ZN(n5485) );
  CLKBUF_X1 U3435 ( .A(n3764), .Z(n4398) );
  BUF_X1 U3436 ( .A(n3641), .Z(n3026) );
  CLKBUF_X2 U3437 ( .A(n3154), .Z(n5266) );
  CLKBUF_X2 U3438 ( .A(n3226), .Z(n4189) );
  CLKBUF_X2 U3439 ( .A(n3135), .Z(n4194) );
  CLKBUF_X2 U3440 ( .A(n3127), .Z(n5276) );
  CLKBUF_X2 U3441 ( .A(n3134), .Z(n5274) );
  CLKBUF_X2 U3442 ( .A(n3095), .Z(n4188) );
  CLKBUF_X2 U3443 ( .A(n3136), .Z(n4187) );
  CLKBUF_X2 U3444 ( .A(n3263), .Z(n2986) );
  CLKBUF_X1 U34450 ( .A(n3593), .Z(n4492) );
  NAND2_X1 U34460 ( .A1(n3029), .A2(n3122), .ZN(n3189) );
  AND2_X2 U34470 ( .A1(n3047), .A2(n3049), .ZN(n3138) );
  AND2_X2 U34480 ( .A1(n3042), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3047) );
  INV_X1 U3449 ( .A(n5258), .ZN(n3193) );
  INV_X1 U3450 ( .A(n3189), .ZN(n3580) );
  INV_X1 U34510 ( .A(n3604), .ZN(n3251) );
  INV_X1 U34520 ( .A(n3032), .ZN(n4204) );
  BUF_X1 U34530 ( .A(n4709), .Z(n3022) );
  NAND2_X1 U3454 ( .A1(n3251), .A2(n3187), .ZN(n3510) );
  NOR2_X1 U34550 ( .A1(n5316), .A2(n5315), .ZN(n5319) );
  AOI21_X1 U34560 ( .B1(n3803), .B2(n3930), .A(n3802), .ZN(n4837) );
  AOI21_X1 U3457 ( .B1(n2982), .B2(n3022), .A(n3643), .ZN(n4458) );
  INV_X2 U3458 ( .A(n3593), .ZN(n3187) );
  AND2_X1 U34590 ( .A1(n3562), .A2(n3561), .ZN(n5404) );
  AND2_X1 U34600 ( .A1(n5526), .A2(n5525), .ZN(n5528) );
  NOR2_X1 U34610 ( .A1(n6425), .A2(n6017), .ZN(n6047) );
  AOI21_X1 U34620 ( .B1(n5408), .B2(n5419), .A(n4207), .ZN(n5594) );
  INV_X1 U34630 ( .A(n5968), .ZN(n5996) );
  XOR2_X1 U34640 ( .A(n3642), .B(n4346), .Z(n2982) );
  AND2_X2 U34650 ( .A1(n3177), .A2(n4300), .ZN(n3214) );
  AOI22_X2 U3466 ( .A1(n3411), .A2(n3410), .B1(n3409), .B2(n4960), .ZN(n4932)
         );
  NAND2_X2 U3467 ( .A1(n4207), .A2(n4208), .ZN(n5316) );
  NAND2_X2 U34680 ( .A1(n3066), .A2(n3065), .ZN(n3176) );
  AND2_X2 U34700 ( .A1(n3182), .A2(n3218), .ZN(n3592) );
  AND2_X4 U34710 ( .A1(n3048), .A2(n3047), .ZN(n3129) );
  AND2_X2 U34720 ( .A1(n3040), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3048) );
  NOR2_X4 U34730 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4423) );
  CLKBUF_X1 U34740 ( .A(n5650), .Z(n3000) );
  AND2_X1 U3475 ( .A1(n5653), .A2(n5651), .ZN(n5650) );
  NAND2_X1 U3476 ( .A1(n3501), .A2(n3027), .ZN(n5653) );
  AND2_X1 U3477 ( .A1(n2996), .A2(n2997), .ZN(n2989) );
  AND2_X1 U3478 ( .A1(n5068), .A2(n2997), .ZN(n2988) );
  INV_X1 U3479 ( .A(n5427), .ZN(n3001) );
  NAND2_X1 U3480 ( .A1(n4934), .A2(n3434), .ZN(n6063) );
  NAND2_X1 U3481 ( .A1(n5672), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5034)
         );
  INV_X2 U3482 ( .A(n3477), .ZN(n5672) );
  NAND2_X1 U3483 ( .A1(n6069), .A2(n6070), .ZN(n4960) );
  NAND2_X1 U3484 ( .A1(n4452), .A2(n4460), .ZN(n4580) );
  OR2_X1 U3485 ( .A1(n3764), .A2(n3763), .ZN(n4454) );
  CLKBUF_X1 U3486 ( .A(n4470), .Z(n5805) );
  CLKBUF_X2 U3487 ( .A(n3751), .Z(n5046) );
  CLKBUF_X1 U3488 ( .A(n3290), .Z(n3320) );
  NAND2_X1 U3489 ( .A1(n3586), .A2(n3188), .ZN(n5903) );
  CLKBUF_X1 U3490 ( .A(n3592), .Z(n2995) );
  AND2_X1 U3491 ( .A1(n3210), .A2(n4499), .ZN(n3125) );
  BUF_X2 U3492 ( .A(n3606), .Z(n5535) );
  INV_X1 U3493 ( .A(n3641), .ZN(n4709) );
  AND2_X1 U3494 ( .A1(n3190), .A2(n3593), .ZN(n3606) );
  NAND2_X1 U3495 ( .A1(n3593), .A2(n3604), .ZN(n3641) );
  CLKBUF_X2 U3496 ( .A(n3218), .Z(n5259) );
  CLKBUF_X2 U3497 ( .A(n3604), .Z(n3602) );
  INV_X2 U3498 ( .A(n3298), .ZN(n5275) );
  BUF_X2 U3499 ( .A(n3129), .Z(n2985) );
  CLKBUF_X2 U3500 ( .A(n5273), .Z(n4121) );
  BUF_X2 U3501 ( .A(n3128), .Z(n5268) );
  OAI21_X1 U3502 ( .B1(n4207), .B2(n4208), .A(n5316), .ZN(n5386) );
  OAI22_X1 U3503 ( .A1(n5621), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5631), .B2(n5620), .ZN(n5622) );
  NAND2_X1 U3504 ( .A1(n3019), .A2(n5619), .ZN(n5631) );
  AND2_X2 U3505 ( .A1(n5441), .A2(n2992), .ZN(n4207) );
  CLKBUF_X1 U3506 ( .A(n5300), .Z(n5517) );
  CLKBUF_X1 U3507 ( .A(n5476), .Z(n5524) );
  CLKBUF_X1 U3508 ( .A(n5531), .Z(n5543) );
  AND2_X1 U3509 ( .A1(n4283), .A2(n4282), .ZN(n4284) );
  XNOR2_X1 U3510 ( .A(n4277), .B(n4276), .ZN(n5331) );
  AOI21_X1 U3511 ( .B1(n4274), .B2(n5369), .A(n4273), .ZN(n4277) );
  NAND2_X1 U3512 ( .A1(n4986), .A2(n4985), .ZN(n4984) );
  NAND2_X1 U3513 ( .A1(n3030), .A2(n4272), .ZN(n5369) );
  CLKBUF_X1 U3514 ( .A(n4971), .Z(n5008) );
  NAND2_X1 U3515 ( .A1(n3477), .A2(n3018), .ZN(n3019) );
  NAND2_X1 U3516 ( .A1(n3004), .A2(n3005), .ZN(n5312) );
  NOR2_X1 U3517 ( .A1(n5407), .A2(n5408), .ZN(n4184) );
  INV_X1 U3518 ( .A(n5444), .ZN(n3004) );
  NAND2_X1 U3519 ( .A1(n4224), .A2(n5458), .ZN(n5444) );
  NOR2_X1 U3520 ( .A1(n4578), .A2(n4588), .ZN(n4586) );
  AND2_X1 U3521 ( .A1(n3414), .A2(n3413), .ZN(n2987) );
  AND2_X1 U3522 ( .A1(n5213), .A2(n5214), .ZN(n5240) );
  OR2_X1 U3523 ( .A1(n4351), .A2(n3757), .ZN(n4352) );
  NAND2_X1 U3524 ( .A1(n3342), .A2(n3341), .ZN(n4480) );
  NAND2_X1 U3525 ( .A1(n4691), .A2(n4690), .ZN(n6538) );
  OR2_X2 U3526 ( .A1(n4691), .A2(n4492), .ZN(n4355) );
  OR2_X1 U3527 ( .A1(n3009), .A2(n3010), .ZN(n5025) );
  INV_X1 U3528 ( .A(n4462), .ZN(n3012) );
  OR2_X1 U3529 ( .A1(n3320), .A2(n3319), .ZN(n3326) );
  OR2_X1 U3530 ( .A1(n3320), .A2(n3291), .ZN(n3296) );
  NAND2_X1 U3531 ( .A1(n3201), .A2(n3202), .ZN(n3288) );
  NAND2_X1 U3532 ( .A1(n4458), .A2(n4457), .ZN(n4462) );
  AND2_X1 U3533 ( .A1(n3203), .A2(n3200), .ZN(n3201) );
  OAI211_X1 U3534 ( .C1(n5396), .C2(n3195), .A(n5903), .B(n3594), .ZN(n3196)
         );
  NAND2_X1 U3535 ( .A1(n3637), .A2(n3034), .ZN(n3642) );
  INV_X1 U3536 ( .A(n3684), .ZN(n4232) );
  AND3_X1 U3537 ( .A1(n3636), .A2(n3675), .A3(n3635), .ZN(n3034) );
  AND2_X2 U3538 ( .A1(n5535), .A2(n4709), .ZN(n4234) );
  AND2_X1 U3539 ( .A1(n3328), .A2(n3327), .ZN(n3552) );
  NOR2_X1 U3540 ( .A1(n3276), .A2(n6536), .ZN(n3279) );
  INV_X1 U3541 ( .A(n3376), .ZN(n3184) );
  AND2_X1 U3542 ( .A1(n3208), .A2(n3191), .ZN(n3192) );
  INV_X1 U3543 ( .A(n3638), .ZN(n4236) );
  AND2_X1 U3544 ( .A1(n3603), .A2(n3602), .ZN(n3024) );
  INV_X2 U3545 ( .A(n3606), .ZN(n5371) );
  AND2_X1 U3546 ( .A1(n3173), .A2(n4499), .ZN(n3183) );
  CLKBUF_X1 U3547 ( .A(n3173), .Z(n3583) );
  OR2_X1 U3548 ( .A1(n3250), .A2(n3249), .ZN(n3479) );
  BUF_X1 U3549 ( .A(n3123), .Z(n4503) );
  INV_X1 U3550 ( .A(n2990), .ZN(n3113) );
  CLKBUF_X1 U3551 ( .A(n3176), .Z(n3218) );
  NAND4_X2 U3552 ( .A1(n3166), .A2(n3165), .A3(n3164), .A4(n3163), .ZN(n3604)
         );
  AND4_X1 U3553 ( .A1(n3158), .A2(n3157), .A3(n3156), .A4(n3155), .ZN(n3164)
         );
  AND4_X1 U3554 ( .A1(n3148), .A2(n3147), .A3(n3146), .A4(n3145), .ZN(n3166)
         );
  NAND2_X1 U3555 ( .A1(n3143), .A2(n3031), .ZN(n3593) );
  AND4_X1 U3556 ( .A1(n3121), .A2(n3120), .A3(n3119), .A4(n3118), .ZN(n3122)
         );
  AND4_X1 U3557 ( .A1(n3152), .A2(n3151), .A3(n3150), .A4(n3149), .ZN(n3165)
         );
  AND4_X1 U3558 ( .A1(n3046), .A2(n3045), .A3(n3044), .A4(n3043), .ZN(n3056)
         );
  AND4_X1 U3559 ( .A1(n3054), .A2(n3053), .A3(n3052), .A4(n3051), .ZN(n3055)
         );
  AND4_X1 U3560 ( .A1(n3094), .A2(n3093), .A3(n3092), .A4(n3091), .ZN(n3111)
         );
  AND4_X1 U3561 ( .A1(n3064), .A2(n3063), .A3(n3062), .A4(n3061), .ZN(n3065)
         );
  AND4_X1 U3562 ( .A1(n3099), .A2(n3098), .A3(n3097), .A4(n3096), .ZN(n3110)
         );
  AND4_X1 U3563 ( .A1(n3162), .A2(n3161), .A3(n3160), .A4(n3159), .ZN(n3163)
         );
  AND4_X1 U3564 ( .A1(n3133), .A2(n3132), .A3(n3131), .A4(n3130), .ZN(n3143)
         );
  AOI21_X1 U3565 ( .B1(n3136), .B2(INSTQUEUE_REG_4__3__SCAN_IN), .A(n3070), 
        .ZN(n3071) );
  INV_X2 U3566 ( .A(n5687), .ZN(n2983) );
  BUF_X2 U3567 ( .A(n3297), .Z(n2984) );
  AND2_X2 U3568 ( .A1(n3050), .A2(n4303), .ZN(n3137) );
  AND2_X2 U3569 ( .A1(n3047), .A2(n4303), .ZN(n3226) );
  INV_X2 U3570 ( .A(n6739), .ZN(n6500) );
  AND2_X2 U3571 ( .A1(n4423), .A2(n4433), .ZN(n3095) );
  AND2_X2 U3572 ( .A1(n3318), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3050)
         );
  AND2_X2 U3573 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4303) );
  AND2_X2 U3574 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4422) );
  CLKBUF_X1 U3575 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n4416) );
  NOR2_X2 U3576 ( .A1(n5404), .A2(n6438), .ZN(n4740) );
  AOI211_X1 U3577 ( .C1(REIP_REG_31__SCAN_IN), .C2(n5335), .A(n5334), .B(n5333), .ZN(n5336) );
  OR2_X2 U3578 ( .A1(n2998), .A2(n5033), .ZN(n2997) );
  CLKBUF_X1 U3579 ( .A(n3178), .Z(n3191) );
  AND2_X2 U3580 ( .A1(n3050), .A2(n4433), .ZN(n3136) );
  NAND2_X1 U3581 ( .A1(n3055), .A2(n3056), .ZN(n2990) );
  OR2_X2 U3582 ( .A1(n3079), .A2(n3078), .ZN(n3190) );
  NAND2_X1 U3583 ( .A1(n3055), .A2(n3056), .ZN(n3123) );
  AND2_X2 U3584 ( .A1(n4423), .A2(n4303), .ZN(n3128) );
  AND2_X1 U3585 ( .A1(n3167), .A2(n3251), .ZN(n2991) );
  NAND2_X2 U3586 ( .A1(n3185), .A2(n3602), .ZN(n5396) );
  AND2_X1 U3587 ( .A1(n5442), .A2(n4184), .ZN(n2992) );
  NAND2_X1 U3588 ( .A1(n5441), .A2(n5442), .ZN(n5307) );
  AND2_X1 U3589 ( .A1(n2994), .A2(STATE2_REG_0__SCAN_IN), .ZN(n2993) );
  OAI211_X1 U3590 ( .C1(n5396), .C2(n3195), .A(n5903), .B(n3594), .ZN(n2994)
         );
  AND2_X2 U3591 ( .A1(n5477), .A2(n5479), .ZN(n5476) );
  XNOR2_X1 U3592 ( .A(n3374), .B(n3373), .ZN(n4471) );
  NAND2_X1 U3593 ( .A1(n4984), .A2(n2999), .ZN(n2996) );
  INV_X1 U3594 ( .A(n5034), .ZN(n2998) );
  AND2_X1 U3595 ( .A1(n3483), .A2(n5034), .ZN(n2999) );
  AND2_X2 U3596 ( .A1(n3050), .A2(n3049), .ZN(n3263) );
  AND2_X2 U3597 ( .A1(n3048), .A2(n4422), .ZN(n3297) );
  AND2_X2 U3598 ( .A1(n3049), .A2(n4422), .ZN(n3153) );
  AND2_X1 U3599 ( .A1(n5372), .A2(n3002), .ZN(n3003) );
  INV_X1 U3600 ( .A(n5409), .ZN(n3002) );
  AND2_X1 U3601 ( .A1(n3001), .A2(n3002), .ZN(n5410) );
  AND2_X1 U3602 ( .A1(n4231), .A2(n3005), .ZN(n3006) );
  INV_X1 U3603 ( .A(n5445), .ZN(n3005) );
  AND2_X1 U3604 ( .A1(n5528), .A2(n3007), .ZN(n4224) );
  AND2_X1 U3605 ( .A1(n5520), .A2(n3008), .ZN(n3007) );
  INV_X1 U3606 ( .A(n3704), .ZN(n3008) );
  NAND2_X1 U3607 ( .A1(n4589), .A2(n4651), .ZN(n3009) );
  OR2_X1 U3608 ( .A1(n3011), .A2(n4839), .ZN(n3010) );
  INV_X1 U3609 ( .A(n4974), .ZN(n3011) );
  AND2_X1 U3610 ( .A1(n4583), .A2(n3013), .ZN(n3014) );
  INV_X1 U3611 ( .A(n4463), .ZN(n3013) );
  AND2_X1 U3612 ( .A1(n3012), .A2(n3013), .ZN(n4461) );
  INV_X1 U3613 ( .A(n2982), .ZN(n3015) );
  CLKBUF_X1 U3614 ( .A(n6061), .Z(n3016) );
  CLKBUF_X1 U3615 ( .A(n6052), .Z(n3017) );
  INV_X1 U3616 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3018) );
  OR2_X1 U3617 ( .A1(n3647), .A2(n3646), .ZN(n4457) );
  AND2_X1 U3618 ( .A1(n3047), .A2(n3049), .ZN(n3020) );
  AND2_X1 U3619 ( .A1(n4433), .A2(n4422), .ZN(n3021) );
  AND2_X1 U3620 ( .A1(n3050), .A2(n4303), .ZN(n3023) );
  OR2_X1 U3621 ( .A1(n3290), .A2(n3181), .ZN(n3202) );
  AND2_X1 U3622 ( .A1(n3603), .A2(n3602), .ZN(n3025) );
  AND2_X1 U3623 ( .A1(n3603), .A2(n3602), .ZN(n3638) );
  XNOR2_X2 U3624 ( .A(n3225), .B(n3224), .ZN(n4465) );
  AOI21_X1 U3625 ( .B1(n3786), .B2(n3930), .A(n3790), .ZN(n4588) );
  NOR2_X4 U3626 ( .A1(n5611), .A2(n3726), .ZN(n5605) );
  AND4_X4 U3627 ( .A1(n3111), .A2(n3110), .A3(n3109), .A4(n3108), .ZN(n3175)
         );
  AOI21_X2 U3628 ( .B1(n3153), .B2(INSTQUEUE_REG_14__4__SCAN_IN), .A(n3103), 
        .ZN(n3109) );
  AND4_X1 U3629 ( .A1(n3107), .A2(n3106), .A3(n3105), .A4(n3104), .ZN(n3108)
         );
  XNOR2_X1 U3630 ( .A(n3363), .B(n6168), .ZN(n4962) );
  NAND2_X1 U3631 ( .A1(n3362), .A2(n3361), .ZN(n3363) );
  NOR2_X2 U3632 ( .A1(n5485), .A2(n3696), .ZN(n5526) );
  NOR2_X2 U3633 ( .A1(n5496), .A2(n5497), .ZN(n5213) );
  INV_X1 U3634 ( .A(n3398), .ZN(n3356) );
  INV_X1 U3635 ( .A(n3176), .ZN(n3178) );
  NAND2_X1 U3636 ( .A1(n3602), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3508) );
  NAND2_X1 U3637 ( .A1(n3182), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3328) );
  NAND2_X1 U3638 ( .A1(n3251), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3327) );
  AND2_X1 U3639 ( .A1(n3477), .A2(n5893), .ZN(n3495) );
  AND2_X2 U3640 ( .A1(n3041), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3049)
         );
  NAND2_X1 U3641 ( .A1(n3258), .A2(n3256), .ZN(n3287) );
  OR2_X1 U3642 ( .A1(n3338), .A2(n3337), .ZN(n3357) );
  INV_X1 U3643 ( .A(n5519), .ZN(n4047) );
  XNOR2_X1 U3644 ( .A(n3476), .B(n3464), .ZN(n3803) );
  OR2_X1 U3645 ( .A1(n3309), .A2(n3308), .ZN(n3398) );
  INV_X1 U3646 ( .A(n5689), .ZN(n3496) );
  INV_X1 U3647 ( .A(n3510), .ZN(n3596) );
  NAND2_X1 U3648 ( .A1(n3238), .A2(n3237), .ZN(n3372) );
  OR2_X1 U3649 ( .A1(n3252), .A2(n3328), .ZN(n3237) );
  OAI211_X1 U3650 ( .C1(n3529), .C2(n3255), .A(n3254), .B(n3253), .ZN(n3370)
         );
  XNOR2_X1 U3651 ( .A(n4435), .B(n4853), .ZN(n4414) );
  OR2_X1 U3652 ( .A1(n3508), .A2(n3175), .ZN(n3529) );
  INV_X1 U3653 ( .A(n6538), .ZN(n4724) );
  NAND2_X1 U3654 ( .A1(n4179), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4696)
         );
  OR2_X1 U3655 ( .A1(n5004), .A2(n3866), .ZN(n3867) );
  NOR2_X2 U3656 ( .A1(n5597), .A2(n4259), .ZN(n4263) );
  AND2_X1 U3657 ( .A1(n5200), .A2(n5196), .ZN(n6134) );
  CLKBUF_X1 U3658 ( .A(n3600), .Z(n3601) );
  AOI21_X1 U3659 ( .B1(n3591), .B2(n3590), .A(n6438), .ZN(n3634) );
  AND2_X1 U3660 ( .A1(n3175), .A2(n3123), .ZN(n3126) );
  NAND2_X1 U3661 ( .A1(n3317), .A2(n3316), .ZN(n4435) );
  INV_X1 U3662 ( .A(n3315), .ZN(n3317) );
  AOI22_X1 U3663 ( .A1(n3135), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3073) );
  AND2_X1 U3664 ( .A1(n4950), .A2(n4707), .ZN(n5968) );
  INV_X1 U3665 ( .A(n5581), .ZN(n6013) );
  OAI211_X1 U3666 ( .C1(n4248), .C2(n4247), .A(n4246), .B(n4245), .ZN(n4249)
         );
  OR2_X1 U3667 ( .A1(n5777), .A2(n3713), .ZN(n5756) );
  XNOR2_X1 U3668 ( .A(n3504), .B(n3503), .ZN(n5302) );
  INV_X1 U3669 ( .A(n6157), .ZN(n6183) );
  INV_X1 U3670 ( .A(n6160), .ZN(n6180) );
  OR2_X1 U3671 ( .A1(n3552), .A2(n3187), .ZN(n3505) );
  AOI22_X1 U3672 ( .A1(n3263), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3051) );
  AOI22_X1 U3673 ( .A1(n3129), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3128), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3052) );
  OR2_X1 U3674 ( .A1(n3236), .A2(n3235), .ZN(n3375) );
  NOR2_X1 U3675 ( .A1(n3216), .A2(n3215), .ZN(n3223) );
  NAND2_X1 U3676 ( .A1(n2993), .A2(n3038), .ZN(n3286) );
  NAND2_X1 U3677 ( .A1(n3180), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3290) );
  NOR2_X1 U3678 ( .A1(n3921), .A2(n3920), .ZN(n3938) );
  OR2_X1 U3679 ( .A1(n3850), .A2(n5007), .ZN(n5004) );
  INV_X1 U3680 ( .A(n4581), .ZN(n3784) );
  AND2_X1 U3681 ( .A1(n5371), .A2(n3022), .ZN(n3684) );
  INV_X1 U3682 ( .A(n3287), .ZN(n3224) );
  NAND2_X1 U3683 ( .A1(n3288), .A2(n3286), .ZN(n3225) );
  INV_X1 U3684 ( .A(n3370), .ZN(n3282) );
  XNOR2_X1 U3685 ( .A(n3313), .B(n3312), .ZN(n3397) );
  AOI21_X1 U3686 ( .B1(n4299), .B2(n6536), .A(n3310), .ZN(n3313) );
  NAND2_X1 U3687 ( .A1(n3592), .A2(n3606), .ZN(n4300) );
  OR2_X1 U3688 ( .A1(n3547), .A2(n3546), .ZN(n3557) );
  NAND2_X1 U3689 ( .A1(n3289), .A2(n3288), .ZN(n3315) );
  NAND2_X1 U3690 ( .A1(n3287), .A2(n3286), .ZN(n3289) );
  CLKBUF_X1 U3691 ( .A(n3318), .Z(n3319) );
  NOR2_X1 U3692 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4478), .ZN(n4658) );
  AOI22_X1 U3693 ( .A1(n3129), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3021), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3116) );
  AOI21_X1 U3694 ( .B1(n3138), .B2(INSTQUEUE_REG_10__7__SCAN_IN), .A(n3080), 
        .ZN(n3081) );
  AND2_X1 U3695 ( .A1(n3154), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3080) );
  AOI21_X1 U3696 ( .B1(n6535), .B2(n4743), .A(n6521), .ZN(n4478) );
  INV_X1 U3697 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5135) );
  INV_X1 U3698 ( .A(n5327), .ZN(n5991) );
  AND2_X1 U3699 ( .A1(n4270), .A2(n5371), .ZN(n4273) );
  NAND2_X1 U3700 ( .A1(n3891), .A2(n3874), .ZN(n3878) );
  AND2_X1 U3701 ( .A1(n5076), .A2(n3891), .ZN(n3876) );
  NAND2_X1 U3702 ( .A1(n5128), .A2(n5127), .ZN(n5126) );
  NAND2_X1 U3703 ( .A1(n3797), .A2(n3796), .ZN(n4648) );
  AND2_X1 U3704 ( .A1(n4742), .A2(n6455), .ZN(n6017) );
  INV_X1 U3705 ( .A(n4395), .ZN(n4373) );
  AND2_X1 U3706 ( .A1(n4178), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4179)
         );
  NOR2_X1 U3707 ( .A1(n4089), .A2(n5466), .ZN(n4090) );
  AND2_X1 U3708 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n4041), .ZN(n4042)
         );
  CLKBUF_X1 U3709 ( .A(n5515), .Z(n5516) );
  NAND2_X1 U3710 ( .A1(n3991), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4040)
         );
  CLKBUF_X1 U3711 ( .A(n5477), .Z(n5478) );
  NOR2_X1 U3712 ( .A1(n3955), .A2(n5680), .ZN(n3956) );
  AND2_X1 U3713 ( .A1(n3956), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3990)
         );
  CLKBUF_X1 U3714 ( .A(n5235), .Z(n5236) );
  CLKBUF_X1 U3715 ( .A(n5207), .Z(n5208) );
  AND2_X1 U3716 ( .A1(n5664), .A2(n3493), .ZN(n3494) );
  OR2_X1 U3717 ( .A1(n5663), .A2(n3495), .ZN(n5688) );
  NAND2_X1 U3718 ( .A1(n3906), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3921)
         );
  CLKBUF_X1 U3719 ( .A(n5186), .Z(n5494) );
  AND2_X1 U3720 ( .A1(n3868), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3869)
         );
  NOR2_X1 U3721 ( .A1(n3851), .A2(n3852), .ZN(n3868) );
  NAND2_X1 U3722 ( .A1(n3845), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3819)
         );
  AND2_X1 U3723 ( .A1(n3798), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3845)
         );
  BUF_X1 U3724 ( .A(n4647), .Z(n4836) );
  NAND2_X1 U3725 ( .A1(n3787), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3792)
         );
  INV_X1 U3726 ( .A(n3768), .ZN(n3779) );
  AND2_X1 U3727 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3779), .ZN(n3787)
         );
  INV_X1 U3728 ( .A(n3760), .ZN(n3769) );
  NAND2_X1 U3729 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3760) );
  NAND2_X1 U3730 ( .A1(n3731), .A2(n5714), .ZN(n4220) );
  NAND2_X1 U3731 ( .A1(n5605), .A2(n3727), .ZN(n5597) );
  NAND2_X1 U3732 ( .A1(n5240), .A2(n5241), .ZN(n5538) );
  NAND2_X1 U3733 ( .A1(n5129), .A2(n5189), .ZN(n5496) );
  CLKBUF_X1 U3734 ( .A(n5191), .Z(n5192) );
  AND2_X1 U3735 ( .A1(n3477), .A2(n3485), .ZN(n3488) );
  NOR2_X1 U3736 ( .A1(n3477), .A2(n5118), .ZN(n5109) );
  NOR2_X2 U3737 ( .A1(n5025), .A2(n5026), .ZN(n5024) );
  OR2_X1 U3738 ( .A1(n3656), .A2(n3655), .ZN(n4651) );
  NAND2_X1 U3739 ( .A1(n3194), .A2(n3193), .ZN(n3594) );
  CLKBUF_X1 U3740 ( .A(n3563), .Z(n4313) );
  XNOR2_X1 U3741 ( .A(n3371), .B(n3370), .ZN(n3374) );
  CLKBUF_X1 U3742 ( .A(n4465), .Z(n4466) );
  XNOR2_X1 U3743 ( .A(n3315), .B(n3316), .ZN(n4299) );
  NOR2_X1 U3744 ( .A1(n6517), .A2(n4478), .ZN(n4508) );
  INV_X1 U3745 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6409) );
  CLKBUF_X1 U3746 ( .A(n4414), .Z(n4415) );
  NAND2_X1 U3747 ( .A1(n4414), .A2(n6536), .ZN(n3342) );
  INV_X1 U3748 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5978) );
  NOR2_X1 U3749 ( .A1(n6470), .A2(n4841), .ZN(n5981) );
  INV_X1 U3750 ( .A(n5938), .ZN(n5987) );
  AND2_X1 U3751 ( .A1(n4950), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5956) );
  AND2_X1 U3752 ( .A1(n5861), .A2(n4700), .ZN(n5989) );
  AND2_X1 U3753 ( .A1(n6009), .A2(n5387), .ZN(n6005) );
  AND2_X1 U3754 ( .A1(n4350), .A2(n6426), .ZN(n6009) );
  INV_X1 U3755 ( .A(n6005), .ZN(n5549) );
  NAND2_X1 U3756 ( .A1(n4390), .A2(n4395), .ZN(n5581) );
  BUF_X1 U3757 ( .A(n6047), .Z(n6038) );
  CLKBUF_X2 U3758 ( .A(n6540), .Z(n6425) );
  OR2_X1 U3759 ( .A1(n5264), .A2(n5263), .ZN(n4698) );
  INV_X1 U3760 ( .A(n5386), .ZN(n4210) );
  CLKBUF_X1 U3761 ( .A(n5453), .Z(n5455) );
  OAI211_X1 U3762 ( .C1(n4280), .C2(n4279), .A(n4278), .B(n3028), .ZN(n4281)
         );
  OR2_X1 U3763 ( .A1(n5873), .A2(n3629), .ZN(n5774) );
  CLKBUF_X1 U3764 ( .A(n4471), .Z(n4472) );
  CLKBUF_X1 U3765 ( .A(n4299), .Z(n5806) );
  CLKBUF_X1 U3766 ( .A(n3767), .Z(n5810) );
  NOR2_X1 U3768 ( .A1(n6519), .A2(n5404), .ZN(n6521) );
  INV_X1 U3769 ( .A(n6232), .ZN(n6218) );
  INV_X1 U3770 ( .A(n6228), .ZN(n4927) );
  INV_X1 U3771 ( .A(n4521), .ZN(n6317) );
  OR2_X1 U3772 ( .A1(n4598), .A2(n4597), .ZN(n6393) );
  INV_X1 U3773 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6536) );
  AND2_X1 U3774 ( .A1(n4261), .A2(n4260), .ZN(n4262) );
  OR2_X1 U3775 ( .A1(n3715), .A2(n3714), .ZN(n3716) );
  BUF_X1 U3776 ( .A(n3175), .Z(n3182) );
  NOR2_X1 U3777 ( .A1(n3190), .A2(n3189), .ZN(n3208) );
  OR2_X1 U3778 ( .A1(n5662), .A2(n3711), .ZN(n3027) );
  INV_X1 U3779 ( .A(n3190), .ZN(n3603) );
  NAND2_X4 U3780 ( .A1(n3476), .A2(n3475), .ZN(n3477) );
  OR2_X1 U3781 ( .A1(n5331), .A2(n6160), .ZN(n3028) );
  AND4_X1 U3782 ( .A1(n3117), .A2(n3116), .A3(n3115), .A4(n3114), .ZN(n3029)
         );
  OR2_X1 U3783 ( .A1(n4270), .A2(n5535), .ZN(n3030) );
  AND4_X1 U3784 ( .A1(n3142), .A2(n3141), .A3(n3140), .A4(n3139), .ZN(n3031)
         );
  OR2_X1 U3785 ( .A1(n4499), .A2(n6534), .ZN(n3032) );
  NAND2_X1 U3786 ( .A1(n5528), .A2(n5520), .ZN(n3703) );
  INV_X1 U3787 ( .A(n4416), .ZN(n3291) );
  NOR2_X2 U3788 ( .A1(n5080), .A2(n5130), .ZN(n5129) );
  INV_X2 U3789 ( .A(n6159), .ZN(n6185) );
  OR2_X2 U3790 ( .A1(n4211), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6159) );
  CLKBUF_X1 U3791 ( .A(n4578), .Z(n4587) );
  INV_X1 U3792 ( .A(n5346), .ZN(n5362) );
  XNOR2_X1 U3793 ( .A(n3396), .B(n3397), .ZN(n4470) );
  NAND2_X1 U3794 ( .A1(n3385), .A2(n3384), .ZN(n3751) );
  NAND2_X1 U3795 ( .A1(n3385), .A2(n3474), .ZN(n3371) );
  XOR2_X1 U3796 ( .A(n5315), .B(n5316), .Z(n5346) );
  CLKBUF_X1 U3797 ( .A(n5662), .Z(n5671) );
  NOR2_X2 U3798 ( .A1(n5531), .A2(n5532), .ZN(n5477) );
  AOI22_X1 U3799 ( .A1(n3127), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5273), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3077) );
  NOR2_X2 U3800 ( .A1(n5585), .A2(n5612), .ZN(n5611) );
  NOR2_X2 U3801 ( .A1(n5300), .A2(n5301), .ZN(n5453) );
  AND2_X1 U3802 ( .A1(n5330), .A2(n5329), .ZN(n3033) );
  NAND2_X1 U3803 ( .A1(n3003), .A2(n3001), .ZN(n4270) );
  XNOR2_X1 U3804 ( .A(n3435), .B(n3436), .ZN(n3786) );
  AND2_X2 U3805 ( .A1(n4433), .A2(n4422), .ZN(n3154) );
  AND2_X1 U3806 ( .A1(n3191), .A2(n3182), .ZN(n3035) );
  OR2_X1 U3807 ( .A1(n4266), .A2(n4265), .ZN(n3036) );
  NOR2_X1 U3808 ( .A1(n5688), .A2(n3492), .ZN(n3037) );
  OR2_X1 U3809 ( .A1(n3204), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3038)
         );
  AND2_X1 U3810 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3039) );
  NAND2_X1 U3811 ( .A1(n3067), .A2(n3176), .ZN(n3171) );
  NAND2_X1 U3812 ( .A1(n3171), .A2(n3190), .ZN(n3210) );
  INV_X1 U3813 ( .A(n2995), .ZN(n3509) );
  NOR2_X1 U3814 ( .A1(n3577), .A2(n3182), .ZN(n3172) );
  AND2_X1 U3815 ( .A1(n3297), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3070) );
  INV_X1 U3816 ( .A(n3372), .ZN(n3283) );
  AOI22_X1 U3817 ( .A1(n3137), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3153), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3044) );
  AND2_X1 U3818 ( .A1(n6398), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3525)
         );
  OR2_X1 U3819 ( .A1(n3552), .A2(n3571), .ZN(n3532) );
  INV_X1 U3820 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3318) );
  INV_X1 U3821 ( .A(n3529), .ZN(n3545) );
  OR2_X1 U3822 ( .A1(n3523), .A2(n3522), .ZN(n3535) );
  INV_X1 U3823 ( .A(n3452), .ZN(n3450) );
  INV_X1 U3824 ( .A(n3153), .ZN(n3299) );
  OR2_X1 U3825 ( .A1(n3269), .A2(n3268), .ZN(n3387) );
  AND2_X1 U3826 ( .A1(n3449), .A2(n3448), .ZN(n3452) );
  AND2_X1 U3827 ( .A1(n4144), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4154)
         );
  AND2_X1 U3828 ( .A1(n3722), .A2(n5766), .ZN(n3723) );
  AND2_X1 U3829 ( .A1(n6051), .A2(n3486), .ZN(n3487) );
  NAND2_X1 U3830 ( .A1(n3296), .A2(n3295), .ZN(n3316) );
  INV_X1 U3831 ( .A(n3892), .ZN(n3906) );
  OR2_X1 U3832 ( .A1(n4696), .A2(n4695), .ZN(n5264) );
  NAND2_X1 U3833 ( .A1(n4154), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4177)
         );
  AND2_X1 U3834 ( .A1(n3990), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3991)
         );
  NOR2_X1 U3835 ( .A1(n3819), .A2(n5963), .ZN(n3814) );
  AND2_X1 U3836 ( .A1(n3410), .A2(n4961), .ZN(n3409) );
  AND2_X1 U3837 ( .A1(n3477), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3727)
         );
  NAND2_X1 U3838 ( .A1(n3278), .A2(n3381), .ZN(n3385) );
  NAND2_X1 U3839 ( .A1(n3326), .A2(n3325), .ZN(n4853) );
  NAND2_X1 U3840 ( .A1(n3557), .A2(n3556), .ZN(n3562) );
  INV_X1 U3841 ( .A(n5956), .ZN(n5997) );
  NAND2_X1 U3842 ( .A1(n4703), .A2(n4702), .ZN(n5327) );
  INV_X1 U3843 ( .A(n4234), .ZN(n4271) );
  NAND2_X1 U3844 ( .A1(n4042), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4089)
         );
  OR2_X1 U3845 ( .A1(n3495), .A2(n3494), .ZN(n5689) );
  NAND2_X1 U3846 ( .A1(n3814), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3851)
         );
  NAND2_X1 U3847 ( .A1(n3477), .A2(n3481), .ZN(n3482) );
  NOR2_X1 U3848 ( .A1(n5672), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3726)
         );
  INV_X1 U3849 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3503) );
  OR2_X1 U3850 ( .A1(n6134), .A2(n4446), .ZN(n4252) );
  AND2_X1 U3851 ( .A1(n3640), .A2(n3639), .ZN(n4346) );
  CLKBUF_X1 U3852 ( .A(n4303), .Z(n5818) );
  INV_X1 U3853 ( .A(n4480), .ZN(n4542) );
  INV_X1 U3854 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6403) );
  OAI211_X1 U3855 ( .C1(n6682), .C2(n5357), .A(n5356), .B(n5355), .ZN(n5358)
         );
  NOR2_X1 U3856 ( .A1(n6493), .A2(n5481), .ZN(n5852) );
  NOR2_X1 U3857 ( .A1(n6490), .A2(n5332), .ZN(n5925) );
  NOR2_X1 U3858 ( .A1(n6485), .A2(n5234), .ZN(n5498) );
  OR3_X1 U3859 ( .A1(n6538), .A2(n6185), .A3(n4694), .ZN(n4950) );
  INV_X1 U3860 ( .A(n5861), .ZN(n5983) );
  INV_X1 U3861 ( .A(n4950), .ZN(n4993) );
  INV_X1 U3862 ( .A(n4393), .ZN(n4372) );
  AOI22_X1 U3863 ( .A1(n5642), .A2(n5643), .B1(n3477), .B2(n3718), .ZN(n5637)
         );
  NAND2_X1 U3864 ( .A1(n3869), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3892)
         );
  NOR2_X1 U3865 ( .A1(n3792), .A2(n5978), .ZN(n3798) );
  NAND2_X1 U3866 ( .A1(n3769), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3768)
         );
  NOR2_X1 U3867 ( .A1(n5756), .A2(n4258), .ZN(n5751) );
  NOR2_X1 U3868 ( .A1(n5878), .A2(n3711), .ZN(n5789) );
  INV_X1 U3869 ( .A(n4252), .ZN(n6186) );
  AND2_X1 U3870 ( .A1(n3393), .A2(n3394), .ZN(n4444) );
  INV_X1 U3871 ( .A(n4658), .ZN(n4515) );
  INV_X1 U3872 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3205) );
  OR2_X1 U3873 ( .A1(n4520), .A2(n4519), .ZN(n6319) );
  INV_X1 U3874 ( .A(n6384), .ZN(n6369) );
  INV_X1 U3875 ( .A(n6396), .ZN(n6376) );
  INV_X1 U3876 ( .A(n5172), .ZN(n6388) );
  NAND2_X1 U3877 ( .A1(n4740), .A2(n4291), .ZN(n4691) );
  INV_X1 U3878 ( .A(n5986), .ZN(n5974) );
  NAND2_X1 U3879 ( .A1(n4950), .A2(n4699), .ZN(n5861) );
  INV_X1 U3880 ( .A(n6006), .ZN(n5553) );
  INV_X1 U3881 ( .A(n6017), .ZN(n6049) );
  NAND2_X1 U3882 ( .A1(n5302), .A2(n6081), .ZN(n5306) );
  OR2_X1 U3883 ( .A1(n5023), .A2(n5022), .ZN(n5966) );
  OR2_X1 U3884 ( .A1(n6076), .A2(n4408), .ZN(n6085) );
  AOI21_X1 U3885 ( .B1(n5302), .B2(n6183), .A(n3716), .ZN(n3717) );
  INV_X1 U3886 ( .A(n6087), .ZN(n5901) );
  INV_X1 U3887 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6398) );
  OR2_X1 U3888 ( .A1(n5136), .A2(n5810), .ZN(n6224) );
  OR2_X1 U3889 ( .A1(n6234), .A2(n6233), .ZN(n6311) );
  OR2_X1 U3890 ( .A1(n6329), .A2(n4859), .ZN(n4830) );
  INV_X1 U3891 ( .A(n3717), .ZN(U2995) );
  INV_X1 U3892 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3040) );
  NOR2_X4 U3893 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4433) );
  AOI22_X1 U3894 ( .A1(n3297), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3046) );
  AND2_X2 U3895 ( .A1(n3050), .A2(n3048), .ZN(n3135) );
  AND2_X2 U3896 ( .A1(n3048), .A2(n4423), .ZN(n3134) );
  AOI22_X1 U3897 ( .A1(n3135), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3045) );
  INV_X1 U3898 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3041) );
  INV_X1 U3899 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3042) );
  AOI22_X1 U3900 ( .A1(n3138), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3154), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3043) );
  AND2_X4 U3901 ( .A1(n3047), .A2(n4433), .ZN(n5273) );
  AND2_X2 U3902 ( .A1(n3049), .A2(n4423), .ZN(n3127) );
  AOI22_X1 U3903 ( .A1(n5273), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3054) );
  AOI22_X1 U3904 ( .A1(n3226), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3053) );
  AND2_X4 U3905 ( .A1(n4303), .A2(n4422), .ZN(n3244) );
  INV_X1 U3906 ( .A(n3123), .ZN(n3067) );
  AOI22_X1 U3907 ( .A1(n3129), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5273), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3060) );
  AOI22_X1 U3908 ( .A1(n3297), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3153), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3059) );
  AOI22_X1 U3909 ( .A1(n3263), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3058) );
  AOI22_X1 U3910 ( .A1(n3226), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3057) );
  AOI22_X1 U3911 ( .A1(n3137), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3064) );
  AOI22_X1 U3912 ( .A1(n3127), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3128), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3063) );
  AOI22_X1 U3913 ( .A1(n3138), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3154), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3062) );
  AOI22_X1 U3914 ( .A1(n3135), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3061) );
  AOI22_X1 U3915 ( .A1(n3137), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3153), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3069) );
  AOI22_X1 U3916 ( .A1(n3138), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3154), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3068) );
  AND2_X1 U3917 ( .A1(n3069), .A2(n3068), .ZN(n3072) );
  NAND3_X1 U3918 ( .A1(n3073), .A2(n3072), .A3(n3071), .ZN(n3079) );
  AOI22_X1 U3919 ( .A1(n3226), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3076) );
  AOI22_X1 U3920 ( .A1(n3129), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3128), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3075) );
  AOI22_X1 U3921 ( .A1(n3263), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3074) );
  NAND4_X1 U3922 ( .A1(n3077), .A2(n3076), .A3(n3075), .A4(n3074), .ZN(n3078)
         );
  AOI22_X1 U3923 ( .A1(n3137), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3153), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3084) );
  AOI22_X1 U3924 ( .A1(n3297), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3083) );
  AOI22_X1 U3925 ( .A1(n3135), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3082) );
  NAND4_X1 U3926 ( .A1(n3084), .A2(n3083), .A3(n3082), .A4(n3081), .ZN(n3090)
         );
  AOI22_X1 U3927 ( .A1(n3127), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5273), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3088) );
  AOI22_X1 U3928 ( .A1(n3226), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3087) );
  AOI22_X1 U3929 ( .A1(n3129), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3128), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3086) );
  AOI22_X1 U3930 ( .A1(n3263), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3085) );
  NAND4_X1 U3931 ( .A1(n3088), .A2(n3087), .A3(n3086), .A4(n3085), .ZN(n3089)
         );
  OR2_X2 U3932 ( .A1(n3090), .A2(n3089), .ZN(n4499) );
  NAND2_X1 U3933 ( .A1(n3297), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3094)
         );
  NAND2_X1 U3934 ( .A1(n3135), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3093) );
  NAND2_X1 U3935 ( .A1(n3134), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3092) );
  NAND2_X1 U3936 ( .A1(n3136), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3091) );
  NAND2_X1 U3937 ( .A1(n3226), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3099)
         );
  NAND2_X1 U3938 ( .A1(n3263), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3098) );
  NAND2_X1 U3939 ( .A1(n3095), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3097) );
  NAND2_X1 U3940 ( .A1(n3244), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3096)
         );
  NAND2_X1 U3941 ( .A1(n3020), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3102)
         );
  NAND2_X1 U3942 ( .A1(n3023), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3101) );
  NAND2_X1 U3943 ( .A1(n3021), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3100)
         );
  NAND3_X1 U3944 ( .A1(n3102), .A2(n3101), .A3(n3100), .ZN(n3103) );
  NAND2_X1 U3945 ( .A1(n3129), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3107) );
  NAND2_X1 U3946 ( .A1(n5273), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3106) );
  NAND2_X1 U3947 ( .A1(n3127), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3105) );
  NAND2_X1 U3948 ( .A1(n3128), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3104) );
  INV_X1 U3949 ( .A(n3175), .ZN(n3112) );
  NAND2_X1 U3950 ( .A1(n3113), .A2(n3112), .ZN(n3207) );
  AOI22_X1 U3951 ( .A1(n5273), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3128), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3117) );
  AOI22_X1 U3952 ( .A1(n3134), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3153), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3115) );
  AOI22_X1 U3953 ( .A1(n3263), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3114) );
  AOI22_X1 U3954 ( .A1(n3137), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3121) );
  AOI22_X1 U3955 ( .A1(n3138), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3120) );
  AOI22_X1 U3956 ( .A1(n3226), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3119) );
  AOI22_X1 U3957 ( .A1(n3297), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3118) );
  NAND2_X2 U3958 ( .A1(n3178), .A2(n2990), .ZN(n3173) );
  NAND3_X1 U3959 ( .A1(n3207), .A2(n3580), .A3(n3173), .ZN(n3124) );
  AND2_X2 U3960 ( .A1(n3125), .A2(n3124), .ZN(n3586) );
  NAND2_X1 U3961 ( .A1(n3126), .A2(n3173), .ZN(n3587) );
  AOI22_X1 U3962 ( .A1(n5273), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3133) );
  AOI22_X1 U3963 ( .A1(n3226), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3132) );
  AOI22_X1 U3964 ( .A1(n3129), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3128), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3131) );
  AOI22_X1 U3965 ( .A1(n3263), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3130) );
  AOI22_X1 U3966 ( .A1(n3135), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3142) );
  AOI22_X1 U3967 ( .A1(n3297), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3136), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3141) );
  AOI22_X1 U3968 ( .A1(n3137), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3153), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3140) );
  AOI22_X1 U3969 ( .A1(n3138), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3154), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3139) );
  AOI21_X1 U3970 ( .B1(n3587), .B2(n3189), .A(n4492), .ZN(n3144) );
  NAND2_X1 U3971 ( .A1(n3586), .A2(n3144), .ZN(n3167) );
  NAND2_X1 U3972 ( .A1(n3138), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3148)
         );
  NAND2_X1 U3973 ( .A1(n3135), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3147) );
  NAND2_X1 U3974 ( .A1(n3297), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3146)
         );
  NAND2_X1 U3975 ( .A1(n3137), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3145) );
  NAND2_X1 U3976 ( .A1(n3226), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3152)
         );
  NAND2_X1 U3977 ( .A1(n3129), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3151) );
  NAND2_X1 U3978 ( .A1(n3263), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3150) );
  NAND2_X1 U3979 ( .A1(n3244), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3149)
         );
  NAND2_X1 U3980 ( .A1(n3134), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3158) );
  NAND2_X1 U3981 ( .A1(n3136), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3157) );
  NAND2_X1 U3982 ( .A1(n3153), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3156)
         );
  NAND2_X1 U3983 ( .A1(n3154), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3155)
         );
  NAND2_X1 U3984 ( .A1(n5273), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3162) );
  NAND2_X1 U3985 ( .A1(n3127), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3161) );
  NAND2_X1 U3986 ( .A1(n3095), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3160) );
  NAND2_X1 U3987 ( .A1(n3128), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3159) );
  NAND2_X1 U3988 ( .A1(n3167), .A2(n3251), .ZN(n3217) );
  INV_X1 U3989 ( .A(n3171), .ZN(n3168) );
  NAND2_X1 U3990 ( .A1(n3168), .A2(n3175), .ZN(n3169) );
  NAND2_X1 U3991 ( .A1(n3183), .A2(n3169), .ZN(n3605) );
  INV_X1 U3992 ( .A(n3605), .ZN(n3170) );
  NAND2_X1 U3993 ( .A1(n3170), .A2(n3190), .ZN(n3579) );
  INV_X1 U3994 ( .A(n3171), .ZN(n3577) );
  NOR2_X2 U3995 ( .A1(n3579), .A2(n3172), .ZN(n3220) );
  NAND3_X1 U3996 ( .A1(n3583), .A2(n3182), .A3(n4499), .ZN(n3174) );
  AND2_X4 U3997 ( .A1(n3187), .A2(n3604), .ZN(n3359) );
  NAND2_X1 U3998 ( .A1(n3174), .A2(n3359), .ZN(n3177) );
  NAND2_X1 U3999 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6457) );
  OAI21_X1 U4000 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6457), .ZN(n3564) );
  NAND2_X1 U4001 ( .A1(n3187), .A2(n3564), .ZN(n3186) );
  AOI21_X1 U4002 ( .B1(n3186), .B2(n3191), .A(n3189), .ZN(n3179) );
  NAND4_X1 U4003 ( .A1(n3217), .A2(n3214), .A3(n3220), .A4(n3179), .ZN(n3180)
         );
  INV_X1 U4004 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3181) );
  NAND2_X1 U4005 ( .A1(n3580), .A2(n3190), .ZN(n3376) );
  NAND3_X1 U4006 ( .A1(n3035), .A2(n3184), .A3(n3183), .ZN(n3563) );
  INV_X1 U4007 ( .A(n3563), .ZN(n3185) );
  INV_X1 U4008 ( .A(n3186), .ZN(n3195) );
  NOR2_X1 U4009 ( .A1(n3587), .A2(n3510), .ZN(n3188) );
  NAND2_X1 U4010 ( .A1(n3192), .A2(n3596), .ZN(n3600) );
  INV_X1 U4011 ( .A(n3600), .ZN(n3194) );
  NAND2_X1 U4012 ( .A1(n4503), .A2(n4499), .ZN(n5258) );
  NAND2_X1 U4013 ( .A1(n3196), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3203) );
  NOR2_X1 U4014 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6522) );
  NAND2_X1 U4015 ( .A1(n6522), .A2(n6536), .ZN(n4211) );
  INV_X1 U4016 ( .A(n4211), .ZN(n3324) );
  NAND2_X1 U4017 ( .A1(n6398), .A2(n6403), .ZN(n3197) );
  NAND2_X1 U4018 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3293) );
  AND2_X1 U4019 ( .A1(n3197), .A2(n3293), .ZN(n4654) );
  NAND2_X1 U4020 ( .A1(n3324), .A2(n4654), .ZN(n3199) );
  INV_X1 U4021 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5340) );
  AND2_X1 U4022 ( .A1(n5340), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3589) );
  INV_X1 U4023 ( .A(n3589), .ZN(n3323) );
  NAND2_X1 U4024 ( .A1(n3323), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3198) );
  NAND2_X1 U4025 ( .A1(n3199), .A2(n3198), .ZN(n3204) );
  INV_X1 U4026 ( .A(n3204), .ZN(n3200) );
  MUX2_X1 U4027 ( .A(n3589), .B(n4211), .S(n6398), .Z(n3206) );
  OAI21_X2 U4028 ( .B1(n3290), .B2(n3205), .A(n3206), .ZN(n3258) );
  NAND2_X1 U4029 ( .A1(n6522), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6439) );
  AOI21_X1 U4030 ( .B1(n3189), .B2(n3602), .A(n6439), .ZN(n3213) );
  INV_X1 U4031 ( .A(n3207), .ZN(n3209) );
  NAND2_X1 U4032 ( .A1(n3209), .A2(n3208), .ZN(n3212) );
  NAND2_X1 U4033 ( .A1(n3210), .A2(n3359), .ZN(n3211) );
  NAND3_X1 U4034 ( .A1(n3213), .A2(n3212), .A3(n3211), .ZN(n3216) );
  INV_X1 U4035 ( .A(n3214), .ZN(n3215) );
  AND2_X2 U4036 ( .A1(n4492), .A2(n5259), .ZN(n3520) );
  NAND2_X1 U4037 ( .A1(n3520), .A2(n3175), .ZN(n3219) );
  NAND2_X1 U4038 ( .A1(n2991), .A2(n3219), .ZN(n3612) );
  INV_X1 U4039 ( .A(n3220), .ZN(n3221) );
  NAND2_X1 U4040 ( .A1(n3221), .A2(n4492), .ZN(n3222) );
  NAND3_X1 U4041 ( .A1(n3223), .A2(n3612), .A3(n3222), .ZN(n3256) );
  NAND2_X1 U4042 ( .A1(n4465), .A2(n6536), .ZN(n3238) );
  AOI22_X1 U4043 ( .A1(n2985), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3230) );
  AOI22_X1 U4044 ( .A1(n5274), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3229) );
  AOI22_X1 U4046 ( .A1(n5277), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3228) );
  AOI22_X1 U4048 ( .A1(n4189), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3227) );
  NAND4_X1 U4049 ( .A1(n3230), .A2(n3229), .A3(n3228), .A4(n3227), .ZN(n3236)
         );
  AOI22_X1 U4050 ( .A1(n2984), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3234) );
  AOI22_X1 U4051 ( .A1(n2986), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3233) );
  AOI22_X1 U4052 ( .A1(n4121), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3232) );
  INV_X1 U4053 ( .A(n3137), .ZN(n3298) );
  AOI22_X1 U4054 ( .A1(n5275), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3231) );
  NAND4_X1 U4055 ( .A1(n3234), .A2(n3233), .A3(n3232), .A4(n3231), .ZN(n3235)
         );
  INV_X1 U4056 ( .A(n3375), .ZN(n3252) );
  INV_X1 U4057 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3255) );
  AOI22_X1 U4058 ( .A1(n2984), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3243) );
  AOI22_X1 U4059 ( .A1(n4194), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3242) );
  AOI22_X1 U4060 ( .A1(n3137), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3241) );
  AOI22_X1 U4061 ( .A1(n3239), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3240) );
  NAND4_X1 U4062 ( .A1(n3243), .A2(n3242), .A3(n3241), .A4(n3240), .ZN(n3250)
         );
  AOI22_X1 U4063 ( .A1(n4121), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3248) );
  AOI22_X1 U4064 ( .A1(n4189), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3247) );
  AOI22_X1 U4065 ( .A1(n3129), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3128), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3246) );
  AOI22_X1 U4066 ( .A1(n2986), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3245) );
  NAND4_X1 U4067 ( .A1(n3248), .A2(n3247), .A3(n3246), .A4(n3245), .ZN(n3249)
         );
  NOR2_X1 U4068 ( .A1(n3328), .A2(n3479), .ZN(n3270) );
  INV_X1 U4069 ( .A(n3270), .ZN(n3254) );
  OR2_X1 U4070 ( .A1(n3327), .A2(n3252), .ZN(n3253) );
  NAND2_X1 U4071 ( .A1(n3372), .A2(n3370), .ZN(n3281) );
  INV_X1 U4072 ( .A(n3256), .ZN(n3257) );
  XNOR2_X1 U4073 ( .A(n3258), .B(n3257), .ZN(n3753) );
  NAND2_X1 U4074 ( .A1(n3753), .A2(n6536), .ZN(n3274) );
  AOI22_X1 U4075 ( .A1(n4194), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3262) );
  AOI22_X1 U4076 ( .A1(n4121), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3261) );
  AOI22_X1 U4077 ( .A1(n2985), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3260) );
  AOI22_X1 U4078 ( .A1(n3137), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3259) );
  NAND4_X1 U4079 ( .A1(n3262), .A2(n3261), .A3(n3260), .A4(n3259), .ZN(n3269)
         );
  AOI22_X1 U4080 ( .A1(n2984), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3267) );
  BUF_X1 U4081 ( .A(n3138), .Z(n5277) );
  AOI22_X1 U4082 ( .A1(n5277), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3266) );
  AOI22_X1 U4083 ( .A1(n4189), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3265) );
  AOI22_X1 U4084 ( .A1(n2986), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3264) );
  NAND4_X1 U4085 ( .A1(n3267), .A2(n3266), .A3(n3265), .A4(n3264), .ZN(n3268)
         );
  NAND2_X1 U4086 ( .A1(n3270), .A2(n3387), .ZN(n3382) );
  NAND2_X1 U4087 ( .A1(n3175), .A2(n3479), .ZN(n3276) );
  INV_X1 U4088 ( .A(n3387), .ZN(n3271) );
  NAND2_X1 U4089 ( .A1(n3279), .A2(n3271), .ZN(n3272) );
  AND2_X1 U4090 ( .A1(n3382), .A2(n3272), .ZN(n3273) );
  NAND2_X1 U4091 ( .A1(n3274), .A2(n3273), .ZN(n3278) );
  INV_X1 U4092 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3277) );
  OAI21_X1 U4093 ( .B1(n3387), .B2(n6536), .A(n3508), .ZN(n3275) );
  OAI211_X1 U4094 ( .C1(n3529), .C2(n3277), .A(n3276), .B(n3275), .ZN(n3381)
         );
  INV_X1 U4095 ( .A(n3279), .ZN(n3474) );
  INV_X1 U4096 ( .A(n3371), .ZN(n3280) );
  NAND2_X1 U4097 ( .A1(n3281), .A2(n3280), .ZN(n3285) );
  NAND2_X1 U4098 ( .A1(n3283), .A2(n3282), .ZN(n3284) );
  NAND2_X1 U4099 ( .A1(n3285), .A2(n3284), .ZN(n3396) );
  INV_X1 U4100 ( .A(n3396), .ZN(n3314) );
  INV_X1 U4101 ( .A(n3293), .ZN(n3292) );
  NAND2_X1 U4102 ( .A1(n3292), .A2(n5135), .ZN(n6324) );
  NAND2_X1 U4103 ( .A1(n3293), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3294) );
  NAND2_X1 U4104 ( .A1(n6324), .A2(n3294), .ZN(n4514) );
  AOI22_X1 U4105 ( .A1(n3324), .A2(n4514), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3323), .ZN(n3295) );
  AOI22_X1 U4106 ( .A1(n2984), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U4107 ( .A1(n4194), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3302) );
  INV_X2 U4108 ( .A(n3299), .ZN(n5265) );
  AOI22_X1 U4109 ( .A1(n5275), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4110 ( .A1(n5277), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3300) );
  NAND4_X1 U4111 ( .A1(n3303), .A2(n3302), .A3(n3301), .A4(n3300), .ZN(n3309)
         );
  AOI22_X1 U4112 ( .A1(n5273), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U4113 ( .A1(n4189), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4114 ( .A1(n3129), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3305) );
  AOI22_X1 U4115 ( .A1(n2986), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3304) );
  NAND4_X1 U4116 ( .A1(n3307), .A2(n3306), .A3(n3305), .A4(n3304), .ZN(n3308)
         );
  NOR2_X1 U4117 ( .A1(n3328), .A2(n3356), .ZN(n3310) );
  INV_X1 U4118 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3311) );
  OAI22_X1 U4119 ( .A1(n3529), .A2(n3311), .B1(n3327), .B2(n3356), .ZN(n3312)
         );
  NAND2_X1 U4120 ( .A1(n3314), .A2(n3397), .ZN(n3364) );
  INV_X1 U4121 ( .A(n3364), .ZN(n3343) );
  NAND3_X1 U4122 ( .A1(n6409), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6280) );
  INV_X1 U4123 ( .A(n6280), .ZN(n3321) );
  NAND2_X1 U4124 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3321), .ZN(n6272) );
  NAND2_X1 U4125 ( .A1(n6409), .A2(n6272), .ZN(n3322) );
  NOR3_X1 U4126 ( .A1(n6409), .A2(n5135), .A3(n6403), .ZN(n4544) );
  NAND2_X1 U4127 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4544), .ZN(n4467) );
  AND2_X1 U4128 ( .A1(n3322), .A2(n4467), .ZN(n4653) );
  AOI22_X1 U4129 ( .A1(n3324), .A2(n4653), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3323), .ZN(n3325) );
  AOI22_X1 U4130 ( .A1(n5277), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5275), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3332) );
  AOI22_X1 U4131 ( .A1(n5274), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4132 ( .A1(n2986), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4133 ( .A1(n4189), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3329) );
  NAND4_X1 U4134 ( .A1(n3332), .A2(n3331), .A3(n3330), .A4(n3329), .ZN(n3338)
         );
  AOI22_X1 U4135 ( .A1(n2984), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4136 ( .A1(n4121), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4137 ( .A1(n2985), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4138 ( .A1(n5265), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3333) );
  NAND4_X1 U4139 ( .A1(n3336), .A2(n3335), .A3(n3334), .A4(n3333), .ZN(n3337)
         );
  INV_X1 U4140 ( .A(n3357), .ZN(n3365) );
  INV_X1 U4141 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3339) );
  OAI22_X1 U4142 ( .A1(n3552), .A2(n3365), .B1(n3339), .B2(n3529), .ZN(n3340)
         );
  INV_X1 U4143 ( .A(n3340), .ZN(n3341) );
  NAND2_X1 U4144 ( .A1(n3343), .A2(n4480), .ZN(n3412) );
  AOI22_X1 U4145 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n2984), .B1(n4187), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3347) );
  AOI22_X1 U4146 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4194), .B1(n5274), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3346) );
  AOI22_X1 U4147 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n5275), .B1(n5265), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3345) );
  AOI22_X1 U4148 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n5277), .B1(n5266), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3344) );
  NAND4_X1 U4149 ( .A1(n3347), .A2(n3346), .A3(n3345), .A4(n3344), .ZN(n3353)
         );
  AOI22_X1 U4150 ( .A1(n4121), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3351) );
  AOI22_X1 U4151 ( .A1(n4189), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3350) );
  AOI22_X1 U4152 ( .A1(n2985), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3349) );
  AOI22_X1 U4153 ( .A1(n2986), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3348) );
  NAND4_X1 U4154 ( .A1(n3351), .A2(n3350), .A3(n3349), .A4(n3348), .ZN(n3352)
         );
  OR2_X1 U4155 ( .A1(n3353), .A2(n3352), .ZN(n3358) );
  INV_X1 U4156 ( .A(n3358), .ZN(n3428) );
  OR2_X1 U4157 ( .A1(n3552), .A2(n3428), .ZN(n3355) );
  NAND2_X1 U4158 ( .A1(n3545), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3354) );
  NAND2_X1 U4159 ( .A1(n3355), .A2(n3354), .ZN(n3413) );
  XNOR2_X1 U4160 ( .A(n3412), .B(n3413), .ZN(n3775) );
  NAND2_X1 U4161 ( .A1(n3775), .A2(n3520), .ZN(n3362) );
  NAND2_X1 U4162 ( .A1(n3375), .A2(n3387), .ZN(n3399) );
  NAND2_X1 U4163 ( .A1(n3399), .A2(n3356), .ZN(n3366) );
  NAND2_X1 U4164 ( .A1(n3366), .A2(n3357), .ZN(n3429) );
  XNOR2_X1 U4165 ( .A(n3429), .B(n3358), .ZN(n3360) );
  NAND2_X1 U4166 ( .A1(n3360), .A2(n3359), .ZN(n3361) );
  INV_X1 U4167 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6168) );
  INV_X1 U4168 ( .A(n4962), .ZN(n3411) );
  NAND2_X1 U4169 ( .A1(n3363), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3410)
         );
  XNOR2_X1 U4170 ( .A(n3364), .B(n4480), .ZN(n3767) );
  NAND2_X1 U4171 ( .A1(n3767), .A2(n3520), .ZN(n3369) );
  XNOR2_X1 U4172 ( .A(n3366), .B(n3365), .ZN(n3367) );
  NAND2_X1 U4173 ( .A1(n3367), .A2(n3359), .ZN(n3368) );
  NAND2_X1 U4174 ( .A1(n3369), .A2(n3368), .ZN(n3408) );
  NAND2_X1 U4175 ( .A1(n3408), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4961)
         );
  NAND2_X1 U4177 ( .A1(n4471), .A2(n3520), .ZN(n3380) );
  OAI21_X1 U4178 ( .B1(n3387), .B2(n3375), .A(n3399), .ZN(n3377) );
  INV_X1 U4179 ( .A(n3359), .ZN(n3631) );
  OAI211_X1 U4180 ( .C1(n3377), .C2(n3631), .A(n3184), .B(n5259), .ZN(n3378)
         );
  INV_X1 U4181 ( .A(n3378), .ZN(n3379) );
  NAND2_X1 U4182 ( .A1(n3380), .A2(n3379), .ZN(n4445) );
  INV_X1 U4183 ( .A(n3381), .ZN(n3383) );
  NAND2_X1 U4184 ( .A1(n3383), .A2(n3382), .ZN(n3384) );
  INV_X1 U4185 ( .A(n3751), .ZN(n3386) );
  NAND2_X1 U4186 ( .A1(n3386), .A2(n3520), .ZN(n3390) );
  NAND2_X1 U4187 ( .A1(n3251), .A2(n3190), .ZN(n3400) );
  OAI21_X1 U4188 ( .B1(n3631), .B2(n3387), .A(n3400), .ZN(n3388) );
  INV_X1 U4189 ( .A(n3388), .ZN(n3389) );
  NAND2_X1 U4190 ( .A1(n3390), .A2(n3389), .ZN(n4402) );
  NAND2_X1 U4191 ( .A1(n4402), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3391)
         );
  INV_X1 U4192 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4447) );
  NAND2_X1 U4193 ( .A1(n3391), .A2(n4447), .ZN(n3393) );
  AND2_X1 U4194 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3392) );
  NAND2_X1 U4195 ( .A1(n4402), .A2(n3392), .ZN(n3394) );
  NAND2_X1 U4196 ( .A1(n4445), .A2(n4444), .ZN(n3395) );
  NAND2_X1 U4197 ( .A1(n3395), .A2(n3394), .ZN(n6077) );
  NAND2_X1 U4198 ( .A1(n6077), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3403)
         );
  XNOR2_X1 U4199 ( .A(n3399), .B(n3398), .ZN(n3401) );
  OAI21_X1 U4200 ( .B1(n3401), .B2(n3631), .A(n3400), .ZN(n3402) );
  AOI21_X1 U4201 ( .B1(n4470), .B2(n3520), .A(n3402), .ZN(n6078) );
  NAND2_X1 U4202 ( .A1(n3403), .A2(n6078), .ZN(n3407) );
  INV_X1 U4203 ( .A(n6077), .ZN(n3405) );
  INV_X1 U4204 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3404) );
  NAND2_X1 U4205 ( .A1(n3405), .A2(n3404), .ZN(n3406) );
  AND2_X1 U4206 ( .A1(n3407), .A2(n3406), .ZN(n6069) );
  INV_X1 U4207 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6174) );
  XNOR2_X1 U4208 ( .A(n3408), .B(n6174), .ZN(n6070) );
  INV_X1 U4209 ( .A(n3412), .ZN(n3414) );
  NAND2_X1 U4210 ( .A1(n3414), .A2(n3413), .ZN(n3435) );
  AOI22_X1 U4211 ( .A1(n4189), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n2986), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3418) );
  AOI22_X1 U4212 ( .A1(n2984), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3417) );
  AOI22_X1 U4213 ( .A1(n5275), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3416) );
  AOI22_X1 U4214 ( .A1(n4121), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3415) );
  NAND4_X1 U4215 ( .A1(n3418), .A2(n3417), .A3(n3416), .A4(n3415), .ZN(n3424)
         );
  AOI22_X1 U4216 ( .A1(n5277), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3422) );
  AOI22_X1 U4217 ( .A1(n5276), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3421) );
  AOI22_X1 U4218 ( .A1(n2985), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3420) );
  AOI22_X1 U4219 ( .A1(n4188), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3419) );
  NAND4_X1 U4220 ( .A1(n3422), .A2(n3421), .A3(n3420), .A4(n3419), .ZN(n3423)
         );
  OR2_X1 U4221 ( .A1(n3424), .A2(n3423), .ZN(n3455) );
  INV_X1 U4222 ( .A(n3455), .ZN(n3425) );
  OR2_X1 U4223 ( .A1(n3552), .A2(n3425), .ZN(n3427) );
  NAND2_X1 U4224 ( .A1(n3545), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3426) );
  NAND2_X1 U4225 ( .A1(n3427), .A2(n3426), .ZN(n3436) );
  NAND2_X1 U4226 ( .A1(n3786), .A2(n3520), .ZN(n3432) );
  OR2_X1 U4227 ( .A1(n3429), .A2(n3428), .ZN(n3454) );
  XNOR2_X1 U4228 ( .A(n3454), .B(n3455), .ZN(n3430) );
  NAND2_X1 U4229 ( .A1(n3430), .A2(n3359), .ZN(n3431) );
  NAND2_X1 U4230 ( .A1(n3432), .A2(n3431), .ZN(n3433) );
  INV_X1 U4231 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6144) );
  XNOR2_X1 U4232 ( .A(n3433), .B(n6144), .ZN(n4935) );
  NAND2_X1 U4233 ( .A1(n4932), .A2(n4935), .ZN(n4934) );
  NAND2_X1 U4234 ( .A1(n3433), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3434)
         );
  NAND2_X1 U4235 ( .A1(n2987), .A2(n3436), .ZN(n3453) );
  INV_X1 U4236 ( .A(n3453), .ZN(n3451) );
  AOI22_X1 U4237 ( .A1(n2984), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3440) );
  AOI22_X1 U4238 ( .A1(n4194), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3439) );
  AOI22_X1 U4239 ( .A1(n5275), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3438) );
  AOI22_X1 U4240 ( .A1(n5277), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3437) );
  NAND4_X1 U4241 ( .A1(n3440), .A2(n3439), .A3(n3438), .A4(n3437), .ZN(n3446)
         );
  AOI22_X1 U4242 ( .A1(n4121), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4243 ( .A1(n4189), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4244 ( .A1(n2985), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3442) );
  AOI22_X1 U4245 ( .A1(n2986), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3441) );
  NAND4_X1 U4246 ( .A1(n3444), .A2(n3443), .A3(n3442), .A4(n3441), .ZN(n3445)
         );
  OR2_X1 U4247 ( .A1(n3446), .A2(n3445), .ZN(n3466) );
  INV_X1 U4248 ( .A(n3466), .ZN(n3447) );
  OR2_X1 U4249 ( .A1(n3552), .A2(n3447), .ZN(n3449) );
  NAND2_X1 U4250 ( .A1(n3545), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3448) );
  NAND2_X2 U4251 ( .A1(n3451), .A2(n3450), .ZN(n3476) );
  NAND2_X1 U4252 ( .A1(n3453), .A2(n3452), .ZN(n3791) );
  NAND3_X1 U4253 ( .A1(n3476), .A2(n3791), .A3(n3520), .ZN(n3459) );
  INV_X1 U4254 ( .A(n3454), .ZN(n3456) );
  NAND2_X1 U4255 ( .A1(n3456), .A2(n3455), .ZN(n3465) );
  XNOR2_X1 U4256 ( .A(n3465), .B(n3466), .ZN(n3457) );
  NAND2_X1 U4257 ( .A1(n3457), .A2(n3359), .ZN(n3458) );
  NAND2_X1 U4258 ( .A1(n3459), .A2(n3458), .ZN(n3460) );
  INV_X1 U4259 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6143) );
  XNOR2_X1 U4260 ( .A(n3460), .B(n6143), .ZN(n6062) );
  NAND2_X1 U4261 ( .A1(n6063), .A2(n6062), .ZN(n6061) );
  NAND2_X1 U4262 ( .A1(n3460), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3461)
         );
  NAND2_X1 U4263 ( .A1(n6061), .A2(n3461), .ZN(n4943) );
  INV_X1 U4264 ( .A(n3479), .ZN(n3463) );
  INV_X1 U4265 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3462) );
  OAI22_X1 U4266 ( .A1(n3552), .A2(n3463), .B1(n3462), .B2(n3529), .ZN(n3464)
         );
  NAND2_X1 U4267 ( .A1(n3803), .A2(n3520), .ZN(n3470) );
  INV_X1 U4268 ( .A(n3465), .ZN(n3467) );
  NAND2_X1 U4269 ( .A1(n3467), .A2(n3466), .ZN(n3478) );
  XNOR2_X1 U4270 ( .A(n3478), .B(n3479), .ZN(n3468) );
  NAND2_X1 U4271 ( .A1(n3468), .A2(n3359), .ZN(n3469) );
  NAND2_X1 U4272 ( .A1(n3470), .A2(n3469), .ZN(n3471) );
  INV_X1 U4273 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6130) );
  XNOR2_X1 U4274 ( .A(n3471), .B(n6130), .ZN(n4942) );
  NAND2_X1 U4275 ( .A1(n4943), .A2(n4942), .ZN(n4941) );
  NAND2_X1 U4276 ( .A1(n3471), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3472)
         );
  NAND2_X1 U4277 ( .A1(n4941), .A2(n3472), .ZN(n4986) );
  INV_X1 U4278 ( .A(n3520), .ZN(n3473) );
  NOR2_X1 U4279 ( .A1(n3474), .A2(n3473), .ZN(n3475) );
  INV_X1 U4280 ( .A(n3478), .ZN(n3480) );
  NAND3_X1 U4281 ( .A1(n3480), .A2(n3359), .A3(n3479), .ZN(n3481) );
  INV_X1 U4282 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6121) );
  XNOR2_X1 U4283 ( .A(n3482), .B(n6121), .ZN(n4985) );
  NAND2_X1 U4284 ( .A1(n3482), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3483)
         );
  NAND2_X1 U4285 ( .A1(n4984), .A2(n3483), .ZN(n5032) );
  INV_X1 U4286 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U4287 ( .A1(n3477), .A2(n6093), .ZN(n5033) );
  INV_X1 U4288 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3484) );
  NAND2_X1 U4289 ( .A1(n3477), .A2(n3484), .ZN(n5068) );
  NAND2_X1 U4290 ( .A1(n2988), .A2(n2996), .ZN(n6052) );
  INV_X1 U4291 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3485) );
  NAND2_X1 U4292 ( .A1(n5672), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U4293 ( .A1(n5672), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3486) );
  OAI21_X2 U4294 ( .B1(n6052), .B2(n3488), .A(n3487), .ZN(n5105) );
  INV_X1 U4295 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5118) );
  NAND2_X1 U4296 ( .A1(n3477), .A2(n5118), .ZN(n5107) );
  OAI21_X1 U4297 ( .B1(n5105), .B2(n5109), .A(n5107), .ZN(n5868) );
  XNOR2_X1 U4298 ( .A(n3477), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5869)
         );
  NAND2_X1 U4299 ( .A1(n5868), .A2(n5869), .ZN(n3491) );
  INV_X1 U4300 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3489) );
  NAND2_X1 U4301 ( .A1(n3477), .A2(n3489), .ZN(n3490) );
  NAND2_X1 U4302 ( .A1(n3491), .A2(n3490), .ZN(n5191) );
  INV_X1 U4303 ( .A(n5191), .ZN(n3497) );
  INV_X1 U4304 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5193) );
  AND2_X1 U4305 ( .A1(n3477), .A2(n5193), .ZN(n5663) );
  INV_X1 U4306 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5893) );
  INV_X1 U4307 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3498) );
  AND2_X1 U4308 ( .A1(n3477), .A2(n3498), .ZN(n3492) );
  NAND2_X1 U4309 ( .A1(n5672), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5664) );
  XNOR2_X1 U4310 ( .A(n3477), .B(n5893), .ZN(n5698) );
  INV_X1 U4311 ( .A(n5698), .ZN(n3493) );
  AOI21_X1 U4312 ( .B1(n3497), .B2(n3037), .A(n3496), .ZN(n5662) );
  INV_X1 U4313 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5796) );
  INV_X1 U4314 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5801) );
  AND3_X1 U4315 ( .A1(n3498), .A2(n5796), .A3(n5801), .ZN(n3499) );
  AOI21_X1 U4316 ( .B1(n5662), .B2(n3499), .A(n3477), .ZN(n3500) );
  INV_X1 U4317 ( .A(n3500), .ZN(n3501) );
  NAND2_X1 U4318 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3711) );
  INV_X1 U4319 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U4320 ( .A1(n3477), .A2(n5788), .ZN(n5651) );
  NOR2_X1 U4321 ( .A1(n3477), .A2(n5788), .ZN(n5655) );
  NOR2_X1 U4322 ( .A1(n5650), .A2(n5655), .ZN(n5642) );
  XNOR2_X1 U4323 ( .A(n3477), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5643)
         );
  INV_X1 U4324 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3718) );
  XNOR2_X1 U4325 ( .A(n3477), .B(n3018), .ZN(n5636) );
  NOR2_X1 U4326 ( .A1(n5637), .A2(n5636), .ZN(n5635) );
  NOR2_X1 U4327 ( .A1(n3477), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5629)
         );
  NAND2_X1 U4328 ( .A1(n5635), .A2(n5629), .ZN(n5621) );
  AND2_X1 U4329 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5766) );
  NAND4_X1 U4330 ( .A1(n3000), .A2(n5766), .A3(INSTADDRPOINTER_REG_20__SCAN_IN), .A4(n3477), .ZN(n3502) );
  NAND2_X1 U4331 ( .A1(n5621), .A2(n3502), .ZN(n3504) );
  NAND2_X1 U4332 ( .A1(n3505), .A2(n5259), .ZN(n3515) );
  XNOR2_X1 U4333 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3524) );
  INV_X1 U4334 ( .A(n3524), .ZN(n3506) );
  XNOR2_X1 U4335 ( .A(n3506), .B(n3525), .ZN(n3569) );
  AND2_X1 U4336 ( .A1(n3569), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3516) );
  AND2_X1 U4337 ( .A1(n3205), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3507)
         );
  NOR2_X1 U4338 ( .A1(n3525), .A2(n3507), .ZN(n3513) );
  AOI21_X1 U4339 ( .B1(n3509), .B2(n3513), .A(n3508), .ZN(n3512) );
  NAND2_X1 U4340 ( .A1(n3187), .A2(n5259), .ZN(n3511) );
  NAND2_X1 U4341 ( .A1(n3510), .A2(n3511), .ZN(n3528) );
  OAI22_X1 U4342 ( .A1(n3515), .A2(n3516), .B1(n3512), .B2(n3528), .ZN(n3521)
         );
  INV_X1 U4343 ( .A(n3513), .ZN(n3514) );
  OR2_X1 U4344 ( .A1(n3552), .A2(n3514), .ZN(n3519) );
  INV_X1 U4345 ( .A(n3515), .ZN(n3518) );
  INV_X1 U4346 ( .A(n3516), .ZN(n3517) );
  OAI22_X1 U4347 ( .A1(n3521), .A2(n3519), .B1(n3518), .B2(n3517), .ZN(n3523)
         );
  NAND2_X1 U4348 ( .A1(n3545), .A2(n3520), .ZN(n3558) );
  AOI21_X1 U4349 ( .B1(n3521), .B2(n3569), .A(n3558), .ZN(n3522) );
  NAND2_X1 U4350 ( .A1(n3525), .A2(n3524), .ZN(n3527) );
  NAND2_X1 U4351 ( .A1(n6403), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3526) );
  NAND2_X1 U4352 ( .A1(n3527), .A2(n3526), .ZN(n3537) );
  XNOR2_X1 U4353 ( .A(n4416), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3536)
         );
  XNOR2_X1 U4354 ( .A(n3537), .B(n3536), .ZN(n3571) );
  INV_X1 U4355 ( .A(n3571), .ZN(n3530) );
  INV_X1 U4356 ( .A(n3528), .ZN(n3531) );
  OAI211_X1 U4357 ( .C1(n3530), .C2(n3529), .A(n3532), .B(n3531), .ZN(n3534)
         );
  NOR2_X1 U4358 ( .A1(n3532), .A2(n3531), .ZN(n3533) );
  AOI21_X1 U4359 ( .B1(n3535), .B2(n3534), .A(n3533), .ZN(n3547) );
  NAND2_X1 U4360 ( .A1(n3537), .A2(n3536), .ZN(n3539) );
  NAND2_X1 U4361 ( .A1(n5135), .A2(n4416), .ZN(n3538) );
  NAND2_X1 U4362 ( .A1(n3539), .A2(n3538), .ZN(n3542) );
  XNOR2_X1 U4363 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3541) );
  NOR2_X1 U4364 ( .A1(n3319), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3540)
         );
  AOI21_X1 U4365 ( .B1(n3542), .B2(n3541), .A(n3540), .ZN(n3549) );
  AND2_X1 U4366 ( .A1(n3549), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3548)
         );
  INV_X1 U4367 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5908) );
  AND2_X1 U4368 ( .A1(n3548), .A2(n5908), .ZN(n3544) );
  XNOR2_X1 U4369 ( .A(n3542), .B(n3541), .ZN(n3543) );
  NOR2_X1 U4370 ( .A1(n3544), .A2(n3543), .ZN(n3568) );
  NOR2_X1 U4371 ( .A1(n3568), .A2(n3545), .ZN(n3546) );
  INV_X1 U4372 ( .A(n3548), .ZN(n3551) );
  OAI21_X1 U4373 ( .B1(n3549), .B2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n5908), 
        .ZN(n3550) );
  NAND2_X1 U4374 ( .A1(n3551), .A2(n3550), .ZN(n3573) );
  NOR2_X1 U4375 ( .A1(n3552), .A2(n3573), .ZN(n3553) );
  AOI21_X1 U4376 ( .B1(n6536), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n3553), 
        .ZN(n3554) );
  OAI21_X1 U4377 ( .B1(n3568), .B2(n3558), .A(n3554), .ZN(n3555) );
  INV_X1 U4378 ( .A(n3555), .ZN(n3556) );
  INV_X1 U4379 ( .A(n3558), .ZN(n3560) );
  INV_X1 U4380 ( .A(n3573), .ZN(n3559) );
  NAND2_X1 U4381 ( .A1(n3560), .A2(n3559), .ZN(n3561) );
  INV_X1 U4382 ( .A(n5404), .ZN(n3567) );
  OR2_X1 U4383 ( .A1(n3564), .A2(STATE_REG_0__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U4384 ( .A1(n3187), .A2(n4710), .ZN(n4703) );
  NAND2_X1 U4385 ( .A1(n4703), .A2(n6638), .ZN(n3565) );
  OAI211_X1 U4386 ( .C1(n4313), .C2(n3565), .A(n3602), .B(n5258), .ZN(n3566)
         );
  NAND2_X1 U4387 ( .A1(n3567), .A2(n3566), .ZN(n3576) );
  NAND2_X1 U4388 ( .A1(n4492), .A2(n4710), .ZN(n3574) );
  NAND2_X1 U4389 ( .A1(n3569), .A2(n3568), .ZN(n3570) );
  OR2_X1 U4390 ( .A1(n3571), .A2(n3570), .ZN(n3572) );
  NAND2_X1 U4391 ( .A1(n3573), .A2(n3572), .ZN(n5399) );
  NOR2_X1 U4392 ( .A1(READY_N), .A2(n5399), .ZN(n4321) );
  NAND2_X1 U4393 ( .A1(n3574), .A2(n4321), .ZN(n3575) );
  MUX2_X1 U4394 ( .A(n3576), .B(n3575), .S(n3189), .Z(n3591) );
  INV_X1 U4395 ( .A(n4499), .ZN(n5387) );
  NOR2_X1 U4396 ( .A1(n5387), .A2(n3175), .ZN(n3578) );
  NAND2_X1 U4397 ( .A1(n3578), .A2(n3577), .ZN(n5817) );
  NOR2_X1 U4398 ( .A1(n5817), .A2(n3187), .ZN(n3618) );
  NAND2_X1 U4399 ( .A1(n5817), .A2(n3251), .ZN(n3581) );
  NAND2_X1 U4400 ( .A1(n3581), .A2(n3580), .ZN(n3582) );
  NOR2_X1 U4401 ( .A1(n3579), .A2(n3582), .ZN(n3597) );
  OR2_X1 U4402 ( .A1(n3577), .A2(n5387), .ZN(n4391) );
  NAND2_X1 U4403 ( .A1(n3583), .A2(n3175), .ZN(n3585) );
  AOI21_X1 U4404 ( .B1(n3577), .B2(n4492), .A(n3251), .ZN(n3584) );
  OAI21_X1 U4405 ( .B1(n4391), .B2(n3585), .A(n3584), .ZN(n3610) );
  NOR2_X1 U4406 ( .A1(n3587), .A2(n3602), .ZN(n3588) );
  NAND2_X1 U4407 ( .A1(n3586), .A2(n3588), .ZN(n4285) );
  INV_X1 U4408 ( .A(n4285), .ZN(n5400) );
  AOI21_X1 U4409 ( .B1(n3597), .B2(n3610), .A(n5400), .ZN(n4318) );
  AOI21_X1 U4410 ( .B1(n5404), .B2(n3618), .A(n4318), .ZN(n3590) );
  NAND2_X1 U4411 ( .A1(n3589), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6438) );
  AND2_X1 U4412 ( .A1(n3597), .A2(n2995), .ZN(n6417) );
  INV_X1 U4413 ( .A(n6417), .ZN(n5397) );
  OAI22_X1 U4414 ( .A1(n3175), .A2(n3594), .B1(n4313), .B2(n3026), .ZN(n3595)
         );
  INV_X1 U4415 ( .A(n3595), .ZN(n3598) );
  NAND2_X1 U4416 ( .A1(n3597), .A2(n3596), .ZN(n5395) );
  NAND4_X1 U4417 ( .A1(n5397), .A2(n3598), .A3(n5903), .A4(n5395), .ZN(n3599)
         );
  NAND2_X1 U4418 ( .A1(n3634), .A2(n3599), .ZN(n6157) );
  NOR2_X1 U4419 ( .A1(n4285), .A2(n3187), .ZN(n6399) );
  NAND2_X1 U4420 ( .A1(n3634), .A2(n6399), .ZN(n5200) );
  NAND2_X1 U4421 ( .A1(n3251), .A2(n4492), .ZN(n5392) );
  NOR2_X1 U4422 ( .A1(n5392), .A2(n3189), .ZN(n4317) );
  NAND2_X2 U4423 ( .A1(n5371), .A2(n4236), .ZN(n4344) );
  OAI21_X1 U4424 ( .B1(n4317), .B2(n4344), .A(n3376), .ZN(n3609) );
  OAI21_X1 U4425 ( .B1(n5258), .B2(n3604), .A(n3189), .ZN(n3608) );
  NAND2_X1 U4426 ( .A1(n3605), .A2(n5535), .ZN(n3607) );
  AND4_X1 U4427 ( .A1(n3610), .A2(n3609), .A3(n3608), .A4(n3607), .ZN(n3611)
         );
  AND2_X1 U4428 ( .A1(n3612), .A2(n3611), .ZN(n4302) );
  INV_X1 U4429 ( .A(n3208), .ZN(n3613) );
  OR2_X1 U4430 ( .A1(n5817), .A2(n3613), .ZN(n4418) );
  OAI21_X1 U4431 ( .B1(n4300), .B2(n3602), .A(n4418), .ZN(n3614) );
  INV_X1 U4432 ( .A(n3614), .ZN(n3615) );
  OAI211_X1 U4433 ( .C1(n4503), .C2(n3601), .A(n4302), .B(n3615), .ZN(n3616)
         );
  NAND2_X1 U4434 ( .A1(n3634), .A2(n3616), .ZN(n5196) );
  NOR2_X1 U4435 ( .A1(n3404), .A2(n4447), .ZN(n6133) );
  INV_X1 U4436 ( .A(n6133), .ZN(n3617) );
  NAND2_X1 U4437 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6165) );
  NOR2_X1 U4438 ( .A1(n3617), .A2(n6165), .ZN(n6148) );
  NAND3_X1 U4439 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6148), .ZN(n6099) );
  NAND2_X1 U4440 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6118) );
  INV_X1 U4441 ( .A(n6118), .ZN(n6101) );
  NAND3_X1 U4442 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6101), .ZN(n3620) );
  NOR2_X1 U4443 ( .A1(n6099), .A2(n3620), .ZN(n3708) );
  AND2_X1 U4444 ( .A1(n4302), .A2(n3618), .ZN(n4316) );
  NAND2_X1 U4445 ( .A1(n3634), .A2(n4316), .ZN(n6146) );
  NAND2_X1 U4446 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3619) );
  NAND2_X1 U4447 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U4448 ( .A1(n3404), .A2(n6177), .ZN(n6176) );
  NAND3_X1 U4449 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n6176), .ZN(n6145) );
  NOR2_X1 U4450 ( .A1(n3619), .A2(n6145), .ZN(n6096) );
  INV_X1 U4451 ( .A(n6096), .ZN(n6092) );
  NOR2_X1 U4452 ( .A1(n3620), .A2(n6092), .ZN(n3709) );
  OR2_X1 U4453 ( .A1(n5196), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3622)
         );
  OR2_X1 U4454 ( .A1(n3634), .A2(n6185), .ZN(n3621) );
  AND2_X1 U4455 ( .A1(n3622), .A2(n3621), .ZN(n6132) );
  OAI21_X1 U4456 ( .B1(n6146), .B2(n3709), .A(n6132), .ZN(n3623) );
  INV_X1 U4457 ( .A(n3623), .ZN(n3624) );
  OAI21_X1 U4458 ( .B1(n6134), .B2(n3708), .A(n3624), .ZN(n6088) );
  NAND2_X1 U4459 ( .A1(n6134), .A2(n6146), .ZN(n6136) );
  NAND2_X1 U4460 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5895) );
  NOR2_X1 U4461 ( .A1(n3489), .A2(n5895), .ZN(n5199) );
  NAND2_X1 U4462 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5199), .ZN(n3710) );
  AND2_X1 U4463 ( .A1(n6136), .A2(n3710), .ZN(n3625) );
  NOR2_X1 U4464 ( .A1(n6088), .A2(n3625), .ZN(n5894) );
  NOR2_X1 U4465 ( .A1(n5893), .A2(n3498), .ZN(n5880) );
  INV_X1 U4466 ( .A(n5880), .ZN(n3626) );
  NAND2_X1 U4467 ( .A1(n6136), .A2(n3626), .ZN(n3627) );
  NAND2_X1 U4468 ( .A1(n5894), .A2(n3627), .ZN(n5873) );
  NAND2_X1 U4469 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3721) );
  OAI21_X1 U4470 ( .B1(n3721), .B2(n3711), .A(n6136), .ZN(n3628) );
  INV_X1 U4471 ( .A(n3628), .ZN(n3629) );
  INV_X1 U4472 ( .A(n5766), .ZN(n3713) );
  AND2_X1 U4473 ( .A1(n6136), .A2(n3713), .ZN(n3630) );
  NOR2_X1 U4474 ( .A1(n5774), .A2(n3630), .ZN(n4254) );
  NAND2_X1 U4475 ( .A1(n3193), .A2(n3175), .ZN(n3632) );
  OR2_X1 U4476 ( .A1(n4313), .A2(n3631), .ZN(n6424) );
  OAI21_X1 U4477 ( .B1(n3601), .B2(n3632), .A(n6424), .ZN(n3633) );
  NAND2_X1 U4478 ( .A1(n3634), .A2(n3633), .ZN(n6160) );
  INV_X1 U4479 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4995) );
  NAND2_X1 U4480 ( .A1(n4234), .A2(n4995), .ZN(n3637) );
  NAND3_X1 U4481 ( .A1(n5371), .A2(n3641), .A3(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n3636) );
  NAND2_X1 U4482 ( .A1(n3024), .A2(n3641), .ZN(n3675) );
  NAND2_X1 U4483 ( .A1(n3025), .A2(EBX_REG_1__SCAN_IN), .ZN(n3635) );
  OR2_X1 U4484 ( .A1(n3025), .A2(n4725), .ZN(n3640) );
  INV_X1 U4485 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4725) );
  NAND2_X1 U4486 ( .A1(n5371), .A2(n4725), .ZN(n3639) );
  INV_X1 U4487 ( .A(n3642), .ZN(n3643) );
  NAND2_X1 U4488 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n3026), .ZN(n3644)
         );
  OAI21_X1 U4489 ( .B1(n4271), .B2(EBX_REG_2__SCAN_IN), .A(n3644), .ZN(n3647)
         );
  NAND2_X1 U4490 ( .A1(n3638), .A2(EBX_REG_2__SCAN_IN), .ZN(n3645) );
  NAND2_X1 U4491 ( .A1(n3675), .A2(n3645), .ZN(n3646) );
  MUX2_X1 U4492 ( .A(n4232), .B(n5371), .S(EBX_REG_3__SCAN_IN), .Z(n3648) );
  OAI21_X1 U4493 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n4344), .A(n3648), 
        .ZN(n4463) );
  INV_X1 U4494 ( .A(EBX_REG_4__SCAN_IN), .ZN(n3649) );
  NAND2_X1 U4495 ( .A1(n3022), .A2(n3649), .ZN(n3650) );
  OAI211_X1 U4496 ( .C1(n3638), .C2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n5371), 
        .B(n3650), .ZN(n3651) );
  OAI21_X1 U4497 ( .B1(EBX_REG_4__SCAN_IN), .B2(n4271), .A(n3651), .ZN(n4583)
         );
  NAND2_X1 U4498 ( .A1(n3014), .A2(n3012), .ZN(n4582) );
  MUX2_X1 U4499 ( .A(n4232), .B(n5371), .S(EBX_REG_5__SCAN_IN), .Z(n3652) );
  OAI21_X1 U4500 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4344), .A(n3652), 
        .ZN(n4590) );
  NOR2_X2 U4501 ( .A1(n4582), .A2(n4590), .ZN(n4589) );
  NAND2_X1 U4502 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n3026), .ZN(n3653)
         );
  OAI21_X1 U4503 ( .B1(n4271), .B2(EBX_REG_6__SCAN_IN), .A(n3653), .ZN(n3656)
         );
  NAND2_X1 U4504 ( .A1(n3638), .A2(EBX_REG_6__SCAN_IN), .ZN(n3654) );
  NAND2_X1 U4505 ( .A1(n3675), .A2(n3654), .ZN(n3655) );
  NAND2_X1 U4506 ( .A1(n4589), .A2(n4651), .ZN(n4650) );
  MUX2_X1 U4507 ( .A(n4232), .B(n5371), .S(EBX_REG_7__SCAN_IN), .Z(n3657) );
  OAI21_X1 U4508 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n4344), .A(n3657), 
        .ZN(n4839) );
  NOR2_X1 U4509 ( .A1(n4650), .A2(n4839), .ZN(n4838) );
  INV_X1 U4510 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4975) );
  NAND2_X1 U4511 ( .A1(n3022), .A2(n4975), .ZN(n3658) );
  OAI211_X1 U4512 ( .C1(n3638), .C2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n5371), 
        .B(n3658), .ZN(n3659) );
  OAI21_X1 U4513 ( .B1(EBX_REG_8__SCAN_IN), .B2(n4271), .A(n3659), .ZN(n4974)
         );
  MUX2_X1 U4514 ( .A(n4232), .B(n5371), .S(EBX_REG_9__SCAN_IN), .Z(n3660) );
  OAI21_X1 U4515 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n4344), .A(n3660), 
        .ZN(n5026) );
  INV_X1 U4516 ( .A(n3675), .ZN(n3661) );
  AOI21_X1 U4517 ( .B1(n3638), .B2(EBX_REG_10__SCAN_IN), .A(n3661), .ZN(n3663)
         );
  NAND2_X1 U4518 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n3026), .ZN(n3662) );
  OAI211_X1 U4519 ( .C1(EBX_REG_10__SCAN_IN), .C2(n4271), .A(n3663), .B(n3662), 
        .ZN(n5013) );
  NAND2_X1 U4520 ( .A1(n5024), .A2(n5013), .ZN(n5950) );
  INV_X1 U4521 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U4522 ( .A1(n3684), .A2(n6008), .ZN(n3666) );
  NAND2_X1 U4523 ( .A1(n3022), .A2(n6008), .ZN(n3664) );
  OAI211_X1 U4524 ( .C1(n5535), .C2(n3485), .A(n4236), .B(n3664), .ZN(n3665)
         );
  NAND2_X1 U4525 ( .A1(n3666), .A2(n3665), .ZN(n5951) );
  NOR2_X2 U4526 ( .A1(n5950), .A2(n5951), .ZN(n5078) );
  INV_X1 U4527 ( .A(EBX_REG_12__SCAN_IN), .ZN(n3667) );
  NAND2_X1 U4528 ( .A1(n4234), .A2(n3667), .ZN(n3670) );
  NAND2_X1 U4529 ( .A1(n3638), .A2(EBX_REG_12__SCAN_IN), .ZN(n3669) );
  NAND2_X1 U4530 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n3026), .ZN(n3668) );
  NAND4_X1 U4531 ( .A1(n3670), .A2(n3675), .A3(n3669), .A4(n3668), .ZN(n5079)
         );
  NAND2_X1 U4532 ( .A1(n5078), .A2(n5079), .ZN(n5080) );
  INV_X1 U4533 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U4534 ( .A1(n3022), .A2(n5948), .ZN(n3671) );
  OAI211_X1 U4535 ( .C1(n5535), .C2(n3489), .A(n4236), .B(n3671), .ZN(n3672)
         );
  OAI21_X1 U4536 ( .B1(n4232), .B2(EBX_REG_13__SCAN_IN), .A(n3672), .ZN(n5130)
         );
  NAND2_X1 U4537 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n3026), .ZN(n3673) );
  OAI21_X1 U4538 ( .B1(n4271), .B2(EBX_REG_14__SCAN_IN), .A(n3673), .ZN(n3677)
         );
  NAND2_X1 U4539 ( .A1(n3638), .A2(EBX_REG_14__SCAN_IN), .ZN(n3674) );
  NAND2_X1 U4540 ( .A1(n3675), .A2(n3674), .ZN(n3676) );
  OR2_X1 U4541 ( .A1(n3677), .A2(n3676), .ZN(n5189) );
  INV_X1 U4542 ( .A(EBX_REG_15__SCAN_IN), .ZN(n3678) );
  NAND2_X1 U4543 ( .A1(n3684), .A2(n3678), .ZN(n3681) );
  NAND2_X1 U4544 ( .A1(n3022), .A2(n3678), .ZN(n3679) );
  OAI211_X1 U4545 ( .C1(n5535), .C2(n5893), .A(n4236), .B(n3679), .ZN(n3680)
         );
  NAND2_X1 U4546 ( .A1(n3681), .A2(n3680), .ZN(n5497) );
  NAND2_X1 U4547 ( .A1(n3026), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3683) );
  NAND2_X1 U4548 ( .A1(n3638), .A2(EBX_REG_16__SCAN_IN), .ZN(n3682) );
  OAI211_X1 U4549 ( .C1(n4271), .C2(EBX_REG_16__SCAN_IN), .A(n3683), .B(n3682), 
        .ZN(n5214) );
  INV_X1 U4550 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U4551 ( .A1(n3684), .A2(n5243), .ZN(n3687) );
  NAND2_X1 U4552 ( .A1(n3022), .A2(n5243), .ZN(n3685) );
  OAI211_X1 U4553 ( .C1(n5535), .C2(n5796), .A(n3685), .B(n4236), .ZN(n3686)
         );
  AND2_X1 U4554 ( .A1(n3687), .A2(n3686), .ZN(n5241) );
  INV_X1 U4555 ( .A(EBX_REG_19__SCAN_IN), .ZN(n3688) );
  NAND2_X1 U4556 ( .A1(n4234), .A2(n3688), .ZN(n3692) );
  NAND2_X1 U4557 ( .A1(n4236), .A2(n5788), .ZN(n3690) );
  NAND2_X1 U4558 ( .A1(n3022), .A2(n3688), .ZN(n3689) );
  NAND3_X1 U4559 ( .A1(n3690), .A2(n5371), .A3(n3689), .ZN(n3691) );
  AND2_X1 U4560 ( .A1(n3692), .A2(n3691), .ZN(n5539) );
  OR2_X1 U4561 ( .A1(n4344), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3693)
         );
  INV_X1 U4562 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U4563 ( .A1(n3022), .A2(n5550), .ZN(n5534) );
  AND2_X1 U4564 ( .A1(n3693), .A2(n5534), .ZN(n5537) );
  OAI22_X1 U4565 ( .A1(n4344), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n3026), .ZN(n5487) );
  NAND2_X1 U4566 ( .A1(n5537), .A2(n5487), .ZN(n3695) );
  NAND2_X1 U4567 ( .A1(n5535), .A2(EBX_REG_20__SCAN_IN), .ZN(n3694) );
  OAI211_X1 U4568 ( .C1(n5537), .C2(n5535), .A(n3695), .B(n3694), .ZN(n3696)
         );
  MUX2_X1 U4569 ( .A(n4232), .B(n5371), .S(EBX_REG_21__SCAN_IN), .Z(n3698) );
  INV_X1 U4570 ( .A(n4344), .ZN(n4242) );
  NAND2_X1 U4571 ( .A1(n4242), .A2(n3018), .ZN(n3697) );
  AND2_X1 U4572 ( .A1(n3698), .A2(n3697), .ZN(n5525) );
  NAND2_X1 U4573 ( .A1(n3026), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3700) );
  NAND2_X1 U4574 ( .A1(n3638), .A2(EBX_REG_22__SCAN_IN), .ZN(n3699) );
  OAI211_X1 U4575 ( .C1(n4271), .C2(EBX_REG_22__SCAN_IN), .A(n3700), .B(n3699), 
        .ZN(n5520) );
  INV_X1 U4576 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U4577 ( .A1(n3022), .A2(n5467), .ZN(n3701) );
  OAI211_X1 U4578 ( .C1(n5535), .C2(n3503), .A(n3701), .B(n4236), .ZN(n3702)
         );
  OAI21_X1 U4579 ( .B1(n4232), .B2(EBX_REG_23__SCAN_IN), .A(n3702), .ZN(n3704)
         );
  AND2_X1 U4580 ( .A1(n3703), .A2(n3704), .ZN(n3705) );
  OR2_X1 U4581 ( .A1(n4224), .A2(n3705), .ZN(n5468) );
  INV_X1 U4582 ( .A(n5468), .ZN(n5513) );
  INV_X1 U4583 ( .A(REIP_REG_23__SCAN_IN), .ZN(n3706) );
  NOR2_X1 U4584 ( .A1(n6159), .A2(n3706), .ZN(n5304) );
  AOI21_X1 U4585 ( .B1(n6180), .B2(n5513), .A(n5304), .ZN(n3707) );
  OAI21_X1 U4586 ( .B1(n4254), .B2(n3503), .A(n3707), .ZN(n3715) );
  INV_X1 U4587 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4309) );
  AND2_X1 U4588 ( .A1(n5200), .A2(n4309), .ZN(n4446) );
  NAND2_X1 U4589 ( .A1(n3708), .A2(n6186), .ZN(n5116) );
  INV_X1 U4590 ( .A(n6146), .ZN(n6179) );
  NAND2_X1 U4591 ( .A1(n6179), .A2(n3709), .ZN(n5195) );
  NAND2_X1 U4592 ( .A1(n5116), .A2(n5195), .ZN(n6087) );
  NOR2_X1 U4593 ( .A1(n3710), .A2(n5901), .ZN(n5879) );
  NAND2_X1 U4594 ( .A1(n5880), .A2(n5879), .ZN(n5878) );
  INV_X1 U4595 ( .A(n3721), .ZN(n3712) );
  NAND2_X1 U4596 ( .A1(n5789), .A2(n3712), .ZN(n5777) );
  NOR2_X1 U4597 ( .A1(n5756), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3714)
         );
  NOR2_X1 U4598 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5765) );
  NOR2_X1 U4599 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3719) );
  NAND4_X1 U4600 ( .A1(n5765), .A2(n3719), .A3(n5788), .A4(n3718), .ZN(n3720)
         );
  OAI21_X1 U4601 ( .B1(n5653), .B2(n3720), .A(n5672), .ZN(n3725) );
  NAND2_X1 U4602 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4258) );
  NOR2_X1 U4603 ( .A1(n4258), .A2(n3721), .ZN(n3722) );
  NAND2_X1 U4604 ( .A1(n5653), .A2(n3723), .ZN(n3724) );
  NAND2_X1 U4605 ( .A1(n3725), .A2(n3724), .ZN(n5585) );
  XOR2_X1 U4606 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(n3477), .Z(n5612) );
  INV_X1 U4607 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U4608 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4259) );
  INV_X1 U4609 ( .A(n5605), .ZN(n3729) );
  NOR2_X1 U4610 ( .A1(n3477), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5586)
         );
  NOR2_X1 U4611 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5725) );
  AND2_X1 U4612 ( .A1(n5586), .A2(n5725), .ZN(n3728) );
  NAND2_X1 U4613 ( .A1(n3729), .A2(n3728), .ZN(n3731) );
  INV_X1 U4614 ( .A(n3731), .ZN(n3730) );
  OAI21_X1 U4615 ( .B1(n4263), .B2(n3730), .A(INSTADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n3732) );
  INV_X1 U4616 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5714) );
  AOI22_X1 U4617 ( .A1(n3732), .A2(n4220), .B1(n4263), .B2(n5714), .ZN(n5717)
         );
  NAND2_X2 U4618 ( .A1(n4740), .A2(n6417), .ZN(n6060) );
  AOI22_X1 U4619 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n2985), .B1(n5275), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4620 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4194), .B1(n4187), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4621 ( .A1(n4121), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4622 ( .A1(n2986), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3733) );
  NAND4_X1 U4623 ( .A1(n3736), .A2(n3735), .A3(n3734), .A4(n3733), .ZN(n3742)
         );
  AOI22_X1 U4624 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n2984), .B1(n5274), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4625 ( .A1(n3239), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4626 ( .A1(n4189), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4627 ( .A1(n5268), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3737) );
  NAND4_X1 U4628 ( .A1(n3740), .A2(n3739), .A3(n3738), .A4(n3737), .ZN(n3741)
         );
  NOR2_X1 U4629 ( .A1(n3742), .A2(n3741), .ZN(n3745) );
  INV_X2 U4630 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6534) );
  NOR2_X2 U4631 ( .A1(n4503), .A2(n6534), .ZN(n3930) );
  INV_X1 U4632 ( .A(n3930), .ZN(n3817) );
  INV_X1 U4633 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5963) );
  INV_X1 U4634 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3852) );
  XNOR2_X1 U4635 ( .A(n3868), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5112)
         );
  INV_X1 U4636 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6604) );
  NAND2_X1 U4637 ( .A1(n6534), .A2(n6604), .ZN(n5294) );
  INV_X2 U4638 ( .A(n5294), .ZN(n5288) );
  NAND2_X1 U4639 ( .A1(n5112), .A2(n5288), .ZN(n3744) );
  NAND2_X1 U4640 ( .A1(n6534), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3871) );
  INV_X1 U4641 ( .A(n3871), .ZN(n5317) );
  AOI22_X1 U4642 ( .A1(n4204), .A2(EAX_REG_12__SCAN_IN), .B1(n5317), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3743) );
  OAI211_X1 U4643 ( .C1(n3745), .C2(n3817), .A(n3744), .B(n3743), .ZN(n5076)
         );
  NAND2_X1 U4644 ( .A1(n4471), .A2(n3930), .ZN(n3750) );
  NAND2_X1 U4645 ( .A1(n3193), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3778) );
  NAND2_X1 U4646 ( .A1(n4204), .A2(EAX_REG_1__SCAN_IN), .ZN(n3747) );
  NAND2_X1 U4647 ( .A1(n6534), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3746)
         );
  OAI211_X1 U4648 ( .C1(n3778), .C2(n3181), .A(n3747), .B(n3746), .ZN(n3748)
         );
  INV_X1 U4649 ( .A(n3748), .ZN(n3749) );
  NAND2_X1 U4650 ( .A1(n3750), .A2(n3749), .ZN(n4397) );
  NAND2_X1 U4651 ( .A1(n5046), .A2(n3113), .ZN(n3752) );
  NAND2_X1 U4652 ( .A1(n3752), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4351) );
  NAND2_X1 U4654 ( .A1(n4204), .A2(EAX_REG_0__SCAN_IN), .ZN(n3755) );
  NAND2_X1 U4655 ( .A1(n6534), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3754)
         );
  OAI211_X1 U4656 ( .C1(n3778), .C2(n3205), .A(n3755), .B(n3754), .ZN(n3756)
         );
  AOI21_X1 U4657 ( .B1(n6330), .B2(n3930), .A(n3756), .ZN(n3757) );
  INV_X1 U4658 ( .A(n3757), .ZN(n4353) );
  OR2_X1 U4659 ( .A1(n4353), .A2(n5294), .ZN(n3758) );
  NAND2_X1 U4660 ( .A1(n4352), .A2(n3758), .ZN(n4400) );
  AND2_X2 U4661 ( .A1(n4397), .A2(n4400), .ZN(n3764) );
  NAND2_X1 U4662 ( .A1(n4470), .A2(n3930), .ZN(n3759) );
  NAND2_X1 U4663 ( .A1(n3759), .A2(n3871), .ZN(n3763) );
  OAI21_X1 U4664 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3760), .ZN(n6084) );
  AOI22_X1 U4665 ( .A1(n5317), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n5288), 
        .B2(n6084), .ZN(n3762) );
  NAND2_X1 U4666 ( .A1(n4204), .A2(EAX_REG_2__SCAN_IN), .ZN(n3761) );
  OAI211_X1 U4667 ( .C1(n3778), .C2(n3291), .A(n3762), .B(n3761), .ZN(n4455)
         );
  NAND2_X1 U4668 ( .A1(n4454), .A2(n4455), .ZN(n3766) );
  NAND2_X1 U4669 ( .A1(n3763), .A2(n4398), .ZN(n3765) );
  NAND2_X1 U4670 ( .A1(n3766), .A2(n3765), .ZN(n4452) );
  NAND2_X1 U4671 ( .A1(n3767), .A2(n3930), .ZN(n3774) );
  OAI21_X1 U4672 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3769), .A(n3768), 
        .ZN(n6075) );
  AOI22_X1 U4673 ( .A1(n5288), .A2(n6075), .B1(n5317), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3771) );
  NAND2_X1 U4674 ( .A1(n4204), .A2(EAX_REG_3__SCAN_IN), .ZN(n3770) );
  OAI211_X1 U4675 ( .C1(n3778), .C2(n3319), .A(n3771), .B(n3770), .ZN(n3772)
         );
  INV_X1 U4676 ( .A(n3772), .ZN(n3773) );
  NAND2_X1 U4677 ( .A1(n3774), .A2(n3773), .ZN(n4460) );
  INV_X1 U4678 ( .A(n4580), .ZN(n3785) );
  NAND2_X1 U4679 ( .A1(n4204), .A2(EAX_REG_4__SCAN_IN), .ZN(n3777) );
  OAI21_X1 U4680 ( .B1(n6604), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6534), 
        .ZN(n3776) );
  OAI211_X1 U4681 ( .C1(n3778), .C2(n5908), .A(n3777), .B(n3776), .ZN(n3782)
         );
  NOR2_X1 U4682 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3779), .ZN(n3780)
         );
  NOR2_X1 U4683 ( .A1(n3787), .A2(n3780), .ZN(n4968) );
  NAND2_X1 U4684 ( .A1(n4968), .A2(n5288), .ZN(n3781) );
  AND2_X1 U4685 ( .A1(n3782), .A2(n3781), .ZN(n3783) );
  AOI21_X1 U4686 ( .B1(n3775), .B2(n3930), .A(n3783), .ZN(n4581) );
  NAND2_X1 U4687 ( .A1(n3785), .A2(n3784), .ZN(n4578) );
  INV_X1 U4688 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3789) );
  XNOR2_X1 U4689 ( .A(n3787), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4937) );
  AOI22_X1 U4690 ( .A1(n4937), .A2(n5288), .B1(n5317), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3788) );
  OAI21_X1 U4691 ( .B1(n3032), .B2(n3789), .A(n3788), .ZN(n3790) );
  NAND2_X1 U4692 ( .A1(n3791), .A2(n3930), .ZN(n3797) );
  AND2_X1 U4693 ( .A1(n3792), .A2(n5978), .ZN(n3793) );
  OR2_X1 U4694 ( .A1(n3793), .A2(n3798), .ZN(n6068) );
  NAND2_X1 U4695 ( .A1(n6068), .A2(n5288), .ZN(n3794) );
  OAI21_X1 U4696 ( .B1(n5978), .B2(n3871), .A(n3794), .ZN(n3795) );
  AOI21_X1 U4697 ( .B1(n4204), .B2(EAX_REG_6__SCAN_IN), .A(n3795), .ZN(n3796)
         );
  NAND2_X1 U4698 ( .A1(n4586), .A2(n4648), .ZN(n4647) );
  INV_X1 U4699 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3801) );
  XNOR2_X1 U4700 ( .A(n3798), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4945) );
  INV_X1 U4701 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4844) );
  NOR2_X1 U4702 ( .A1(n3871), .A2(n4844), .ZN(n3799) );
  AOI21_X1 U4703 ( .B1(n4945), .B2(n5288), .A(n3799), .ZN(n3800) );
  OAI21_X1 U4704 ( .B1(n3032), .B2(n3801), .A(n3800), .ZN(n3802) );
  OR2_X2 U4705 ( .A1(n4647), .A2(n4837), .ZN(n4971) );
  AOI22_X1 U4706 ( .A1(n4189), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n2986), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4707 ( .A1(n4194), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4708 ( .A1(n2984), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4709 ( .A1(n5277), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3804) );
  NAND4_X1 U4710 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3813)
         );
  AOI22_X1 U4711 ( .A1(n5275), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4712 ( .A1(n4121), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4713 ( .A1(n4188), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4714 ( .A1(n2985), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3808) );
  NAND4_X1 U4715 ( .A1(n3811), .A2(n3810), .A3(n3809), .A4(n3808), .ZN(n3812)
         );
  NOR2_X1 U4716 ( .A1(n3813), .A2(n3812), .ZN(n3818) );
  XNOR2_X1 U4717 ( .A(n3814), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5070)
         );
  NAND2_X1 U4718 ( .A1(n5070), .A2(n5288), .ZN(n3816) );
  AOI22_X1 U4719 ( .A1(n4204), .A2(EAX_REG_10__SCAN_IN), .B1(n5317), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3815) );
  OAI211_X1 U4720 ( .C1(n3818), .C2(n3817), .A(n3816), .B(n3815), .ZN(n5009)
         );
  INV_X1 U4721 ( .A(n5009), .ZN(n3850) );
  XOR2_X1 U4722 ( .A(n5963), .B(n3819), .Z(n5967) );
  INV_X1 U4723 ( .A(n5967), .ZN(n3834) );
  AOI22_X1 U4724 ( .A1(n2985), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5277), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4725 ( .A1(n4194), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4726 ( .A1(n4189), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4727 ( .A1(n5276), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3820) );
  NAND4_X1 U4728 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3829)
         );
  AOI22_X1 U4729 ( .A1(n2984), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4730 ( .A1(n5275), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4731 ( .A1(n2986), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4732 ( .A1(n4121), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3824) );
  NAND4_X1 U4733 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3828)
         );
  OAI21_X1 U4734 ( .B1(n3829), .B2(n3828), .A(n3930), .ZN(n3832) );
  NAND2_X1 U4735 ( .A1(n4204), .A2(EAX_REG_9__SCAN_IN), .ZN(n3831) );
  NAND2_X1 U4736 ( .A1(n5317), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3830)
         );
  NAND3_X1 U4737 ( .A1(n3832), .A2(n3831), .A3(n3830), .ZN(n3833) );
  AOI21_X1 U4738 ( .B1(n3834), .B2(n5288), .A(n3833), .ZN(n5020) );
  AOI22_X1 U4739 ( .A1(n5274), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n5275), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4740 ( .A1(n4121), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4741 ( .A1(n2986), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4742 ( .A1(n5265), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3835) );
  NAND4_X1 U4743 ( .A1(n3838), .A2(n3837), .A3(n3836), .A4(n3835), .ZN(n3844)
         );
  AOI22_X1 U4744 ( .A1(n2984), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4745 ( .A1(n3239), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4746 ( .A1(n4189), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4747 ( .A1(n2985), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3839) );
  NAND4_X1 U4748 ( .A1(n3842), .A2(n3841), .A3(n3840), .A4(n3839), .ZN(n3843)
         );
  OAI21_X1 U4749 ( .B1(n3844), .B2(n3843), .A(n3930), .ZN(n3849) );
  NAND2_X1 U4750 ( .A1(n4204), .A2(EAX_REG_8__SCAN_IN), .ZN(n3848) );
  XNOR2_X1 U4751 ( .A(n3845), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4988) );
  NAND2_X1 U4752 ( .A1(n4988), .A2(n5288), .ZN(n3847) );
  NAND2_X1 U4753 ( .A1(n5317), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3846)
         );
  AND4_X1 U4754 ( .A1(n3849), .A2(n3848), .A3(n3847), .A4(n3846), .ZN(n4973)
         );
  OR2_X1 U4755 ( .A1(n5020), .A2(n4973), .ZN(n5007) );
  XOR2_X1 U4756 ( .A(n3852), .B(n3851), .Z(n6055) );
  AOI22_X1 U4757 ( .A1(n5275), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4758 ( .A1(n2984), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4759 ( .A1(n3239), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4760 ( .A1(n5276), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3853) );
  NAND4_X1 U4761 ( .A1(n3856), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(n3862)
         );
  AOI22_X1 U4762 ( .A1(n2985), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4121), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4763 ( .A1(n4189), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4764 ( .A1(n5274), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4765 ( .A1(n2986), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3857) );
  NAND4_X1 U4766 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3861)
         );
  OR2_X1 U4767 ( .A1(n3862), .A2(n3861), .ZN(n3863) );
  AOI22_X1 U4768 ( .A1(n3930), .A2(n3863), .B1(n5317), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3865) );
  NAND2_X1 U4769 ( .A1(n4204), .A2(EAX_REG_11__SCAN_IN), .ZN(n3864) );
  OAI211_X1 U4770 ( .C1(n6055), .C2(n5294), .A(n3865), .B(n3864), .ZN(n5005)
         );
  INV_X1 U4771 ( .A(n5005), .ZN(n3866) );
  NOR2_X2 U4772 ( .A1(n4971), .A2(n3867), .ZN(n5075) );
  AND2_X2 U4773 ( .A1(n5075), .A2(n5076), .ZN(n3875) );
  INV_X1 U4774 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3872) );
  OAI21_X1 U4775 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3869), .A(n3892), 
        .ZN(n5939) );
  NAND2_X1 U4776 ( .A1(n5939), .A2(n5288), .ZN(n3870) );
  OAI21_X1 U4777 ( .B1(n3872), .B2(n3871), .A(n3870), .ZN(n3873) );
  AOI21_X1 U4778 ( .B1(n4204), .B2(EAX_REG_13__SCAN_IN), .A(n3873), .ZN(n3877)
         );
  INV_X1 U4779 ( .A(n3877), .ZN(n3874) );
  NAND2_X2 U4780 ( .A1(n3875), .A2(n3874), .ZN(n3891) );
  NAND2_X1 U4781 ( .A1(n3876), .A2(n5075), .ZN(n3879) );
  NAND2_X1 U4782 ( .A1(n3879), .A2(n3878), .ZN(n5128) );
  AOI22_X1 U4783 ( .A1(n4121), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4784 ( .A1(n2984), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4785 ( .A1(n5277), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4786 ( .A1(n2985), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3880) );
  NAND4_X1 U4787 ( .A1(n3883), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3889)
         );
  AOI22_X1 U4788 ( .A1(n5274), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4789 ( .A1(n4189), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4790 ( .A1(n5275), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4791 ( .A1(n2986), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3884) );
  NAND4_X1 U4792 ( .A1(n3887), .A2(n3886), .A3(n3885), .A4(n3884), .ZN(n3888)
         );
  OR2_X1 U4793 ( .A1(n3889), .A2(n3888), .ZN(n3890) );
  AND2_X1 U4794 ( .A1(n3930), .A2(n3890), .ZN(n5127) );
  NAND2_X1 U4795 ( .A1(n5126), .A2(n3891), .ZN(n5188) );
  XOR2_X1 U4796 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3906), .Z(n5251) );
  AOI22_X1 U4797 ( .A1(n4121), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4798 ( .A1(n5275), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4799 ( .A1(n3239), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4800 ( .A1(n5268), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3893) );
  NAND4_X1 U4801 ( .A1(n3896), .A2(n3895), .A3(n3894), .A4(n3893), .ZN(n3902)
         );
  AOI22_X1 U4802 ( .A1(n2985), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4803 ( .A1(n4194), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4804 ( .A1(n4189), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4805 ( .A1(n2986), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3897) );
  NAND4_X1 U4806 ( .A1(n3900), .A2(n3899), .A3(n3898), .A4(n3897), .ZN(n3901)
         );
  OR2_X1 U4807 ( .A1(n3902), .A2(n3901), .ZN(n3903) );
  AOI22_X1 U4808 ( .A1(n3930), .A2(n3903), .B1(n5317), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3905) );
  NAND2_X1 U4809 ( .A1(n4204), .A2(EAX_REG_14__SCAN_IN), .ZN(n3904) );
  OAI211_X1 U4810 ( .C1(n5251), .C2(n5294), .A(n3905), .B(n3904), .ZN(n5187)
         );
  NAND2_X1 U4811 ( .A1(n5188), .A2(n5187), .ZN(n5186) );
  INV_X1 U4812 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3920) );
  XOR2_X1 U4813 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3938), .Z(n5218) );
  INV_X1 U4814 ( .A(n5218), .ZN(n5695) );
  OR2_X1 U4815 ( .A1(n5817), .A2(n6536), .ZN(n5291) );
  AOI22_X1 U4816 ( .A1(n2984), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4817 ( .A1(n4121), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n2986), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4818 ( .A1(n4189), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4819 ( .A1(n2985), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3907) );
  NAND4_X1 U4820 ( .A1(n3910), .A2(n3909), .A3(n3908), .A4(n3907), .ZN(n3916)
         );
  AOI22_X1 U4821 ( .A1(n4194), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4822 ( .A1(n5275), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4823 ( .A1(n5276), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4824 ( .A1(n3239), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3911) );
  NAND4_X1 U4825 ( .A1(n3914), .A2(n3913), .A3(n3912), .A4(n3911), .ZN(n3915)
         );
  NOR2_X1 U4826 ( .A1(n3916), .A2(n3915), .ZN(n3918) );
  AOI22_X1 U4827 ( .A1(n4204), .A2(EAX_REG_16__SCAN_IN), .B1(n5317), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3917) );
  OAI21_X1 U4828 ( .B1(n5291), .B2(n3918), .A(n3917), .ZN(n3919) );
  AOI21_X1 U4829 ( .B1(n5695), .B2(n5288), .A(n3919), .ZN(n5206) );
  XNOR2_X1 U4830 ( .A(n3921), .B(n3920), .ZN(n5703) );
  AOI22_X1 U4831 ( .A1(n4194), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4832 ( .A1(n2985), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4833 ( .A1(n2986), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4834 ( .A1(n5276), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3922) );
  NAND4_X1 U4835 ( .A1(n3925), .A2(n3924), .A3(n3923), .A4(n3922), .ZN(n3932)
         );
  AOI22_X1 U4836 ( .A1(n2984), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n5275), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4837 ( .A1(n5277), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4838 ( .A1(n4189), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4839 ( .A1(n4121), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3926) );
  NAND4_X1 U4840 ( .A1(n3929), .A2(n3928), .A3(n3927), .A4(n3926), .ZN(n3931)
         );
  OAI21_X1 U4841 ( .B1(n3932), .B2(n3931), .A(n3930), .ZN(n3935) );
  NAND2_X1 U4842 ( .A1(n4204), .A2(EAX_REG_15__SCAN_IN), .ZN(n3934) );
  NAND2_X1 U4843 ( .A1(n5317), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3933)
         );
  NAND3_X1 U4844 ( .A1(n3935), .A2(n3934), .A3(n3933), .ZN(n3936) );
  AOI21_X1 U4845 ( .B1(n5703), .B2(n5288), .A(n3936), .ZN(n5495) );
  OR2_X1 U4846 ( .A1(n5206), .A2(n5495), .ZN(n3937) );
  NOR2_X2 U4847 ( .A1(n5186), .A2(n3937), .ZN(n5207) );
  NAND2_X1 U4848 ( .A1(n3938), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3955)
         );
  XNOR2_X1 U4849 ( .A(n3955), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5683)
         );
  NAND2_X1 U4850 ( .A1(n5291), .A2(n5294), .ZN(n4022) );
  AOI22_X1 U4851 ( .A1(n2985), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4852 ( .A1(n4189), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4853 ( .A1(n5276), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3942) );
  NAND2_X1 U4854 ( .A1(n5274), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3940) );
  AOI21_X1 U4855 ( .B1(n3244), .B2(INSTQUEUE_REG_2__1__SCAN_IN), .A(n5288), 
        .ZN(n3939) );
  AND2_X1 U4856 ( .A1(n3940), .A2(n3939), .ZN(n3941) );
  NAND4_X1 U4857 ( .A1(n3944), .A2(n3943), .A3(n3942), .A4(n3941), .ZN(n3950)
         );
  AOI22_X1 U4858 ( .A1(n2986), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5275), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4859 ( .A1(n4121), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4860 ( .A1(n4194), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4861 ( .A1(n3239), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3945) );
  NAND4_X1 U4862 ( .A1(n3948), .A2(n3947), .A3(n3946), .A4(n3945), .ZN(n3949)
         );
  OR2_X1 U4863 ( .A1(n3950), .A2(n3949), .ZN(n3953) );
  INV_X1 U4864 ( .A(EAX_REG_17__SCAN_IN), .ZN(n3951) );
  INV_X1 U4865 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5680) );
  OAI22_X1 U4866 ( .A1(n3032), .A2(n3951), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5680), .ZN(n3952) );
  AOI21_X1 U4867 ( .B1(n4022), .B2(n3953), .A(n3952), .ZN(n3954) );
  AOI21_X1 U4868 ( .B1(n5683), .B2(n5288), .A(n3954), .ZN(n5237) );
  NAND2_X1 U4869 ( .A1(n5207), .A2(n5237), .ZN(n5235) );
  NOR2_X1 U4870 ( .A1(n3956), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3957)
         );
  OR2_X1 U4871 ( .A1(n3990), .A2(n3957), .ZN(n5928) );
  AOI22_X1 U4872 ( .A1(n5275), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4873 ( .A1(n2984), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4874 ( .A1(n4189), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4875 ( .A1(n5265), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3958) );
  NAND4_X1 U4876 ( .A1(n3961), .A2(n3960), .A3(n3959), .A4(n3958), .ZN(n3967)
         );
  AOI22_X1 U4877 ( .A1(n3239), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4878 ( .A1(n4121), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n2986), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4879 ( .A1(n4188), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4880 ( .A1(n2985), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3962) );
  NAND4_X1 U4881 ( .A1(n3965), .A2(n3964), .A3(n3963), .A4(n3962), .ZN(n3966)
         );
  NOR2_X1 U4882 ( .A1(n3967), .A2(n3966), .ZN(n3968) );
  NOR2_X1 U4883 ( .A1(n5291), .A2(n3968), .ZN(n3972) );
  INV_X1 U4884 ( .A(EAX_REG_18__SCAN_IN), .ZN(n3970) );
  NAND2_X1 U4885 ( .A1(n6534), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3969)
         );
  OAI211_X1 U4886 ( .C1(n3032), .C2(n3970), .A(n5294), .B(n3969), .ZN(n3971)
         );
  OAI22_X1 U4887 ( .A1(n5928), .A2(n5294), .B1(n3972), .B2(n3971), .ZN(n5542)
         );
  NOR2_X1 U4888 ( .A1(n5235), .A2(n5542), .ZN(n3973) );
  INV_X1 U4889 ( .A(n3973), .ZN(n5531) );
  INV_X1 U4890 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5859) );
  XNOR2_X1 U4891 ( .A(n3990), .B(n5859), .ZN(n5857) );
  NAND2_X1 U4892 ( .A1(n5857), .A2(n5288), .ZN(n3989) );
  AOI22_X1 U4893 ( .A1(n4194), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5275), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4894 ( .A1(n4189), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4895 ( .A1(n2984), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4896 ( .A1(n5266), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3974) );
  NAND4_X1 U4897 ( .A1(n3977), .A2(n3976), .A3(n3975), .A4(n3974), .ZN(n3985)
         );
  AOI22_X1 U4898 ( .A1(n5277), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n2986), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3983) );
  NAND2_X1 U4899 ( .A1(n5273), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3979)
         );
  NAND2_X1 U4900 ( .A1(n4187), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3978) );
  AND3_X1 U4901 ( .A1(n3979), .A2(n3978), .A3(n5294), .ZN(n3982) );
  AOI22_X1 U4902 ( .A1(n2985), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4903 ( .A1(n4188), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3980) );
  NAND4_X1 U4904 ( .A1(n3983), .A2(n3982), .A3(n3981), .A4(n3980), .ZN(n3984)
         );
  OAI21_X1 U4905 ( .B1(n3985), .B2(n3984), .A(n4022), .ZN(n3987) );
  AOI22_X1 U4906 ( .A1(n4204), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6534), .ZN(n3986) );
  NAND2_X1 U4907 ( .A1(n3987), .A2(n3986), .ZN(n3988) );
  NAND2_X1 U4908 ( .A1(n3989), .A2(n3988), .ZN(n5532) );
  OR2_X1 U4909 ( .A1(n3991), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3992)
         );
  NAND2_X1 U4910 ( .A1(n3992), .A2(n4040), .ZN(n5646) );
  INV_X1 U4911 ( .A(n5646), .ZN(n4008) );
  INV_X1 U4912 ( .A(n5291), .ZN(n4201) );
  AOI22_X1 U4913 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4194), .B1(n5274), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4914 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4121), .B1(n2986), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4915 ( .A1(n4189), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4916 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n5275), .B1(n5268), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3993) );
  NAND4_X1 U4917 ( .A1(n3996), .A2(n3995), .A3(n3994), .A4(n3993), .ZN(n4002)
         );
  AOI22_X1 U4918 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n2984), .B1(n4187), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4919 ( .A1(n5277), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4920 ( .A1(n5276), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4921 ( .A1(n2985), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3997) );
  NAND4_X1 U4922 ( .A1(n4000), .A2(n3999), .A3(n3998), .A4(n3997), .ZN(n4001)
         );
  OR2_X1 U4923 ( .A1(n4002), .A2(n4001), .ZN(n4006) );
  INV_X1 U4924 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4004) );
  NAND2_X1 U4925 ( .A1(n6534), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4003)
         );
  OAI211_X1 U4926 ( .C1(n3032), .C2(n4004), .A(n5294), .B(n4003), .ZN(n4005)
         );
  AOI21_X1 U4927 ( .B1(n4201), .B2(n4006), .A(n4005), .ZN(n4007) );
  AOI21_X1 U4928 ( .B1(n4008), .B2(n5288), .A(n4007), .ZN(n5479) );
  AOI22_X1 U4929 ( .A1(n3239), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4014) );
  NAND2_X1 U4930 ( .A1(n5274), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4010) );
  NAND2_X1 U4931 ( .A1(n4189), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4009)
         );
  AND3_X1 U4932 ( .A1(n4010), .A2(n4009), .A3(n5294), .ZN(n4013) );
  AOI22_X1 U4933 ( .A1(n5266), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4934 ( .A1(n5275), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4011) );
  NAND4_X1 U4935 ( .A1(n4014), .A2(n4013), .A3(n4012), .A4(n4011), .ZN(n4020)
         );
  AOI22_X1 U4936 ( .A1(n2985), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U4937 ( .A1(n2986), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4938 ( .A1(n4121), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U4939 ( .A1(n5276), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4015) );
  NAND4_X1 U4940 ( .A1(n4018), .A2(n4017), .A3(n4016), .A4(n4015), .ZN(n4019)
         );
  OR2_X1 U4941 ( .A1(n4020), .A2(n4019), .ZN(n4021) );
  NAND2_X1 U4942 ( .A1(n4022), .A2(n4021), .ZN(n4025) );
  AOI22_X1 U4943 ( .A1(n4204), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6534), .ZN(n4024) );
  XNOR2_X1 U4944 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n4040), .ZN(n5847)
         );
  AND2_X1 U4945 ( .A1(n5847), .A2(n5288), .ZN(n4023) );
  AOI21_X1 U4946 ( .B1(n4025), .B2(n4024), .A(n4023), .ZN(n5523) );
  NAND2_X1 U4947 ( .A1(n5476), .A2(n5523), .ZN(n5515) );
  INV_X1 U4948 ( .A(n5515), .ZN(n4048) );
  AOI22_X1 U4949 ( .A1(n5275), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U4950 ( .A1(n4194), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U4951 ( .A1(n5276), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U4952 ( .A1(n4189), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4026) );
  NAND4_X1 U4953 ( .A1(n4029), .A2(n4028), .A3(n4027), .A4(n4026), .ZN(n4035)
         );
  AOI22_X1 U4954 ( .A1(n5277), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U4955 ( .A1(n5273), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U4956 ( .A1(n3129), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U4957 ( .A1(n2986), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4030) );
  NAND4_X1 U4958 ( .A1(n4033), .A2(n4032), .A3(n4031), .A4(n4030), .ZN(n4034)
         );
  NOR2_X1 U4959 ( .A1(n4035), .A2(n4034), .ZN(n4039) );
  NAND2_X1 U4960 ( .A1(n6534), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4036)
         );
  NAND2_X1 U4961 ( .A1(n5294), .A2(n4036), .ZN(n4037) );
  AOI21_X1 U4962 ( .B1(n4204), .B2(EAX_REG_22__SCAN_IN), .A(n4037), .ZN(n4038)
         );
  OAI21_X1 U4963 ( .B1(n5291), .B2(n4039), .A(n4038), .ZN(n4046) );
  INV_X1 U4964 ( .A(n4040), .ZN(n4041) );
  INV_X1 U4965 ( .A(n4042), .ZN(n4043) );
  INV_X1 U4966 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U4967 ( .A1(n4043), .A2(n5840), .ZN(n4044) );
  AND2_X1 U4968 ( .A1(n4089), .A2(n4044), .ZN(n5838) );
  NAND2_X1 U4969 ( .A1(n5838), .A2(n5288), .ZN(n4045) );
  NAND2_X1 U4970 ( .A1(n4046), .A2(n4045), .ZN(n5519) );
  NAND2_X1 U4971 ( .A1(n4048), .A2(n4047), .ZN(n5300) );
  AOI22_X1 U4972 ( .A1(n2986), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U4973 ( .A1(n5274), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U4974 ( .A1(n5275), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4050) );
  AOI22_X1 U4975 ( .A1(n2985), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4049) );
  NAND4_X1 U4976 ( .A1(n4052), .A2(n4051), .A3(n4050), .A4(n4049), .ZN(n4058)
         );
  AOI22_X1 U4977 ( .A1(n4194), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U4978 ( .A1(n4189), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U4979 ( .A1(n3239), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U4980 ( .A1(n4121), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4053) );
  NAND4_X1 U4981 ( .A1(n4056), .A2(n4055), .A3(n4054), .A4(n4053), .ZN(n4057)
         );
  NOR2_X1 U4982 ( .A1(n4058), .A2(n4057), .ZN(n4075) );
  AOI22_X1 U4983 ( .A1(n5277), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U4984 ( .A1(n4189), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U4985 ( .A1(n5276), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U4986 ( .A1(n5273), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4059) );
  NAND4_X1 U4987 ( .A1(n4062), .A2(n4061), .A3(n4060), .A4(n4059), .ZN(n4068)
         );
  AOI22_X1 U4988 ( .A1(n2985), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n2986), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U4989 ( .A1(n4194), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U4990 ( .A1(n5275), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U4991 ( .A1(n5265), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4063) );
  NAND4_X1 U4992 ( .A1(n4066), .A2(n4065), .A3(n4064), .A4(n4063), .ZN(n4067)
         );
  NOR2_X1 U4993 ( .A1(n4068), .A2(n4067), .ZN(n4076) );
  XOR2_X1 U4994 ( .A(n4075), .B(n4076), .Z(n4069) );
  NAND2_X1 U4995 ( .A1(n4069), .A2(n4201), .ZN(n4072) );
  INV_X1 U4996 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5466) );
  OAI21_X1 U4997 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5466), .A(n5294), .ZN(
        n4070) );
  AOI21_X1 U4998 ( .B1(n4204), .B2(EAX_REG_23__SCAN_IN), .A(n4070), .ZN(n4071)
         );
  NAND2_X1 U4999 ( .A1(n4072), .A2(n4071), .ZN(n4074) );
  XNOR2_X1 U5000 ( .A(n4089), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5471)
         );
  NAND2_X1 U5001 ( .A1(n5471), .A2(n5288), .ZN(n4073) );
  NAND2_X1 U5002 ( .A1(n4074), .A2(n4073), .ZN(n5301) );
  INV_X1 U5003 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4096) );
  NOR2_X1 U5004 ( .A1(n4076), .A2(n4075), .ZN(n4108) );
  AOI22_X1 U5005 ( .A1(n2984), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4080) );
  AOI22_X1 U5006 ( .A1(n4194), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4079) );
  AOI22_X1 U5007 ( .A1(n5275), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U5008 ( .A1(n3239), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4077) );
  NAND4_X1 U5009 ( .A1(n4080), .A2(n4079), .A3(n4078), .A4(n4077), .ZN(n4086)
         );
  AOI22_X1 U5010 ( .A1(n4121), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U5011 ( .A1(n4189), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U5012 ( .A1(n2985), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U5013 ( .A1(n2986), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4081) );
  NAND4_X1 U5014 ( .A1(n4084), .A2(n4083), .A3(n4082), .A4(n4081), .ZN(n4085)
         );
  OR2_X1 U5015 ( .A1(n4086), .A2(n4085), .ZN(n4107) );
  INV_X1 U5016 ( .A(n4107), .ZN(n4087) );
  XNOR2_X1 U5017 ( .A(n4108), .B(n4087), .ZN(n4088) );
  NAND2_X1 U5018 ( .A1(n4088), .A2(n4201), .ZN(n4095) );
  NAND2_X1 U5019 ( .A1(n4090), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4143)
         );
  INV_X1 U5020 ( .A(n4090), .ZN(n4092) );
  INV_X1 U5021 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4091) );
  NAND2_X1 U5022 ( .A1(n4092), .A2(n4091), .ZN(n4093) );
  NAND2_X1 U5023 ( .A1(n4143), .A2(n4093), .ZN(n5625) );
  AOI22_X1 U5024 ( .A1(n5625), .A2(n5288), .B1(PHYADDRPOINTER_REG_24__SCAN_IN), 
        .B2(n5317), .ZN(n4094) );
  OAI211_X1 U5025 ( .C1(n3032), .C2(n4096), .A(n4095), .B(n4094), .ZN(n5454)
         );
  AND2_X2 U5026 ( .A1(n5453), .A2(n5454), .ZN(n5441) );
  AOI22_X1 U5027 ( .A1(n4121), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U5028 ( .A1(n4189), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4099) );
  AOI22_X1 U5029 ( .A1(n2985), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4098) );
  AOI22_X1 U5030 ( .A1(n2986), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4097) );
  NAND4_X1 U5031 ( .A1(n4100), .A2(n4099), .A3(n4098), .A4(n4097), .ZN(n4106)
         );
  AOI22_X1 U5032 ( .A1(n2984), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5033 ( .A1(n4194), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U5034 ( .A1(n5275), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5035 ( .A1(n5277), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4101) );
  NAND4_X1 U5036 ( .A1(n4104), .A2(n4103), .A3(n4102), .A4(n4101), .ZN(n4105)
         );
  NOR2_X1 U5037 ( .A1(n4106), .A2(n4105), .ZN(n4116) );
  NAND2_X1 U5038 ( .A1(n4108), .A2(n4107), .ZN(n4115) );
  XOR2_X1 U5039 ( .A(n4116), .B(n4115), .Z(n4109) );
  NAND2_X1 U5040 ( .A1(n4109), .A2(n4201), .ZN(n4114) );
  NAND2_X1 U5041 ( .A1(n6534), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4110)
         );
  NAND2_X1 U5042 ( .A1(n5294), .A2(n4110), .ZN(n4111) );
  AOI21_X1 U5043 ( .B1(n4204), .B2(EAX_REG_25__SCAN_IN), .A(n4111), .ZN(n4113)
         );
  XNOR2_X1 U5044 ( .A(n4143), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5613)
         );
  AND2_X1 U5045 ( .A1(n5613), .A2(n5288), .ZN(n4112) );
  AOI21_X1 U5046 ( .B1(n4114), .B2(n4113), .A(n4112), .ZN(n5442) );
  NOR2_X1 U5047 ( .A1(n4116), .A2(n4115), .ZN(n4149) );
  AOI22_X1 U5048 ( .A1(n2984), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U5049 ( .A1(n4194), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4119) );
  AOI22_X1 U5050 ( .A1(n5275), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U5051 ( .A1(n5277), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4117) );
  NAND4_X1 U5052 ( .A1(n4120), .A2(n4119), .A3(n4118), .A4(n4117), .ZN(n4127)
         );
  AOI22_X1 U5053 ( .A1(n4121), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5054 ( .A1(n4189), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5055 ( .A1(n2985), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5056 ( .A1(n2986), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4122) );
  NAND4_X1 U5057 ( .A1(n4125), .A2(n4124), .A3(n4123), .A4(n4122), .ZN(n4126)
         );
  OR2_X1 U5058 ( .A1(n4127), .A2(n4126), .ZN(n4147) );
  NAND2_X1 U5059 ( .A1(n4149), .A2(n4147), .ZN(n4160) );
  AOI22_X1 U5060 ( .A1(n4189), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n2986), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U5061 ( .A1(n2984), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U5062 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n5275), .B1(n5265), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U5063 ( .A1(n2985), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4128) );
  NAND4_X1 U5064 ( .A1(n4131), .A2(n4130), .A3(n4129), .A4(n4128), .ZN(n4137)
         );
  AOI22_X1 U5065 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4194), .B1(n4187), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U5066 ( .A1(n5273), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U5067 ( .A1(n4188), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U5068 ( .A1(n3239), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4132) );
  NAND4_X1 U5069 ( .A1(n4135), .A2(n4134), .A3(n4133), .A4(n4132), .ZN(n4136)
         );
  NOR2_X1 U5070 ( .A1(n4137), .A2(n4136), .ZN(n4161) );
  XOR2_X1 U5071 ( .A(n4160), .B(n4161), .Z(n4138) );
  NAND2_X1 U5072 ( .A1(n4138), .A2(n4201), .ZN(n4142) );
  NAND2_X1 U5073 ( .A1(n6534), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4139)
         );
  NAND2_X1 U5074 ( .A1(n5294), .A2(n4139), .ZN(n4140) );
  AOI21_X1 U5075 ( .B1(n4204), .B2(EAX_REG_27__SCAN_IN), .A(n4140), .ZN(n4141)
         );
  NAND2_X1 U5076 ( .A1(n4142), .A2(n4141), .ZN(n4146) );
  INV_X1 U5077 ( .A(n4143), .ZN(n4144) );
  XNOR2_X1 U5078 ( .A(n4177), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5423)
         );
  NAND2_X1 U5079 ( .A1(n5423), .A2(n5288), .ZN(n4145) );
  NAND2_X1 U5080 ( .A1(n4146), .A2(n4145), .ZN(n5422) );
  INV_X1 U5081 ( .A(n4147), .ZN(n4148) );
  XNOR2_X1 U5082 ( .A(n4149), .B(n4148), .ZN(n4153) );
  INV_X1 U5083 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4151) );
  NAND2_X1 U5084 ( .A1(n6534), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4150)
         );
  OAI211_X1 U5085 ( .C1(n3032), .C2(n4151), .A(n5294), .B(n4150), .ZN(n4152)
         );
  AOI21_X1 U5086 ( .B1(n4153), .B2(n4201), .A(n4152), .ZN(n4159) );
  INV_X1 U5087 ( .A(n4154), .ZN(n4156) );
  INV_X1 U5088 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4155) );
  NAND2_X1 U5089 ( .A1(n4156), .A2(n4155), .ZN(n4157) );
  NAND2_X1 U5090 ( .A1(n4177), .A2(n4157), .ZN(n5607) );
  NOR2_X1 U5091 ( .A1(n5607), .A2(n5294), .ZN(n4158) );
  OR2_X1 U5092 ( .A1(n4159), .A2(n4158), .ZN(n5308) );
  OR2_X1 U5093 ( .A1(n5422), .A2(n5308), .ZN(n5407) );
  NOR2_X1 U5094 ( .A1(n4161), .A2(n4160), .ZN(n4186) );
  AOI22_X1 U5095 ( .A1(n2984), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4165) );
  AOI22_X1 U5096 ( .A1(n4194), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U5097 ( .A1(n5275), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4163) );
  AOI22_X1 U5098 ( .A1(n3239), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4162) );
  NAND4_X1 U5099 ( .A1(n4165), .A2(n4164), .A3(n4163), .A4(n4162), .ZN(n4171)
         );
  AOI22_X1 U5100 ( .A1(n5273), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U5101 ( .A1(n4189), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U5102 ( .A1(n2985), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4167) );
  AOI22_X1 U5103 ( .A1(n2986), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4166) );
  NAND4_X1 U5104 ( .A1(n4169), .A2(n4168), .A3(n4167), .A4(n4166), .ZN(n4170)
         );
  OR2_X1 U5105 ( .A1(n4171), .A2(n4170), .ZN(n4185) );
  INV_X1 U5106 ( .A(n4185), .ZN(n4172) );
  XNOR2_X1 U5107 ( .A(n4186), .B(n4172), .ZN(n4176) );
  INV_X1 U5108 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4174) );
  NAND2_X1 U5109 ( .A1(n6534), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4173)
         );
  OAI211_X1 U5110 ( .C1(n3032), .C2(n4174), .A(n5294), .B(n4173), .ZN(n4175)
         );
  AOI21_X1 U5111 ( .B1(n4176), .B2(n4201), .A(n4175), .ZN(n4183) );
  INV_X1 U5112 ( .A(n4177), .ZN(n4178) );
  INV_X1 U5113 ( .A(n4179), .ZN(n4180) );
  INV_X1 U5114 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U5115 ( .A1(n4180), .A2(n5412), .ZN(n4181) );
  NAND2_X1 U5116 ( .A1(n4696), .A2(n4181), .ZN(n5592) );
  NOR2_X1 U5117 ( .A1(n5592), .A2(n5294), .ZN(n4182) );
  OR2_X1 U5118 ( .A1(n4183), .A2(n4182), .ZN(n5408) );
  NAND2_X1 U5119 ( .A1(n4186), .A2(n4185), .ZN(n5284) );
  AOI22_X1 U5120 ( .A1(n2985), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n2986), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4193) );
  AOI22_X1 U5121 ( .A1(n3239), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5275), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4192) );
  AOI22_X1 U5122 ( .A1(n2984), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4191) );
  AOI22_X1 U5123 ( .A1(n4189), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4190) );
  NAND4_X1 U5124 ( .A1(n4193), .A2(n4192), .A3(n4191), .A4(n4190), .ZN(n4200)
         );
  AOI22_X1 U5125 ( .A1(n4194), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4198) );
  AOI22_X1 U5126 ( .A1(n5276), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5268), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4197) );
  AOI22_X1 U5127 ( .A1(n5265), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4196) );
  AOI22_X1 U5128 ( .A1(n5273), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4195) );
  NAND4_X1 U5129 ( .A1(n4198), .A2(n4197), .A3(n4196), .A4(n4195), .ZN(n4199)
         );
  NOR2_X1 U5130 ( .A1(n4200), .A2(n4199), .ZN(n5285) );
  XOR2_X1 U5131 ( .A(n5284), .B(n5285), .Z(n4202) );
  NAND2_X1 U5132 ( .A1(n4202), .A2(n4201), .ZN(n4206) );
  INV_X1 U5133 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4695) );
  NOR2_X1 U5134 ( .A1(n4695), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4203) );
  AOI211_X1 U5135 ( .C1(n4204), .C2(EAX_REG_29__SCAN_IN), .A(n5288), .B(n4203), 
        .ZN(n4205) );
  XNOR2_X1 U5136 ( .A(n4696), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5376)
         );
  AOI22_X1 U5137 ( .A1(n4206), .A2(n4205), .B1(n5288), .B2(n5376), .ZN(n4208)
         );
  NAND3_X1 U5138 ( .A1(n6536), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6445) );
  INV_X1 U5139 ( .A(n6445), .ZN(n4209) );
  NOR2_X2 U5140 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6327) );
  NAND2_X1 U5141 ( .A1(n4209), .A2(n6327), .ZN(n5687) );
  NAND2_X1 U5142 ( .A1(n4210), .A2(n2983), .ZN(n4219) );
  INV_X1 U5143 ( .A(n6327), .ZN(n6332) );
  NAND2_X1 U5144 ( .A1(n6332), .A2(n4211), .ZN(n6539) );
  NAND2_X1 U5145 ( .A1(n6539), .A2(n6536), .ZN(n4212) );
  AND2_X2 U5146 ( .A1(n6060), .A2(n4212), .ZN(n6076) );
  NAND2_X1 U5147 ( .A1(n6536), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4214) );
  NAND2_X1 U5148 ( .A1(n6604), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4213) );
  AND2_X1 U5149 ( .A1(n4214), .A2(n4213), .ZN(n4408) );
  INV_X1 U5150 ( .A(n5376), .ZN(n4216) );
  INV_X1 U5151 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6738) );
  NOR2_X1 U5152 ( .A1(n6159), .A2(n6738), .ZN(n5709) );
  AOI21_X1 U5153 ( .B1(n6076), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5709), 
        .ZN(n4215) );
  OAI21_X1 U5154 ( .B1(n6085), .B2(n4216), .A(n4215), .ZN(n4217) );
  INV_X1 U5155 ( .A(n4217), .ZN(n4218) );
  OAI211_X1 U5156 ( .C1(n5717), .C2(n6060), .A(n4219), .B(n4218), .ZN(U2957)
         );
  OAI21_X1 U5157 ( .B1(n4263), .B2(n5714), .A(n4220), .ZN(n4221) );
  INV_X1 U5158 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4264) );
  XNOR2_X1 U5159 ( .A(n4221), .B(n4264), .ZN(n5299) );
  NAND2_X1 U5160 ( .A1(n3026), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4223) );
  NAND2_X1 U5161 ( .A1(n3638), .A2(EBX_REG_24__SCAN_IN), .ZN(n4222) );
  OAI211_X1 U5162 ( .C1(n4271), .C2(EBX_REG_24__SCAN_IN), .A(n4223), .B(n4222), 
        .ZN(n5458) );
  MUX2_X1 U5163 ( .A(n4232), .B(n5371), .S(EBX_REG_25__SCAN_IN), .Z(n4226) );
  NAND2_X1 U5164 ( .A1(n4242), .A2(n5750), .ZN(n4225) );
  NAND2_X1 U5165 ( .A1(n4226), .A2(n4225), .ZN(n5445) );
  INV_X1 U5166 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U5167 ( .A1(n4234), .A2(n5434), .ZN(n4230) );
  INV_X1 U5168 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U5169 ( .A1(n4236), .A2(n5588), .ZN(n4228) );
  NAND2_X1 U5170 ( .A1(n3022), .A2(n5434), .ZN(n4227) );
  NAND3_X1 U5171 ( .A1(n4228), .A2(n5371), .A3(n4227), .ZN(n4229) );
  AND2_X1 U5172 ( .A1(n4230), .A2(n4229), .ZN(n5313) );
  INV_X1 U5173 ( .A(n5313), .ZN(n4231) );
  NAND2_X1 U5174 ( .A1(n3006), .A2(n3004), .ZN(n5425) );
  MUX2_X1 U5175 ( .A(n4232), .B(n5371), .S(EBX_REG_27__SCAN_IN), .Z(n4233) );
  OAI21_X1 U5176 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n4344), .A(n4233), 
        .ZN(n5424) );
  OR2_X2 U5177 ( .A1(n5425), .A2(n5424), .ZN(n5427) );
  INV_X1 U5178 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U5179 ( .A1(n4234), .A2(n5510), .ZN(n4240) );
  INV_X1 U5180 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4235) );
  NAND2_X1 U5181 ( .A1(n4236), .A2(n4235), .ZN(n4238) );
  NAND2_X1 U5182 ( .A1(n3022), .A2(n5510), .ZN(n4237) );
  NAND3_X1 U5183 ( .A1(n4238), .A2(n5371), .A3(n4237), .ZN(n4239) );
  AND2_X1 U5184 ( .A1(n4240), .A2(n4239), .ZN(n5409) );
  INV_X1 U5185 ( .A(n5410), .ZN(n4248) );
  INV_X1 U5186 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5385) );
  AND2_X1 U5187 ( .A1(n3022), .A2(n5385), .ZN(n4241) );
  AOI21_X1 U5188 ( .B1(n4242), .B2(n5714), .A(n4241), .ZN(n5372) );
  INV_X1 U5189 ( .A(n4270), .ZN(n4247) );
  NAND2_X1 U5190 ( .A1(n4344), .A2(EBX_REG_30__SCAN_IN), .ZN(n4244) );
  NAND2_X1 U5191 ( .A1(n3026), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4243) );
  AND2_X1 U5192 ( .A1(n4244), .A2(n4243), .ZN(n4274) );
  INV_X1 U5193 ( .A(n4274), .ZN(n4246) );
  INV_X1 U5194 ( .A(n4273), .ZN(n4245) );
  INV_X1 U5195 ( .A(n4249), .ZN(n4251) );
  AOI211_X1 U5196 ( .C1(n5535), .C2(n4248), .A(n4246), .B(n4247), .ZN(n4250)
         );
  NOR2_X1 U5197 ( .A1(n4251), .A2(n4250), .ZN(n5349) );
  INV_X1 U5198 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6682) );
  NOR2_X1 U5199 ( .A1(n6159), .A2(n6682), .ZN(n5295) );
  INV_X1 U5200 ( .A(n4259), .ZN(n5724) );
  AND2_X1 U5201 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5718) );
  NAND2_X1 U5202 ( .A1(n5724), .A2(n5718), .ZN(n4255) );
  NAND2_X1 U5203 ( .A1(n4252), .A2(n6146), .ZN(n5778) );
  NAND2_X1 U5204 ( .A1(n5778), .A2(n4258), .ZN(n4253) );
  NAND2_X1 U5205 ( .A1(n4254), .A2(n4253), .ZN(n5760) );
  AOI21_X1 U5206 ( .B1(n6136), .B2(n4255), .A(n5760), .ZN(n5712) );
  OAI21_X1 U5207 ( .B1(n5760), .B2(n6136), .A(INSTADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n4256) );
  AOI21_X1 U5208 ( .B1(n5712), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n4256), 
        .ZN(n4257) );
  AOI211_X1 U5209 ( .C1(n6180), .C2(n5349), .A(n5295), .B(n4257), .ZN(n4261)
         );
  NAND2_X1 U5210 ( .A1(n5751), .A2(n5718), .ZN(n5734) );
  NOR2_X1 U5211 ( .A1(n5734), .A2(n4259), .ZN(n5715) );
  NAND3_X1 U5212 ( .A1(n5715), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n4264), .ZN(n4260) );
  OAI21_X1 U5213 ( .B1(n5299), .B2(n6157), .A(n4262), .ZN(U2988) );
  NAND2_X1 U5214 ( .A1(n4263), .A2(n3039), .ZN(n4267) );
  INV_X1 U5215 ( .A(n5611), .ZN(n4266) );
  NAND4_X1 U5216 ( .A1(n5586), .A2(n5725), .A3(n4264), .A4(n5714), .ZN(n4265)
         );
  NAND2_X1 U5217 ( .A1(n4267), .A2(n3036), .ZN(n4268) );
  XNOR2_X1 U5218 ( .A(n4268), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5368)
         );
  INV_X1 U5219 ( .A(n6136), .ZN(n6102) );
  OAI21_X1 U5220 ( .B1(n6102), .B2(n3039), .A(n5712), .ZN(n4269) );
  INV_X1 U5221 ( .A(n4269), .ZN(n4280) );
  INV_X1 U5222 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4279) );
  INV_X1 U5223 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6655) );
  NOR2_X1 U5224 ( .A1(n6159), .A2(n6655), .ZN(n5363) );
  INV_X1 U5225 ( .A(n5363), .ZN(n4278) );
  NOR2_X1 U5226 ( .A1(n4271), .A2(EBX_REG_29__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U5227 ( .A1(n5410), .A2(n5370), .ZN(n4272) );
  OAI22_X1 U5228 ( .A1(n4344), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n3026), .ZN(n4275) );
  INV_X1 U5229 ( .A(n4275), .ZN(n4276) );
  INV_X1 U5230 ( .A(n4281), .ZN(n4283) );
  NAND3_X1 U5231 ( .A1(n5715), .A2(n3039), .A3(n4279), .ZN(n4282) );
  OAI21_X1 U5232 ( .B1(n5368), .B2(n6157), .A(n4284), .ZN(U2987) );
  NOR2_X1 U5233 ( .A1(n4285), .A2(n5399), .ZN(n4290) );
  INV_X1 U5234 ( .A(n4290), .ZN(n4286) );
  AOI22_X1 U5235 ( .A1(n5404), .A2(n3510), .B1(n5396), .B2(n4286), .ZN(n5406)
         );
  INV_X1 U5236 ( .A(n6438), .ZN(n6426) );
  AND2_X1 U5237 ( .A1(n5406), .A2(n6426), .ZN(n4289) );
  INV_X1 U5238 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n4288) );
  NOR2_X1 U5239 ( .A1(n6332), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4292) );
  NAND2_X1 U5240 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4292), .ZN(n4287) );
  OAI21_X1 U5241 ( .B1(n4289), .B2(n4288), .A(n4287), .ZN(U2790) );
  NAND2_X1 U5242 ( .A1(n4290), .A2(n6426), .ZN(n4690) );
  INV_X1 U5243 ( .A(n4690), .ZN(n4294) );
  INV_X1 U5244 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n4293) );
  INV_X1 U5245 ( .A(n5396), .ZN(n4291) );
  INV_X1 U5246 ( .A(n4292), .ZN(n5391) );
  OAI211_X1 U5247 ( .C1(n4294), .C2(n4293), .A(n4691), .B(n5391), .ZN(U2788)
         );
  INV_X1 U5248 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6029) );
  INV_X1 U5249 ( .A(READY_N), .ZN(n6638) );
  INV_X1 U5250 ( .A(n4691), .ZN(n4295) );
  OAI21_X1 U5251 ( .B1(n3359), .B2(n6638), .A(n4295), .ZN(n4327) );
  NAND2_X1 U5252 ( .A1(n4327), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4297) );
  NAND2_X1 U5253 ( .A1(n3022), .A2(n6638), .ZN(n4296) );
  NOR2_X1 U5254 ( .A1(n4313), .A2(n4296), .ZN(n4315) );
  NAND2_X1 U5255 ( .A1(n4740), .A2(n4315), .ZN(n4395) );
  NAND2_X1 U5256 ( .A1(n4373), .A2(DATAI_10_), .ZN(n4340) );
  OAI211_X1 U5257 ( .C1(n6029), .C2(n4355), .A(n4297), .B(n4340), .ZN(U2949)
         );
  INV_X1 U5258 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U5259 ( .A1(n4327), .A2(LWORD_REG_9__SCAN_IN), .ZN(n4298) );
  NAND2_X1 U5260 ( .A1(n4373), .A2(DATAI_9_), .ZN(n4337) );
  OAI211_X1 U5261 ( .C1(n6031), .C2(n4355), .A(n4298), .B(n4337), .ZN(U2948)
         );
  AND4_X1 U5262 ( .A1(n4300), .A2(n5903), .A3(n4313), .A4(n3601), .ZN(n4301)
         );
  AND2_X1 U5263 ( .A1(n4302), .A2(n4301), .ZN(n5823) );
  INV_X1 U5264 ( .A(n5823), .ZN(n5339) );
  XNOR2_X1 U5265 ( .A(n5818), .B(n4416), .ZN(n4307) );
  INV_X1 U5266 ( .A(n4316), .ZN(n5403) );
  NAND2_X1 U5267 ( .A1(n5403), .A2(n5395), .ZN(n4427) );
  NAND2_X1 U5268 ( .A1(n4427), .A2(n4307), .ZN(n4306) );
  NAND2_X1 U5269 ( .A1(n6399), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4304) );
  NAND2_X1 U5270 ( .A1(n6399), .A2(n3181), .ZN(n5822) );
  MUX2_X1 U5271 ( .A(n4304), .B(n5822), .S(n4416), .Z(n4305) );
  OAI211_X1 U5272 ( .C1(n4307), .C2(n4418), .A(n4306), .B(n4305), .ZN(n4308)
         );
  AOI21_X1 U5273 ( .B1(n5806), .B2(n5339), .A(n4308), .ZN(n4430) );
  INV_X1 U5274 ( .A(n4430), .ZN(n4312) );
  NOR2_X1 U5275 ( .A1(n5340), .A2(n4309), .ZN(n5826) );
  INV_X1 U5276 ( .A(n5826), .ZN(n5341) );
  AOI22_X1 U5277 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4279), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4447), .ZN(n5825) );
  INV_X1 U5278 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6519) );
  NAND3_X1 U5279 ( .A1(n5818), .A2(n6521), .A3(n3291), .ZN(n4310) );
  OAI21_X1 U5280 ( .B1(n5341), .B2(n5825), .A(n4310), .ZN(n4311) );
  AOI21_X1 U5281 ( .B1(n4312), .B2(n6522), .A(n4311), .ZN(n4326) );
  NAND2_X1 U5282 ( .A1(n6536), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6517) );
  INV_X1 U5283 ( .A(n4710), .ZN(n6455) );
  AND2_X1 U5284 ( .A1(n6455), .A2(n6638), .ZN(n4314) );
  OAI22_X1 U5285 ( .A1(n6399), .A2(n3185), .B1(n4315), .B2(n4314), .ZN(n4320)
         );
  NAND2_X1 U5286 ( .A1(n5404), .A2(n4316), .ZN(n4349) );
  NOR2_X1 U5287 ( .A1(n4318), .A2(n4317), .ZN(n4319) );
  OAI211_X1 U5288 ( .C1(n5404), .C2(n4320), .A(n4349), .B(n4319), .ZN(n4323)
         );
  INV_X1 U5289 ( .A(n4321), .ZN(n4322) );
  OAI22_X1 U5290 ( .A1(n5404), .A2(n5395), .B1(n5903), .B2(n4322), .ZN(n4388)
         );
  OR2_X1 U5291 ( .A1(n4323), .A2(n4388), .ZN(n6404) );
  INV_X1 U5292 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6551) );
  NAND2_X1 U5293 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4743) );
  NOR2_X1 U5294 ( .A1(n6536), .A2(n4743), .ZN(n4439) );
  INV_X1 U5295 ( .A(n4439), .ZN(n6516) );
  NOR2_X1 U5296 ( .A1(n6551), .A2(n6516), .ZN(n4324) );
  AOI21_X1 U5297 ( .B1(n6404), .B2(n6426), .A(n4324), .ZN(n5902) );
  NAND2_X1 U5298 ( .A1(n6517), .A2(n5902), .ZN(n6525) );
  INV_X1 U5299 ( .A(n6525), .ZN(n5343) );
  INV_X1 U5300 ( .A(n6521), .ZN(n6433) );
  NOR2_X1 U5301 ( .A1(n5818), .A2(n6433), .ZN(n5828) );
  OAI21_X1 U5302 ( .B1(n5343), .B2(n5828), .A(n4416), .ZN(n4325) );
  OAI21_X1 U5303 ( .B1(n4326), .B2(n5343), .A(n4325), .ZN(U3459) );
  INV_X1 U5304 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6036) );
  INV_X1 U5305 ( .A(n4327), .ZN(n4393) );
  NAND2_X1 U5306 ( .A1(n4372), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4328) );
  NAND2_X1 U5307 ( .A1(n4373), .A2(DATAI_6_), .ZN(n4342) );
  OAI211_X1 U5308 ( .C1(n6036), .C2(n4355), .A(n4328), .B(n4342), .ZN(U2945)
         );
  INV_X1 U5309 ( .A(EAX_REG_23__SCAN_IN), .ZN(n5099) );
  NAND2_X1 U5310 ( .A1(n4327), .A2(UWORD_REG_7__SCAN_IN), .ZN(n4329) );
  NAND2_X1 U5311 ( .A1(n4373), .A2(DATAI_7_), .ZN(n4356) );
  OAI211_X1 U5312 ( .C1(n5099), .C2(n4355), .A(n4329), .B(n4356), .ZN(U2931)
         );
  INV_X1 U5313 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6025) );
  NAND2_X1 U5314 ( .A1(n4372), .A2(LWORD_REG_12__SCAN_IN), .ZN(n4330) );
  NAND2_X1 U5315 ( .A1(n4373), .A2(DATAI_12_), .ZN(n4366) );
  OAI211_X1 U5316 ( .C1(n6025), .C2(n4355), .A(n4330), .B(n4366), .ZN(U2951)
         );
  INV_X1 U5317 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U5318 ( .A1(n4327), .A2(LWORD_REG_11__SCAN_IN), .ZN(n4331) );
  NAND2_X1 U5319 ( .A1(n4373), .A2(DATAI_11_), .ZN(n4361) );
  OAI211_X1 U5320 ( .C1(n6027), .C2(n4355), .A(n4331), .B(n4361), .ZN(U2950)
         );
  INV_X1 U5321 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U5322 ( .A1(n4372), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4332) );
  NAND2_X1 U5323 ( .A1(n4373), .A2(DATAI_8_), .ZN(n4333) );
  OAI211_X1 U5324 ( .C1(n6033), .C2(n4355), .A(n4332), .B(n4333), .ZN(U2947)
         );
  NAND2_X1 U5325 ( .A1(n4327), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4334) );
  OAI211_X1 U5326 ( .C1(n4096), .C2(n4355), .A(n4334), .B(n4333), .ZN(U2932)
         );
  INV_X1 U5327 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U5328 ( .A1(n4372), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4335) );
  NAND2_X1 U5329 ( .A1(n4373), .A2(DATAI_14_), .ZN(n4363) );
  OAI211_X1 U5330 ( .C1(n6021), .C2(n4355), .A(n4335), .B(n4363), .ZN(U2953)
         );
  INV_X1 U5331 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U5332 ( .A1(n4327), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4336) );
  NAND2_X1 U5333 ( .A1(n4373), .A2(DATAI_13_), .ZN(n4358) );
  OAI211_X1 U5334 ( .C1(n6023), .C2(n4355), .A(n4336), .B(n4358), .ZN(U2952)
         );
  INV_X1 U5335 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4754) );
  NAND2_X1 U5336 ( .A1(n4327), .A2(UWORD_REG_9__SCAN_IN), .ZN(n4338) );
  OAI211_X1 U5337 ( .C1(n4754), .C2(n4355), .A(n4338), .B(n4337), .ZN(U2933)
         );
  NAND2_X1 U5338 ( .A1(n4372), .A2(LWORD_REG_5__SCAN_IN), .ZN(n4339) );
  NAND2_X1 U5339 ( .A1(n4373), .A2(DATAI_5_), .ZN(n4381) );
  OAI211_X1 U5340 ( .C1(n3789), .C2(n4355), .A(n4339), .B(n4381), .ZN(U2944)
         );
  NAND2_X1 U5341 ( .A1(n4327), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4341) );
  OAI211_X1 U5342 ( .C1(n4151), .C2(n4355), .A(n4341), .B(n4340), .ZN(U2934)
         );
  INV_X1 U5343 ( .A(EAX_REG_22__SCAN_IN), .ZN(n5102) );
  NAND2_X1 U5344 ( .A1(n4327), .A2(UWORD_REG_6__SCAN_IN), .ZN(n4343) );
  OAI211_X1 U5345 ( .C1(n5102), .C2(n4355), .A(n4343), .B(n4342), .ZN(U2930)
         );
  NOR2_X1 U5346 ( .A1(n4344), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4345)
         );
  NOR2_X1 U5347 ( .A1(n4346), .A2(n4345), .ZN(n4404) );
  INV_X1 U5348 ( .A(n4404), .ZN(n4726) );
  INV_X1 U5349 ( .A(n3583), .ZN(n4347) );
  AND2_X1 U5350 ( .A1(n5387), .A2(n3175), .ZN(n4385) );
  NAND4_X1 U5351 ( .A1(n4347), .A2(n3208), .A3(n3022), .A4(n4385), .ZN(n4348)
         );
  NAND2_X1 U5352 ( .A1(n4349), .A2(n4348), .ZN(n4350) );
  INV_X1 U5353 ( .A(n4351), .ZN(n4354) );
  OAI21_X1 U5354 ( .B1(n4354), .B2(n4353), .A(n4352), .ZN(n4731) );
  AND2_X1 U5355 ( .A1(n6009), .A2(n4499), .ZN(n6006) );
  OAI222_X1 U5356 ( .A1(n4726), .A2(n5549), .B1(n4725), .B2(n6009), .C1(n4731), 
        .C2(n5553), .ZN(U2859) );
  NAND2_X1 U5357 ( .A1(n4372), .A2(LWORD_REG_7__SCAN_IN), .ZN(n4357) );
  OAI211_X1 U5358 ( .C1(n3801), .C2(n4355), .A(n4357), .B(n4356), .ZN(U2946)
         );
  INV_X1 U5359 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4751) );
  NAND2_X1 U5360 ( .A1(n4372), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4359) );
  OAI211_X1 U5361 ( .C1(n4751), .C2(n4355), .A(n4359), .B(n4358), .ZN(U2937)
         );
  INV_X1 U5362 ( .A(EAX_REG_16__SCAN_IN), .ZN(n5090) );
  NAND2_X1 U5363 ( .A1(n4327), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4360) );
  NAND2_X1 U5364 ( .A1(n4373), .A2(DATAI_0_), .ZN(n4370) );
  OAI211_X1 U5365 ( .C1(n5090), .C2(n4355), .A(n4360), .B(n4370), .ZN(U2924)
         );
  INV_X1 U5366 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4748) );
  NAND2_X1 U5367 ( .A1(n4372), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4362) );
  OAI211_X1 U5368 ( .C1(n4748), .C2(n4355), .A(n4362), .B(n4361), .ZN(U2935)
         );
  INV_X1 U5369 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4745) );
  NAND2_X1 U5370 ( .A1(n4372), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4364) );
  OAI211_X1 U5371 ( .C1(n4745), .C2(n4355), .A(n4364), .B(n4363), .ZN(U2938)
         );
  INV_X1 U5372 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U5373 ( .A1(n4372), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4365) );
  NAND2_X1 U5374 ( .A1(n4373), .A2(DATAI_4_), .ZN(n4375) );
  OAI211_X1 U5375 ( .C1(n6040), .C2(n4355), .A(n4365), .B(n4375), .ZN(U2943)
         );
  NAND2_X1 U5376 ( .A1(n4372), .A2(UWORD_REG_12__SCAN_IN), .ZN(n4367) );
  OAI211_X1 U5377 ( .C1(n4174), .C2(n4355), .A(n4367), .B(n4366), .ZN(U2936)
         );
  INV_X1 U5378 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U5379 ( .A1(n4372), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4368) );
  NAND2_X1 U5380 ( .A1(n4373), .A2(DATAI_2_), .ZN(n4379) );
  OAI211_X1 U5381 ( .C1(n6044), .C2(n4355), .A(n4368), .B(n4379), .ZN(U2941)
         );
  INV_X1 U5382 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U5383 ( .A1(n4372), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4369) );
  NAND2_X1 U5384 ( .A1(n4373), .A2(DATAI_1_), .ZN(n4383) );
  OAI211_X1 U5385 ( .C1(n6046), .C2(n4355), .A(n4369), .B(n4383), .ZN(U2940)
         );
  INV_X1 U5386 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U5387 ( .A1(n4372), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4371) );
  OAI211_X1 U5388 ( .C1(n6050), .C2(n4355), .A(n4371), .B(n4370), .ZN(U2939)
         );
  INV_X1 U5389 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U5390 ( .A1(n4372), .A2(LWORD_REG_3__SCAN_IN), .ZN(n4374) );
  NAND2_X1 U5391 ( .A1(n4373), .A2(DATAI_3_), .ZN(n4377) );
  OAI211_X1 U5392 ( .C1(n6042), .C2(n4355), .A(n4374), .B(n4377), .ZN(U2942)
         );
  NAND2_X1 U5393 ( .A1(n4372), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4376) );
  OAI211_X1 U5394 ( .C1(n4004), .C2(n4355), .A(n4376), .B(n4375), .ZN(U2928)
         );
  INV_X1 U5395 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U5396 ( .A1(n4372), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4378) );
  OAI211_X1 U5397 ( .C1(n5094), .C2(n4355), .A(n4378), .B(n4377), .ZN(U2927)
         );
  NAND2_X1 U5398 ( .A1(n4372), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4380) );
  OAI211_X1 U5399 ( .C1(n3970), .C2(n4355), .A(n4380), .B(n4379), .ZN(U2926)
         );
  INV_X1 U5400 ( .A(EAX_REG_21__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U5401 ( .A1(n4372), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4382) );
  OAI211_X1 U5402 ( .C1(n5097), .C2(n4355), .A(n4382), .B(n4381), .ZN(U2929)
         );
  NAND2_X1 U5403 ( .A1(n4372), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4384) );
  OAI211_X1 U5404 ( .C1(n3951), .C2(n4355), .A(n4384), .B(n4383), .ZN(U2925)
         );
  NAND2_X1 U5405 ( .A1(n4385), .A2(n4503), .ZN(n4386) );
  NOR2_X1 U5406 ( .A1(n3601), .A2(n4386), .ZN(n4387) );
  OR2_X1 U5407 ( .A1(n4388), .A2(n4387), .ZN(n4389) );
  NAND2_X1 U5408 ( .A1(n4389), .A2(n6426), .ZN(n4390) );
  AND2_X1 U5409 ( .A1(n5581), .A2(n4391), .ZN(n6011) );
  INV_X2 U5410 ( .A(n6011), .ZN(n5583) );
  INV_X1 U5411 ( .A(n4391), .ZN(n4392) );
  NAND2_X1 U5412 ( .A1(n5581), .A2(n4392), .ZN(n5582) );
  INV_X1 U5413 ( .A(DATAI_0_), .ZN(n6643) );
  OAI222_X1 U5414 ( .A1(n4731), .A2(n5583), .B1(n5582), .B2(n6643), .C1(n5581), 
        .C2(n6050), .ZN(U2891) );
  INV_X1 U5415 ( .A(DATAI_15_), .ZN(n4396) );
  INV_X1 U5416 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6019) );
  INV_X1 U5417 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4394) );
  OAI222_X1 U5418 ( .A1(n4396), .A2(n4395), .B1(n4355), .B2(n6019), .C1(n4394), 
        .C2(n4393), .ZN(U2954) );
  INV_X1 U5419 ( .A(n4398), .ZN(n4399) );
  OAI21_X1 U5420 ( .B1(n4400), .B2(n4397), .A(n4399), .ZN(n5003) );
  INV_X1 U5421 ( .A(n6006), .ZN(n5348) );
  XNOR2_X1 U5422 ( .A(n3015), .B(n3026), .ZN(n4997) );
  INV_X1 U5423 ( .A(n4997), .ZN(n4401) );
  OAI222_X1 U5424 ( .A1(n5003), .A2(n5348), .B1(n6009), .B2(n4995), .C1(n4401), 
        .C2(n5549), .ZN(U2858) );
  INV_X1 U5425 ( .A(DATAI_1_), .ZN(n4491) );
  OAI222_X1 U5426 ( .A1(n5003), .A2(n5583), .B1(n5582), .B2(n4491), .C1(n5581), 
        .C2(n6046), .ZN(U2890) );
  XNOR2_X1 U5427 ( .A(n4402), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4413)
         );
  NAND2_X1 U5428 ( .A1(n6146), .A2(n5196), .ZN(n5197) );
  INV_X1 U5429 ( .A(n5200), .ZN(n4403) );
  OAI21_X1 U5430 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n6146), .A(n6132), 
        .ZN(n4449) );
  OAI22_X1 U5431 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5197), .B1(n4403), 
        .B2(n4449), .ZN(n4406) );
  AND2_X1 U5432 ( .A1(n6185), .A2(REIP_REG_0__SCAN_IN), .ZN(n4410) );
  AOI21_X1 U5433 ( .B1(n6180), .B2(n4404), .A(n4410), .ZN(n4405) );
  OAI211_X1 U5434 ( .C1(n4413), .C2(n6157), .A(n4406), .B(n4405), .ZN(U3018)
         );
  INV_X1 U5435 ( .A(n4731), .ZN(n4411) );
  INV_X1 U5436 ( .A(n6076), .ZN(n5681) );
  INV_X1 U5437 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4407) );
  AOI21_X1 U5438 ( .B1(n5681), .B2(n4408), .A(n4407), .ZN(n4409) );
  AOI211_X1 U5439 ( .C1(n4411), .C2(n2983), .A(n4410), .B(n4409), .ZN(n4412)
         );
  OAI21_X1 U5440 ( .B1(n4413), .B2(n6060), .A(n4412), .ZN(U2986) );
  INV_X1 U5441 ( .A(n4415), .ZN(n5993) );
  NAND2_X1 U5442 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n4416), .ZN(n4417) );
  NAND2_X1 U5443 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n4417), .ZN(n4419) );
  OAI21_X1 U5444 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n4417), .A(n4419), 
        .ZN(n4421) );
  INV_X1 U5445 ( .A(n4418), .ZN(n4420) );
  NAND3_X1 U5446 ( .A1(n3298), .A2(n3299), .A3(n4419), .ZN(n6520) );
  AOI22_X1 U5447 ( .A1(n6399), .A2(n4421), .B1(n4420), .B2(n6520), .ZN(n4429)
         );
  INV_X1 U5448 ( .A(n4422), .ZN(n4426) );
  INV_X1 U5449 ( .A(n4423), .ZN(n4424) );
  MUX2_X1 U5450 ( .A(n4424), .B(n3319), .S(n5818), .Z(n4425) );
  NAND3_X1 U5451 ( .A1(n4427), .A2(n4426), .A3(n4425), .ZN(n4428) );
  OAI211_X1 U5452 ( .C1(n5993), .C2(n5823), .A(n4429), .B(n4428), .ZN(n6523)
         );
  MUX2_X1 U5453 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6523), .S(n6404), 
        .Z(n6410) );
  MUX2_X1 U5454 ( .A(n3291), .B(n4430), .S(n6404), .Z(n6408) );
  NOR2_X1 U5455 ( .A1(n6408), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4432) );
  NOR2_X1 U5456 ( .A1(FLUSH_REG_SCAN_IN), .A2(n5340), .ZN(n4431) );
  AOI22_X1 U5457 ( .A1(n6410), .A2(n4432), .B1(n4422), .B2(n4431), .ZN(n6421)
         );
  INV_X1 U5458 ( .A(n6404), .ZN(n4434) );
  MUX2_X1 U5459 ( .A(n6551), .B(n4434), .S(n5340), .Z(n4438) );
  INV_X1 U5460 ( .A(n4853), .ZN(n6239) );
  NOR2_X1 U5461 ( .A1(n4435), .A2(n6239), .ZN(n4436) );
  XNOR2_X1 U5462 ( .A(n4436), .B(n5908), .ZN(n5904) );
  NOR2_X1 U5463 ( .A1(n5903), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4437) );
  AOI22_X1 U5464 ( .A1(n4438), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(n5904), .B2(n4437), .ZN(n6420) );
  OAI21_X1 U5465 ( .B1(n6421), .B2(n4433), .A(n6420), .ZN(n4441) );
  OAI21_X1 U5466 ( .B1(n4441), .B2(FLUSH_REG_SCAN_IN), .A(n4439), .ZN(n4440)
         );
  NOR2_X1 U5467 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6447) );
  INV_X1 U5468 ( .A(n6447), .ZN(n6535) );
  NAND2_X1 U5469 ( .A1(n4440), .A2(n4515), .ZN(n6191) );
  NOR2_X1 U5470 ( .A1(n4441), .A2(n4743), .ZN(n6432) );
  INV_X1 U5471 ( .A(n6330), .ZN(n4857) );
  AND2_X1 U5472 ( .A1(n6519), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5812) );
  OAI22_X1 U5473 ( .A1(n5046), .A2(n6332), .B1(n4857), .B2(n5812), .ZN(n4442)
         );
  OAI21_X1 U5474 ( .B1(n6432), .B2(n4442), .A(n6191), .ZN(n4443) );
  OAI21_X1 U5475 ( .B1(n6191), .B2(n6398), .A(n4443), .ZN(U3465) );
  XNOR2_X1 U5476 ( .A(n4445), .B(n4444), .ZN(n4897) );
  INV_X1 U5477 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6527) );
  NOR2_X1 U5478 ( .A1(n6159), .A2(n6527), .ZN(n4892) );
  NOR2_X1 U5479 ( .A1(n6102), .A2(n4446), .ZN(n4448) );
  MUX2_X1 U5480 ( .A(n4449), .B(n4448), .S(n4447), .Z(n4450) );
  AOI211_X1 U5481 ( .C1(n6180), .C2(n4997), .A(n4892), .B(n4450), .ZN(n4451)
         );
  OAI21_X1 U5482 ( .B1(n4897), .B2(n6157), .A(n4451), .ZN(U3017) );
  CLKBUF_X1 U5483 ( .A(n4452), .Z(n4453) );
  NOR2_X1 U5484 ( .A1(n4454), .A2(n4455), .ZN(n4456) );
  NOR2_X1 U5485 ( .A1(n4453), .A2(n4456), .ZN(n6080) );
  INV_X1 U5486 ( .A(n6080), .ZN(n4959) );
  XOR2_X1 U5487 ( .A(n4458), .B(n4457), .Z(n6181) );
  INV_X1 U5488 ( .A(n6009), .ZN(n5551) );
  AOI22_X1 U5489 ( .A1(n6181), .A2(n6005), .B1(EBX_REG_2__SCAN_IN), .B2(n5551), 
        .ZN(n4459) );
  OAI21_X1 U5490 ( .B1(n4959), .B2(n5348), .A(n4459), .ZN(U2857) );
  INV_X1 U5491 ( .A(DATAI_2_), .ZN(n4469) );
  OAI222_X1 U5492 ( .A1(n4959), .A2(n5583), .B1(n5582), .B2(n4469), .C1(n5581), 
        .C2(n6044), .ZN(U2889) );
  OAI21_X1 U5493 ( .B1(n4453), .B2(n4460), .A(n4580), .ZN(n5988) );
  AOI21_X1 U5494 ( .B1(n4463), .B2(n4462), .A(n4461), .ZN(n6169) );
  AOI22_X1 U5495 ( .A1(n6005), .A2(n6169), .B1(n5551), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4464) );
  OAI21_X1 U5496 ( .B1(n5988), .B2(n5348), .A(n4464), .ZN(U2856) );
  INV_X1 U5497 ( .A(DATAI_3_), .ZN(n6688) );
  OAI222_X1 U5498 ( .A1(n5988), .A2(n5583), .B1(n5582), .B2(n6688), .C1(n5581), 
        .C2(n6042), .ZN(U2888) );
  AND2_X1 U5499 ( .A1(n4415), .A2(n6330), .ZN(n4757) );
  AND2_X1 U5500 ( .A1(n4466), .A2(n5806), .ZN(n6240) );
  INV_X1 U5501 ( .A(n4467), .ZN(n4510) );
  AOI21_X1 U5502 ( .B1(n4757), .B2(n6240), .A(n4510), .ZN(n4475) );
  INV_X1 U5503 ( .A(n4475), .ZN(n4468) );
  AOI22_X1 U5504 ( .A1(n4468), .A2(n6327), .B1(n4544), .B2(
        STATE2_REG_2__SCAN_IN), .ZN(n4513) );
  NOR2_X1 U5505 ( .A1(n4469), .A2(n4515), .ZN(n6350) );
  INV_X1 U5506 ( .A(n6350), .ZN(n5166) );
  AOI21_X1 U5507 ( .B1(n6398), .B2(STATE2_REG_3__SCAN_IN), .A(n4515), .ZN(
        n6278) );
  INV_X1 U5508 ( .A(n5805), .ZN(n6194) );
  INV_X1 U5509 ( .A(n4472), .ZN(n4473) );
  NOR3_X1 U5510 ( .A1(n6194), .A2(n4542), .A3(n4473), .ZN(n4474) );
  NAND2_X1 U5511 ( .A1(n6327), .A2(n6604), .ZN(n5815) );
  OAI21_X1 U5512 ( .B1(n4474), .B2(n5687), .A(n5815), .ZN(n4476) );
  NAND2_X1 U5513 ( .A1(n4476), .A2(n4475), .ZN(n4477) );
  OAI211_X1 U5514 ( .C1(n4544), .C2(n6327), .A(n6278), .B(n4477), .ZN(n4507)
         );
  NAND2_X1 U5515 ( .A1(n4507), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4484)
         );
  NAND2_X1 U5516 ( .A1(n4508), .A2(n3189), .ZN(n5162) );
  INV_X1 U5517 ( .A(n5162), .ZN(n6349) );
  NAND2_X1 U5518 ( .A1(n2983), .A2(DATAI_18_), .ZN(n6353) );
  NAND2_X1 U5519 ( .A1(n4472), .A2(n3386), .ZN(n4902) );
  INV_X1 U5520 ( .A(n4902), .ZN(n4479) );
  NAND3_X1 U5521 ( .A1(n4479), .A2(n5805), .A3(n4480), .ZN(n4683) );
  NAND2_X1 U5522 ( .A1(n4472), .A2(n5046), .ZN(n6233) );
  INV_X1 U5523 ( .A(n6233), .ZN(n4481) );
  NAND3_X1 U5524 ( .A1(n4481), .A2(n5805), .A3(n4480), .ZN(n4570) );
  NAND2_X1 U5525 ( .A1(n2983), .A2(DATAI_26_), .ZN(n6293) );
  OAI22_X1 U5526 ( .A1(n6353), .A2(n4683), .B1(n4570), .B2(n6293), .ZN(n4482)
         );
  AOI21_X1 U5527 ( .B1(n6349), .B2(n4510), .A(n4482), .ZN(n4483) );
  OAI211_X1 U5528 ( .C1(n4513), .C2(n5166), .A(n4484), .B(n4483), .ZN(U3142)
         );
  NOR2_X1 U5529 ( .A1(n6688), .A2(n4515), .ZN(n6390) );
  INV_X1 U5530 ( .A(n6390), .ZN(n5176) );
  NAND2_X1 U5531 ( .A1(n4507), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4487)
         );
  NAND2_X1 U5532 ( .A1(n4508), .A2(n3190), .ZN(n5172) );
  NAND2_X1 U5533 ( .A1(n2983), .A2(DATAI_19_), .ZN(n6255) );
  NAND2_X1 U5534 ( .A1(n2983), .A2(DATAI_27_), .ZN(n6397) );
  OAI22_X1 U5535 ( .A1(n6255), .A2(n4683), .B1(n4570), .B2(n6397), .ZN(n4485)
         );
  AOI21_X1 U5536 ( .B1(n6388), .B2(n4510), .A(n4485), .ZN(n4486) );
  OAI211_X1 U5537 ( .C1(n4513), .C2(n5176), .A(n4487), .B(n4486), .ZN(U3143)
         );
  NOR2_X1 U5538 ( .A1(n6643), .A2(n4515), .ZN(n6338) );
  INV_X1 U5539 ( .A(n6338), .ZN(n5146) );
  NAND2_X1 U5540 ( .A1(n4507), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4490)
         );
  NAND2_X1 U5541 ( .A1(n4508), .A2(n3602), .ZN(n5142) );
  INV_X1 U5542 ( .A(n5142), .ZN(n6326) );
  NAND2_X1 U5543 ( .A1(n2983), .A2(DATAI_16_), .ZN(n6341) );
  NAND2_X1 U5544 ( .A1(n2983), .A2(DATAI_24_), .ZN(n6285) );
  OAI22_X1 U5545 ( .A1(n6341), .A2(n4683), .B1(n4570), .B2(n6285), .ZN(n4488)
         );
  AOI21_X1 U5546 ( .B1(n6326), .B2(n4510), .A(n4488), .ZN(n4489) );
  OAI211_X1 U5547 ( .C1(n4513), .C2(n5146), .A(n4490), .B(n4489), .ZN(U3140)
         );
  NOR2_X1 U5548 ( .A1(n4491), .A2(n4515), .ZN(n6344) );
  INV_X1 U5549 ( .A(n6344), .ZN(n5184) );
  NAND2_X1 U5550 ( .A1(n4507), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4495)
         );
  NAND2_X1 U5551 ( .A1(n4508), .A2(n4492), .ZN(n5179) );
  INV_X1 U5552 ( .A(n5179), .ZN(n6343) );
  NAND2_X1 U5553 ( .A1(n2983), .A2(DATAI_17_), .ZN(n6347) );
  NAND2_X1 U5554 ( .A1(n2983), .A2(DATAI_25_), .ZN(n6289) );
  OAI22_X1 U5555 ( .A1(n6347), .A2(n4683), .B1(n4570), .B2(n6289), .ZN(n4493)
         );
  AOI21_X1 U5556 ( .B1(n6343), .B2(n4510), .A(n4493), .ZN(n4494) );
  OAI211_X1 U5557 ( .C1(n4513), .C2(n5184), .A(n4495), .B(n4494), .ZN(U3141)
         );
  INV_X1 U5558 ( .A(DATAI_5_), .ZN(n6674) );
  NOR2_X1 U5559 ( .A1(n6674), .A2(n4515), .ZN(n6364) );
  INV_X1 U5560 ( .A(n6364), .ZN(n5156) );
  NAND2_X1 U5561 ( .A1(n4507), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4498)
         );
  NAND2_X1 U5562 ( .A1(n4508), .A2(n5259), .ZN(n5152) );
  INV_X1 U5563 ( .A(n5152), .ZN(n6363) );
  NAND2_X1 U5564 ( .A1(n2983), .A2(DATAI_21_), .ZN(n6367) );
  NAND2_X1 U5565 ( .A1(n2983), .A2(DATAI_29_), .ZN(n6323) );
  OAI22_X1 U5566 ( .A1(n6367), .A2(n4683), .B1(n4570), .B2(n6323), .ZN(n4496)
         );
  AOI21_X1 U5567 ( .B1(n6363), .B2(n4510), .A(n4496), .ZN(n4497) );
  OAI211_X1 U5568 ( .C1(n4513), .C2(n5156), .A(n4498), .B(n4497), .ZN(U3145)
         );
  INV_X1 U5569 ( .A(DATAI_7_), .ZN(n4849) );
  NOR2_X1 U5570 ( .A1(n4849), .A2(n4515), .ZN(n6380) );
  INV_X1 U5571 ( .A(n6380), .ZN(n5161) );
  NAND2_X1 U5572 ( .A1(n4507), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4502)
         );
  NAND2_X1 U5573 ( .A1(n4508), .A2(n4499), .ZN(n5157) );
  INV_X1 U5574 ( .A(n5157), .ZN(n6378) );
  NAND2_X1 U5575 ( .A1(n2983), .A2(DATAI_23_), .ZN(n6271) );
  NAND2_X1 U5576 ( .A1(n2983), .A2(DATAI_31_), .ZN(n6385) );
  OAI22_X1 U5577 ( .A1(n6271), .A2(n4683), .B1(n4570), .B2(n6385), .ZN(n4500)
         );
  AOI21_X1 U5578 ( .B1(n6378), .B2(n4510), .A(n4500), .ZN(n4501) );
  OAI211_X1 U5579 ( .C1(n4513), .C2(n5161), .A(n4502), .B(n4501), .ZN(U3147)
         );
  INV_X1 U5580 ( .A(DATAI_6_), .ZN(n6549) );
  NOR2_X1 U5581 ( .A1(n6549), .A2(n4515), .ZN(n6371) );
  INV_X1 U5582 ( .A(n6371), .ZN(n5151) );
  NAND2_X1 U5583 ( .A1(n4507), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4506)
         );
  NAND2_X1 U5584 ( .A1(n4508), .A2(n4503), .ZN(n5147) );
  INV_X1 U5585 ( .A(n5147), .ZN(n6370) );
  NAND2_X1 U5586 ( .A1(n2983), .A2(DATAI_22_), .ZN(n6374) );
  NAND2_X1 U5587 ( .A1(n2983), .A2(DATAI_30_), .ZN(n6304) );
  OAI22_X1 U5588 ( .A1(n6374), .A2(n4683), .B1(n4570), .B2(n6304), .ZN(n4504)
         );
  AOI21_X1 U5589 ( .B1(n6370), .B2(n4510), .A(n4504), .ZN(n4505) );
  OAI211_X1 U5590 ( .C1(n4513), .C2(n5151), .A(n4506), .B(n4505), .ZN(U3146)
         );
  INV_X1 U5591 ( .A(DATAI_4_), .ZN(n6611) );
  NOR2_X1 U5592 ( .A1(n6611), .A2(n4515), .ZN(n6358) );
  INV_X1 U5593 ( .A(n6358), .ZN(n5171) );
  NAND2_X1 U5594 ( .A1(n4507), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4512)
         );
  NAND2_X1 U5595 ( .A1(n4508), .A2(n3112), .ZN(n5167) );
  INV_X1 U5596 ( .A(n5167), .ZN(n6357) );
  NAND2_X1 U5597 ( .A1(n2983), .A2(DATAI_20_), .ZN(n6259) );
  NAND2_X1 U5598 ( .A1(n2983), .A2(DATAI_28_), .ZN(n6361) );
  OAI22_X1 U5599 ( .A1(n6259), .A2(n4683), .B1(n4570), .B2(n6361), .ZN(n4509)
         );
  AOI21_X1 U5600 ( .B1(n6357), .B2(n4510), .A(n4509), .ZN(n4511) );
  OAI211_X1 U5601 ( .C1(n4513), .C2(n5171), .A(n4512), .B(n4511), .ZN(U3144)
         );
  OR2_X1 U5602 ( .A1(n5806), .A2(n4466), .ZN(n4652) );
  NOR2_X1 U5603 ( .A1(n5993), .A2(n4652), .ZN(n4517) );
  NOR2_X1 U5604 ( .A1(n4514), .A2(n6534), .ZN(n5134) );
  INV_X1 U5605 ( .A(n4654), .ZN(n5133) );
  NAND2_X1 U5606 ( .A1(n5133), .A2(n4653), .ZN(n4516) );
  INV_X1 U5607 ( .A(n4516), .ZN(n4592) );
  AOI22_X1 U5608 ( .A1(n4517), .A2(n6327), .B1(n5134), .B2(n4592), .ZN(n6312)
         );
  NAND3_X1 U5609 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5135), .A3(n6403), .ZN(n4625) );
  NOR2_X1 U5610 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4625), .ZN(n6315)
         );
  AND2_X1 U5611 ( .A1(n4514), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4899) );
  INV_X1 U5612 ( .A(n4899), .ZN(n6237) );
  AOI21_X1 U5613 ( .B1(n4516), .B2(STATE2_REG_2__SCAN_IN), .A(n4515), .ZN(
        n4595) );
  OAI211_X1 U5614 ( .C1(n6519), .C2(n6315), .A(n6237), .B(n4595), .ZN(n4520)
         );
  NAND2_X1 U5615 ( .A1(n6194), .A2(n5810), .ZN(n6329) );
  OR2_X1 U5616 ( .A1(n4472), .A2(n3386), .ZN(n4860) );
  OR2_X1 U5617 ( .A1(n6329), .A2(n4860), .ZN(n4521) );
  NAND2_X1 U5618 ( .A1(n5805), .A2(n4542), .ZN(n6234) );
  OR2_X1 U5619 ( .A1(n6234), .A2(n4902), .ZN(n6322) );
  NAND3_X1 U5620 ( .A1(n4521), .A2(n6327), .A3(n6322), .ZN(n4518) );
  AOI21_X1 U5621 ( .B1(n4518), .B2(n5815), .A(n4517), .ZN(n4519) );
  NAND2_X1 U5622 ( .A1(n6319), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4524) );
  INV_X1 U5623 ( .A(n6271), .ZN(n6375) );
  INV_X1 U5624 ( .A(n6315), .ZN(n4537) );
  OAI22_X1 U5625 ( .A1(n5157), .A2(n4537), .B1(n6385), .B2(n6322), .ZN(n4522)
         );
  AOI21_X1 U5626 ( .B1(n6375), .B2(n6317), .A(n4522), .ZN(n4523) );
  OAI211_X1 U5627 ( .C1(n6312), .C2(n5161), .A(n4524), .B(n4523), .ZN(U3091)
         );
  NAND2_X1 U5628 ( .A1(n6319), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4527) );
  INV_X1 U5629 ( .A(n6341), .ZN(n6273) );
  OAI22_X1 U5630 ( .A1(n5142), .A2(n4537), .B1(n6285), .B2(n6322), .ZN(n4525)
         );
  AOI21_X1 U5631 ( .B1(n6273), .B2(n6317), .A(n4525), .ZN(n4526) );
  OAI211_X1 U5632 ( .C1(n6312), .C2(n5146), .A(n4527), .B(n4526), .ZN(U3084)
         );
  NAND2_X1 U5633 ( .A1(n6319), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4530) );
  INV_X1 U5634 ( .A(n6347), .ZN(n6286) );
  OAI22_X1 U5635 ( .A1(n5179), .A2(n4537), .B1(n6289), .B2(n6322), .ZN(n4528)
         );
  AOI21_X1 U5636 ( .B1(n6286), .B2(n6317), .A(n4528), .ZN(n4529) );
  OAI211_X1 U5637 ( .C1(n6312), .C2(n5184), .A(n4530), .B(n4529), .ZN(U3085)
         );
  NAND2_X1 U5638 ( .A1(n6319), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4533) );
  INV_X1 U5639 ( .A(n6353), .ZN(n6290) );
  OAI22_X1 U5640 ( .A1(n5162), .A2(n4537), .B1(n6293), .B2(n6322), .ZN(n4531)
         );
  AOI21_X1 U5641 ( .B1(n6290), .B2(n6317), .A(n4531), .ZN(n4532) );
  OAI211_X1 U5642 ( .C1(n6312), .C2(n5166), .A(n4533), .B(n4532), .ZN(U3086)
         );
  NAND2_X1 U5643 ( .A1(n6319), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4536) );
  INV_X1 U5644 ( .A(n6259), .ZN(n6356) );
  OAI22_X1 U5645 ( .A1(n5167), .A2(n4537), .B1(n6361), .B2(n6322), .ZN(n4534)
         );
  AOI21_X1 U5646 ( .B1(n6356), .B2(n6317), .A(n4534), .ZN(n4535) );
  OAI211_X1 U5647 ( .C1(n6312), .C2(n5171), .A(n4536), .B(n4535), .ZN(U3088)
         );
  NAND2_X1 U5648 ( .A1(n6319), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4540) );
  INV_X1 U5649 ( .A(n6374), .ZN(n6301) );
  OAI22_X1 U5650 ( .A1(n5147), .A2(n4537), .B1(n6304), .B2(n6322), .ZN(n4538)
         );
  AOI21_X1 U5651 ( .B1(n6301), .B2(n6317), .A(n4538), .ZN(n4539) );
  OAI211_X1 U5652 ( .C1(n6312), .C2(n5151), .A(n4540), .B(n4539), .ZN(U3090)
         );
  NAND2_X1 U5653 ( .A1(n6240), .A2(n6327), .ZN(n6238) );
  INV_X1 U5654 ( .A(n6238), .ZN(n4541) );
  NOR2_X1 U5655 ( .A1(n5133), .A2(n6409), .ZN(n4803) );
  AOI22_X1 U5656 ( .A1(n4541), .A2(n4415), .B1(n4899), .B2(n4803), .ZN(n4577)
         );
  INV_X1 U5657 ( .A(n6361), .ZN(n6256) );
  NOR2_X1 U5658 ( .A1(n4472), .A2(n4542), .ZN(n4543) );
  NAND2_X1 U5659 ( .A1(n5805), .A2(n4543), .ZN(n4593) );
  INV_X1 U5660 ( .A(n4593), .ZN(n4758) );
  NAND2_X1 U5661 ( .A1(n4758), .A2(n3386), .ZN(n4796) );
  INV_X1 U5662 ( .A(n4796), .ZN(n4573) );
  NAND2_X1 U5663 ( .A1(n6398), .A2(n4544), .ZN(n4571) );
  OAI22_X1 U5664 ( .A1(n5167), .A2(n4571), .B1(n6259), .B2(n4570), .ZN(n4545)
         );
  AOI21_X1 U5665 ( .B1(n6256), .B2(n4573), .A(n4545), .ZN(n4551) );
  AOI21_X1 U5666 ( .B1(n4796), .B2(n4570), .A(n6604), .ZN(n4549) );
  INV_X1 U5667 ( .A(n6240), .ZN(n4546) );
  NAND2_X1 U5668 ( .A1(n6327), .A2(n4546), .ZN(n4548) );
  OAI21_X1 U5669 ( .B1(n4654), .B2(n6534), .A(n4658), .ZN(n4804) );
  NOR2_X1 U5670 ( .A1(n5134), .A2(n4804), .ZN(n6245) );
  AOI21_X1 U5671 ( .B1(n4571), .B2(STATE2_REG_3__SCAN_IN), .A(n6409), .ZN(
        n4547) );
  OAI211_X1 U5672 ( .C1(n4549), .C2(n4548), .A(n6245), .B(n4547), .ZN(n4574)
         );
  NAND2_X1 U5673 ( .A1(n4574), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4550)
         );
  OAI211_X1 U5674 ( .C1(n5171), .C2(n4577), .A(n4551), .B(n4550), .ZN(U3136)
         );
  INV_X1 U5675 ( .A(n6304), .ZN(n6368) );
  OAI22_X1 U5676 ( .A1(n5147), .A2(n4571), .B1(n6374), .B2(n4570), .ZN(n4552)
         );
  AOI21_X1 U5677 ( .B1(n6368), .B2(n4573), .A(n4552), .ZN(n4554) );
  NAND2_X1 U5678 ( .A1(n4574), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4553)
         );
  OAI211_X1 U5679 ( .C1(n5151), .C2(n4577), .A(n4554), .B(n4553), .ZN(U3138)
         );
  INV_X1 U5680 ( .A(n6323), .ZN(n6362) );
  OAI22_X1 U5681 ( .A1(n5152), .A2(n4571), .B1(n6367), .B2(n4570), .ZN(n4555)
         );
  AOI21_X1 U5682 ( .B1(n6362), .B2(n4573), .A(n4555), .ZN(n4557) );
  NAND2_X1 U5683 ( .A1(n4574), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4556)
         );
  OAI211_X1 U5684 ( .C1(n5156), .C2(n4577), .A(n4557), .B(n4556), .ZN(U3137)
         );
  INV_X1 U5685 ( .A(n6285), .ZN(n6325) );
  OAI22_X1 U5686 ( .A1(n5142), .A2(n4571), .B1(n6341), .B2(n4570), .ZN(n4558)
         );
  AOI21_X1 U5687 ( .B1(n6325), .B2(n4573), .A(n4558), .ZN(n4560) );
  NAND2_X1 U5688 ( .A1(n4574), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4559)
         );
  OAI211_X1 U5689 ( .C1(n5146), .C2(n4577), .A(n4560), .B(n4559), .ZN(U3132)
         );
  INV_X1 U5690 ( .A(n6385), .ZN(n6267) );
  OAI22_X1 U5691 ( .A1(n5157), .A2(n4571), .B1(n6271), .B2(n4570), .ZN(n4561)
         );
  AOI21_X1 U5692 ( .B1(n6267), .B2(n4573), .A(n4561), .ZN(n4563) );
  NAND2_X1 U5693 ( .A1(n4574), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4562)
         );
  OAI211_X1 U5694 ( .C1(n5161), .C2(n4577), .A(n4563), .B(n4562), .ZN(U3139)
         );
  INV_X1 U5695 ( .A(n6293), .ZN(n6348) );
  OAI22_X1 U5696 ( .A1(n5162), .A2(n4571), .B1(n6353), .B2(n4570), .ZN(n4564)
         );
  AOI21_X1 U5697 ( .B1(n6348), .B2(n4573), .A(n4564), .ZN(n4566) );
  NAND2_X1 U5698 ( .A1(n4574), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4565)
         );
  OAI211_X1 U5699 ( .C1(n5166), .C2(n4577), .A(n4566), .B(n4565), .ZN(U3134)
         );
  INV_X1 U5700 ( .A(n6289), .ZN(n6342) );
  OAI22_X1 U5701 ( .A1(n5179), .A2(n4571), .B1(n6347), .B2(n4570), .ZN(n4567)
         );
  AOI21_X1 U5702 ( .B1(n6342), .B2(n4573), .A(n4567), .ZN(n4569) );
  NAND2_X1 U5703 ( .A1(n4574), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4568)
         );
  OAI211_X1 U5704 ( .C1(n5184), .C2(n4577), .A(n4569), .B(n4568), .ZN(U3133)
         );
  INV_X1 U5705 ( .A(n6397), .ZN(n6252) );
  OAI22_X1 U5706 ( .A1(n5172), .A2(n4571), .B1(n6255), .B2(n4570), .ZN(n4572)
         );
  AOI21_X1 U5707 ( .B1(n6252), .B2(n4573), .A(n4572), .ZN(n4576) );
  NAND2_X1 U5708 ( .A1(n4574), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4575)
         );
  OAI211_X1 U5709 ( .C1(n5176), .C2(n4577), .A(n4576), .B(n4575), .ZN(U3135)
         );
  INV_X1 U5710 ( .A(n4587), .ZN(n4579) );
  AOI21_X1 U5711 ( .B1(n4581), .B2(n4580), .A(n4579), .ZN(n4965) );
  INV_X1 U5712 ( .A(n4965), .ZN(n4739) );
  OAI21_X1 U5713 ( .B1(n4583), .B2(n4461), .A(n4582), .ZN(n6161) );
  INV_X1 U5714 ( .A(n6161), .ZN(n4584) );
  AOI22_X1 U5715 ( .A1(n6005), .A2(n4584), .B1(n5551), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4585) );
  OAI21_X1 U5716 ( .B1(n4739), .B2(n5348), .A(n4585), .ZN(U2855) );
  OAI222_X1 U5717 ( .A1(n4739), .A2(n5583), .B1(n5582), .B2(n6611), .C1(n5581), 
        .C2(n6040), .ZN(U2887) );
  CLKBUF_X1 U5718 ( .A(n4586), .Z(n4649) );
  AOI21_X1 U5719 ( .B1(n4588), .B2(n4587), .A(n4649), .ZN(n4939) );
  INV_X1 U5720 ( .A(n4939), .ZN(n4723) );
  AOI21_X1 U5721 ( .B1(n4590), .B2(n4582), .A(n4589), .ZN(n6150) );
  AOI22_X1 U5722 ( .A1(n6005), .A2(n6150), .B1(n5551), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4591) );
  OAI21_X1 U5723 ( .B1(n4723), .B2(n5348), .A(n4591), .ZN(U2854) );
  OAI222_X1 U5724 ( .A1(n4723), .A2(n5583), .B1(n5582), .B2(n6674), .C1(n5581), 
        .C2(n3789), .ZN(U2886) );
  INV_X1 U5725 ( .A(n4466), .ZN(n5824) );
  NAND2_X1 U5726 ( .A1(n5806), .A2(n5824), .ZN(n4854) );
  NOR2_X1 U5727 ( .A1(n4854), .A2(n6332), .ZN(n4900) );
  AOI22_X1 U5728 ( .A1(n4900), .A2(n4415), .B1(n4592), .B2(n4899), .ZN(n6386)
         );
  INV_X1 U5729 ( .A(n4854), .ZN(n4756) );
  OR2_X1 U5730 ( .A1(n6329), .A2(n4902), .ZN(n6396) );
  OR2_X1 U5731 ( .A1(n4593), .A2(n3386), .ZN(n4765) );
  AOI21_X1 U5732 ( .B1(n6396), .B2(n4765), .A(n6604), .ZN(n4594) );
  AOI211_X1 U5733 ( .C1(n4756), .C2(n4853), .A(n6332), .B(n4594), .ZN(n4598)
         );
  NAND2_X1 U5734 ( .A1(n6403), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4855) );
  NOR2_X1 U5735 ( .A1(n6409), .A2(n4855), .ZN(n4755) );
  AND2_X1 U5736 ( .A1(n6398), .A2(n4755), .ZN(n6387) );
  INV_X1 U5737 ( .A(n5134), .ZN(n4596) );
  OAI211_X1 U5738 ( .C1(n6519), .C2(n6387), .A(n4596), .B(n4595), .ZN(n4597)
         );
  NAND2_X1 U5739 ( .A1(n6393), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4601)
         );
  INV_X1 U5740 ( .A(n6387), .ZN(n4617) );
  OAI22_X1 U5741 ( .A1(n5152), .A2(n4617), .B1(n6367), .B2(n4765), .ZN(n4599)
         );
  AOI21_X1 U5742 ( .B1(n6362), .B2(n6376), .A(n4599), .ZN(n4600) );
  OAI211_X1 U5743 ( .C1(n6386), .C2(n5156), .A(n4601), .B(n4600), .ZN(U3121)
         );
  NAND2_X1 U5744 ( .A1(n6393), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4604)
         );
  OAI22_X1 U5745 ( .A1(n5157), .A2(n4617), .B1(n6271), .B2(n4765), .ZN(n4602)
         );
  AOI21_X1 U5746 ( .B1(n6267), .B2(n6376), .A(n4602), .ZN(n4603) );
  OAI211_X1 U5747 ( .C1(n6386), .C2(n5161), .A(n4604), .B(n4603), .ZN(U3123)
         );
  NAND2_X1 U5748 ( .A1(n6393), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4607)
         );
  OAI22_X1 U5749 ( .A1(n5147), .A2(n4617), .B1(n6374), .B2(n4765), .ZN(n4605)
         );
  AOI21_X1 U5750 ( .B1(n6368), .B2(n6376), .A(n4605), .ZN(n4606) );
  OAI211_X1 U5751 ( .C1(n6386), .C2(n5151), .A(n4607), .B(n4606), .ZN(U3122)
         );
  NAND2_X1 U5752 ( .A1(n6393), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4610)
         );
  OAI22_X1 U5753 ( .A1(n5167), .A2(n4617), .B1(n6259), .B2(n4765), .ZN(n4608)
         );
  AOI21_X1 U5754 ( .B1(n6256), .B2(n6376), .A(n4608), .ZN(n4609) );
  OAI211_X1 U5755 ( .C1(n6386), .C2(n5171), .A(n4610), .B(n4609), .ZN(U3120)
         );
  NAND2_X1 U5756 ( .A1(n6393), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4613)
         );
  OAI22_X1 U5757 ( .A1(n5179), .A2(n4617), .B1(n6347), .B2(n4765), .ZN(n4611)
         );
  AOI21_X1 U5758 ( .B1(n6342), .B2(n6376), .A(n4611), .ZN(n4612) );
  OAI211_X1 U5759 ( .C1(n6386), .C2(n5184), .A(n4613), .B(n4612), .ZN(U3117)
         );
  NAND2_X1 U5760 ( .A1(n6393), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4616)
         );
  OAI22_X1 U5761 ( .A1(n5142), .A2(n4617), .B1(n6341), .B2(n4765), .ZN(n4614)
         );
  AOI21_X1 U5762 ( .B1(n6325), .B2(n6376), .A(n4614), .ZN(n4615) );
  OAI211_X1 U5763 ( .C1(n6386), .C2(n5146), .A(n4616), .B(n4615), .ZN(U3116)
         );
  NAND2_X1 U5764 ( .A1(n6393), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4620)
         );
  OAI22_X1 U5765 ( .A1(n5162), .A2(n4617), .B1(n6353), .B2(n4765), .ZN(n4618)
         );
  AOI21_X1 U5766 ( .B1(n6348), .B2(n6376), .A(n4618), .ZN(n4619) );
  OAI211_X1 U5767 ( .C1(n6386), .C2(n5166), .A(n4620), .B(n4619), .ZN(U3118)
         );
  OR2_X1 U5768 ( .A1(n4472), .A2(n5046), .ZN(n4859) );
  OR2_X1 U5769 ( .A1(n4472), .A2(n6604), .ZN(n4851) );
  OR2_X1 U5770 ( .A1(n6329), .A2(n4851), .ZN(n4621) );
  AND2_X1 U5771 ( .A1(n4621), .A2(n6327), .ZN(n4624) );
  INV_X1 U5772 ( .A(n4652), .ZN(n4622) );
  NOR2_X1 U5773 ( .A1(n6398), .A2(n4625), .ZN(n4644) );
  AOI21_X1 U5774 ( .B1(n4757), .B2(n4622), .A(n4644), .ZN(n4627) );
  AOI22_X1 U5775 ( .A1(n4624), .A2(n4627), .B1(n6332), .B2(n4625), .ZN(n4623)
         );
  NAND2_X1 U5776 ( .A1(n6278), .A2(n4623), .ZN(n4643) );
  INV_X1 U5777 ( .A(n4624), .ZN(n4626) );
  OAI22_X1 U5778 ( .A1(n4627), .A2(n4626), .B1(n6534), .B2(n4625), .ZN(n4642)
         );
  AOI22_X1 U5779 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4643), .B1(n6390), 
        .B2(n4642), .ZN(n4629) );
  AOI22_X1 U5780 ( .A1(n6388), .A2(n4644), .B1(n6317), .B2(n6252), .ZN(n4628)
         );
  OAI211_X1 U5781 ( .C1(n4830), .C2(n6255), .A(n4629), .B(n4628), .ZN(U3095)
         );
  AOI22_X1 U5782 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4643), .B1(n6364), 
        .B2(n4642), .ZN(n4631) );
  AOI22_X1 U5783 ( .A1(n6363), .A2(n4644), .B1(n6317), .B2(n6362), .ZN(n4630)
         );
  OAI211_X1 U5784 ( .C1(n4830), .C2(n6367), .A(n4631), .B(n4630), .ZN(U3097)
         );
  AOI22_X1 U5785 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4643), .B1(n6358), 
        .B2(n4642), .ZN(n4633) );
  AOI22_X1 U5786 ( .A1(n6357), .A2(n4644), .B1(n6317), .B2(n6256), .ZN(n4632)
         );
  OAI211_X1 U5787 ( .C1(n4830), .C2(n6259), .A(n4633), .B(n4632), .ZN(U3096)
         );
  AOI22_X1 U5788 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4643), .B1(n6338), 
        .B2(n4642), .ZN(n4635) );
  AOI22_X1 U5789 ( .A1(n6326), .A2(n4644), .B1(n6317), .B2(n6325), .ZN(n4634)
         );
  OAI211_X1 U5790 ( .C1(n4830), .C2(n6341), .A(n4635), .B(n4634), .ZN(U3092)
         );
  AOI22_X1 U5791 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4643), .B1(n6371), 
        .B2(n4642), .ZN(n4637) );
  AOI22_X1 U5792 ( .A1(n6370), .A2(n4644), .B1(n6317), .B2(n6368), .ZN(n4636)
         );
  OAI211_X1 U5793 ( .C1(n4830), .C2(n6374), .A(n4637), .B(n4636), .ZN(U3098)
         );
  AOI22_X1 U5794 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4643), .B1(n6350), 
        .B2(n4642), .ZN(n4639) );
  AOI22_X1 U5795 ( .A1(n6349), .A2(n4644), .B1(n6317), .B2(n6348), .ZN(n4638)
         );
  OAI211_X1 U5796 ( .C1(n4830), .C2(n6353), .A(n4639), .B(n4638), .ZN(U3094)
         );
  AOI22_X1 U5797 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4643), .B1(n6344), 
        .B2(n4642), .ZN(n4641) );
  AOI22_X1 U5798 ( .A1(n6343), .A2(n4644), .B1(n6317), .B2(n6342), .ZN(n4640)
         );
  OAI211_X1 U5799 ( .C1(n4830), .C2(n6347), .A(n4641), .B(n4640), .ZN(U3093)
         );
  AOI22_X1 U5800 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4643), .B1(n6380), 
        .B2(n4642), .ZN(n4646) );
  AOI22_X1 U5801 ( .A1(n6378), .A2(n4644), .B1(n6317), .B2(n6267), .ZN(n4645)
         );
  OAI211_X1 U5802 ( .C1(n4830), .C2(n6271), .A(n4646), .B(n4645), .ZN(U3099)
         );
  OAI21_X1 U5803 ( .B1(n4649), .B2(n4648), .A(n4836), .ZN(n5982) );
  OAI222_X1 U5804 ( .A1(n5982), .A2(n5583), .B1(n5582), .B2(n6549), .C1(n5581), 
        .C2(n6036), .ZN(U2885) );
  OAI21_X1 U5805 ( .B1(n4651), .B2(n4589), .A(n4650), .ZN(n6138) );
  INV_X1 U5806 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5973) );
  OAI222_X1 U5807 ( .A1(n6138), .A2(n5549), .B1(n5973), .B2(n6009), .C1(n5982), 
        .C2(n5553), .ZN(U2853) );
  NOR2_X1 U5808 ( .A1(n4415), .A2(n4652), .ZN(n5039) );
  NOR2_X1 U5809 ( .A1(n4654), .A2(n4653), .ZN(n4898) );
  AOI22_X1 U5810 ( .A1(n5039), .A2(n6327), .B1(n5134), .B2(n4898), .ZN(n4689)
         );
  INV_X1 U5811 ( .A(n4683), .ZN(n4655) );
  NOR2_X1 U5812 ( .A1(n4655), .A2(n6332), .ZN(n4657) );
  OR3_X1 U5813 ( .A1(n5810), .A2(n5805), .A3(n4472), .ZN(n5047) );
  INV_X1 U5814 ( .A(n5047), .ZN(n5040) );
  NAND2_X1 U5815 ( .A1(n5040), .A2(n5046), .ZN(n5067) );
  INV_X1 U5816 ( .A(n5815), .ZN(n4656) );
  AOI21_X1 U5817 ( .B1(n4657), .B2(n5067), .A(n4656), .ZN(n4660) );
  NAND3_X1 U5818 ( .A1(n6409), .A2(n5135), .A3(n6403), .ZN(n5043) );
  OR2_X1 U5819 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5043), .ZN(n4684)
         );
  OAI21_X1 U5820 ( .B1(n4898), .B2(n6534), .A(n4658), .ZN(n4906) );
  AOI211_X1 U5821 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4684), .A(n4899), .B(
        n4906), .ZN(n4659) );
  OAI21_X1 U5822 ( .B1(n5039), .B2(n4660), .A(n4659), .ZN(n4682) );
  NAND2_X1 U5823 ( .A1(n4682), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4663) );
  INV_X1 U5824 ( .A(n5067), .ZN(n4686) );
  OAI22_X1 U5825 ( .A1(n5147), .A2(n4684), .B1(n6304), .B2(n4683), .ZN(n4661)
         );
  AOI21_X1 U5826 ( .B1(n6301), .B2(n4686), .A(n4661), .ZN(n4662) );
  OAI211_X1 U5827 ( .C1(n4689), .C2(n5151), .A(n4663), .B(n4662), .ZN(U3026)
         );
  NAND2_X1 U5828 ( .A1(n4682), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4666) );
  OAI22_X1 U5829 ( .A1(n5162), .A2(n4684), .B1(n6293), .B2(n4683), .ZN(n4664)
         );
  AOI21_X1 U5830 ( .B1(n6290), .B2(n4686), .A(n4664), .ZN(n4665) );
  OAI211_X1 U5831 ( .C1(n4689), .C2(n5166), .A(n4666), .B(n4665), .ZN(U3022)
         );
  NAND2_X1 U5832 ( .A1(n4682), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4669) );
  OAI22_X1 U5833 ( .A1(n5167), .A2(n4684), .B1(n6361), .B2(n4683), .ZN(n4667)
         );
  AOI21_X1 U5834 ( .B1(n6356), .B2(n4686), .A(n4667), .ZN(n4668) );
  OAI211_X1 U5835 ( .C1(n4689), .C2(n5171), .A(n4669), .B(n4668), .ZN(U3024)
         );
  NAND2_X1 U5836 ( .A1(n4682), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4672) );
  INV_X1 U5837 ( .A(n6255), .ZN(n6392) );
  OAI22_X1 U5838 ( .A1(n5172), .A2(n4684), .B1(n6397), .B2(n4683), .ZN(n4670)
         );
  AOI21_X1 U5839 ( .B1(n6392), .B2(n4686), .A(n4670), .ZN(n4671) );
  OAI211_X1 U5840 ( .C1(n4689), .C2(n5176), .A(n4672), .B(n4671), .ZN(U3023)
         );
  NAND2_X1 U5841 ( .A1(n4682), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4675) );
  OAI22_X1 U5842 ( .A1(n5142), .A2(n4684), .B1(n6285), .B2(n4683), .ZN(n4673)
         );
  AOI21_X1 U5843 ( .B1(n6273), .B2(n4686), .A(n4673), .ZN(n4674) );
  OAI211_X1 U5844 ( .C1(n4689), .C2(n5146), .A(n4675), .B(n4674), .ZN(U3020)
         );
  NAND2_X1 U5845 ( .A1(n4682), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4678) );
  OAI22_X1 U5846 ( .A1(n5157), .A2(n4684), .B1(n6385), .B2(n4683), .ZN(n4676)
         );
  AOI21_X1 U5847 ( .B1(n6375), .B2(n4686), .A(n4676), .ZN(n4677) );
  OAI211_X1 U5848 ( .C1(n4689), .C2(n5161), .A(n4678), .B(n4677), .ZN(U3027)
         );
  NAND2_X1 U5849 ( .A1(n4682), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4681) );
  INV_X1 U5850 ( .A(n6367), .ZN(n6318) );
  OAI22_X1 U5851 ( .A1(n5152), .A2(n4684), .B1(n6323), .B2(n4683), .ZN(n4679)
         );
  AOI21_X1 U5852 ( .B1(n6318), .B2(n4686), .A(n4679), .ZN(n4680) );
  OAI211_X1 U5853 ( .C1(n4689), .C2(n5156), .A(n4681), .B(n4680), .ZN(U3025)
         );
  NAND2_X1 U5854 ( .A1(n4682), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4688) );
  OAI22_X1 U5855 ( .A1(n5179), .A2(n4684), .B1(n6289), .B2(n4683), .ZN(n4685)
         );
  AOI21_X1 U5856 ( .B1(n6286), .B2(n4686), .A(n4685), .ZN(n4687) );
  OAI211_X1 U5857 ( .C1(n4689), .C2(n5184), .A(n4688), .B(n4687), .ZN(U3021)
         );
  NOR3_X1 U5858 ( .A1(n6536), .A2(n6519), .A3(n6535), .ZN(n6431) );
  INV_X1 U5859 ( .A(n6431), .ZN(n4693) );
  NAND2_X1 U5860 ( .A1(n6536), .A2(n6534), .ZN(n6444) );
  NOR3_X1 U5861 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6444), .A3(n5340), .ZN(
        n6440) );
  INV_X1 U5862 ( .A(n6440), .ZN(n4692) );
  NAND2_X1 U5863 ( .A1(n4693), .A2(n4692), .ZN(n4694) );
  INV_X1 U5864 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5263) );
  INV_X1 U5865 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4697) );
  XNOR2_X1 U5866 ( .A(n4698), .B(n4697), .ZN(n5365) );
  NOR2_X1 U5867 ( .A1(n5365), .A2(n5340), .ZN(n4699) );
  OR2_X1 U5868 ( .A1(n3510), .A2(n4724), .ZN(n4700) );
  INV_X1 U5869 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U5870 ( .A1(n6638), .A2(n6604), .ZN(n4712) );
  NOR2_X1 U5871 ( .A1(n4724), .A2(n4712), .ZN(n4701) );
  AND2_X1 U5872 ( .A1(n3602), .A2(n4701), .ZN(n4702) );
  INV_X1 U5873 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6158) );
  NAND3_X1 U5874 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5990) );
  NOR2_X1 U5875 ( .A1(n6158), .A2(n5990), .ZN(n4704) );
  NAND2_X1 U5876 ( .A1(n5991), .A2(n4704), .ZN(n4841) );
  NAND2_X1 U5877 ( .A1(n4950), .A2(n5327), .ZN(n5835) );
  INV_X1 U5878 ( .A(n5835), .ZN(n5483) );
  AND3_X1 U5879 ( .A1(n4950), .A2(REIP_REG_5__SCAN_IN), .A3(n4704), .ZN(n5216)
         );
  NOR2_X1 U5880 ( .A1(n5483), .A2(n5216), .ZN(n5980) );
  INV_X1 U5881 ( .A(n5980), .ZN(n4705) );
  AOI21_X1 U5882 ( .B1(n6470), .B2(n4841), .A(n4705), .ZN(n4706) );
  INV_X1 U5883 ( .A(n4706), .ZN(n4722) );
  AND2_X1 U5884 ( .A1(n5365), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4707) );
  INV_X1 U5885 ( .A(n4937), .ZN(n4720) );
  INV_X1 U5886 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4718) );
  AND3_X1 U5887 ( .A1(EBX_REG_31__SCAN_IN), .A2(n6538), .A3(n4712), .ZN(n4708)
         );
  NAND2_X1 U5888 ( .A1(n3022), .A2(n4708), .ZN(n5938) );
  NOR2_X1 U5889 ( .A1(n4710), .A2(n4712), .ZN(n6429) );
  INV_X1 U5890 ( .A(n6429), .ZN(n4711) );
  AND2_X1 U5891 ( .A1(n3359), .A2(n4711), .ZN(n5328) );
  INV_X1 U5892 ( .A(n4712), .ZN(n4713) );
  NOR2_X1 U5893 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4713), .ZN(n4714) );
  AND2_X1 U5894 ( .A1(n3602), .A2(n4714), .ZN(n4715) );
  OR2_X1 U5895 ( .A1(n5328), .A2(n4715), .ZN(n4716) );
  AND2_X1 U5896 ( .A1(n4716), .A2(n6538), .ZN(n5986) );
  AOI22_X1 U5897 ( .A1(n5987), .A2(n6150), .B1(n5986), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4717) );
  OAI211_X1 U5898 ( .C1(n5997), .C2(n4718), .A(n4717), .B(n6159), .ZN(n4719)
         );
  AOI21_X1 U5899 ( .B1(n5968), .B2(n4720), .A(n4719), .ZN(n4721) );
  OAI211_X1 U5900 ( .C1(n5989), .C2(n4723), .A(n4722), .B(n4721), .ZN(U2822)
         );
  OAI21_X1 U5901 ( .B1(n5956), .B2(n5968), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4730) );
  NOR2_X1 U5902 ( .A1(n5392), .A2(n4724), .ZN(n4952) );
  INV_X1 U5903 ( .A(n4952), .ZN(n5992) );
  NOR2_X1 U5904 ( .A1(n4857), .A2(n5992), .ZN(n4728) );
  OAI22_X1 U5905 ( .A1(n4726), .A2(n5938), .B1(n4725), .B2(n5974), .ZN(n4727)
         );
  AOI211_X1 U5906 ( .C1(n5835), .C2(REIP_REG_0__SCAN_IN), .A(n4728), .B(n4727), 
        .ZN(n4729) );
  OAI211_X1 U5907 ( .C1(n5989), .C2(n4731), .A(n4730), .B(n4729), .ZN(U2827)
         );
  NOR3_X1 U5908 ( .A1(n5327), .A2(REIP_REG_4__SCAN_IN), .A3(n5990), .ZN(n4733)
         );
  OAI21_X1 U5909 ( .B1(n4993), .B2(n5990), .A(n5835), .ZN(n6004) );
  INV_X1 U5910 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4966) );
  OAI22_X1 U5911 ( .A1(n6004), .A2(n6158), .B1(n4966), .B2(n5997), .ZN(n4732)
         );
  NOR3_X1 U5912 ( .A1(n4733), .A2(n6185), .A3(n4732), .ZN(n4735) );
  NAND2_X1 U5913 ( .A1(n5986), .A2(EBX_REG_4__SCAN_IN), .ZN(n4734) );
  OAI211_X1 U5914 ( .C1(n6161), .C2(n5938), .A(n4735), .B(n4734), .ZN(n4736)
         );
  AOI21_X1 U5915 ( .B1(n5968), .B2(n4968), .A(n4736), .ZN(n4738) );
  NAND2_X1 U5916 ( .A1(n5904), .A2(n4952), .ZN(n4737) );
  OAI211_X1 U5917 ( .C1(n4739), .C2(n5989), .A(n4738), .B(n4737), .ZN(U2823)
         );
  NAND2_X1 U5918 ( .A1(n4740), .A2(n6399), .ZN(n4741) );
  NAND2_X1 U5919 ( .A1(n4355), .A2(n4741), .ZN(n4742) );
  NAND2_X1 U5920 ( .A1(n6017), .A2(n3602), .ZN(n5101) );
  NOR2_X1 U5921 ( .A1(n4743), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6540) );
  AOI22_X1 U5922 ( .A1(n6540), .A2(UWORD_REG_14__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4744) );
  OAI21_X1 U5923 ( .B1(n4745), .B2(n5101), .A(n4744), .ZN(U2893) );
  AOI22_X1 U5924 ( .A1(n6540), .A2(UWORD_REG_10__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4746) );
  OAI21_X1 U5925 ( .B1(n4151), .B2(n5101), .A(n4746), .ZN(U2897) );
  AOI22_X1 U5926 ( .A1(n6540), .A2(UWORD_REG_11__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4747) );
  OAI21_X1 U5927 ( .B1(n4748), .B2(n5101), .A(n4747), .ZN(U2896) );
  AOI22_X1 U5928 ( .A1(n6540), .A2(UWORD_REG_12__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4749) );
  OAI21_X1 U5929 ( .B1(n4174), .B2(n5101), .A(n4749), .ZN(U2895) );
  AOI22_X1 U5930 ( .A1(n6540), .A2(UWORD_REG_13__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4750) );
  OAI21_X1 U5931 ( .B1(n4751), .B2(n5101), .A(n4750), .ZN(U2894) );
  AOI22_X1 U5932 ( .A1(n6540), .A2(UWORD_REG_8__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4752) );
  OAI21_X1 U5933 ( .B1(n4096), .B2(n5101), .A(n4752), .ZN(U2899) );
  AOI22_X1 U5934 ( .A1(n6540), .A2(UWORD_REG_9__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4753) );
  OAI21_X1 U5935 ( .B1(n4754), .B2(n5101), .A(n4753), .ZN(U2898) );
  INV_X1 U5936 ( .A(n4755), .ZN(n4762) );
  AND2_X1 U5937 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4755), .ZN(n4794)
         );
  AOI21_X1 U5938 ( .B1(n4757), .B2(n4756), .A(n4794), .ZN(n4764) );
  NAND2_X1 U5939 ( .A1(n4758), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5811) );
  NAND2_X1 U5940 ( .A1(n4764), .A2(n5811), .ZN(n4759) );
  NOR2_X1 U5941 ( .A1(n6332), .A2(n4759), .ZN(n4761) );
  INV_X1 U5942 ( .A(n6278), .ZN(n4760) );
  AOI211_X2 U5943 ( .C1(n6332), .C2(n4762), .A(n4761), .B(n4760), .ZN(n4801)
         );
  INV_X1 U5944 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4769) );
  NAND2_X1 U5945 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4763) );
  OAI22_X1 U5946 ( .A1(n4764), .A2(n6332), .B1(n4763), .B2(n4855), .ZN(n4798)
         );
  INV_X1 U5947 ( .A(n4765), .ZN(n6391) );
  AOI22_X1 U5948 ( .A1(n6343), .A2(n4794), .B1(n6342), .B2(n6391), .ZN(n4766)
         );
  OAI21_X1 U5949 ( .B1(n6347), .B2(n4796), .A(n4766), .ZN(n4767) );
  AOI21_X1 U5950 ( .B1(n6344), .B2(n4798), .A(n4767), .ZN(n4768) );
  OAI21_X1 U5951 ( .B1(n4801), .B2(n4769), .A(n4768), .ZN(U3125) );
  INV_X1 U5952 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4773) );
  AOI22_X1 U5953 ( .A1(n6378), .A2(n4794), .B1(n6267), .B2(n6391), .ZN(n4770)
         );
  OAI21_X1 U5954 ( .B1(n6271), .B2(n4796), .A(n4770), .ZN(n4771) );
  AOI21_X1 U5955 ( .B1(n6380), .B2(n4798), .A(n4771), .ZN(n4772) );
  OAI21_X1 U5956 ( .B1(n4801), .B2(n4773), .A(n4772), .ZN(U3131) );
  INV_X1 U5957 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4777) );
  AOI22_X1 U5958 ( .A1(n6363), .A2(n4794), .B1(n6362), .B2(n6391), .ZN(n4774)
         );
  OAI21_X1 U5959 ( .B1(n6367), .B2(n4796), .A(n4774), .ZN(n4775) );
  AOI21_X1 U5960 ( .B1(n6364), .B2(n4798), .A(n4775), .ZN(n4776) );
  OAI21_X1 U5961 ( .B1(n4801), .B2(n4777), .A(n4776), .ZN(U3129) );
  INV_X1 U5962 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4781) );
  AOI22_X1 U5963 ( .A1(n6349), .A2(n4794), .B1(n6348), .B2(n6391), .ZN(n4778)
         );
  OAI21_X1 U5964 ( .B1(n6353), .B2(n4796), .A(n4778), .ZN(n4779) );
  AOI21_X1 U5965 ( .B1(n6350), .B2(n4798), .A(n4779), .ZN(n4780) );
  OAI21_X1 U5966 ( .B1(n4801), .B2(n4781), .A(n4780), .ZN(U3126) );
  INV_X1 U5967 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4785) );
  AOI22_X1 U5968 ( .A1(n6388), .A2(n4794), .B1(n6252), .B2(n6391), .ZN(n4782)
         );
  OAI21_X1 U5969 ( .B1(n6255), .B2(n4796), .A(n4782), .ZN(n4783) );
  AOI21_X1 U5970 ( .B1(n6390), .B2(n4798), .A(n4783), .ZN(n4784) );
  OAI21_X1 U5971 ( .B1(n4801), .B2(n4785), .A(n4784), .ZN(U3127) );
  INV_X1 U5972 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4789) );
  AOI22_X1 U5973 ( .A1(n6326), .A2(n4794), .B1(n6325), .B2(n6391), .ZN(n4786)
         );
  OAI21_X1 U5974 ( .B1(n6341), .B2(n4796), .A(n4786), .ZN(n4787) );
  AOI21_X1 U5975 ( .B1(n6338), .B2(n4798), .A(n4787), .ZN(n4788) );
  OAI21_X1 U5976 ( .B1(n4801), .B2(n4789), .A(n4788), .ZN(U3124) );
  INV_X1 U5977 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4793) );
  AOI22_X1 U5978 ( .A1(n6370), .A2(n4794), .B1(n6368), .B2(n6391), .ZN(n4790)
         );
  OAI21_X1 U5979 ( .B1(n6374), .B2(n4796), .A(n4790), .ZN(n4791) );
  AOI21_X1 U5980 ( .B1(n6371), .B2(n4798), .A(n4791), .ZN(n4792) );
  OAI21_X1 U5981 ( .B1(n4801), .B2(n4793), .A(n4792), .ZN(U3130) );
  INV_X1 U5982 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4800) );
  AOI22_X1 U5983 ( .A1(n6357), .A2(n4794), .B1(n6256), .B2(n6391), .ZN(n4795)
         );
  OAI21_X1 U5984 ( .B1(n6259), .B2(n4796), .A(n4795), .ZN(n4797) );
  AOI21_X1 U5985 ( .B1(n6358), .B2(n4798), .A(n4797), .ZN(n4799) );
  OAI21_X1 U5986 ( .B1(n4801), .B2(n4800), .A(n4799), .ZN(U3128) );
  OR2_X1 U5987 ( .A1(n6329), .A2(n6233), .ZN(n6384) );
  NAND2_X1 U5988 ( .A1(n6384), .A2(n4830), .ZN(n4802) );
  AOI21_X1 U5989 ( .B1(n4802), .B2(STATEBS16_REG_SCAN_IN), .A(n6332), .ZN(
        n4806) );
  NOR2_X1 U5990 ( .A1(n5806), .A2(n5824), .ZN(n5132) );
  AND2_X1 U5991 ( .A1(n5132), .A2(n4415), .ZN(n6331) );
  AOI22_X1 U5992 ( .A1(n4806), .A2(n6331), .B1(n5134), .B2(n4803), .ZN(n4835)
         );
  NOR2_X1 U5993 ( .A1(n4899), .A2(n4804), .ZN(n5139) );
  INV_X1 U5994 ( .A(n6331), .ZN(n4805) );
  NAND3_X1 U5995 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n5135), .ZN(n6335) );
  OR2_X1 U5996 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6335), .ZN(n4831)
         );
  AOI22_X1 U5997 ( .A1(n4806), .A2(n4805), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n4831), .ZN(n4807) );
  OAI211_X1 U5998 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6534), .A(n5139), .B(n4807), .ZN(n4829) );
  NAND2_X1 U5999 ( .A1(n4829), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4810)
         );
  OAI22_X1 U6000 ( .A1(n5152), .A2(n4831), .B1(n4830), .B2(n6323), .ZN(n4808)
         );
  AOI21_X1 U6001 ( .B1(n6369), .B2(n6318), .A(n4808), .ZN(n4809) );
  OAI211_X1 U6002 ( .C1(n4835), .C2(n5156), .A(n4810), .B(n4809), .ZN(U3105)
         );
  NAND2_X1 U6003 ( .A1(n4829), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4813)
         );
  OAI22_X1 U6004 ( .A1(n5142), .A2(n4831), .B1(n4830), .B2(n6285), .ZN(n4811)
         );
  AOI21_X1 U6005 ( .B1(n6369), .B2(n6273), .A(n4811), .ZN(n4812) );
  OAI211_X1 U6006 ( .C1(n4835), .C2(n5146), .A(n4813), .B(n4812), .ZN(U3100)
         );
  NAND2_X1 U6007 ( .A1(n4829), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4816)
         );
  OAI22_X1 U6008 ( .A1(n5157), .A2(n4831), .B1(n4830), .B2(n6385), .ZN(n4814)
         );
  AOI21_X1 U6009 ( .B1(n6369), .B2(n6375), .A(n4814), .ZN(n4815) );
  OAI211_X1 U6010 ( .C1(n4835), .C2(n5161), .A(n4816), .B(n4815), .ZN(U3107)
         );
  NAND2_X1 U6011 ( .A1(n4829), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4819)
         );
  OAI22_X1 U6012 ( .A1(n5147), .A2(n4831), .B1(n4830), .B2(n6304), .ZN(n4817)
         );
  AOI21_X1 U6013 ( .B1(n6369), .B2(n6301), .A(n4817), .ZN(n4818) );
  OAI211_X1 U6014 ( .C1(n4835), .C2(n5151), .A(n4819), .B(n4818), .ZN(U3106)
         );
  NAND2_X1 U6015 ( .A1(n4829), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4822)
         );
  OAI22_X1 U6016 ( .A1(n5162), .A2(n4831), .B1(n4830), .B2(n6293), .ZN(n4820)
         );
  AOI21_X1 U6017 ( .B1(n6369), .B2(n6290), .A(n4820), .ZN(n4821) );
  OAI211_X1 U6018 ( .C1(n4835), .C2(n5166), .A(n4822), .B(n4821), .ZN(U3102)
         );
  NAND2_X1 U6019 ( .A1(n4829), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4825)
         );
  OAI22_X1 U6020 ( .A1(n5167), .A2(n4831), .B1(n4830), .B2(n6361), .ZN(n4823)
         );
  AOI21_X1 U6021 ( .B1(n6369), .B2(n6356), .A(n4823), .ZN(n4824) );
  OAI211_X1 U6022 ( .C1(n4835), .C2(n5171), .A(n4825), .B(n4824), .ZN(U3104)
         );
  NAND2_X1 U6023 ( .A1(n4829), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4828)
         );
  OAI22_X1 U6024 ( .A1(n5172), .A2(n4831), .B1(n4830), .B2(n6397), .ZN(n4826)
         );
  AOI21_X1 U6025 ( .B1(n6369), .B2(n6392), .A(n4826), .ZN(n4827) );
  OAI211_X1 U6026 ( .C1(n4835), .C2(n5176), .A(n4828), .B(n4827), .ZN(U3103)
         );
  NAND2_X1 U6027 ( .A1(n4829), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4834)
         );
  OAI22_X1 U6028 ( .A1(n5179), .A2(n4831), .B1(n4830), .B2(n6289), .ZN(n4832)
         );
  AOI21_X1 U6029 ( .B1(n6369), .B2(n6286), .A(n4832), .ZN(n4833) );
  OAI211_X1 U6030 ( .C1(n4835), .C2(n5184), .A(n4834), .B(n4833), .ZN(U3101)
         );
  XOR2_X1 U6031 ( .A(n4837), .B(n4836), .Z(n4947) );
  INV_X1 U6032 ( .A(n4947), .ZN(n4850) );
  AOI21_X1 U6033 ( .B1(n4839), .B2(n4650), .A(n4838), .ZN(n6124) );
  AOI22_X1 U6034 ( .A1(n6005), .A2(n6124), .B1(n5551), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n4840) );
  OAI21_X1 U6035 ( .B1(n4850), .B2(n5348), .A(n4840), .ZN(U2852) );
  INV_X1 U6036 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6137) );
  INV_X1 U6037 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6473) );
  AOI22_X1 U6038 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .B1(
        n6137), .B2(n6473), .ZN(n4842) );
  AOI22_X1 U6039 ( .A1(n5981), .A2(n4842), .B1(REIP_REG_7__SCAN_IN), .B2(n5980), .ZN(n4848) );
  INV_X1 U6040 ( .A(n4945), .ZN(n4846) );
  AOI22_X1 U6041 ( .A1(n5987), .A2(n6124), .B1(n5986), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n4843) );
  OAI211_X1 U6042 ( .C1(n5997), .C2(n4844), .A(n4843), .B(n6159), .ZN(n4845)
         );
  AOI21_X1 U6043 ( .B1(n5968), .B2(n4846), .A(n4845), .ZN(n4847) );
  OAI211_X1 U6044 ( .C1(n4850), .C2(n5861), .A(n4848), .B(n4847), .ZN(U2820)
         );
  OAI222_X1 U6045 ( .A1(n5583), .A2(n4850), .B1(n5582), .B2(n4849), .C1(n5581), 
        .C2(n3801), .ZN(U2884) );
  OR2_X1 U6046 ( .A1(n6234), .A2(n4851), .ZN(n4852) );
  AND2_X1 U6047 ( .A1(n4852), .A2(n6327), .ZN(n4863) );
  OR2_X1 U6048 ( .A1(n4854), .A2(n4853), .ZN(n4904) );
  OR2_X1 U6049 ( .A1(n4855), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4901)
         );
  NOR2_X1 U6050 ( .A1(n6398), .A2(n4901), .ZN(n4887) );
  INV_X1 U6051 ( .A(n4887), .ZN(n4856) );
  OAI21_X1 U6052 ( .B1(n4904), .B2(n4857), .A(n4856), .ZN(n4861) );
  INV_X1 U6053 ( .A(n4901), .ZN(n4858) );
  AOI22_X1 U6054 ( .A1(n4863), .A2(n4861), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4858), .ZN(n4891) );
  NOR2_X2 U6055 ( .A1(n6234), .A2(n4859), .ZN(n6266) );
  NOR2_X1 U6056 ( .A1(n6234), .A2(n4860), .ZN(n6228) );
  INV_X1 U6057 ( .A(n4861), .ZN(n4862) );
  AOI22_X1 U6058 ( .A1(n4863), .A2(n4862), .B1(n4901), .B2(n6332), .ZN(n4864)
         );
  NAND2_X1 U6059 ( .A1(n6278), .A2(n4864), .ZN(n4886) );
  AOI22_X1 U6060 ( .A1(n6343), .A2(n4887), .B1(INSTQUEUE_REG_5__1__SCAN_IN), 
        .B2(n4886), .ZN(n4865) );
  OAI21_X1 U6061 ( .B1(n6289), .B2(n4927), .A(n4865), .ZN(n4866) );
  AOI21_X1 U6062 ( .B1(n6286), .B2(n6266), .A(n4866), .ZN(n4867) );
  OAI21_X1 U6063 ( .B1(n4891), .B2(n5184), .A(n4867), .ZN(U3061) );
  AOI22_X1 U6064 ( .A1(n6370), .A2(n4887), .B1(INSTQUEUE_REG_5__6__SCAN_IN), 
        .B2(n4886), .ZN(n4868) );
  OAI21_X1 U6065 ( .B1(n6304), .B2(n4927), .A(n4868), .ZN(n4869) );
  AOI21_X1 U6066 ( .B1(n6301), .B2(n6266), .A(n4869), .ZN(n4870) );
  OAI21_X1 U6067 ( .B1(n4891), .B2(n5151), .A(n4870), .ZN(U3066) );
  AOI22_X1 U6068 ( .A1(n6388), .A2(n4887), .B1(INSTQUEUE_REG_5__3__SCAN_IN), 
        .B2(n4886), .ZN(n4871) );
  OAI21_X1 U6069 ( .B1(n6397), .B2(n4927), .A(n4871), .ZN(n4872) );
  AOI21_X1 U6070 ( .B1(n6392), .B2(n6266), .A(n4872), .ZN(n4873) );
  OAI21_X1 U6071 ( .B1(n4891), .B2(n5176), .A(n4873), .ZN(U3063) );
  AOI22_X1 U6072 ( .A1(n6326), .A2(n4887), .B1(INSTQUEUE_REG_5__0__SCAN_IN), 
        .B2(n4886), .ZN(n4874) );
  OAI21_X1 U6073 ( .B1(n6285), .B2(n4927), .A(n4874), .ZN(n4875) );
  AOI21_X1 U6074 ( .B1(n6273), .B2(n6266), .A(n4875), .ZN(n4876) );
  OAI21_X1 U6075 ( .B1(n4891), .B2(n5146), .A(n4876), .ZN(U3060) );
  AOI22_X1 U6076 ( .A1(n6363), .A2(n4887), .B1(INSTQUEUE_REG_5__5__SCAN_IN), 
        .B2(n4886), .ZN(n4877) );
  OAI21_X1 U6077 ( .B1(n6323), .B2(n4927), .A(n4877), .ZN(n4878) );
  AOI21_X1 U6078 ( .B1(n6318), .B2(n6266), .A(n4878), .ZN(n4879) );
  OAI21_X1 U6079 ( .B1(n4891), .B2(n5156), .A(n4879), .ZN(U3065) );
  AOI22_X1 U6080 ( .A1(n6349), .A2(n4887), .B1(INSTQUEUE_REG_5__2__SCAN_IN), 
        .B2(n4886), .ZN(n4880) );
  OAI21_X1 U6081 ( .B1(n6293), .B2(n4927), .A(n4880), .ZN(n4881) );
  AOI21_X1 U6082 ( .B1(n6290), .B2(n6266), .A(n4881), .ZN(n4882) );
  OAI21_X1 U6083 ( .B1(n4891), .B2(n5166), .A(n4882), .ZN(U3062) );
  AOI22_X1 U6084 ( .A1(n6378), .A2(n4887), .B1(INSTQUEUE_REG_5__7__SCAN_IN), 
        .B2(n4886), .ZN(n4883) );
  OAI21_X1 U6085 ( .B1(n6385), .B2(n4927), .A(n4883), .ZN(n4884) );
  AOI21_X1 U6086 ( .B1(n6375), .B2(n6266), .A(n4884), .ZN(n4885) );
  OAI21_X1 U6087 ( .B1(n4891), .B2(n5161), .A(n4885), .ZN(U3067) );
  AOI22_X1 U6088 ( .A1(n6357), .A2(n4887), .B1(INSTQUEUE_REG_5__4__SCAN_IN), 
        .B2(n4886), .ZN(n4888) );
  OAI21_X1 U6089 ( .B1(n6361), .B2(n4927), .A(n4888), .ZN(n4889) );
  AOI21_X1 U6090 ( .B1(n6356), .B2(n6266), .A(n4889), .ZN(n4890) );
  OAI21_X1 U6091 ( .B1(n4891), .B2(n5171), .A(n4890), .ZN(U3064) );
  INV_X1 U6092 ( .A(n5003), .ZN(n4895) );
  AOI21_X1 U6093 ( .B1(n6076), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4892), 
        .ZN(n4893) );
  OAI21_X1 U6094 ( .B1(n6085), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4893), 
        .ZN(n4894) );
  AOI21_X1 U6095 ( .B1(n4895), .B2(n2983), .A(n4894), .ZN(n4896) );
  OAI21_X1 U6096 ( .B1(n4897), .B2(n6060), .A(n4896), .ZN(U2985) );
  AOI22_X1 U6097 ( .A1(n4900), .A2(n5993), .B1(n4899), .B2(n4898), .ZN(n6225)
         );
  NOR2_X1 U6098 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4901), .ZN(n6226)
         );
  OR2_X1 U6099 ( .A1(n5805), .A2(n4902), .ZN(n4903) );
  OR2_X1 U6100 ( .A1(n4903), .A2(n5810), .ZN(n6232) );
  OAI21_X1 U6101 ( .B1(n6228), .B2(n6218), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4905) );
  AND2_X1 U6102 ( .A1(n4905), .A2(n4904), .ZN(n4907) );
  AOI211_X1 U6103 ( .C1(n6327), .C2(n4907), .A(n5134), .B(n4906), .ZN(n4908)
         );
  OAI21_X1 U6104 ( .B1(n6226), .B2(n6519), .A(n4908), .ZN(n6229) );
  NAND2_X1 U6105 ( .A1(n6229), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4911) );
  INV_X1 U6106 ( .A(n6226), .ZN(n4928) );
  OAI22_X1 U6107 ( .A1(n5167), .A2(n4928), .B1(n4927), .B2(n6259), .ZN(n4909)
         );
  AOI21_X1 U6108 ( .B1(n6256), .B2(n6218), .A(n4909), .ZN(n4910) );
  OAI211_X1 U6109 ( .C1(n6225), .C2(n5171), .A(n4911), .B(n4910), .ZN(U3056)
         );
  NAND2_X1 U6110 ( .A1(n6229), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4914) );
  OAI22_X1 U6111 ( .A1(n5152), .A2(n4928), .B1(n4927), .B2(n6367), .ZN(n4912)
         );
  AOI21_X1 U6112 ( .B1(n6362), .B2(n6218), .A(n4912), .ZN(n4913) );
  OAI211_X1 U6113 ( .C1(n6225), .C2(n5156), .A(n4914), .B(n4913), .ZN(U3057)
         );
  NAND2_X1 U6114 ( .A1(n6229), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4917) );
  OAI22_X1 U6115 ( .A1(n5147), .A2(n4928), .B1(n4927), .B2(n6374), .ZN(n4915)
         );
  AOI21_X1 U6116 ( .B1(n6368), .B2(n6218), .A(n4915), .ZN(n4916) );
  OAI211_X1 U6117 ( .C1(n6225), .C2(n5151), .A(n4917), .B(n4916), .ZN(U3058)
         );
  NAND2_X1 U6118 ( .A1(n6229), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4920) );
  OAI22_X1 U6119 ( .A1(n5179), .A2(n4928), .B1(n4927), .B2(n6347), .ZN(n4918)
         );
  AOI21_X1 U6120 ( .B1(n6342), .B2(n6218), .A(n4918), .ZN(n4919) );
  OAI211_X1 U6121 ( .C1(n6225), .C2(n5184), .A(n4920), .B(n4919), .ZN(U3053)
         );
  NAND2_X1 U6122 ( .A1(n6229), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4923) );
  OAI22_X1 U6123 ( .A1(n5162), .A2(n4928), .B1(n4927), .B2(n6353), .ZN(n4921)
         );
  AOI21_X1 U6124 ( .B1(n6348), .B2(n6218), .A(n4921), .ZN(n4922) );
  OAI211_X1 U6125 ( .C1(n6225), .C2(n5166), .A(n4923), .B(n4922), .ZN(U3054)
         );
  NAND2_X1 U6126 ( .A1(n6229), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4926) );
  OAI22_X1 U6127 ( .A1(n5142), .A2(n4928), .B1(n4927), .B2(n6341), .ZN(n4924)
         );
  AOI21_X1 U6128 ( .B1(n6325), .B2(n6218), .A(n4924), .ZN(n4925) );
  OAI211_X1 U6129 ( .C1(n6225), .C2(n5146), .A(n4926), .B(n4925), .ZN(U3052)
         );
  NAND2_X1 U6130 ( .A1(n6229), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4931) );
  OAI22_X1 U6131 ( .A1(n5157), .A2(n4928), .B1(n4927), .B2(n6271), .ZN(n4929)
         );
  AOI21_X1 U6132 ( .B1(n6267), .B2(n6218), .A(n4929), .ZN(n4930) );
  OAI211_X1 U6133 ( .C1(n6225), .C2(n5161), .A(n4931), .B(n4930), .ZN(U3059)
         );
  CLKBUF_X1 U6134 ( .A(n4932), .Z(n4933) );
  OAI21_X1 U6135 ( .B1(n4933), .B2(n4935), .A(n4934), .ZN(n6149) );
  AOI22_X1 U6136 ( .A1(n6076), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n6185), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n4936) );
  OAI21_X1 U6137 ( .B1(n6085), .B2(n4937), .A(n4936), .ZN(n4938) );
  AOI21_X1 U6138 ( .B1(n4939), .B2(n2983), .A(n4938), .ZN(n4940) );
  OAI21_X1 U6139 ( .B1(n6060), .B2(n6149), .A(n4940), .ZN(U2981) );
  OAI21_X1 U6140 ( .B1(n4943), .B2(n4942), .A(n4941), .ZN(n6125) );
  NAND2_X1 U6141 ( .A1(n6185), .A2(REIP_REG_7__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U6142 ( .A1(n6076), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4944)
         );
  OAI211_X1 U6143 ( .C1(n6085), .C2(n4945), .A(n6122), .B(n4944), .ZN(n4946)
         );
  AOI21_X1 U6144 ( .B1(n4947), .B2(n2983), .A(n4946), .ZN(n4948) );
  OAI21_X1 U6145 ( .B1(n6125), .B2(n6060), .A(n4948), .ZN(U2979) );
  OR2_X1 U6146 ( .A1(n5327), .A2(REIP_REG_1__SCAN_IN), .ZN(n4994) );
  AND2_X1 U6147 ( .A1(n4994), .A2(REIP_REG_2__SCAN_IN), .ZN(n4949) );
  NAND2_X1 U6148 ( .A1(n4950), .A2(n4949), .ZN(n5995) );
  INV_X1 U6149 ( .A(n5995), .ZN(n4956) );
  AOI21_X1 U6150 ( .B1(n5991), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n4955) );
  INV_X1 U6151 ( .A(n6084), .ZN(n4951) );
  AOI22_X1 U6152 ( .A1(n5956), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n5968), 
        .B2(n4951), .ZN(n4954) );
  AOI22_X1 U6153 ( .A1(n5806), .A2(n4952), .B1(EBX_REG_2__SCAN_IN), .B2(n5986), 
        .ZN(n4953) );
  OAI211_X1 U6154 ( .C1(n4956), .C2(n4955), .A(n4954), .B(n4953), .ZN(n4957)
         );
  AOI21_X1 U6155 ( .B1(n5987), .B2(n6181), .A(n4957), .ZN(n4958) );
  OAI21_X1 U6156 ( .B1(n4959), .B2(n5989), .A(n4958), .ZN(U2825) );
  NAND2_X1 U6157 ( .A1(n4960), .A2(n4961), .ZN(n4964) );
  NAND2_X1 U6158 ( .A1(n4964), .A2(n4962), .ZN(n4963) );
  OAI21_X1 U6159 ( .B1(n4964), .B2(n4962), .A(n4963), .ZN(n6156) );
  NAND2_X1 U6160 ( .A1(n4965), .A2(n2983), .ZN(n4970) );
  INV_X1 U6161 ( .A(n6085), .ZN(n6056) );
  OAI22_X1 U6162 ( .A1(n5681), .A2(n4966), .B1(n6159), .B2(n6158), .ZN(n4967)
         );
  AOI21_X1 U6163 ( .B1(n4968), .B2(n6056), .A(n4967), .ZN(n4969) );
  OAI211_X1 U6164 ( .C1(n6156), .C2(n6060), .A(n4970), .B(n4969), .ZN(U2982)
         );
  OR2_X1 U6165 ( .A1(n5008), .A2(n4973), .ZN(n5021) );
  INV_X1 U6166 ( .A(n5021), .ZN(n4972) );
  AOI21_X1 U6167 ( .B1(n4973), .B2(n5008), .A(n4972), .ZN(n4990) );
  INV_X1 U6168 ( .A(n4990), .ZN(n4992) );
  INV_X1 U6169 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6475) );
  NAND3_X1 U6170 ( .A1(n5981), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .ZN(n5012) );
  NAND2_X1 U6171 ( .A1(n6475), .A2(n5012), .ZN(n4980) );
  NOR3_X1 U6172 ( .A1(n6475), .A2(n6473), .A3(n6137), .ZN(n5210) );
  AOI21_X1 U6173 ( .B1(n5216), .B2(n5210), .A(n5483), .ZN(n5965) );
  OAI21_X1 U6174 ( .B1(n4974), .B2(n4838), .A(n5025), .ZN(n6116) );
  NOR2_X1 U6175 ( .A1(n6116), .A2(n5938), .ZN(n4977) );
  OAI21_X1 U6176 ( .B1(n5974), .B2(n4975), .A(n6159), .ZN(n4976) );
  AOI211_X1 U6177 ( .C1(n5956), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n4977), 
        .B(n4976), .ZN(n4978) );
  OAI21_X1 U6178 ( .B1(n4988), .B2(n5996), .A(n4978), .ZN(n4979) );
  AOI21_X1 U6179 ( .B1(n4980), .B2(n5965), .A(n4979), .ZN(n4981) );
  OAI21_X1 U6180 ( .B1(n4992), .B2(n5861), .A(n4981), .ZN(U2819) );
  INV_X1 U6181 ( .A(n6116), .ZN(n4982) );
  AOI22_X1 U6182 ( .A1(n6005), .A2(n4982), .B1(n5551), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4983) );
  OAI21_X1 U6183 ( .B1(n4992), .B2(n5348), .A(n4983), .ZN(U2851) );
  OAI21_X1 U6184 ( .B1(n4986), .B2(n4985), .A(n4984), .ZN(n6115) );
  AOI22_X1 U6185 ( .A1(n6076), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6185), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n4987) );
  OAI21_X1 U6186 ( .B1(n6085), .B2(n4988), .A(n4987), .ZN(n4989) );
  AOI21_X1 U6187 ( .B1(n4990), .B2(n2983), .A(n4989), .ZN(n4991) );
  OAI21_X1 U6188 ( .B1(n6115), .B2(n6060), .A(n4991), .ZN(U2978) );
  INV_X1 U6189 ( .A(DATAI_8_), .ZN(n6647) );
  OAI222_X1 U6190 ( .A1(n4992), .A2(n5583), .B1(n5582), .B2(n6647), .C1(n5581), 
        .C2(n6033), .ZN(U2883) );
  NAND2_X1 U6191 ( .A1(n4993), .A2(REIP_REG_1__SCAN_IN), .ZN(n4999) );
  OAI21_X1 U6192 ( .B1(n5974), .B2(n4995), .A(n4994), .ZN(n4996) );
  AOI21_X1 U6193 ( .B1(n4997), .B2(n5987), .A(n4996), .ZN(n4998) );
  OAI211_X1 U6194 ( .C1(n5992), .C2(n5824), .A(n4999), .B(n4998), .ZN(n5001)
         );
  NOR2_X1 U6195 ( .A1(n5996), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5000)
         );
  AOI211_X1 U6196 ( .C1(n5956), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n5001), 
        .B(n5000), .ZN(n5002) );
  OAI21_X1 U6197 ( .B1(n5989), .B2(n5003), .A(n5002), .ZN(U2826) );
  NOR2_X1 U6198 ( .A1(n5008), .A2(n5004), .ZN(n5011) );
  NOR2_X1 U6199 ( .A1(n5011), .A2(n5005), .ZN(n5006) );
  OR2_X1 U6200 ( .A1(n5075), .A2(n5006), .ZN(n5957) );
  INV_X1 U6201 ( .A(DATAI_11_), .ZN(n6598) );
  OAI222_X1 U6202 ( .A1(n5957), .A2(n5583), .B1(n5582), .B2(n6598), .C1(n5581), 
        .C2(n6027), .ZN(U2880) );
  NOR2_X1 U6203 ( .A1(n5008), .A2(n5007), .ZN(n5022) );
  NOR2_X1 U6204 ( .A1(n5022), .A2(n5009), .ZN(n5010) );
  OR2_X1 U6205 ( .A1(n5011), .A2(n5010), .ZN(n5074) );
  NOR2_X1 U6206 ( .A1(n6475), .A2(n5012), .ZN(n5949) );
  NAND2_X1 U6207 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5961) );
  OAI211_X1 U6208 ( .C1(REIP_REG_10__SCAN_IN), .C2(REIP_REG_9__SCAN_IN), .A(
        n5949), .B(n5961), .ZN(n5019) );
  INV_X1 U6209 ( .A(n5070), .ZN(n5017) );
  INV_X1 U6210 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5031) );
  AOI21_X1 U6211 ( .B1(n5956), .B2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6185), 
        .ZN(n5015) );
  XNOR2_X1 U6212 ( .A(n5013), .B(n5024), .ZN(n5030) );
  INV_X1 U6213 ( .A(n5030), .ZN(n6095) );
  AOI22_X1 U6214 ( .A1(n5965), .A2(REIP_REG_10__SCAN_IN), .B1(n5987), .B2(
        n6095), .ZN(n5014) );
  OAI211_X1 U6215 ( .C1(n5031), .C2(n5974), .A(n5015), .B(n5014), .ZN(n5016)
         );
  AOI21_X1 U6216 ( .B1(n5968), .B2(n5017), .A(n5016), .ZN(n5018) );
  OAI211_X1 U6217 ( .C1(n5074), .C2(n5861), .A(n5019), .B(n5018), .ZN(U2817)
         );
  AND2_X1 U6218 ( .A1(n5021), .A2(n5020), .ZN(n5023) );
  AOI21_X1 U6219 ( .B1(n5026), .B2(n5025), .A(n5024), .ZN(n6109) );
  AOI22_X1 U6220 ( .A1(n6005), .A2(n6109), .B1(n5551), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n5027) );
  OAI21_X1 U6221 ( .B1(n5966), .B2(n5348), .A(n5027), .ZN(U2850) );
  INV_X1 U6222 ( .A(DATAI_10_), .ZN(n5028) );
  OAI222_X1 U6223 ( .A1(n5074), .A2(n5583), .B1(n5582), .B2(n5028), .C1(n5581), 
        .C2(n6029), .ZN(U2881) );
  INV_X1 U6224 ( .A(DATAI_9_), .ZN(n5029) );
  OAI222_X1 U6225 ( .A1(n5966), .A2(n5583), .B1(n5582), .B2(n5029), .C1(n5581), 
        .C2(n6031), .ZN(U2882) );
  OAI222_X1 U6226 ( .A1(n5553), .A2(n5074), .B1(n6009), .B2(n5031), .C1(n5549), 
        .C2(n5030), .ZN(U2849) );
  NAND2_X1 U6227 ( .A1(n5034), .A2(n5033), .ZN(n5035) );
  XNOR2_X1 U6228 ( .A(n5032), .B(n5035), .ZN(n6111) );
  INV_X1 U6229 ( .A(n6060), .ZN(n6081) );
  NAND2_X1 U6230 ( .A1(n6111), .A2(n6081), .ZN(n5038) );
  NAND2_X1 U6231 ( .A1(n6185), .A2(REIP_REG_9__SCAN_IN), .ZN(n6107) );
  OAI21_X1 U6232 ( .B1(n5681), .B2(n5963), .A(n6107), .ZN(n5036) );
  AOI21_X1 U6233 ( .B1(n6056), .B2(n5967), .A(n5036), .ZN(n5037) );
  OAI211_X1 U6234 ( .C1(n5687), .C2(n5966), .A(n5038), .B(n5037), .ZN(U2977)
         );
  NOR2_X1 U6235 ( .A1(n6398), .A2(n5043), .ZN(n5064) );
  AOI21_X1 U6236 ( .B1(n5039), .B2(n6330), .A(n5064), .ZN(n5044) );
  AOI21_X1 U6237 ( .B1(n5040), .B2(STATEBS16_REG_SCAN_IN), .A(n6332), .ZN(
        n5042) );
  AOI22_X1 U6238 ( .A1(n5044), .A2(n5042), .B1(n6332), .B2(n5043), .ZN(n5041)
         );
  NAND2_X1 U6239 ( .A1(n6278), .A2(n5041), .ZN(n5063) );
  INV_X1 U6240 ( .A(n5042), .ZN(n5045) );
  OAI22_X1 U6241 ( .A1(n5045), .A2(n5044), .B1(n6534), .B2(n5043), .ZN(n5062)
         );
  AOI22_X1 U6242 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5063), .B1(n6390), 
        .B2(n5062), .ZN(n5049) );
  NOR2_X2 U6243 ( .A1(n5047), .A2(n5046), .ZN(n5181) );
  AOI22_X1 U6244 ( .A1(n6388), .A2(n5064), .B1(n6392), .B2(n5181), .ZN(n5048)
         );
  OAI211_X1 U6245 ( .C1(n6397), .C2(n5067), .A(n5049), .B(n5048), .ZN(U3031)
         );
  AOI22_X1 U6246 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5063), .B1(n6364), 
        .B2(n5062), .ZN(n5051) );
  AOI22_X1 U6247 ( .A1(n6363), .A2(n5064), .B1(n6318), .B2(n5181), .ZN(n5050)
         );
  OAI211_X1 U6248 ( .C1(n6323), .C2(n5067), .A(n5051), .B(n5050), .ZN(U3033)
         );
  AOI22_X1 U6249 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5063), .B1(n6344), 
        .B2(n5062), .ZN(n5053) );
  AOI22_X1 U6250 ( .A1(n6343), .A2(n5064), .B1(n6286), .B2(n5181), .ZN(n5052)
         );
  OAI211_X1 U6251 ( .C1(n6289), .C2(n5067), .A(n5053), .B(n5052), .ZN(U3029)
         );
  AOI22_X1 U6252 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5063), .B1(n6350), 
        .B2(n5062), .ZN(n5055) );
  AOI22_X1 U6253 ( .A1(n6349), .A2(n5064), .B1(n6290), .B2(n5181), .ZN(n5054)
         );
  OAI211_X1 U6254 ( .C1(n6293), .C2(n5067), .A(n5055), .B(n5054), .ZN(U3030)
         );
  AOI22_X1 U6255 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5063), .B1(n6358), 
        .B2(n5062), .ZN(n5057) );
  AOI22_X1 U6256 ( .A1(n6357), .A2(n5064), .B1(n6356), .B2(n5181), .ZN(n5056)
         );
  OAI211_X1 U6257 ( .C1(n6361), .C2(n5067), .A(n5057), .B(n5056), .ZN(U3032)
         );
  AOI22_X1 U6258 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5063), .B1(n6380), 
        .B2(n5062), .ZN(n5059) );
  AOI22_X1 U6259 ( .A1(n6378), .A2(n5064), .B1(n6375), .B2(n5181), .ZN(n5058)
         );
  OAI211_X1 U6260 ( .C1(n6385), .C2(n5067), .A(n5059), .B(n5058), .ZN(U3035)
         );
  AOI22_X1 U6261 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5063), .B1(n6338), 
        .B2(n5062), .ZN(n5061) );
  AOI22_X1 U6262 ( .A1(n6326), .A2(n5064), .B1(n6273), .B2(n5181), .ZN(n5060)
         );
  OAI211_X1 U6263 ( .C1(n6285), .C2(n5067), .A(n5061), .B(n5060), .ZN(U3028)
         );
  AOI22_X1 U6264 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5063), .B1(n6371), 
        .B2(n5062), .ZN(n5066) );
  AOI22_X1 U6265 ( .A1(n6370), .A2(n5064), .B1(n6301), .B2(n5181), .ZN(n5065)
         );
  OAI211_X1 U6266 ( .C1(n6304), .C2(n5067), .A(n5066), .B(n5065), .ZN(U3034)
         );
  NAND2_X1 U6267 ( .A1(n6051), .A2(n5068), .ZN(n5069) );
  XNOR2_X1 U6268 ( .A(n2989), .B(n5069), .ZN(n6103) );
  NAND2_X1 U6269 ( .A1(n6103), .A2(n6081), .ZN(n5073) );
  AND2_X1 U6270 ( .A1(n6185), .A2(REIP_REG_10__SCAN_IN), .ZN(n6094) );
  NOR2_X1 U6271 ( .A1(n6085), .A2(n5070), .ZN(n5071) );
  AOI211_X1 U6272 ( .C1(n6076), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6094), 
        .B(n5071), .ZN(n5072) );
  OAI211_X1 U6273 ( .C1(n5687), .C2(n5074), .A(n5073), .B(n5072), .ZN(U2976)
         );
  XOR2_X1 U6274 ( .A(n5076), .B(n5075), .Z(n5114) );
  INV_X1 U6275 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5084) );
  INV_X1 U6276 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6480) );
  NOR2_X1 U6277 ( .A1(n6480), .A2(n5961), .ZN(n5211) );
  INV_X1 U6278 ( .A(n5211), .ZN(n5077) );
  AOI21_X1 U6279 ( .B1(n5077), .B2(n5835), .A(n5965), .ZN(n5953) );
  INV_X1 U6280 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5085) );
  OR2_X1 U6281 ( .A1(n5079), .A2(n5078), .ZN(n5081) );
  AND2_X1 U6282 ( .A1(n5081), .A2(n5080), .ZN(n5123) );
  INV_X1 U6283 ( .A(n5123), .ZN(n5104) );
  OAI22_X1 U6284 ( .A1(n5953), .A2(n5085), .B1(n5938), .B2(n5104), .ZN(n5082)
         );
  AOI21_X1 U6285 ( .B1(EBX_REG_12__SCAN_IN), .B2(n5986), .A(n5082), .ZN(n5083)
         );
  OAI211_X1 U6286 ( .C1(n5997), .C2(n5084), .A(n5083), .B(n6159), .ZN(n5087)
         );
  NAND3_X1 U6287 ( .A1(n5211), .A2(n5949), .A3(n5085), .ZN(n5942) );
  OAI21_X1 U6288 ( .B1(n5112), .B2(n5996), .A(n5942), .ZN(n5086) );
  AOI211_X1 U6289 ( .C1(n5114), .C2(n5983), .A(n5087), .B(n5086), .ZN(n5088)
         );
  INV_X1 U6290 ( .A(n5088), .ZN(U2815) );
  AOI22_X1 U6291 ( .A1(n6425), .A2(UWORD_REG_0__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5089) );
  OAI21_X1 U6292 ( .B1(n5090), .B2(n5101), .A(n5089), .ZN(U2907) );
  AOI22_X1 U6293 ( .A1(n6425), .A2(UWORD_REG_1__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5091) );
  OAI21_X1 U6294 ( .B1(n3951), .B2(n5101), .A(n5091), .ZN(U2906) );
  AOI22_X1 U6295 ( .A1(n6425), .A2(UWORD_REG_2__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5092) );
  OAI21_X1 U6296 ( .B1(n3970), .B2(n5101), .A(n5092), .ZN(U2905) );
  AOI22_X1 U6297 ( .A1(n6425), .A2(UWORD_REG_3__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5093) );
  OAI21_X1 U6298 ( .B1(n5094), .B2(n5101), .A(n5093), .ZN(U2904) );
  AOI22_X1 U6299 ( .A1(n6425), .A2(UWORD_REG_4__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n5095) );
  OAI21_X1 U6300 ( .B1(n4004), .B2(n5101), .A(n5095), .ZN(U2903) );
  AOI22_X1 U6301 ( .A1(n6425), .A2(UWORD_REG_5__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n5096) );
  OAI21_X1 U6302 ( .B1(n5097), .B2(n5101), .A(n5096), .ZN(U2902) );
  AOI22_X1 U6303 ( .A1(n6540), .A2(UWORD_REG_7__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n5098) );
  OAI21_X1 U6304 ( .B1(n5099), .B2(n5101), .A(n5098), .ZN(U2900) );
  AOI22_X1 U6305 ( .A1(n6540), .A2(UWORD_REG_6__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n5100) );
  OAI21_X1 U6306 ( .B1(n5102), .B2(n5101), .A(n5100), .ZN(U2901) );
  INV_X1 U6307 ( .A(n5114), .ZN(n5103) );
  INV_X1 U6308 ( .A(DATAI_12_), .ZN(n6664) );
  OAI222_X1 U6309 ( .A1(n5583), .A2(n5103), .B1(n5582), .B2(n6664), .C1(n5581), 
        .C2(n6025), .ZN(U2879) );
  OAI222_X1 U6310 ( .A1(n5549), .A2(n5104), .B1(n6009), .B2(n3667), .C1(n5553), 
        .C2(n5103), .ZN(U2847) );
  CLKBUF_X1 U6311 ( .A(n5105), .Z(n5106) );
  INV_X1 U6312 ( .A(n5107), .ZN(n5108) );
  NOR2_X1 U6313 ( .A1(n5109), .A2(n5108), .ZN(n5110) );
  XNOR2_X1 U6314 ( .A(n5106), .B(n5110), .ZN(n5125) );
  NOR2_X1 U6315 ( .A1(n6159), .A2(n5085), .ZN(n5122) );
  AOI21_X1 U6316 ( .B1(n6076), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n5122), 
        .ZN(n5111) );
  OAI21_X1 U6317 ( .B1(n6085), .B2(n5112), .A(n5111), .ZN(n5113) );
  AOI21_X1 U6318 ( .B1(n5114), .B2(n2983), .A(n5113), .ZN(n5115) );
  OAI21_X1 U6319 ( .B1(n5125), .B2(n6060), .A(n5115), .ZN(U2974) );
  AOI21_X1 U6321 ( .B1(n5116), .B2(n6146), .A(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n5117) );
  NOR2_X1 U6322 ( .A1(n5117), .A2(n6088), .ZN(n5119) );
  OAI33_X1 U6323 ( .A1(1'b0), .A2(n5119), .A3(n5118), .B1(
        INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n5901), .B3(n3485), .ZN(n5121)
         );
  AOI211_X1 U6324 ( .C1(n6180), .C2(n5123), .A(n5122), .B(n5121), .ZN(n5124)
         );
  OAI21_X1 U6325 ( .B1(n5125), .B2(n6157), .A(n5124), .ZN(U3006) );
  OAI21_X1 U6326 ( .B1(n5128), .B2(n5127), .A(n5126), .ZN(n5870) );
  AOI21_X1 U6327 ( .B1(n5130), .B2(n5080), .A(n5129), .ZN(n5936) );
  AOI22_X1 U6328 ( .A1(n6005), .A2(n5936), .B1(n5551), .B2(EBX_REG_13__SCAN_IN), .ZN(n5131) );
  OAI21_X1 U6329 ( .B1(n5870), .B2(n5348), .A(n5131), .ZN(U2846) );
  AND2_X1 U6330 ( .A1(n5993), .A2(n5132), .ZN(n6197) );
  NOR2_X1 U6331 ( .A1(n5133), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6235)
         );
  AOI22_X1 U6332 ( .A1(n6197), .A2(n6327), .B1(n5134), .B2(n6235), .ZN(n5185)
         );
  NAND3_X1 U6333 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6409), .A3(n5135), .ZN(n6200) );
  NOR2_X1 U6334 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6200), .ZN(n5141)
         );
  OR2_X1 U6335 ( .A1(n5805), .A2(n6233), .ZN(n5136) );
  INV_X1 U6336 ( .A(n6224), .ZN(n6207) );
  OAI21_X1 U6337 ( .B1(n5181), .B2(n6207), .A(n5815), .ZN(n5138) );
  INV_X1 U6338 ( .A(n6197), .ZN(n5137) );
  NAND2_X1 U6339 ( .A1(n5138), .A2(n5137), .ZN(n5140) );
  OAI221_X1 U6340 ( .B1(n5141), .B2(n6519), .C1(n5141), .C2(n5140), .A(n5139), 
        .ZN(n5177) );
  NAND2_X1 U6341 ( .A1(n5177), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5145) );
  INV_X1 U6342 ( .A(n5141), .ZN(n5178) );
  OAI22_X1 U6343 ( .A1(n5142), .A2(n5178), .B1(n6341), .B2(n6224), .ZN(n5143)
         );
  AOI21_X1 U6344 ( .B1(n6325), .B2(n5181), .A(n5143), .ZN(n5144) );
  OAI211_X1 U6345 ( .C1(n5185), .C2(n5146), .A(n5145), .B(n5144), .ZN(U3036)
         );
  NAND2_X1 U6346 ( .A1(n5177), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5150) );
  OAI22_X1 U6347 ( .A1(n5147), .A2(n5178), .B1(n6374), .B2(n6224), .ZN(n5148)
         );
  AOI21_X1 U6348 ( .B1(n6368), .B2(n5181), .A(n5148), .ZN(n5149) );
  OAI211_X1 U6349 ( .C1(n5185), .C2(n5151), .A(n5150), .B(n5149), .ZN(U3042)
         );
  NAND2_X1 U6350 ( .A1(n5177), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5155) );
  OAI22_X1 U6351 ( .A1(n5152), .A2(n5178), .B1(n6367), .B2(n6224), .ZN(n5153)
         );
  AOI21_X1 U6352 ( .B1(n6362), .B2(n5181), .A(n5153), .ZN(n5154) );
  OAI211_X1 U6353 ( .C1(n5185), .C2(n5156), .A(n5155), .B(n5154), .ZN(U3041)
         );
  NAND2_X1 U6354 ( .A1(n5177), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5160) );
  OAI22_X1 U6355 ( .A1(n5157), .A2(n5178), .B1(n6271), .B2(n6224), .ZN(n5158)
         );
  AOI21_X1 U6356 ( .B1(n6267), .B2(n5181), .A(n5158), .ZN(n5159) );
  OAI211_X1 U6357 ( .C1(n5185), .C2(n5161), .A(n5160), .B(n5159), .ZN(U3043)
         );
  NAND2_X1 U6358 ( .A1(n5177), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5165) );
  OAI22_X1 U6359 ( .A1(n5162), .A2(n5178), .B1(n6353), .B2(n6224), .ZN(n5163)
         );
  AOI21_X1 U6360 ( .B1(n6348), .B2(n5181), .A(n5163), .ZN(n5164) );
  OAI211_X1 U6361 ( .C1(n5185), .C2(n5166), .A(n5165), .B(n5164), .ZN(U3038)
         );
  NAND2_X1 U6362 ( .A1(n5177), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5170) );
  OAI22_X1 U6363 ( .A1(n5167), .A2(n5178), .B1(n6259), .B2(n6224), .ZN(n5168)
         );
  AOI21_X1 U6364 ( .B1(n6256), .B2(n5181), .A(n5168), .ZN(n5169) );
  OAI211_X1 U6365 ( .C1(n5185), .C2(n5171), .A(n5170), .B(n5169), .ZN(U3040)
         );
  NAND2_X1 U6366 ( .A1(n5177), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5175) );
  OAI22_X1 U6367 ( .A1(n5172), .A2(n5178), .B1(n6255), .B2(n6224), .ZN(n5173)
         );
  AOI21_X1 U6368 ( .B1(n6252), .B2(n5181), .A(n5173), .ZN(n5174) );
  OAI211_X1 U6369 ( .C1(n5185), .C2(n5176), .A(n5175), .B(n5174), .ZN(U3039)
         );
  NAND2_X1 U6370 ( .A1(n5177), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5183) );
  OAI22_X1 U6371 ( .A1(n5179), .A2(n5178), .B1(n6347), .B2(n6224), .ZN(n5180)
         );
  AOI21_X1 U6372 ( .B1(n6342), .B2(n5181), .A(n5180), .ZN(n5182) );
  OAI211_X1 U6373 ( .C1(n5185), .C2(n5184), .A(n5183), .B(n5182), .ZN(U3037)
         );
  INV_X1 U6374 ( .A(DATAI_13_), .ZN(n6601) );
  OAI222_X1 U6375 ( .A1(n5870), .A2(n5583), .B1(n5582), .B2(n6601), .C1(n5581), 
        .C2(n6023), .ZN(U2878) );
  OAI21_X1 U6376 ( .B1(n5188), .B2(n5187), .A(n5494), .ZN(n5226) );
  INV_X1 U6377 ( .A(DATAI_14_), .ZN(n6547) );
  OAI222_X1 U6378 ( .A1(n5226), .A2(n5583), .B1(n5582), .B2(n6547), .C1(n5581), 
        .C2(n6021), .ZN(U2877) );
  INV_X1 U6379 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5190) );
  OAI21_X1 U6380 ( .B1(n5189), .B2(n5129), .A(n5496), .ZN(n5229) );
  OAI222_X1 U6381 ( .A1(n5226), .A2(n5553), .B1(n6009), .B2(n5190), .C1(n5229), 
        .C2(n5549), .ZN(U2845) );
  XNOR2_X1 U6382 ( .A(n3477), .B(n5193), .ZN(n5194) );
  XNOR2_X1 U6383 ( .A(n5192), .B(n5194), .ZN(n5257) );
  NAND3_X1 U6384 ( .A1(n5199), .A2(n5193), .A3(n6087), .ZN(n5205) );
  AOI21_X1 U6385 ( .B1(n5196), .B2(n5195), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5201) );
  AOI21_X1 U6386 ( .B1(n5197), .B2(n5895), .A(n6088), .ZN(n5198) );
  OAI21_X1 U6387 ( .B1(n5200), .B2(n5199), .A(n5198), .ZN(n5896) );
  OR2_X1 U6388 ( .A1(n5201), .A2(n5896), .ZN(n5203) );
  INV_X1 U6389 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6485) );
  OAI22_X1 U6390 ( .A1(n6160), .A2(n5229), .B1(n6485), .B2(n6159), .ZN(n5202)
         );
  AOI21_X1 U6391 ( .B1(n5203), .B2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n5202), 
        .ZN(n5204) );
  OAI211_X1 U6392 ( .C1(n5257), .C2(n6157), .A(n5205), .B(n5204), .ZN(U3004)
         );
  OR2_X1 U6393 ( .A1(n5494), .A2(n5495), .ZN(n5492) );
  AND2_X1 U6394 ( .A1(n5492), .A2(n5206), .ZN(n5209) );
  OR2_X1 U6395 ( .A1(n5209), .A2(n5208), .ZN(n5693) );
  INV_X1 U6396 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6482) );
  INV_X1 U6397 ( .A(n5210), .ZN(n5212) );
  NAND2_X1 U6398 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5211), .ZN(n5941) );
  NOR3_X1 U6399 ( .A1(n6482), .A2(n5212), .A3(n5941), .ZN(n5217) );
  NAND2_X1 U6400 ( .A1(n5981), .A2(n5217), .ZN(n5234) );
  NAND2_X1 U6401 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n5239) );
  OAI211_X1 U6402 ( .C1(REIP_REG_16__SCAN_IN), .C2(REIP_REG_15__SCAN_IN), .A(
        n5498), .B(n5239), .ZN(n5224) );
  NOR2_X1 U6403 ( .A1(n5214), .A2(n5213), .ZN(n5215) );
  OR2_X1 U6404 ( .A1(n5240), .A2(n5215), .ZN(n5881) );
  INV_X1 U6405 ( .A(n5881), .ZN(n5222) );
  INV_X1 U6406 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6488) );
  NAND3_X1 U6407 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5217), .A3(n5216), .ZN(
        n5238) );
  NAND2_X1 U6408 ( .A1(n5835), .A2(n5238), .ZN(n5507) );
  AOI21_X1 U6409 ( .B1(n5956), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6185), 
        .ZN(n5220) );
  AOI22_X1 U6410 ( .A1(EBX_REG_16__SCAN_IN), .A2(n5986), .B1(n5218), .B2(n5968), .ZN(n5219) );
  OAI211_X1 U6411 ( .C1(n6488), .C2(n5507), .A(n5220), .B(n5219), .ZN(n5221)
         );
  AOI21_X1 U6412 ( .B1(n5222), .B2(n5987), .A(n5221), .ZN(n5223) );
  OAI211_X1 U6413 ( .C1(n5693), .C2(n5861), .A(n5224), .B(n5223), .ZN(U2811)
         );
  INV_X1 U6414 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5225) );
  OAI222_X1 U6415 ( .A1(n5693), .A2(n5348), .B1(n5225), .B2(n6009), .C1(n5549), 
        .C2(n5881), .ZN(U2843) );
  INV_X1 U6416 ( .A(n5226), .ZN(n5255) );
  NAND2_X1 U6417 ( .A1(n5255), .A2(n5983), .ZN(n5233) );
  AOI22_X1 U6418 ( .A1(EBX_REG_14__SCAN_IN), .A2(n5986), .B1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n5956), .ZN(n5227) );
  OAI211_X1 U6419 ( .C1(n6485), .C2(n5507), .A(n5227), .B(n6159), .ZN(n5231)
         );
  NAND2_X1 U6420 ( .A1(n5968), .A2(n5251), .ZN(n5228) );
  OAI21_X1 U6421 ( .B1(n5229), .B2(n5938), .A(n5228), .ZN(n5230) );
  NOR2_X1 U6422 ( .A1(n5231), .A2(n5230), .ZN(n5232) );
  OAI211_X1 U6423 ( .C1(REIP_REG_14__SCAN_IN), .C2(n5234), .A(n5233), .B(n5232), .ZN(U2813) );
  OAI21_X1 U6424 ( .B1(n5208), .B2(n5237), .A(n5236), .ZN(n5686) );
  INV_X1 U6425 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6490) );
  NAND3_X1 U6426 ( .A1(n5498), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U6427 ( .A1(n6490), .A2(n5332), .ZN(n5248) );
  NOR3_X1 U6428 ( .A1(n6490), .A2(n5239), .A3(n5238), .ZN(n5320) );
  NOR2_X1 U6429 ( .A1(n5320), .A2(n5483), .ZN(n5926) );
  INV_X1 U6430 ( .A(n5683), .ZN(n5246) );
  OR2_X1 U6431 ( .A1(n5241), .A2(n5240), .ZN(n5242) );
  AND2_X1 U6432 ( .A1(n5538), .A2(n5242), .ZN(n5874) );
  OAI22_X1 U6433 ( .A1(n5243), .A2(n5974), .B1(n5680), .B2(n5997), .ZN(n5244)
         );
  AOI211_X1 U6434 ( .C1(n5874), .C2(n5987), .A(n5244), .B(n6185), .ZN(n5245)
         );
  OAI21_X1 U6435 ( .B1(n5996), .B2(n5246), .A(n5245), .ZN(n5247) );
  AOI21_X1 U6436 ( .B1(n5248), .B2(n5926), .A(n5247), .ZN(n5249) );
  OAI21_X1 U6437 ( .B1(n5686), .B2(n5861), .A(n5249), .ZN(U2810) );
  AOI22_X1 U6438 ( .A1(n6005), .A2(n5874), .B1(n5551), .B2(EBX_REG_17__SCAN_IN), .ZN(n5250) );
  OAI21_X1 U6439 ( .B1(n5686), .B2(n5553), .A(n5250), .ZN(U2842) );
  INV_X1 U6440 ( .A(n5251), .ZN(n5253) );
  AOI22_X1 U6441 ( .A1(n6076), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6185), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5252) );
  OAI21_X1 U6442 ( .B1(n6085), .B2(n5253), .A(n5252), .ZN(n5254) );
  AOI21_X1 U6443 ( .B1(n5255), .B2(n2983), .A(n5254), .ZN(n5256) );
  OAI21_X1 U6444 ( .B1(n5257), .B2(n6060), .A(n5256), .ZN(U2972) );
  NOR2_X2 U6445 ( .A1(n6013), .A2(n5258), .ZN(n6010) );
  AOI22_X1 U6446 ( .A1(n6010), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n6013), .ZN(n5261) );
  NOR3_X4 U6447 ( .A1(n6013), .A2(n5387), .A3(n5259), .ZN(n6014) );
  NAND2_X1 U6448 ( .A1(n6014), .A2(DATAI_1_), .ZN(n5260) );
  OAI211_X1 U6449 ( .C1(n5686), .C2(n5583), .A(n5261), .B(n5260), .ZN(U2874)
         );
  INV_X1 U6450 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5262) );
  OAI22_X1 U6451 ( .A1(n5331), .A2(n5549), .B1(n6009), .B2(n5262), .ZN(U2828)
         );
  XNOR2_X1 U6452 ( .A(n5264), .B(n5263), .ZN(n5352) );
  AOI22_X1 U6453 ( .A1(n2984), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n5265), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5272) );
  AOI22_X1 U6454 ( .A1(n4189), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5271) );
  AOI22_X1 U6455 ( .A1(n3129), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5266), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5270) );
  AOI22_X1 U6456 ( .A1(n5268), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5267), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5269) );
  NAND4_X1 U6457 ( .A1(n5272), .A2(n5271), .A3(n5270), .A4(n5269), .ZN(n5283)
         );
  AOI22_X1 U6458 ( .A1(n5273), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n2986), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5281) );
  AOI22_X1 U6459 ( .A1(n4194), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5274), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5280) );
  AOI22_X1 U6460 ( .A1(n5275), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5279) );
  AOI22_X1 U6461 ( .A1(n5277), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n5276), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5278) );
  NAND4_X1 U6462 ( .A1(n5281), .A2(n5280), .A3(n5279), .A4(n5278), .ZN(n5282)
         );
  NOR2_X1 U6463 ( .A1(n5283), .A2(n5282), .ZN(n5287) );
  NOR2_X1 U6464 ( .A1(n5285), .A2(n5284), .ZN(n5286) );
  XOR2_X1 U6465 ( .A(n5287), .B(n5286), .Z(n5292) );
  AOI21_X1 U6466 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6534), .A(n5288), 
        .ZN(n5290) );
  NAND2_X1 U6467 ( .A1(n4204), .A2(EAX_REG_30__SCAN_IN), .ZN(n5289) );
  OAI211_X1 U6468 ( .C1(n5292), .C2(n5291), .A(n5290), .B(n5289), .ZN(n5293)
         );
  OAI21_X1 U6469 ( .B1(n5294), .B2(n5352), .A(n5293), .ZN(n5315) );
  AOI21_X1 U6470 ( .B1(n6076), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5295), 
        .ZN(n5296) );
  OAI21_X1 U6471 ( .B1(n6085), .B2(n5352), .A(n5296), .ZN(n5297) );
  AOI21_X1 U6472 ( .B1(n5346), .B2(n2983), .A(n5297), .ZN(n5298) );
  OAI21_X1 U6473 ( .B1(n5299), .B2(n6060), .A(n5298), .ZN(U2956) );
  XNOR2_X1 U6474 ( .A(n5517), .B(n5301), .ZN(n5569) );
  NOR2_X1 U6475 ( .A1(n5681), .A2(n5466), .ZN(n5303) );
  AOI211_X1 U6476 ( .C1(n6056), .C2(n5471), .A(n5304), .B(n5303), .ZN(n5305)
         );
  OAI211_X1 U6477 ( .C1(n5687), .C2(n5569), .A(n5306), .B(n5305), .ZN(U2963)
         );
  INV_X1 U6478 ( .A(n5308), .ZN(n5310) );
  INV_X1 U6479 ( .A(n5307), .ZN(n5309) );
  OAI21_X2 U6480 ( .B1(n5310), .B2(n5309), .A(n5421), .ZN(n5311) );
  INV_X1 U6481 ( .A(n5311), .ZN(n5609) );
  NAND2_X1 U6482 ( .A1(n5312), .A2(n5313), .ZN(n5314) );
  NAND2_X1 U6483 ( .A1(n5425), .A2(n5314), .ZN(n5740) );
  OAI222_X1 U6484 ( .A1(n5553), .A2(n5311), .B1(n5434), .B2(n6009), .C1(n5740), 
        .C2(n5549), .ZN(U2833) );
  AOI22_X1 U6485 ( .A1(n4204), .A2(EAX_REG_31__SCAN_IN), .B1(n5317), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5318) );
  XNOR2_X1 U6486 ( .A(n5319), .B(n5318), .ZN(n5388) );
  INV_X1 U6487 ( .A(n5388), .ZN(n5337) );
  NAND3_X1 U6488 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5321) );
  NAND4_X1 U6489 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(n5320), .ZN(n5834) );
  NOR2_X1 U6490 ( .A1(n5321), .A2(n5834), .ZN(n5322) );
  OR2_X1 U6491 ( .A1(n5322), .A2(n5483), .ZN(n5457) );
  INV_X1 U6492 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6683) );
  INV_X1 U6493 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6612) );
  INV_X1 U6494 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6658) );
  OR3_X1 U6495 ( .A1(n6683), .A2(n6612), .A3(n6658), .ZN(n5430) );
  NAND2_X1 U6496 ( .A1(n5835), .A2(n5430), .ZN(n5323) );
  NAND2_X1 U6497 ( .A1(n5457), .A2(n5323), .ZN(n5437) );
  INV_X1 U6498 ( .A(n5437), .ZN(n5326) );
  NAND2_X1 U6499 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5324) );
  NAND2_X1 U6500 ( .A1(n5991), .A2(n5324), .ZN(n5325) );
  NAND2_X1 U6501 ( .A1(n5326), .A2(n5325), .ZN(n5415) );
  AOI21_X1 U6502 ( .B1(n5991), .B2(n6738), .A(n5415), .ZN(n5357) );
  OAI21_X1 U6503 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5327), .A(n5357), .ZN(n5335) );
  NAND2_X1 U6504 ( .A1(n5956), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5330)
         );
  NAND3_X1 U6505 ( .A1(n5328), .A2(n6538), .A3(EBX_REG_31__SCAN_IN), .ZN(n5329) );
  OAI21_X1 U6506 ( .B1(n5331), .B2(n5938), .A(n3033), .ZN(n5334) );
  INV_X1 U6507 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6493) );
  NAND3_X1 U6508 ( .A1(n5925), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n5481) );
  NAND4_X1 U6509 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5852), .ZN(n5462) );
  INV_X1 U6510 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6667) );
  NOR3_X1 U6511 ( .A1(n5462), .A2(n6667), .A3(n5430), .ZN(n5416) );
  NAND2_X1 U6512 ( .A1(n5416), .A2(REIP_REG_28__SCAN_IN), .ZN(n5379) );
  NOR4_X1 U6513 ( .A1(n5379), .A2(REIP_REG_31__SCAN_IN), .A3(n6682), .A4(n6738), .ZN(n5333) );
  OAI21_X1 U6514 ( .B1(n5337), .B2(n5861), .A(n5336), .ZN(U2796) );
  AOI21_X1 U6515 ( .B1(n6522), .B2(n6399), .A(n5343), .ZN(n5345) );
  NOR2_X1 U6516 ( .A1(n5817), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5338)
         );
  AOI21_X1 U6517 ( .B1(n6330), .B2(n5339), .A(n5338), .ZN(n6401) );
  OAI21_X1 U6518 ( .B1(n6401), .B2(STATE2_REG_3__SCAN_IN), .A(n5340), .ZN(
        n5342) );
  AOI22_X1 U6519 ( .A1(n5342), .A2(n5341), .B1(n6521), .B2(n3205), .ZN(n5344)
         );
  OAI22_X1 U6520 ( .A1(n5345), .A2(n3205), .B1(n5344), .B2(n5343), .ZN(U3461)
         );
  AOI22_X1 U6521 ( .A1(n5349), .A2(n6005), .B1(EBX_REG_30__SCAN_IN), .B2(n5551), .ZN(n5347) );
  OAI21_X1 U6522 ( .B1(n5362), .B2(n5348), .A(n5347), .ZN(U2829) );
  NAND2_X1 U6523 ( .A1(n5349), .A2(n5987), .ZN(n5351) );
  AOI22_X1 U6524 ( .A1(n5956), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        EBX_REG_30__SCAN_IN), .B2(n5986), .ZN(n5350) );
  OAI211_X1 U6525 ( .C1(n5352), .C2(n5996), .A(n5351), .B(n5350), .ZN(n5353)
         );
  INV_X1 U6526 ( .A(n5353), .ZN(n5356) );
  NOR3_X1 U6527 ( .A1(n5379), .A2(REIP_REG_30__SCAN_IN), .A3(n6738), .ZN(n5354) );
  INV_X1 U6528 ( .A(n5354), .ZN(n5355) );
  INV_X1 U6529 ( .A(n5358), .ZN(n5359) );
  OAI21_X1 U6530 ( .B1(n5362), .B2(n5861), .A(n5359), .ZN(U2797) );
  AOI22_X1 U6531 ( .A1(n6010), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6013), .ZN(n5361) );
  NAND2_X1 U6532 ( .A1(n6014), .A2(DATAI_14_), .ZN(n5360) );
  OAI211_X1 U6533 ( .C1(n5362), .C2(n5583), .A(n5361), .B(n5360), .ZN(U2861)
         );
  AOI21_X1 U6534 ( .B1(n6076), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5363), 
        .ZN(n5364) );
  OAI21_X1 U6535 ( .B1(n6085), .B2(n5365), .A(n5364), .ZN(n5366) );
  AOI21_X1 U6536 ( .B1(n5388), .B2(n2983), .A(n5366), .ZN(n5367) );
  OAI21_X1 U6537 ( .B1(n5368), .B2(n6060), .A(n5367), .ZN(U2955) );
  INV_X1 U6538 ( .A(n5369), .ZN(n5375) );
  AOI21_X1 U6539 ( .B1(n5372), .B2(n5371), .A(n5370), .ZN(n5373) );
  NAND2_X1 U6540 ( .A1(n4248), .A2(n5373), .ZN(n5374) );
  NAND2_X1 U6541 ( .A1(n5375), .A2(n5374), .ZN(n5708) );
  AOI22_X1 U6542 ( .A1(n5956), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .B1(n5986), 
        .B2(EBX_REG_29__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U6543 ( .A1(n5968), .A2(n5376), .ZN(n5377) );
  OAI211_X1 U6544 ( .C1(n5708), .C2(n5938), .A(n5378), .B(n5377), .ZN(n5381)
         );
  NOR2_X1 U6545 ( .A1(n5379), .A2(REIP_REG_29__SCAN_IN), .ZN(n5380) );
  AOI211_X1 U6546 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5415), .A(n5381), .B(n5380), .ZN(n5382) );
  OAI21_X1 U6547 ( .B1(n5386), .B2(n5861), .A(n5382), .ZN(U2798) );
  AOI22_X1 U6548 ( .A1(n6010), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6013), .ZN(n5384) );
  NAND2_X1 U6549 ( .A1(n6014), .A2(DATAI_13_), .ZN(n5383) );
  OAI211_X1 U6550 ( .C1(n5386), .C2(n5583), .A(n5384), .B(n5383), .ZN(U2862)
         );
  OAI222_X1 U6551 ( .A1(n5553), .A2(n5386), .B1(n5385), .B2(n6009), .C1(n5708), 
        .C2(n5549), .ZN(U2830) );
  NAND3_X1 U6552 ( .A1(n5388), .A2(n5387), .A3(n5581), .ZN(n5390) );
  AOI22_X1 U6553 ( .A1(n6010), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6013), .ZN(n5389) );
  NAND2_X1 U6554 ( .A1(n5390), .A2(n5389), .ZN(U2860) );
  INV_X1 U6555 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6670) );
  NAND2_X1 U6556 ( .A1(n5391), .A2(n6670), .ZN(n5394) );
  INV_X1 U6557 ( .A(n5392), .ZN(n5393) );
  NOR2_X1 U6558 ( .A1(n5393), .A2(n3359), .ZN(n5405) );
  MUX2_X1 U6559 ( .A(n5394), .B(n5405), .S(n6538), .Z(U3474) );
  NAND3_X1 U6560 ( .A1(n5397), .A2(n5396), .A3(n5395), .ZN(n5398) );
  NAND2_X1 U6561 ( .A1(n5404), .A2(n5398), .ZN(n5402) );
  NAND2_X1 U6562 ( .A1(n5400), .A2(n5399), .ZN(n5401) );
  OAI211_X1 U6563 ( .C1(n5404), .C2(n5403), .A(n5402), .B(n5401), .ZN(n6416)
         );
  OAI21_X1 U6564 ( .B1(n5405), .B2(n6455), .A(n6638), .ZN(n6533) );
  NAND2_X1 U6565 ( .A1(n5406), .A2(n6533), .ZN(n6415) );
  AND2_X1 U6566 ( .A1(n6415), .A2(n6426), .ZN(n5911) );
  MUX2_X1 U6567 ( .A(MORE_REG_SCAN_IN), .B(n6416), .S(n5911), .Z(U3471) );
  INV_X1 U6568 ( .A(n5594), .ZN(n5556) );
  AND2_X1 U6569 ( .A1(n5427), .A2(n5409), .ZN(n5411) );
  OR2_X1 U6570 ( .A1(n5411), .A2(n5410), .ZN(n5720) );
  OAI22_X1 U6571 ( .A1(n5720), .A2(n5938), .B1(n5974), .B2(n5510), .ZN(n5414)
         );
  OAI22_X1 U6572 ( .A1(n5412), .A2(n5997), .B1(n5996), .B2(n5592), .ZN(n5413)
         );
  AOI211_X1 U6573 ( .C1(n5415), .C2(REIP_REG_28__SCAN_IN), .A(n5414), .B(n5413), .ZN(n5418) );
  INV_X1 U6574 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6614) );
  NAND2_X1 U6575 ( .A1(n5416), .A2(n6614), .ZN(n5417) );
  OAI211_X1 U6576 ( .C1(n5556), .C2(n5861), .A(n5418), .B(n5417), .ZN(U2799)
         );
  INV_X1 U6577 ( .A(n5419), .ZN(n5420) );
  INV_X1 U6578 ( .A(n5602), .ZN(n5559) );
  INV_X1 U6579 ( .A(n5423), .ZN(n5600) );
  NAND2_X1 U6580 ( .A1(n5425), .A2(n5424), .ZN(n5426) );
  AND2_X1 U6581 ( .A1(n5427), .A2(n5426), .ZN(n5733) );
  AOI22_X1 U6582 ( .A1(n5733), .A2(n5987), .B1(n5986), .B2(EBX_REG_27__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U6583 ( .A1(n5956), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5428)
         );
  OAI211_X1 U6584 ( .C1(n5996), .C2(n5600), .A(n5429), .B(n5428), .ZN(n5432)
         );
  NOR3_X1 U6585 ( .A1(n5462), .A2(REIP_REG_27__SCAN_IN), .A3(n5430), .ZN(n5431) );
  AOI211_X1 U6586 ( .C1(REIP_REG_27__SCAN_IN), .C2(n5437), .A(n5432), .B(n5431), .ZN(n5433) );
  OAI21_X1 U6587 ( .B1(n5559), .B2(n5861), .A(n5433), .ZN(U2800) );
  OAI22_X1 U6588 ( .A1(n5740), .A2(n5938), .B1(n5974), .B2(n5434), .ZN(n5436)
         );
  NOR2_X1 U6589 ( .A1(n5996), .A2(n5607), .ZN(n5435) );
  AOI211_X1 U6590 ( .C1(n5956), .C2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5436), 
        .B(n5435), .ZN(n5440) );
  NOR3_X1 U6591 ( .A1(n5462), .A2(n6683), .A3(n6658), .ZN(n5438) );
  OAI21_X1 U6592 ( .B1(n5438), .B2(REIP_REG_26__SCAN_IN), .A(n5437), .ZN(n5439) );
  OAI211_X1 U6593 ( .C1(n5311), .C2(n5861), .A(n5440), .B(n5439), .ZN(U2801)
         );
  OAI21_X1 U6594 ( .B1(n5441), .B2(n5442), .A(n5307), .ZN(n5564) );
  INV_X1 U6595 ( .A(n5564), .ZN(n5617) );
  XNOR2_X1 U6596 ( .A(REIP_REG_24__SCAN_IN), .B(REIP_REG_25__SCAN_IN), .ZN(
        n5443) );
  NOR2_X1 U6597 ( .A1(n5462), .A2(n5443), .ZN(n5451) );
  NAND2_X1 U6598 ( .A1(n5444), .A2(n5445), .ZN(n5446) );
  NAND2_X1 U6599 ( .A1(n5312), .A2(n5446), .ZN(n5748) );
  INV_X1 U6600 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5512) );
  OAI22_X1 U6601 ( .A1(n5748), .A2(n5938), .B1(n5974), .B2(n5512), .ZN(n5447)
         );
  AOI21_X1 U6602 ( .B1(n5956), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5447), 
        .ZN(n5449) );
  NAND2_X1 U6603 ( .A1(n5968), .A2(n5613), .ZN(n5448) );
  OAI211_X1 U6604 ( .C1(n5457), .C2(n6658), .A(n5449), .B(n5448), .ZN(n5450)
         );
  AOI211_X1 U6605 ( .C1(n5617), .C2(n5983), .A(n5451), .B(n5450), .ZN(n5452)
         );
  INV_X1 U6606 ( .A(n5452), .ZN(U2802) );
  NOR2_X1 U6607 ( .A1(n5455), .A2(n5454), .ZN(n5456) );
  OR2_X1 U6608 ( .A1(n5441), .A2(n5456), .ZN(n5623) );
  INV_X1 U6609 ( .A(n5457), .ZN(n5472) );
  OAI21_X1 U6610 ( .B1(n4224), .B2(n5458), .A(n5444), .ZN(n5758) );
  INV_X1 U6611 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5459) );
  OAI22_X1 U6612 ( .A1(n5758), .A2(n5938), .B1(n5459), .B2(n5974), .ZN(n5460)
         );
  AOI21_X1 U6613 ( .B1(n5956), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5460), 
        .ZN(n5461) );
  OAI21_X1 U6614 ( .B1(n5996), .B2(n5625), .A(n5461), .ZN(n5464) );
  NOR2_X1 U6615 ( .A1(n5462), .A2(REIP_REG_24__SCAN_IN), .ZN(n5463) );
  AOI211_X1 U6616 ( .C1(n5472), .C2(REIP_REG_24__SCAN_IN), .A(n5464), .B(n5463), .ZN(n5465) );
  OAI21_X1 U6617 ( .B1(n5623), .B2(n5861), .A(n5465), .ZN(U2803) );
  OAI22_X1 U6618 ( .A1(n5467), .A2(n5974), .B1(n5466), .B2(n5997), .ZN(n5470)
         );
  NOR2_X1 U6619 ( .A1(n5468), .A2(n5938), .ZN(n5469) );
  AOI211_X1 U6620 ( .C1(n5968), .C2(n5471), .A(n5470), .B(n5469), .ZN(n5475)
         );
  INV_X1 U6621 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6498) );
  NAND2_X1 U6622 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5852), .ZN(n5845) );
  OAI21_X1 U6623 ( .B1(n6498), .B2(n5845), .A(n3706), .ZN(n5473) );
  NAND2_X1 U6624 ( .A1(n5473), .A2(n5472), .ZN(n5474) );
  OAI211_X1 U6625 ( .C1(n5569), .C2(n5861), .A(n5475), .B(n5474), .ZN(U2804)
         );
  NOR2_X1 U6626 ( .A1(n5478), .A2(n5479), .ZN(n5480) );
  OR2_X1 U6627 ( .A1(n5524), .A2(n5480), .ZN(n5644) );
  NAND2_X1 U6628 ( .A1(n6493), .A2(n5481), .ZN(n5490) );
  INV_X1 U6629 ( .A(n5834), .ZN(n5482) );
  NOR2_X1 U6630 ( .A1(n5483), .A2(n5482), .ZN(n5846) );
  INV_X1 U6631 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5484) );
  OAI22_X1 U6632 ( .A1(n5484), .A2(n5997), .B1(n5646), .B2(n5996), .ZN(n5489)
         );
  MUX2_X1 U6633 ( .A(n5537), .B(n5535), .S(n5485), .Z(n5486) );
  XOR2_X1 U6634 ( .A(n5487), .B(n5486), .Z(n5782) );
  INV_X1 U6635 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5530) );
  OAI22_X1 U6636 ( .A1(n5782), .A2(n5938), .B1(n5530), .B2(n5974), .ZN(n5488)
         );
  AOI211_X1 U6637 ( .C1(n5490), .C2(n5846), .A(n5489), .B(n5488), .ZN(n5491)
         );
  OAI21_X1 U6638 ( .B1(n5644), .B2(n5861), .A(n5491), .ZN(U2807) );
  INV_X1 U6639 ( .A(n5492), .ZN(n5493) );
  AOI21_X1 U6640 ( .B1(n5495), .B2(n5494), .A(n5493), .ZN(n5705) );
  INV_X1 U6641 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5506) );
  AOI21_X1 U6642 ( .B1(n5497), .B2(n5496), .A(n5213), .ZN(n5887) );
  NAND2_X1 U6643 ( .A1(n5887), .A2(n5987), .ZN(n5501) );
  NAND2_X1 U6644 ( .A1(n5986), .A2(EBX_REG_15__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U6645 ( .A1(n5506), .A2(n5498), .ZN(n5499) );
  NAND4_X1 U6646 ( .A1(n5501), .A2(n6159), .A3(n5500), .A4(n5499), .ZN(n5502)
         );
  AOI21_X1 U6647 ( .B1(n5956), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5502), 
        .ZN(n5505) );
  INV_X1 U6648 ( .A(n5703), .ZN(n5503) );
  NAND2_X1 U6649 ( .A1(n5968), .A2(n5503), .ZN(n5504) );
  OAI211_X1 U6650 ( .C1(n5507), .C2(n5506), .A(n5505), .B(n5504), .ZN(n5508)
         );
  AOI21_X1 U6651 ( .B1(n5705), .B2(n5983), .A(n5508), .ZN(n5509) );
  INV_X1 U6652 ( .A(n5509), .ZN(U2812) );
  OAI222_X1 U6653 ( .A1(n5553), .A2(n5556), .B1(n5510), .B2(n6009), .C1(n5720), 
        .C2(n5549), .ZN(U2831) );
  AOI22_X1 U6654 ( .A1(n5733), .A2(n6005), .B1(EBX_REG_27__SCAN_IN), .B2(n5551), .ZN(n5511) );
  OAI21_X1 U6655 ( .B1(n5559), .B2(n5553), .A(n5511), .ZN(U2832) );
  OAI222_X1 U6656 ( .A1(n5564), .A2(n5553), .B1(n5512), .B2(n6009), .C1(n5748), 
        .C2(n5549), .ZN(U2834) );
  OAI222_X1 U6657 ( .A1(n5553), .A2(n5623), .B1(n6009), .B2(n5459), .C1(n5758), 
        .C2(n5549), .ZN(U2835) );
  AOI22_X1 U6658 ( .A1(n6005), .A2(n5513), .B1(n5551), .B2(EBX_REG_23__SCAN_IN), .ZN(n5514) );
  OAI21_X1 U6659 ( .B1(n5569), .B2(n5553), .A(n5514), .ZN(U2836) );
  INV_X1 U6660 ( .A(n5517), .ZN(n5518) );
  AOI21_X1 U6661 ( .B1(n5519), .B2(n5516), .A(n5518), .ZN(n5842) );
  INV_X1 U6662 ( .A(n5842), .ZN(n5572) );
  INV_X1 U6663 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5522) );
  OR2_X1 U6664 ( .A1(n5528), .A2(n5520), .ZN(n5521) );
  NAND2_X1 U6665 ( .A1(n3703), .A2(n5521), .ZN(n5836) );
  OAI222_X1 U6666 ( .A1(n5553), .A2(n5572), .B1(n6009), .B2(n5522), .C1(n5836), 
        .C2(n5549), .ZN(U2837) );
  OAI21_X1 U6667 ( .B1(n5524), .B2(n5523), .A(n5516), .ZN(n5848) );
  INV_X1 U6668 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5529) );
  NOR2_X1 U6669 ( .A1(n5526), .A2(n5525), .ZN(n5527) );
  OR2_X1 U6670 ( .A1(n5528), .A2(n5527), .ZN(n5849) );
  OAI222_X1 U6671 ( .A1(n5553), .A2(n5848), .B1(n5529), .B2(n6009), .C1(n5849), 
        .C2(n5549), .ZN(U2838) );
  OAI222_X1 U6672 ( .A1(n5549), .A2(n5782), .B1(n5530), .B2(n6009), .C1(n5644), 
        .C2(n5553), .ZN(U2839) );
  AND2_X1 U6673 ( .A1(n5543), .A2(n5532), .ZN(n5533) );
  NOR2_X1 U6674 ( .A1(n5478), .A2(n5533), .ZN(n5659) );
  INV_X1 U6675 ( .A(n5659), .ZN(n5862) );
  INV_X1 U6676 ( .A(n5534), .ZN(n5536) );
  MUX2_X1 U6677 ( .A(n5537), .B(n5536), .S(n5535), .Z(n5547) );
  INV_X1 U6678 ( .A(n5538), .ZN(n5548) );
  NAND2_X1 U6679 ( .A1(n5547), .A2(n5548), .ZN(n5546) );
  XNOR2_X1 U6680 ( .A(n5546), .B(n5539), .ZN(n5860) );
  INV_X1 U6681 ( .A(n5860), .ZN(n5540) );
  AOI22_X1 U6682 ( .A1(n6005), .A2(n5540), .B1(n5551), .B2(EBX_REG_19__SCAN_IN), .ZN(n5541) );
  OAI21_X1 U6683 ( .B1(n5862), .B2(n5553), .A(n5541), .ZN(U2840) );
  INV_X1 U6684 ( .A(n5236), .ZN(n5545) );
  INV_X1 U6685 ( .A(n5542), .ZN(n5544) );
  OAI21_X1 U6686 ( .B1(n5545), .B2(n5544), .A(n5543), .ZN(n5930) );
  OAI21_X1 U6687 ( .B1(n5548), .B2(n5547), .A(n5546), .ZN(n5795) );
  OAI222_X1 U6688 ( .A1(n5930), .A2(n5553), .B1(n5550), .B2(n6009), .C1(n5549), 
        .C2(n5795), .ZN(U2841) );
  INV_X1 U6689 ( .A(n5705), .ZN(n5584) );
  AOI22_X1 U6690 ( .A1(n6005), .A2(n5887), .B1(n5551), .B2(EBX_REG_15__SCAN_IN), .ZN(n5552) );
  OAI21_X1 U6691 ( .B1(n5584), .B2(n5553), .A(n5552), .ZN(U2844) );
  AOI22_X1 U6692 ( .A1(n6010), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6013), .ZN(n5555) );
  NAND2_X1 U6693 ( .A1(n6014), .A2(DATAI_12_), .ZN(n5554) );
  OAI211_X1 U6694 ( .C1(n5556), .C2(n5583), .A(n5555), .B(n5554), .ZN(U2863)
         );
  AOI22_X1 U6695 ( .A1(n6010), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6013), .ZN(n5558) );
  NAND2_X1 U6696 ( .A1(n6014), .A2(DATAI_11_), .ZN(n5557) );
  OAI211_X1 U6697 ( .C1(n5559), .C2(n5583), .A(n5558), .B(n5557), .ZN(U2864)
         );
  AOI22_X1 U6698 ( .A1(n6010), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6013), .ZN(n5561) );
  NAND2_X1 U6699 ( .A1(n6014), .A2(DATAI_10_), .ZN(n5560) );
  OAI211_X1 U6700 ( .C1(n5311), .C2(n5583), .A(n5561), .B(n5560), .ZN(U2865)
         );
  AOI22_X1 U6701 ( .A1(n6010), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6013), .ZN(n5563) );
  NAND2_X1 U6702 ( .A1(n6014), .A2(DATAI_9_), .ZN(n5562) );
  OAI211_X1 U6703 ( .C1(n5564), .C2(n5583), .A(n5563), .B(n5562), .ZN(U2866)
         );
  AOI22_X1 U6704 ( .A1(n6010), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6013), .ZN(n5566) );
  NAND2_X1 U6705 ( .A1(n6014), .A2(DATAI_8_), .ZN(n5565) );
  OAI211_X1 U6706 ( .C1(n5623), .C2(n5583), .A(n5566), .B(n5565), .ZN(U2867)
         );
  AOI22_X1 U6707 ( .A1(n6010), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6013), .ZN(n5568) );
  NAND2_X1 U6708 ( .A1(n6014), .A2(DATAI_7_), .ZN(n5567) );
  OAI211_X1 U6709 ( .C1(n5569), .C2(n5583), .A(n5568), .B(n5567), .ZN(U2868)
         );
  AOI22_X1 U6710 ( .A1(n6010), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n6013), .ZN(n5571) );
  NAND2_X1 U6711 ( .A1(n6014), .A2(DATAI_6_), .ZN(n5570) );
  OAI211_X1 U6712 ( .C1(n5572), .C2(n5583), .A(n5571), .B(n5570), .ZN(U2869)
         );
  AOI22_X1 U6713 ( .A1(n6010), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n6013), .ZN(n5574) );
  NAND2_X1 U6714 ( .A1(n6014), .A2(DATAI_5_), .ZN(n5573) );
  OAI211_X1 U6715 ( .C1(n5848), .C2(n5583), .A(n5574), .B(n5573), .ZN(U2870)
         );
  AOI22_X1 U6716 ( .A1(n6010), .A2(DATAI_20_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n6013), .ZN(n5576) );
  NAND2_X1 U6717 ( .A1(n6014), .A2(DATAI_4_), .ZN(n5575) );
  OAI211_X1 U6718 ( .C1(n5644), .C2(n5583), .A(n5576), .B(n5575), .ZN(U2871)
         );
  AOI22_X1 U6719 ( .A1(n6010), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6013), .ZN(n5578) );
  NAND2_X1 U6720 ( .A1(n6014), .A2(DATAI_3_), .ZN(n5577) );
  OAI211_X1 U6721 ( .C1(n5862), .C2(n5583), .A(n5578), .B(n5577), .ZN(U2872)
         );
  AOI22_X1 U6722 ( .A1(n6010), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n6013), .ZN(n5580) );
  NAND2_X1 U6723 ( .A1(n6014), .A2(DATAI_2_), .ZN(n5579) );
  OAI211_X1 U6724 ( .C1(n5930), .C2(n5583), .A(n5580), .B(n5579), .ZN(U2873)
         );
  OAI222_X1 U6725 ( .A1(n5584), .A2(n5583), .B1(n5582), .B2(n4396), .C1(n5581), 
        .C2(n6019), .ZN(U2876) );
  NAND3_X1 U6726 ( .A1(n5605), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n3477), .ZN(n5589) );
  NAND2_X1 U6727 ( .A1(n5586), .A2(n5750), .ZN(n5587) );
  OR2_X1 U6728 ( .A1(n5585), .A2(n5587), .ZN(n5596) );
  AOI22_X1 U6729 ( .A1(n5589), .A2(n5596), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5588), .ZN(n5590) );
  XNOR2_X1 U6730 ( .A(n5590), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5728)
         );
  NOR2_X1 U6731 ( .A1(n6159), .A2(n6614), .ZN(n5722) );
  AOI21_X1 U6732 ( .B1(n6076), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5722), 
        .ZN(n5591) );
  OAI21_X1 U6733 ( .B1(n6085), .B2(n5592), .A(n5591), .ZN(n5593) );
  AOI21_X1 U6734 ( .B1(n5594), .B2(n2983), .A(n5593), .ZN(n5595) );
  OAI21_X1 U6735 ( .B1(n6060), .B2(n5728), .A(n5595), .ZN(U2958) );
  NAND2_X1 U6736 ( .A1(n5597), .A2(n5596), .ZN(n5598) );
  XNOR2_X1 U6737 ( .A(n5598), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5737)
         );
  NOR2_X1 U6738 ( .A1(n6159), .A2(n6667), .ZN(n5732) );
  AOI21_X1 U6739 ( .B1(n6076), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5732), 
        .ZN(n5599) );
  OAI21_X1 U6740 ( .B1(n6085), .B2(n5600), .A(n5599), .ZN(n5601) );
  AOI21_X1 U6741 ( .B1(n5602), .B2(n2983), .A(n5601), .ZN(n5603) );
  OAI21_X1 U6742 ( .B1(n5737), .B2(n6060), .A(n5603), .ZN(U2959) );
  XNOR2_X1 U6743 ( .A(n3477), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5604)
         );
  XNOR2_X1 U6744 ( .A(n5605), .B(n5604), .ZN(n5745) );
  NOR2_X1 U6745 ( .A1(n6159), .A2(n6612), .ZN(n5738) );
  AOI21_X1 U6746 ( .B1(n6076), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5738), 
        .ZN(n5606) );
  OAI21_X1 U6747 ( .B1(n6085), .B2(n5607), .A(n5606), .ZN(n5608) );
  OAI21_X1 U6748 ( .B1(n6060), .B2(n5745), .A(n5610), .ZN(U2960) );
  AOI21_X1 U6749 ( .B1(n5612), .B2(n5585), .A(n5611), .ZN(n5754) );
  INV_X1 U6750 ( .A(n5613), .ZN(n5615) );
  NOR2_X1 U6751 ( .A1(n6159), .A2(n6658), .ZN(n5746) );
  AOI21_X1 U6752 ( .B1(n6076), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5746), 
        .ZN(n5614) );
  OAI21_X1 U6753 ( .B1(n6085), .B2(n5615), .A(n5614), .ZN(n5616) );
  AOI21_X1 U6754 ( .B1(n5617), .B2(n2983), .A(n5616), .ZN(n5618) );
  OAI21_X1 U6755 ( .B1(n5754), .B2(n6060), .A(n5618), .ZN(U2961) );
  INV_X1 U6756 ( .A(n5635), .ZN(n5619) );
  NAND3_X1 U6757 ( .A1(n3477), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5620) );
  XNOR2_X1 U6758 ( .A(n5622), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5763)
         );
  INV_X1 U6759 ( .A(n5623), .ZN(n5627) );
  NAND2_X1 U6760 ( .A1(n6185), .A2(REIP_REG_24__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U6761 ( .A1(n6076), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5624)
         );
  OAI211_X1 U6762 ( .C1(n6085), .C2(n5625), .A(n5757), .B(n5624), .ZN(n5626)
         );
  AOI21_X1 U6763 ( .B1(n5627), .B2(n2983), .A(n5626), .ZN(n5628) );
  OAI21_X1 U6764 ( .B1(n5763), .B2(n6060), .A(n5628), .ZN(U2962) );
  AOI21_X1 U6765 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n3477), .A(n5629), 
        .ZN(n5630) );
  XNOR2_X1 U6766 ( .A(n5631), .B(n5630), .ZN(n5770) );
  NAND2_X1 U6767 ( .A1(n6056), .A2(n5838), .ZN(n5632) );
  NAND2_X1 U6768 ( .A1(n6185), .A2(REIP_REG_22__SCAN_IN), .ZN(n5764) );
  OAI211_X1 U6769 ( .C1(n5681), .C2(n5840), .A(n5632), .B(n5764), .ZN(n5633)
         );
  AOI21_X1 U6770 ( .B1(n5842), .B2(n2983), .A(n5633), .ZN(n5634) );
  OAI21_X1 U6771 ( .B1(n5770), .B2(n6060), .A(n5634), .ZN(U2964) );
  AOI21_X1 U6772 ( .B1(n5637), .B2(n5636), .A(n5635), .ZN(n5771) );
  INV_X1 U6773 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5638) );
  INV_X1 U6774 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6496) );
  OR2_X1 U6775 ( .A1(n6159), .A2(n6496), .ZN(n5772) );
  OAI21_X1 U6776 ( .B1(n5681), .B2(n5638), .A(n5772), .ZN(n5640) );
  NOR2_X1 U6777 ( .A1(n5848), .A2(n5687), .ZN(n5639) );
  AOI211_X1 U6778 ( .C1(n6056), .C2(n5847), .A(n5640), .B(n5639), .ZN(n5641)
         );
  OAI21_X1 U6779 ( .B1(n5771), .B2(n6060), .A(n5641), .ZN(U2965) );
  XOR2_X1 U6780 ( .A(n5643), .B(n5642), .Z(n5785) );
  INV_X1 U6781 ( .A(n5644), .ZN(n5648) );
  NAND2_X1 U6782 ( .A1(n6185), .A2(REIP_REG_20__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U6783 ( .A1(n6076), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5645)
         );
  OAI211_X1 U6784 ( .C1(n6085), .C2(n5646), .A(n5780), .B(n5645), .ZN(n5647)
         );
  AOI21_X1 U6785 ( .B1(n5648), .B2(n2983), .A(n5647), .ZN(n5649) );
  OAI21_X1 U6786 ( .B1(n5785), .B2(n6060), .A(n5649), .ZN(U2966) );
  INV_X1 U6787 ( .A(n3000), .ZN(n5656) );
  INV_X1 U6788 ( .A(n5651), .ZN(n5652) );
  NOR2_X1 U6789 ( .A1(n5655), .A2(n5652), .ZN(n5654) );
  OAI22_X1 U6790 ( .A1(n5656), .A2(n5655), .B1(n5654), .B2(n5653), .ZN(n5793)
         );
  INV_X1 U6791 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5657) );
  NOR2_X1 U6792 ( .A1(n6159), .A2(n5657), .ZN(n5786) );
  NOR2_X1 U6793 ( .A1(n5681), .A2(n5859), .ZN(n5658) );
  AOI211_X1 U6794 ( .C1(n6056), .C2(n5857), .A(n5786), .B(n5658), .ZN(n5661)
         );
  NAND2_X1 U6795 ( .A1(n5659), .A2(n2983), .ZN(n5660) );
  OAI211_X1 U6796 ( .C1(n5793), .C2(n6060), .A(n5661), .B(n5660), .ZN(U2967)
         );
  NOR3_X1 U6797 ( .A1(n5671), .A2(n5672), .A3(n5796), .ZN(n5679) );
  OR2_X1 U6798 ( .A1(n5192), .A2(n5663), .ZN(n5665) );
  NAND2_X1 U6799 ( .A1(n5665), .A2(n5664), .ZN(n5699) );
  OR2_X1 U6800 ( .A1(n5699), .A2(n5698), .ZN(n5701) );
  NAND2_X1 U6801 ( .A1(n5672), .A2(n5796), .ZN(n5674) );
  NOR3_X1 U6802 ( .A1(n5701), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5674), 
        .ZN(n5676) );
  NOR2_X1 U6803 ( .A1(n5679), .A2(n5676), .ZN(n5666) );
  XNOR2_X1 U6804 ( .A(n5666), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5794)
         );
  NAND2_X1 U6805 ( .A1(n5794), .A2(n6081), .ZN(n5670) );
  INV_X1 U6806 ( .A(REIP_REG_18__SCAN_IN), .ZN(n5667) );
  NOR2_X1 U6807 ( .A1(n6159), .A2(n5667), .ZN(n5798) );
  NOR2_X1 U6808 ( .A1(n6085), .A2(n5928), .ZN(n5668) );
  AOI211_X1 U6809 ( .C1(n6076), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5798), 
        .B(n5668), .ZN(n5669) );
  OAI211_X1 U6810 ( .C1(n5687), .C2(n5930), .A(n5670), .B(n5669), .ZN(U2968)
         );
  INV_X1 U6811 ( .A(n5671), .ZN(n5675) );
  AOI21_X1 U6812 ( .B1(n5672), .B2(n3498), .A(n5796), .ZN(n5673) );
  AOI21_X1 U6813 ( .B1(n5675), .B2(n5674), .A(n5673), .ZN(n5678) );
  INV_X1 U6814 ( .A(n5676), .ZN(n5677) );
  OAI21_X1 U6815 ( .B1(n5679), .B2(n5678), .A(n5677), .ZN(n5875) );
  NAND2_X1 U6816 ( .A1(n5875), .A2(n6081), .ZN(n5685) );
  OAI22_X1 U6817 ( .A1(n5681), .A2(n5680), .B1(n6159), .B2(n6490), .ZN(n5682)
         );
  AOI21_X1 U6818 ( .B1(n6056), .B2(n5683), .A(n5682), .ZN(n5684) );
  OAI211_X1 U6819 ( .C1(n5687), .C2(n5686), .A(n5685), .B(n5684), .ZN(U2969)
         );
  OR2_X1 U6820 ( .A1(n5192), .A2(n5688), .ZN(n5690) );
  AND2_X1 U6821 ( .A1(n5690), .A2(n5689), .ZN(n5692) );
  MUX2_X1 U6822 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .B(n3498), .S(n3477), 
        .Z(n5691) );
  XNOR2_X1 U6823 ( .A(n5692), .B(n5691), .ZN(n5882) );
  INV_X1 U6824 ( .A(n5693), .ZN(n6012) );
  AOI22_X1 U6825 ( .A1(n6076), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6185), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5694) );
  OAI21_X1 U6826 ( .B1(n6085), .B2(n5695), .A(n5694), .ZN(n5696) );
  AOI21_X1 U6827 ( .B1(n6012), .B2(n2983), .A(n5696), .ZN(n5697) );
  OAI21_X1 U6828 ( .B1(n5882), .B2(n6060), .A(n5697), .ZN(U2970) );
  NAND2_X1 U6829 ( .A1(n5699), .A2(n5698), .ZN(n5700) );
  NAND2_X1 U6830 ( .A1(n5701), .A2(n5700), .ZN(n5891) );
  INV_X1 U6831 ( .A(n5891), .ZN(n5707) );
  AOI22_X1 U6832 ( .A1(n6076), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6185), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5702) );
  OAI21_X1 U6833 ( .B1(n6085), .B2(n5703), .A(n5702), .ZN(n5704) );
  AOI21_X1 U6834 ( .B1(n5705), .B2(n2983), .A(n5704), .ZN(n5706) );
  OAI21_X1 U6835 ( .B1(n5707), .B2(n6060), .A(n5706), .ZN(U2971) );
  INV_X1 U6836 ( .A(n5708), .ZN(n5710) );
  AOI21_X1 U6837 ( .B1(n5710), .B2(n6180), .A(n5709), .ZN(n5711) );
  OAI21_X1 U6838 ( .B1(n5712), .B2(n5714), .A(n5711), .ZN(n5713) );
  AOI21_X1 U6839 ( .B1(n5715), .B2(n5714), .A(n5713), .ZN(n5716) );
  OAI21_X1 U6840 ( .B1(n5717), .B2(n6157), .A(n5716), .ZN(U2989) );
  INV_X1 U6841 ( .A(n5718), .ZN(n5719) );
  AOI21_X1 U6842 ( .B1(n5719), .B2(n6136), .A(n5760), .ZN(n5730) );
  INV_X1 U6843 ( .A(n5730), .ZN(n5723) );
  NOR2_X1 U6844 ( .A1(n5720), .A2(n6160), .ZN(n5721) );
  AOI211_X1 U6845 ( .C1(n5723), .C2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5722), .B(n5721), .ZN(n5727) );
  OR3_X1 U6846 ( .A1(n5734), .A2(n5725), .A3(n5724), .ZN(n5726) );
  OAI211_X1 U6847 ( .C1(n5728), .C2(n6157), .A(n5727), .B(n5726), .ZN(U2990)
         );
  INV_X1 U6848 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5729) );
  NOR2_X1 U6849 ( .A1(n5730), .A2(n5729), .ZN(n5731) );
  AOI211_X1 U6850 ( .C1(n6180), .C2(n5733), .A(n5732), .B(n5731), .ZN(n5736)
         );
  OR2_X1 U6851 ( .A1(n5734), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5735)
         );
  OAI211_X1 U6852 ( .C1(n5737), .C2(n6157), .A(n5736), .B(n5735), .ZN(U2991)
         );
  INV_X1 U6853 ( .A(n5738), .ZN(n5739) );
  OAI21_X1 U6854 ( .B1(n6160), .B2(n5740), .A(n5739), .ZN(n5741) );
  AOI21_X1 U6855 ( .B1(n5760), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5741), 
        .ZN(n5744) );
  XNOR2_X1 U6856 ( .A(n5750), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5742)
         );
  NAND2_X1 U6857 ( .A1(n5751), .A2(n5742), .ZN(n5743) );
  OAI211_X1 U6858 ( .C1(n5745), .C2(n6157), .A(n5744), .B(n5743), .ZN(U2992)
         );
  INV_X1 U6859 ( .A(n5746), .ZN(n5747) );
  OAI21_X1 U6860 ( .B1(n6160), .B2(n5748), .A(n5747), .ZN(n5749) );
  AOI21_X1 U6861 ( .B1(n5760), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5749), 
        .ZN(n5753) );
  NAND2_X1 U6862 ( .A1(n5751), .A2(n5750), .ZN(n5752) );
  OAI211_X1 U6863 ( .C1(n5754), .C2(n6157), .A(n5753), .B(n5752), .ZN(U2993)
         );
  INV_X1 U6864 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5755) );
  OAI21_X1 U6865 ( .B1(n5756), .B2(n3503), .A(n5755), .ZN(n5761) );
  OAI21_X1 U6866 ( .B1(n6160), .B2(n5758), .A(n5757), .ZN(n5759) );
  AOI21_X1 U6867 ( .B1(n5761), .B2(n5760), .A(n5759), .ZN(n5762) );
  OAI21_X1 U6868 ( .B1(n5763), .B2(n6157), .A(n5762), .ZN(U2994) );
  OAI21_X1 U6869 ( .B1(n6160), .B2(n5836), .A(n5764), .ZN(n5768) );
  NOR3_X1 U6870 ( .A1(n5777), .A2(n5766), .A3(n5765), .ZN(n5767) );
  AOI211_X1 U6871 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5774), .A(n5768), .B(n5767), .ZN(n5769) );
  OAI21_X1 U6872 ( .B1(n5770), .B2(n6157), .A(n5769), .ZN(U2996) );
  OR2_X1 U6873 ( .A1(n5771), .A2(n6157), .ZN(n5776) );
  OAI21_X1 U6874 ( .B1(n6160), .B2(n5849), .A(n5772), .ZN(n5773) );
  AOI21_X1 U6875 ( .B1(n5774), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5773), 
        .ZN(n5775) );
  OAI211_X1 U6876 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5777), .A(n5776), .B(n5775), .ZN(U2997) );
  AOI21_X1 U6877 ( .B1(n5796), .B2(n5778), .A(n5873), .ZN(n5802) );
  OAI21_X1 U6878 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6102), .A(n5802), 
        .ZN(n5790) );
  XNOR2_X1 U6879 ( .A(n5788), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5779)
         );
  NAND2_X1 U6880 ( .A1(n5789), .A2(n5779), .ZN(n5781) );
  OAI211_X1 U6881 ( .C1(n6160), .C2(n5782), .A(n5781), .B(n5780), .ZN(n5783)
         );
  AOI21_X1 U6882 ( .B1(n5790), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5783), 
        .ZN(n5784) );
  OAI21_X1 U6883 ( .B1(n5785), .B2(n6157), .A(n5784), .ZN(U2998) );
  NOR2_X1 U6884 ( .A1(n6160), .A2(n5860), .ZN(n5787) );
  AOI211_X1 U6885 ( .C1(n5789), .C2(n5788), .A(n5787), .B(n5786), .ZN(n5792)
         );
  NAND2_X1 U6886 ( .A1(n5790), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5791) );
  OAI211_X1 U6887 ( .C1(n5793), .C2(n6157), .A(n5792), .B(n5791), .ZN(U2999)
         );
  NAND2_X1 U6888 ( .A1(n5794), .A2(n6183), .ZN(n5800) );
  INV_X1 U6889 ( .A(n5795), .ZN(n5931) );
  NOR3_X1 U6890 ( .A1(n5878), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n5796), 
        .ZN(n5797) );
  AOI211_X1 U6891 ( .C1(n6180), .C2(n5931), .A(n5798), .B(n5797), .ZN(n5799)
         );
  OAI211_X1 U6892 ( .C1(n5802), .C2(n5801), .A(n5800), .B(n5799), .ZN(U3000)
         );
  AND2_X1 U6893 ( .A1(n4472), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6193) );
  INV_X1 U6894 ( .A(n6193), .ZN(n6328) );
  OAI211_X1 U6895 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4472), .A(n6328), .B(
        n6327), .ZN(n5803) );
  OAI21_X1 U6896 ( .B1(n5812), .B2(n5824), .A(n5803), .ZN(n5804) );
  MUX2_X1 U6897 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5804), .S(n6191), 
        .Z(U3464) );
  XNOR2_X1 U6898 ( .A(n5805), .B(n6193), .ZN(n5808) );
  INV_X1 U6899 ( .A(n5806), .ZN(n5807) );
  OAI22_X1 U6900 ( .A1(n5808), .A2(n6332), .B1(n5807), .B2(n5812), .ZN(n5809)
         );
  MUX2_X1 U6901 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5809), .S(n6191), 
        .Z(U3463) );
  INV_X1 U6902 ( .A(n5810), .ZN(n5814) );
  NAND2_X1 U6903 ( .A1(n5811), .A2(n6329), .ZN(n6196) );
  NOR2_X1 U6904 ( .A1(n6234), .A2(n6328), .ZN(n6274) );
  NOR2_X1 U6905 ( .A1(n6196), .A2(n6274), .ZN(n5813) );
  OAI222_X1 U6906 ( .A1(n5815), .A2(n5814), .B1(n6332), .B2(n5813), .C1(n5812), 
        .C2(n5993), .ZN(n5816) );
  MUX2_X1 U6907 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5816), .S(n6191), 
        .Z(U3462) );
  INV_X1 U6908 ( .A(n5817), .ZN(n5820) );
  INV_X1 U6909 ( .A(n5818), .ZN(n5819) );
  INV_X1 U6910 ( .A(n4433), .ZN(n5827) );
  NAND3_X1 U6911 ( .A1(n5820), .A2(n5819), .A3(n5827), .ZN(n5821) );
  OAI211_X1 U6912 ( .C1(n5824), .C2(n5823), .A(n5822), .B(n5821), .ZN(n6405)
         );
  INV_X1 U6913 ( .A(n6405), .ZN(n5831) );
  INV_X1 U6914 ( .A(n6522), .ZN(n5830) );
  AOI22_X1 U6915 ( .A1(n5828), .A2(n5827), .B1(n5826), .B2(n5825), .ZN(n5829)
         );
  OAI21_X1 U6916 ( .B1(n5831), .B2(n5830), .A(n5829), .ZN(n5832) );
  MUX2_X1 U6917 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n5832), .S(n6525), 
        .Z(U3460) );
  AND2_X1 U6918 ( .A1(n6038), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6919 ( .A1(n5852), .A2(n6496), .B1(n5835), .B2(n5834), .ZN(n5844)
         );
  OAI22_X1 U6920 ( .A1(n5836), .A2(n5938), .B1(n5522), .B2(n5974), .ZN(n5837)
         );
  AOI21_X1 U6921 ( .B1(n5968), .B2(n5838), .A(n5837), .ZN(n5839) );
  OAI21_X1 U6922 ( .B1(n5997), .B2(n5840), .A(n5839), .ZN(n5841) );
  AOI21_X1 U6923 ( .B1(n5842), .B2(n5983), .A(n5841), .ZN(n5843) );
  OAI221_X1 U6924 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5845), .C1(n6498), .C2(
        n5844), .A(n5843), .ZN(U2805) );
  AOI22_X1 U6925 ( .A1(EBX_REG_21__SCAN_IN), .A2(n5986), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n5956), .ZN(n5856) );
  AOI22_X1 U6926 ( .A1(n5847), .A2(n5968), .B1(REIP_REG_21__SCAN_IN), .B2(
        n5846), .ZN(n5855) );
  INV_X1 U6927 ( .A(n5848), .ZN(n5851) );
  INV_X1 U6928 ( .A(n5849), .ZN(n5850) );
  AOI22_X1 U6929 ( .A1(n5851), .A2(n5983), .B1(n5987), .B2(n5850), .ZN(n5854)
         );
  NAND2_X1 U6930 ( .A1(n5852), .A2(n6496), .ZN(n5853) );
  NAND4_X1 U6931 ( .A1(n5856), .A2(n5855), .A3(n5854), .A4(n5853), .ZN(U2806)
         );
  AOI22_X1 U6932 ( .A1(n5857), .A2(n5968), .B1(REIP_REG_19__SCAN_IN), .B2(
        n5926), .ZN(n5858) );
  OAI211_X1 U6933 ( .C1(n5997), .C2(n5859), .A(n5858), .B(n6159), .ZN(n5864)
         );
  OAI22_X1 U6934 ( .A1(n5862), .A2(n5861), .B1(n5860), .B2(n5938), .ZN(n5863)
         );
  AOI211_X1 U6935 ( .C1(EBX_REG_19__SCAN_IN), .C2(n5986), .A(n5864), .B(n5863), 
        .ZN(n5867) );
  NAND2_X1 U6936 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5865) );
  OAI211_X1 U6937 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n5925), .B(n5865), .ZN(n5866) );
  NAND2_X1 U6938 ( .A1(n5867), .A2(n5866), .ZN(U2808) );
  AOI22_X1 U6939 ( .A1(n6185), .A2(REIP_REG_13__SCAN_IN), .B1(n6076), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5872) );
  XNOR2_X1 U6940 ( .A(n5868), .B(n5869), .ZN(n5897) );
  INV_X1 U6941 ( .A(n5870), .ZN(n5945) );
  AOI22_X1 U6942 ( .A1(n5897), .A2(n6081), .B1(n2983), .B2(n5945), .ZN(n5871)
         );
  OAI211_X1 U6943 ( .C1(n6085), .C2(n5939), .A(n5872), .B(n5871), .ZN(U2973)
         );
  AOI22_X1 U6944 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5873), .B1(n6185), .B2(REIP_REG_17__SCAN_IN), .ZN(n5877) );
  AOI22_X1 U6945 ( .A1(n5875), .A2(n6183), .B1(n6180), .B2(n5874), .ZN(n5876)
         );
  OAI211_X1 U6946 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5878), .A(n5877), .B(n5876), .ZN(U3001) );
  INV_X1 U6947 ( .A(n5879), .ZN(n5889) );
  AOI211_X1 U6948 ( .C1(n5893), .C2(n3498), .A(n5880), .B(n5889), .ZN(n5884)
         );
  OAI22_X1 U6949 ( .A1(n5882), .A2(n6157), .B1(n6160), .B2(n5881), .ZN(n5883)
         );
  NOR2_X1 U6950 ( .A1(n5884), .A2(n5883), .ZN(n5886) );
  NAND2_X1 U6951 ( .A1(n6185), .A2(REIP_REG_16__SCAN_IN), .ZN(n5885) );
  OAI211_X1 U6952 ( .C1(n5894), .C2(n3498), .A(n5886), .B(n5885), .ZN(U3002)
         );
  AOI22_X1 U6953 ( .A1(n6180), .A2(n5887), .B1(n6185), .B2(
        REIP_REG_15__SCAN_IN), .ZN(n5888) );
  OAI21_X1 U6954 ( .B1(n5889), .B2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5888), 
        .ZN(n5890) );
  AOI21_X1 U6955 ( .B1(n5891), .B2(n6183), .A(n5890), .ZN(n5892) );
  OAI21_X1 U6956 ( .B1(n5894), .B2(n5893), .A(n5892), .ZN(U3003) );
  OR2_X1 U6957 ( .A1(n5895), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5900)
         );
  AOI22_X1 U6958 ( .A1(n6180), .A2(n5936), .B1(n6185), .B2(
        REIP_REG_13__SCAN_IN), .ZN(n5899) );
  AOI22_X1 U6959 ( .A1(n5897), .A2(n6183), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5896), .ZN(n5898) );
  OAI211_X1 U6960 ( .C1(n5901), .C2(n5900), .A(n5899), .B(n5898), .ZN(U3005)
         );
  INV_X1 U6961 ( .A(n5902), .ZN(n5906) );
  INV_X1 U6962 ( .A(n5903), .ZN(n5905) );
  NAND4_X1 U6963 ( .A1(n5906), .A2(n5905), .A3(n6522), .A4(n5904), .ZN(n5907)
         );
  OAI21_X1 U6964 ( .B1(n6525), .B2(n5908), .A(n5907), .ZN(U3455) );
  INV_X1 U6965 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6461) );
  NOR2_X1 U6966 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6461), .ZN(n6739) );
  INV_X1 U6967 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6562) );
  AOI221_X1 U6968 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_0__SCAN_IN), .C1(
        n6461), .C2(STATE_REG_0__SCAN_IN), .A(n6739), .ZN(n6515) );
  INV_X1 U6969 ( .A(n6515), .ZN(n6448) );
  OAI21_X1 U6970 ( .B1(n6739), .B2(n6562), .A(n6448), .ZN(U2789) );
  INV_X1 U6971 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6665) );
  NOR2_X1 U6972 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5910) );
  NOR2_X1 U6973 ( .A1(n6739), .A2(n5910), .ZN(n5909) );
  AOI22_X1 U6974 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n6739), .B1(n6665), .B2(
        n5909), .ZN(U2791) );
  OAI21_X1 U6975 ( .B1(BS16_N), .B2(n5910), .A(n6515), .ZN(n6513) );
  OAI21_X1 U6976 ( .B1(n6515), .B2(n6604), .A(n6513), .ZN(U2792) );
  OAI21_X1 U6977 ( .B1(n5911), .B2(n6551), .A(n6060), .ZN(U2793) );
  NOR4_X1 U6978 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5915) );
  NOR4_X1 U6979 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n5914) );
  NOR4_X1 U6980 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5913) );
  NOR4_X1 U6981 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5912) );
  NAND4_X1 U6982 ( .A1(n5915), .A2(n5914), .A3(n5913), .A4(n5912), .ZN(n5921)
         );
  NOR4_X1 U6983 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n5919) );
  AOI211_X1 U6984 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_2__SCAN_IN), .B(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n5918) );
  NOR4_X1 U6985 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n5917) );
  NOR4_X1 U6986 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n5916) );
  NAND4_X1 U6987 ( .A1(n5919), .A2(n5918), .A3(n5917), .A4(n5916), .ZN(n5920)
         );
  NOR2_X1 U6988 ( .A1(n5921), .A2(n5920), .ZN(n6532) );
  INV_X1 U6989 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6640) );
  NOR3_X1 U6990 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5923) );
  OAI21_X1 U6991 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5923), .A(n6532), .ZN(n5922)
         );
  OAI21_X1 U6992 ( .B1(n6532), .B2(n6640), .A(n5922), .ZN(U2794) );
  INV_X1 U6993 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6514) );
  AOI21_X1 U6994 ( .B1(n6527), .B2(n6514), .A(n5923), .ZN(n5924) );
  INV_X1 U6995 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6603) );
  INV_X1 U6996 ( .A(n6532), .ZN(n6529) );
  AOI22_X1 U6997 ( .A1(n6532), .A2(n5924), .B1(n6603), .B2(n6529), .ZN(U2795)
         );
  INV_X1 U6998 ( .A(n5925), .ZN(n5935) );
  AOI22_X1 U6999 ( .A1(EBX_REG_18__SCAN_IN), .A2(n5986), .B1(
        REIP_REG_18__SCAN_IN), .B2(n5926), .ZN(n5927) );
  OAI21_X1 U7000 ( .B1(n5928), .B2(n5996), .A(n5927), .ZN(n5929) );
  AOI211_X1 U7001 ( .C1(n5956), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6185), 
        .B(n5929), .ZN(n5934) );
  INV_X1 U7002 ( .A(n5930), .ZN(n5932) );
  AOI22_X1 U7003 ( .A1(n5932), .A2(n5983), .B1(n5987), .B2(n5931), .ZN(n5933)
         );
  OAI211_X1 U7004 ( .C1(REIP_REG_18__SCAN_IN), .C2(n5935), .A(n5934), .B(n5933), .ZN(U2809) );
  INV_X1 U7005 ( .A(n5936), .ZN(n5937) );
  OAI22_X1 U7006 ( .A1(n5996), .A2(n5939), .B1(n5938), .B2(n5937), .ZN(n5940)
         );
  AOI211_X1 U7007 ( .C1(n5956), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6185), 
        .B(n5940), .ZN(n5947) );
  INV_X1 U7008 ( .A(n5949), .ZN(n5972) );
  NOR3_X1 U7009 ( .A1(REIP_REG_13__SCAN_IN), .A2(n5941), .A3(n5972), .ZN(n5944) );
  AOI21_X1 U7010 ( .B1(n5953), .B2(n5942), .A(n6482), .ZN(n5943) );
  AOI211_X1 U7011 ( .C1(n5945), .C2(n5983), .A(n5944), .B(n5943), .ZN(n5946)
         );
  OAI211_X1 U7012 ( .C1(n5948), .C2(n5974), .A(n5947), .B(n5946), .ZN(U2814)
         );
  NAND2_X1 U7013 ( .A1(n5949), .A2(n6480), .ZN(n5960) );
  AOI21_X1 U7014 ( .B1(n5951), .B2(n5950), .A(n5078), .ZN(n6086) );
  NAND2_X1 U7015 ( .A1(n6086), .A2(n5987), .ZN(n5952) );
  OAI211_X1 U7016 ( .C1(n6008), .C2(n5974), .A(n5952), .B(n6159), .ZN(n5955)
         );
  NOR2_X1 U7017 ( .A1(n5953), .A2(n6480), .ZN(n5954) );
  AOI211_X1 U7018 ( .C1(n5956), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n5955), 
        .B(n5954), .ZN(n5959) );
  INV_X1 U7019 ( .A(n5957), .ZN(n6057) );
  AOI22_X1 U7020 ( .A1(n6057), .A2(n5983), .B1(n5968), .B2(n6055), .ZN(n5958)
         );
  OAI211_X1 U7021 ( .C1(n5961), .C2(n5960), .A(n5959), .B(n5958), .ZN(U2816)
         );
  AOI22_X1 U7022 ( .A1(n6109), .A2(n5987), .B1(n5986), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n5962) );
  OAI211_X1 U7023 ( .C1(n5997), .C2(n5963), .A(n5962), .B(n6159), .ZN(n5964)
         );
  AOI21_X1 U7024 ( .B1(REIP_REG_9__SCAN_IN), .B2(n5965), .A(n5964), .ZN(n5971)
         );
  INV_X1 U7025 ( .A(n5966), .ZN(n5969) );
  AOI22_X1 U7026 ( .A1(n5969), .A2(n5983), .B1(n5968), .B2(n5967), .ZN(n5970)
         );
  OAI211_X1 U7027 ( .C1(REIP_REG_9__SCAN_IN), .C2(n5972), .A(n5971), .B(n5970), 
        .ZN(U2818) );
  INV_X1 U7028 ( .A(n6138), .ZN(n5976) );
  OAI21_X1 U7029 ( .B1(n5974), .B2(n5973), .A(n6159), .ZN(n5975) );
  AOI21_X1 U7030 ( .B1(n5987), .B2(n5976), .A(n5975), .ZN(n5977) );
  OAI21_X1 U7031 ( .B1(n5997), .B2(n5978), .A(n5977), .ZN(n5979) );
  AOI221_X1 U7032 ( .B1(n5981), .B2(n6137), .C1(n5980), .C2(
        REIP_REG_6__SCAN_IN), .A(n5979), .ZN(n5985) );
  INV_X1 U7033 ( .A(n5982), .ZN(n6065) );
  NAND2_X1 U7034 ( .A1(n6065), .A2(n5983), .ZN(n5984) );
  OAI211_X1 U7035 ( .C1(n5996), .C2(n6068), .A(n5985), .B(n5984), .ZN(U2821)
         );
  INV_X1 U7036 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6467) );
  AOI22_X1 U7037 ( .A1(n6169), .A2(n5987), .B1(n5986), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n6003) );
  INV_X1 U7038 ( .A(n5988), .ZN(n6072) );
  INV_X1 U7039 ( .A(n5989), .ZN(n6001) );
  NAND2_X1 U7040 ( .A1(n5991), .A2(n5990), .ZN(n5994) );
  OAI22_X1 U7041 ( .A1(n5995), .A2(n5994), .B1(n5993), .B2(n5992), .ZN(n6000)
         );
  INV_X1 U7042 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5998) );
  OAI22_X1 U7043 ( .A1(n5998), .A2(n5997), .B1(n5996), .B2(n6075), .ZN(n5999)
         );
  AOI211_X1 U7044 ( .C1(n6072), .C2(n6001), .A(n6000), .B(n5999), .ZN(n6002)
         );
  OAI211_X1 U7045 ( .C1(n6004), .C2(n6467), .A(n6003), .B(n6002), .ZN(U2824)
         );
  AOI22_X1 U7046 ( .A1(n6057), .A2(n6006), .B1(n6005), .B2(n6086), .ZN(n6007)
         );
  OAI21_X1 U7047 ( .B1(n6009), .B2(n6008), .A(n6007), .ZN(U2848) );
  AOI22_X1 U7048 ( .A1(n6012), .A2(n6011), .B1(n6010), .B2(DATAI_16_), .ZN(
        n6016) );
  AOI22_X1 U7049 ( .A1(n6014), .A2(DATAI_0_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n6013), .ZN(n6015) );
  NAND2_X1 U7050 ( .A1(n6016), .A2(n6015), .ZN(U2875) );
  AOI22_X1 U7051 ( .A1(n6425), .A2(LWORD_REG_15__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6018) );
  OAI21_X1 U7052 ( .B1(n6019), .B2(n6049), .A(n6018), .ZN(U2908) );
  AOI22_X1 U7053 ( .A1(n6425), .A2(LWORD_REG_14__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6020) );
  OAI21_X1 U7054 ( .B1(n6021), .B2(n6049), .A(n6020), .ZN(U2909) );
  AOI22_X1 U7055 ( .A1(n6425), .A2(LWORD_REG_13__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6022) );
  OAI21_X1 U7056 ( .B1(n6023), .B2(n6049), .A(n6022), .ZN(U2910) );
  AOI22_X1 U7057 ( .A1(n6425), .A2(LWORD_REG_12__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6024) );
  OAI21_X1 U7058 ( .B1(n6025), .B2(n6049), .A(n6024), .ZN(U2911) );
  AOI22_X1 U7059 ( .A1(n6425), .A2(LWORD_REG_11__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6026) );
  OAI21_X1 U7060 ( .B1(n6027), .B2(n6049), .A(n6026), .ZN(U2912) );
  AOI22_X1 U7061 ( .A1(n6425), .A2(LWORD_REG_10__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6028) );
  OAI21_X1 U7062 ( .B1(n6029), .B2(n6049), .A(n6028), .ZN(U2913) );
  AOI22_X1 U7063 ( .A1(n6425), .A2(LWORD_REG_9__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6030) );
  OAI21_X1 U7064 ( .B1(n6031), .B2(n6049), .A(n6030), .ZN(U2914) );
  AOI22_X1 U7065 ( .A1(n6425), .A2(LWORD_REG_8__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6032) );
  OAI21_X1 U7066 ( .B1(n6033), .B2(n6049), .A(n6032), .ZN(U2915) );
  AOI22_X1 U7067 ( .A1(n6425), .A2(LWORD_REG_7__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6034) );
  OAI21_X1 U7068 ( .B1(n3801), .B2(n6049), .A(n6034), .ZN(U2916) );
  AOI22_X1 U7069 ( .A1(n6425), .A2(LWORD_REG_6__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6035) );
  OAI21_X1 U7070 ( .B1(n6036), .B2(n6049), .A(n6035), .ZN(U2917) );
  AOI22_X1 U7071 ( .A1(n6425), .A2(LWORD_REG_5__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6037) );
  OAI21_X1 U7072 ( .B1(n3789), .B2(n6049), .A(n6037), .ZN(U2918) );
  AOI22_X1 U7073 ( .A1(n6425), .A2(LWORD_REG_4__SCAN_IN), .B1(n6038), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6039) );
  OAI21_X1 U7074 ( .B1(n6040), .B2(n6049), .A(n6039), .ZN(U2919) );
  AOI22_X1 U7075 ( .A1(n6425), .A2(LWORD_REG_3__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6041) );
  OAI21_X1 U7076 ( .B1(n6042), .B2(n6049), .A(n6041), .ZN(U2920) );
  AOI22_X1 U7077 ( .A1(n6425), .A2(LWORD_REG_2__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6043) );
  OAI21_X1 U7078 ( .B1(n6044), .B2(n6049), .A(n6043), .ZN(U2921) );
  AOI22_X1 U7079 ( .A1(n6425), .A2(LWORD_REG_1__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6045) );
  OAI21_X1 U7080 ( .B1(n6046), .B2(n6049), .A(n6045), .ZN(U2922) );
  AOI22_X1 U7081 ( .A1(n6425), .A2(LWORD_REG_0__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6048) );
  OAI21_X1 U7082 ( .B1(n6050), .B2(n6049), .A(n6048), .ZN(U2923) );
  NAND2_X1 U7083 ( .A1(n3017), .A2(n6051), .ZN(n6054) );
  XNOR2_X1 U7084 ( .A(n3477), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6053)
         );
  XNOR2_X1 U7085 ( .A(n6054), .B(n6053), .ZN(n6091) );
  AOI22_X1 U7086 ( .A1(n6185), .A2(REIP_REG_11__SCAN_IN), .B1(n6076), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6059) );
  AOI22_X1 U7087 ( .A1(n6057), .A2(n2983), .B1(n6056), .B2(n6055), .ZN(n6058)
         );
  OAI211_X1 U7088 ( .C1(n6091), .C2(n6060), .A(n6059), .B(n6058), .ZN(U2975)
         );
  AOI22_X1 U7089 ( .A1(n6185), .A2(REIP_REG_6__SCAN_IN), .B1(n6076), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6067) );
  OAI21_X1 U7090 ( .B1(n6063), .B2(n6062), .A(n3016), .ZN(n6064) );
  INV_X1 U7091 ( .A(n6064), .ZN(n6141) );
  AOI22_X1 U7092 ( .A1(n6141), .A2(n6081), .B1(n2983), .B2(n6065), .ZN(n6066)
         );
  OAI211_X1 U7093 ( .C1(n6085), .C2(n6068), .A(n6067), .B(n6066), .ZN(U2980)
         );
  AOI22_X1 U7094 ( .A1(n6185), .A2(REIP_REG_3__SCAN_IN), .B1(n6076), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6074) );
  OAI21_X1 U7095 ( .B1(n6070), .B2(n6069), .A(n4960), .ZN(n6071) );
  INV_X1 U7096 ( .A(n6071), .ZN(n6170) );
  AOI22_X1 U7097 ( .A1(n6081), .A2(n6170), .B1(n6072), .B2(n2983), .ZN(n6073)
         );
  OAI211_X1 U7098 ( .C1(n6085), .C2(n6075), .A(n6074), .B(n6073), .ZN(U2983)
         );
  AOI22_X1 U7099 ( .A1(n6185), .A2(REIP_REG_2__SCAN_IN), .B1(n6076), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6083) );
  XOR2_X1 U7100 ( .A(n6077), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n6079) );
  XNOR2_X1 U7101 ( .A(n6079), .B(n6078), .ZN(n6184) );
  AOI22_X1 U7102 ( .A1(n6184), .A2(n6081), .B1(n6080), .B2(n2983), .ZN(n6082)
         );
  OAI211_X1 U7103 ( .C1(n6085), .C2(n6084), .A(n6083), .B(n6082), .ZN(U2984)
         );
  AOI22_X1 U7104 ( .A1(n6180), .A2(n6086), .B1(n6185), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n6090) );
  AOI22_X1 U7105 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6088), .B1(n6087), .B2(n3485), .ZN(n6089) );
  OAI211_X1 U7106 ( .C1(n6091), .C2(n6157), .A(n6090), .B(n6089), .ZN(U3007)
         );
  AOI21_X1 U7107 ( .B1(n6133), .B2(n6186), .A(n6179), .ZN(n6163) );
  NOR2_X1 U7108 ( .A1(n6092), .A2(n6163), .ZN(n6126) );
  NAND2_X1 U7109 ( .A1(n6101), .A2(n6126), .ZN(n6114) );
  AOI22_X1 U7110 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n3484), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6093), .ZN(n6106) );
  AOI21_X1 U7111 ( .B1(n6180), .B2(n6095), .A(n6094), .ZN(n6105) );
  INV_X1 U7112 ( .A(n6134), .ZN(n6100) );
  NOR2_X1 U7113 ( .A1(n6096), .A2(n6146), .ZN(n6098) );
  INV_X1 U7114 ( .A(n6132), .ZN(n6097) );
  AOI211_X1 U7115 ( .C1(n6100), .C2(n6099), .A(n6098), .B(n6097), .ZN(n6131)
         );
  OAI21_X1 U7116 ( .B1(n6102), .B2(n6101), .A(n6131), .ZN(n6110) );
  AOI22_X1 U7117 ( .A1(n6103), .A2(n6183), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6110), .ZN(n6104) );
  OAI211_X1 U7118 ( .C1(n6114), .C2(n6106), .A(n6105), .B(n6104), .ZN(U3008)
         );
  INV_X1 U7119 ( .A(n6107), .ZN(n6108) );
  AOI21_X1 U7120 ( .B1(n6180), .B2(n6109), .A(n6108), .ZN(n6113) );
  AOI22_X1 U7121 ( .A1(n6111), .A2(n6183), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6110), .ZN(n6112) );
  OAI211_X1 U7122 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6114), .A(n6113), 
        .B(n6112), .ZN(U3009) );
  OAI222_X1 U7123 ( .A1(n6116), .A2(n6160), .B1(n6159), .B2(n6475), .C1(n6157), 
        .C2(n6115), .ZN(n6117) );
  INV_X1 U7124 ( .A(n6117), .ZN(n6120) );
  OAI211_X1 U7125 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6126), .B(n6118), .ZN(n6119) );
  OAI211_X1 U7126 ( .C1(n6131), .C2(n6121), .A(n6120), .B(n6119), .ZN(U3010)
         );
  INV_X1 U7127 ( .A(n6122), .ZN(n6123) );
  AOI21_X1 U7128 ( .B1(n6180), .B2(n6124), .A(n6123), .ZN(n6129) );
  INV_X1 U7129 ( .A(n6125), .ZN(n6127) );
  AOI22_X1 U7130 ( .A1(n6127), .A2(n6183), .B1(n6126), .B2(n6130), .ZN(n6128)
         );
  OAI211_X1 U7131 ( .C1(n6131), .C2(n6130), .A(n6129), .B(n6128), .ZN(U3011)
         );
  OR2_X1 U7132 ( .A1(n6144), .A2(n6145), .ZN(n6135) );
  OAI21_X1 U7133 ( .B1(n6134), .B2(n6133), .A(n6132), .ZN(n6182) );
  AOI21_X1 U7134 ( .B1(n6136), .B2(n6135), .A(n6182), .ZN(n6155) );
  OAI22_X1 U7135 ( .A1(n6160), .A2(n6138), .B1(n6137), .B2(n6159), .ZN(n6140)
         );
  NOR4_X1 U7136 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6144), .A3(n6145), 
        .A4(n6163), .ZN(n6139) );
  AOI211_X1 U7137 ( .C1(n6141), .C2(n6183), .A(n6140), .B(n6139), .ZN(n6142)
         );
  OAI21_X1 U7138 ( .B1(n6155), .B2(n6143), .A(n6142), .ZN(U3012) );
  OAI21_X1 U7139 ( .B1(n6146), .B2(n6145), .A(n6144), .ZN(n6147) );
  AOI21_X1 U7140 ( .B1(n6148), .B2(n6186), .A(n6147), .ZN(n6154) );
  INV_X1 U7141 ( .A(n6149), .ZN(n6151) );
  AOI22_X1 U7142 ( .A1(n6151), .A2(n6183), .B1(n6180), .B2(n6150), .ZN(n6153)
         );
  NAND2_X1 U7143 ( .A1(n6185), .A2(REIP_REG_5__SCAN_IN), .ZN(n6152) );
  OAI211_X1 U7144 ( .C1(n6155), .C2(n6154), .A(n6153), .B(n6152), .ZN(U3013)
         );
  INV_X1 U7145 ( .A(n6176), .ZN(n6164) );
  AOI21_X1 U7146 ( .B1(n6179), .B2(n6164), .A(n6182), .ZN(n6175) );
  OAI222_X1 U7147 ( .A1(n6161), .A2(n6160), .B1(n6159), .B2(n6158), .C1(n6157), 
        .C2(n6156), .ZN(n6162) );
  INV_X1 U7148 ( .A(n6162), .ZN(n6167) );
  NOR2_X1 U7149 ( .A1(n6164), .A2(n6163), .ZN(n6171) );
  OAI211_X1 U7150 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6171), .B(n6165), .ZN(n6166) );
  OAI211_X1 U7151 ( .C1(n6175), .C2(n6168), .A(n6167), .B(n6166), .ZN(U3014)
         );
  AOI22_X1 U7152 ( .A1(n6180), .A2(n6169), .B1(n6185), .B2(REIP_REG_3__SCAN_IN), .ZN(n6173) );
  AOI22_X1 U7153 ( .A1(n6171), .A2(n6174), .B1(n6170), .B2(n6183), .ZN(n6172)
         );
  OAI211_X1 U7154 ( .C1(n6175), .C2(n6174), .A(n6173), .B(n6172), .ZN(U3015)
         );
  OAI21_X1 U7155 ( .B1(n6177), .B2(n3404), .A(n6176), .ZN(n6178) );
  AOI22_X1 U7156 ( .A1(n6181), .A2(n6180), .B1(n6179), .B2(n6178), .ZN(n6190)
         );
  AOI22_X1 U7157 ( .A1(n6184), .A2(n6183), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6182), .ZN(n6189) );
  NAND2_X1 U7158 ( .A1(n6185), .A2(REIP_REG_2__SCAN_IN), .ZN(n6188) );
  NAND3_X1 U7159 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6186), .A3(n3404), 
        .ZN(n6187) );
  NAND4_X1 U7160 ( .A1(n6190), .A2(n6189), .A3(n6188), .A4(n6187), .ZN(U3016)
         );
  INV_X1 U7161 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6192) );
  NOR2_X1 U7162 ( .A1(n6192), .A2(n6191), .ZN(U3019) );
  NOR2_X1 U7163 ( .A1(n6324), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6219)
         );
  AOI22_X1 U7164 ( .A1(n6326), .A2(n6219), .B1(n6273), .B2(n6218), .ZN(n6204)
         );
  NAND2_X1 U7165 ( .A1(n6194), .A2(n6193), .ZN(n6195) );
  OAI21_X1 U7166 ( .B1(n6196), .B2(n6195), .A(n6327), .ZN(n6202) );
  AOI21_X1 U7167 ( .B1(n6197), .B2(n6330), .A(n6219), .ZN(n6201) );
  INV_X1 U7168 ( .A(n6201), .ZN(n6199) );
  AOI21_X1 U7169 ( .B1(n6332), .B2(n6200), .A(n4760), .ZN(n6198) );
  OAI21_X1 U7170 ( .B1(n6202), .B2(n6199), .A(n6198), .ZN(n6221) );
  OAI22_X1 U7171 ( .A1(n6202), .A2(n6201), .B1(n6200), .B2(n6534), .ZN(n6220)
         );
  AOI22_X1 U7172 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6221), .B1(n6338), 
        .B2(n6220), .ZN(n6203) );
  OAI211_X1 U7173 ( .C1(n6285), .C2(n6224), .A(n6204), .B(n6203), .ZN(U3044)
         );
  AOI22_X1 U7174 ( .A1(n6343), .A2(n6219), .B1(n6342), .B2(n6207), .ZN(n6206)
         );
  AOI22_X1 U7175 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6221), .B1(n6344), 
        .B2(n6220), .ZN(n6205) );
  OAI211_X1 U7176 ( .C1(n6347), .C2(n6232), .A(n6206), .B(n6205), .ZN(U3045)
         );
  AOI22_X1 U7177 ( .A1(n6349), .A2(n6219), .B1(n6348), .B2(n6207), .ZN(n6209)
         );
  AOI22_X1 U7178 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6221), .B1(n6350), 
        .B2(n6220), .ZN(n6208) );
  OAI211_X1 U7179 ( .C1(n6353), .C2(n6232), .A(n6209), .B(n6208), .ZN(U3046)
         );
  AOI22_X1 U7180 ( .A1(n6388), .A2(n6219), .B1(n6392), .B2(n6218), .ZN(n6211)
         );
  AOI22_X1 U7181 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6221), .B1(n6390), 
        .B2(n6220), .ZN(n6210) );
  OAI211_X1 U7182 ( .C1(n6224), .C2(n6397), .A(n6211), .B(n6210), .ZN(U3047)
         );
  AOI22_X1 U7183 ( .A1(n6357), .A2(n6219), .B1(n6356), .B2(n6218), .ZN(n6213)
         );
  AOI22_X1 U7184 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6221), .B1(n6358), 
        .B2(n6220), .ZN(n6212) );
  OAI211_X1 U7185 ( .C1(n6224), .C2(n6361), .A(n6213), .B(n6212), .ZN(U3048)
         );
  AOI22_X1 U7186 ( .A1(n6363), .A2(n6219), .B1(n6318), .B2(n6218), .ZN(n6215)
         );
  AOI22_X1 U7187 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6221), .B1(n6364), 
        .B2(n6220), .ZN(n6214) );
  OAI211_X1 U7188 ( .C1(n6224), .C2(n6323), .A(n6215), .B(n6214), .ZN(U3049)
         );
  AOI22_X1 U7189 ( .A1(n6370), .A2(n6219), .B1(n6301), .B2(n6218), .ZN(n6217)
         );
  AOI22_X1 U7190 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6221), .B1(n6371), 
        .B2(n6220), .ZN(n6216) );
  OAI211_X1 U7191 ( .C1(n6224), .C2(n6304), .A(n6217), .B(n6216), .ZN(U3050)
         );
  AOI22_X1 U7192 ( .A1(n6378), .A2(n6219), .B1(n6375), .B2(n6218), .ZN(n6223)
         );
  AOI22_X1 U7193 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6221), .B1(n6380), 
        .B2(n6220), .ZN(n6222) );
  OAI211_X1 U7194 ( .C1(n6224), .C2(n6385), .A(n6223), .B(n6222), .ZN(U3051)
         );
  INV_X1 U7195 ( .A(n6225), .ZN(n6227) );
  AOI22_X1 U7196 ( .A1(n6390), .A2(n6227), .B1(n6388), .B2(n6226), .ZN(n6231)
         );
  AOI22_X1 U7197 ( .A1(n6229), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6392), 
        .B2(n6228), .ZN(n6230) );
  OAI211_X1 U7198 ( .C1(n6397), .C2(n6232), .A(n6231), .B(n6230), .ZN(U3055)
         );
  INV_X1 U7199 ( .A(n6235), .ZN(n6236) );
  OAI22_X1 U7200 ( .A1(n6238), .A2(n4415), .B1(n6237), .B2(n6236), .ZN(n6265)
         );
  NOR2_X1 U7201 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6280), .ZN(n6264)
         );
  AOI22_X1 U7202 ( .A1(n6338), .A2(n6265), .B1(n6326), .B2(n6264), .ZN(n6247)
         );
  INV_X1 U7203 ( .A(n6311), .ZN(n6298) );
  OAI21_X1 U7204 ( .B1(n6298), .B2(n6266), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6241) );
  NAND2_X1 U7205 ( .A1(n6240), .A2(n6239), .ZN(n6275) );
  NAND3_X1 U7206 ( .A1(n6241), .A2(n6327), .A3(n6275), .ZN(n6244) );
  OAI21_X1 U7207 ( .B1(n6519), .B2(n6264), .A(n6409), .ZN(n6242) );
  INV_X1 U7208 ( .A(n6242), .ZN(n6243) );
  NAND3_X1 U7209 ( .A1(n6245), .A2(n6244), .A3(n6243), .ZN(n6268) );
  AOI22_X1 U7210 ( .A1(n6268), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6325), 
        .B2(n6266), .ZN(n6246) );
  OAI211_X1 U7211 ( .C1(n6341), .C2(n6311), .A(n6247), .B(n6246), .ZN(U3068)
         );
  AOI22_X1 U7212 ( .A1(n6344), .A2(n6265), .B1(n6343), .B2(n6264), .ZN(n6249)
         );
  AOI22_X1 U7213 ( .A1(n6268), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6342), 
        .B2(n6266), .ZN(n6248) );
  OAI211_X1 U7214 ( .C1(n6347), .C2(n6311), .A(n6249), .B(n6248), .ZN(U3069)
         );
  AOI22_X1 U7215 ( .A1(n6350), .A2(n6265), .B1(n6349), .B2(n6264), .ZN(n6251)
         );
  AOI22_X1 U7216 ( .A1(n6268), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6348), 
        .B2(n6266), .ZN(n6250) );
  OAI211_X1 U7217 ( .C1(n6353), .C2(n6311), .A(n6251), .B(n6250), .ZN(U3070)
         );
  AOI22_X1 U7218 ( .A1(n6390), .A2(n6265), .B1(n6388), .B2(n6264), .ZN(n6254)
         );
  AOI22_X1 U7219 ( .A1(n6268), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6252), 
        .B2(n6266), .ZN(n6253) );
  OAI211_X1 U7220 ( .C1(n6255), .C2(n6311), .A(n6254), .B(n6253), .ZN(U3071)
         );
  AOI22_X1 U7221 ( .A1(n6358), .A2(n6265), .B1(n6357), .B2(n6264), .ZN(n6258)
         );
  AOI22_X1 U7222 ( .A1(n6268), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6256), 
        .B2(n6266), .ZN(n6257) );
  OAI211_X1 U7223 ( .C1(n6259), .C2(n6311), .A(n6258), .B(n6257), .ZN(U3072)
         );
  AOI22_X1 U7224 ( .A1(n6364), .A2(n6265), .B1(n6363), .B2(n6264), .ZN(n6261)
         );
  AOI22_X1 U7225 ( .A1(n6268), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6362), 
        .B2(n6266), .ZN(n6260) );
  OAI211_X1 U7226 ( .C1(n6367), .C2(n6311), .A(n6261), .B(n6260), .ZN(U3073)
         );
  AOI22_X1 U7227 ( .A1(n6371), .A2(n6265), .B1(n6370), .B2(n6264), .ZN(n6263)
         );
  AOI22_X1 U7228 ( .A1(n6268), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6368), 
        .B2(n6266), .ZN(n6262) );
  OAI211_X1 U7229 ( .C1(n6374), .C2(n6311), .A(n6263), .B(n6262), .ZN(U3074)
         );
  AOI22_X1 U7230 ( .A1(n6380), .A2(n6265), .B1(n6378), .B2(n6264), .ZN(n6270)
         );
  AOI22_X1 U7231 ( .A1(n6268), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6267), 
        .B2(n6266), .ZN(n6269) );
  OAI211_X1 U7232 ( .C1(n6271), .C2(n6311), .A(n6270), .B(n6269), .ZN(U3075)
         );
  INV_X1 U7233 ( .A(n6272), .ZN(n6306) );
  INV_X1 U7234 ( .A(n6322), .ZN(n6305) );
  AOI22_X1 U7235 ( .A1(n6326), .A2(n6306), .B1(n6273), .B2(n6305), .ZN(n6284)
         );
  NOR2_X1 U7236 ( .A1(n6274), .A2(n6332), .ZN(n6279) );
  INV_X1 U7237 ( .A(n6275), .ZN(n6276) );
  AOI21_X1 U7238 ( .B1(n6276), .B2(n6330), .A(n6306), .ZN(n6281) );
  AOI22_X1 U7239 ( .A1(n6279), .A2(n6281), .B1(n6280), .B2(n6332), .ZN(n6277)
         );
  NAND2_X1 U7240 ( .A1(n6278), .A2(n6277), .ZN(n6308) );
  INV_X1 U7241 ( .A(n6279), .ZN(n6282) );
  OAI22_X1 U7242 ( .A1(n6282), .A2(n6281), .B1(n6280), .B2(n6534), .ZN(n6307)
         );
  AOI22_X1 U7243 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6308), .B1(n6338), 
        .B2(n6307), .ZN(n6283) );
  OAI211_X1 U7244 ( .C1(n6285), .C2(n6311), .A(n6284), .B(n6283), .ZN(U3076)
         );
  AOI22_X1 U7245 ( .A1(n6343), .A2(n6306), .B1(n6286), .B2(n6305), .ZN(n6288)
         );
  AOI22_X1 U7246 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6308), .B1(n6344), 
        .B2(n6307), .ZN(n6287) );
  OAI211_X1 U7247 ( .C1(n6289), .C2(n6311), .A(n6288), .B(n6287), .ZN(U3077)
         );
  AOI22_X1 U7248 ( .A1(n6349), .A2(n6306), .B1(n6290), .B2(n6305), .ZN(n6292)
         );
  AOI22_X1 U7249 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6308), .B1(n6350), 
        .B2(n6307), .ZN(n6291) );
  OAI211_X1 U7250 ( .C1(n6293), .C2(n6311), .A(n6292), .B(n6291), .ZN(U3078)
         );
  AOI22_X1 U7251 ( .A1(n6388), .A2(n6306), .B1(n6392), .B2(n6305), .ZN(n6295)
         );
  AOI22_X1 U7252 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6308), .B1(n6390), 
        .B2(n6307), .ZN(n6294) );
  OAI211_X1 U7253 ( .C1(n6397), .C2(n6311), .A(n6295), .B(n6294), .ZN(U3079)
         );
  AOI22_X1 U7254 ( .A1(n6357), .A2(n6306), .B1(n6356), .B2(n6305), .ZN(n6297)
         );
  AOI22_X1 U7255 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6308), .B1(n6358), 
        .B2(n6307), .ZN(n6296) );
  OAI211_X1 U7256 ( .C1(n6361), .C2(n6311), .A(n6297), .B(n6296), .ZN(U3080)
         );
  AOI22_X1 U7257 ( .A1(n6363), .A2(n6306), .B1(n6362), .B2(n6298), .ZN(n6300)
         );
  AOI22_X1 U7258 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6308), .B1(n6364), 
        .B2(n6307), .ZN(n6299) );
  OAI211_X1 U7259 ( .C1(n6367), .C2(n6322), .A(n6300), .B(n6299), .ZN(U3081)
         );
  AOI22_X1 U7260 ( .A1(n6370), .A2(n6306), .B1(n6301), .B2(n6305), .ZN(n6303)
         );
  AOI22_X1 U7261 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6308), .B1(n6371), 
        .B2(n6307), .ZN(n6302) );
  OAI211_X1 U7262 ( .C1(n6304), .C2(n6311), .A(n6303), .B(n6302), .ZN(U3082)
         );
  AOI22_X1 U7263 ( .A1(n6378), .A2(n6306), .B1(n6375), .B2(n6305), .ZN(n6310)
         );
  AOI22_X1 U7264 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6308), .B1(n6380), 
        .B2(n6307), .ZN(n6309) );
  OAI211_X1 U7265 ( .C1(n6385), .C2(n6311), .A(n6310), .B(n6309), .ZN(U3083)
         );
  INV_X1 U7266 ( .A(n6312), .ZN(n6316) );
  AOI22_X1 U7267 ( .A1(n6390), .A2(n6316), .B1(n6388), .B2(n6315), .ZN(n6314)
         );
  AOI22_X1 U7268 ( .A1(n6319), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6392), 
        .B2(n6317), .ZN(n6313) );
  OAI211_X1 U7269 ( .C1(n6397), .C2(n6322), .A(n6314), .B(n6313), .ZN(U3087)
         );
  AOI22_X1 U7270 ( .A1(n6364), .A2(n6316), .B1(n6363), .B2(n6315), .ZN(n6321)
         );
  AOI22_X1 U7271 ( .A1(n6319), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6318), 
        .B2(n6317), .ZN(n6320) );
  OAI211_X1 U7272 ( .C1(n6323), .C2(n6322), .A(n6321), .B(n6320), .ZN(U3089)
         );
  NOR2_X1 U7273 ( .A1(n6324), .A2(n6409), .ZN(n6377) );
  AOI22_X1 U7274 ( .A1(n6326), .A2(n6377), .B1(n6369), .B2(n6325), .ZN(n6340)
         );
  OAI21_X1 U7275 ( .B1(n6329), .B2(n6328), .A(n6327), .ZN(n6337) );
  AOI21_X1 U7276 ( .B1(n6331), .B2(n6330), .A(n6377), .ZN(n6336) );
  INV_X1 U7277 ( .A(n6336), .ZN(n6334) );
  AOI21_X1 U7278 ( .B1(n6332), .B2(n6335), .A(n4760), .ZN(n6333) );
  OAI21_X1 U7279 ( .B1(n6337), .B2(n6334), .A(n6333), .ZN(n6381) );
  OAI22_X1 U7280 ( .A1(n6337), .A2(n6336), .B1(n6335), .B2(n6534), .ZN(n6379)
         );
  AOI22_X1 U7281 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6381), .B1(n6338), 
        .B2(n6379), .ZN(n6339) );
  OAI211_X1 U7282 ( .C1(n6341), .C2(n6396), .A(n6340), .B(n6339), .ZN(U3108)
         );
  AOI22_X1 U7283 ( .A1(n6343), .A2(n6377), .B1(n6369), .B2(n6342), .ZN(n6346)
         );
  AOI22_X1 U7284 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6381), .B1(n6344), 
        .B2(n6379), .ZN(n6345) );
  OAI211_X1 U7285 ( .C1(n6347), .C2(n6396), .A(n6346), .B(n6345), .ZN(U3109)
         );
  AOI22_X1 U7286 ( .A1(n6349), .A2(n6377), .B1(n6369), .B2(n6348), .ZN(n6352)
         );
  AOI22_X1 U7287 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6381), .B1(n6350), 
        .B2(n6379), .ZN(n6351) );
  OAI211_X1 U7288 ( .C1(n6353), .C2(n6396), .A(n6352), .B(n6351), .ZN(U3110)
         );
  AOI22_X1 U7289 ( .A1(n6388), .A2(n6377), .B1(n6376), .B2(n6392), .ZN(n6355)
         );
  AOI22_X1 U7290 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6381), .B1(n6390), 
        .B2(n6379), .ZN(n6354) );
  OAI211_X1 U7291 ( .C1(n6397), .C2(n6384), .A(n6355), .B(n6354), .ZN(U3111)
         );
  AOI22_X1 U7292 ( .A1(n6357), .A2(n6377), .B1(n6376), .B2(n6356), .ZN(n6360)
         );
  AOI22_X1 U7293 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6381), .B1(n6358), 
        .B2(n6379), .ZN(n6359) );
  OAI211_X1 U7294 ( .C1(n6361), .C2(n6384), .A(n6360), .B(n6359), .ZN(U3112)
         );
  AOI22_X1 U7295 ( .A1(n6363), .A2(n6377), .B1(n6369), .B2(n6362), .ZN(n6366)
         );
  AOI22_X1 U7296 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6381), .B1(n6364), 
        .B2(n6379), .ZN(n6365) );
  OAI211_X1 U7297 ( .C1(n6367), .C2(n6396), .A(n6366), .B(n6365), .ZN(U3113)
         );
  AOI22_X1 U7298 ( .A1(n6370), .A2(n6377), .B1(n6369), .B2(n6368), .ZN(n6373)
         );
  AOI22_X1 U7299 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6381), .B1(n6371), 
        .B2(n6379), .ZN(n6372) );
  OAI211_X1 U7300 ( .C1(n6374), .C2(n6396), .A(n6373), .B(n6372), .ZN(U3114)
         );
  AOI22_X1 U7301 ( .A1(n6378), .A2(n6377), .B1(n6376), .B2(n6375), .ZN(n6383)
         );
  AOI22_X1 U7302 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6381), .B1(n6380), 
        .B2(n6379), .ZN(n6382) );
  OAI211_X1 U7303 ( .C1(n6385), .C2(n6384), .A(n6383), .B(n6382), .ZN(U3115)
         );
  INV_X1 U7304 ( .A(n6386), .ZN(n6389) );
  AOI22_X1 U7305 ( .A1(n6390), .A2(n6389), .B1(n6388), .B2(n6387), .ZN(n6395)
         );
  AOI22_X1 U7306 ( .A1(n6393), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n6392), 
        .B2(n6391), .ZN(n6394) );
  OAI211_X1 U7307 ( .C1(n6397), .C2(n6396), .A(n6395), .B(n6394), .ZN(U3119)
         );
  INV_X1 U7308 ( .A(n6410), .ZN(n6414) );
  AOI21_X1 U7309 ( .B1(n6399), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n6398), 
        .ZN(n6400) );
  NAND2_X1 U7310 ( .A1(n6401), .A2(n6400), .ZN(n6402) );
  NOR2_X1 U7311 ( .A1(n6402), .A2(n6403), .ZN(n6407) );
  AOI22_X1 U7312 ( .A1(n6405), .A2(n6404), .B1(n6403), .B2(n6402), .ZN(n6406)
         );
  AOI211_X1 U7313 ( .C1(n6408), .C2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(n6407), .B(n6406), .ZN(n6412) );
  NOR2_X1 U7314 ( .A1(n6408), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6411)
         );
  OAI22_X1 U7315 ( .A1(n6412), .A2(n6411), .B1(n6410), .B2(n6409), .ZN(n6413)
         );
  OAI21_X1 U7316 ( .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6414), .A(n6413), 
        .ZN(n6423) );
  INV_X1 U7317 ( .A(MORE_REG_SCAN_IN), .ZN(n6656) );
  AOI21_X1 U7318 ( .B1(n6551), .B2(n6656), .A(n6415), .ZN(n6418) );
  NOR3_X1 U7319 ( .A1(n6418), .A2(n6417), .A3(n6416), .ZN(n6419) );
  NAND3_X1 U7320 ( .A1(n6421), .A2(n6420), .A3(n6419), .ZN(n6422) );
  AOI21_X1 U7321 ( .B1(n6423), .B2(n6192), .A(n6422), .ZN(n6436) );
  INV_X1 U7322 ( .A(n6424), .ZN(n6428) );
  AOI22_X1 U7323 ( .A1(n6436), .A2(n6426), .B1(READY_N), .B2(n6425), .ZN(n6427) );
  AOI21_X1 U7324 ( .B1(n6429), .B2(n6428), .A(n6427), .ZN(n6430) );
  INV_X1 U7325 ( .A(n6430), .ZN(n6518) );
  OAI21_X1 U7326 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6638), .A(n6518), .ZN(
        n6437) );
  AOI221_X1 U7327 ( .B1(n6432), .B2(STATE2_REG_0__SCAN_IN), .C1(n6437), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6431), .ZN(n6435) );
  OAI211_X1 U7328 ( .C1(n6535), .C2(n6433), .A(n6536), .B(n6518), .ZN(n6434)
         );
  OAI211_X1 U7329 ( .C1(n6436), .C2(n6438), .A(n6435), .B(n6434), .ZN(U3148)
         );
  NAND3_X1 U7330 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6444), .A3(n6437), .ZN(
        n6443) );
  OAI21_X1 U7331 ( .B1(READY_N), .B2(n6439), .A(n6438), .ZN(n6441) );
  AOI21_X1 U7332 ( .B1(n6441), .B2(n6518), .A(n6440), .ZN(n6442) );
  NAND2_X1 U7333 ( .A1(n6443), .A2(n6442), .ZN(U3149) );
  OAI211_X1 U7334 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6638), .A(n6516), .B(
        n6444), .ZN(n6446) );
  OAI21_X1 U7335 ( .B1(n6447), .B2(n6446), .A(n6445), .ZN(U3150) );
  AND2_X1 U7336 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6448), .ZN(U3151) );
  AND2_X1 U7337 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6448), .ZN(U3152) );
  AND2_X1 U7338 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6448), .ZN(U3153) );
  AND2_X1 U7339 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6448), .ZN(U3154) );
  AND2_X1 U7340 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6448), .ZN(U3155) );
  AND2_X1 U7341 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6448), .ZN(U3156) );
  AND2_X1 U7342 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6448), .ZN(U3157) );
  AND2_X1 U7343 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6448), .ZN(U3158) );
  AND2_X1 U7344 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6448), .ZN(U3159) );
  AND2_X1 U7345 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6448), .ZN(U3160) );
  AND2_X1 U7346 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6448), .ZN(U3161) );
  AND2_X1 U7347 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6448), .ZN(U3162) );
  AND2_X1 U7348 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6448), .ZN(U3163) );
  AND2_X1 U7349 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6448), .ZN(U3164) );
  AND2_X1 U7350 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6448), .ZN(U3165) );
  AND2_X1 U7351 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6448), .ZN(U3166) );
  AND2_X1 U7352 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6448), .ZN(U3167) );
  AND2_X1 U7353 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6448), .ZN(U3168) );
  AND2_X1 U7354 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6448), .ZN(U3169) );
  AND2_X1 U7355 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6448), .ZN(U3170) );
  AND2_X1 U7356 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6448), .ZN(U3171) );
  AND2_X1 U7357 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6448), .ZN(U3172) );
  AND2_X1 U7358 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6448), .ZN(U3173) );
  AND2_X1 U7359 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6448), .ZN(U3174) );
  AND2_X1 U7360 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6448), .ZN(U3175) );
  AND2_X1 U7361 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6448), .ZN(U3176) );
  AND2_X1 U7362 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6448), .ZN(U3177) );
  AND2_X1 U7363 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6448), .ZN(U3178) );
  AND2_X1 U7364 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6448), .ZN(U3179) );
  AND2_X1 U7365 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6448), .ZN(U3180) );
  NAND2_X1 U7366 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6451) );
  AND2_X1 U7367 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6450) );
  NOR2_X1 U7368 ( .A1(n6638), .A2(n6461), .ZN(n6454) );
  INV_X1 U7369 ( .A(NA_N), .ZN(n6671) );
  AOI221_X1 U7370 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6671), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6462) );
  AOI221_X1 U7371 ( .B1(n6450), .B2(n6457), .C1(n6454), .C2(n6457), .A(n6462), 
        .ZN(n6449) );
  OAI221_X1 U7372 ( .B1(n6739), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n6739), 
        .C2(n6451), .A(n6449), .ZN(U3181) );
  NAND2_X1 U7373 ( .A1(STATE_REG_0__SCAN_IN), .A2(REQUESTPENDING_REG_SCAN_IN), 
        .ZN(n6452) );
  AOI21_X1 U7374 ( .B1(n6452), .B2(n6451), .A(n6450), .ZN(n6453) );
  OR3_X1 U7375 ( .A1(n6455), .A2(n6454), .A3(n6453), .ZN(U3182) );
  NAND2_X1 U7376 ( .A1(READY_N), .A2(n6671), .ZN(n6456) );
  AOI21_X1 U7377 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6456), .A(
        REQUESTPENDING_REG_SCAN_IN), .ZN(n6459) );
  OAI21_X1 U7378 ( .B1(n6638), .B2(n6457), .A(STATE_REG_0__SCAN_IN), .ZN(n6458) );
  AOI221_X1 U7379 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6459), .C2(HOLD), .A(n6458), .ZN(n6463) );
  NAND4_X1 U7380 ( .A1(STATE_REG_0__SCAN_IN), .A2(READY_N), .A3(
        REQUESTPENDING_REG_SCAN_IN), .A4(n6671), .ZN(n6460) );
  OAI22_X1 U7381 ( .A1(n6463), .A2(n6462), .B1(n6461), .B2(n6460), .ZN(U3183)
         );
  NAND2_X1 U7382 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6739), .ZN(n6508) );
  NOR2_X2 U7383 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6500), .ZN(n6506) );
  AOI22_X1 U7384 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6500), .ZN(n6464) );
  OAI21_X1 U7385 ( .B1(n6527), .B2(n6508), .A(n6464), .ZN(U3184) );
  INV_X1 U7386 ( .A(n6506), .ZN(n6511) );
  INV_X1 U7387 ( .A(n6508), .ZN(n6509) );
  AOI22_X1 U7388 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6509), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6500), .ZN(n6465) );
  OAI21_X1 U7389 ( .B1(n6467), .B2(n6511), .A(n6465), .ZN(U3185) );
  AOI22_X1 U7390 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6500), .ZN(n6466) );
  OAI21_X1 U7391 ( .B1(n6467), .B2(n6508), .A(n6466), .ZN(U3186) );
  AOI22_X1 U7392 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6509), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6500), .ZN(n6468) );
  OAI21_X1 U7393 ( .B1(n6470), .B2(n6511), .A(n6468), .ZN(U3187) );
  AOI22_X1 U7394 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6500), .ZN(n6469) );
  OAI21_X1 U7395 ( .B1(n6470), .B2(n6508), .A(n6469), .ZN(U3188) );
  AOI22_X1 U7396 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6509), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6500), .ZN(n6471) );
  OAI21_X1 U7397 ( .B1(n6473), .B2(n6511), .A(n6471), .ZN(U3189) );
  AOI22_X1 U7398 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6500), .ZN(n6472) );
  OAI21_X1 U7399 ( .B1(n6473), .B2(n6508), .A(n6472), .ZN(U3190) );
  AOI22_X1 U7400 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6500), .ZN(n6474) );
  OAI21_X1 U7401 ( .B1(n6475), .B2(n6508), .A(n6474), .ZN(U3191) );
  INV_X1 U7402 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6477) );
  AOI22_X1 U7403 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6500), .ZN(n6476) );
  OAI21_X1 U7404 ( .B1(n6477), .B2(n6508), .A(n6476), .ZN(U3192) );
  AOI22_X1 U7405 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6509), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6500), .ZN(n6478) );
  OAI21_X1 U7406 ( .B1(n6480), .B2(n6511), .A(n6478), .ZN(U3193) );
  AOI22_X1 U7407 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6500), .ZN(n6479) );
  OAI21_X1 U7408 ( .B1(n6480), .B2(n6508), .A(n6479), .ZN(U3194) );
  AOI22_X1 U7409 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6509), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6500), .ZN(n6481) );
  OAI21_X1 U7410 ( .B1(n6482), .B2(n6511), .A(n6481), .ZN(U3195) );
  AOI22_X1 U7411 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6509), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6500), .ZN(n6483) );
  OAI21_X1 U7412 ( .B1(n6485), .B2(n6511), .A(n6483), .ZN(U3196) );
  AOI22_X1 U7413 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6500), .ZN(n6484) );
  OAI21_X1 U7414 ( .B1(n6485), .B2(n6508), .A(n6484), .ZN(U3197) );
  AOI22_X1 U7415 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6509), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6500), .ZN(n6486) );
  OAI21_X1 U7416 ( .B1(n6488), .B2(n6511), .A(n6486), .ZN(U3198) );
  AOI22_X1 U7417 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6500), .ZN(n6487) );
  OAI21_X1 U7418 ( .B1(n6488), .B2(n6508), .A(n6487), .ZN(U3199) );
  AOI22_X1 U7419 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6500), .ZN(n6489) );
  OAI21_X1 U7420 ( .B1(n6490), .B2(n6508), .A(n6489), .ZN(U3200) );
  AOI22_X1 U7421 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6509), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6500), .ZN(n6491) );
  OAI21_X1 U7422 ( .B1(n5657), .B2(n6511), .A(n6491), .ZN(U3201) );
  AOI22_X1 U7423 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6509), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6500), .ZN(n6492) );
  OAI21_X1 U7424 ( .B1(n6493), .B2(n6511), .A(n6492), .ZN(U3202) );
  AOI22_X1 U7425 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6509), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6500), .ZN(n6494) );
  OAI21_X1 U7426 ( .B1(n6496), .B2(n6511), .A(n6494), .ZN(U3203) );
  AOI22_X1 U7427 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6500), .ZN(n6495) );
  OAI21_X1 U7428 ( .B1(n6496), .B2(n6508), .A(n6495), .ZN(U3204) );
  AOI22_X1 U7429 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6500), .ZN(n6497) );
  OAI21_X1 U7430 ( .B1(n6498), .B2(n6508), .A(n6497), .ZN(U3205) );
  AOI22_X1 U7431 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6500), .ZN(n6499) );
  OAI21_X1 U7432 ( .B1(n3706), .B2(n6508), .A(n6499), .ZN(U3206) );
  AOI22_X1 U7433 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6500), .ZN(n6501) );
  OAI21_X1 U7434 ( .B1(n6683), .B2(n6508), .A(n6501), .ZN(U3207) );
  AOI22_X1 U7435 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6509), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6500), .ZN(n6502) );
  OAI21_X1 U7436 ( .B1(n6612), .B2(n6511), .A(n6502), .ZN(U3208) );
  AOI22_X1 U7437 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6500), .ZN(n6503) );
  OAI21_X1 U7438 ( .B1(n6612), .B2(n6508), .A(n6503), .ZN(U3209) );
  AOI22_X1 U7439 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6500), .ZN(n6504) );
  OAI21_X1 U7440 ( .B1(n6667), .B2(n6508), .A(n6504), .ZN(U3210) );
  AOI22_X1 U7441 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6509), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6500), .ZN(n6505) );
  OAI21_X1 U7442 ( .B1(n6738), .B2(n6511), .A(n6505), .ZN(U3211) );
  AOI22_X1 U7443 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6500), .ZN(n6507) );
  OAI21_X1 U7444 ( .B1(n6738), .B2(n6508), .A(n6507), .ZN(U3212) );
  AOI22_X1 U7445 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6509), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6500), .ZN(n6510) );
  OAI21_X1 U7446 ( .B1(n6655), .B2(n6511), .A(n6510), .ZN(U3213) );
  MUX2_X1 U7447 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6500), .Z(U3446) );
  MUX2_X1 U7448 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6500), .Z(U3447) );
  MUX2_X1 U7449 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6500), .Z(U3448) );
  OAI21_X1 U7450 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6515), .A(n6513), .ZN(
        n6512) );
  INV_X1 U7451 ( .A(n6512), .ZN(U3451) );
  OAI21_X1 U7452 ( .B1(n6515), .B2(n6514), .A(n6513), .ZN(U3452) );
  OAI211_X1 U7453 ( .C1(n6519), .C2(n6518), .A(n6517), .B(n6516), .ZN(U3453)
         );
  AOI22_X1 U7454 ( .A1(n6523), .A2(n6522), .B1(n6521), .B2(n6520), .ZN(n6524)
         );
  INV_X1 U7455 ( .A(n6524), .ZN(n6526) );
  MUX2_X1 U7456 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6526), .S(n6525), 
        .Z(U3456) );
  AOI21_X1 U7457 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6528) );
  AOI22_X1 U7458 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6528), .B2(n6527), .ZN(n6530) );
  INV_X1 U7459 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6641) );
  AOI22_X1 U7460 ( .A1(n6532), .A2(n6530), .B1(n6641), .B2(n6529), .ZN(U3468)
         );
  INV_X1 U7461 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6600) );
  OAI21_X1 U7462 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6532), .ZN(n6531) );
  OAI21_X1 U7463 ( .B1(n6532), .B2(n6600), .A(n6531), .ZN(U3469) );
  INV_X1 U7464 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6644) );
  AOI22_X1 U7465 ( .A1(n6739), .A2(READREQUEST_REG_SCAN_IN), .B1(n6644), .B2(
        n6500), .ZN(U3470) );
  AOI211_X1 U7466 ( .C1(n3359), .C2(n6604), .A(n6534), .B(n6533), .ZN(n6537)
         );
  OAI21_X1 U7467 ( .B1(n6537), .B2(n6536), .A(n6535), .ZN(n6542) );
  AOI211_X1 U7468 ( .C1(n6540), .C2(n6638), .A(n6539), .B(n6538), .ZN(n6541)
         );
  MUX2_X1 U7469 ( .A(n6542), .B(REQUESTPENDING_REG_SCAN_IN), .S(n6541), .Z(
        U3472) );
  OAI22_X1 U7470 ( .A1(n6500), .A2(MEMORYFETCH_REG_SCAN_IN), .B1(
        M_IO_N_REG_SCAN_IN), .B2(n6739), .ZN(n6543) );
  INV_X1 U7471 ( .A(n6543), .ZN(U3473) );
  INV_X1 U7472 ( .A(keyinput_f53), .ZN(n6636) );
  INV_X1 U7473 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6545) );
  AOI22_X1 U7474 ( .A1(n6667), .A2(keyinput_f55), .B1(keyinput_f42), .B2(n6545), .ZN(n6544) );
  OAI221_X1 U7475 ( .B1(n6667), .B2(keyinput_f55), .C1(n6545), .C2(
        keyinput_f42), .A(n6544), .ZN(n6634) );
  AOI22_X1 U7476 ( .A1(n6547), .A2(keyinput_f17), .B1(n3706), .B2(keyinput_f59), .ZN(n6546) );
  OAI221_X1 U7477 ( .B1(n6547), .B2(keyinput_f17), .C1(n3706), .C2(
        keyinput_f59), .A(n6546), .ZN(n6633) );
  OAI22_X1 U7478 ( .A1(n6647), .A2(keyinput_f23), .B1(n6549), .B2(keyinput_f25), .ZN(n6548) );
  AOI221_X1 U7479 ( .B1(n6647), .B2(keyinput_f23), .C1(keyinput_f25), .C2(
        n6549), .A(n6548), .ZN(n6566) );
  INV_X1 U7480 ( .A(DATAI_31_), .ZN(n6689) );
  AOI22_X1 U7481 ( .A1(n6551), .A2(keyinput_f45), .B1(n6689), .B2(keyinput_f0), 
        .ZN(n6550) );
  OAI221_X1 U7482 ( .B1(n6551), .B2(keyinput_f45), .C1(n6689), .C2(keyinput_f0), .A(n6550), .ZN(n6561) );
  INV_X1 U7483 ( .A(DATAI_25_), .ZN(n6706) );
  AOI22_X1 U7484 ( .A1(n6706), .A2(keyinput_f6), .B1(n6658), .B2(keyinput_f57), 
        .ZN(n6552) );
  OAI221_X1 U7485 ( .B1(n6706), .B2(keyinput_f6), .C1(n6658), .C2(keyinput_f57), .A(n6552), .ZN(n6560) );
  INV_X1 U7486 ( .A(DATAI_18_), .ZN(n6555) );
  INV_X1 U7487 ( .A(DATAI_16_), .ZN(n6554) );
  AOI22_X1 U7488 ( .A1(n6555), .A2(keyinput_f13), .B1(keyinput_f15), .B2(n6554), .ZN(n6553) );
  OAI221_X1 U7489 ( .B1(n6555), .B2(keyinput_f13), .C1(n6554), .C2(
        keyinput_f15), .A(n6553), .ZN(n6559) );
  INV_X1 U7490 ( .A(DATAI_28_), .ZN(n6557) );
  AOI22_X1 U7491 ( .A1(n6638), .A2(keyinput_f35), .B1(keyinput_f3), .B2(n6557), 
        .ZN(n6556) );
  OAI221_X1 U7492 ( .B1(n6638), .B2(keyinput_f35), .C1(n6557), .C2(keyinput_f3), .A(n6556), .ZN(n6558) );
  NOR4_X1 U7493 ( .A1(n6561), .A2(n6560), .A3(n6559), .A4(n6558), .ZN(n6565)
         );
  XOR2_X1 U7494 ( .A(keyinput_f38), .B(n6562), .Z(n6564) );
  XOR2_X1 U7495 ( .A(keyinput_f48), .B(n6640), .Z(n6563) );
  NAND4_X1 U7496 ( .A1(n6566), .A2(n6565), .A3(n6564), .A4(n6563), .ZN(n6632)
         );
  OAI22_X1 U7497 ( .A1(DATAI_1_), .A2(keyinput_f30), .B1(keyinput_f44), .B2(
        MORE_REG_SCAN_IN), .ZN(n6567) );
  AOI221_X1 U7498 ( .B1(DATAI_1_), .B2(keyinput_f30), .C1(MORE_REG_SCAN_IN), 
        .C2(keyinput_f44), .A(n6567), .ZN(n6630) );
  OAI22_X1 U7499 ( .A1(DATAI_0_), .A2(keyinput_f31), .B1(NA_N), .B2(
        keyinput_f33), .ZN(n6568) );
  AOI221_X1 U7500 ( .B1(DATAI_0_), .B2(keyinput_f31), .C1(keyinput_f33), .C2(
        NA_N), .A(n6568), .ZN(n6629) );
  AOI22_X1 U7501 ( .A1(DATAI_20_), .A2(keyinput_f11), .B1(REIP_REG_20__SCAN_IN), .B2(keyinput_f62), .ZN(n6569) );
  OAI221_X1 U7502 ( .B1(DATAI_20_), .B2(keyinput_f11), .C1(
        REIP_REG_20__SCAN_IN), .C2(keyinput_f62), .A(n6569), .ZN(n6576) );
  AOI22_X1 U7503 ( .A1(DATAI_27_), .A2(keyinput_f4), .B1(DATAI_29_), .B2(
        keyinput_f2), .ZN(n6570) );
  OAI221_X1 U7504 ( .B1(DATAI_27_), .B2(keyinput_f4), .C1(DATAI_29_), .C2(
        keyinput_f2), .A(n6570), .ZN(n6575) );
  AOI22_X1 U7505 ( .A1(DATAI_17_), .A2(keyinput_f14), .B1(DATAI_7_), .B2(
        keyinput_f24), .ZN(n6571) );
  OAI221_X1 U7506 ( .B1(DATAI_17_), .B2(keyinput_f14), .C1(DATAI_7_), .C2(
        keyinput_f24), .A(n6571), .ZN(n6574) );
  AOI22_X1 U7507 ( .A1(keyinput_f40), .A2(M_IO_N_REG_SCAN_IN), .B1(DATAI_2_), 
        .B2(keyinput_f29), .ZN(n6572) );
  OAI221_X1 U7508 ( .B1(keyinput_f40), .B2(M_IO_N_REG_SCAN_IN), .C1(DATAI_2_), 
        .C2(keyinput_f29), .A(n6572), .ZN(n6573) );
  NOR4_X1 U7509 ( .A1(n6576), .A2(n6575), .A3(n6574), .A4(n6573), .ZN(n6579)
         );
  INV_X1 U7510 ( .A(HOLD), .ZN(n6668) );
  OAI22_X1 U7511 ( .A1(keyinput_f36), .A2(n6668), .B1(DATAI_15_), .B2(
        keyinput_f16), .ZN(n6577) );
  AOI221_X1 U7512 ( .B1(n6668), .B2(keyinput_f36), .C1(DATAI_15_), .C2(
        keyinput_f16), .A(n6577), .ZN(n6578) );
  OAI211_X1 U7513 ( .C1(REIP_REG_21__SCAN_IN), .C2(keyinput_f61), .A(n6579), 
        .B(n6578), .ZN(n6580) );
  AOI21_X1 U7514 ( .B1(REIP_REG_21__SCAN_IN), .B2(keyinput_f61), .A(n6580), 
        .ZN(n6628) );
  OAI22_X1 U7515 ( .A1(DATAI_9_), .A2(keyinput_f22), .B1(keyinput_f46), .B2(
        W_R_N_REG_SCAN_IN), .ZN(n6581) );
  AOI221_X1 U7516 ( .B1(DATAI_9_), .B2(keyinput_f22), .C1(W_R_N_REG_SCAN_IN), 
        .C2(keyinput_f46), .A(n6581), .ZN(n6588) );
  OAI22_X1 U7517 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(DATAI_24_), .B2(
        keyinput_f7), .ZN(n6582) );
  AOI221_X1 U7518 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(keyinput_f7), .C2(
        DATAI_24_), .A(n6582), .ZN(n6587) );
  OAI22_X1 U7519 ( .A1(DATAI_5_), .A2(keyinput_f26), .B1(DATAI_19_), .B2(
        keyinput_f12), .ZN(n6583) );
  AOI221_X1 U7520 ( .B1(DATAI_5_), .B2(keyinput_f26), .C1(keyinput_f12), .C2(
        DATAI_19_), .A(n6583), .ZN(n6586) );
  OAI22_X1 U7521 ( .A1(REIP_REG_24__SCAN_IN), .A2(keyinput_f58), .B1(
        keyinput_f60), .B2(REIP_REG_22__SCAN_IN), .ZN(n6584) );
  AOI221_X1 U7522 ( .B1(REIP_REG_24__SCAN_IN), .B2(keyinput_f58), .C1(
        REIP_REG_22__SCAN_IN), .C2(keyinput_f60), .A(n6584), .ZN(n6585) );
  NAND4_X1 U7523 ( .A1(n6588), .A2(n6587), .A3(n6586), .A4(n6585), .ZN(n6626)
         );
  OAI22_X1 U7524 ( .A1(DATAI_26_), .A2(keyinput_f5), .B1(
        READREQUEST_REG_SCAN_IN), .B2(keyinput_f37), .ZN(n6589) );
  AOI221_X1 U7525 ( .B1(DATAI_26_), .B2(keyinput_f5), .C1(keyinput_f37), .C2(
        READREQUEST_REG_SCAN_IN), .A(n6589), .ZN(n6596) );
  OAI22_X1 U7526 ( .A1(DATAI_10_), .A2(keyinput_f21), .B1(DATAI_23_), .B2(
        keyinput_f8), .ZN(n6590) );
  AOI221_X1 U7527 ( .B1(DATAI_10_), .B2(keyinput_f21), .C1(keyinput_f8), .C2(
        DATAI_23_), .A(n6590), .ZN(n6595) );
  OAI22_X1 U7528 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput_f51), .B1(
        keyinput_f39), .B2(CODEFETCH_REG_SCAN_IN), .ZN(n6591) );
  AOI221_X1 U7529 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_f51), .C1(
        CODEFETCH_REG_SCAN_IN), .C2(keyinput_f39), .A(n6591), .ZN(n6594) );
  OAI22_X1 U7530 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_f32), .B1(BS16_N), .B2(keyinput_f34), .ZN(n6592) );
  AOI221_X1 U7531 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_f32), .C1(
        keyinput_f34), .C2(BS16_N), .A(n6592), .ZN(n6593) );
  NAND4_X1 U7532 ( .A1(n6596), .A2(n6595), .A3(n6594), .A4(n6593), .ZN(n6625)
         );
  OAI22_X1 U7533 ( .A1(n6664), .A2(keyinput_f19), .B1(n6598), .B2(keyinput_f20), .ZN(n6597) );
  AOI221_X1 U7534 ( .B1(n6664), .B2(keyinput_f19), .C1(keyinput_f20), .C2(
        n6598), .A(n6597), .ZN(n6609) );
  OAI22_X1 U7535 ( .A1(n6601), .A2(keyinput_f18), .B1(n6600), .B2(keyinput_f47), .ZN(n6599) );
  AOI221_X1 U7536 ( .B1(n6601), .B2(keyinput_f18), .C1(keyinput_f47), .C2(
        n6600), .A(n6599), .ZN(n6608) );
  OAI22_X1 U7537 ( .A1(n6604), .A2(keyinput_f43), .B1(n6603), .B2(keyinput_f50), .ZN(n6602) );
  AOI221_X1 U7538 ( .B1(n6604), .B2(keyinput_f43), .C1(keyinput_f50), .C2(
        n6603), .A(n6602), .ZN(n6607) );
  OAI22_X1 U7539 ( .A1(n5657), .A2(keyinput_f63), .B1(n6688), .B2(keyinput_f28), .ZN(n6605) );
  AOI221_X1 U7540 ( .B1(n5657), .B2(keyinput_f63), .C1(keyinput_f28), .C2(
        n6688), .A(n6605), .ZN(n6606) );
  NAND4_X1 U7541 ( .A1(n6609), .A2(n6608), .A3(n6607), .A4(n6606), .ZN(n6624)
         );
  OAI22_X1 U7542 ( .A1(n6612), .A2(keyinput_f56), .B1(n6611), .B2(keyinput_f27), .ZN(n6610) );
  AOI221_X1 U7543 ( .B1(n6612), .B2(keyinput_f56), .C1(keyinput_f27), .C2(
        n6611), .A(n6610), .ZN(n6622) );
  OAI22_X1 U7544 ( .A1(n6614), .A2(keyinput_f54), .B1(keyinput_f9), .B2(
        DATAI_22_), .ZN(n6613) );
  AOI221_X1 U7545 ( .B1(n6614), .B2(keyinput_f54), .C1(DATAI_22_), .C2(
        keyinput_f9), .A(n6613), .ZN(n6621) );
  INV_X1 U7546 ( .A(DATAI_21_), .ZN(n6616) );
  OAI22_X1 U7547 ( .A1(n6682), .A2(keyinput_f52), .B1(n6616), .B2(keyinput_f10), .ZN(n6615) );
  AOI221_X1 U7548 ( .B1(n6682), .B2(keyinput_f52), .C1(keyinput_f10), .C2(
        n6616), .A(n6615), .ZN(n6620) );
  INV_X1 U7549 ( .A(keyinput_f49), .ZN(n6618) );
  OAI22_X1 U7550 ( .A1(n6665), .A2(keyinput_f41), .B1(n6618), .B2(
        BYTEENABLE_REG_2__SCAN_IN), .ZN(n6617) );
  AOI221_X1 U7551 ( .B1(n6665), .B2(keyinput_f41), .C1(
        BYTEENABLE_REG_2__SCAN_IN), .C2(n6618), .A(n6617), .ZN(n6619) );
  NAND4_X1 U7552 ( .A1(n6622), .A2(n6621), .A3(n6620), .A4(n6619), .ZN(n6623)
         );
  NOR4_X1 U7553 ( .A1(n6626), .A2(n6625), .A3(n6624), .A4(n6623), .ZN(n6627)
         );
  NAND4_X1 U7554 ( .A1(n6630), .A2(n6629), .A3(n6628), .A4(n6627), .ZN(n6631)
         );
  NOR4_X1 U7555 ( .A1(n6634), .A2(n6633), .A3(n6632), .A4(n6631), .ZN(n6635)
         );
  AOI221_X1 U7556 ( .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_f53), .C1(n6738), 
        .C2(n6636), .A(n6635), .ZN(n6737) );
  AOI22_X1 U7557 ( .A1(n6638), .A2(keyinput_g35), .B1(keyinput_g63), .B2(n5657), .ZN(n6637) );
  OAI221_X1 U7558 ( .B1(n6638), .B2(keyinput_g35), .C1(n5657), .C2(
        keyinput_g63), .A(n6637), .ZN(n6651) );
  AOI22_X1 U7559 ( .A1(n6641), .A2(keyinput_g49), .B1(keyinput_g48), .B2(n6640), .ZN(n6639) );
  OAI221_X1 U7560 ( .B1(n6641), .B2(keyinput_g49), .C1(n6640), .C2(
        keyinput_g48), .A(n6639), .ZN(n6650) );
  AOI22_X1 U7561 ( .A1(n6644), .A2(keyinput_g46), .B1(n6643), .B2(keyinput_g31), .ZN(n6642) );
  OAI221_X1 U7562 ( .B1(n6644), .B2(keyinput_g46), .C1(n6643), .C2(
        keyinput_g31), .A(n6642), .ZN(n6649) );
  INV_X1 U7563 ( .A(DATAI_19_), .ZN(n6646) );
  AOI22_X1 U7564 ( .A1(n6647), .A2(keyinput_g23), .B1(keyinput_g12), .B2(n6646), .ZN(n6645) );
  OAI221_X1 U7565 ( .B1(n6647), .B2(keyinput_g23), .C1(n6646), .C2(
        keyinput_g12), .A(n6645), .ZN(n6648) );
  NOR4_X1 U7566 ( .A1(n6651), .A2(n6650), .A3(n6649), .A4(n6648), .ZN(n6697)
         );
  AOI22_X1 U7567 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_g32), .B1(
        STATEBS16_REG_SCAN_IN), .B2(keyinput_g43), .ZN(n6652) );
  OAI221_X1 U7568 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_g32), .C1(
        STATEBS16_REG_SCAN_IN), .C2(keyinput_g43), .A(n6652), .ZN(n6662) );
  AOI22_X1 U7569 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_g50), .B1(
        DATAI_2_), .B2(keyinput_g29), .ZN(n6653) );
  OAI221_X1 U7570 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_g50), .C1(
        DATAI_2_), .C2(keyinput_g29), .A(n6653), .ZN(n6661) );
  AOI22_X1 U7571 ( .A1(n6656), .A2(keyinput_g44), .B1(n6655), .B2(keyinput_g51), .ZN(n6654) );
  OAI221_X1 U7572 ( .B1(n6656), .B2(keyinput_g44), .C1(n6655), .C2(
        keyinput_g51), .A(n6654), .ZN(n6660) );
  AOI22_X1 U7573 ( .A1(DATAI_26_), .A2(keyinput_g5), .B1(n6658), .B2(
        keyinput_g57), .ZN(n6657) );
  OAI221_X1 U7574 ( .B1(DATAI_26_), .B2(keyinput_g5), .C1(n6658), .C2(
        keyinput_g57), .A(n6657), .ZN(n6659) );
  NOR4_X1 U7575 ( .A1(n6662), .A2(n6661), .A3(n6660), .A4(n6659), .ZN(n6696)
         );
  AOI22_X1 U7576 ( .A1(n6665), .A2(keyinput_g41), .B1(n6664), .B2(keyinput_g19), .ZN(n6663) );
  OAI221_X1 U7577 ( .B1(n6665), .B2(keyinput_g41), .C1(n6664), .C2(
        keyinput_g19), .A(n6663), .ZN(n6678) );
  AOI22_X1 U7578 ( .A1(n6668), .A2(keyinput_g36), .B1(n6667), .B2(keyinput_g55), .ZN(n6666) );
  OAI221_X1 U7579 ( .B1(n6668), .B2(keyinput_g36), .C1(n6667), .C2(
        keyinput_g55), .A(n6666), .ZN(n6677) );
  AOI22_X1 U7580 ( .A1(n6671), .A2(keyinput_g33), .B1(n6670), .B2(keyinput_g37), .ZN(n6669) );
  OAI221_X1 U7581 ( .B1(n6671), .B2(keyinput_g33), .C1(n6670), .C2(
        keyinput_g37), .A(n6669), .ZN(n6676) );
  INV_X1 U7582 ( .A(DATAI_20_), .ZN(n6673) );
  AOI22_X1 U7583 ( .A1(n6674), .A2(keyinput_g26), .B1(keyinput_g11), .B2(n6673), .ZN(n6672) );
  OAI221_X1 U7584 ( .B1(n6674), .B2(keyinput_g26), .C1(n6673), .C2(
        keyinput_g11), .A(n6672), .ZN(n6675) );
  NOR4_X1 U7585 ( .A1(n6678), .A2(n6677), .A3(n6676), .A4(n6675), .ZN(n6695)
         );
  INV_X1 U7586 ( .A(DATAI_17_), .ZN(n6680) );
  AOI22_X1 U7587 ( .A1(n6680), .A2(keyinput_g14), .B1(keyinput_g16), .B2(n4396), .ZN(n6679) );
  OAI221_X1 U7588 ( .B1(n6680), .B2(keyinput_g14), .C1(n4396), .C2(
        keyinput_g16), .A(n6679), .ZN(n6693) );
  AOI22_X1 U7589 ( .A1(n6683), .A2(keyinput_g58), .B1(n6682), .B2(keyinput_g52), .ZN(n6681) );
  OAI221_X1 U7590 ( .B1(n6683), .B2(keyinput_g58), .C1(n6682), .C2(
        keyinput_g52), .A(n6681), .ZN(n6692) );
  INV_X1 U7591 ( .A(DATAI_24_), .ZN(n6686) );
  INV_X1 U7592 ( .A(DATAI_23_), .ZN(n6685) );
  AOI22_X1 U7593 ( .A1(n6686), .A2(keyinput_g7), .B1(keyinput_g8), .B2(n6685), 
        .ZN(n6684) );
  OAI221_X1 U7594 ( .B1(n6686), .B2(keyinput_g7), .C1(n6685), .C2(keyinput_g8), 
        .A(n6684), .ZN(n6691) );
  AOI22_X1 U7595 ( .A1(n6689), .A2(keyinput_g0), .B1(keyinput_g28), .B2(n6688), 
        .ZN(n6687) );
  OAI221_X1 U7596 ( .B1(n6689), .B2(keyinput_g0), .C1(n6688), .C2(keyinput_g28), .A(n6687), .ZN(n6690) );
  NOR4_X1 U7597 ( .A1(n6693), .A2(n6692), .A3(n6691), .A4(n6690), .ZN(n6694)
         );
  NAND4_X1 U7598 ( .A1(n6697), .A2(n6696), .A3(n6695), .A4(n6694), .ZN(n6735)
         );
  AOI22_X1 U7599 ( .A1(BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_g47), .B1(
        DATAI_21_), .B2(keyinput_g10), .ZN(n6698) );
  OAI221_X1 U7600 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_g47), .C1(
        DATAI_21_), .C2(keyinput_g10), .A(n6698), .ZN(n6705) );
  AOI22_X1 U7601 ( .A1(DATAI_10_), .A2(keyinput_g21), .B1(DATAI_29_), .B2(
        keyinput_g2), .ZN(n6699) );
  OAI221_X1 U7602 ( .B1(DATAI_10_), .B2(keyinput_g21), .C1(DATAI_29_), .C2(
        keyinput_g2), .A(n6699), .ZN(n6704) );
  AOI22_X1 U7603 ( .A1(DATAI_16_), .A2(keyinput_g15), .B1(REIP_REG_26__SCAN_IN), .B2(keyinput_g56), .ZN(n6700) );
  OAI221_X1 U7604 ( .B1(DATAI_16_), .B2(keyinput_g15), .C1(
        REIP_REG_26__SCAN_IN), .C2(keyinput_g56), .A(n6700), .ZN(n6703) );
  AOI22_X1 U7605 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(keyinput_g39), .B1(
        DATAI_18_), .B2(keyinput_g13), .ZN(n6701) );
  OAI221_X1 U7606 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_g39), .C1(
        DATAI_18_), .C2(keyinput_g13), .A(n6701), .ZN(n6702) );
  NOR4_X1 U7607 ( .A1(n6705), .A2(n6704), .A3(n6703), .A4(n6702), .ZN(n6733)
         );
  XNOR2_X1 U7608 ( .A(n6706), .B(keyinput_g6), .ZN(n6713) );
  AOI22_X1 U7609 ( .A1(DATAI_7_), .A2(keyinput_g24), .B1(DATAI_11_), .B2(
        keyinput_g20), .ZN(n6707) );
  OAI221_X1 U7610 ( .B1(DATAI_7_), .B2(keyinput_g24), .C1(DATAI_11_), .C2(
        keyinput_g20), .A(n6707), .ZN(n6712) );
  AOI22_X1 U7611 ( .A1(ADS_N_REG_SCAN_IN), .A2(keyinput_g38), .B1(
        M_IO_N_REG_SCAN_IN), .B2(keyinput_g40), .ZN(n6708) );
  OAI221_X1 U7612 ( .B1(ADS_N_REG_SCAN_IN), .B2(keyinput_g38), .C1(
        M_IO_N_REG_SCAN_IN), .C2(keyinput_g40), .A(n6708), .ZN(n6711) );
  AOI22_X1 U7613 ( .A1(DATAI_22_), .A2(keyinput_g9), .B1(REIP_REG_22__SCAN_IN), 
        .B2(keyinput_g60), .ZN(n6709) );
  OAI221_X1 U7614 ( .B1(DATAI_22_), .B2(keyinput_g9), .C1(REIP_REG_22__SCAN_IN), .C2(keyinput_g60), .A(n6709), .ZN(n6710) );
  NOR4_X1 U7615 ( .A1(n6713), .A2(n6712), .A3(n6711), .A4(n6710), .ZN(n6732)
         );
  AOI22_X1 U7616 ( .A1(DATAI_4_), .A2(keyinput_g27), .B1(DATAI_30_), .B2(
        keyinput_g1), .ZN(n6714) );
  OAI221_X1 U7617 ( .B1(DATAI_4_), .B2(keyinput_g27), .C1(DATAI_30_), .C2(
        keyinput_g1), .A(n6714), .ZN(n6721) );
  AOI22_X1 U7618 ( .A1(DATAI_28_), .A2(keyinput_g3), .B1(DATAI_14_), .B2(
        keyinput_g17), .ZN(n6715) );
  OAI221_X1 U7619 ( .B1(DATAI_28_), .B2(keyinput_g3), .C1(DATAI_14_), .C2(
        keyinput_g17), .A(n6715), .ZN(n6720) );
  AOI22_X1 U7620 ( .A1(FLUSH_REG_SCAN_IN), .A2(keyinput_g45), .B1(
        REIP_REG_20__SCAN_IN), .B2(keyinput_g62), .ZN(n6716) );
  OAI221_X1 U7621 ( .B1(FLUSH_REG_SCAN_IN), .B2(keyinput_g45), .C1(
        REIP_REG_20__SCAN_IN), .C2(keyinput_g62), .A(n6716), .ZN(n6719) );
  AOI22_X1 U7622 ( .A1(DATAI_9_), .A2(keyinput_g22), .B1(DATAI_13_), .B2(
        keyinput_g18), .ZN(n6717) );
  OAI221_X1 U7623 ( .B1(DATAI_9_), .B2(keyinput_g22), .C1(DATAI_13_), .C2(
        keyinput_g18), .A(n6717), .ZN(n6718) );
  NOR4_X1 U7624 ( .A1(n6721), .A2(n6720), .A3(n6719), .A4(n6718), .ZN(n6731)
         );
  AOI22_X1 U7625 ( .A1(REIP_REG_21__SCAN_IN), .A2(keyinput_g61), .B1(
        REIP_REG_23__SCAN_IN), .B2(keyinput_g59), .ZN(n6722) );
  OAI221_X1 U7626 ( .B1(REIP_REG_21__SCAN_IN), .B2(keyinput_g61), .C1(
        REIP_REG_23__SCAN_IN), .C2(keyinput_g59), .A(n6722), .ZN(n6729) );
  AOI22_X1 U7627 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_g42), .B1(
        DATAI_27_), .B2(keyinput_g4), .ZN(n6723) );
  OAI221_X1 U7628 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_g42), .C1(
        DATAI_27_), .C2(keyinput_g4), .A(n6723), .ZN(n6728) );
  AOI22_X1 U7629 ( .A1(DATAI_1_), .A2(keyinput_g30), .B1(DATAI_6_), .B2(
        keyinput_g25), .ZN(n6724) );
  OAI221_X1 U7630 ( .B1(DATAI_1_), .B2(keyinput_g30), .C1(DATAI_6_), .C2(
        keyinput_g25), .A(n6724), .ZN(n6727) );
  AOI22_X1 U7631 ( .A1(BS16_N), .A2(keyinput_g34), .B1(REIP_REG_28__SCAN_IN), 
        .B2(keyinput_g54), .ZN(n6725) );
  OAI221_X1 U7632 ( .B1(BS16_N), .B2(keyinput_g34), .C1(REIP_REG_28__SCAN_IN), 
        .C2(keyinput_g54), .A(n6725), .ZN(n6726) );
  NOR4_X1 U7633 ( .A1(n6729), .A2(n6728), .A3(n6727), .A4(n6726), .ZN(n6730)
         );
  NAND4_X1 U7634 ( .A1(n6733), .A2(n6732), .A3(n6731), .A4(n6730), .ZN(n6734)
         );
  OAI22_X1 U7635 ( .A1(keyinput_g53), .A2(n6738), .B1(n6735), .B2(n6734), .ZN(
        n6736) );
  AOI211_X1 U7636 ( .C1(keyinput_g53), .C2(n6738), .A(n6737), .B(n6736), .ZN(
        n6741) );
  AOI22_X1 U7637 ( .A1(n6739), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6500), .ZN(n6740) );
  XNOR2_X1 U7638 ( .A(n6741), .B(n6740), .ZN(U3445) );
  CLKBUF_X1 U34690 ( .A(n3138), .Z(n3239) );
  AND4_X1 U3767 ( .A1(n3060), .A2(n3059), .A3(n3058), .A4(n3057), .ZN(n3066)
         );
  CLKBUF_X1 U4045 ( .A(n3244), .Z(n5267) );
  CLKBUF_X1 U4047 ( .A(n3372), .Z(n3373) );
  CLKBUF_X1 U4176 ( .A(n3753), .Z(n6330) );
endmodule

