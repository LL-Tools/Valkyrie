

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960;

  INV_X2 U4765 ( .A(n8178), .ZN(n9844) );
  INV_X2 U4766 ( .A(n6912), .ZN(n6919) );
  XNOR2_X1 U4769 ( .A(n4964), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6396) );
  AND2_X1 U4770 ( .A1(n4856), .A2(n4862), .ZN(n4942) );
  NOR2_X1 U4771 ( .A1(n8471), .A2(n4615), .ZN(n4614) );
  INV_X1 U4772 ( .A(n5743), .ZN(n5899) );
  OR2_X1 U4773 ( .A1(n8438), .A2(n4296), .ZN(n8424) );
  INV_X1 U4774 ( .A(n6760), .ZN(n6734) );
  INV_X1 U4775 ( .A(n4960), .ZN(n5008) );
  OAI211_X1 U4776 ( .C1(n5008), .C2(n6766), .A(n4968), .B(n4967), .ZN(n7051)
         );
  NAND2_X1 U4777 ( .A1(n5208), .A2(n5066), .ZN(n5071) );
  INV_X1 U4778 ( .A(n9827), .ZN(n6763) );
  AND3_X1 U4780 ( .A1(n6438), .A2(n6440), .A3(n6439), .ZN(n4794) );
  XNOR2_X1 U4781 ( .A(n4354), .B(n8469), .ZN(n8473) );
  AND2_X1 U4782 ( .A1(n4745), .A2(n4748), .ZN(n6760) );
  INV_X1 U4783 ( .A(n7711), .ZN(n9850) );
  INV_X1 U4784 ( .A(n5026), .ZN(n5482) );
  INV_X1 U4785 ( .A(n5355), .ZN(n5340) );
  XNOR2_X1 U4786 ( .A(n7497), .B(n7496), .ZN(n7280) );
  INV_X1 U4787 ( .A(n7523), .ZN(n7380) );
  INV_X1 U4788 ( .A(n5683), .ZN(n9664) );
  INV_X1 U4789 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9535) );
  INV_X1 U4790 ( .A(n8461), .ZN(n8455) );
  NOR2_X1 U4791 ( .A1(n4426), .A2(n4425), .ZN(n4424) );
  INV_X4 U4792 ( .A(n6442), .ZN(n6445) );
  INV_X1 U4793 ( .A(n6456), .ZN(n8389) );
  INV_X2 U4794 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  AOI22_X2 U4795 ( .A1(n8555), .A2(n8554), .B1(n8761), .B2(n8581), .ZN(n8543)
         );
  INV_X2 U4796 ( .A(n6219), .ZN(n6224) );
  NOR2_X2 U4797 ( .A1(n7262), .A2(n8017), .ZN(n4560) );
  NAND2_X2 U4798 ( .A1(n4931), .A2(n4930), .ZN(n5683) );
  NAND2_X1 U4799 ( .A1(n4726), .A2(n4725), .ZN(n8965) );
  AND2_X1 U4800 ( .A1(n5846), .A2(n5845), .ZN(n8956) );
  NAND2_X1 U4801 ( .A1(n8414), .A2(n4349), .ZN(n8525) );
  AOI21_X1 U4802 ( .B1(n4606), .B2(n4294), .A(n4607), .ZN(n8439) );
  AOI21_X1 U4803 ( .B1(n4822), .B2(n4825), .A(n8469), .ZN(n4821) );
  INV_X1 U4804 ( .A(n8499), .ZN(n4606) );
  OAI21_X1 U4805 ( .B1(n4263), .B2(n8461), .A(n4608), .ZN(n4607) );
  NAND2_X1 U4806 ( .A1(n9071), .A2(n4830), .ZN(n9285) );
  AND2_X1 U4807 ( .A1(n8562), .A2(n8247), .ZN(n8548) );
  XNOR2_X1 U4808 ( .A(n5440), .B(n5439), .ZN(n8827) );
  NAND2_X1 U4809 ( .A1(n5416), .A2(n5415), .ZN(n5440) );
  AOI21_X1 U4810 ( .B1(n9063), .B2(n4291), .A(n4784), .ZN(n9320) );
  NAND2_X1 U4811 ( .A1(n8684), .A2(n4292), .ZN(n8673) );
  NAND2_X1 U4812 ( .A1(n8686), .A2(n8685), .ZN(n8684) );
  NAND2_X1 U4813 ( .A1(n5414), .A2(n5413), .ZN(n5416) );
  AND2_X1 U4814 ( .A1(n8402), .A2(n8401), .ZN(n8686) );
  NAND2_X1 U4815 ( .A1(n7508), .A2(n4827), .ZN(n9727) );
  NAND2_X1 U4816 ( .A1(n4350), .A2(n7337), .ZN(n7508) );
  NAND2_X1 U4817 ( .A1(n5272), .A2(n5271), .ZN(n9463) );
  NAND2_X1 U4818 ( .A1(n5256), .A2(n5255), .ZN(n9468) );
  AND2_X1 U4819 ( .A1(n8635), .A2(n8640), .ZN(n8636) );
  NOR2_X1 U4820 ( .A1(n7214), .A2(n7711), .ZN(n9751) );
  OR3_X1 U4821 ( .A1(n7116), .A2(n7115), .A3(n7114), .ZN(n8185) );
  INV_X2 U4822 ( .A(n9910), .ZN(n4260) );
  NAND2_X1 U4823 ( .A1(n8154), .A2(n8149), .ZN(n8121) );
  OAI211_X1 U4824 ( .C1(n6926), .C2(n5008), .A(n5007), .B(n5006), .ZN(n7523)
         );
  INV_X1 U4825 ( .A(n7051), .ZN(n5706) );
  XNOR2_X1 U4826 ( .A(n4381), .B(n5004), .ZN(n6926) );
  INV_X8 U4827 ( .A(n4261), .ZN(n7689) );
  AND4_X1 U4828 ( .A1(n4988), .A2(n4987), .A3(n4986), .A4(n4985), .ZN(n7379)
         );
  NAND3_X2 U4829 ( .A1(n4953), .A2(n4952), .A3(n4951), .ZN(n8948) );
  AND4_X1 U4830 ( .A1(n4959), .A2(n4958), .A3(n4957), .A4(n4956), .ZN(n7032)
         );
  AND4_X1 U4831 ( .A1(n5003), .A2(n5002), .A3(n5001), .A4(n5000), .ZN(n7438)
         );
  OAI211_X1 U4832 ( .C1(n5008), .C2(n6816), .A(n4981), .B(n4980), .ZN(n7059)
         );
  BUF_X2 U4833 ( .A(n5707), .Z(n4261) );
  NOR2_X2 U4834 ( .A1(n7234), .A2(n7204), .ZN(n7261) );
  INV_X1 U4835 ( .A(n9834), .ZN(n7021) );
  INV_X1 U4836 ( .A(n8318), .ZN(n9702) );
  NAND2_X1 U4837 ( .A1(n4794), .A2(n6437), .ZN(n6724) );
  BUF_X2 U4838 ( .A(n7916), .Z(n7141) );
  OAI211_X1 U4839 ( .C1(n6768), .C2(n6728), .A(n6727), .B(n6726), .ZN(n9827)
         );
  INV_X4 U4840 ( .A(n9207), .ZN(n9250) );
  NAND2_X1 U4841 ( .A1(n5519), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5070) );
  AND2_X1 U4842 ( .A1(n4855), .A2(n9536), .ZN(n9543) );
  NAND2_X1 U4843 ( .A1(n5519), .A2(n5518), .ZN(n5670) );
  NAND2_X1 U4844 ( .A1(n4348), .A2(n5916), .ZN(n5954) );
  XNOR2_X1 U4845 ( .A(n4852), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9540) );
  NAND2_X1 U4846 ( .A1(n6768), .A2(n6442), .ZN(n6815) );
  NOR2_X1 U4847 ( .A1(n7352), .A2(n7472), .ZN(n4348) );
  XNOR2_X1 U4848 ( .A(n5660), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5916) );
  AOI21_X1 U4849 ( .B1(n5071), .B2(P1_IR_REG_31__SCAN_IN), .A(n4732), .ZN(
        n4731) );
  OR2_X1 U4850 ( .A1(n4854), .A2(n9535), .ZN(n4852) );
  NAND2_X1 U4851 ( .A1(n5664), .A2(n5663), .ZN(n7472) );
  AND2_X1 U4852 ( .A1(n4873), .A2(n4791), .ZN(n4854) );
  MUX2_X1 U4853 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6215), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n6217) );
  NAND2_X1 U4854 ( .A1(n5663), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U4855 ( .A1(n6079), .A2(n4427), .ZN(n8828) );
  NAND2_X1 U4856 ( .A1(n6079), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4428) );
  NAND2_X2 U4857 ( .A1(n6445), .A2(P1_U3084), .ZN(n9552) );
  NOR2_X1 U4858 ( .A1(n6445), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9549) );
  NOR2_X1 U4859 ( .A1(n4812), .A2(n4645), .ZN(n4644) );
  AND2_X1 U4860 ( .A1(n4729), .A2(n5064), .ZN(n4728) );
  NAND2_X1 U4861 ( .A1(n4733), .A2(n5068), .ZN(n4732) );
  AND2_X1 U4862 ( .A1(n4790), .A2(n4600), .ZN(n4599) );
  AND2_X1 U4863 ( .A1(n4730), .A2(n5063), .ZN(n4729) );
  INV_X1 U4864 ( .A(n4978), .ZN(n4841) );
  NOR2_X1 U4865 ( .A1(n4844), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n4730) );
  NAND2_X1 U4866 ( .A1(n4734), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4733) );
  NAND3_X1 U4867 ( .A1(n9040), .A2(n4650), .A3(n4649), .ZN(n4533) );
  INV_X4 U4868 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U4869 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4839) );
  INV_X1 U4870 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6072) );
  INV_X1 U4871 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6078) );
  NOR2_X1 U4872 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4845) );
  NOR2_X1 U4873 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n4600) );
  INV_X1 U4874 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5211) );
  INV_X1 U4875 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5978) );
  INV_X1 U4876 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4877) );
  INV_X1 U4877 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5067) );
  NOR2_X1 U4878 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5955) );
  NOR2_X1 U4879 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5956) );
  INV_X1 U4880 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5068) );
  INV_X1 U4881 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9040) );
  INV_X1 U4882 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4781) );
  INV_X1 U4883 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4840) );
  NOR2_X2 U4884 ( .A1(n8658), .A2(n8659), .ZN(n8657) );
  NAND2_X2 U4885 ( .A1(n4949), .A2(n6442), .ZN(n5050) );
  XNOR2_X1 U4886 ( .A(n5683), .B(n5682), .ZN(n5529) );
  NOR2_X2 U4887 ( .A1(n5173), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n5208) );
  INV_X1 U4888 ( .A(n5699), .ZN(n5707) );
  AND2_X1 U4889 ( .A1(n4700), .A2(n5954), .ZN(n4262) );
  OAI21_X2 U4890 ( .B1(n7243), .B2(n5738), .A(n5737), .ZN(n7375) );
  NAND2_X2 U4891 ( .A1(n7028), .A2(n5727), .ZN(n7243) );
  INV_X2 U4892 ( .A(n4949), .ZN(n5982) );
  CLKBUF_X3 U4893 ( .A(n6817), .Z(n8111) );
  AOI21_X2 U4894 ( .B1(n8845), .B2(n8843), .A(n8842), .ZN(n8905) );
  NOR2_X2 U4895 ( .A1(n5886), .A2(n5885), .ZN(n8842) );
  NOR3_X2 U4896 ( .A1(n8965), .A2(n5913), .A3(n5912), .ZN(n7704) );
  INV_X1 U4897 ( .A(SI_16_), .ZN(n5186) );
  OR2_X1 U4898 ( .A1(n9423), .A2(n9089), .ZN(n5548) );
  NAND2_X1 U4899 ( .A1(n5470), .A2(n5469), .ZN(n5497) );
  AND2_X1 U4900 ( .A1(n5431), .A2(n5430), .ZN(n9143) );
  NAND2_X1 U4901 ( .A1(n4524), .A2(n4522), .ZN(n8207) );
  AOI21_X1 U4902 ( .B1(n8201), .B2(n8295), .A(n4523), .ZN(n4522) );
  NAND2_X1 U4903 ( .A1(n4525), .A2(n8195), .ZN(n4524) );
  AND2_X1 U4904 ( .A1(n8200), .A2(n8280), .ZN(n4523) );
  INV_X1 U4905 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4880) );
  INV_X1 U4906 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4650) );
  INV_X1 U4907 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4649) );
  NOR2_X1 U4908 ( .A1(n4475), .A2(n4471), .ZN(n4470) );
  INV_X1 U4909 ( .A(n7575), .ZN(n4471) );
  INV_X1 U4910 ( .A(n4760), .ZN(n4475) );
  OR2_X1 U4911 ( .A1(n8745), .A2(n8751), .ZN(n4559) );
  AND2_X1 U4912 ( .A1(n4410), .A2(n4409), .ZN(n4408) );
  INV_X1 U4913 ( .A(n4806), .ZN(n4413) );
  NOR2_X1 U4914 ( .A1(n8660), .A2(n8786), .ZN(n8090) );
  NAND2_X1 U4915 ( .A1(n4564), .A2(n9888), .ZN(n4563) );
  NOR2_X1 U4916 ( .A1(n4565), .A2(n8797), .ZN(n4564) );
  AND2_X1 U4917 ( .A1(n9749), .A2(n8182), .ZN(n4642) );
  AND2_X1 U4918 ( .A1(n7509), .A2(n7507), .ZN(n4827) );
  INV_X1 U4919 ( .A(n9737), .ZN(n7509) );
  OR2_X1 U4920 ( .A1(n8720), .A2(n8420), .ZN(n8279) );
  NOR2_X1 U4921 ( .A1(n8740), .A2(n4559), .ZN(n4558) );
  AND3_X1 U4922 ( .A1(n4330), .A2(n4502), .A3(n4813), .ZN(n6298) );
  INV_X1 U4923 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4501) );
  INV_X1 U4924 ( .A(n9540), .ZN(n4856) );
  AND2_X1 U4925 ( .A1(n6999), .A2(n6998), .ZN(n7002) );
  OAI21_X1 U4926 ( .B1(n5390), .B2(n5389), .A(n5388), .ZN(n5414) );
  AND2_X1 U4927 ( .A1(n5205), .A2(n5189), .ZN(n5203) );
  INV_X1 U4928 ( .A(n4685), .ZN(n4684) );
  AOI21_X1 U4929 ( .B1(n4685), .B2(n4683), .A(n4682), .ZN(n4681) );
  INV_X1 U4930 ( .A(n4888), .ZN(n6442) );
  AND2_X1 U4931 ( .A1(n7709), .A2(n7128), .ZN(n4755) );
  OR2_X1 U4932 ( .A1(n8041), .A2(n4483), .ZN(n4482) );
  INV_X1 U4933 ( .A(n7807), .ZN(n4483) );
  NAND2_X1 U4934 ( .A1(n7012), .A2(n4276), .ZN(n7017) );
  AND2_X1 U4935 ( .A1(n6931), .A2(n6925), .ZN(n4505) );
  NAND2_X1 U4936 ( .A1(n6449), .A2(n8389), .ZN(n6679) );
  AOI21_X1 U4937 ( .B1(n8424), .B2(n4634), .A(n4629), .ZN(n8116) );
  NOR2_X1 U4938 ( .A1(n8119), .A2(n4635), .ZN(n4634) );
  NAND2_X1 U4939 ( .A1(n4630), .A2(n4298), .ZN(n4629) );
  AOI21_X1 U4940 ( .B1(n8299), .B2(n8298), .A(n8297), .ZN(n4541) );
  OR2_X1 U4941 ( .A1(n6470), .A2(n6877), .ZN(n6676) );
  NAND2_X1 U4942 ( .A1(n4801), .A2(n4799), .ZN(n4798) );
  NAND2_X1 U4943 ( .A1(n8421), .A2(n4804), .ZN(n4799) );
  OR2_X1 U4944 ( .A1(n4801), .A2(n8422), .ZN(n4797) );
  AND2_X1 U4945 ( .A1(n8456), .A2(n8448), .ZN(n8444) );
  AOI21_X1 U4946 ( .B1(n4824), .B2(n4823), .A(n4306), .ZN(n4822) );
  AOI22_X1 U4947 ( .A1(n8525), .A2(n8417), .B1(n8416), .B2(n8530), .ZN(n8520)
         );
  INV_X2 U4948 ( .A(n6815), .ZN(n8110) );
  INV_X1 U4949 ( .A(n8111), .ZN(n7795) );
  INV_X1 U4950 ( .A(n6768), .ZN(n7794) );
  NAND2_X1 U4951 ( .A1(n6768), .A2(n6445), .ZN(n6817) );
  AND2_X1 U4952 ( .A1(n4819), .A2(n5973), .ZN(n4553) );
  NAND2_X1 U4953 ( .A1(n5954), .A2(n6759), .ZN(n4699) );
  NAND2_X1 U4954 ( .A1(n5496), .A2(n5504), .ZN(n5610) );
  NAND2_X1 U4955 ( .A1(n9540), .A2(n4862), .ZN(n5355) );
  NAND2_X1 U4956 ( .A1(n5502), .A2(n5501), .ZN(n9417) );
  NOR2_X1 U4957 ( .A1(n5550), .A2(n5646), .ZN(n9120) );
  NOR2_X1 U4958 ( .A1(n9139), .A2(n4764), .ZN(n4763) );
  INV_X1 U4959 ( .A(n9087), .ZN(n4764) );
  AOI21_X1 U4960 ( .B1(n9168), .B2(n9085), .A(n9084), .ZN(n9153) );
  NAND2_X1 U4961 ( .A1(n9082), .A2(n9081), .ZN(n9183) );
  INV_X1 U4962 ( .A(n9235), .ZN(n9203) );
  NAND2_X1 U4963 ( .A1(n9588), .A2(n9095), .ZN(n4577) );
  NAND2_X1 U4964 ( .A1(n7002), .A2(n7001), .ZN(n7091) );
  OR2_X1 U4965 ( .A1(n5947), .A2(n6707), .ZN(n9510) );
  NOR2_X1 U4966 ( .A1(n4492), .A2(n4491), .ZN(n4490) );
  INV_X1 U4967 ( .A(n7977), .ZN(n4491) );
  NOR2_X1 U4968 ( .A1(n4494), .A2(n4493), .ZN(n4492) );
  NAND2_X1 U4969 ( .A1(n9699), .A2(n9700), .ZN(n9698) );
  NAND2_X1 U4970 ( .A1(n6768), .A2(n4746), .ZN(n4745) );
  NAND2_X1 U4971 ( .A1(n4314), .A2(n4747), .ZN(n4746) );
  AND2_X1 U4972 ( .A1(n4665), .A2(n5657), .ZN(n4377) );
  NAND2_X1 U4973 ( .A1(n5604), .A2(n9250), .ZN(n4665) );
  OAI21_X1 U4974 ( .B1(n8168), .B2(n8280), .A(n8167), .ZN(n4510) );
  NAND2_X1 U4975 ( .A1(n4358), .A2(n4355), .ZN(n5157) );
  AND2_X1 U4976 ( .A1(n9579), .A2(n4356), .ZN(n4355) );
  NAND2_X1 U4977 ( .A1(n4359), .A2(n5511), .ZN(n4358) );
  NAND2_X1 U4978 ( .A1(n4357), .A2(n5947), .ZN(n4356) );
  AOI21_X1 U4979 ( .B1(n8207), .B2(n8204), .A(n8203), .ZN(n8206) );
  NAND2_X1 U4980 ( .A1(n4369), .A2(n4366), .ZN(n4365) );
  OAI21_X1 U4981 ( .B1(n5159), .B2(n5577), .A(n4370), .ZN(n4369) );
  AOI21_X1 U4982 ( .B1(n5156), .B2(n4368), .A(n4367), .ZN(n4366) );
  NOR2_X1 U4983 ( .A1(n4371), .A2(n5947), .ZN(n4370) );
  NAND2_X1 U4984 ( .A1(n4518), .A2(n4516), .ZN(n4515) );
  NOR2_X1 U4985 ( .A1(n8643), .A2(n4517), .ZN(n4516) );
  NAND2_X1 U4986 ( .A1(n4519), .A2(n4301), .ZN(n4518) );
  INV_X1 U4987 ( .A(n8220), .ZN(n4517) );
  NAND2_X1 U4988 ( .A1(n4364), .A2(n4363), .ZN(n5381) );
  NAND2_X1 U4989 ( .A1(n5286), .A2(n5947), .ZN(n4363) );
  NAND2_X1 U4990 ( .A1(n5285), .A2(n5511), .ZN(n4364) );
  INV_X1 U4991 ( .A(n8276), .ZN(n4550) );
  NAND2_X1 U4992 ( .A1(n4361), .A2(n5589), .ZN(n5384) );
  INV_X1 U4993 ( .A(n4533), .ZN(n4531) );
  INV_X1 U4994 ( .A(n8579), .ZN(n4409) );
  INV_X1 U4995 ( .A(n5503), .ZN(n5510) );
  INV_X1 U4996 ( .A(n4656), .ZN(n4655) );
  OAI21_X1 U4997 ( .B1(n4989), .B2(n4657), .A(n5004), .ZN(n4656) );
  INV_X1 U4998 ( .A(n4900), .ZN(n4657) );
  INV_X1 U4999 ( .A(n7990), .ZN(n4478) );
  INV_X1 U5000 ( .A(n4482), .ZN(n4479) );
  INV_X1 U5001 ( .A(n7719), .ZN(n4474) );
  NAND2_X1 U5002 ( .A1(n4636), .A2(n8285), .ZN(n4635) );
  NAND2_X1 U5003 ( .A1(n8396), .A2(n4637), .ZN(n4636) );
  NAND2_X1 U5004 ( .A1(n4562), .A2(n8460), .ZN(n4561) );
  NOR2_X1 U5005 ( .A1(n8720), .A2(n8391), .ZN(n4562) );
  OR2_X1 U5006 ( .A1(n8751), .A2(n8416), .ZN(n8238) );
  OR2_X1 U5007 ( .A1(n8761), .A2(n8092), .ZN(n8247) );
  OR2_X1 U5008 ( .A1(n8791), .A2(n8668), .ZN(n8218) );
  NAND2_X1 U5009 ( .A1(n7340), .A2(n4642), .ZN(n9761) );
  NAND2_X1 U5010 ( .A1(n7181), .A2(n8315), .ZN(n8150) );
  NAND2_X1 U5011 ( .A1(n4558), .A2(n8491), .ZN(n4557) );
  XNOR2_X1 U5012 ( .A(n8317), .B(n8147), .ZN(n6837) );
  OR2_X1 U5013 ( .A1(n6414), .A2(n7569), .ZN(n6433) );
  AND2_X1 U5014 ( .A1(n7469), .A2(n6413), .ZN(n6414) );
  INV_X1 U5015 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6231) );
  NOR2_X1 U5016 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4817) );
  NAND2_X1 U5017 ( .A1(n7432), .A2(n4717), .ZN(n4716) );
  INV_X1 U5018 ( .A(n5742), .ZN(n4717) );
  OR2_X1 U5019 ( .A1(n9427), .A2(n9143), .ZN(n9140) );
  OR2_X1 U5020 ( .A1(n9430), .A2(n9158), .ZN(n5641) );
  AND2_X1 U5021 ( .A1(n9430), .A2(n9158), .ZN(n9116) );
  NOR2_X1 U5022 ( .A1(n4585), .A2(n9105), .ZN(n4579) );
  NAND2_X1 U5023 ( .A1(n4586), .A2(n4587), .ZN(n4585) );
  NOR2_X1 U5024 ( .A1(n9458), .A2(n4441), .ZN(n4440) );
  INV_X1 U5025 ( .A(n4442), .ZN(n4441) );
  INV_X1 U5026 ( .A(n4770), .ZN(n4768) );
  NAND2_X1 U5027 ( .A1(n4588), .A2(n9106), .ZN(n4587) );
  INV_X1 U5028 ( .A(n9272), .ZN(n4588) );
  NAND2_X1 U5029 ( .A1(n4590), .A2(n9106), .ZN(n4589) );
  NOR2_X1 U5030 ( .A1(n9352), .A2(n4788), .ZN(n4787) );
  INV_X1 U5031 ( .A(n9062), .ZN(n4788) );
  NAND2_X1 U5032 ( .A1(n6861), .A2(n4941), .ZN(n6711) );
  NOR2_X1 U5033 ( .A1(n9159), .A2(n9423), .ZN(n9145) );
  NOR2_X1 U5034 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4793) );
  NAND2_X1 U5035 ( .A1(n4869), .A2(n4352), .ZN(n4871) );
  NOR2_X1 U5036 ( .A1(n4870), .A2(n9535), .ZN(n4352) );
  INV_X1 U5037 ( .A(n5439), .ZN(n4664) );
  AOI21_X1 U5038 ( .B1(n5439), .B2(n4663), .A(n4662), .ZN(n4661) );
  INV_X1 U5039 ( .A(n5441), .ZN(n4662) );
  INV_X1 U5040 ( .A(n5415), .ZN(n4663) );
  INV_X1 U5041 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5659) );
  OAI21_X1 U5042 ( .B1(n5360), .B2(n4690), .A(n5363), .ZN(n5390) );
  INV_X1 U5043 ( .A(n5361), .ZN(n4690) );
  OAI21_X1 U5044 ( .B1(n5307), .B2(n5306), .A(n5305), .ZN(n5324) );
  OAI21_X1 U5045 ( .B1(n5265), .B2(n5264), .A(n5266), .ZN(n5288) );
  AND2_X1 U5046 ( .A1(n5289), .A2(n5270), .ZN(n5287) );
  INV_X1 U5047 ( .A(n4695), .ZN(n4694) );
  NOR2_X1 U5048 ( .A1(n5183), .A2(n4698), .ZN(n4697) );
  INV_X1 U5049 ( .A(n5163), .ZN(n4698) );
  AOI21_X1 U5050 ( .B1(n4697), .B2(n5164), .A(n4696), .ZN(n4695) );
  INV_X1 U5051 ( .A(n5185), .ZN(n4696) );
  AND2_X1 U5052 ( .A1(n4781), .A2(n4840), .ZN(n4598) );
  NAND2_X1 U5053 ( .A1(n4430), .A2(n4429), .ZN(n4783) );
  INV_X1 U5054 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4430) );
  INV_X1 U5055 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4429) );
  OAI211_X1 U5056 ( .C1(n4533), .C2(n4375), .A(n4374), .B(n4372), .ZN(n4887)
         );
  NAND2_X1 U5057 ( .A1(n4373), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4372) );
  XNOR2_X1 U5058 ( .A(n4887), .B(SI_2_), .ZN(n4947) );
  AND2_X1 U5059 ( .A1(n7734), .A2(n7724), .ZN(n4760) );
  INV_X1 U5060 ( .A(n4481), .ZN(n4480) );
  OAI21_X1 U5061 ( .B1(n4756), .B2(n4482), .A(n7825), .ZN(n4481) );
  NAND2_X1 U5062 ( .A1(n8060), .A2(n8061), .ZN(n4758) );
  OAI21_X1 U5063 ( .B1(n8051), .B2(n4736), .A(n4304), .ZN(n7877) );
  OR2_X1 U5064 ( .A1(n7851), .A2(n4738), .ZN(n4736) );
  NOR2_X1 U5065 ( .A1(n7864), .A2(n4739), .ZN(n4738) );
  AND2_X1 U5066 ( .A1(n6219), .A2(n6218), .ZN(n6462) );
  NOR2_X1 U5067 ( .A1(n6574), .A2(n6573), .ZN(n6572) );
  OR2_X1 U5068 ( .A1(n6572), .A2(n4457), .ZN(n4456) );
  AND2_X1 U5069 ( .A1(n6522), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4457) );
  NAND2_X1 U5070 ( .A1(n4456), .A2(n4455), .ZN(n4454) );
  INV_X1 U5071 ( .A(n6603), .ZN(n4455) );
  NOR2_X1 U5072 ( .A1(n6584), .A2(n6583), .ZN(n6582) );
  OR2_X1 U5073 ( .A1(n6582), .A2(n4452), .ZN(n4451) );
  NOR2_X1 U5074 ( .A1(n7112), .A2(n6527), .ZN(n4452) );
  AND2_X1 U5075 ( .A1(n4451), .A2(n4450), .ZN(n6622) );
  INV_X1 U5076 ( .A(n6623), .ZN(n4450) );
  NAND2_X1 U5077 ( .A1(n7417), .A2(n4461), .ZN(n8321) );
  OR2_X1 U5078 ( .A1(n7726), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4461) );
  NOR3_X1 U5079 ( .A1(n8474), .A2(n4561), .A3(n8396), .ZN(n8395) );
  AOI21_X1 U5080 ( .B1(n4803), .B2(n4264), .A(n4308), .ZN(n4801) );
  NAND2_X1 U5081 ( .A1(n4614), .A2(n8500), .ZN(n4613) );
  INV_X1 U5082 ( .A(n4617), .ZN(n4616) );
  OAI21_X1 U5083 ( .B1(n8471), .B2(n8272), .A(n8273), .ZN(n4617) );
  NAND2_X1 U5084 ( .A1(n8418), .A2(n8500), .ZN(n4826) );
  INV_X1 U5085 ( .A(n4612), .ZN(n4610) );
  NAND2_X1 U5086 ( .A1(n8521), .A2(n4332), .ZN(n8495) );
  NOR2_X1 U5087 ( .A1(n8527), .A2(n8751), .ZN(n8526) );
  NAND2_X1 U5088 ( .A1(n8546), .A2(n8536), .ZN(n4349) );
  OR2_X1 U5089 ( .A1(n8546), .A2(n8536), .ZN(n4835) );
  NAND2_X1 U5090 ( .A1(n4315), .A2(n4413), .ZN(n4410) );
  NOR2_X1 U5091 ( .A1(n8412), .A2(n8620), .ZN(n4412) );
  NAND2_X1 U5092 ( .A1(n4413), .A2(n4414), .ZN(n4411) );
  AND2_X1 U5093 ( .A1(n4623), .A2(n4620), .ZN(n4619) );
  NAND2_X1 U5094 ( .A1(n4284), .A2(n8643), .ZN(n4620) );
  NAND2_X1 U5095 ( .A1(n4810), .A2(n8619), .ZN(n4809) );
  INV_X1 U5096 ( .A(n8778), .ZN(n4810) );
  INV_X1 U5097 ( .A(n8090), .ZN(n4627) );
  AOI21_X1 U5098 ( .B1(n8621), .B2(n8620), .A(n8412), .ZN(n8604) );
  NAND2_X1 U5099 ( .A1(n8604), .A2(n8603), .ZN(n8602) );
  AND2_X1 U5100 ( .A1(n8216), .A2(n8215), .ZN(n8670) );
  OR2_X1 U5101 ( .A1(n8400), .A2(n7516), .ZN(n4565) );
  NAND2_X1 U5102 ( .A1(n6483), .A2(n6461), .ZN(n8692) );
  NAND2_X1 U5103 ( .A1(n4640), .A2(n8191), .ZN(n4639) );
  NAND2_X1 U5104 ( .A1(n7512), .A2(n4641), .ZN(n4640) );
  NAND2_X1 U5105 ( .A1(n7508), .A2(n7507), .ZN(n9725) );
  OR2_X1 U5106 ( .A1(n9753), .A2(n9864), .ZN(n9728) );
  NAND2_X1 U5107 ( .A1(n9751), .A2(n9858), .ZN(n9753) );
  NAND2_X1 U5108 ( .A1(n7021), .A2(n8316), .ZN(n8149) );
  AND2_X1 U5109 ( .A1(n8117), .A2(n6730), .ZN(n8690) );
  INV_X1 U5110 ( .A(n8694), .ZN(n9764) );
  INV_X1 U5111 ( .A(n8690), .ZN(n9769) );
  NAND2_X1 U5112 ( .A1(n7738), .A2(n7737), .ZN(n8781) );
  NAND2_X1 U5113 ( .A1(n4313), .A2(n4819), .ZN(n4818) );
  INV_X1 U5114 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6077) );
  INV_X1 U5115 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6417) );
  INV_X1 U5116 ( .A(n4500), .ZN(n4499) );
  OAI21_X1 U5117 ( .B1(n6378), .B2(n6071), .A(n6415), .ZN(n4500) );
  INV_X1 U5118 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6297) );
  NOR2_X1 U5119 ( .A1(n6044), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6057) );
  NOR2_X1 U5120 ( .A1(n4706), .A2(n4703), .ZN(n4702) );
  NOR2_X1 U5121 ( .A1(n8924), .A2(n8923), .ZN(n4706) );
  INV_X1 U5122 ( .A(n8874), .ZN(n4703) );
  AND2_X1 U5123 ( .A1(n5892), .A2(n8904), .ZN(n4727) );
  INV_X1 U5124 ( .A(n5195), .ZN(n5193) );
  AND2_X1 U5125 ( .A1(n5889), .A2(n5888), .ZN(n5890) );
  NAND2_X1 U5126 ( .A1(n4712), .A2(n5764), .ZN(n7628) );
  INV_X1 U5127 ( .A(n7627), .ZN(n4712) );
  AOI21_X1 U5128 ( .B1(n5674), .B2(n5710), .A(n5673), .ZN(n6252) );
  INV_X1 U5129 ( .A(n8865), .ZN(n4724) );
  NAND2_X1 U5130 ( .A1(n8913), .A2(n8915), .ZN(n4721) );
  NOR2_X1 U5131 ( .A1(n4724), .A2(n5865), .ZN(n4723) );
  AND2_X1 U5132 ( .A1(n4671), .A2(n4669), .ZN(n5608) );
  NAND2_X1 U5133 ( .A1(n5508), .A2(n5947), .ZN(n4671) );
  NOR2_X1 U5134 ( .A1(n4670), .A2(n5516), .ZN(n4669) );
  INV_X1 U5135 ( .A(n4955), .ZN(n5481) );
  INV_X1 U5136 ( .A(n4969), .ZN(n5459) );
  NAND2_X1 U5137 ( .A1(n9612), .A2(n4385), .ZN(n6691) );
  NAND2_X1 U5138 ( .A1(n4387), .A2(n4386), .ZN(n4385) );
  INV_X1 U5139 ( .A(n9609), .ZN(n4387) );
  NOR2_X1 U5140 ( .A1(n6691), .A2(n6692), .ZN(n6690) );
  NOR2_X1 U5141 ( .A1(n6307), .A2(n4399), .ZN(n6309) );
  AND2_X1 U5142 ( .A1(n6308), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4399) );
  OR2_X1 U5143 ( .A1(n6309), .A2(n6310), .ZN(n4398) );
  NOR2_X1 U5144 ( .A1(n6953), .A2(n4400), .ZN(n7270) );
  AND2_X1 U5145 ( .A1(n6954), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4400) );
  NAND2_X1 U5146 ( .A1(n9145), .A2(n9129), .ZN(n9125) );
  OR2_X1 U5147 ( .A1(n9435), .A2(n9204), .ZN(n9173) );
  AND2_X1 U5148 ( .A1(n9447), .A2(n9235), .ZN(n9078) );
  INV_X1 U5149 ( .A(n4587), .ZN(n4581) );
  INV_X1 U5150 ( .A(n4589), .ZN(n4582) );
  AOI21_X1 U5151 ( .B1(n4772), .B2(n4277), .A(n4771), .ZN(n4770) );
  NOR2_X1 U5152 ( .A1(n9282), .A2(n9263), .ZN(n4771) );
  INV_X1 U5153 ( .A(n9072), .ZN(n4772) );
  NOR2_X1 U5154 ( .A1(n9294), .A2(n9072), .ZN(n4773) );
  AOI21_X1 U5155 ( .B1(n4593), .B2(n9103), .A(n4591), .ZN(n4590) );
  INV_X1 U5156 ( .A(n9104), .ZN(n4591) );
  AND2_X1 U5157 ( .A1(n5524), .A2(n9106), .ZN(n9272) );
  AND2_X1 U5158 ( .A1(n9098), .A2(n5558), .ZN(n9352) );
  NAND2_X1 U5159 ( .A1(n9063), .A2(n4787), .ZN(n9349) );
  NOR2_X1 U5160 ( .A1(n9368), .A2(n4576), .ZN(n4575) );
  INV_X1 U5161 ( .A(n9096), .ZN(n4576) );
  NAND2_X1 U5162 ( .A1(n4577), .A2(n9096), .ZN(n9369) );
  NOR2_X1 U5163 ( .A1(n9579), .A2(n4776), .ZN(n4775) );
  INV_X1 U5164 ( .A(n9054), .ZN(n4776) );
  NAND2_X1 U5165 ( .A1(n9094), .A2(n9093), .ZN(n9588) );
  NOR2_X1 U5166 ( .A1(n7478), .A2(n4779), .ZN(n4778) );
  INV_X1 U5167 ( .A(n7475), .ZN(n4779) );
  NAND2_X1 U5168 ( .A1(n7095), .A2(n7094), .ZN(n7476) );
  INV_X1 U5169 ( .A(n7359), .ZN(n7092) );
  AND2_X1 U5170 ( .A1(n5624), .A2(n7085), .ZN(n7359) );
  INV_X1 U5171 ( .A(n5670), .ZN(n6284) );
  INV_X1 U5172 ( .A(n9311), .ZN(n9638) );
  INV_X1 U5173 ( .A(n5529), .ZN(n6699) );
  NAND2_X1 U5174 ( .A1(n9125), .A2(n4438), .ZN(n9415) );
  OR2_X1 U5175 ( .A1(n9145), .A2(n9129), .ZN(n4438) );
  AND2_X1 U5176 ( .A1(n9417), .A2(n9568), .ZN(n4436) );
  INV_X1 U5177 ( .A(n9172), .ZN(n9430) );
  NAND2_X1 U5178 ( .A1(n5130), .A2(n5129), .ZN(n9499) );
  NAND2_X1 U5179 ( .A1(n5106), .A2(n5105), .ZN(n9506) );
  NAND2_X1 U5180 ( .A1(n5678), .A2(n5670), .ZN(n6881) );
  AOI21_X1 U5181 ( .B1(n4675), .B2(n4679), .A(n4673), .ZN(n4672) );
  INV_X1 U5182 ( .A(n5488), .ZN(n4673) );
  NAND2_X1 U5183 ( .A1(n4677), .A2(n4678), .ZN(n5490) );
  OR2_X1 U5184 ( .A1(n5497), .A2(n4679), .ZN(n4677) );
  NAND2_X1 U5185 ( .A1(n4434), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4602) );
  XNOR2_X1 U5186 ( .A(n5414), .B(n5413), .ZN(n7894) );
  NAND2_X1 U5187 ( .A1(n4281), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U5188 ( .A1(n4850), .A2(n4599), .ZN(n4433) );
  NAND2_X1 U5189 ( .A1(n5661), .A2(n5659), .ZN(n5663) );
  AND2_X1 U5190 ( .A1(n5330), .A2(n5329), .ZN(n5344) );
  NAND2_X1 U5191 ( .A1(n5067), .A2(n4735), .ZN(n4734) );
  NAND2_X1 U5192 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n4735) );
  OAI21_X1 U5193 ( .B1(n5165), .B2(n5164), .A(n5163), .ZN(n5184) );
  NOR2_X1 U5194 ( .A1(n5116), .A2(n4688), .ZN(n4687) );
  INV_X1 U5195 ( .A(n5097), .ZN(n4688) );
  AOI21_X1 U5196 ( .B1(n4687), .B2(n5098), .A(n4686), .ZN(n4685) );
  INV_X1 U5197 ( .A(n5118), .ZN(n4686) );
  AND2_X1 U5198 ( .A1(n4879), .A2(n5085), .ZN(n6404) );
  OR3_X1 U5199 ( .A1(n7354), .A2(n7569), .A3(n7469), .ZN(n6480) );
  AND2_X1 U5200 ( .A1(n6910), .A2(n6911), .ZN(n7014) );
  NAND2_X1 U5201 ( .A1(n7797), .A2(n7796), .ZN(n8767) );
  NOR2_X1 U5202 ( .A1(n4486), .A2(n4488), .ZN(n4485) );
  NOR2_X1 U5203 ( .A1(n4489), .A2(n7978), .ZN(n4488) );
  INV_X1 U5204 ( .A(n4490), .ZN(n4486) );
  INV_X1 U5205 ( .A(n7976), .ZN(n4493) );
  NAND2_X1 U5206 ( .A1(n7129), .A2(n4755), .ZN(n7708) );
  INV_X1 U5207 ( .A(n4751), .ZN(n4750) );
  AND2_X1 U5208 ( .A1(n6733), .A2(n6732), .ZN(n9700) );
  INV_X1 U5209 ( .A(n7181), .ZN(n8017) );
  NAND2_X1 U5210 ( .A1(n7013), .A2(n7014), .ZN(n7012) );
  NAND2_X1 U5211 ( .A1(n7580), .A2(n7579), .ZN(n8797) );
  NOR2_X1 U5212 ( .A1(n8071), .A2(n8692), .ZN(n7985) );
  INV_X1 U5213 ( .A(n8085), .ZN(n9709) );
  NOR2_X1 U5214 ( .A1(n6941), .A2(P2_U3152), .ZN(n8073) );
  NAND2_X1 U5215 ( .A1(n6678), .A2(n6677), .ZN(n8085) );
  INV_X1 U5216 ( .A(n8692), .ZN(n9762) );
  OAI21_X1 U5217 ( .B1(n4541), .B2(n4540), .A(n4539), .ZN(n4538) );
  INV_X1 U5218 ( .A(n8301), .ZN(n4540) );
  NAND2_X1 U5219 ( .A1(n8303), .A2(n8302), .ZN(n4539) );
  INV_X1 U5220 ( .A(n9716), .ZN(n9714) );
  NAND2_X1 U5221 ( .A1(n8113), .A2(n8112), .ZN(n8705) );
  OR2_X1 U5222 ( .A1(n9782), .A2(n6674), .ZN(n8613) );
  INV_X1 U5223 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n4423) );
  INV_X1 U5224 ( .A(n8722), .ZN(n4425) );
  NAND2_X1 U5225 ( .A1(n8451), .A2(n4264), .ZN(n4419) );
  OR2_X1 U5226 ( .A1(n6081), .A2(n6080), .ZN(n4427) );
  AND3_X1 U5227 ( .A1(n5022), .A2(n5021), .A3(n5020), .ZN(n9675) );
  INV_X1 U5228 ( .A(n9225), .ZN(n9447) );
  AND4_X1 U5229 ( .A1(n5114), .A2(n5113), .A3(n5112), .A4(n5111), .ZN(n9589)
         );
  AND4_X1 U5230 ( .A1(n5299), .A2(n5298), .A3(n5297), .A4(n5296), .ZN(n9262)
         );
  NAND2_X1 U5231 ( .A1(n5233), .A2(n5232), .ZN(n9471) );
  AND2_X1 U5232 ( .A1(n5950), .A2(n9245), .ZN(n8977) );
  AND4_X1 U5233 ( .A1(n5154), .A2(n5153), .A3(n5152), .A4(n5151), .ZN(n9373)
         );
  NAND2_X1 U5234 ( .A1(n4668), .A2(n4667), .ZN(n4666) );
  NOR2_X1 U5235 ( .A1(n5601), .A2(n9250), .ZN(n4667) );
  NAND2_X1 U5236 ( .A1(n5608), .A2(n6717), .ZN(n4668) );
  AOI21_X1 U5237 ( .B1(n4838), .B2(n6759), .A(n7151), .ZN(n5657) );
  INV_X1 U5238 ( .A(n7379), .ZN(n9000) );
  NAND2_X1 U5239 ( .A1(n4393), .A2(n4392), .ZN(n4391) );
  NAND2_X1 U5240 ( .A1(n9034), .A2(n9623), .ZN(n4392) );
  OR2_X1 U5241 ( .A1(n9534), .A2(n6442), .ZN(n4652) );
  NAND2_X1 U5242 ( .A1(n9136), .A2(n9091), .ZN(n9092) );
  AND2_X1 U5243 ( .A1(n9136), .A2(n9135), .ZN(n9420) );
  NAND2_X1 U5244 ( .A1(n9088), .A2(n9087), .ZN(n9134) );
  NAND2_X1 U5245 ( .A1(n4597), .A2(n4594), .ZN(n9421) );
  NOR2_X1 U5246 ( .A1(n4596), .A2(n4595), .ZN(n4594) );
  OAI21_X1 U5247 ( .B1(n9141), .B2(n9142), .A(n9640), .ZN(n4597) );
  NOR2_X1 U5248 ( .A1(n9144), .A2(n9635), .ZN(n4596) );
  NAND2_X1 U5249 ( .A1(n4507), .A2(n4506), .ZN(n8196) );
  AND2_X1 U5250 ( .A1(n8181), .A2(n8180), .ZN(n4506) );
  NAND2_X1 U5251 ( .A1(n4509), .A2(n4508), .ZN(n4507) );
  INV_X1 U5252 ( .A(n5533), .ZN(n4357) );
  INV_X1 U5253 ( .A(n4360), .ZN(n4359) );
  AOI21_X1 U5254 ( .B1(n5062), .B2(n7610), .A(n7616), .ZN(n4360) );
  NAND2_X1 U5255 ( .A1(n4527), .A2(n4526), .ZN(n4525) );
  AOI21_X1 U5256 ( .B1(n8187), .B2(n8295), .A(n8189), .ZN(n4526) );
  NAND2_X1 U5257 ( .A1(n8188), .A2(n8280), .ZN(n4527) );
  AND2_X1 U5258 ( .A1(n9098), .A2(n5947), .ZN(n4368) );
  NAND2_X1 U5259 ( .A1(n5157), .A2(n9095), .ZN(n5158) );
  NAND2_X1 U5260 ( .A1(n4521), .A2(n4520), .ZN(n4519) );
  AOI21_X1 U5261 ( .B1(n8213), .B2(n8295), .A(n8667), .ZN(n4521) );
  NAND2_X1 U5262 ( .A1(n8214), .A2(n8280), .ZN(n4520) );
  AOI21_X1 U5263 ( .B1(n4365), .B2(n5222), .A(n5221), .ZN(n5245) );
  AOI21_X1 U5264 ( .B1(n4515), .B2(n8223), .A(n8620), .ZN(n8232) );
  OAI22_X1 U5265 ( .A1(n4362), .A2(n5383), .B1(n5382), .B2(n9110), .ZN(n4361)
         );
  AOI21_X1 U5266 ( .B1(n5381), .B2(n5523), .A(n9109), .ZN(n4362) );
  NAND2_X1 U5267 ( .A1(n4311), .A2(n4267), .ZN(n4545) );
  NOR2_X1 U5268 ( .A1(n4549), .A2(n4547), .ZN(n4546) );
  NAND2_X1 U5269 ( .A1(n8273), .A2(n8295), .ZN(n4547) );
  NOR2_X1 U5270 ( .A1(n4549), .A2(n4303), .ZN(n4548) );
  NOR2_X1 U5271 ( .A1(n4638), .A2(n6877), .ZN(n4637) );
  NAND2_X1 U5272 ( .A1(n8606), .A2(n4809), .ZN(n4807) );
  INV_X1 U5273 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5970) );
  INV_X1 U5274 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5959) );
  AND2_X1 U5275 ( .A1(n5458), .A2(n5457), .ZN(n5503) );
  AOI21_X1 U5276 ( .B1(n5416), .B2(n4661), .A(n4659), .ZN(n4658) );
  NAND2_X1 U5277 ( .A1(n4660), .A2(n5465), .ZN(n4659) );
  NAND2_X1 U5278 ( .A1(n4661), .A2(n4664), .ZN(n4660) );
  INV_X1 U5279 ( .A(n4599), .ZN(n4345) );
  NAND2_X1 U5280 ( .A1(n4695), .A2(n4693), .ZN(n4692) );
  INV_X1 U5281 ( .A(n4697), .ZN(n4693) );
  INV_X1 U5282 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5207) );
  INV_X1 U5283 ( .A(SI_15_), .ZN(n5166) );
  INV_X1 U5284 ( .A(n4836), .ZN(n4682) );
  INV_X1 U5285 ( .A(n4687), .ZN(n4683) );
  NAND2_X1 U5286 ( .A1(n4843), .A2(n4877), .ZN(n4844) );
  INV_X1 U5287 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n4843) );
  NAND2_X1 U5288 ( .A1(n4531), .A2(n4534), .ZN(n4530) );
  NAND2_X1 U5289 ( .A1(n4373), .A2(n4534), .ZN(n4528) );
  NAND2_X1 U5290 ( .A1(n4532), .A2(n4533), .ZN(n4888) );
  INV_X1 U5291 ( .A(n7949), .ZN(n4739) );
  NOR2_X1 U5292 ( .A1(n7960), .A2(n4757), .ZN(n4756) );
  INV_X1 U5293 ( .A(n7792), .ZN(n4757) );
  OR2_X1 U5294 ( .A1(n4631), .A2(n8119), .ZN(n4630) );
  NAND2_X1 U5295 ( .A1(n4633), .A2(n4632), .ZN(n4631) );
  INV_X1 U5296 ( .A(n4637), .ZN(n4632) );
  INV_X1 U5297 ( .A(n8289), .ZN(n4633) );
  OR2_X1 U5298 ( .A1(n8461), .A2(n4264), .ZN(n4805) );
  INV_X1 U5299 ( .A(n8281), .ZN(n4608) );
  INV_X1 U5300 ( .A(n4613), .ZN(n4609) );
  NAND2_X1 U5301 ( .A1(n8495), .A2(n4822), .ZN(n4403) );
  NOR2_X1 U5302 ( .A1(n8740), .A2(n8256), .ZN(n4612) );
  NAND2_X1 U5303 ( .A1(n4624), .A2(n8091), .ZN(n4623) );
  NAND2_X1 U5304 ( .A1(n8606), .A2(n8224), .ZN(n4624) );
  INV_X1 U5305 ( .A(n6676), .ZN(n6483) );
  INV_X1 U5306 ( .A(n8183), .ZN(n4641) );
  NAND2_X1 U5307 ( .A1(n4560), .A2(n9844), .ZN(n7214) );
  NAND2_X1 U5308 ( .A1(n7182), .A2(n8017), .ZN(n8155) );
  NAND2_X1 U5309 ( .A1(n9702), .A2(n9827), .ZN(n8171) );
  NAND2_X1 U5310 ( .A1(n6668), .A2(n6734), .ZN(n6452) );
  AOI21_X1 U5311 ( .B1(n6431), .B2(n6430), .A(n6433), .ZN(n7158) );
  INV_X1 U5312 ( .A(n9818), .ZN(n7154) );
  INV_X1 U5313 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4820) );
  NAND2_X1 U5314 ( .A1(n6019), .A2(n4816), .ZN(n6026) );
  NOR2_X1 U5315 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n4816) );
  INV_X1 U5316 ( .A(n5954), .ZN(n5675) );
  AND2_X1 U5317 ( .A1(n5509), .A2(n5511), .ZN(n4670) );
  NAND2_X1 U5318 ( .A1(n4383), .A2(n5547), .ZN(n5509) );
  NAND2_X1 U5319 ( .A1(n5503), .A2(n4384), .ZN(n4383) );
  NOR2_X1 U5320 ( .A1(n5597), .A2(n9144), .ZN(n4384) );
  NAND2_X1 U5321 ( .A1(n4651), .A2(n5486), .ZN(n5504) );
  NAND2_X1 U5322 ( .A1(n4942), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4934) );
  AND2_X1 U5323 ( .A1(n9417), .A2(n9144), .ZN(n5646) );
  OR2_X1 U5324 ( .A1(n5371), .A2(n5370), .ZN(n5400) );
  OR2_X1 U5325 ( .A1(n9442), .A2(n9218), .ZN(n5589) );
  OR2_X1 U5326 ( .A1(n5315), .A2(n5314), .ZN(n5351) );
  NOR2_X1 U5327 ( .A1(n9463), .A2(n9468), .ZN(n4442) );
  OR2_X1 U5328 ( .A1(n9458), .A2(n9262), .ZN(n9108) );
  NOR2_X1 U5329 ( .A1(n9487), .A2(n9495), .ZN(n4446) );
  INV_X1 U5330 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n4860) );
  OR2_X1 U5331 ( .A1(n4568), .A2(n4566), .ZN(n7611) );
  NAND2_X1 U5332 ( .A1(n4569), .A2(n4295), .ZN(n4566) );
  NOR2_X1 U5333 ( .A1(n7603), .A2(n7635), .ZN(n4435) );
  INV_X1 U5334 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5042) );
  OR2_X1 U5335 ( .A1(n5043), .A2(n5042), .ZN(n5045) );
  INV_X1 U5336 ( .A(n4570), .ZN(n4569) );
  OAI21_X1 U5337 ( .B1(n4571), .B2(n5569), .A(n7609), .ZN(n4570) );
  NOR2_X1 U5338 ( .A1(n7086), .A2(n4571), .ZN(n4568) );
  NOR2_X1 U5339 ( .A1(n7363), .A2(n7098), .ZN(n7484) );
  NOR2_X1 U5340 ( .A1(n7047), .A2(n7051), .ZN(n6971) );
  NAND2_X1 U5341 ( .A1(n6712), .A2(n6284), .ZN(n6292) );
  INV_X1 U5342 ( .A(n8948), .ZN(n6960) );
  NAND2_X1 U5343 ( .A1(n6858), .A2(n5529), .ZN(n6861) );
  NAND2_X1 U5344 ( .A1(n9287), .A2(n9282), .ZN(n9276) );
  NOR2_X1 U5345 ( .A1(n5489), .A2(n4676), .ZN(n4675) );
  INV_X1 U5346 ( .A(n4678), .ZN(n4676) );
  NOR2_X1 U5347 ( .A1(n5499), .A2(SI_29_), .ZN(n4679) );
  NAND2_X1 U5348 ( .A1(n5499), .A2(SI_29_), .ZN(n4678) );
  AND2_X1 U5349 ( .A1(n5441), .A2(n5421), .ZN(n5439) );
  NAND2_X1 U5350 ( .A1(n4689), .A2(n5250), .ZN(n5265) );
  AND2_X1 U5351 ( .A1(n5051), .A2(n4729), .ZN(n5124) );
  AOI21_X1 U5352 ( .B1(n4655), .B2(n4657), .A(n4312), .ZN(n4654) );
  NAND2_X1 U5353 ( .A1(n7922), .A2(n7909), .ZN(n4743) );
  NAND2_X1 U5354 ( .A1(n7720), .A2(n7719), .ZN(n4761) );
  OR2_X1 U5355 ( .A1(n7783), .A2(n8359), .ZN(n7815) );
  INV_X1 U5356 ( .A(n4494), .ZN(n4489) );
  NOR2_X1 U5357 ( .A1(n4495), .A2(n7966), .ZN(n4494) );
  INV_X1 U5358 ( .A(n4743), .ZN(n4495) );
  OAI21_X1 U5359 ( .B1(n4755), .B2(n4752), .A(n7146), .ZN(n4751) );
  NAND2_X1 U5360 ( .A1(n4758), .A2(n4756), .ZN(n7958) );
  AOI21_X1 U5361 ( .B1(n4476), .B2(n4269), .A(n4477), .ZN(n7848) );
  INV_X1 U5362 ( .A(n4758), .ZN(n4476) );
  AOI21_X1 U5363 ( .B1(n4760), .B2(n4474), .A(n4473), .ZN(n4472) );
  INV_X1 U5364 ( .A(n7735), .ZN(n4473) );
  AND2_X1 U5365 ( .A1(n6669), .A2(n8305), .ZN(n6678) );
  AOI21_X1 U5366 ( .B1(n6515), .B2(P2_REG1_REG_1__SCAN_IN), .A(n6560), .ZN(
        n9557) );
  NAND2_X1 U5367 ( .A1(n6524), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4453) );
  AOI21_X1 U5368 ( .B1(n6526), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6540), .ZN(
        n6584) );
  NOR2_X1 U5369 ( .A1(n6622), .A2(n4447), .ZN(n6551) );
  NOR2_X1 U5370 ( .A1(n4449), .A2(n4448), .ZN(n4447) );
  NOR2_X1 U5371 ( .A1(n6789), .A2(n4460), .ZN(n6532) );
  AND2_X1 U5372 ( .A1(n7453), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4460) );
  NAND2_X1 U5373 ( .A1(n6532), .A2(n6531), .ZN(n6804) );
  NAND2_X1 U5374 ( .A1(n6804), .A2(n4459), .ZN(n6805) );
  OR2_X1 U5375 ( .A1(n7539), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4459) );
  NAND2_X1 U5376 ( .A1(n6805), .A2(n6806), .ZN(n6978) );
  NOR2_X1 U5377 ( .A1(n8323), .A2(n8324), .ZN(n8326) );
  AOI21_X1 U5378 ( .B1(n8363), .B2(P2_REG1_REG_17__SCAN_IN), .A(n8362), .ZN(
        n8364) );
  OR2_X1 U5379 ( .A1(n8474), .A2(n4561), .ZN(n8430) );
  NAND2_X1 U5380 ( .A1(n8104), .A2(n8103), .ZN(n8396) );
  OR2_X1 U5381 ( .A1(n7899), .A2(n7898), .ZN(n7914) );
  OR2_X1 U5382 ( .A1(n7870), .A2(n8035), .ZN(n7899) );
  NOR2_X1 U5383 ( .A1(n8527), .A2(n4559), .ZN(n8513) );
  NAND2_X1 U5384 ( .A1(n8548), .A2(n8547), .ZN(n8531) );
  AND2_X1 U5385 ( .A1(n8246), .A2(n8533), .ZN(n8547) );
  AND2_X1 U5386 ( .A1(n4406), .A2(n4321), .ZN(n4405) );
  NAND2_X1 U5387 ( .A1(n8578), .A2(n8579), .ZN(n8577) );
  OAI21_X1 U5388 ( .B1(n8687), .B2(n8203), .A(n8210), .ZN(n8666) );
  AND2_X1 U5389 ( .A1(n8210), .A2(n8209), .ZN(n8688) );
  OR2_X1 U5390 ( .A1(n7319), .A2(n7318), .ZN(n7457) );
  NOR2_X1 U5391 ( .A1(n9728), .A2(n7516), .ZN(n9729) );
  AND2_X1 U5392 ( .A1(n8197), .A2(n8199), .ZN(n9737) );
  INV_X1 U5393 ( .A(n7338), .ZN(n4350) );
  NAND2_X1 U5394 ( .A1(n9761), .A2(n8183), .ZN(n7513) );
  NAND2_X1 U5395 ( .A1(n7340), .A2(n8182), .ZN(n9759) );
  NAND2_X1 U5396 ( .A1(n4605), .A2(n8153), .ZN(n7254) );
  INV_X1 U5397 ( .A(n8153), .ZN(n4604) );
  NAND2_X1 U5398 ( .A1(n6814), .A2(n6813), .ZN(n7260) );
  NAND2_X1 U5399 ( .A1(n6763), .A2(n4554), .ZN(n7234) );
  NAND2_X1 U5400 ( .A1(n6762), .A2(n6761), .ZN(n7233) );
  NAND2_X1 U5401 ( .A1(n6445), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4747) );
  OR2_X1 U5402 ( .A1(n9856), .A2(n6421), .ZN(n6674) );
  NAND2_X1 U5403 ( .A1(n7971), .A2(n7970), .ZN(n8720) );
  NOR2_X1 U5404 ( .A1(n8451), .A2(n4264), .ZN(n4420) );
  INV_X1 U5405 ( .A(n4558), .ZN(n4556) );
  NAND2_X1 U5406 ( .A1(n6679), .A2(n9822), .ZN(n9887) );
  INV_X1 U5407 ( .A(n9889), .ZN(n9836) );
  INV_X1 U5408 ( .A(n9887), .ZN(n9835) );
  INV_X1 U5409 ( .A(n6729), .ZN(n9822) );
  INV_X1 U5410 ( .A(n6433), .ZN(n9783) );
  INV_X1 U5411 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U5412 ( .A1(n5962), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U5413 ( .A1(n6084), .A2(n6083), .ZN(n5962) );
  XNOR2_X1 U5414 ( .A(n5979), .B(n5978), .ZN(n6670) );
  OAI21_X1 U5415 ( .B1(n6085), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6084) );
  INV_X1 U5416 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6083) );
  INV_X1 U5417 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5958) );
  AND2_X1 U5418 ( .A1(n4811), .A2(n4503), .ZN(n4502) );
  INV_X1 U5419 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4503) );
  INV_X1 U5420 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5961) );
  AND2_X1 U5421 ( .A1(n5905), .A2(n5904), .ZN(n5913) );
  OR2_X1 U5422 ( .A1(n5177), .A2(n7276), .ZN(n5195) );
  NAND2_X1 U5423 ( .A1(n4347), .A2(n4346), .ZN(n5841) );
  INV_X1 U5424 ( .A(n8894), .ZN(n4346) );
  INV_X1 U5425 ( .A(n7432), .ZN(n4718) );
  NOR2_X1 U5426 ( .A1(n8914), .A2(n8915), .ZN(n8912) );
  XNOR2_X1 U5427 ( .A(n5878), .B(n5900), .ZN(n8936) );
  CLKBUF_X1 U5428 ( .A(n6889), .Z(n6890) );
  NAND2_X1 U5429 ( .A1(n4280), .A2(n4316), .ZN(n4725) );
  OR2_X1 U5430 ( .A1(n6292), .A2(n5934), .ZN(n6253) );
  INV_X1 U5431 ( .A(n5678), .ZN(n6712) );
  OR2_X1 U5432 ( .A1(n7694), .A2(n5459), .ZN(n5454) );
  NOR2_X1 U5433 ( .A1(n4273), .A2(n4389), .ZN(n4388) );
  INV_X1 U5434 ( .A(n5988), .ZN(n4389) );
  INV_X1 U5435 ( .A(n6359), .ZN(n9615) );
  AND2_X1 U5436 ( .A1(n4398), .A2(n4397), .ZN(n6405) );
  NAND2_X1 U5437 ( .A1(n6404), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4397) );
  NAND2_X1 U5438 ( .A1(n6405), .A2(n6406), .ZN(n6640) );
  NOR2_X1 U5439 ( .A1(n7271), .A2(n7272), .ZN(n7490) );
  NAND2_X1 U5440 ( .A1(n9153), .A2(n9086), .ZN(n9088) );
  NOR2_X1 U5441 ( .A1(n9143), .A2(n9638), .ZN(n4595) );
  AND2_X1 U5442 ( .A1(n5407), .A2(n5406), .ZN(n9158) );
  OR2_X1 U5443 ( .A1(n8972), .A2(n5459), .ZN(n5407) );
  AOI21_X1 U5444 ( .B1(n9174), .B2(n9117), .A(n9116), .ZN(n9155) );
  NAND2_X1 U5445 ( .A1(n9155), .A2(n9154), .ZN(n9138) );
  NOR2_X1 U5446 ( .A1(n9184), .A2(n9430), .ZN(n9169) );
  NOR2_X1 U5447 ( .A1(n9219), .A2(n9442), .ZN(n9205) );
  AND2_X1 U5448 ( .A1(n5333), .A2(n5332), .ZN(n9080) );
  AOI21_X1 U5449 ( .B1(n9214), .B2(n9112), .A(n9111), .ZN(n9201) );
  NOR2_X1 U5450 ( .A1(n9201), .A2(n9200), .ZN(n9199) );
  AND2_X1 U5451 ( .A1(n9287), .A2(n4319), .ZN(n9229) );
  AND2_X1 U5452 ( .A1(n4584), .A2(n9107), .ZN(n4583) );
  NAND2_X1 U5453 ( .A1(n9287), .A2(n4440), .ZN(n9241) );
  OR2_X1 U5454 ( .A1(n4767), .A2(n9074), .ZN(n4766) );
  NOR2_X1 U5455 ( .A1(n4290), .A2(n4768), .ZN(n4767) );
  OR2_X1 U5456 ( .A1(n5236), .A2(n5235), .ZN(n5258) );
  AND2_X1 U5457 ( .A1(n9304), .A2(n9291), .ZN(n9287) );
  AND2_X1 U5458 ( .A1(n5242), .A2(n9292), .ZN(n9308) );
  AND2_X1 U5459 ( .A1(n9377), .A2(n4444), .ZN(n9304) );
  AND2_X1 U5460 ( .A1(n4265), .A2(n9069), .ZN(n4444) );
  AOI21_X1 U5461 ( .B1(n9335), .B2(n9101), .A(n9100), .ZN(n9317) );
  OAI21_X1 U5462 ( .B1(n9065), .B2(n4786), .A(n4785), .ZN(n4784) );
  INV_X1 U5463 ( .A(n9066), .ZN(n4785) );
  NAND2_X1 U5464 ( .A1(n9377), .A2(n4265), .ZN(n9324) );
  AND2_X1 U5465 ( .A1(n9377), .A2(n9361), .ZN(n9356) );
  NAND2_X1 U5466 ( .A1(n9377), .A2(n4446), .ZN(n9342) );
  NAND2_X1 U5467 ( .A1(n9349), .A2(n9065), .ZN(n9332) );
  NAND2_X1 U5468 ( .A1(n4574), .A2(n4572), .ZN(n9353) );
  OR2_X1 U5469 ( .A1(n4575), .A2(n4573), .ZN(n4572) );
  NOR2_X1 U5470 ( .A1(n9399), .A2(n9499), .ZN(n9377) );
  OR2_X1 U5471 ( .A1(n9583), .A2(n9506), .ZN(n9399) );
  NAND2_X1 U5472 ( .A1(n9053), .A2(n9052), .ZN(n4777) );
  NAND3_X1 U5473 ( .A1(n7484), .A2(n4266), .A3(n9600), .ZN(n9583) );
  AND2_X1 U5474 ( .A1(n7484), .A2(n4266), .ZN(n9581) );
  NAND2_X1 U5475 ( .A1(n7484), .A2(n4435), .ZN(n9629) );
  AND4_X1 U5476 ( .A1(n4866), .A2(n4865), .A3(n4864), .A4(n4863), .ZN(n9636)
         );
  NAND2_X1 U5477 ( .A1(n7086), .A2(n5569), .ZN(n7608) );
  INV_X1 U5478 ( .A(n9675), .ZN(n7098) );
  OAI21_X1 U5479 ( .B1(n6995), .B2(n5090), .A(n5561), .ZN(n7355) );
  NAND2_X1 U5480 ( .A1(n7003), .A2(n6709), .ZN(n9643) );
  AND2_X1 U5481 ( .A1(n5623), .A2(n5561), .ZN(n7000) );
  NAND2_X1 U5482 ( .A1(n4601), .A2(n5622), .ZN(n6995) );
  NAND2_X1 U5483 ( .A1(n5089), .A2(n5620), .ZN(n4601) );
  NAND2_X1 U5484 ( .A1(n4942), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n4958) );
  AND4_X2 U5485 ( .A1(n4974), .A2(n4973), .A3(n4972), .A4(n4971), .ZN(n7246)
         );
  NAND2_X1 U5486 ( .A1(n4942), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n4973) );
  INV_X1 U5487 ( .A(n9635), .ZN(n9309) );
  OR2_X1 U5488 ( .A1(n6870), .A2(n6869), .ZN(n7097) );
  NAND2_X1 U5489 ( .A1(n5423), .A2(n5422), .ZN(n9427) );
  INV_X1 U5490 ( .A(n9055), .ZN(n9600) );
  INV_X1 U5491 ( .A(n9682), .ZN(n9500) );
  NAND2_X1 U5492 ( .A1(n6253), .A2(n9654), .ZN(n6870) );
  AND2_X1 U5493 ( .A1(n6288), .A2(n6287), .ZN(n6663) );
  AND2_X1 U5494 ( .A1(n4793), .A2(n4792), .ZN(n4791) );
  INV_X1 U5495 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4792) );
  XNOR2_X1 U5496 ( .A(n5497), .B(n5500), .ZN(n8097) );
  CLKBUF_X1 U5497 ( .A(n5658), .Z(n6356) );
  XNOR2_X1 U5498 ( .A(n5466), .B(n5465), .ZN(n7968) );
  OAI21_X1 U5499 ( .B1(n5416), .B2(n4664), .A(n4661), .ZN(n5466) );
  XNOR2_X1 U5500 ( .A(n5665), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5932) );
  XNOR2_X1 U5501 ( .A(n5656), .B(n5655), .ZN(n5953) );
  NAND2_X1 U5502 ( .A1(n4691), .A2(n4695), .ZN(n5204) );
  NAND2_X1 U5503 ( .A1(n5165), .A2(n4697), .ZN(n4691) );
  INV_X1 U5504 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5065) );
  OAI21_X1 U5505 ( .B1(n5099), .B2(n5098), .A(n5097), .ZN(n5117) );
  INV_X1 U5506 ( .A(n4991), .ZN(n4780) );
  AOI21_X1 U5507 ( .B1(n4886), .B2(n4512), .A(n4300), .ZN(n4511) );
  OR2_X1 U5508 ( .A1(n4950), .A2(n9535), .ZN(n4964) );
  NAND2_X1 U5509 ( .A1(n4514), .A2(n4885), .ZN(n4948) );
  NAND2_X1 U5510 ( .A1(n4882), .A2(n4928), .ZN(n4514) );
  NOR2_X1 U5511 ( .A1(n4754), .A2(n4753), .ZN(n7710) );
  INV_X1 U5512 ( .A(n7128), .ZN(n4753) );
  INV_X1 U5513 ( .A(n7129), .ZN(n4754) );
  AND2_X1 U5514 ( .A1(n4744), .A2(n4743), .ZN(n7967) );
  NAND2_X1 U5515 ( .A1(n8067), .A2(n7910), .ZN(n7923) );
  NAND2_X1 U5516 ( .A1(n4761), .A2(n7724), .ZN(n7939) );
  NAND2_X1 U5517 ( .A1(n7728), .A2(n7727), .ZN(n8791) );
  NAND2_X1 U5518 ( .A1(n4740), .A2(n4737), .ZN(n7947) );
  NOR2_X1 U5519 ( .A1(n7851), .A2(n4741), .ZN(n4737) );
  AND3_X1 U5520 ( .A1(n4648), .A2(n4647), .A3(n4646), .ZN(n8147) );
  OR2_X1 U5521 ( .A1(n6768), .A2(n6767), .ZN(n4646) );
  OR2_X1 U5522 ( .A1(n6815), .A2(n6766), .ZN(n4648) );
  OR2_X1 U5523 ( .A1(n8111), .A2(n6765), .ZN(n4647) );
  AND4_X1 U5524 ( .A1(n7846), .A2(n7845), .A3(n7844), .A4(n7843), .ZN(n8416)
         );
  INV_X1 U5525 ( .A(n9735), .ZN(n8691) );
  INV_X1 U5526 ( .A(n8405), .ZN(n8693) );
  NAND2_X1 U5527 ( .A1(n7017), .A2(n4759), .ZN(n8020) );
  AND2_X1 U5528 ( .A1(n8021), .A2(n6918), .ZN(n4759) );
  AND2_X1 U5529 ( .A1(n7017), .A2(n6918), .ZN(n8022) );
  XNOR2_X1 U5530 ( .A(n7877), .B(n7869), .ZN(n8033) );
  NAND2_X1 U5531 ( .A1(n7958), .A2(n7807), .ZN(n8042) );
  NAND2_X1 U5532 ( .A1(n7811), .A2(n7810), .ZN(n8761) );
  INV_X1 U5533 ( .A(n8501), .ZN(n8537) );
  NAND2_X1 U5534 ( .A1(n7842), .A2(n7841), .ZN(n8751) );
  INV_X1 U5535 ( .A(n8403), .ZN(n8669) );
  NAND2_X1 U5536 ( .A1(n6903), .A2(n6744), .ZN(n6745) );
  NAND2_X1 U5537 ( .A1(n9698), .A2(n6738), .ZN(n6746) );
  NAND2_X1 U5538 ( .A1(n7782), .A2(n7781), .ZN(n8771) );
  NAND2_X1 U5539 ( .A1(n8020), .A2(n4505), .ZN(n7129) );
  AND2_X1 U5540 ( .A1(n8020), .A2(n6925), .ZN(n6932) );
  AND2_X1 U5541 ( .A1(n7893), .A2(n7892), .ZN(n8069) );
  INV_X1 U5542 ( .A(n7985), .ZN(n9704) );
  INV_X1 U5543 ( .A(n7986), .ZN(n9703) );
  NAND2_X1 U5544 ( .A1(n7746), .A2(n7745), .ZN(n8786) );
  INV_X1 U5545 ( .A(n9701), .ZN(n8083) );
  INV_X1 U5546 ( .A(n8309), .ZN(n4537) );
  NAND4_X2 U5547 ( .A1(n6467), .A2(n6466), .A3(n6465), .A4(n6464), .ZN(n8318)
         );
  INV_X2 U5548 ( .A(P2_U3966), .ZN(n8319) );
  CLKBUF_X1 U5549 ( .A(n6724), .Z(n8320) );
  NOR2_X1 U5550 ( .A1(n6561), .A2(n6562), .ZN(n6560) );
  INV_X1 U5551 ( .A(n4456), .ZN(n6604) );
  INV_X1 U5552 ( .A(n4454), .ZN(n6602) );
  INV_X1 U5553 ( .A(n4451), .ZN(n6624) );
  XNOR2_X1 U5554 ( .A(n8321), .B(n8322), .ZN(n7419) );
  NOR2_X1 U5555 ( .A1(n7419), .A2(n7418), .ZN(n8323) );
  NAND2_X1 U5556 ( .A1(n6088), .A2(n6087), .ZN(n9715) );
  NAND2_X1 U5557 ( .A1(n8384), .A2(n6510), .ZN(n9716) );
  NAND2_X1 U5558 ( .A1(n9715), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4465) );
  INV_X1 U5559 ( .A(n8390), .ZN(n4464) );
  OAI21_X1 U5560 ( .B1(n8386), .B2(n9718), .A(n4286), .ZN(n4468) );
  OAI22_X1 U5561 ( .A1(n8387), .A2(n9718), .B1(n8388), .B2(n9716), .ZN(n4466)
         );
  NAND2_X1 U5562 ( .A1(n4801), .A2(n8421), .ZN(n4800) );
  NAND2_X1 U5563 ( .A1(n4798), .A2(n4797), .ZN(n4796) );
  OAI21_X1 U5564 ( .B1(n8499), .B2(n4613), .A(n4263), .ZN(n8462) );
  NAND2_X1 U5565 ( .A1(n4618), .A2(n8272), .ZN(n4354) );
  OAI21_X1 U5566 ( .B1(n8495), .B2(n4825), .A(n4822), .ZN(n8470) );
  NAND2_X1 U5567 ( .A1(n4404), .A2(n4410), .ZN(n8572) );
  OR2_X1 U5568 ( .A1(n8621), .A2(n4411), .ZN(n4404) );
  NAND2_X1 U5569 ( .A1(n8602), .A2(n4809), .ZN(n8587) );
  NAND2_X1 U5570 ( .A1(n7766), .A2(n7765), .ZN(n8778) );
  NAND2_X1 U5571 ( .A1(n4498), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6416) );
  INV_X1 U5572 ( .A(n4622), .ZN(n8607) );
  OAI21_X1 U5573 ( .B1(n8641), .B2(n4626), .A(n8224), .ZN(n4622) );
  NAND2_X1 U5574 ( .A1(n8684), .A2(n8404), .ZN(n8671) );
  NOR2_X1 U5575 ( .A1(n9728), .A2(n4565), .ZN(n8695) );
  INV_X1 U5576 ( .A(n8613), .ZN(n9773) );
  NAND2_X1 U5577 ( .A1(n7288), .A2(n7287), .ZN(n9864) );
  AND2_X1 U5578 ( .A1(n6833), .A2(n4551), .ZN(n7181) );
  INV_X1 U5579 ( .A(n4552), .ZN(n4551) );
  OAI22_X1 U5580 ( .A1(n6831), .A2(n6815), .B1(n6768), .B2(n6834), .ZN(n4552)
         );
  OR2_X1 U5581 ( .A1(n7165), .A2(n8118), .ZN(n9754) );
  INV_X1 U5582 ( .A(n8147), .ZN(n7204) );
  NAND2_X1 U5583 ( .A1(n9779), .A2(n7162), .ZN(n8703) );
  INV_X1 U5584 ( .A(n9777), .ZN(n8698) );
  INV_X1 U5585 ( .A(n9754), .ZN(n9733) );
  INV_X1 U5586 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6212) );
  CLKBUF_X1 U5587 ( .A(n6459), .Z(n6460) );
  XNOR2_X1 U5588 ( .A(n5974), .B(n6077), .ZN(n7569) );
  XNOR2_X1 U5589 ( .A(n5965), .B(n5964), .ZN(n7354) );
  INV_X1 U5590 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U5591 ( .A1(n5963), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U5592 ( .A1(n5979), .A2(n5978), .ZN(n5963) );
  INV_X1 U5593 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7853) );
  INV_X1 U5594 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7840) );
  INV_X1 U5595 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7827) );
  INV_X1 U5596 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7809) );
  XNOR2_X1 U5597 ( .A(n6418), .B(n6417), .ZN(n6449) );
  NAND2_X1 U5598 ( .A1(n4497), .A2(n4496), .ZN(n6418) );
  AOI21_X1 U5599 ( .B1(n4499), .B2(n6071), .A(n6071), .ZN(n4496) );
  INV_X1 U5600 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6380) );
  INV_X1 U5601 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6248) );
  INV_X1 U5602 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6241) );
  INV_X1 U5603 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6074) );
  INV_X1 U5604 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6068) );
  INV_X1 U5605 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6055) );
  INV_X1 U5606 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6927) );
  INV_X1 U5607 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6832) );
  INV_X1 U5608 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6818) );
  NAND2_X1 U5609 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4458) );
  OR2_X1 U5610 ( .A1(n5954), .A2(n5980), .ZN(n6012) );
  NAND2_X1 U5611 ( .A1(n4701), .A2(n4704), .ZN(n8835) );
  AOI21_X1 U5612 ( .B1(n4287), .B2(n8923), .A(n4705), .ZN(n4704) );
  AND2_X1 U5613 ( .A1(n8924), .A2(n4707), .ZN(n4705) );
  NAND2_X1 U5614 ( .A1(n7628), .A2(n5769), .ZN(n7655) );
  AOI21_X1 U5615 ( .B1(n4977), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n4828), .ZN(
        n4931) );
  AND4_X1 U5616 ( .A1(n5080), .A2(n5079), .A3(n5078), .A4(n5077), .ZN(n9391)
         );
  NOR2_X1 U5617 ( .A1(n8903), .A2(n5893), .ZN(n8886) );
  NAND2_X1 U5618 ( .A1(n5369), .A2(n5368), .ZN(n9435) );
  AND4_X1 U5619 ( .A1(n5200), .A2(n5199), .A3(n5198), .A4(n5197), .ZN(n9336)
         );
  NOR2_X1 U5620 ( .A1(n8905), .A2(n8904), .ZN(n8903) );
  AND4_X1 U5621 ( .A1(n5033), .A2(n5032), .A3(n5031), .A4(n5030), .ZN(n9637)
         );
  NAND2_X1 U5622 ( .A1(n8873), .A2(n8874), .ZN(n4708) );
  INV_X1 U5623 ( .A(n4720), .ZN(n4719) );
  OAI21_X1 U5624 ( .B1(n4724), .B2(n4721), .A(n8866), .ZN(n4720) );
  AOI21_X1 U5625 ( .B1(n4711), .B2(n7630), .A(n4309), .ZN(n4710) );
  INV_X1 U5626 ( .A(n8991), .ZN(n8970) );
  INV_X1 U5627 ( .A(n8977), .ZN(n8989) );
  INV_X1 U5628 ( .A(n9143), .ZN(n9178) );
  INV_X1 U5629 ( .A(n9158), .ZN(n9193) );
  OR2_X1 U5630 ( .A1(n5357), .A2(n5356), .ZN(n9235) );
  INV_X1 U5631 ( .A(n9391), .ZN(n9056) );
  INV_X1 U5632 ( .A(n9637), .ZN(n8997) );
  CLKBUF_X1 U5633 ( .A(n5689), .Z(n9005) );
  NAND2_X1 U5634 ( .A1(n4942), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n4938) );
  CLKBUF_X2 U5635 ( .A(P1_U4006), .Z(n9004) );
  OR2_X1 U5636 ( .A1(n6010), .A2(n5982), .ZN(n6264) );
  NAND2_X1 U5637 ( .A1(n6279), .A2(n6280), .ZN(n6278) );
  NOR2_X1 U5638 ( .A1(n6690), .A2(n4282), .ZN(n6330) );
  NAND2_X1 U5639 ( .A1(n6330), .A2(n6331), .ZN(n6329) );
  INV_X1 U5640 ( .A(n4398), .ZN(n6403) );
  INV_X1 U5641 ( .A(n9030), .ZN(n9623) );
  XNOR2_X1 U5642 ( .A(n7270), .B(n7269), .ZN(n6956) );
  NOR2_X1 U5643 ( .A1(n6956), .A2(n6955), .ZN(n7271) );
  NAND2_X1 U5644 ( .A1(n5477), .A2(n5476), .ZN(n9410) );
  INV_X1 U5645 ( .A(n9417), .ZN(n9129) );
  AND2_X1 U5646 ( .A1(n5447), .A2(n5425), .ZN(n9162) );
  AND2_X1 U5647 ( .A1(n5397), .A2(n5396), .ZN(n9172) );
  INV_X1 U5648 ( .A(n9080), .ZN(n9442) );
  AND2_X1 U5649 ( .A1(n5347), .A2(n5346), .ZN(n9225) );
  INV_X1 U5650 ( .A(n4580), .ZN(n9260) );
  AOI21_X1 U5651 ( .B1(n4592), .B2(n4582), .A(n4581), .ZN(n4580) );
  NAND2_X1 U5652 ( .A1(n4769), .A2(n4770), .ZN(n9258) );
  NAND2_X1 U5653 ( .A1(n9285), .A2(n4773), .ZN(n4769) );
  NAND2_X1 U5654 ( .A1(n4592), .A2(n4590), .ZN(n9271) );
  AOI21_X1 U5655 ( .B1(n9285), .B2(n9286), .A(n4277), .ZN(n9270) );
  CLKBUF_X1 U5656 ( .A(n9321), .Z(n9322) );
  NAND2_X1 U5657 ( .A1(n9063), .A2(n9062), .ZN(n9351) );
  NAND2_X1 U5658 ( .A1(n4577), .A2(n4575), .ZN(n9372) );
  CLKBUF_X1 U5659 ( .A(n7605), .Z(n7477) );
  NAND2_X1 U5660 ( .A1(n7476), .A2(n7475), .ZN(n7479) );
  NAND2_X1 U5661 ( .A1(n7091), .A2(n7090), .ZN(n7358) );
  OR2_X1 U5662 ( .A1(n9510), .A2(n5949), .ZN(n9245) );
  INV_X1 U5663 ( .A(n9584), .ZN(n9631) );
  NAND2_X1 U5664 ( .A1(n7097), .A2(n9245), .ZN(n9650) );
  AND2_X1 U5665 ( .A1(n4437), .A2(n4320), .ZN(n9418) );
  OR2_X1 U5666 ( .A1(n9415), .A2(n9682), .ZN(n4437) );
  NAND2_X1 U5667 ( .A1(n9424), .A2(n4353), .ZN(n9514) );
  NOR2_X1 U5668 ( .A1(n9421), .A2(n4268), .ZN(n4353) );
  INV_X1 U5669 ( .A(n9659), .ZN(n9660) );
  XNOR2_X1 U5670 ( .A(n5494), .B(n5493), .ZN(n9534) );
  NAND2_X1 U5671 ( .A1(n4674), .A2(n4672), .ZN(n5494) );
  INV_X1 U5672 ( .A(n5661), .ZN(n5662) );
  INV_X1 U5673 ( .A(n5932), .ZN(n7352) );
  INV_X1 U5674 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7057) );
  INV_X1 U5675 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7706) );
  OR2_X1 U5676 ( .A1(n5517), .A2(n5068), .ZN(n5518) );
  OAI21_X1 U5677 ( .B1(n5071), .B2(n4734), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5517) );
  INV_X1 U5678 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6758) );
  INV_X1 U5679 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6381) );
  AND2_X1 U5680 ( .A1(n5213), .A2(n5230), .ZN(n9015) );
  INV_X1 U5681 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6230) );
  INV_X1 U5682 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6075) );
  INV_X1 U5683 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U5684 ( .A1(n4680), .A2(n4685), .ZN(n5140) );
  NAND2_X1 U5685 ( .A1(n5099), .A2(n4687), .ZN(n4680) );
  INV_X1 U5686 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6064) );
  INV_X1 U5687 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6062) );
  INV_X1 U5688 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6186) );
  INV_X1 U5689 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U5690 ( .A1(n4382), .A2(n4900), .ZN(n4381) );
  NAND2_X1 U5691 ( .A1(n4990), .A2(n4989), .ZN(n4382) );
  NOR2_X1 U5692 ( .A1(n7410), .A2(n9950), .ZN(n9941) );
  AOI21_X1 U5693 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9939), .ZN(n9938) );
  NOR2_X1 U5694 ( .A1(n9938), .A2(n9937), .ZN(n9936) );
  AOI21_X1 U5695 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9936), .ZN(n9935) );
  OAI21_X1 U5696 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9933), .ZN(n9931) );
  NAND2_X1 U5697 ( .A1(n4490), .A2(n4493), .ZN(n4487) );
  NAND2_X1 U5698 ( .A1(n7708), .A2(n7140), .ZN(n7147) );
  NAND2_X1 U5699 ( .A1(n7012), .A2(n6911), .ZN(n7019) );
  NAND2_X1 U5700 ( .A1(n4536), .A2(n8308), .ZN(P2_U3244) );
  OAI21_X1 U5701 ( .B1(n4538), .B2(n4299), .A(n4537), .ZN(n4536) );
  NAND2_X1 U5702 ( .A1(n4467), .A2(n4462), .ZN(P2_U3264) );
  AOI21_X1 U5703 ( .B1(n4466), .B2(n8389), .A(n4463), .ZN(n4462) );
  NAND2_X1 U5704 ( .A1(n4468), .A2(n6456), .ZN(n4467) );
  NAND2_X1 U5705 ( .A1(n4465), .A2(n4464), .ZN(n4463) );
  NAND2_X1 U5706 ( .A1(n4260), .A2(n9894), .ZN(n4421) );
  INV_X1 U5707 ( .A(n4416), .ZN(n4415) );
  OAI21_X1 U5708 ( .B1(n4424), .B2(n9910), .A(n4422), .ZN(n4416) );
  NAND2_X1 U5709 ( .A1(n4379), .A2(n4378), .ZN(P1_U3240) );
  NAND2_X1 U5710 ( .A1(n4666), .A2(n4377), .ZN(n4378) );
  INV_X1 U5711 ( .A(n5669), .ZN(n4380) );
  INV_X1 U5712 ( .A(n4395), .ZN(n4394) );
  XNOR2_X1 U5713 ( .A(n6086), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6421) );
  INV_X4 U5714 ( .A(n5050), .ZN(n4977) );
  AND2_X1 U5715 ( .A1(n8781), .A2(n8411), .ZN(n8412) );
  OR2_X1 U5716 ( .A1(n6679), .A2(n6729), .ZN(n6739) );
  OR2_X1 U5717 ( .A1(n8732), .A2(n8274), .ZN(n8273) );
  XNOR2_X1 U5718 ( .A(n6084), .B(n6083), .ZN(n6470) );
  OAI21_X1 U5719 ( .B1(n4808), .B2(n4807), .A(n4279), .ZN(n4806) );
  AND2_X1 U5720 ( .A1(n4616), .A2(n4611), .ZN(n4263) );
  AND2_X1 U5721 ( .A1(n8460), .A2(n8440), .ZN(n4264) );
  AND2_X1 U5722 ( .A1(n4446), .A2(n4445), .ZN(n4265) );
  AND2_X1 U5723 ( .A1(n4435), .A2(n9570), .ZN(n4266) );
  NAND2_X1 U5724 ( .A1(n6217), .A2(n6216), .ZN(n6219) );
  NAND3_X1 U5725 ( .A1(n4880), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4532) );
  INV_X1 U5726 ( .A(n4532), .ZN(n4373) );
  OR2_X1 U5727 ( .A1(n8277), .A2(n8280), .ZN(n4267) );
  OR2_X1 U5728 ( .A1(n9422), .A2(n4331), .ZN(n4268) );
  AND2_X1 U5729 ( .A1(n4479), .A2(n7990), .ZN(n4269) );
  AND3_X1 U5730 ( .A1(n4781), .A2(n4840), .A3(n4842), .ZN(n4270) );
  NAND2_X1 U5731 ( .A1(n4780), .A2(n4782), .ZN(n5037) );
  OR2_X1 U5732 ( .A1(n8527), .A2(n4556), .ZN(n4271) );
  NAND3_X1 U5733 ( .A1(n4841), .A2(n4782), .A3(n4270), .ZN(n4875) );
  INV_X1 U5734 ( .A(n7512), .ZN(n7337) );
  AND2_X1 U5735 ( .A1(n8190), .A2(n8191), .ZN(n7512) );
  INV_X1 U5736 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4870) );
  NAND2_X1 U5737 ( .A1(n4652), .A2(n4342), .ZN(n9046) );
  INV_X1 U5738 ( .A(n9046), .ZN(n4651) );
  AOI21_X1 U5739 ( .B1(n4740), .B2(n4742), .A(n7864), .ZN(n7946) );
  NAND2_X1 U5740 ( .A1(n4834), .A2(n4809), .ZN(n4272) );
  INV_X1 U5741 ( .A(n8418), .ZN(n4823) );
  NAND2_X1 U5742 ( .A1(n9287), .A2(n4442), .ZN(n4443) );
  INV_X1 U5743 ( .A(n8643), .ZN(n4628) );
  INV_X1 U5744 ( .A(n8115), .ZN(n4638) );
  XOR2_X1 U5745 ( .A(n6032), .B(n5989), .Z(n4273) );
  INV_X1 U5746 ( .A(n5355), .ZN(n4954) );
  INV_X1 U5747 ( .A(n6462), .ZN(n7931) );
  AND2_X1 U5748 ( .A1(n6224), .A2(n6218), .ZN(n7916) );
  OR2_X1 U5749 ( .A1(n9728), .A2(n4563), .ZN(n4274) );
  AND2_X1 U5750 ( .A1(n8286), .A2(n8285), .ZN(n8421) );
  OR2_X1 U5751 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4275) );
  INV_X1 U5752 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5655) );
  INV_X1 U5753 ( .A(n4825), .ZN(n4824) );
  NAND2_X1 U5754 ( .A1(n4615), .A2(n4826), .ZN(n4825) );
  AND2_X1 U5755 ( .A1(n6913), .A2(n6911), .ZN(n4276) );
  NAND2_X1 U5756 ( .A1(n4278), .A2(n5960), .ZN(n4812) );
  OR2_X1 U5757 ( .A1(n8737), .A2(n8094), .ZN(n8272) );
  AND2_X1 U5758 ( .A1(n9471), .A2(n9310), .ZN(n4277) );
  AND2_X1 U5759 ( .A1(n5959), .A2(n4814), .ZN(n4278) );
  NOR2_X1 U5760 ( .A1(n4991), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n4993) );
  NAND2_X1 U5761 ( .A1(n8771), .A2(n8580), .ZN(n4279) );
  OR2_X1 U5762 ( .A1(n8740), .A2(n8511), .ZN(n8418) );
  XNOR2_X1 U5763 ( .A(n4458), .B(n6029), .ZN(n6571) );
  NOR2_X1 U5764 ( .A1(n8966), .A2(n8967), .ZN(n4280) );
  OR2_X1 U5765 ( .A1(n4433), .A2(n4875), .ZN(n4281) );
  NOR2_X1 U5766 ( .A1(n8494), .A2(n4823), .ZN(n8482) );
  INV_X1 U5767 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5957) );
  AND2_X1 U5768 ( .A1(n6695), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4282) );
  NAND2_X1 U5769 ( .A1(n6470), .A2(n6877), .ZN(n6729) );
  INV_X1 U5770 ( .A(n9259), .ZN(n4586) );
  NOR2_X1 U5771 ( .A1(n8912), .A2(n5865), .ZN(n4283) );
  AND2_X1 U5772 ( .A1(n8091), .A2(n4625), .ZN(n4284) );
  AND3_X1 U5773 ( .A1(n6072), .A2(n6231), .A3(n5961), .ZN(n4285) );
  INV_X1 U5774 ( .A(n9097), .ZN(n4573) );
  NAND2_X1 U5775 ( .A1(n7718), .A2(n7717), .ZN(n8725) );
  AND2_X1 U5776 ( .A1(n8385), .A2(n9717), .ZN(n4286) );
  INV_X1 U5777 ( .A(n9067), .ZN(n4786) );
  OR2_X1 U5778 ( .A1(n8924), .A2(n4707), .ZN(n4287) );
  NAND2_X1 U5779 ( .A1(n5313), .A2(n5312), .ZN(n9450) );
  INV_X1 U5780 ( .A(n9450), .ZN(n4439) );
  XNOR2_X1 U5781 ( .A(n8725), .B(n8440), .ZN(n8461) );
  INV_X1 U5782 ( .A(n5558), .ZN(n4371) );
  INV_X1 U5783 ( .A(n8875), .ZN(n4707) );
  AND2_X1 U5784 ( .A1(n4454), .A2(n4453), .ZN(n4288) );
  NOR2_X1 U5785 ( .A1(n9307), .A2(n9103), .ZN(n4289) );
  AND2_X1 U5786 ( .A1(n9463), .A2(n9073), .ZN(n4290) );
  AND2_X1 U5787 ( .A1(n4787), .A2(n9067), .ZN(n4291) );
  NAND2_X1 U5788 ( .A1(n8273), .A2(n8095), .ZN(n8471) );
  AND2_X1 U5789 ( .A1(n8667), .A2(n8404), .ZN(n4292) );
  INV_X1 U5790 ( .A(n4813), .ZN(n6044) );
  AND2_X1 U5791 ( .A1(n9758), .A2(n7334), .ZN(n4293) );
  NAND2_X1 U5792 ( .A1(n7868), .A2(n7867), .ZN(n8740) );
  NAND2_X1 U5793 ( .A1(n6019), .A2(n5957), .ZN(n6024) );
  AND2_X1 U5794 ( .A1(n4609), .A2(n8455), .ZN(n4294) );
  NAND2_X1 U5795 ( .A1(n5176), .A2(n5175), .ZN(n9487) );
  NAND2_X1 U5796 ( .A1(n8996), .A2(n9681), .ZN(n4295) );
  NAND2_X1 U5797 ( .A1(n5292), .A2(n5291), .ZN(n9458) );
  NAND2_X1 U5798 ( .A1(n8421), .A2(n8279), .ZN(n4296) );
  INV_X1 U5799 ( .A(n7140), .ZN(n4752) );
  AND2_X1 U5800 ( .A1(n4642), .A2(n7512), .ZN(n4297) );
  NAND2_X1 U5801 ( .A1(n8705), .A2(n8115), .ZN(n4298) );
  NOR2_X1 U5802 ( .A1(n8527), .A2(n4557), .ZN(n4555) );
  NAND2_X1 U5803 ( .A1(n5444), .A2(n5443), .ZN(n9423) );
  AND2_X1 U5804 ( .A1(n4541), .A2(n8300), .ZN(n4299) );
  AND2_X1 U5805 ( .A1(n4887), .A2(SI_2_), .ZN(n4300) );
  AND2_X1 U5806 ( .A1(n8217), .A2(n8653), .ZN(n4301) );
  AND2_X1 U5807 ( .A1(n9387), .A2(n9385), .ZN(n9579) );
  AND2_X1 U5808 ( .A1(n4548), .A2(n8270), .ZN(n4302) );
  AND2_X1 U5809 ( .A1(n5548), .A2(n9118), .ZN(n9139) );
  INV_X1 U5810 ( .A(n8391), .ZN(n8714) );
  OR2_X1 U5811 ( .A1(n9066), .A2(n4786), .ZN(n9334) );
  INV_X1 U5812 ( .A(n9334), .ZN(n4367) );
  INV_X1 U5813 ( .A(n4804), .ZN(n4803) );
  NAND2_X1 U5814 ( .A1(n8450), .A2(n4805), .ZN(n4804) );
  NAND2_X1 U5815 ( .A1(n8269), .A2(n8273), .ZN(n4303) );
  OR2_X1 U5816 ( .A1(n4741), .A2(n7949), .ZN(n4304) );
  OR3_X1 U5817 ( .A1(n4875), .A2(n4789), .A3(P1_IR_REG_23__SCAN_IN), .ZN(n4305) );
  NOR2_X1 U5818 ( .A1(n8737), .A2(n8502), .ZN(n4306) );
  NAND2_X1 U5819 ( .A1(n7838), .A2(n7837), .ZN(n4307) );
  AND2_X1 U5820 ( .A1(n8272), .A2(n8260), .ZN(n8483) );
  INV_X1 U5821 ( .A(n8483), .ZN(n4615) );
  AND2_X1 U5822 ( .A1(n8448), .A2(n8420), .ZN(n4308) );
  INV_X1 U5823 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4874) );
  INV_X1 U5824 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n4842) );
  NAND2_X1 U5825 ( .A1(n4841), .A2(n4840), .ZN(n4991) );
  AND2_X1 U5826 ( .A1(n5774), .A2(n7652), .ZN(n4309) );
  AND2_X1 U5827 ( .A1(n7922), .A2(n8068), .ZN(n4310) );
  OR2_X1 U5828 ( .A1(n4549), .A2(n4550), .ZN(n4311) );
  AND2_X1 U5829 ( .A1(n4902), .A2(SI_6_), .ZN(n4312) );
  OAI21_X1 U5830 ( .B1(n4480), .B2(n4478), .A(n4307), .ZN(n4477) );
  NOR2_X1 U5831 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n4313) );
  OR2_X1 U5832 ( .A1(n6443), .A2(n6445), .ZN(n4314) );
  OR2_X1 U5833 ( .A1(n4272), .A2(n4412), .ZN(n4315) );
  INV_X1 U5834 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4375) );
  INV_X1 U5835 ( .A(n4834), .ZN(n4808) );
  NAND2_X1 U5836 ( .A1(n8279), .A2(n8096), .ZN(n8450) );
  OR2_X1 U5837 ( .A1(n8885), .A2(n4727), .ZN(n4316) );
  NAND2_X1 U5838 ( .A1(n5755), .A2(n5754), .ZN(n4317) );
  AND2_X1 U5839 ( .A1(n9095), .A2(n9097), .ZN(n4318) );
  AND2_X1 U5840 ( .A1(n4440), .A2(n4439), .ZN(n4319) );
  NOR2_X1 U5841 ( .A1(n9416), .A2(n4436), .ZN(n4320) );
  INV_X1 U5842 ( .A(n8745), .ZN(n8517) );
  NAND2_X1 U5843 ( .A1(n7855), .A2(n7854), .ZN(n8745) );
  INV_X1 U5844 ( .A(n8720), .ZN(n8448) );
  OR2_X1 U5845 ( .A1(n8576), .A2(n8413), .ZN(n4321) );
  AND2_X1 U5846 ( .A1(n8218), .A2(n8219), .ZN(n8653) );
  AND2_X1 U5847 ( .A1(n4774), .A2(n4773), .ZN(n4322) );
  NAND2_X1 U5848 ( .A1(n7653), .A2(n5773), .ZN(n4323) );
  INV_X1 U5849 ( .A(n9074), .ZN(n4774) );
  NOR2_X1 U5850 ( .A1(n9463), .A2(n9073), .ZN(n9074) );
  AND2_X1 U5851 ( .A1(n7092), .A2(n7090), .ZN(n4324) );
  AND2_X1 U5852 ( .A1(n4803), .A2(n8422), .ZN(n4325) );
  NAND2_X1 U5853 ( .A1(n5659), .A2(n4851), .ZN(n4326) );
  AND2_X1 U5854 ( .A1(n4505), .A2(n7140), .ZN(n4327) );
  AND2_X1 U5855 ( .A1(n4692), .A2(n5203), .ZN(n4328) );
  AND2_X1 U5856 ( .A1(n4280), .A2(n5892), .ZN(n4329) );
  AND2_X1 U5857 ( .A1(n4285), .A2(n4501), .ZN(n4330) );
  INV_X1 U5858 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5063) );
  AND2_X1 U5859 ( .A1(n4820), .A2(n6077), .ZN(n4819) );
  INV_X1 U5860 ( .A(n4812), .ZN(n4811) );
  AND2_X1 U5861 ( .A1(n4323), .A2(n5769), .ZN(n4711) );
  INV_X1 U5862 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n4535) );
  NAND2_X1 U5863 ( .A1(n6452), .A2(n8170), .ZN(n6447) );
  AND3_X1 U5864 ( .A1(n4841), .A2(n4598), .A3(n4782), .ZN(n5051) );
  INV_X1 U5865 ( .A(n7619), .ZN(n9570) );
  NAND2_X1 U5866 ( .A1(n4469), .A2(n4472), .ZN(n8006) );
  INV_X1 U5867 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4376) );
  OAI21_X1 U5868 ( .B1(n4758), .B2(n4482), .A(n4480), .ZN(n7989) );
  NAND2_X1 U5869 ( .A1(n7576), .A2(n7575), .ZN(n7720) );
  NAND2_X1 U5870 ( .A1(n4708), .A2(n8875), .ZN(n8922) );
  INV_X1 U5871 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4814) );
  NAND2_X1 U5872 ( .A1(n5192), .A2(n5191), .ZN(n9483) );
  INV_X1 U5873 ( .A(n9483), .ZN(n4445) );
  AND2_X1 U5874 ( .A1(n9423), .A2(n9568), .ZN(n4331) );
  AND2_X1 U5875 ( .A1(n5051), .A2(n4728), .ZN(n5170) );
  NAND2_X1 U5876 ( .A1(n4813), .A2(n4811), .ZN(n6065) );
  NAND2_X1 U5877 ( .A1(n4758), .A2(n7792), .ZN(n7957) );
  NAND2_X1 U5878 ( .A1(n7829), .A2(n7828), .ZN(n8756) );
  NAND2_X1 U5879 ( .A1(n4777), .A2(n9054), .ZN(n9578) );
  NAND2_X1 U5880 ( .A1(n4813), .A2(n4278), .ZN(n6047) );
  OR2_X1 U5881 ( .A1(n8517), .A2(n8537), .ZN(n4332) );
  AND2_X1 U5882 ( .A1(n4761), .A2(n4760), .ZN(n4333) );
  INV_X1 U5883 ( .A(n8412), .ZN(n4414) );
  NAND2_X1 U5884 ( .A1(n5215), .A2(n5214), .ZN(n9476) );
  INV_X1 U5885 ( .A(n4626), .ZN(n4625) );
  NAND2_X1 U5886 ( .A1(n4627), .A2(n8225), .ZN(n4626) );
  INV_X1 U5887 ( .A(n7607), .ZN(n4571) );
  AND2_X1 U5888 ( .A1(n5051), .A2(n4730), .ZN(n4334) );
  AND2_X1 U5889 ( .A1(n4502), .A2(n4813), .ZN(n4335) );
  OR2_X1 U5890 ( .A1(n6476), .A2(n7153), .ZN(n9910) );
  AND2_X1 U5891 ( .A1(n7484), .A2(n7557), .ZN(n4336) );
  NAND2_X1 U5892 ( .A1(n6299), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6379) );
  INV_X2 U5893 ( .A(n6905), .ZN(n8118) );
  INV_X1 U5894 ( .A(n6739), .ZN(n6905) );
  OR3_X1 U5895 ( .A1(n9728), .A2(n8697), .A3(n4565), .ZN(n4337) );
  NAND2_X1 U5896 ( .A1(n9747), .A2(n7335), .ZN(n7338) );
  NAND2_X1 U5897 ( .A1(n4815), .A2(n4293), .ZN(n9747) );
  NAND2_X1 U5898 ( .A1(n4815), .A2(n7334), .ZN(n9748) );
  OR2_X1 U5899 ( .A1(n5975), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4338) );
  INV_X1 U5900 ( .A(n4560), .ZN(n7185) );
  OR2_X1 U5901 ( .A1(n4875), .A2(n4789), .ZN(n4339) );
  AND2_X1 U5902 ( .A1(n7987), .A2(n7988), .ZN(n4340) );
  NAND2_X1 U5903 ( .A1(n6741), .A2(n6740), .ZN(n6903) );
  NAND2_X1 U5904 ( .A1(n5678), .A2(n9207), .ZN(n5947) );
  NAND2_X1 U5905 ( .A1(n6760), .A2(n8160), .ZN(n7236) );
  INV_X1 U5906 ( .A(n7236), .ZN(n4554) );
  OR2_X1 U5907 ( .A1(n6445), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n4341) );
  INV_X1 U5908 ( .A(n6421), .ZN(n6877) );
  AND2_X1 U5909 ( .A1(n4949), .A2(n4341), .ZN(n4342) );
  INV_X1 U5910 ( .A(n7286), .ZN(n4449) );
  INV_X1 U5911 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n4448) );
  XNOR2_X1 U5912 ( .A(n6416), .B(P2_IR_REG_19__SCAN_IN), .ZN(n6456) );
  NAND2_X1 U5913 ( .A1(n6278), .A2(n5988), .ZN(n4343) );
  INV_X1 U5914 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n4386) );
  INV_X1 U5915 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4534) );
  OR2_X1 U5916 ( .A1(n8177), .A2(n8295), .ZN(n4508) );
  NAND3_X2 U5917 ( .A1(n6470), .A2(n6456), .A3(n6421), .ZN(n8295) );
  AND2_X1 U5918 ( .A1(n4344), .A2(n6891), .ZN(n8943) );
  NAND2_X1 U5919 ( .A1(n5704), .A2(n5705), .ZN(n4344) );
  NAND2_X1 U5920 ( .A1(n7430), .A2(n5757), .ZN(n7554) );
  INV_X1 U5921 ( .A(n8892), .ZN(n4347) );
  OAI21_X1 U5922 ( .B1(n8858), .B2(n8855), .A(n8854), .ZN(n8914) );
  NOR2_X1 U5923 ( .A1(n4345), .A2(n4326), .ZN(n4431) );
  NAND2_X2 U5924 ( .A1(n5841), .A2(n8893), .ZN(n8953) );
  INV_X1 U5925 ( .A(n4844), .ZN(n4790) );
  NAND2_X1 U5926 ( .A1(n7431), .A2(n7432), .ZN(n7430) );
  INV_X1 U5927 ( .A(n4434), .ZN(n4873) );
  NAND2_X1 U5928 ( .A1(n5688), .A2(n5687), .ZN(n6370) );
  NAND2_X1 U5929 ( .A1(n6895), .A2(n5719), .ZN(n7029) );
  NOR2_X1 U5930 ( .A1(n5836), .A2(n5835), .ZN(n5847) );
  OAI21_X2 U5931 ( .B1(n5071), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5606) );
  NOR2_X2 U5932 ( .A1(n5670), .A2(n4699), .ZN(n5699) );
  NAND2_X1 U5933 ( .A1(n5718), .A2(n6892), .ZN(n6895) );
  NOR2_X2 U5934 ( .A1(n4849), .A2(n4848), .ZN(n4850) );
  NAND2_X1 U5935 ( .A1(n7332), .A2(n7331), .ZN(n4815) );
  OR2_X2 U5936 ( .A1(n4802), .A2(n8450), .ZN(n4418) );
  NAND2_X1 U5937 ( .A1(n9727), .A2(n7510), .ZN(n7511) );
  NAND2_X1 U5938 ( .A1(n4403), .A2(n4821), .ZN(n4402) );
  NAND2_X1 U5939 ( .A1(n8673), .A2(n8406), .ZN(n8652) );
  NAND2_X2 U5940 ( .A1(n8650), .A2(n8408), .ZN(n8634) );
  NAND2_X1 U5941 ( .A1(n4813), .A2(n4644), .ZN(n5975) );
  NOR2_X2 U5942 ( .A1(n4351), .A2(n5972), .ZN(n5973) );
  NAND4_X1 U5943 ( .A1(n5966), .A2(n5968), .A3(n5967), .A4(n5969), .ZN(n4351)
         );
  NAND2_X1 U5944 ( .A1(n4407), .A2(n4405), .ZN(n8555) );
  OAI21_X1 U5945 ( .B1(n7212), .B2(n9844), .A(n8179), .ZN(n4401) );
  NAND2_X1 U5946 ( .A1(n9252), .A2(n9251), .ZN(n9253) );
  NAND2_X1 U5947 ( .A1(n7356), .A2(n7093), .ZN(n7095) );
  NAND2_X1 U5948 ( .A1(n5331), .A2(n5330), .ZN(n5360) );
  NAND2_X1 U5949 ( .A1(n5290), .A2(n5289), .ZN(n5307) );
  NAND2_X1 U5950 ( .A1(n4919), .A2(n4918), .ZN(n5081) );
  NAND2_X1 U5951 ( .A1(n4614), .A2(n4612), .ZN(n4611) );
  NAND2_X1 U5952 ( .A1(n5248), .A2(n5247), .ZN(n4689) );
  NAND2_X1 U5953 ( .A1(n5142), .A2(n5141), .ZN(n5165) );
  OAI21_X1 U5954 ( .B1(n5324), .B2(n5323), .A(n5325), .ZN(n5345) );
  OAI21_X1 U5955 ( .B1(n8724), .B2(n8796), .A(n4424), .ZN(n8805) );
  INV_X1 U5956 ( .A(n8723), .ZN(n4426) );
  NAND2_X1 U5957 ( .A1(n5206), .A2(n5205), .ZN(n5223) );
  NAND2_X1 U5958 ( .A1(n7255), .A2(n8145), .ZN(n7188) );
  NAND2_X1 U5959 ( .A1(n4603), .A2(n4605), .ZN(n7255) );
  AOI211_X2 U5960 ( .C1(n9835), .C2(n8732), .A(n8731), .B(n8730), .ZN(n8733)
         );
  AOI21_X2 U5961 ( .B1(n7218), .B2(n8130), .A(n8156), .ZN(n7219) );
  AND4_X4 U5962 ( .A1(n4817), .A2(n6019), .A3(n5958), .A4(n5957), .ZN(n4813)
         );
  NAND2_X1 U5963 ( .A1(n8484), .A2(n8483), .ZN(n4618) );
  NOR2_X1 U5964 ( .A1(n8657), .A2(n8089), .ZN(n8642) );
  NAND2_X1 U5965 ( .A1(n6838), .A2(n8165), .ZN(n4605) );
  NAND2_X1 U5966 ( .A1(n6214), .A2(n6212), .ZN(n6216) );
  INV_X1 U5967 ( .A(n5973), .ZN(n4645) );
  NAND2_X2 U5968 ( .A1(n7219), .A2(n8181), .ZN(n7340) );
  NAND2_X2 U5969 ( .A1(n8509), .A2(n8253), .ZN(n8499) );
  NAND2_X1 U5970 ( .A1(n4722), .A2(n4719), .ZN(n8934) );
  NAND2_X1 U5971 ( .A1(n4850), .A2(n4790), .ZN(n4789) );
  NAND3_X1 U5972 ( .A1(n4533), .A2(P1_DATAO_REG_2__SCAN_IN), .A3(n4532), .ZN(
        n4374) );
  AOI21_X1 U5973 ( .B1(n5609), .B2(n5657), .A(n4380), .ZN(n4379) );
  NAND2_X1 U5974 ( .A1(n6278), .A2(n4388), .ZN(n6359) );
  NAND3_X1 U5975 ( .A1(n4396), .A2(n4394), .A3(n4390), .ZN(P1_U3260) );
  NAND2_X1 U5976 ( .A1(n4391), .A2(n9250), .ZN(n4390) );
  NAND2_X1 U5977 ( .A1(n9035), .A2(n9616), .ZN(n4393) );
  XNOR2_X1 U5978 ( .A(n9024), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9035) );
  OAI21_X1 U5979 ( .B1(n9039), .B2(n9040), .A(n9038), .ZN(n4395) );
  OR2_X1 U5980 ( .A1(n9036), .A2(n9250), .ZN(n4396) );
  OR2_X2 U5981 ( .A1(n8652), .A2(n8653), .ZN(n8650) );
  NAND2_X1 U5982 ( .A1(n7213), .A2(n4401), .ZN(n7332) );
  NAND2_X1 U5983 ( .A1(n7184), .A2(n7183), .ZN(n7212) );
  NAND2_X2 U5984 ( .A1(n4402), .A2(n8419), .ZN(n8454) );
  NAND2_X1 U5985 ( .A1(n8621), .A2(n4408), .ZN(n4407) );
  NAND3_X1 U5986 ( .A1(n4410), .A2(n4411), .A3(n4409), .ZN(n4406) );
  NAND2_X1 U5987 ( .A1(n4802), .A2(n4420), .ZN(n4417) );
  OAI21_X1 U5988 ( .B1(n8724), .B2(n4421), .A(n4415), .ZN(P2_U3548) );
  NAND3_X1 U5989 ( .A1(n4418), .A2(n4417), .A3(n4419), .ZN(n8724) );
  OR2_X1 U5990 ( .A1(n4260), .A2(n4423), .ZN(n4422) );
  NAND2_X4 U5991 ( .A1(n6459), .A2(n8828), .ZN(n6768) );
  XNOR2_X2 U5992 ( .A(n4428), .B(n6078), .ZN(n6459) );
  NOR2_X2 U5993 ( .A1(n4783), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n4782) );
  INV_X1 U5994 ( .A(n4875), .ZN(n4432) );
  NAND3_X1 U5995 ( .A1(n4432), .A2(n4431), .A3(n4850), .ZN(n4434) );
  INV_X1 U5996 ( .A(n4443), .ZN(n9240) );
  MUX2_X1 U5997 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6479), .S(n6571), .Z(n6561)
         );
  NAND4_X1 U5998 ( .A1(n9698), .A2(n6738), .A3(n6744), .A4(n6903), .ZN(n6904)
         );
  NAND2_X1 U5999 ( .A1(n7576), .A2(n4470), .ZN(n4469) );
  NAND2_X1 U6000 ( .A1(n4744), .A2(n4485), .ZN(n4484) );
  OAI211_X1 U6001 ( .C1(n4744), .C2(n4487), .A(n4484), .B(n4340), .ZN(P2_U3222) );
  NAND2_X1 U6002 ( .A1(n6379), .A2(n4499), .ZN(n4497) );
  NAND2_X1 U6003 ( .A1(n6379), .A2(n6378), .ZN(n4498) );
  NAND3_X1 U6004 ( .A1(n4502), .A2(n4813), .A3(n4285), .ZN(n6238) );
  NAND2_X1 U6005 ( .A1(n8020), .A2(n4327), .ZN(n4504) );
  NAND2_X1 U6006 ( .A1(n4504), .A2(n4750), .ZN(n7297) );
  NAND2_X1 U6007 ( .A1(n7297), .A2(n7296), .ZN(n7310) );
  NAND3_X1 U6008 ( .A1(n4510), .A2(n8175), .A3(n8176), .ZN(n4509) );
  INV_X1 U6009 ( .A(n4885), .ZN(n4512) );
  NAND2_X1 U6010 ( .A1(n4513), .A2(n4511), .ZN(n4961) );
  NAND3_X1 U6011 ( .A1(n4882), .A2(n4928), .A3(n4886), .ZN(n4513) );
  NAND4_X1 U6012 ( .A1(n4530), .A2(n4529), .A3(SI_0_), .A4(n4528), .ZN(n4883)
         );
  NAND3_X1 U6013 ( .A1(n4533), .A2(n4532), .A3(n4535), .ZN(n4529) );
  NAND2_X1 U6014 ( .A1(n8262), .A2(n4546), .ZN(n4544) );
  NAND2_X1 U6015 ( .A1(n8271), .A2(n4548), .ZN(n4543) );
  NAND3_X1 U6016 ( .A1(n4544), .A2(n4543), .A3(n4542), .ZN(n8278) );
  NOR2_X1 U6017 ( .A1(n4545), .A2(n4302), .ZN(n4542) );
  NAND2_X1 U6018 ( .A1(n8455), .A2(n8275), .ZN(n4549) );
  NAND3_X1 U6019 ( .A1(n4811), .A2(n4813), .A3(n4553), .ZN(n4643) );
  AND2_X2 U6020 ( .A1(n5955), .A2(n5956), .ZN(n6019) );
  MUX2_X1 U6021 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8831), .S(n6768), .Z(n9821) );
  INV_X1 U6022 ( .A(n4555), .ZN(n8487) );
  NOR2_X1 U6023 ( .A1(n8474), .A2(n8725), .ZN(n8456) );
  NAND2_X1 U6024 ( .A1(n4567), .A2(n4569), .ZN(n9634) );
  INV_X1 U6025 ( .A(n4568), .ZN(n4567) );
  NAND2_X1 U6026 ( .A1(n9588), .A2(n4318), .ZN(n4574) );
  NAND2_X1 U6027 ( .A1(n9307), .A2(n4579), .ZN(n4578) );
  NAND2_X1 U6028 ( .A1(n9307), .A2(n4593), .ZN(n4592) );
  NAND2_X1 U6029 ( .A1(n4578), .A2(n4583), .ZN(n9246) );
  NAND3_X1 U6030 ( .A1(n4586), .A2(n4587), .A3(n4589), .ZN(n4584) );
  INV_X1 U6031 ( .A(n9105), .ZN(n4593) );
  NAND2_X2 U6032 ( .A1(n5658), .A2(n5667), .ZN(n4949) );
  XNOR2_X2 U6033 ( .A(n4602), .B(n4874), .ZN(n5667) );
  OAI21_X1 U6034 ( .B1(n9246), .B2(n9109), .A(n9108), .ZN(n9233) );
  NOR2_X1 U6035 ( .A1(n9199), .A2(n9114), .ZN(n9191) );
  OAI21_X1 U6036 ( .B1(n9317), .B2(n9319), .A(n9102), .ZN(n9307) );
  NAND2_X1 U6037 ( .A1(n9191), .A2(n9115), .ZN(n9174) );
  AOI21_X1 U6038 ( .B1(n9353), .B2(n9352), .A(n9099), .ZN(n9335) );
  NOR2_X1 U6039 ( .A1(n8121), .A2(n4604), .ZN(n4603) );
  OAI21_X1 U6040 ( .B1(n8499), .B2(n8270), .A(n4610), .ZN(n8484) );
  NOR2_X1 U6041 ( .A1(n8642), .A2(n8643), .ZN(n8641) );
  NAND2_X1 U6042 ( .A1(n4621), .A2(n4619), .ZN(n8595) );
  NAND2_X1 U6043 ( .A1(n8642), .A2(n4284), .ZN(n4621) );
  NOR2_X1 U6044 ( .A1(n8641), .A2(n8090), .ZN(n8618) );
  AOI21_X2 U6045 ( .B1(n7340), .B2(n4297), .A(n4639), .ZN(n9738) );
  NAND2_X1 U6046 ( .A1(n4643), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U6047 ( .A1(n4990), .A2(n4655), .ZN(n4653) );
  NAND2_X1 U6048 ( .A1(n4653), .A2(n4654), .ZN(n5017) );
  INV_X1 U6049 ( .A(n4658), .ZN(n5470) );
  NAND2_X1 U6050 ( .A1(n5497), .A2(n4675), .ZN(n4674) );
  OAI21_X1 U6051 ( .B1(n5099), .B2(n4684), .A(n4681), .ZN(n5142) );
  OAI21_X1 U6052 ( .B1(n5165), .B2(n4694), .A(n4328), .ZN(n5206) );
  NAND2_X1 U6053 ( .A1(n6370), .A2(n6373), .ZN(n5694) );
  OR2_X2 U6054 ( .A1(n5670), .A2(n6707), .ZN(n4700) );
  AND2_X4 U6055 ( .A1(n4700), .A2(n5954), .ZN(n5743) );
  NOR2_X1 U6056 ( .A1(n4700), .A2(n9250), .ZN(n6871) );
  NAND2_X1 U6057 ( .A1(n5679), .A2(n4700), .ZN(n5746) );
  AOI21_X1 U6058 ( .B1(n5678), .B2(n4700), .A(n9207), .ZN(n6709) );
  NAND2_X1 U6059 ( .A1(n8873), .A2(n4702), .ZN(n4701) );
  NAND2_X1 U6060 ( .A1(n7627), .A2(n4711), .ZN(n4709) );
  NAND2_X1 U6061 ( .A1(n4709), .A2(n4710), .ZN(n7669) );
  NAND2_X1 U6062 ( .A1(n4713), .A2(n4714), .ZN(n7553) );
  NAND2_X1 U6063 ( .A1(n7375), .A2(n4715), .ZN(n4713) );
  NAND2_X1 U6064 ( .A1(n7375), .A2(n5742), .ZN(n7431) );
  AOI21_X1 U6065 ( .B1(n4715), .B2(n4718), .A(n4317), .ZN(n4714) );
  AND2_X1 U6066 ( .A1(n4716), .A2(n7434), .ZN(n4715) );
  NAND2_X1 U6067 ( .A1(n8914), .A2(n4723), .ZN(n4722) );
  NAND2_X1 U6068 ( .A1(n8905), .A2(n4329), .ZN(n4726) );
  AOI21_X1 U6069 ( .B1(n8905), .B2(n5892), .A(n4316), .ZN(n8968) );
  INV_X1 U6070 ( .A(n4731), .ZN(n5519) );
  INV_X1 U6071 ( .A(n8051), .ZN(n4740) );
  INV_X1 U6072 ( .A(n7864), .ZN(n4741) );
  INV_X1 U6073 ( .A(n7851), .ZN(n4742) );
  NAND3_X1 U6074 ( .A1(n7893), .A2(n7892), .A3(n4310), .ZN(n4744) );
  NAND3_X1 U6075 ( .A1(n7893), .A2(n7892), .A3(n8068), .ZN(n8067) );
  NAND3_X1 U6076 ( .A1(n6460), .A2(n8828), .A3(n6515), .ZN(n4748) );
  NAND3_X1 U6077 ( .A1(n6019), .A2(n4817), .A3(n5957), .ZN(n4749) );
  NAND2_X1 U6078 ( .A1(n4749), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U6079 ( .A1(n4762), .A2(n6700), .ZN(n6702) );
  OAI21_X1 U6080 ( .B1(n6859), .B2(n6857), .A(n4762), .ZN(n9661) );
  NAND2_X1 U6081 ( .A1(n6857), .A2(n6699), .ZN(n4762) );
  NAND2_X1 U6082 ( .A1(n9088), .A2(n4763), .ZN(n9136) );
  NAND2_X1 U6083 ( .A1(n9285), .A2(n4322), .ZN(n4765) );
  NAND2_X1 U6084 ( .A1(n4765), .A2(n4766), .ZN(n9252) );
  NAND2_X1 U6085 ( .A1(n4777), .A2(n4775), .ZN(n9577) );
  NAND2_X1 U6086 ( .A1(n7476), .A2(n4778), .ZN(n7605) );
  NAND2_X1 U6087 ( .A1(n7091), .A2(n4324), .ZN(n7356) );
  NOR2_X1 U6088 ( .A1(n4991), .A2(n4783), .ZN(n5018) );
  NAND2_X1 U6089 ( .A1(n4873), .A2(n4793), .ZN(n4867) );
  NAND2_X1 U6090 ( .A1(n4873), .A2(n4874), .ZN(n4869) );
  NAND2_X1 U6091 ( .A1(n6724), .A2(n6760), .ZN(n8170) );
  INV_X1 U6092 ( .A(n6724), .ZN(n6668) );
  NAND2_X1 U6093 ( .A1(n8454), .A2(n4325), .ZN(n4795) );
  OAI211_X1 U6094 ( .C1(n8454), .C2(n4800), .A(n4796), .B(n4795), .ZN(n8713)
         );
  NAND2_X1 U6095 ( .A1(n8454), .A2(n8461), .ZN(n4802) );
  NOR2_X2 U6096 ( .A1(n5975), .A2(n4818), .ZN(n6214) );
  NOR2_X1 U6097 ( .A1(n8495), .A2(n8500), .ZN(n8494) );
  NAND2_X1 U6098 ( .A1(n8944), .A2(n8943), .ZN(n6889) );
  NAND2_X1 U6099 ( .A1(n5847), .A2(n8956), .ZN(n8858) );
  NOR2_X2 U6100 ( .A1(n8588), .A2(n8767), .ZN(n8573) );
  NAND3_X1 U6101 ( .A1(n8577), .A2(n8563), .A3(n8564), .ZN(n8562) );
  NAND3_X1 U6102 ( .A1(n8531), .A2(n8532), .A3(n8533), .ZN(n8507) );
  NAND2_X1 U6103 ( .A1(n6452), .A2(n6454), .ZN(n8162) );
  OR2_X1 U6104 ( .A1(n7226), .A2(n8120), .ZN(n7228) );
  CLKBUF_X1 U6105 ( .A(n9365), .Z(n9367) );
  NAND2_X1 U6106 ( .A1(n6298), .A2(n4837), .ZN(n6085) );
  OR2_X1 U6107 ( .A1(n6214), .A2(n6071), .ZN(n6215) );
  NAND2_X1 U6108 ( .A1(n6449), .A2(n6420), .ZN(n9856) );
  NAND2_X2 U6109 ( .A1(n8173), .A2(n8171), .ZN(n8120) );
  XNOR2_X1 U6110 ( .A(n6213), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U6111 ( .A1(n6216), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6213) );
  NAND2_X1 U6112 ( .A1(n6750), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6465) );
  NOR2_X1 U6113 ( .A1(n4949), .A2(n4927), .ZN(n4828) );
  AND2_X1 U6114 ( .A1(n5082), .A2(n4923), .ZN(n4829) );
  OR2_X1 U6115 ( .A1(n9069), .A2(n9068), .ZN(n4830) );
  OR2_X1 U6116 ( .A1(n9041), .A2(n9262), .ZN(n4831) );
  OR2_X1 U6117 ( .A1(n4439), .A2(n9248), .ZN(n4832) );
  OR2_X1 U6118 ( .A1(n9165), .A2(n8977), .ZN(n4833) );
  OR2_X1 U6119 ( .A1(n8771), .A2(n8580), .ZN(n4834) );
  INV_X1 U6120 ( .A(n8409), .ZN(n8660) );
  INV_X1 U6121 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5131) );
  AND2_X1 U6122 ( .A1(n5141), .A2(n5123), .ZN(n4836) );
  AND2_X1 U6123 ( .A1(n5454), .A2(n5453), .ZN(n9089) );
  INV_X1 U6124 ( .A(n9697), .ZN(n9694) );
  AND2_X2 U6125 ( .A1(n6663), .A2(n6289), .ZN(n9697) );
  INV_X2 U6126 ( .A(n9688), .ZN(n9530) );
  AND3_X1 U6127 ( .A1(n5375), .A2(n5374), .A3(n5373), .ZN(n9204) );
  AND3_X1 U6128 ( .A1(n5343), .A2(n5342), .A3(n5341), .ZN(n9218) );
  INV_X1 U6129 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6071) );
  INV_X1 U6130 ( .A(n9073), .ZN(n9274) );
  AND3_X1 U6131 ( .A1(n5969), .A2(n6417), .A3(n6415), .ZN(n4837) );
  INV_X1 U6132 ( .A(n8580), .ZN(n8609) );
  INV_X1 U6133 ( .A(n9435), .ZN(n9189) );
  INV_X1 U6134 ( .A(n9476), .ZN(n9069) );
  OR2_X1 U6135 ( .A1(n6476), .A2(n6436), .ZN(n9895) );
  NAND2_X1 U6136 ( .A1(n7165), .A2(n8613), .ZN(n9779) );
  INV_X1 U6137 ( .A(n9458), .ZN(n9041) );
  XOR2_X1 U6138 ( .A(n5654), .B(n9207), .Z(n4838) );
  INV_X1 U6139 ( .A(n6707), .ZN(n6759) );
  INV_X1 U6140 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4851) );
  INV_X1 U6141 ( .A(n7848), .ZN(n7849) );
  INV_X1 U6142 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6415) );
  INV_X1 U6143 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6378) );
  NOR2_X1 U6144 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5960) );
  INV_X1 U6145 ( .A(n9296), .ZN(n9068) );
  NOR2_X1 U6146 ( .A1(n7850), .A2(n7849), .ZN(n7851) );
  INV_X1 U6147 ( .A(n7876), .ZN(n7869) );
  INV_X1 U6148 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7117) );
  OR2_X1 U6149 ( .A1(n8732), .A2(n8464), .ZN(n8419) );
  NAND2_X1 U6150 ( .A1(n8307), .A2(n6456), .ZN(n6730) );
  INV_X1 U6151 ( .A(n7630), .ZN(n5764) );
  INV_X1 U6152 ( .A(n5715), .ZN(n5713) );
  INV_X1 U6153 ( .A(n5258), .ZN(n5257) );
  INV_X1 U6154 ( .A(n9089), .ZN(n9090) );
  OR2_X1 U6155 ( .A1(n5294), .A2(n5293), .ZN(n5315) );
  INV_X1 U6156 ( .A(SI_22_), .ZN(n5308) );
  INV_X1 U6157 ( .A(n7940), .ZN(n7734) );
  INV_X1 U6158 ( .A(n7020), .ZN(n6913) );
  OR2_X1 U6159 ( .A1(n7830), .A2(n7991), .ZN(n7858) );
  OR2_X1 U6160 ( .A1(n7118), .A2(n7117), .ZN(n7120) );
  INV_X1 U6161 ( .A(n8913), .ZN(n5865) );
  OR2_X1 U6162 ( .A1(n5045), .A2(n4860), .ZN(n5075) );
  INV_X1 U6163 ( .A(n9543), .ZN(n4862) );
  OR2_X1 U6164 ( .A1(n5132), .A2(n5131), .ZN(n5149) );
  NAND2_X1 U6165 ( .A1(n4955), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4935) );
  AND2_X1 U6166 ( .A1(n6759), .A2(n9250), .ZN(n5934) );
  INV_X1 U6167 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5069) );
  INV_X1 U6168 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5126) );
  INV_X1 U6169 ( .A(n8463), .ZN(n8420) );
  OR3_X1 U6170 ( .A1(n7583), .A2(n7582), .A3(n7581), .ZN(n7747) );
  OR2_X1 U6171 ( .A1(n7754), .A2(n7753), .ZN(n7763) );
  INV_X1 U6172 ( .A(n8073), .ZN(n8080) );
  AND3_X1 U6173 ( .A1(n6222), .A2(n6221), .A3(n6220), .ZN(n8115) );
  INV_X1 U6174 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7582) );
  INV_X1 U6175 ( .A(n8411), .ZN(n8644) );
  INV_X1 U6176 ( .A(n8407), .ZN(n8668) );
  OR2_X1 U6177 ( .A1(n6817), .A2(n4376), .ZN(n6727) );
  INV_X1 U6178 ( .A(n8185), .ZN(n9858) );
  OR2_X1 U6179 ( .A1(n5424), .A2(n5943), .ZN(n5447) );
  NAND2_X1 U6180 ( .A1(n5193), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5236) );
  INV_X1 U6181 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7276) );
  NOR2_X1 U6182 ( .A1(n6010), .A2(n9551), .ZN(n9032) );
  INV_X1 U6183 ( .A(n5934), .ZN(n6880) );
  INV_X1 U6184 ( .A(n9427), .ZN(n9165) );
  NOR2_X1 U6185 ( .A1(n9435), .A2(n9177), .ZN(n9083) );
  INV_X1 U6186 ( .A(n9075), .ZN(n9248) );
  INV_X1 U6187 ( .A(n9297), .ZN(n9263) );
  OR2_X1 U6188 ( .A1(n6292), .A2(n6880), .ZN(n7003) );
  AND2_X1 U6189 ( .A1(n7473), .A2(n7609), .ZN(n7478) );
  OR2_X1 U6190 ( .A1(n6292), .A2(n6716), .ZN(n9635) );
  AND2_X1 U6191 ( .A1(n6714), .A2(n6713), .ZN(n9370) );
  INV_X1 U6192 ( .A(n9568), .ZN(n9680) );
  AND2_X1 U6193 ( .A1(n5415), .A2(n5395), .ZN(n5413) );
  OAI21_X1 U6194 ( .B1(n8006), .B2(n7763), .A(n7762), .ZN(n8027) );
  INV_X1 U6195 ( .A(n6750), .ZN(n7984) );
  NAND2_X1 U6196 ( .A1(n6514), .A2(n6513), .ZN(n9718) );
  INV_X1 U6197 ( .A(n9718), .ZN(n9713) );
  AND2_X1 U6198 ( .A1(n8241), .A2(n8564), .ZN(n8579) );
  NAND2_X1 U6199 ( .A1(n9815), .A2(n6435), .ZN(n7153) );
  NAND2_X1 U6200 ( .A1(n9822), .A2(n6449), .ZN(n9889) );
  INV_X1 U6201 ( .A(n9894), .ZN(n8796) );
  NAND2_X1 U6202 ( .A1(n9757), .A2(n9856), .ZN(n9894) );
  OR2_X1 U6203 ( .A1(n6432), .A2(n7158), .ZN(n6476) );
  NAND2_X1 U6204 ( .A1(n6480), .A2(n7154), .ZN(n9782) );
  AND2_X1 U6205 ( .A1(n6054), .A2(n6053), .ZN(n7313) );
  INV_X1 U6206 ( .A(n8912), .ZN(n8917) );
  NAND2_X1 U6207 ( .A1(n5940), .A2(n6256), .ZN(n8982) );
  AND2_X2 U6208 ( .A1(n5915), .A2(n6880), .ZN(n9568) );
  AND2_X1 U6209 ( .A1(n5464), .A2(n5463), .ZN(n9144) );
  AND4_X1 U6210 ( .A1(n5241), .A2(n5240), .A3(n5239), .A4(n5238), .ZN(n9275)
         );
  NOR2_X1 U6211 ( .A1(n5993), .A2(n6356), .ZN(n9616) );
  INV_X1 U6212 ( .A(n9616), .ZN(n9017) );
  INV_X1 U6213 ( .A(n9029), .ZN(n9610) );
  INV_X1 U6214 ( .A(n9086), .ZN(n9154) );
  AND2_X1 U6215 ( .A1(n7003), .A2(n5900), .ZN(n7004) );
  AND2_X1 U6216 ( .A1(n6717), .A2(n6716), .ZN(n9311) );
  INV_X1 U6217 ( .A(n9370), .ZN(n9640) );
  INV_X1 U6218 ( .A(n9595), .ZN(n9254) );
  OR2_X1 U6219 ( .A1(n6881), .A2(n6707), .ZN(n9682) );
  INV_X1 U6220 ( .A(n9678), .ZN(n9497) );
  NAND2_X1 U6221 ( .A1(n9643), .A2(n9510), .ZN(n9678) );
  NOR2_X1 U6222 ( .A1(n6870), .A2(n9533), .ZN(n6662) );
  NAND2_X1 U6223 ( .A1(n5916), .A2(n5918), .ZN(n9653) );
  AND2_X1 U6224 ( .A1(n5128), .A2(n5143), .ZN(n6954) );
  AND2_X1 U6225 ( .A1(n4995), .A2(n4994), .ZN(n9609) );
  NAND2_X1 U6226 ( .A1(n6670), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9818) );
  AND2_X1 U6227 ( .A1(n6675), .A2(n8613), .ZN(n9701) );
  NAND2_X1 U6228 ( .A1(n8384), .A2(n6460), .ZN(n9717) );
  NAND2_X1 U6229 ( .A1(n9779), .A2(n7164), .ZN(n9777) );
  INV_X2 U6230 ( .A(n9779), .ZN(n9775) );
  NOR2_X1 U6231 ( .A1(n9783), .A2(n9782), .ZN(n9799) );
  CLKBUF_X1 U6232 ( .A(n9799), .Z(n9819) );
  INV_X1 U6233 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6236) );
  INV_X1 U6234 ( .A(n8982), .ZN(n8906) );
  OR3_X1 U6235 ( .A1(n9568), .A2(n5942), .A3(n6717), .ZN(n8991) );
  INV_X1 U6236 ( .A(n9218), .ZN(n9192) );
  OR2_X1 U6237 ( .A1(n6010), .A2(n6009), .ZN(n9030) );
  NAND2_X1 U6238 ( .A1(n6013), .A2(n6012), .ZN(n9039) );
  NAND2_X1 U6239 ( .A1(n9650), .A2(n7004), .ZN(n9364) );
  INV_X2 U6240 ( .A(n9650), .ZN(n9647) );
  OR2_X1 U6241 ( .A1(n9492), .A2(n9491), .ZN(n9527) );
  NAND2_X1 U6242 ( .A1(n6663), .A2(n6662), .ZN(n9688) );
  AND2_X1 U6243 ( .A1(n9654), .A2(n9653), .ZN(n9659) );
  AND2_X1 U6244 ( .A1(n5954), .A2(n5666), .ZN(n9654) );
  INV_X1 U6245 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7470) );
  INV_X1 U6246 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6244) );
  INV_X1 U6247 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6050) );
  NOR2_X1 U6248 ( .A1(n9941), .A2(n9940), .ZN(n9939) );
  OAI21_X1 U6249 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9930), .ZN(n9928) );
  NOR2_X1 U6250 ( .A1(n6480), .A2(n9818), .ZN(P2_U3966) );
  NOR2_X1 U6251 ( .A1(n6012), .A2(P1_U3084), .ZN(P1_U4006) );
  NOR2_X2 U6252 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4950) );
  NAND2_X1 U6253 ( .A1(n4950), .A2(n4839), .ZN(n4978) );
  NOR2_X1 U6254 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4847) );
  NOR2_X1 U6255 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4846) );
  NAND4_X1 U6256 ( .A1(n4847), .A2(n4846), .A3(n4845), .A4(n5063), .ZN(n4849)
         );
  NAND4_X1 U6257 ( .A1(n5068), .A2(n5211), .A3(n5126), .A4(n5067), .ZN(n4848)
         );
  NAND2_X1 U6258 ( .A1(n4867), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4853) );
  MUX2_X1 U6259 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4853), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n4855) );
  INV_X1 U6260 ( .A(n4854), .ZN(n9536) );
  AND2_X4 U6261 ( .A1(n9543), .A2(n4856), .ZN(n4955) );
  NAND2_X1 U6262 ( .A1(n4955), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4866) );
  INV_X1 U6263 ( .A(n4942), .ZN(n5026) );
  NAND2_X1 U6264 ( .A1(n5482), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n4865) );
  AND2_X2 U6265 ( .A1(n9540), .A2(n9543), .ZN(n4969) );
  NAND3_X1 U6266 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n4998) );
  INV_X1 U6267 ( .A(n4998), .ZN(n4857) );
  NAND2_X1 U6268 ( .A1(n4857), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5010) );
  INV_X1 U6269 ( .A(n5010), .ZN(n4858) );
  NAND2_X1 U6270 ( .A1(n4858), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5028) );
  INV_X1 U6271 ( .A(n5028), .ZN(n4859) );
  NAND2_X1 U6272 ( .A1(n4859), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U6273 ( .A1(n5045), .A2(n4860), .ZN(n4861) );
  AND2_X1 U6274 ( .A1(n5075), .A2(n4861), .ZN(n7656) );
  NAND2_X1 U6275 ( .A1(n5277), .A2(n7656), .ZN(n4864) );
  NAND2_X1 U6276 ( .A1(n5340), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4863) );
  INV_X1 U6277 ( .A(n4867), .ZN(n4868) );
  AOI21_X1 U6278 ( .B1(n4870), .B2(n9535), .A(n4868), .ZN(n4872) );
  NAND2_X1 U6279 ( .A1(n4872), .A2(n4871), .ZN(n5658) );
  NAND2_X1 U6280 ( .A1(n4875), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4878) );
  INV_X1 U6281 ( .A(n4878), .ZN(n4876) );
  NAND2_X1 U6282 ( .A1(n4876), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n4879) );
  NAND2_X1 U6283 ( .A1(n4878), .A2(n4877), .ZN(n5085) );
  INV_X1 U6284 ( .A(n6404), .ZN(n6400) );
  INV_X1 U6285 ( .A(SI_1_), .ZN(n4881) );
  XNOR2_X1 U6286 ( .A(n4883), .B(n4881), .ZN(n4929) );
  INV_X1 U6287 ( .A(n4929), .ZN(n4882) );
  MUX2_X1 U6288 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4888), .Z(n4928) );
  INV_X1 U6289 ( .A(n4883), .ZN(n4884) );
  NAND2_X1 U6290 ( .A1(n4884), .A2(SI_1_), .ZN(n4885) );
  INV_X1 U6291 ( .A(n4947), .ZN(n4886) );
  MUX2_X1 U6292 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n4888), .Z(n4890) );
  INV_X1 U6293 ( .A(SI_3_), .ZN(n4889) );
  XNOR2_X1 U6294 ( .A(n4890), .B(n4889), .ZN(n4962) );
  NAND2_X1 U6295 ( .A1(n4961), .A2(n4962), .ZN(n4892) );
  NAND2_X1 U6296 ( .A1(n4890), .A2(SI_3_), .ZN(n4891) );
  NAND2_X1 U6297 ( .A1(n4892), .A2(n4891), .ZN(n4975) );
  INV_X1 U6298 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6033) );
  MUX2_X1 U6299 ( .A(n6818), .B(n6033), .S(n4888), .Z(n4893) );
  XNOR2_X1 U6300 ( .A(n4893), .B(SI_4_), .ZN(n4976) );
  NAND2_X1 U6301 ( .A1(n4975), .A2(n4976), .ZN(n4896) );
  INV_X1 U6302 ( .A(n4893), .ZN(n4894) );
  NAND2_X1 U6303 ( .A1(n4894), .A2(SI_4_), .ZN(n4895) );
  NAND2_X1 U6304 ( .A1(n4896), .A2(n4895), .ZN(n4990) );
  INV_X1 U6305 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n4897) );
  MUX2_X1 U6306 ( .A(n6832), .B(n4897), .S(n4888), .Z(n4898) );
  XNOR2_X1 U6307 ( .A(n4898), .B(SI_5_), .ZN(n4989) );
  INV_X1 U6308 ( .A(n4898), .ZN(n4899) );
  NAND2_X1 U6309 ( .A1(n4899), .A2(SI_5_), .ZN(n4900) );
  MUX2_X1 U6310 ( .A(n6927), .B(n6037), .S(n4888), .Z(n4901) );
  XNOR2_X1 U6311 ( .A(n4901), .B(SI_6_), .ZN(n5004) );
  INV_X1 U6312 ( .A(n4901), .ZN(n4902) );
  MUX2_X1 U6313 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6445), .Z(n4908) );
  XNOR2_X1 U6314 ( .A(n4908), .B(SI_7_), .ZN(n5016) );
  INV_X1 U6315 ( .A(n5016), .ZN(n4903) );
  NAND2_X1 U6316 ( .A1(n5017), .A2(n4903), .ZN(n5035) );
  INV_X1 U6317 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6059) );
  INV_X1 U6318 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6060) );
  MUX2_X1 U6319 ( .A(n6059), .B(n6060), .S(n6445), .Z(n4905) );
  INV_X1 U6320 ( .A(SI_9_), .ZN(n4904) );
  NAND2_X1 U6321 ( .A1(n4905), .A2(n4904), .ZN(n4915) );
  INV_X1 U6322 ( .A(n4905), .ZN(n4906) );
  NAND2_X1 U6323 ( .A1(n4906), .A2(SI_9_), .ZN(n4907) );
  NAND2_X1 U6324 ( .A1(n4915), .A2(n4907), .ZN(n4912) );
  NAND2_X1 U6325 ( .A1(n4908), .A2(SI_7_), .ZN(n5034) );
  INV_X1 U6326 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7113) );
  MUX2_X1 U6327 ( .A(n7113), .B(n6186), .S(n6445), .Z(n4914) );
  INV_X1 U6328 ( .A(n4914), .ZN(n4909) );
  NAND2_X1 U6329 ( .A1(n4909), .A2(SI_8_), .ZN(n5036) );
  NAND2_X1 U6330 ( .A1(n5034), .A2(n5036), .ZN(n4910) );
  NOR2_X1 U6331 ( .A1(n4912), .A2(n4910), .ZN(n4911) );
  NAND2_X1 U6332 ( .A1(n5035), .A2(n4911), .ZN(n4919) );
  INV_X1 U6333 ( .A(n4912), .ZN(n5057) );
  INV_X1 U6334 ( .A(SI_8_), .ZN(n4913) );
  NAND2_X1 U6335 ( .A1(n4914), .A2(n4913), .ZN(n5054) );
  INV_X1 U6336 ( .A(n5054), .ZN(n4917) );
  INV_X1 U6337 ( .A(n4915), .ZN(n4916) );
  AOI21_X1 U6338 ( .B1(n5057), .B2(n4917), .A(n4916), .ZN(n4918) );
  MUX2_X1 U6339 ( .A(n6055), .B(n6050), .S(n6445), .Z(n4921) );
  INV_X1 U6340 ( .A(SI_10_), .ZN(n4920) );
  NAND2_X1 U6341 ( .A1(n4921), .A2(n4920), .ZN(n5082) );
  INV_X1 U6342 ( .A(n4921), .ZN(n4922) );
  NAND2_X1 U6343 ( .A1(n4922), .A2(SI_10_), .ZN(n4923) );
  XNOR2_X1 U6344 ( .A(n5081), .B(n4829), .ZN(n7314) );
  AND2_X4 U6345 ( .A1(n4949), .A2(n6445), .ZN(n4960) );
  NAND2_X1 U6346 ( .A1(n7314), .A2(n4960), .ZN(n4925) );
  NAND2_X1 U6347 ( .A1(n4977), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n4924) );
  OAI211_X1 U6348 ( .C1(n4949), .C2(n6400), .A(n4925), .B(n4924), .ZN(n7619)
         );
  NAND2_X1 U6349 ( .A1(n9636), .A2(n7619), .ZN(n5533) );
  NAND2_X1 U6350 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4926) );
  XNOR2_X1 U6351 ( .A(n4926), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6034) );
  INV_X1 U6352 ( .A(n6034), .ZN(n4927) );
  XNOR2_X1 U6353 ( .A(n4929), .B(n4928), .ZN(n6028) );
  NAND2_X1 U6354 ( .A1(n4960), .A2(n6028), .ZN(n4930) );
  NAND2_X1 U6355 ( .A1(n4954), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4933) );
  NAND2_X1 U6356 ( .A1(n4969), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4932) );
  NAND4_X1 U6357 ( .A1(n4935), .A2(n4934), .A3(n4933), .A4(n4932), .ZN(n5682)
         );
  NAND2_X1 U6358 ( .A1(n4955), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4939) );
  NAND2_X1 U6359 ( .A1(n4954), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4937) );
  NAND2_X1 U6360 ( .A1(n4969), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4936) );
  NAND4_X2 U6361 ( .A1(n4939), .A2(n4938), .A3(n4937), .A4(n4936), .ZN(n5674)
         );
  NAND2_X1 U6362 ( .A1(n6445), .A2(SI_0_), .ZN(n4940) );
  XNOR2_X1 U6363 ( .A(n4940), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9554) );
  MUX2_X1 U6364 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9554), .S(n4949), .Z(n6883) );
  INV_X1 U6365 ( .A(n6883), .ZN(n6704) );
  NOR2_X1 U6366 ( .A1(n5674), .A2(n6704), .ZN(n6858) );
  CLKBUF_X1 U6367 ( .A(n5682), .Z(n5689) );
  INV_X1 U6368 ( .A(n5689), .ZN(n6698) );
  NAND2_X1 U6369 ( .A1(n6698), .A2(n5683), .ZN(n4941) );
  NAND2_X1 U6370 ( .A1(n4942), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n4946) );
  NAND2_X1 U6371 ( .A1(n4955), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4945) );
  NAND2_X1 U6372 ( .A1(n4954), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4944) );
  NAND2_X1 U6373 ( .A1(n4969), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n4943) );
  NAND4_X1 U6374 ( .A1(n4946), .A2(n4945), .A3(n4944), .A4(n4943), .ZN(n5698)
         );
  INV_X2 U6375 ( .A(n5698), .ZN(n7043) );
  XNOR2_X1 U6376 ( .A(n4948), .B(n4947), .ZN(n6017) );
  NAND2_X1 U6377 ( .A1(n4960), .A2(n6017), .ZN(n4953) );
  NAND2_X1 U6378 ( .A1(n5982), .A2(n6396), .ZN(n4952) );
  NAND2_X1 U6379 ( .A1(n4977), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4951) );
  XNOR2_X2 U6380 ( .A(n7043), .B(n8948), .ZN(n6701) );
  INV_X1 U6381 ( .A(n6701), .ZN(n6710) );
  NAND2_X1 U6382 ( .A1(n6711), .A2(n6710), .ZN(n5560) );
  INV_X1 U6383 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7050) );
  NAND2_X1 U6384 ( .A1(n4969), .A2(n7050), .ZN(n4959) );
  NAND2_X1 U6385 ( .A1(n4954), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4957) );
  NAND2_X1 U6386 ( .A1(n4955), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4956) );
  XNOR2_X1 U6387 ( .A(n4961), .B(n4962), .ZN(n6766) );
  NAND2_X1 U6388 ( .A1(n4977), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4968) );
  INV_X1 U6389 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4963) );
  NAND2_X1 U6390 ( .A1(n4964), .A2(n4963), .ZN(n4965) );
  NAND2_X1 U6391 ( .A1(n4965), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4966) );
  XNOR2_X1 U6392 ( .A(n4966), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U6393 ( .A1(n5982), .A2(n6270), .ZN(n4967) );
  NAND2_X1 U6394 ( .A1(n7032), .A2(n7051), .ZN(n5564) );
  NAND2_X1 U6395 ( .A1(n7043), .A2(n8948), .ZN(n5559) );
  AND2_X1 U6396 ( .A1(n5564), .A2(n5559), .ZN(n5618) );
  NAND2_X1 U6397 ( .A1(n5560), .A2(n5618), .ZN(n5089) );
  INV_X1 U6398 ( .A(n7032), .ZN(n9002) );
  NAND2_X1 U6399 ( .A1(n9002), .A2(n5706), .ZN(n5527) );
  NAND2_X1 U6400 ( .A1(n5089), .A2(n5527), .ZN(n6967) );
  NAND2_X1 U6401 ( .A1(n4955), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n4974) );
  BUF_X1 U6402 ( .A(n4969), .Z(n5277) );
  INV_X1 U6403 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n4970) );
  XNOR2_X1 U6404 ( .A(n4970), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7027) );
  NAND2_X1 U6405 ( .A1(n5277), .A2(n7027), .ZN(n4972) );
  NAND2_X1 U6406 ( .A1(n4954), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4971) );
  XNOR2_X1 U6407 ( .A(n4975), .B(n4976), .ZN(n6816) );
  NAND2_X1 U6408 ( .A1(n4977), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4981) );
  NAND2_X1 U6409 ( .A1(n4978), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4979) );
  XNOR2_X1 U6410 ( .A(n4979), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U6411 ( .A1(n5982), .A2(n6032), .ZN(n4980) );
  NAND2_X1 U6412 ( .A1(n7246), .A2(n7059), .ZN(n5622) );
  NAND2_X1 U6413 ( .A1(n4942), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n4988) );
  NAND2_X1 U6414 ( .A1(n5340), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4987) );
  INV_X1 U6415 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n4983) );
  NAND2_X1 U6416 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n4982) );
  NAND2_X1 U6417 ( .A1(n4983), .A2(n4982), .ZN(n4984) );
  AND2_X1 U6418 ( .A1(n4998), .A2(n4984), .ZN(n7250) );
  NAND2_X1 U6419 ( .A1(n5277), .A2(n7250), .ZN(n4986) );
  NAND2_X1 U6420 ( .A1(n4955), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4985) );
  XNOR2_X1 U6421 ( .A(n4990), .B(n4989), .ZN(n6831) );
  NAND2_X1 U6422 ( .A1(n4977), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n4997) );
  NAND2_X1 U6423 ( .A1(n4991), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4992) );
  MUX2_X1 U6424 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4992), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n4995) );
  INV_X1 U6425 ( .A(n4993), .ZN(n4994) );
  NAND2_X1 U6426 ( .A1(n5982), .A2(n9609), .ZN(n4996) );
  OAI211_X1 U6427 ( .C1(n5008), .C2(n6831), .A(n4997), .B(n4996), .ZN(n7089)
         );
  INV_X1 U6428 ( .A(n7089), .ZN(n7247) );
  NAND2_X1 U6429 ( .A1(n9000), .A2(n7247), .ZN(n5561) );
  INV_X1 U6430 ( .A(n7246), .ZN(n9001) );
  INV_X1 U6431 ( .A(n7059), .ZN(n7033) );
  NAND2_X1 U6432 ( .A1(n9001), .A2(n7033), .ZN(n5526) );
  NAND2_X1 U6433 ( .A1(n5561), .A2(n5526), .ZN(n5565) );
  AOI21_X1 U6434 ( .B1(n6967), .B2(n5622), .A(n5565), .ZN(n5025) );
  NAND2_X1 U6435 ( .A1(n4942), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U6436 ( .A1(n4955), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5002) );
  INV_X1 U6437 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U6438 ( .A1(n4998), .A2(n6136), .ZN(n4999) );
  AND2_X1 U6439 ( .A1(n5010), .A2(n4999), .ZN(n7370) );
  NAND2_X1 U6440 ( .A1(n5277), .A2(n7370), .ZN(n5001) );
  NAND2_X1 U6441 ( .A1(n5340), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5000) );
  NAND2_X1 U6442 ( .A1(n4977), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5007) );
  OR2_X1 U6443 ( .A1(n4993), .A2(n9535), .ZN(n5005) );
  XNOR2_X1 U6444 ( .A(n5005), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6695) );
  NAND2_X1 U6445 ( .A1(n5982), .A2(n6695), .ZN(n5006) );
  NAND2_X1 U6446 ( .A1(n7438), .A2(n7523), .ZN(n5624) );
  INV_X1 U6447 ( .A(n7438), .ZN(n8999) );
  NAND2_X1 U6448 ( .A1(n8999), .A2(n7380), .ZN(n7085) );
  NAND2_X1 U6449 ( .A1(n7379), .A2(n7089), .ZN(n5623) );
  NAND2_X1 U6450 ( .A1(n7359), .A2(n5623), .ZN(n5024) );
  NAND2_X1 U6451 ( .A1(n4955), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5015) );
  NAND2_X1 U6452 ( .A1(n4942), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5014) );
  INV_X1 U6453 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5009) );
  NAND2_X1 U6454 ( .A1(n5010), .A2(n5009), .ZN(n5011) );
  AND2_X1 U6455 ( .A1(n5028), .A2(n5011), .ZN(n7442) );
  NAND2_X1 U6456 ( .A1(n4969), .A2(n7442), .ZN(n5013) );
  NAND2_X1 U6457 ( .A1(n5340), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5012) );
  NAND4_X1 U6458 ( .A1(n5015), .A2(n5014), .A3(n5013), .A4(n5012), .ZN(n8998)
         );
  XNOR2_X1 U6459 ( .A(n5017), .B(n5016), .ZN(n6039) );
  NAND2_X1 U6460 ( .A1(n4960), .A2(n6039), .ZN(n5022) );
  NAND2_X1 U6461 ( .A1(n4977), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n5021) );
  OR2_X1 U6462 ( .A1(n5018), .A2(n9535), .ZN(n5019) );
  XNOR2_X1 U6463 ( .A(n5019), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U6464 ( .A1(n5982), .A2(n6335), .ZN(n5020) );
  NAND2_X1 U6465 ( .A1(n8998), .A2(n9675), .ZN(n5023) );
  AND2_X1 U6466 ( .A1(n7085), .A2(n5023), .ZN(n5569) );
  OAI21_X1 U6467 ( .B1(n5025), .B2(n5024), .A(n5569), .ZN(n5041) );
  NAND2_X1 U6468 ( .A1(n4955), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5033) );
  NAND2_X1 U6469 ( .A1(n5482), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5032) );
  INV_X1 U6470 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5027) );
  NAND2_X1 U6471 ( .A1(n5028), .A2(n5027), .ZN(n5029) );
  AND2_X1 U6472 ( .A1(n5043), .A2(n5029), .ZN(n7558) );
  NAND2_X1 U6473 ( .A1(n4969), .A2(n7558), .ZN(n5031) );
  NAND2_X1 U6474 ( .A1(n5340), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5030) );
  NAND2_X1 U6475 ( .A1(n5035), .A2(n5034), .ZN(n5056) );
  NAND2_X1 U6476 ( .A1(n5054), .A2(n5036), .ZN(n5055) );
  XNOR2_X1 U6477 ( .A(n5056), .B(n5055), .ZN(n7111) );
  NAND2_X1 U6478 ( .A1(n4960), .A2(n7111), .ZN(n5040) );
  NAND2_X1 U6479 ( .A1(n5037), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5038) );
  XNOR2_X1 U6480 ( .A(n5038), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6322) );
  NAND2_X1 U6481 ( .A1(n5982), .A2(n6322), .ZN(n5039) );
  OAI211_X1 U6482 ( .C1(n5050), .C2(n6186), .A(n5040), .B(n5039), .ZN(n7603)
         );
  NAND2_X1 U6483 ( .A1(n9637), .A2(n7603), .ZN(n7473) );
  INV_X1 U6484 ( .A(n8998), .ZN(n7563) );
  NAND2_X1 U6485 ( .A1(n7563), .A2(n7098), .ZN(n5091) );
  AND2_X1 U6486 ( .A1(n7473), .A2(n5091), .ZN(n7607) );
  NAND2_X1 U6487 ( .A1(n5041), .A2(n7607), .ZN(n5061) );
  NAND2_X1 U6488 ( .A1(n5043), .A2(n5042), .ZN(n5044) );
  AND2_X1 U6489 ( .A1(n5045), .A2(n5044), .ZN(n9646) );
  NAND2_X1 U6490 ( .A1(n4969), .A2(n9646), .ZN(n5049) );
  NAND2_X1 U6491 ( .A1(n5482), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5048) );
  NAND2_X1 U6492 ( .A1(n5340), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5047) );
  NAND2_X1 U6493 ( .A1(n4955), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5046) );
  NAND4_X1 U6494 ( .A1(n5049), .A2(n5048), .A3(n5047), .A4(n5046), .ZN(n8996)
         );
  INV_X1 U6495 ( .A(n5051), .ZN(n5052) );
  NAND2_X1 U6496 ( .A1(n5052), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5053) );
  XNOR2_X1 U6497 ( .A(n5053), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6308) );
  AOI22_X1 U6498 ( .A1(n4977), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5982), .B2(
        n6308), .ZN(n5060) );
  OAI21_X1 U6499 ( .B1(n5056), .B2(n5055), .A(n5054), .ZN(n5058) );
  XNOR2_X1 U6500 ( .A(n5058), .B(n5057), .ZN(n7285) );
  NAND2_X1 U6501 ( .A1(n7285), .A2(n4960), .ZN(n5059) );
  NAND2_X1 U6502 ( .A1(n5060), .A2(n5059), .ZN(n7635) );
  INV_X1 U6503 ( .A(n7635), .ZN(n9681) );
  INV_X1 U6504 ( .A(n7603), .ZN(n7557) );
  NAND2_X1 U6505 ( .A1(n8997), .A2(n7557), .ZN(n7609) );
  AND2_X1 U6506 ( .A1(n4295), .A2(n7609), .ZN(n5573) );
  NAND2_X1 U6507 ( .A1(n5061), .A2(n5573), .ZN(n5062) );
  INV_X1 U6508 ( .A(n8996), .ZN(n7661) );
  NAND2_X1 U6509 ( .A1(n7661), .A2(n7635), .ZN(n7612) );
  AND2_X1 U6510 ( .A1(n7612), .A2(n5533), .ZN(n7610) );
  INV_X1 U6511 ( .A(n9636), .ZN(n8995) );
  NAND2_X1 U6512 ( .A1(n8995), .A2(n9570), .ZN(n9093) );
  INV_X1 U6513 ( .A(n9093), .ZN(n7616) );
  NOR2_X1 U6514 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5064) );
  NAND2_X1 U6515 ( .A1(n5170), .A2(n5065), .ZN(n5173) );
  NOR2_X1 U6516 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5066) );
  XNOR2_X2 U6517 ( .A(n5070), .B(n5069), .ZN(n5678) );
  NAND2_X1 U6518 ( .A1(n5071), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5072) );
  XNOR2_X2 U6519 ( .A(n5072), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9207) );
  INV_X1 U6520 ( .A(n5947), .ZN(n5511) );
  NAND2_X1 U6521 ( .A1(n5482), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U6522 ( .A1(n4954), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5079) );
  INV_X1 U6523 ( .A(n5075), .ZN(n5073) );
  NAND2_X1 U6524 ( .A1(n5073), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5109) );
  INV_X1 U6525 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5074) );
  NAND2_X1 U6526 ( .A1(n5075), .A2(n5074), .ZN(n5076) );
  AND2_X1 U6527 ( .A1(n5109), .A2(n5076), .ZN(n9593) );
  NAND2_X1 U6528 ( .A1(n4969), .A2(n9593), .ZN(n5078) );
  NAND2_X1 U6529 ( .A1(n4955), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5077) );
  NAND2_X1 U6530 ( .A1(n5081), .A2(n4829), .ZN(n5083) );
  NAND2_X1 U6531 ( .A1(n5083), .A2(n5082), .ZN(n5099) );
  INV_X1 U6532 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5084) );
  MUX2_X1 U6533 ( .A(n5084), .B(n6062), .S(n6445), .Z(n5095) );
  XNOR2_X1 U6534 ( .A(n5095), .B(SI_11_), .ZN(n5094) );
  XNOR2_X1 U6535 ( .A(n5099), .B(n5094), .ZN(n7452) );
  NAND2_X1 U6536 ( .A1(n7452), .A2(n4960), .ZN(n5088) );
  NAND2_X1 U6537 ( .A1(n5085), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5086) );
  XNOR2_X1 U6538 ( .A(n5086), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6641) );
  AOI22_X1 U6539 ( .A1(n4977), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5982), .B2(
        n6641), .ZN(n5087) );
  NAND2_X1 U6540 ( .A1(n5088), .A2(n5087), .ZN(n9055) );
  NAND2_X1 U6541 ( .A1(n9391), .A2(n9055), .ZN(n9387) );
  NAND2_X1 U6542 ( .A1(n9056), .A2(n9600), .ZN(n9385) );
  AND2_X1 U6543 ( .A1(n5526), .A2(n5527), .ZN(n5620) );
  INV_X1 U6544 ( .A(n5623), .ZN(n5090) );
  NAND2_X1 U6545 ( .A1(n7355), .A2(n5624), .ZN(n7086) );
  NAND2_X1 U6546 ( .A1(n7608), .A2(n5091), .ZN(n7474) );
  NAND2_X1 U6547 ( .A1(n7474), .A2(n7609), .ZN(n5092) );
  NAND3_X1 U6548 ( .A1(n5092), .A2(n7612), .A3(n7473), .ZN(n5093) );
  NAND3_X1 U6549 ( .A1(n5093), .A2(n9093), .A3(n4295), .ZN(n5115) );
  INV_X1 U6550 ( .A(n5094), .ZN(n5098) );
  INV_X1 U6551 ( .A(n5095), .ZN(n5096) );
  NAND2_X1 U6552 ( .A1(n5096), .A2(SI_11_), .ZN(n5097) );
  MUX2_X1 U6553 ( .A(n6068), .B(n6064), .S(n6445), .Z(n5101) );
  INV_X1 U6554 ( .A(SI_12_), .ZN(n5100) );
  NAND2_X1 U6555 ( .A1(n5101), .A2(n5100), .ZN(n5118) );
  INV_X1 U6556 ( .A(n5101), .ZN(n5102) );
  NAND2_X1 U6557 ( .A1(n5102), .A2(SI_12_), .ZN(n5103) );
  NAND2_X1 U6558 ( .A1(n5118), .A2(n5103), .ZN(n5116) );
  XNOR2_X1 U6559 ( .A(n5117), .B(n5116), .ZN(n7538) );
  NAND2_X1 U6560 ( .A1(n7538), .A2(n4960), .ZN(n5106) );
  OR2_X1 U6561 ( .A1(n4334), .A2(n9535), .ZN(n5104) );
  XNOR2_X1 U6562 ( .A(n5104), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6642) );
  AOI22_X1 U6563 ( .A1(n4977), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5982), .B2(
        n6642), .ZN(n5105) );
  NAND2_X1 U6564 ( .A1(n4942), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5114) );
  NAND2_X1 U6565 ( .A1(n4955), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5113) );
  INV_X1 U6566 ( .A(n5109), .ZN(n5107) );
  NAND2_X1 U6567 ( .A1(n5107), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5132) );
  INV_X1 U6568 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U6569 ( .A1(n5109), .A2(n5108), .ZN(n5110) );
  AND2_X1 U6570 ( .A1(n5132), .A2(n5110), .ZN(n9401) );
  NAND2_X1 U6571 ( .A1(n4969), .A2(n9401), .ZN(n5112) );
  NAND2_X1 U6572 ( .A1(n5340), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5111) );
  NAND2_X1 U6573 ( .A1(n9506), .A2(n9589), .ZN(n5536) );
  NAND2_X1 U6574 ( .A1(n5115), .A2(n5536), .ZN(n5139) );
  INV_X1 U6575 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n5119) );
  MUX2_X1 U6576 ( .A(n5119), .B(n6070), .S(n6445), .Z(n5121) );
  INV_X1 U6577 ( .A(SI_13_), .ZN(n5120) );
  NAND2_X1 U6578 ( .A1(n5121), .A2(n5120), .ZN(n5141) );
  INV_X1 U6579 ( .A(n5121), .ZN(n5122) );
  NAND2_X1 U6580 ( .A1(n5122), .A2(SI_13_), .ZN(n5123) );
  XNOR2_X1 U6581 ( .A(n5140), .B(n4836), .ZN(n7577) );
  NAND2_X1 U6582 ( .A1(n7577), .A2(n4960), .ZN(n5130) );
  OR2_X1 U6583 ( .A1(n5124), .A2(n9535), .ZN(n5127) );
  INV_X1 U6584 ( .A(n5127), .ZN(n5125) );
  NAND2_X1 U6585 ( .A1(n5125), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5128) );
  NAND2_X1 U6586 ( .A1(n5127), .A2(n5126), .ZN(n5143) );
  AOI22_X1 U6587 ( .A1(n4977), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5982), .B2(
        n6954), .ZN(n5129) );
  NAND2_X1 U6588 ( .A1(n4942), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U6589 ( .A1(n5340), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5136) );
  NAND2_X1 U6590 ( .A1(n5132), .A2(n5131), .ZN(n5133) );
  AND2_X1 U6591 ( .A1(n5149), .A2(n5133), .ZN(n9378) );
  NAND2_X1 U6592 ( .A1(n5277), .A2(n9378), .ZN(n5135) );
  NAND2_X1 U6593 ( .A1(n4955), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5134) );
  NAND4_X1 U6594 ( .A1(n5137), .A2(n5136), .A3(n5135), .A4(n5134), .ZN(n9061)
         );
  INV_X1 U6595 ( .A(n9061), .ZN(n9390) );
  OR2_X1 U6596 ( .A1(n9499), .A2(n9390), .ZN(n5535) );
  OR2_X1 U6597 ( .A1(n9589), .A2(n9506), .ZN(n5537) );
  NAND2_X1 U6598 ( .A1(n5537), .A2(n9385), .ZN(n5138) );
  NAND2_X1 U6599 ( .A1(n5138), .A2(n5536), .ZN(n9096) );
  OAI211_X1 U6600 ( .C1(n5157), .C2(n5139), .A(n5535), .B(n9096), .ZN(n5155)
         );
  NAND2_X1 U6601 ( .A1(n9499), .A2(n9390), .ZN(n9097) );
  MUX2_X1 U6602 ( .A(n6074), .B(n6075), .S(n6445), .Z(n5161) );
  XNOR2_X1 U6603 ( .A(n5161), .B(SI_14_), .ZN(n5160) );
  XNOR2_X1 U6604 ( .A(n5165), .B(n5160), .ZN(n7725) );
  NAND2_X1 U6605 ( .A1(n7725), .A2(n4960), .ZN(n5146) );
  NAND2_X1 U6606 ( .A1(n5143), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5144) );
  XNOR2_X1 U6607 ( .A(n5144), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7278) );
  AOI22_X1 U6608 ( .A1(n4977), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5982), .B2(
        n7278), .ZN(n5145) );
  NAND2_X1 U6609 ( .A1(n5146), .A2(n5145), .ZN(n9495) );
  NAND2_X1 U6610 ( .A1(n4955), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U6611 ( .A1(n5482), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5153) );
  INV_X1 U6612 ( .A(n5149), .ZN(n5147) );
  NAND2_X1 U6613 ( .A1(n5147), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5177) );
  INV_X1 U6614 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U6615 ( .A1(n5149), .A2(n5148), .ZN(n5150) );
  AND2_X1 U6616 ( .A1(n5177), .A2(n5150), .ZN(n9358) );
  NAND2_X1 U6617 ( .A1(n4969), .A2(n9358), .ZN(n5152) );
  NAND2_X1 U6618 ( .A1(n5340), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5151) );
  NAND2_X1 U6619 ( .A1(n9495), .A2(n9373), .ZN(n5558) );
  NAND3_X1 U6620 ( .A1(n5155), .A2(n9097), .A3(n5558), .ZN(n5156) );
  OR2_X1 U6621 ( .A1(n9495), .A2(n9373), .ZN(n9098) );
  AND2_X1 U6622 ( .A1(n5536), .A2(n9387), .ZN(n9095) );
  AOI21_X1 U6623 ( .B1(n5158), .B2(n5537), .A(n4573), .ZN(n5159) );
  NAND2_X1 U6624 ( .A1(n9098), .A2(n5535), .ZN(n5577) );
  INV_X1 U6625 ( .A(n5160), .ZN(n5164) );
  INV_X1 U6626 ( .A(n5161), .ZN(n5162) );
  NAND2_X1 U6627 ( .A1(n5162), .A2(SI_14_), .ZN(n5163) );
  MUX2_X1 U6628 ( .A(n6236), .B(n6230), .S(n6445), .Z(n5167) );
  NAND2_X1 U6629 ( .A1(n5167), .A2(n5166), .ZN(n5185) );
  INV_X1 U6630 ( .A(n5167), .ZN(n5168) );
  NAND2_X1 U6631 ( .A1(n5168), .A2(SI_15_), .ZN(n5169) );
  NAND2_X1 U6632 ( .A1(n5185), .A2(n5169), .ZN(n5183) );
  XNOR2_X1 U6633 ( .A(n5184), .B(n5183), .ZN(n7744) );
  NAND2_X1 U6634 ( .A1(n7744), .A2(n4960), .ZN(n5176) );
  NOR2_X1 U6635 ( .A1(n5170), .A2(n9535), .ZN(n5171) );
  MUX2_X1 U6636 ( .A(n9535), .B(n5171), .S(P1_IR_REG_15__SCAN_IN), .Z(n5172)
         );
  INV_X1 U6637 ( .A(n5172), .ZN(n5174) );
  NAND2_X1 U6638 ( .A1(n5174), .A2(n5173), .ZN(n7497) );
  INV_X1 U6639 ( .A(n7497), .ZN(n7282) );
  AOI22_X1 U6640 ( .A1(n4977), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5982), .B2(
        n7282), .ZN(n5175) );
  NAND2_X1 U6641 ( .A1(n4955), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U6642 ( .A1(n4942), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5181) );
  NAND2_X1 U6643 ( .A1(n5177), .A2(n7276), .ZN(n5178) );
  AND2_X1 U6644 ( .A1(n5195), .A2(n5178), .ZN(n9343) );
  NAND2_X1 U6645 ( .A1(n5277), .A2(n9343), .ZN(n5180) );
  NAND2_X1 U6646 ( .A1(n5340), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5179) );
  NAND4_X1 U6647 ( .A1(n5182), .A2(n5181), .A3(n5180), .A4(n5179), .ZN(n8994)
         );
  NOR2_X1 U6648 ( .A1(n9487), .A2(n8994), .ZN(n9066) );
  NAND2_X1 U6649 ( .A1(n9487), .A2(n8994), .ZN(n9067) );
  MUX2_X1 U6650 ( .A(n6241), .B(n6244), .S(n6445), .Z(n5187) );
  NAND2_X1 U6651 ( .A1(n5187), .A2(n5186), .ZN(n5205) );
  INV_X1 U6652 ( .A(n5187), .ZN(n5188) );
  NAND2_X1 U6653 ( .A1(n5188), .A2(SI_16_), .ZN(n5189) );
  XNOR2_X1 U6654 ( .A(n5204), .B(n5203), .ZN(n7736) );
  NAND2_X1 U6655 ( .A1(n7736), .A2(n4960), .ZN(n5192) );
  NAND2_X1 U6656 ( .A1(n5173), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5190) );
  XNOR2_X1 U6657 ( .A(n5190), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7644) );
  AOI22_X1 U6658 ( .A1(n4977), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5982), .B2(
        n7644), .ZN(n5191) );
  NAND2_X1 U6659 ( .A1(n4955), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U6660 ( .A1(n5482), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5199) );
  INV_X1 U6661 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U6662 ( .A1(n5195), .A2(n5194), .ZN(n5196) );
  AND2_X1 U6663 ( .A1(n5236), .A2(n5196), .ZN(n9326) );
  NAND2_X1 U6664 ( .A1(n5277), .A2(n9326), .ZN(n5198) );
  NAND2_X1 U6665 ( .A1(n5340), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5197) );
  OR2_X1 U6666 ( .A1(n9483), .A2(n9336), .ZN(n5579) );
  NAND2_X1 U6667 ( .A1(n9483), .A2(n9336), .ZN(n9102) );
  NAND2_X1 U6668 ( .A1(n5579), .A2(n9102), .ZN(n9319) );
  INV_X1 U6669 ( .A(n8994), .ZN(n9355) );
  OR2_X1 U6670 ( .A1(n9487), .A2(n9355), .ZN(n9101) );
  INV_X1 U6671 ( .A(n9101), .ZN(n5201) );
  AND2_X1 U6672 ( .A1(n9487), .A2(n9355), .ZN(n9100) );
  MUX2_X1 U6673 ( .A(n5201), .B(n9100), .S(n5511), .Z(n5202) );
  NOR2_X1 U6674 ( .A1(n9319), .A2(n5202), .ZN(n5222) );
  MUX2_X1 U6675 ( .A(n6248), .B(n5207), .S(n6445), .Z(n5226) );
  XNOR2_X1 U6676 ( .A(n5226), .B(SI_17_), .ZN(n5224) );
  XNOR2_X1 U6677 ( .A(n5223), .B(n5224), .ZN(n7764) );
  NAND2_X1 U6678 ( .A1(n7764), .A2(n4960), .ZN(n5215) );
  INV_X1 U6679 ( .A(n5208), .ZN(n5209) );
  NAND2_X1 U6680 ( .A1(n5209), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5212) );
  INV_X1 U6681 ( .A(n5212), .ZN(n5210) );
  NAND2_X1 U6682 ( .A1(n5210), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U6683 ( .A1(n5212), .A2(n5211), .ZN(n5230) );
  AOI22_X1 U6684 ( .A1(n4977), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5982), .B2(
        n9015), .ZN(n5214) );
  NAND2_X1 U6685 ( .A1(n4942), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5219) );
  NAND2_X1 U6686 ( .A1(n4955), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5218) );
  XNOR2_X1 U6687 ( .A(n5236), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n9305) );
  NAND2_X1 U6688 ( .A1(n4969), .A2(n9305), .ZN(n5217) );
  NAND2_X1 U6689 ( .A1(n5340), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5216) );
  NAND4_X1 U6690 ( .A1(n5219), .A2(n5218), .A3(n5217), .A4(n5216), .ZN(n9296)
         );
  AND2_X1 U6691 ( .A1(n9476), .A2(n9068), .ZN(n9103) );
  INV_X1 U6692 ( .A(n9103), .ZN(n5242) );
  OR2_X1 U6693 ( .A1(n9476), .A2(n9068), .ZN(n9292) );
  MUX2_X1 U6694 ( .A(n5579), .B(n9102), .S(n5947), .Z(n5220) );
  NAND2_X1 U6695 ( .A1(n9308), .A2(n5220), .ZN(n5221) );
  INV_X1 U6696 ( .A(n5223), .ZN(n5225) );
  NAND2_X1 U6697 ( .A1(n5225), .A2(n5224), .ZN(n5229) );
  INV_X1 U6698 ( .A(n5226), .ZN(n5227) );
  NAND2_X1 U6699 ( .A1(n5227), .A2(SI_17_), .ZN(n5228) );
  NAND2_X1 U6700 ( .A1(n5229), .A2(n5228), .ZN(n5248) );
  MUX2_X1 U6701 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6445), .Z(n5249) );
  XNOR2_X1 U6702 ( .A(n5249), .B(SI_18_), .ZN(n5246) );
  XNOR2_X1 U6703 ( .A(n5248), .B(n5246), .ZN(n7780) );
  NAND2_X1 U6704 ( .A1(n7780), .A2(n4960), .ZN(n5233) );
  NAND2_X1 U6705 ( .A1(n5230), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5231) );
  XNOR2_X1 U6706 ( .A(n5231), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9026) );
  AOI22_X1 U6707 ( .A1(n4977), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5982), .B2(
        n9026), .ZN(n5232) );
  NAND2_X1 U6708 ( .A1(n5482), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U6709 ( .A1(n4955), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5240) );
  INV_X1 U6710 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7638) );
  INV_X1 U6711 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5234) );
  OAI21_X1 U6712 ( .B1(n5236), .B2(n7638), .A(n5234), .ZN(n5237) );
  NAND2_X1 U6713 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n5235) );
  AND2_X1 U6714 ( .A1(n5237), .A2(n5258), .ZN(n9289) );
  NAND2_X1 U6715 ( .A1(n5277), .A2(n9289), .ZN(n5239) );
  NAND2_X1 U6716 ( .A1(n5340), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U6717 ( .A1(n9471), .A2(n9275), .ZN(n9104) );
  NAND2_X1 U6718 ( .A1(n9104), .A2(n5242), .ZN(n5243) );
  OR2_X1 U6719 ( .A1(n9471), .A2(n9275), .ZN(n5525) );
  NAND2_X1 U6720 ( .A1(n5525), .A2(n9292), .ZN(n9105) );
  MUX2_X1 U6721 ( .A(n5243), .B(n9105), .S(n5947), .Z(n5244) );
  OR2_X1 U6722 ( .A1(n5245), .A2(n5244), .ZN(n5283) );
  INV_X1 U6723 ( .A(n5246), .ZN(n5247) );
  NAND2_X1 U6724 ( .A1(n5249), .A2(SI_18_), .ZN(n5250) );
  MUX2_X1 U6725 ( .A(n6380), .B(n6381), .S(n6445), .Z(n5252) );
  INV_X1 U6726 ( .A(SI_19_), .ZN(n5251) );
  NAND2_X1 U6727 ( .A1(n5252), .A2(n5251), .ZN(n5266) );
  INV_X1 U6728 ( .A(n5252), .ZN(n5253) );
  NAND2_X1 U6729 ( .A1(n5253), .A2(SI_19_), .ZN(n5254) );
  NAND2_X1 U6730 ( .A1(n5266), .A2(n5254), .ZN(n5264) );
  XNOR2_X1 U6731 ( .A(n5265), .B(n5264), .ZN(n7793) );
  NAND2_X1 U6732 ( .A1(n7793), .A2(n4960), .ZN(n5256) );
  AOI22_X1 U6733 ( .A1(n4977), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5982), .B2(
        n9207), .ZN(n5255) );
  NAND2_X1 U6734 ( .A1(n4955), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5263) );
  NAND2_X1 U6735 ( .A1(n5482), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U6736 ( .A1(n5257), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5275) );
  INV_X1 U6737 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8859) );
  NAND2_X1 U6738 ( .A1(n5258), .A2(n8859), .ZN(n5259) );
  AND2_X1 U6739 ( .A1(n5275), .A2(n5259), .ZN(n9279) );
  NAND2_X1 U6740 ( .A1(n5277), .A2(n9279), .ZN(n5261) );
  NAND2_X1 U6741 ( .A1(n5340), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5260) );
  NAND4_X1 U6742 ( .A1(n5263), .A2(n5262), .A3(n5261), .A4(n5260), .ZN(n9297)
         );
  NAND2_X1 U6743 ( .A1(n9468), .A2(n9263), .ZN(n9106) );
  AND2_X1 U6744 ( .A1(n9106), .A2(n9104), .ZN(n5553) );
  NAND2_X1 U6745 ( .A1(n5283), .A2(n5553), .ZN(n5282) );
  MUX2_X1 U6746 ( .A(n7809), .B(n6758), .S(n6445), .Z(n5268) );
  INV_X1 U6747 ( .A(SI_20_), .ZN(n5267) );
  NAND2_X1 U6748 ( .A1(n5268), .A2(n5267), .ZN(n5289) );
  INV_X1 U6749 ( .A(n5268), .ZN(n5269) );
  NAND2_X1 U6750 ( .A1(n5269), .A2(SI_20_), .ZN(n5270) );
  XNOR2_X1 U6751 ( .A(n5288), .B(n5287), .ZN(n7808) );
  NAND2_X1 U6752 ( .A1(n7808), .A2(n4960), .ZN(n5272) );
  NAND2_X1 U6753 ( .A1(n4977), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6754 ( .A1(n5482), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6755 ( .A1(n5340), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5280) );
  INV_X1 U6756 ( .A(n5275), .ZN(n5273) );
  NAND2_X1 U6757 ( .A1(n5273), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5294) );
  INV_X1 U6758 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5274) );
  NAND2_X1 U6759 ( .A1(n5275), .A2(n5274), .ZN(n5276) );
  AND2_X1 U6760 ( .A1(n5294), .A2(n5276), .ZN(n9264) );
  NAND2_X1 U6761 ( .A1(n5277), .A2(n9264), .ZN(n5279) );
  NAND2_X1 U6762 ( .A1(n4955), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5278) );
  NAND4_X1 U6763 ( .A1(n5281), .A2(n5280), .A3(n5279), .A4(n5278), .ZN(n9073)
         );
  OR2_X1 U6764 ( .A1(n9463), .A2(n9274), .ZN(n5523) );
  OR2_X1 U6765 ( .A1(n9468), .A2(n9263), .ZN(n5524) );
  AND2_X1 U6766 ( .A1(n5523), .A2(n5524), .ZN(n5554) );
  NAND2_X1 U6767 ( .A1(n5282), .A2(n5554), .ZN(n5286) );
  NAND3_X1 U6768 ( .A1(n5283), .A2(n5525), .A3(n5524), .ZN(n5284) );
  NAND2_X1 U6769 ( .A1(n9463), .A2(n9274), .ZN(n9107) );
  NAND3_X1 U6770 ( .A1(n5284), .A2(n9106), .A3(n9107), .ZN(n5285) );
  INV_X1 U6771 ( .A(n5381), .ZN(n5322) );
  NAND2_X1 U6772 ( .A1(n5288), .A2(n5287), .ZN(n5290) );
  MUX2_X1 U6773 ( .A(n7827), .B(n7706), .S(n6445), .Z(n5303) );
  XNOR2_X1 U6774 ( .A(n5303), .B(SI_21_), .ZN(n5302) );
  XNOR2_X1 U6775 ( .A(n5307), .B(n5302), .ZN(n7826) );
  NAND2_X1 U6776 ( .A1(n7826), .A2(n4960), .ZN(n5292) );
  NAND2_X1 U6777 ( .A1(n4977), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6778 ( .A1(n5482), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U6779 ( .A1(n5340), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5298) );
  INV_X1 U6780 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6781 ( .A1(n5294), .A2(n5293), .ZN(n5295) );
  AND2_X1 U6782 ( .A1(n5315), .A2(n5295), .ZN(n9243) );
  NAND2_X1 U6783 ( .A1(n5277), .A2(n9243), .ZN(n5297) );
  NAND2_X1 U6784 ( .A1(n4955), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5296) );
  INV_X1 U6785 ( .A(n9107), .ZN(n5300) );
  NAND2_X1 U6786 ( .A1(n9108), .A2(n5300), .ZN(n5301) );
  NAND2_X1 U6787 ( .A1(n9458), .A2(n9262), .ZN(n5522) );
  AND2_X1 U6788 ( .A1(n5301), .A2(n5522), .ZN(n5321) );
  INV_X1 U6789 ( .A(n5302), .ZN(n5306) );
  INV_X1 U6790 ( .A(n5303), .ZN(n5304) );
  NAND2_X1 U6791 ( .A1(n5304), .A2(SI_21_), .ZN(n5305) );
  MUX2_X1 U6792 ( .A(n7840), .B(n7057), .S(n6445), .Z(n5309) );
  NAND2_X1 U6793 ( .A1(n5309), .A2(n5308), .ZN(n5325) );
  INV_X1 U6794 ( .A(n5309), .ZN(n5310) );
  NAND2_X1 U6795 ( .A1(n5310), .A2(SI_22_), .ZN(n5311) );
  NAND2_X1 U6796 ( .A1(n5325), .A2(n5311), .ZN(n5323) );
  XNOR2_X1 U6797 ( .A(n5324), .B(n5323), .ZN(n7839) );
  NAND2_X1 U6798 ( .A1(n7839), .A2(n4960), .ZN(n5313) );
  NAND2_X1 U6799 ( .A1(n4977), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5312) );
  NAND2_X1 U6800 ( .A1(n5482), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6801 ( .A1(n4955), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5319) );
  INV_X1 U6802 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6803 ( .A1(n5315), .A2(n5314), .ZN(n5316) );
  AND2_X1 U6804 ( .A1(n5351), .A2(n5316), .ZN(n9230) );
  NAND2_X1 U6805 ( .A1(n4969), .A2(n9230), .ZN(n5318) );
  NAND2_X1 U6806 ( .A1(n5340), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5317) );
  NAND4_X1 U6807 ( .A1(n5320), .A2(n5319), .A3(n5318), .A4(n5317), .ZN(n9075)
         );
  NAND2_X1 U6808 ( .A1(n9450), .A2(n9248), .ZN(n9110) );
  NAND2_X1 U6809 ( .A1(n5321), .A2(n9110), .ZN(n5635) );
  AOI21_X1 U6810 ( .B1(n5322), .B2(n9108), .A(n5635), .ZN(n5359) );
  OR2_X1 U6811 ( .A1(n9450), .A2(n9248), .ZN(n9213) );
  INV_X1 U6812 ( .A(n9213), .ZN(n5358) );
  INV_X1 U6813 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5326) );
  MUX2_X1 U6814 ( .A(n7853), .B(n5326), .S(n6445), .Z(n5327) );
  INV_X1 U6815 ( .A(SI_23_), .ZN(n6170) );
  NAND2_X1 U6816 ( .A1(n5327), .A2(n6170), .ZN(n5330) );
  INV_X1 U6817 ( .A(n5327), .ZN(n5328) );
  NAND2_X1 U6818 ( .A1(n5328), .A2(SI_23_), .ZN(n5329) );
  NAND2_X1 U6819 ( .A1(n5345), .A2(n5344), .ZN(n5331) );
  MUX2_X1 U6820 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n6445), .Z(n5362) );
  INV_X1 U6821 ( .A(SI_24_), .ZN(n6152) );
  XNOR2_X1 U6822 ( .A(n5362), .B(n6152), .ZN(n5361) );
  XNOR2_X1 U6823 ( .A(n5360), .B(n5361), .ZN(n7865) );
  NAND2_X1 U6824 ( .A1(n7865), .A2(n4960), .ZN(n5333) );
  NAND2_X1 U6825 ( .A1(n4977), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5332) );
  INV_X1 U6826 ( .A(n5351), .ZN(n5334) );
  NAND2_X1 U6827 ( .A1(n5334), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5353) );
  INV_X1 U6828 ( .A(n5353), .ZN(n5335) );
  NAND2_X1 U6829 ( .A1(n5335), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5371) );
  INV_X1 U6830 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U6831 ( .A1(n5353), .A2(n5336), .ZN(n5337) );
  NAND2_X1 U6832 ( .A1(n5371), .A2(n5337), .ZN(n9206) );
  OR2_X1 U6833 ( .A1(n9206), .A2(n5459), .ZN(n5343) );
  NAND2_X1 U6834 ( .A1(n5482), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6835 ( .A1(n4955), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5338) );
  AND2_X1 U6836 ( .A1(n5339), .A2(n5338), .ZN(n5342) );
  NAND2_X1 U6837 ( .A1(n5340), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U6838 ( .A1(n9442), .A2(n9218), .ZN(n9113) );
  XNOR2_X1 U6839 ( .A(n5345), .B(n5344), .ZN(n7852) );
  NAND2_X1 U6840 ( .A1(n7852), .A2(n4960), .ZN(n5347) );
  NAND2_X1 U6841 ( .A1(n4977), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5346) );
  INV_X1 U6842 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U6843 ( .A1(n5482), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5348) );
  OAI21_X1 U6844 ( .B1(n5349), .B2(n5481), .A(n5348), .ZN(n5357) );
  INV_X1 U6845 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U6846 ( .A1(n5351), .A2(n5350), .ZN(n5352) );
  NAND2_X1 U6847 ( .A1(n5353), .A2(n5352), .ZN(n8847) );
  INV_X1 U6848 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5354) );
  OAI22_X1 U6849 ( .A1(n8847), .A2(n5459), .B1(n5355), .B2(n5354), .ZN(n5356)
         );
  AND2_X1 U6850 ( .A1(n9447), .A2(n9203), .ZN(n9111) );
  INV_X1 U6851 ( .A(n9111), .ZN(n5592) );
  AND2_X1 U6852 ( .A1(n9113), .A2(n5592), .ZN(n5638) );
  OAI21_X1 U6853 ( .B1(n5359), .B2(n5358), .A(n5638), .ZN(n5380) );
  NAND2_X1 U6854 ( .A1(n5362), .A2(SI_24_), .ZN(n5363) );
  INV_X1 U6855 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7881) );
  MUX2_X1 U6856 ( .A(n7881), .B(n7470), .S(n6445), .Z(n5365) );
  INV_X1 U6857 ( .A(SI_25_), .ZN(n5364) );
  NAND2_X1 U6858 ( .A1(n5365), .A2(n5364), .ZN(n5388) );
  INV_X1 U6859 ( .A(n5365), .ZN(n5366) );
  NAND2_X1 U6860 ( .A1(n5366), .A2(SI_25_), .ZN(n5367) );
  NAND2_X1 U6861 ( .A1(n5388), .A2(n5367), .ZN(n5389) );
  XNOR2_X1 U6862 ( .A(n5390), .B(n5389), .ZN(n7880) );
  NAND2_X1 U6863 ( .A1(n7880), .A2(n4960), .ZN(n5369) );
  NAND2_X1 U6864 ( .A1(n4977), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5368) );
  INV_X1 U6865 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6866 ( .A1(n5371), .A2(n5370), .ZN(n5372) );
  AND2_X1 U6867 ( .A1(n5400), .A2(n5372), .ZN(n9187) );
  NAND2_X1 U6868 ( .A1(n9187), .A2(n4969), .ZN(n5375) );
  AOI22_X1 U6869 ( .A1(n4955), .A2(P1_REG1_REG_25__SCAN_IN), .B1(n5482), .B2(
        P1_REG0_REG_25__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6870 ( .A1(n5340), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5373) );
  AND2_X1 U6871 ( .A1(n9173), .A2(n5589), .ZN(n5613) );
  NAND2_X1 U6872 ( .A1(n5589), .A2(n9203), .ZN(n5377) );
  NAND2_X1 U6873 ( .A1(n9113), .A2(n9225), .ZN(n5376) );
  AND2_X1 U6874 ( .A1(n5377), .A2(n5376), .ZN(n5385) );
  INV_X1 U6875 ( .A(n5385), .ZN(n5378) );
  NAND2_X1 U6876 ( .A1(n5378), .A2(n9235), .ZN(n5379) );
  NAND3_X1 U6877 ( .A1(n5380), .A2(n5613), .A3(n5379), .ZN(n5387) );
  INV_X1 U6878 ( .A(n5522), .ZN(n9109) );
  NAND2_X1 U6879 ( .A1(n9225), .A2(n9235), .ZN(n5521) );
  AND2_X1 U6880 ( .A1(n5521), .A2(n9213), .ZN(n9112) );
  NAND2_X1 U6881 ( .A1(n9112), .A2(n9108), .ZN(n5383) );
  INV_X1 U6882 ( .A(n5521), .ZN(n5382) );
  NAND2_X1 U6883 ( .A1(n9435), .A2(n9204), .ZN(n9115) );
  AND2_X1 U6884 ( .A1(n9115), .A2(n9113), .ZN(n5593) );
  OAI211_X1 U6885 ( .C1(n9225), .C2(n5385), .A(n5384), .B(n5593), .ZN(n5386)
         );
  MUX2_X1 U6886 ( .A(n5387), .B(n5386), .S(n5511), .Z(n5436) );
  INV_X1 U6887 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7895) );
  INV_X1 U6888 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5391) );
  MUX2_X1 U6889 ( .A(n7895), .B(n5391), .S(n6445), .Z(n5393) );
  INV_X1 U6890 ( .A(SI_26_), .ZN(n5392) );
  NAND2_X1 U6891 ( .A1(n5393), .A2(n5392), .ZN(n5415) );
  INV_X1 U6892 ( .A(n5393), .ZN(n5394) );
  NAND2_X1 U6893 ( .A1(n5394), .A2(SI_26_), .ZN(n5395) );
  NAND2_X1 U6894 ( .A1(n7894), .A2(n4960), .ZN(n5397) );
  NAND2_X1 U6895 ( .A1(n4977), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5396) );
  OR2_X1 U6896 ( .A1(n9172), .A2(n5947), .ZN(n5434) );
  INV_X1 U6897 ( .A(n5400), .ZN(n5398) );
  NAND2_X1 U6898 ( .A1(n5398), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5424) );
  INV_X1 U6899 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U6900 ( .A1(n5400), .A2(n5399), .ZN(n5401) );
  NAND2_X1 U6901 ( .A1(n5424), .A2(n5401), .ZN(n8972) );
  INV_X1 U6902 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U6903 ( .A1(n5340), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U6904 ( .A1(n5482), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5402) );
  OAI211_X1 U6905 ( .C1(n5481), .C2(n5404), .A(n5403), .B(n5402), .ZN(n5405)
         );
  INV_X1 U6906 ( .A(n5405), .ZN(n5406) );
  NAND2_X1 U6907 ( .A1(n5434), .A2(n9158), .ZN(n5412) );
  INV_X1 U6908 ( .A(n9173), .ZN(n5433) );
  AOI21_X1 U6909 ( .B1(n9172), .B2(n5433), .A(n9193), .ZN(n5410) );
  NAND2_X1 U6910 ( .A1(n9172), .A2(n9115), .ZN(n5408) );
  NAND2_X1 U6911 ( .A1(n5408), .A2(n5641), .ZN(n5409) );
  MUX2_X1 U6912 ( .A(n5410), .B(n5409), .S(n5947), .Z(n5411) );
  OAI21_X1 U6913 ( .B1(n5436), .B2(n5412), .A(n5411), .ZN(n5438) );
  INV_X1 U6914 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8829) );
  INV_X1 U6915 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5417) );
  MUX2_X1 U6916 ( .A(n8829), .B(n5417), .S(n6445), .Z(n5419) );
  INV_X1 U6917 ( .A(SI_27_), .ZN(n5418) );
  NAND2_X1 U6918 ( .A1(n5419), .A2(n5418), .ZN(n5441) );
  INV_X1 U6919 ( .A(n5419), .ZN(n5420) );
  NAND2_X1 U6920 ( .A1(n5420), .A2(SI_27_), .ZN(n5421) );
  NAND2_X1 U6921 ( .A1(n8827), .A2(n4960), .ZN(n5423) );
  NAND2_X1 U6922 ( .A1(n4977), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5422) );
  INV_X1 U6923 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U6924 ( .A1(n5424), .A2(n5943), .ZN(n5425) );
  NAND2_X1 U6925 ( .A1(n9162), .A2(n5277), .ZN(n5431) );
  INV_X1 U6926 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U6927 ( .A1(n5482), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U6928 ( .A1(n5340), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5426) );
  OAI211_X1 U6929 ( .C1(n5481), .C2(n5428), .A(n5427), .B(n5426), .ZN(n5429)
         );
  INV_X1 U6930 ( .A(n5429), .ZN(n5430) );
  NAND2_X1 U6931 ( .A1(n9427), .A2(n9143), .ZN(n5552) );
  NAND2_X1 U6932 ( .A1(n9140), .A2(n5552), .ZN(n9086) );
  NAND3_X1 U6933 ( .A1(n9115), .A2(n9193), .A3(n5947), .ZN(n5432) );
  OAI21_X1 U6934 ( .B1(n5434), .B2(n5433), .A(n5432), .ZN(n5435) );
  NAND2_X1 U6935 ( .A1(n5436), .A2(n5435), .ZN(n5437) );
  NAND3_X1 U6936 ( .A1(n5438), .A2(n9154), .A3(n5437), .ZN(n5456) );
  INV_X1 U6937 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7969) );
  INV_X1 U6938 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5442) );
  MUX2_X1 U6939 ( .A(n7969), .B(n5442), .S(n6445), .Z(n5468) );
  XNOR2_X1 U6940 ( .A(n5468), .B(SI_28_), .ZN(n5465) );
  NAND2_X1 U6941 ( .A1(n7968), .A2(n4960), .ZN(n5444) );
  NAND2_X1 U6942 ( .A1(n4977), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5443) );
  INV_X1 U6943 ( .A(n5447), .ZN(n5445) );
  NAND2_X1 U6944 ( .A1(n5445), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9126) );
  INV_X1 U6945 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5446) );
  NAND2_X1 U6946 ( .A1(n5447), .A2(n5446), .ZN(n5448) );
  NAND2_X1 U6947 ( .A1(n9126), .A2(n5448), .ZN(n7694) );
  INV_X1 U6948 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5451) );
  NAND2_X1 U6949 ( .A1(n5340), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U6950 ( .A1(n5482), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5449) );
  OAI211_X1 U6951 ( .C1(n5481), .C2(n5451), .A(n5450), .B(n5449), .ZN(n5452)
         );
  INV_X1 U6952 ( .A(n5452), .ZN(n5453) );
  NAND2_X1 U6953 ( .A1(n9423), .A2(n9089), .ZN(n9118) );
  MUX2_X1 U6954 ( .A(n9140), .B(n5552), .S(n5947), .Z(n5455) );
  NAND3_X1 U6955 ( .A1(n5456), .A2(n9139), .A3(n5455), .ZN(n5458) );
  MUX2_X1 U6956 ( .A(n9118), .B(n5548), .S(n5947), .Z(n5457) );
  OR2_X1 U6957 ( .A1(n9126), .A2(n5459), .ZN(n5464) );
  INV_X1 U6958 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U6959 ( .A1(n4955), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U6960 ( .A1(n5340), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5460) );
  OAI211_X1 U6961 ( .C1(n5026), .C2(n6141), .A(n5461), .B(n5460), .ZN(n5462)
         );
  INV_X1 U6962 ( .A(n5462), .ZN(n5463) );
  INV_X1 U6963 ( .A(SI_28_), .ZN(n5467) );
  NAND2_X1 U6964 ( .A1(n5468), .A2(n5467), .ZN(n5469) );
  INV_X1 U6965 ( .A(SI_29_), .ZN(n5498) );
  MUX2_X1 U6966 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6445), .Z(n5499) );
  INV_X1 U6967 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8102) );
  INV_X1 U6968 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n5471) );
  MUX2_X1 U6969 ( .A(n8102), .B(n5471), .S(n6445), .Z(n5473) );
  INV_X1 U6970 ( .A(SI_30_), .ZN(n5472) );
  NAND2_X1 U6971 ( .A1(n5473), .A2(n5472), .ZN(n5488) );
  INV_X1 U6972 ( .A(n5473), .ZN(n5474) );
  NAND2_X1 U6973 ( .A1(n5474), .A2(SI_30_), .ZN(n5475) );
  NAND2_X1 U6974 ( .A1(n5488), .A2(n5475), .ZN(n5489) );
  XNOR2_X1 U6975 ( .A(n5490), .B(n5489), .ZN(n8101) );
  NAND2_X1 U6976 ( .A1(n8101), .A2(n4960), .ZN(n5477) );
  NAND2_X1 U6977 ( .A1(n4977), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5476) );
  INV_X1 U6978 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U6979 ( .A1(n5340), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U6980 ( .A1(n5482), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5478) );
  OAI211_X1 U6981 ( .C1(n5481), .C2(n5480), .A(n5479), .B(n5478), .ZN(n9121)
         );
  INV_X1 U6982 ( .A(n9121), .ZN(n5495) );
  NAND2_X1 U6983 ( .A1(n9410), .A2(n5495), .ZN(n5648) );
  NAND2_X1 U6984 ( .A1(n4955), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U6985 ( .A1(n4954), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U6986 ( .A1(n5482), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5483) );
  NAND3_X1 U6987 ( .A1(n5485), .A2(n5484), .A3(n5483), .ZN(n9045) );
  INV_X1 U6988 ( .A(n9045), .ZN(n5486) );
  NAND2_X1 U6989 ( .A1(n9410), .A2(n5486), .ZN(n5487) );
  AND2_X1 U6990 ( .A1(n5648), .A2(n5487), .ZN(n5506) );
  INV_X1 U6991 ( .A(n5506), .ZN(n5597) );
  INV_X1 U6992 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8822) );
  INV_X1 U6993 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5491) );
  MUX2_X1 U6994 ( .A(n8822), .B(n5491), .S(n6445), .Z(n5492) );
  XNOR2_X1 U6995 ( .A(n5492), .B(SI_31_), .ZN(n5493) );
  OR2_X1 U6996 ( .A1(n9410), .A2(n5495), .ZN(n5496) );
  NAND2_X1 U6997 ( .A1(n5610), .A2(n4651), .ZN(n5547) );
  XNOR2_X1 U6998 ( .A(n5499), .B(n5498), .ZN(n5500) );
  NAND2_X1 U6999 ( .A1(n8097), .A2(n4960), .ZN(n5502) );
  NAND2_X1 U7000 ( .A1(n4977), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5501) );
  NAND3_X1 U7001 ( .A1(n5503), .A2(n9417), .A3(n5547), .ZN(n5507) );
  INV_X1 U7002 ( .A(n5504), .ZN(n5505) );
  AOI21_X1 U7003 ( .B1(n5507), .B2(n5506), .A(n5505), .ZN(n5508) );
  NAND3_X1 U7004 ( .A1(n5510), .A2(n9129), .A3(n9144), .ZN(n5514) );
  INV_X1 U7005 ( .A(n9144), .ZN(n8993) );
  MUX2_X1 U7006 ( .A(n8993), .B(n9417), .S(n5511), .Z(n5512) );
  NOR2_X1 U7007 ( .A1(n5597), .A2(n5512), .ZN(n5513) );
  NAND3_X1 U7008 ( .A1(n5514), .A2(n5513), .A3(n5547), .ZN(n5515) );
  NAND2_X1 U7009 ( .A1(n9046), .A2(n9045), .ZN(n5605) );
  NAND2_X1 U7010 ( .A1(n5515), .A2(n5605), .ZN(n5516) );
  INV_X1 U7011 ( .A(n6292), .ZN(n6717) );
  INV_X1 U7012 ( .A(n5605), .ZN(n5651) );
  INV_X1 U7013 ( .A(n5648), .ZN(n5545) );
  NOR2_X1 U7014 ( .A1(n9417), .A2(n9144), .ZN(n5550) );
  INV_X1 U7015 ( .A(n9116), .ZN(n5520) );
  NAND2_X1 U7016 ( .A1(n5520), .A2(n5641), .ZN(n9175) );
  NAND2_X1 U7017 ( .A1(n9173), .A2(n9115), .ZN(n9190) );
  NAND2_X1 U7018 ( .A1(n5589), .A2(n9113), .ZN(n9200) );
  NAND2_X1 U7019 ( .A1(n5592), .A2(n5521), .ZN(n9216) );
  NAND2_X1 U7020 ( .A1(n9213), .A2(n9110), .ZN(n9232) );
  NAND2_X1 U7021 ( .A1(n9108), .A2(n5522), .ZN(n9251) );
  NAND2_X1 U7022 ( .A1(n5523), .A2(n9107), .ZN(n9259) );
  NAND2_X1 U7023 ( .A1(n5525), .A2(n9104), .ZN(n9286) );
  INV_X1 U7024 ( .A(n9286), .ZN(n9294) );
  INV_X1 U7025 ( .A(n9308), .ZN(n9302) );
  NAND2_X1 U7026 ( .A1(n5622), .A2(n5526), .ZN(n6964) );
  INV_X1 U7027 ( .A(n6964), .ZN(n6966) );
  AND2_X1 U7028 ( .A1(n5674), .A2(n6704), .ZN(n5614) );
  NOR2_X1 U7029 ( .A1(n6858), .A2(n5614), .ZN(n6291) );
  NAND2_X1 U7030 ( .A1(n5564), .A2(n5527), .ZN(n7041) );
  INV_X1 U7031 ( .A(n7041), .ZN(n5528) );
  NAND4_X1 U7032 ( .A1(n6966), .A2(n6291), .A3(n5528), .A4(n7000), .ZN(n5531)
         );
  INV_X1 U7033 ( .A(n5529), .ZN(n6859) );
  INV_X1 U7034 ( .A(n5624), .ZN(n5530) );
  NOR4_X1 U7035 ( .A1(n5531), .A2(n6859), .A3(n5530), .A4(n6701), .ZN(n5532)
         );
  NAND4_X1 U7036 ( .A1(n5532), .A2(n5569), .A3(n7607), .A4(n7609), .ZN(n5534)
         );
  INV_X1 U7037 ( .A(n9579), .ZN(n9587) );
  NAND2_X1 U7038 ( .A1(n4295), .A2(n7612), .ZN(n9633) );
  NAND2_X1 U7039 ( .A1(n5533), .A2(n9093), .ZN(n9052) );
  NOR4_X1 U7040 ( .A1(n5534), .A2(n9587), .A3(n9633), .A4(n9052), .ZN(n5538)
         );
  NAND2_X1 U7041 ( .A1(n5535), .A2(n9097), .ZN(n9368) );
  INV_X1 U7042 ( .A(n9368), .ZN(n9366) );
  NAND2_X1 U7043 ( .A1(n5537), .A2(n5536), .ZN(n9392) );
  INV_X1 U7044 ( .A(n9392), .ZN(n9388) );
  NAND4_X1 U7045 ( .A1(n5538), .A2(n9352), .A3(n9366), .A4(n9388), .ZN(n5539)
         );
  NOR4_X1 U7046 ( .A1(n9302), .A2(n5539), .A3(n4367), .A4(n9319), .ZN(n5540)
         );
  NAND4_X1 U7047 ( .A1(n4586), .A2(n9272), .A3(n9294), .A4(n5540), .ZN(n5541)
         );
  OR4_X1 U7048 ( .A1(n9216), .A2(n9232), .A3(n9251), .A4(n5541), .ZN(n5542) );
  NOR4_X1 U7049 ( .A1(n9175), .A2(n9190), .A3(n9200), .A4(n5542), .ZN(n5543)
         );
  NAND4_X1 U7050 ( .A1(n9120), .A2(n9154), .A3(n9139), .A4(n5543), .ZN(n5544)
         );
  NOR4_X1 U7051 ( .A1(n5610), .A2(n5651), .A3(n5545), .A4(n5544), .ZN(n5546)
         );
  NOR2_X1 U7052 ( .A1(n5546), .A2(n6284), .ZN(n5601) );
  INV_X1 U7053 ( .A(n5547), .ZN(n5600) );
  INV_X1 U7054 ( .A(n5548), .ZN(n5549) );
  NOR2_X1 U7055 ( .A1(n5550), .A2(n5549), .ZN(n5611) );
  NAND2_X1 U7056 ( .A1(n9140), .A2(n9116), .ZN(n5551) );
  AND3_X1 U7057 ( .A1(n9118), .A2(n5552), .A3(n5551), .ZN(n5612) );
  INV_X1 U7058 ( .A(n5553), .ZN(n5555) );
  OAI211_X1 U7059 ( .C1(n4593), .C2(n5555), .A(n9108), .B(n5554), .ZN(n5634)
         );
  INV_X1 U7060 ( .A(n9102), .ZN(n5556) );
  NOR2_X1 U7061 ( .A1(n9103), .A2(n5556), .ZN(n5557) );
  NAND2_X1 U7062 ( .A1(n9104), .A2(n5557), .ZN(n5584) );
  OAI211_X1 U7063 ( .C1(n7610), .C2(n7616), .A(n9095), .B(n9097), .ZN(n5576)
         );
  OR2_X1 U7064 ( .A1(n9100), .A2(n4371), .ZN(n5581) );
  OR4_X1 U7065 ( .A1(n5584), .A2(n5576), .A3(n5581), .A4(n4571), .ZN(n5631) );
  NAND2_X1 U7066 ( .A1(n5560), .A2(n5559), .ZN(n7039) );
  INV_X1 U7067 ( .A(n5561), .ZN(n5562) );
  NAND2_X1 U7068 ( .A1(n5562), .A2(n5624), .ZN(n5563) );
  AND2_X1 U7069 ( .A1(n5563), .A2(n5569), .ZN(n5625) );
  NAND3_X1 U7070 ( .A1(n7039), .A2(n5625), .A3(n5620), .ZN(n5572) );
  NAND2_X1 U7071 ( .A1(n5622), .A2(n5564), .ZN(n5567) );
  INV_X1 U7072 ( .A(n5565), .ZN(n5566) );
  NAND2_X1 U7073 ( .A1(n5567), .A2(n5566), .ZN(n5568) );
  NAND3_X1 U7074 ( .A1(n5568), .A2(n5624), .A3(n5623), .ZN(n5570) );
  NAND2_X1 U7075 ( .A1(n5570), .A2(n5569), .ZN(n5571) );
  NAND2_X1 U7076 ( .A1(n5572), .A2(n5571), .ZN(n5585) );
  INV_X1 U7077 ( .A(n5573), .ZN(n5574) );
  NOR2_X1 U7078 ( .A1(n5574), .A2(n7616), .ZN(n5575) );
  OAI22_X1 U7079 ( .A1(n5576), .A2(n5575), .B1(n4573), .B2(n9096), .ZN(n5578)
         );
  NOR2_X1 U7080 ( .A1(n5578), .A2(n5577), .ZN(n5580) );
  OAI211_X1 U7081 ( .C1(n5581), .C2(n5580), .A(n9101), .B(n5579), .ZN(n5582)
         );
  INV_X1 U7082 ( .A(n5582), .ZN(n5583) );
  OR2_X1 U7083 ( .A1(n5584), .A2(n5583), .ZN(n5629) );
  OAI21_X1 U7084 ( .B1(n5631), .B2(n5585), .A(n5629), .ZN(n5586) );
  AND2_X1 U7085 ( .A1(n5586), .A2(n9106), .ZN(n5587) );
  NOR2_X1 U7086 ( .A1(n5634), .A2(n5587), .ZN(n5588) );
  OAI21_X1 U7087 ( .B1(n5588), .B2(n5635), .A(n9112), .ZN(n5591) );
  INV_X1 U7088 ( .A(n5589), .ZN(n5590) );
  AOI21_X1 U7089 ( .B1(n5592), .B2(n5591), .A(n5590), .ZN(n5595) );
  INV_X1 U7090 ( .A(n5593), .ZN(n5594) );
  AND2_X1 U7091 ( .A1(n5641), .A2(n9173), .ZN(n9117) );
  OAI211_X1 U7092 ( .C1(n5595), .C2(n5594), .A(n9140), .B(n9117), .ZN(n5596)
         );
  NAND2_X1 U7093 ( .A1(n5612), .A2(n5596), .ZN(n5598) );
  AOI211_X1 U7094 ( .C1(n5611), .C2(n5598), .A(n5646), .B(n5597), .ZN(n5599)
         );
  OAI211_X1 U7095 ( .C1(n5600), .C2(n5599), .A(n6284), .B(n5605), .ZN(n5603)
         );
  INV_X1 U7096 ( .A(n5601), .ZN(n5602) );
  NAND2_X1 U7097 ( .A1(n5603), .A2(n5602), .ZN(n5604) );
  NAND3_X1 U7098 ( .A1(n5605), .A2(n6284), .A3(n5678), .ZN(n5607) );
  XNOR2_X2 U7099 ( .A(n5606), .B(P1_IR_REG_20__SCAN_IN), .ZN(n6707) );
  OAI21_X1 U7100 ( .B1(n5608), .B2(n5607), .A(n6707), .ZN(n5609) );
  INV_X1 U7101 ( .A(n5610), .ZN(n5653) );
  INV_X1 U7102 ( .A(n5611), .ZN(n5650) );
  INV_X1 U7103 ( .A(n5612), .ZN(n5645) );
  INV_X1 U7104 ( .A(n5613), .ZN(n5640) );
  AOI21_X1 U7105 ( .B1(n9005), .B2(n9664), .A(n5670), .ZN(n5616) );
  INV_X1 U7106 ( .A(n5614), .ZN(n5615) );
  AND2_X1 U7107 ( .A1(n5616), .A2(n5615), .ZN(n5617) );
  OAI22_X1 U7108 ( .A1(n6711), .A2(n5617), .B1(n7043), .B2(n8948), .ZN(n5619)
         );
  NAND2_X1 U7109 ( .A1(n5619), .A2(n5618), .ZN(n5621) );
  NAND2_X1 U7110 ( .A1(n5621), .A2(n5620), .ZN(n5628) );
  AND3_X1 U7111 ( .A1(n5624), .A2(n5623), .A3(n5622), .ZN(n5627) );
  INV_X1 U7112 ( .A(n5625), .ZN(n5626) );
  AOI21_X1 U7113 ( .B1(n5628), .B2(n5627), .A(n5626), .ZN(n5630) );
  OAI21_X1 U7114 ( .B1(n5631), .B2(n5630), .A(n5629), .ZN(n5632) );
  AND2_X1 U7115 ( .A1(n5632), .A2(n9106), .ZN(n5633) );
  NOR2_X1 U7116 ( .A1(n5634), .A2(n5633), .ZN(n5636) );
  OAI21_X1 U7117 ( .B1(n5636), .B2(n5635), .A(n9112), .ZN(n5637) );
  AND2_X1 U7118 ( .A1(n5638), .A2(n5637), .ZN(n5639) );
  OAI21_X1 U7119 ( .B1(n5640), .B2(n5639), .A(n9115), .ZN(n5642) );
  NAND2_X1 U7120 ( .A1(n5642), .A2(n5641), .ZN(n5643) );
  NOR2_X1 U7121 ( .A1(n9086), .A2(n5643), .ZN(n5644) );
  NOR2_X1 U7122 ( .A1(n5645), .A2(n5644), .ZN(n5649) );
  INV_X1 U7123 ( .A(n5646), .ZN(n5647) );
  OAI211_X1 U7124 ( .C1(n5650), .C2(n5649), .A(n5648), .B(n5647), .ZN(n5652)
         );
  AOI21_X1 U7125 ( .B1(n5653), .B2(n5652), .A(n5651), .ZN(n5654) );
  NAND2_X1 U7126 ( .A1(n4339), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5656) );
  OR2_X1 U7127 ( .A1(n5953), .A2(P1_U3084), .ZN(n7151) );
  NOR2_X1 U7128 ( .A1(n7003), .A2(n6356), .ZN(n5941) );
  NAND2_X1 U7129 ( .A1(n5662), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U7130 ( .A1(n4305), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5665) );
  AND2_X1 U7131 ( .A1(n5953), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5666) );
  INV_X1 U7132 ( .A(n5667), .ZN(n9043) );
  NAND3_X1 U7133 ( .A1(n5941), .A2(n9654), .A3(n9043), .ZN(n5668) );
  OAI211_X1 U7134 ( .C1(n6712), .C2(n7151), .A(n5668), .B(P1_B_REG_SCAN_IN), 
        .ZN(n5669) );
  NAND2_X1 U7135 ( .A1(n5678), .A2(n5934), .ZN(n5671) );
  AND2_X4 U7136 ( .A1(n4262), .A2(n5671), .ZN(n5710) );
  AOI22_X1 U7137 ( .A1(n9447), .A2(n7689), .B1(n5710), .B2(n9235), .ZN(n8845)
         );
  AOI22_X1 U7138 ( .A1(n5699), .A2(n6883), .B1(n5675), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5672) );
  INV_X1 U7139 ( .A(n5672), .ZN(n5673) );
  NAND2_X1 U7140 ( .A1(n5674), .A2(n5699), .ZN(n5677) );
  AOI22_X1 U7141 ( .A1(n5743), .A2(n6883), .B1(n5675), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U7142 ( .A1(n5677), .A2(n5676), .ZN(n6250) );
  NAND2_X1 U7143 ( .A1(n6252), .A2(n6250), .ZN(n6251) );
  INV_X1 U7144 ( .A(n6250), .ZN(n5680) );
  OR2_X1 U7145 ( .A1(n5678), .A2(n9207), .ZN(n5679) );
  NAND2_X1 U7146 ( .A1(n5680), .A2(n5900), .ZN(n5681) );
  NAND2_X1 U7147 ( .A1(n6251), .A2(n5681), .ZN(n5693) );
  INV_X1 U7148 ( .A(n5693), .ZN(n5688) );
  NAND2_X1 U7149 ( .A1(n5689), .A2(n5699), .ZN(n5685) );
  NAND2_X1 U7150 ( .A1(n5683), .A2(n5743), .ZN(n5684) );
  NAND2_X1 U7151 ( .A1(n5685), .A2(n5684), .ZN(n5686) );
  INV_X2 U7152 ( .A(n5746), .ZN(n5708) );
  XNOR2_X1 U7153 ( .A(n5686), .B(n5708), .ZN(n5692) );
  INV_X1 U7154 ( .A(n5692), .ZN(n5687) );
  NAND2_X1 U7155 ( .A1(n5710), .A2(n5689), .ZN(n5691) );
  NAND2_X1 U7156 ( .A1(n5683), .A2(n5699), .ZN(n5690) );
  AND2_X1 U7157 ( .A1(n5691), .A2(n5690), .ZN(n6373) );
  NAND2_X1 U7158 ( .A1(n5693), .A2(n5692), .ZN(n6371) );
  NAND2_X1 U7159 ( .A1(n5694), .A2(n6371), .ZN(n8944) );
  NAND2_X1 U7160 ( .A1(n5698), .A2(n5699), .ZN(n5696) );
  NAND2_X1 U7161 ( .A1(n8948), .A2(n5743), .ZN(n5695) );
  NAND2_X1 U7162 ( .A1(n5696), .A2(n5695), .ZN(n5697) );
  XNOR2_X1 U7163 ( .A(n5697), .B(n5708), .ZN(n5702) );
  CLKBUF_X1 U7164 ( .A(n5698), .Z(n9003) );
  NAND2_X1 U7165 ( .A1(n5710), .A2(n9003), .ZN(n5701) );
  NAND2_X1 U7166 ( .A1(n8948), .A2(n5699), .ZN(n5700) );
  AND2_X1 U7167 ( .A1(n5701), .A2(n5700), .ZN(n5703) );
  NAND2_X1 U7168 ( .A1(n5702), .A2(n5703), .ZN(n6891) );
  INV_X1 U7169 ( .A(n5702), .ZN(n5705) );
  INV_X1 U7170 ( .A(n5703), .ZN(n5704) );
  NAND2_X1 U7171 ( .A1(n6889), .A2(n6891), .ZN(n5718) );
  OAI22_X1 U7172 ( .A1(n7032), .A2(n5707), .B1(n5706), .B2(n5899), .ZN(n5709)
         );
  XNOR2_X1 U7173 ( .A(n5709), .B(n5708), .ZN(n5714) );
  INV_X2 U7174 ( .A(n5710), .ZN(n5721) );
  OR2_X1 U7175 ( .A1(n7032), .A2(n5721), .ZN(n5712) );
  NAND2_X1 U7176 ( .A1(n5699), .A2(n7051), .ZN(n5711) );
  NAND2_X1 U7177 ( .A1(n5712), .A2(n5711), .ZN(n5715) );
  NAND2_X1 U7178 ( .A1(n5714), .A2(n5713), .ZN(n5719) );
  INV_X1 U7179 ( .A(n5714), .ZN(n5716) );
  NAND2_X1 U7180 ( .A1(n5716), .A2(n5715), .ZN(n5717) );
  AND2_X1 U7181 ( .A1(n5719), .A2(n5717), .ZN(n6892) );
  OAI22_X1 U7182 ( .A1(n7246), .A2(n4261), .B1(n7033), .B2(n5899), .ZN(n5720)
         );
  XNOR2_X1 U7183 ( .A(n5720), .B(n5708), .ZN(n5726) );
  OR2_X1 U7184 ( .A1(n7246), .A2(n5721), .ZN(n5723) );
  NAND2_X1 U7185 ( .A1(n7689), .A2(n7059), .ZN(n5722) );
  NAND2_X1 U7186 ( .A1(n5723), .A2(n5722), .ZN(n5724) );
  XNOR2_X1 U7187 ( .A(n5726), .B(n5724), .ZN(n7030) );
  NAND2_X1 U7188 ( .A1(n7029), .A2(n7030), .ZN(n7028) );
  INV_X1 U7189 ( .A(n5724), .ZN(n5725) );
  NAND2_X1 U7190 ( .A1(n5726), .A2(n5725), .ZN(n5727) );
  OAI22_X1 U7191 ( .A1(n7379), .A2(n4261), .B1(n7247), .B2(n5899), .ZN(n5728)
         );
  XNOR2_X1 U7192 ( .A(n5728), .B(n5708), .ZN(n7242) );
  OR2_X1 U7193 ( .A1(n7379), .A2(n5721), .ZN(n5730) );
  NAND2_X1 U7194 ( .A1(n7689), .A2(n7089), .ZN(n5729) );
  AND2_X1 U7195 ( .A1(n5730), .A2(n5729), .ZN(n5734) );
  AND2_X1 U7196 ( .A1(n7242), .A2(n5734), .ZN(n5738) );
  OAI22_X1 U7197 ( .A1(n7438), .A2(n4261), .B1(n7380), .B2(n5899), .ZN(n5731)
         );
  XNOR2_X1 U7198 ( .A(n5731), .B(n5708), .ZN(n5741) );
  OR2_X1 U7199 ( .A1(n7438), .A2(n5721), .ZN(n5733) );
  NAND2_X1 U7200 ( .A1(n7689), .A2(n7523), .ZN(n5732) );
  NAND2_X1 U7201 ( .A1(n5733), .A2(n5732), .ZN(n5739) );
  XNOR2_X1 U7202 ( .A(n5741), .B(n5739), .ZN(n7373) );
  INV_X1 U7203 ( .A(n7242), .ZN(n5735) );
  INV_X1 U7204 ( .A(n5734), .ZN(n7245) );
  NAND2_X1 U7205 ( .A1(n5735), .A2(n7245), .ZN(n5736) );
  AND2_X1 U7206 ( .A1(n7373), .A2(n5736), .ZN(n5737) );
  INV_X1 U7207 ( .A(n5739), .ZN(n5740) );
  NAND2_X1 U7208 ( .A1(n5741), .A2(n5740), .ZN(n5742) );
  NAND2_X1 U7209 ( .A1(n8998), .A2(n7689), .ZN(n5745) );
  NAND2_X1 U7210 ( .A1(n7098), .A2(n5743), .ZN(n5744) );
  NAND2_X1 U7211 ( .A1(n5745), .A2(n5744), .ZN(n5747) );
  XNOR2_X1 U7212 ( .A(n5747), .B(n5900), .ZN(n5750) );
  NAND2_X1 U7213 ( .A1(n5710), .A2(n8998), .ZN(n5749) );
  NAND2_X1 U7214 ( .A1(n7098), .A2(n7689), .ZN(n5748) );
  NAND2_X1 U7215 ( .A1(n5749), .A2(n5748), .ZN(n5751) );
  NAND2_X1 U7216 ( .A1(n5750), .A2(n5751), .ZN(n7432) );
  INV_X1 U7217 ( .A(n5750), .ZN(n5753) );
  INV_X1 U7218 ( .A(n5751), .ZN(n5752) );
  NAND2_X1 U7219 ( .A1(n5753), .A2(n5752), .ZN(n7434) );
  OR2_X1 U7220 ( .A1(n9637), .A2(n5721), .ZN(n5755) );
  NAND2_X1 U7221 ( .A1(n7689), .A2(n7603), .ZN(n5754) );
  OAI22_X1 U7222 ( .A1(n9637), .A2(n4261), .B1(n7557), .B2(n5899), .ZN(n5756)
         );
  XNOR2_X1 U7223 ( .A(n5756), .B(n5900), .ZN(n7555) );
  NAND2_X1 U7224 ( .A1(n7553), .A2(n7555), .ZN(n5758) );
  AND2_X1 U7225 ( .A1(n7434), .A2(n4317), .ZN(n5757) );
  NAND2_X1 U7226 ( .A1(n5758), .A2(n7554), .ZN(n7627) );
  NAND2_X1 U7227 ( .A1(n8996), .A2(n7689), .ZN(n5760) );
  NAND2_X1 U7228 ( .A1(n7635), .A2(n5743), .ZN(n5759) );
  NAND2_X1 U7229 ( .A1(n5760), .A2(n5759), .ZN(n5761) );
  XNOR2_X1 U7230 ( .A(n5761), .B(n5900), .ZN(n5765) );
  NAND2_X1 U7231 ( .A1(n5710), .A2(n8996), .ZN(n5763) );
  NAND2_X1 U7232 ( .A1(n7689), .A2(n7635), .ZN(n5762) );
  NAND2_X1 U7233 ( .A1(n5763), .A2(n5762), .ZN(n5766) );
  XNOR2_X1 U7234 ( .A(n5765), .B(n5766), .ZN(n7630) );
  INV_X1 U7235 ( .A(n5765), .ZN(n5768) );
  INV_X1 U7236 ( .A(n5766), .ZN(n5767) );
  NAND2_X1 U7237 ( .A1(n5768), .A2(n5767), .ZN(n5769) );
  OAI22_X1 U7238 ( .A1(n9636), .A2(n4261), .B1(n9570), .B2(n5899), .ZN(n5770)
         );
  XNOR2_X1 U7239 ( .A(n5770), .B(n5708), .ZN(n7653) );
  OR2_X1 U7240 ( .A1(n9636), .A2(n5721), .ZN(n5772) );
  NAND2_X1 U7241 ( .A1(n7689), .A2(n7619), .ZN(n5771) );
  AND2_X1 U7242 ( .A1(n5772), .A2(n5771), .ZN(n5773) );
  INV_X1 U7243 ( .A(n7653), .ZN(n5774) );
  INV_X1 U7244 ( .A(n5773), .ZN(n7652) );
  OAI22_X1 U7245 ( .A1(n9391), .A2(n4261), .B1(n9600), .B2(n5899), .ZN(n5775)
         );
  XNOR2_X1 U7246 ( .A(n5775), .B(n5708), .ZN(n5778) );
  OR2_X1 U7247 ( .A1(n9391), .A2(n5721), .ZN(n5777) );
  NAND2_X1 U7248 ( .A1(n9055), .A2(n7689), .ZN(n5776) );
  NAND2_X1 U7249 ( .A1(n5777), .A2(n5776), .ZN(n5779) );
  XNOR2_X1 U7250 ( .A(n5778), .B(n5779), .ZN(n7670) );
  NAND2_X1 U7251 ( .A1(n7669), .A2(n7670), .ZN(n5782) );
  INV_X1 U7252 ( .A(n5778), .ZN(n5780) );
  NAND2_X1 U7253 ( .A1(n5780), .A2(n5779), .ZN(n5781) );
  NAND2_X1 U7254 ( .A1(n5782), .A2(n5781), .ZN(n8873) );
  NAND2_X1 U7255 ( .A1(n9506), .A2(n5743), .ZN(n5784) );
  OR2_X1 U7256 ( .A1(n9589), .A2(n4261), .ZN(n5783) );
  NAND2_X1 U7257 ( .A1(n5784), .A2(n5783), .ZN(n5785) );
  XNOR2_X1 U7258 ( .A(n5785), .B(n5708), .ZN(n5788) );
  OR2_X1 U7259 ( .A1(n9589), .A2(n5721), .ZN(n5787) );
  NAND2_X1 U7260 ( .A1(n9506), .A2(n7689), .ZN(n5786) );
  AND2_X1 U7261 ( .A1(n5787), .A2(n5786), .ZN(n5789) );
  NAND2_X1 U7262 ( .A1(n5788), .A2(n5789), .ZN(n8874) );
  INV_X1 U7263 ( .A(n5788), .ZN(n5791) );
  INV_X1 U7264 ( .A(n5789), .ZN(n5790) );
  NAND2_X1 U7265 ( .A1(n5791), .A2(n5790), .ZN(n8875) );
  NAND2_X1 U7266 ( .A1(n9499), .A2(n5743), .ZN(n5793) );
  NAND2_X1 U7267 ( .A1(n9061), .A2(n7689), .ZN(n5792) );
  NAND2_X1 U7268 ( .A1(n5793), .A2(n5792), .ZN(n5794) );
  XNOR2_X1 U7269 ( .A(n5794), .B(n5900), .ZN(n8924) );
  NAND2_X1 U7270 ( .A1(n9499), .A2(n7689), .ZN(n5796) );
  NAND2_X1 U7271 ( .A1(n5710), .A2(n9061), .ZN(n5795) );
  NAND2_X1 U7272 ( .A1(n5796), .A2(n5795), .ZN(n8923) );
  NAND2_X1 U7273 ( .A1(n9495), .A2(n7689), .ZN(n5798) );
  OR2_X1 U7274 ( .A1(n9373), .A2(n5721), .ZN(n5797) );
  NAND2_X1 U7275 ( .A1(n5798), .A2(n5797), .ZN(n8833) );
  NAND2_X1 U7276 ( .A1(n9495), .A2(n5743), .ZN(n5800) );
  OR2_X1 U7277 ( .A1(n9373), .A2(n4261), .ZN(n5799) );
  NAND2_X1 U7278 ( .A1(n5800), .A2(n5799), .ZN(n5801) );
  XNOR2_X1 U7279 ( .A(n5801), .B(n5900), .ZN(n8832) );
  OAI21_X1 U7280 ( .B1(n8835), .B2(n8833), .A(n8832), .ZN(n5803) );
  NAND2_X1 U7281 ( .A1(n8835), .A2(n8833), .ZN(n5802) );
  NAND2_X1 U7282 ( .A1(n5803), .A2(n5802), .ZN(n8981) );
  NAND2_X1 U7283 ( .A1(n9487), .A2(n5743), .ZN(n5805) );
  NAND2_X1 U7284 ( .A1(n8994), .A2(n7689), .ZN(n5804) );
  NAND2_X1 U7285 ( .A1(n5805), .A2(n5804), .ZN(n5806) );
  XNOR2_X1 U7286 ( .A(n5806), .B(n5708), .ZN(n8979) );
  AND2_X1 U7287 ( .A1(n5710), .A2(n8994), .ZN(n5807) );
  AOI21_X1 U7288 ( .B1(n9487), .B2(n7689), .A(n5807), .ZN(n5809) );
  NAND2_X1 U7289 ( .A1(n8979), .A2(n5809), .ZN(n5808) );
  NAND2_X1 U7290 ( .A1(n8981), .A2(n5808), .ZN(n5812) );
  INV_X1 U7291 ( .A(n8979), .ZN(n5810) );
  INV_X1 U7292 ( .A(n5809), .ZN(n8978) );
  NAND2_X1 U7293 ( .A1(n5810), .A2(n8978), .ZN(n5811) );
  NAND2_X1 U7294 ( .A1(n5812), .A2(n5811), .ZN(n8892) );
  NAND2_X1 U7295 ( .A1(n9483), .A2(n5743), .ZN(n5814) );
  OR2_X1 U7296 ( .A1(n9336), .A2(n4261), .ZN(n5813) );
  NAND2_X1 U7297 ( .A1(n5814), .A2(n5813), .ZN(n5815) );
  XNOR2_X1 U7298 ( .A(n5815), .B(n5900), .ZN(n5818) );
  NAND2_X1 U7299 ( .A1(n9483), .A2(n7689), .ZN(n5817) );
  OR2_X1 U7300 ( .A1(n9336), .A2(n5721), .ZN(n5816) );
  NAND2_X1 U7301 ( .A1(n5817), .A2(n5816), .ZN(n5819) );
  AND2_X1 U7302 ( .A1(n5818), .A2(n5819), .ZN(n8894) );
  INV_X1 U7303 ( .A(n5818), .ZN(n5821) );
  INV_X1 U7304 ( .A(n5819), .ZN(n5820) );
  NAND2_X1 U7305 ( .A1(n5821), .A2(n5820), .ZN(n8893) );
  NAND2_X1 U7306 ( .A1(n9476), .A2(n5743), .ZN(n5823) );
  NAND2_X1 U7307 ( .A1(n9296), .A2(n7689), .ZN(n5822) );
  NAND2_X1 U7308 ( .A1(n5823), .A2(n5822), .ZN(n5824) );
  XNOR2_X1 U7309 ( .A(n5824), .B(n5708), .ZN(n7678) );
  AND2_X1 U7310 ( .A1(n5710), .A2(n9296), .ZN(n5825) );
  AOI21_X1 U7311 ( .B1(n9476), .B2(n7689), .A(n5825), .ZN(n7677) );
  AND2_X1 U7312 ( .A1(n7678), .A2(n7677), .ZN(n8952) );
  NAND2_X1 U7313 ( .A1(n9471), .A2(n7689), .ZN(n5827) );
  OR2_X1 U7314 ( .A1(n9275), .A2(n5721), .ZN(n5826) );
  NAND2_X1 U7315 ( .A1(n5827), .A2(n5826), .ZN(n8959) );
  INV_X1 U7316 ( .A(n8959), .ZN(n5834) );
  OR2_X1 U7317 ( .A1(n8952), .A2(n5834), .ZN(n5828) );
  NOR2_X1 U7318 ( .A1(n8953), .A2(n5828), .ZN(n5836) );
  NAND2_X1 U7319 ( .A1(n9471), .A2(n5743), .ZN(n5830) );
  OR2_X1 U7320 ( .A1(n9275), .A2(n4261), .ZN(n5829) );
  NAND2_X1 U7321 ( .A1(n5830), .A2(n5829), .ZN(n5831) );
  XNOR2_X1 U7322 ( .A(n5831), .B(n5708), .ZN(n5837) );
  INV_X1 U7323 ( .A(n7678), .ZN(n5833) );
  INV_X1 U7324 ( .A(n7677), .ZN(n5832) );
  NAND2_X1 U7325 ( .A1(n5833), .A2(n5832), .ZN(n5843) );
  AND2_X1 U7326 ( .A1(n5837), .A2(n5843), .ZN(n8954) );
  NOR2_X1 U7327 ( .A1(n5834), .A2(n8954), .ZN(n5835) );
  INV_X1 U7328 ( .A(n5837), .ZN(n5839) );
  INV_X1 U7329 ( .A(n8952), .ZN(n5838) );
  AND2_X1 U7330 ( .A1(n5839), .A2(n5838), .ZN(n5842) );
  AND2_X1 U7331 ( .A1(n8893), .A2(n5842), .ZN(n5840) );
  NAND2_X1 U7332 ( .A1(n5841), .A2(n5840), .ZN(n5846) );
  INV_X1 U7333 ( .A(n5842), .ZN(n5844) );
  OR2_X1 U7334 ( .A1(n5844), .A2(n5843), .ZN(n5845) );
  NAND2_X1 U7335 ( .A1(n9468), .A2(n5743), .ZN(n5849) );
  NAND2_X1 U7336 ( .A1(n9297), .A2(n7689), .ZN(n5848) );
  NAND2_X1 U7337 ( .A1(n5849), .A2(n5848), .ZN(n5850) );
  XNOR2_X1 U7338 ( .A(n5850), .B(n5900), .ZN(n5853) );
  NAND2_X1 U7339 ( .A1(n9468), .A2(n7689), .ZN(n5852) );
  NAND2_X1 U7340 ( .A1(n5710), .A2(n9297), .ZN(n5851) );
  NAND2_X1 U7341 ( .A1(n5852), .A2(n5851), .ZN(n5854) );
  AND2_X1 U7342 ( .A1(n5853), .A2(n5854), .ZN(n8855) );
  INV_X1 U7343 ( .A(n5853), .ZN(n5856) );
  INV_X1 U7344 ( .A(n5854), .ZN(n5855) );
  NAND2_X1 U7345 ( .A1(n5856), .A2(n5855), .ZN(n8854) );
  NAND2_X1 U7346 ( .A1(n9463), .A2(n5743), .ZN(n5858) );
  NAND2_X1 U7347 ( .A1(n9073), .A2(n7689), .ZN(n5857) );
  NAND2_X1 U7348 ( .A1(n5858), .A2(n5857), .ZN(n5859) );
  XNOR2_X1 U7349 ( .A(n5859), .B(n5708), .ZN(n5861) );
  AND2_X1 U7350 ( .A1(n5710), .A2(n9073), .ZN(n5860) );
  AOI21_X1 U7351 ( .B1(n9463), .B2(n7689), .A(n5860), .ZN(n5862) );
  AND2_X1 U7352 ( .A1(n5861), .A2(n5862), .ZN(n8915) );
  INV_X1 U7353 ( .A(n5861), .ZN(n5864) );
  INV_X1 U7354 ( .A(n5862), .ZN(n5863) );
  NAND2_X1 U7355 ( .A1(n5864), .A2(n5863), .ZN(n8913) );
  NAND2_X1 U7356 ( .A1(n9458), .A2(n5743), .ZN(n5867) );
  OR2_X1 U7357 ( .A1(n9262), .A2(n4261), .ZN(n5866) );
  NAND2_X1 U7358 ( .A1(n5867), .A2(n5866), .ZN(n5868) );
  XNOR2_X1 U7359 ( .A(n5868), .B(n5900), .ZN(n5871) );
  NAND2_X1 U7360 ( .A1(n9458), .A2(n7689), .ZN(n5870) );
  OR2_X1 U7361 ( .A1(n9262), .A2(n5721), .ZN(n5869) );
  NAND2_X1 U7362 ( .A1(n5870), .A2(n5869), .ZN(n5872) );
  NAND2_X1 U7363 ( .A1(n5871), .A2(n5872), .ZN(n8865) );
  INV_X1 U7364 ( .A(n5871), .ZN(n5874) );
  INV_X1 U7365 ( .A(n5872), .ZN(n5873) );
  NAND2_X1 U7366 ( .A1(n5874), .A2(n5873), .ZN(n8866) );
  AND2_X1 U7367 ( .A1(n5710), .A2(n9075), .ZN(n5875) );
  AOI21_X1 U7368 ( .B1(n9450), .B2(n7689), .A(n5875), .ZN(n5880) );
  NAND2_X1 U7369 ( .A1(n8934), .A2(n5880), .ZN(n5879) );
  NAND2_X1 U7370 ( .A1(n9450), .A2(n5743), .ZN(n5877) );
  NAND2_X1 U7371 ( .A1(n9075), .A2(n7689), .ZN(n5876) );
  NAND2_X1 U7372 ( .A1(n5877), .A2(n5876), .ZN(n5878) );
  NAND2_X1 U7373 ( .A1(n5879), .A2(n8936), .ZN(n5883) );
  INV_X1 U7374 ( .A(n8934), .ZN(n5881) );
  INV_X1 U7375 ( .A(n5880), .ZN(n8935) );
  NAND2_X1 U7376 ( .A1(n5881), .A2(n8935), .ZN(n5882) );
  NAND2_X1 U7377 ( .A1(n5883), .A2(n5882), .ZN(n5886) );
  OAI22_X1 U7378 ( .A1(n9225), .A2(n5899), .B1(n9203), .B2(n4261), .ZN(n5884)
         );
  XNOR2_X1 U7379 ( .A(n5884), .B(n5900), .ZN(n5885) );
  NAND2_X1 U7380 ( .A1(n5886), .A2(n5885), .ZN(n8843) );
  OAI22_X1 U7381 ( .A1(n9080), .A2(n5899), .B1(n9218), .B2(n4261), .ZN(n5887)
         );
  XNOR2_X1 U7382 ( .A(n5887), .B(n5708), .ZN(n5891) );
  OR2_X1 U7383 ( .A1(n9080), .A2(n4261), .ZN(n5889) );
  NAND2_X1 U7384 ( .A1(n9192), .A2(n5710), .ZN(n5888) );
  NAND2_X1 U7385 ( .A1(n5891), .A2(n5890), .ZN(n5892) );
  OAI21_X1 U7386 ( .B1(n5891), .B2(n5890), .A(n5892), .ZN(n8904) );
  INV_X1 U7387 ( .A(n5892), .ZN(n5893) );
  NAND2_X1 U7388 ( .A1(n9435), .A2(n5743), .ZN(n5895) );
  INV_X1 U7389 ( .A(n9204), .ZN(n9177) );
  NAND2_X1 U7390 ( .A1(n9177), .A2(n7689), .ZN(n5894) );
  NAND2_X1 U7391 ( .A1(n5895), .A2(n5894), .ZN(n5896) );
  XNOR2_X1 U7392 ( .A(n5896), .B(n5900), .ZN(n5898) );
  OAI22_X1 U7393 ( .A1(n9189), .A2(n4261), .B1(n9204), .B2(n5721), .ZN(n5897)
         );
  XNOR2_X1 U7394 ( .A(n5898), .B(n5897), .ZN(n8885) );
  NOR2_X1 U7395 ( .A1(n5898), .A2(n5897), .ZN(n8967) );
  OAI22_X1 U7396 ( .A1(n9172), .A2(n5899), .B1(n9158), .B2(n4261), .ZN(n5901)
         );
  XNOR2_X1 U7397 ( .A(n5901), .B(n5900), .ZN(n5905) );
  OR2_X1 U7398 ( .A1(n9172), .A2(n4261), .ZN(n5903) );
  NAND2_X1 U7399 ( .A1(n9193), .A2(n5710), .ZN(n5902) );
  NAND2_X1 U7400 ( .A1(n5903), .A2(n5902), .ZN(n5904) );
  XNOR2_X1 U7401 ( .A(n5905), .B(n5904), .ZN(n8966) );
  NAND2_X1 U7402 ( .A1(n9427), .A2(n5743), .ZN(n5907) );
  NAND2_X1 U7403 ( .A1(n9178), .A2(n7689), .ZN(n5906) );
  NAND2_X1 U7404 ( .A1(n5907), .A2(n5906), .ZN(n5908) );
  XNOR2_X1 U7405 ( .A(n5908), .B(n5708), .ZN(n5911) );
  NOR2_X1 U7406 ( .A1(n9143), .A2(n5721), .ZN(n5909) );
  AOI21_X1 U7407 ( .B1(n9427), .B2(n7689), .A(n5909), .ZN(n5910) );
  NAND2_X1 U7408 ( .A1(n5911), .A2(n5910), .ZN(n7697) );
  OAI21_X1 U7409 ( .B1(n5911), .B2(n5910), .A(n7697), .ZN(n5912) );
  OAI21_X1 U7410 ( .B1(n8965), .B2(n5913), .A(n5912), .ZN(n5914) );
  INV_X1 U7411 ( .A(n5914), .ZN(n5933) );
  INV_X1 U7412 ( .A(n6881), .ZN(n5915) );
  NAND2_X1 U7413 ( .A1(n7472), .A2(P1_B_REG_SCAN_IN), .ZN(n5917) );
  MUX2_X1 U7414 ( .A(n5917), .B(P1_B_REG_SCAN_IN), .S(n5932), .Z(n5918) );
  INV_X1 U7415 ( .A(n5916), .ZN(n5919) );
  NAND2_X1 U7416 ( .A1(n5919), .A2(n7472), .ZN(n5920) );
  OAI21_X1 U7417 ( .B1(n9653), .B2(P1_D_REG_1__SCAN_IN), .A(n5920), .ZN(n6286)
         );
  INV_X1 U7418 ( .A(n6286), .ZN(n9532) );
  NOR4_X1 U7419 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n5924) );
  NOR4_X1 U7420 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n5923) );
  NOR4_X1 U7421 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5922) );
  NOR4_X1 U7422 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5921) );
  NAND4_X1 U7423 ( .A1(n5924), .A2(n5923), .A3(n5922), .A4(n5921), .ZN(n5931)
         );
  NOR2_X1 U7424 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .ZN(
        n5928) );
  NOR4_X1 U7425 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n5927) );
  NOR4_X1 U7426 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n5926) );
  NOR4_X1 U7427 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n5925) );
  NAND4_X1 U7428 ( .A1(n5928), .A2(n5927), .A3(n5926), .A4(n5925), .ZN(n5930)
         );
  INV_X1 U7429 ( .A(n9653), .ZN(n5929) );
  OAI21_X1 U7430 ( .B1(n5931), .B2(n5930), .A(n5929), .ZN(n6285) );
  NAND2_X1 U7431 ( .A1(n9532), .A2(n6285), .ZN(n6868) );
  OAI22_X1 U7432 ( .A1(n9653), .A2(P1_D_REG_0__SCAN_IN), .B1(n5916), .B2(n5932), .ZN(n6661) );
  NOR2_X1 U7433 ( .A1(n6868), .A2(n6661), .ZN(n5937) );
  NAND2_X1 U7434 ( .A1(n5937), .A2(n9654), .ZN(n5942) );
  OAI21_X1 U7435 ( .B1(n7704), .B2(n5933), .A(n8970), .ZN(n5952) );
  AND3_X1 U7436 ( .A1(n6253), .A2(n5954), .A3(n5953), .ZN(n5935) );
  OR2_X1 U7437 ( .A1(n9568), .A2(n5937), .ZN(n6254) );
  NAND2_X1 U7438 ( .A1(n5935), .A2(n6254), .ZN(n5936) );
  NAND2_X1 U7439 ( .A1(n5936), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5940) );
  NOR2_X1 U7440 ( .A1(n6881), .A2(n6759), .ZN(n6872) );
  INV_X1 U7441 ( .A(n5937), .ZN(n5938) );
  AND2_X1 U7442 ( .A1(n5938), .A2(n9654), .ZN(n5939) );
  NAND2_X1 U7443 ( .A1(n6872), .A2(n5939), .ZN(n6256) );
  INV_X1 U7444 ( .A(n5942), .ZN(n5946) );
  NAND2_X2 U7445 ( .A1(n5941), .A2(n5946), .ZN(n8987) );
  NOR2_X1 U7446 ( .A1(n9158), .A2(n8987), .ZN(n5945) );
  INV_X1 U7447 ( .A(n6356), .ZN(n6716) );
  OR3_X1 U7448 ( .A1(n7003), .A2(n6716), .A3(n5942), .ZN(n6374) );
  OAI22_X1 U7449 ( .A1(n9089), .A2(n6374), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5943), .ZN(n5944) );
  AOI211_X1 U7450 ( .C1(n9162), .C2(n8982), .A(n5945), .B(n5944), .ZN(n5951)
         );
  NAND2_X1 U7451 ( .A1(n5946), .A2(n6872), .ZN(n5950) );
  INV_X1 U7452 ( .A(n9654), .ZN(n5948) );
  OR2_X1 U7453 ( .A1(n6284), .A2(n5948), .ZN(n5949) );
  NAND3_X1 U7454 ( .A1(n5952), .A2(n5951), .A3(n4833), .ZN(P1_U3212) );
  INV_X1 U7455 ( .A(n5953), .ZN(n5980) );
  NOR2_X2 U7456 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5969) );
  NOR2_X1 U7457 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5968) );
  NOR2_X1 U7458 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5967) );
  NOR2_X1 U7459 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5966) );
  NOR2_X1 U7460 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5971) );
  NAND4_X1 U7461 ( .A1(n5971), .A2(n6072), .A3(n5970), .A4(n5978), .ZN(n5972)
         );
  NAND2_X1 U7462 ( .A1(n4338), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U7463 ( .A1(n5975), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5976) );
  MUX2_X1 U7464 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5976), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5977) );
  NAND2_X1 U7465 ( .A1(n5977), .A2(n4338), .ZN(n7469) );
  OR2_X1 U7466 ( .A1(n6292), .A2(n5980), .ZN(n5981) );
  NAND2_X1 U7467 ( .A1(n5981), .A2(n6012), .ZN(n6010) );
  NAND2_X1 U7468 ( .A1(n6264), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AND2_X1 U7469 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7631) );
  INV_X1 U7470 ( .A(n6322), .ZN(n6043) );
  INV_X1 U7471 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5983) );
  AOI22_X1 U7472 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n6322), .B1(n6043), .B2(
        n5983), .ZN(n6318) );
  INV_X1 U7473 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5984) );
  MUX2_X1 U7474 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n5984), .S(n6396), .Z(n6392)
         );
  INV_X1 U7475 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6873) );
  MUX2_X1 U7476 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6873), .S(n6034), .Z(n6344)
         );
  NAND2_X1 U7477 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6354) );
  INV_X1 U7478 ( .A(n6354), .ZN(n6343) );
  NAND2_X1 U7479 ( .A1(n6344), .A2(n6343), .ZN(n6342) );
  NAND2_X1 U7480 ( .A1(n6034), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U7481 ( .A1(n6342), .A2(n5985), .ZN(n6391) );
  NAND2_X1 U7482 ( .A1(n6392), .A2(n6391), .ZN(n6390) );
  NAND2_X1 U7483 ( .A1(n6396), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7484 ( .A1(n6390), .A2(n5986), .ZN(n6279) );
  INV_X1 U7485 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5987) );
  XNOR2_X1 U7486 ( .A(n6270), .B(n5987), .ZN(n6280) );
  NAND2_X1 U7487 ( .A1(n6270), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5988) );
  INV_X1 U7488 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5989) );
  NOR2_X1 U7489 ( .A1(n6032), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9614) );
  NOR2_X1 U7490 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9609), .ZN(n5990) );
  AOI21_X1 U7491 ( .B1(n9609), .B2(P1_REG2_REG_5__SCAN_IN), .A(n5990), .ZN(
        n9613) );
  OAI21_X1 U7492 ( .B1(n9615), .B2(n9614), .A(n9613), .ZN(n9612) );
  XNOR2_X1 U7493 ( .A(n6695), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n6692) );
  NOR2_X1 U7494 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6335), .ZN(n5991) );
  AOI21_X1 U7495 ( .B1(n6335), .B2(P1_REG2_REG_7__SCAN_IN), .A(n5991), .ZN(
        n6331) );
  OAI21_X1 U7496 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6335), .A(n6329), .ZN(
        n6317) );
  NAND2_X1 U7497 ( .A1(n6318), .A2(n6317), .ZN(n6316) );
  OAI21_X1 U7498 ( .B1(n6322), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6316), .ZN(
        n5995) );
  NAND2_X1 U7499 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n6308), .ZN(n5992) );
  OAI21_X1 U7500 ( .B1(n6308), .B2(P1_REG2_REG_9__SCAN_IN), .A(n5992), .ZN(
        n5994) );
  NOR2_X1 U7501 ( .A1(n5994), .A2(n5995), .ZN(n6307) );
  OR2_X1 U7502 ( .A1(n5667), .A2(P1_U3084), .ZN(n9551) );
  INV_X1 U7503 ( .A(n9032), .ZN(n5993) );
  AOI211_X1 U7504 ( .C1(n5995), .C2(n5994), .A(n6307), .B(n9017), .ZN(n6016)
         );
  INV_X1 U7505 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7599) );
  NOR2_X1 U7506 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6335), .ZN(n6006) );
  INV_X1 U7507 ( .A(n6695), .ZN(n6036) );
  INV_X1 U7508 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U7509 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9609), .ZN(n6004) );
  INV_X1 U7510 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5996) );
  MUX2_X1 U7511 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n5996), .S(n6396), .Z(n5999)
         );
  INV_X1 U7512 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5997) );
  MUX2_X1 U7513 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n5997), .S(n6034), .Z(n6346)
         );
  AND2_X1 U7514 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6347) );
  NAND2_X1 U7515 ( .A1(n6346), .A2(n6347), .ZN(n6384) );
  NAND2_X1 U7516 ( .A1(n6034), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6383) );
  NAND2_X1 U7517 ( .A1(n6384), .A2(n6383), .ZN(n5998) );
  NAND2_X1 U7518 ( .A1(n5999), .A2(n5998), .ZN(n6387) );
  NAND2_X1 U7519 ( .A1(n6396), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U7520 ( .A1(n6387), .A2(n6271), .ZN(n6002) );
  INV_X1 U7521 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6000) );
  MUX2_X1 U7522 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6000), .S(n6270), .Z(n6001)
         );
  NAND2_X1 U7523 ( .A1(n6002), .A2(n6001), .ZN(n6274) );
  NAND2_X1 U7524 ( .A1(n6270), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6003) );
  AND2_X1 U7525 ( .A1(n6274), .A2(n6003), .ZN(n6363) );
  INV_X1 U7526 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7065) );
  MUX2_X1 U7527 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n7065), .S(n6032), .Z(n6362)
         );
  NAND2_X1 U7528 ( .A1(n6363), .A2(n6362), .ZN(n6361) );
  OAI21_X1 U7529 ( .B1(n6032), .B2(P1_REG1_REG_4__SCAN_IN), .A(n6361), .ZN(
        n9620) );
  INV_X1 U7530 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7074) );
  MUX2_X1 U7531 ( .A(n7074), .B(P1_REG1_REG_5__SCAN_IN), .S(n9609), .Z(n9619)
         );
  OR2_X1 U7532 ( .A1(n9620), .A2(n9619), .ZN(n9622) );
  NAND2_X1 U7533 ( .A1(n6004), .A2(n9622), .ZN(n6688) );
  MUX2_X1 U7534 ( .A(n6005), .B(P1_REG1_REG_6__SCAN_IN), .S(n6695), .Z(n6687)
         );
  NOR2_X1 U7535 ( .A1(n6688), .A2(n6687), .ZN(n6686) );
  AOI21_X1 U7536 ( .B1(n6036), .B2(n6005), .A(n6686), .ZN(n6334) );
  INV_X1 U7537 ( .A(n6335), .ZN(n6042) );
  INV_X1 U7538 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9692) );
  AOI22_X1 U7539 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6042), .B1(n6335), .B2(
        n9692), .ZN(n6333) );
  NOR2_X1 U7540 ( .A1(n6334), .A2(n6333), .ZN(n6332) );
  NOR2_X1 U7541 ( .A1(n6006), .A2(n6332), .ZN(n6321) );
  AOI22_X1 U7542 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n6043), .B1(n6322), .B2(
        n7599), .ZN(n6320) );
  NOR2_X1 U7543 ( .A1(n6321), .A2(n6320), .ZN(n6319) );
  AOI21_X1 U7544 ( .B1(n7599), .B2(n6043), .A(n6319), .ZN(n6008) );
  INV_X1 U7545 ( .A(n6308), .ZN(n6303) );
  INV_X1 U7546 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9695) );
  AOI22_X1 U7547 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n6303), .B1(n6308), .B2(
        n9695), .ZN(n6007) );
  NOR2_X1 U7548 ( .A1(n6008), .A2(n6007), .ZN(n6302) );
  AOI21_X1 U7549 ( .B1(n6008), .B2(n6007), .A(n6302), .ZN(n6011) );
  NOR2_X1 U7550 ( .A1(n6356), .A2(P1_U3084), .ZN(n9546) );
  NAND2_X1 U7551 ( .A1(n9546), .A2(n5667), .ZN(n6009) );
  NOR2_X1 U7552 ( .A1(n6011), .A2(n9030), .ZN(n6015) );
  INV_X1 U7553 ( .A(P1_U3083), .ZN(n6013) );
  INV_X1 U7554 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U7555 ( .A1(n9032), .A2(n6356), .ZN(n9029) );
  OAI22_X1 U7556 ( .A1(n9039), .A2(n9952), .B1(n9029), .B2(n6303), .ZN(n6014)
         );
  OR4_X1 U7557 ( .A1(n7631), .A2(n6016), .A3(n6015), .A4(n6014), .ZN(P1_U3250)
         );
  INV_X1 U7558 ( .A(n6017), .ZN(n6725) );
  AOI22_X1 U7559 ( .A1(n9549), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n6396), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6018) );
  OAI21_X1 U7560 ( .B1(n6725), .B2(n9552), .A(n6018), .ZN(P1_U3351) );
  AND2_X1 U7561 ( .A1(n6445), .A2(P2_U3152), .ZN(n6090) );
  INV_X2 U7562 ( .A(n6090), .ZN(n8830) );
  NOR2_X1 U7563 ( .A1(n6445), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8825) );
  INV_X2 U7564 ( .A(n8825), .ZN(n7667) );
  OR2_X1 U7565 ( .A1(n6019), .A2(n6071), .ZN(n6020) );
  XNOR2_X1 U7566 ( .A(n6020), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6520) );
  INV_X1 U7567 ( .A(n6520), .ZN(n6821) );
  OAI222_X1 U7568 ( .A1(n8830), .A2(n6818), .B1(n7667), .B2(n6816), .C1(
        P2_U3152), .C2(n6821), .ZN(P2_U3354) );
  OAI21_X1 U7569 ( .B1(P2_IR_REG_2__SCAN_IN), .B2(n4275), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6021) );
  XNOR2_X1 U7570 ( .A(n6021), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6518) );
  INV_X1 U7571 ( .A(n6518), .ZN(n6767) );
  INV_X1 U7572 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6765) );
  OAI222_X1 U7573 ( .A1(P2_U3152), .A2(n6767), .B1(n7667), .B2(n6766), .C1(
        n6765), .C2(n8830), .ZN(P2_U3355) );
  INV_X1 U7574 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7575 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4275), .ZN(n6022) );
  XNOR2_X1 U7576 ( .A(n6023), .B(n6022), .ZN(n6728) );
  OAI222_X1 U7577 ( .A1(P2_U3152), .A2(n6728), .B1(n7667), .B2(n6725), .C1(
        n4376), .C2(n8830), .ZN(P2_U3356) );
  NAND2_X1 U7578 ( .A1(n6024), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6025) );
  MUX2_X1 U7579 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6025), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n6027) );
  AND2_X1 U7580 ( .A1(n6027), .A2(n6026), .ZN(n6522) );
  INV_X1 U7581 ( .A(n6522), .ZN(n6834) );
  OAI222_X1 U7582 ( .A1(n8830), .A2(n6832), .B1(n7667), .B2(n6831), .C1(
        P2_U3152), .C2(n6834), .ZN(P2_U3353) );
  INV_X1 U7583 ( .A(n6028), .ZN(n6443) );
  INV_X1 U7584 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6441) );
  INV_X1 U7585 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6029) );
  OAI222_X1 U7586 ( .A1(n7667), .A2(n6443), .B1(n8830), .B2(n6441), .C1(
        P2_U3152), .C2(n6571), .ZN(P2_U3357) );
  AOI22_X1 U7587 ( .A1(n9609), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9549), .ZN(n6030) );
  OAI21_X1 U7588 ( .B1(n6831), .B2(n9552), .A(n6030), .ZN(P1_U3348) );
  NAND2_X1 U7589 ( .A1(n6026), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6031) );
  XNOR2_X1 U7590 ( .A(n6031), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6524) );
  INV_X1 U7591 ( .A(n6524), .ZN(n6930) );
  OAI222_X1 U7592 ( .A1(n8830), .A2(n6927), .B1(n7667), .B2(n6926), .C1(
        P2_U3152), .C2(n6930), .ZN(P2_U3352) );
  INV_X1 U7593 ( .A(n9549), .ZN(n7705) );
  INV_X1 U7594 ( .A(n6032), .ZN(n6367) );
  OAI222_X1 U7595 ( .A1(n7705), .A2(n6033), .B1(n9552), .B2(n6816), .C1(n6367), 
        .C2(P1_U3084), .ZN(P1_U3349) );
  INV_X1 U7596 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6035) );
  OAI222_X1 U7597 ( .A1(n7705), .A2(n6035), .B1(n9552), .B2(n6443), .C1(
        P1_U3084), .C2(n4927), .ZN(P1_U3352) );
  OAI222_X1 U7598 ( .A1(n7705), .A2(n6037), .B1(n9552), .B2(n6926), .C1(n6036), 
        .C2(P1_U3084), .ZN(P1_U3347) );
  INV_X1 U7599 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6038) );
  INV_X1 U7600 ( .A(n6270), .ZN(n6276) );
  OAI222_X1 U7601 ( .A1(n7705), .A2(n6038), .B1(n9552), .B2(n6766), .C1(n6276), 
        .C2(P1_U3084), .ZN(P1_U3350) );
  INV_X1 U7602 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7131) );
  INV_X1 U7603 ( .A(n6039), .ZN(n7130) );
  XNOR2_X1 U7604 ( .A(n6040), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6526) );
  INV_X1 U7605 ( .A(n6526), .ZN(n7134) );
  OAI222_X1 U7606 ( .A1(n8830), .A2(n7131), .B1(n7667), .B2(n7130), .C1(
        P2_U3152), .C2(n7134), .ZN(P2_U3351) );
  INV_X1 U7607 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6041) );
  OAI222_X1 U7608 ( .A1(n6042), .A2(P1_U3084), .B1(n9552), .B2(n7130), .C1(
        n6041), .C2(n7705), .ZN(P1_U3346) );
  INV_X1 U7609 ( .A(n7111), .ZN(n6046) );
  OAI222_X1 U7610 ( .A1(n6043), .A2(P1_U3084), .B1(n9552), .B2(n6046), .C1(
        n6186), .C2(n7705), .ZN(P1_U3345) );
  NAND2_X1 U7611 ( .A1(n6044), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6045) );
  XNOR2_X1 U7612 ( .A(n6045), .B(n4814), .ZN(n7112) );
  OAI222_X1 U7613 ( .A1(n8830), .A2(n7113), .B1(n7667), .B2(n6046), .C1(
        P2_U3152), .C2(n7112), .ZN(P2_U3350) );
  INV_X1 U7614 ( .A(n7452), .ZN(n6063) );
  NAND2_X1 U7615 ( .A1(n6047), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6052) );
  INV_X1 U7616 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7617 ( .A1(n6052), .A2(n6051), .ZN(n6054) );
  NAND2_X1 U7618 ( .A1(n6054), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6048) );
  XNOR2_X1 U7619 ( .A(n6048), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7453) );
  AOI22_X1 U7620 ( .A1(n7453), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n6090), .ZN(n6049) );
  OAI21_X1 U7621 ( .B1(n6063), .B2(n7667), .A(n6049), .ZN(P2_U3347) );
  INV_X1 U7622 ( .A(n7314), .ZN(n6056) );
  OAI222_X1 U7623 ( .A1(P1_U3084), .A2(n6400), .B1(n9552), .B2(n6056), .C1(
        n6050), .C2(n7705), .ZN(P1_U3343) );
  OR2_X1 U7624 ( .A1(n6052), .A2(n6051), .ZN(n6053) );
  INV_X1 U7625 ( .A(n7313), .ZN(n6559) );
  OAI222_X1 U7626 ( .A1(P2_U3152), .A2(n6559), .B1(n7667), .B2(n6056), .C1(
        n6055), .C2(n8830), .ZN(P2_U3348) );
  INV_X1 U7627 ( .A(n7285), .ZN(n6061) );
  OR2_X1 U7628 ( .A1(n6057), .A2(n6071), .ZN(n6058) );
  XNOR2_X1 U7629 ( .A(n6058), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7286) );
  OAI222_X1 U7630 ( .A1(n8830), .A2(n6059), .B1(n7667), .B2(n6061), .C1(n4449), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  OAI222_X1 U7631 ( .A1(P1_U3084), .A2(n6303), .B1(n9552), .B2(n6061), .C1(
        n6060), .C2(n7705), .ZN(P1_U3344) );
  INV_X1 U7632 ( .A(n6641), .ZN(n6408) );
  OAI222_X1 U7633 ( .A1(P1_U3084), .A2(n6408), .B1(n9552), .B2(n6063), .C1(
        n6062), .C2(n7705), .ZN(P1_U3342) );
  INV_X1 U7634 ( .A(n6642), .ZN(n6653) );
  INV_X1 U7635 ( .A(n7538), .ZN(n6067) );
  OAI222_X1 U7636 ( .A1(n6653), .A2(P1_U3084), .B1(n9552), .B2(n6067), .C1(
        n6064), .C2(n7705), .ZN(P1_U3341) );
  NAND2_X1 U7637 ( .A1(n6065), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6066) );
  XNOR2_X1 U7638 ( .A(n6066), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7539) );
  INV_X1 U7639 ( .A(n7539), .ZN(n6539) );
  OAI222_X1 U7640 ( .A1(n8830), .A2(n6068), .B1(n7667), .B2(n6067), .C1(
        P2_U3152), .C2(n6539), .ZN(P2_U3346) );
  INV_X1 U7641 ( .A(n7577), .ZN(n6069) );
  INV_X1 U7642 ( .A(n6954), .ZN(n6638) );
  OAI222_X1 U7643 ( .A1(n7705), .A2(n6070), .B1(n9552), .B2(n6069), .C1(
        P1_U3084), .C2(n6638), .ZN(P1_U3340) );
  INV_X1 U7644 ( .A(n7725), .ZN(n6076) );
  OR2_X1 U7645 ( .A1(n4335), .A2(n6071), .ZN(n6089) );
  NAND2_X1 U7646 ( .A1(n6089), .A2(n6072), .ZN(n6073) );
  NAND2_X1 U7647 ( .A1(n6073), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6232) );
  XNOR2_X1 U7648 ( .A(n6232), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7726) );
  INV_X1 U7649 ( .A(n7726), .ZN(n7422) );
  OAI222_X1 U7650 ( .A1(n8830), .A2(n6074), .B1(n7667), .B2(n6076), .C1(n7422), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U7651 ( .A(n7278), .ZN(n7269) );
  OAI222_X1 U7652 ( .A1(P1_U3084), .A2(n7269), .B1(n9552), .B2(n6076), .C1(
        n6075), .C2(n7705), .ZN(P1_U3339) );
  OR2_X1 U7653 ( .A1(n6670), .A2(P2_U3152), .ZN(n8309) );
  NAND2_X1 U7654 ( .A1(n9782), .A2(n8309), .ZN(n6082) );
  NAND2_X1 U7655 ( .A1(n6081), .A2(n6080), .ZN(n6079) );
  NAND2_X1 U7656 ( .A1(n6082), .A2(n7794), .ZN(n6088) );
  NAND2_X1 U7657 ( .A1(n6085), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6086) );
  OR2_X1 U7658 ( .A1(n9782), .A2(n6676), .ZN(n6087) );
  NOR2_X1 U7659 ( .A1(n9715), .A2(P2_U3966), .ZN(P2_U3151) );
  XNOR2_X1 U7660 ( .A(n6089), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7578) );
  AOI222_X1 U7661 ( .A1(n7577), .A2(n8825), .B1(n7578), .B2(
        P2_STATE_REG_SCAN_IN), .C1(P1_DATAO_REG_13__SCAN_IN), .C2(n6090), .ZN(
        n6211) );
  INV_X1 U7662 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9879) );
  AOI22_X1 U7663 ( .A1(n7582), .A2(keyinput55), .B1(keyinput6), .B2(n9879), 
        .ZN(n6091) );
  OAI221_X1 U7664 ( .B1(n7582), .B2(keyinput55), .C1(n9879), .C2(keyinput6), 
        .A(n6091), .ZN(n6101) );
  INV_X1 U7665 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n6093) );
  AOI22_X1 U7666 ( .A1(n6093), .A2(keyinput51), .B1(n5009), .B2(keyinput3), 
        .ZN(n6092) );
  OAI221_X1 U7667 ( .B1(n6093), .B2(keyinput51), .C1(n5009), .C2(keyinput3), 
        .A(n6092), .ZN(n6100) );
  INV_X1 U7668 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n6095) );
  AOI22_X1 U7669 ( .A1(n6095), .A2(keyinput10), .B1(n6241), .B2(keyinput18), 
        .ZN(n6094) );
  OAI221_X1 U7670 ( .B1(n6095), .B2(keyinput10), .C1(n6241), .C2(keyinput18), 
        .A(n6094), .ZN(n6099) );
  XNOR2_X1 U7671 ( .A(P2_REG1_REG_20__SCAN_IN), .B(keyinput63), .ZN(n6097) );
  XNOR2_X1 U7672 ( .A(SI_3_), .B(keyinput36), .ZN(n6096) );
  NAND2_X1 U7673 ( .A1(n6097), .A2(n6096), .ZN(n6098) );
  NOR4_X1 U7674 ( .A1(n6101), .A2(n6100), .A3(n6099), .A4(n6098), .ZN(n6134)
         );
  INV_X1 U7675 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n9795) );
  INV_X1 U7676 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9608) );
  AOI22_X1 U7677 ( .A1(n9795), .A2(keyinput44), .B1(keyinput49), .B2(n9608), 
        .ZN(n6102) );
  OAI221_X1 U7678 ( .B1(n9795), .B2(keyinput44), .C1(n9608), .C2(keyinput49), 
        .A(n6102), .ZN(n6111) );
  INV_X1 U7679 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6105) );
  INV_X1 U7680 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n6104) );
  AOI22_X1 U7681 ( .A1(n6105), .A2(keyinput22), .B1(keyinput9), .B2(n6104), 
        .ZN(n6103) );
  OAI221_X1 U7682 ( .B1(n6105), .B2(keyinput22), .C1(n6104), .C2(keyinput9), 
        .A(n6103), .ZN(n6110) );
  AOI22_X1 U7683 ( .A1(n7638), .A2(keyinput39), .B1(n8859), .B2(keyinput1), 
        .ZN(n6106) );
  OAI221_X1 U7684 ( .B1(n7638), .B2(keyinput39), .C1(n8859), .C2(keyinput1), 
        .A(n6106), .ZN(n6109) );
  INV_X1 U7685 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n9655) );
  AOI22_X1 U7686 ( .A1(n9655), .A2(keyinput26), .B1(keyinput61), .B2(n4448), 
        .ZN(n6107) );
  OAI221_X1 U7687 ( .B1(n9655), .B2(keyinput26), .C1(n4448), .C2(keyinput61), 
        .A(n6107), .ZN(n6108) );
  NOR4_X1 U7688 ( .A1(n6111), .A2(n6110), .A3(n6109), .A4(n6108), .ZN(n6133)
         );
  INV_X1 U7689 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n9794) );
  AOI22_X1 U7690 ( .A1(n8829), .A2(keyinput30), .B1(keyinput8), .B2(n9794), 
        .ZN(n6112) );
  OAI221_X1 U7691 ( .B1(n8829), .B2(keyinput30), .C1(n9794), .C2(keyinput8), 
        .A(n6112), .ZN(n6120) );
  AOI22_X1 U7692 ( .A1(P2_U3152), .A2(keyinput14), .B1(n7470), .B2(keyinput21), 
        .ZN(n6113) );
  OAI221_X1 U7693 ( .B1(P2_U3152), .B2(keyinput14), .C1(n7470), .C2(keyinput21), .A(n6113), .ZN(n6119) );
  INV_X1 U7694 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6185) );
  AOI22_X1 U7695 ( .A1(n6185), .A2(keyinput35), .B1(n5131), .B2(keyinput31), 
        .ZN(n6114) );
  OAI221_X1 U7696 ( .B1(n6185), .B2(keyinput35), .C1(n5131), .C2(keyinput31), 
        .A(n6114), .ZN(n6118) );
  INV_X1 U7697 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n9798) );
  INV_X1 U7698 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6116) );
  AOI22_X1 U7699 ( .A1(n9798), .A2(keyinput0), .B1(keyinput46), .B2(n6116), 
        .ZN(n6115) );
  OAI221_X1 U7700 ( .B1(n9798), .B2(keyinput0), .C1(n6116), .C2(keyinput46), 
        .A(n6115), .ZN(n6117) );
  NOR4_X1 U7701 ( .A1(n6120), .A2(n6119), .A3(n6118), .A4(n6117), .ZN(n6132)
         );
  INV_X1 U7702 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9855) );
  INV_X1 U7703 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9911) );
  AOI22_X1 U7704 ( .A1(n9855), .A2(keyinput23), .B1(n9911), .B2(keyinput54), 
        .ZN(n6121) );
  OAI221_X1 U7705 ( .B1(n9855), .B2(keyinput23), .C1(n9911), .C2(keyinput54), 
        .A(n6121), .ZN(n6130) );
  INV_X1 U7706 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9656) );
  INV_X1 U7707 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n6123) );
  AOI22_X1 U7708 ( .A1(n9656), .A2(keyinput29), .B1(keyinput58), .B2(n6123), 
        .ZN(n6122) );
  OAI221_X1 U7709 ( .B1(n9656), .B2(keyinput29), .C1(n6123), .C2(keyinput58), 
        .A(n6122), .ZN(n6129) );
  INV_X1 U7710 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9657) );
  XNOR2_X1 U7711 ( .A(n9657), .B(keyinput20), .ZN(n6128) );
  XNOR2_X1 U7712 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput4), .ZN(n6126) );
  XNOR2_X1 U7713 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput13), .ZN(n6125) );
  XNOR2_X1 U7714 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput47), .ZN(n6124) );
  NAND3_X1 U7715 ( .A1(n6126), .A2(n6125), .A3(n6124), .ZN(n6127) );
  NOR4_X1 U7716 ( .A1(n6130), .A2(n6129), .A3(n6128), .A4(n6127), .ZN(n6131)
         );
  NAND4_X1 U7717 ( .A1(n6134), .A2(n6133), .A3(n6132), .A4(n6131), .ZN(n6184)
         );
  INV_X1 U7718 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n9803) );
  AOI22_X1 U7719 ( .A1(n6136), .A2(keyinput48), .B1(keyinput19), .B2(n9803), 
        .ZN(n6135) );
  OAI221_X1 U7720 ( .B1(n6136), .B2(keyinput48), .C1(n9803), .C2(keyinput19), 
        .A(n6135), .ZN(n6146) );
  INV_X1 U7721 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n6139) );
  INV_X1 U7722 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n6138) );
  AOI22_X1 U7723 ( .A1(n6139), .A2(keyinput12), .B1(keyinput43), .B2(n6138), 
        .ZN(n6137) );
  OAI221_X1 U7724 ( .B1(n6139), .B2(keyinput12), .C1(n6138), .C2(keyinput43), 
        .A(n6137), .ZN(n6145) );
  INV_X1 U7725 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9027) );
  AOI22_X1 U7726 ( .A1(n9027), .A2(keyinput41), .B1(keyinput11), .B2(n6141), 
        .ZN(n6140) );
  OAI221_X1 U7727 ( .B1(n9027), .B2(keyinput41), .C1(n6141), .C2(keyinput11), 
        .A(n6140), .ZN(n6144) );
  INV_X1 U7728 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9658) );
  INV_X1 U7729 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9863) );
  AOI22_X1 U7730 ( .A1(n9658), .A2(keyinput45), .B1(keyinput25), .B2(n9863), 
        .ZN(n6142) );
  OAI221_X1 U7731 ( .B1(n9658), .B2(keyinput45), .C1(n9863), .C2(keyinput25), 
        .A(n6142), .ZN(n6143) );
  NOR4_X1 U7732 ( .A1(n6146), .A2(n6145), .A3(n6144), .A4(n6143), .ZN(n6182)
         );
  INV_X1 U7733 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9711) );
  INV_X1 U7734 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6148) );
  AOI22_X1 U7735 ( .A1(n9711), .A2(keyinput7), .B1(n6148), .B2(keyinput24), 
        .ZN(n6147) );
  OAI221_X1 U7736 ( .B1(n9711), .B2(keyinput7), .C1(n6148), .C2(keyinput24), 
        .A(n6147), .ZN(n6158) );
  INV_X1 U7737 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6150) );
  AOI22_X1 U7738 ( .A1(n6150), .A2(keyinput16), .B1(n6381), .B2(keyinput60), 
        .ZN(n6149) );
  OAI221_X1 U7739 ( .B1(n6150), .B2(keyinput16), .C1(n6381), .C2(keyinput60), 
        .A(n6149), .ZN(n6157) );
  AOI22_X1 U7740 ( .A1(n6186), .A2(keyinput37), .B1(n6152), .B2(keyinput59), 
        .ZN(n6151) );
  OAI221_X1 U7741 ( .B1(n6186), .B2(keyinput37), .C1(n6152), .C2(keyinput59), 
        .A(n6151), .ZN(n6156) );
  XNOR2_X1 U7742 ( .A(P2_REG0_REG_23__SCAN_IN), .B(keyinput40), .ZN(n6154) );
  XNOR2_X1 U7743 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput33), .ZN(n6153) );
  NAND2_X1 U7744 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  NOR4_X1 U7745 ( .A1(n6158), .A2(n6157), .A3(n6156), .A4(n6155), .ZN(n6181)
         );
  AOI22_X1 U7746 ( .A1(n6378), .A2(keyinput52), .B1(n4535), .B2(keyinput15), 
        .ZN(n6159) );
  OAI221_X1 U7747 ( .B1(n6378), .B2(keyinput52), .C1(n4535), .C2(keyinput15), 
        .A(n6159), .ZN(n6168) );
  INV_X1 U7748 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n9804) );
  AOI22_X1 U7749 ( .A1(n4983), .A2(keyinput32), .B1(keyinput53), .B2(n9804), 
        .ZN(n6160) );
  OAI221_X1 U7750 ( .B1(n4983), .B2(keyinput32), .C1(n9804), .C2(keyinput53), 
        .A(n6160), .ZN(n6167) );
  INV_X1 U7751 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6162) );
  INV_X1 U7752 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7530) );
  AOI22_X1 U7753 ( .A1(n6162), .A2(keyinput34), .B1(n7530), .B2(keyinput56), 
        .ZN(n6161) );
  OAI221_X1 U7754 ( .B1(n6162), .B2(keyinput34), .C1(n7530), .C2(keyinput56), 
        .A(n6161), .ZN(n6166) );
  XNOR2_X1 U7755 ( .A(P2_REG1_REG_22__SCAN_IN), .B(keyinput17), .ZN(n6164) );
  XNOR2_X1 U7756 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput5), .ZN(n6163) );
  NAND2_X1 U7757 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  NOR4_X1 U7758 ( .A1(n6168), .A2(n6167), .A3(n6166), .A4(n6165), .ZN(n6180)
         );
  INV_X1 U7759 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n9788) );
  AOI22_X1 U7760 ( .A1(n9788), .A2(keyinput62), .B1(n6170), .B2(keyinput27), 
        .ZN(n6169) );
  OAI221_X1 U7761 ( .B1(n9788), .B2(keyinput62), .C1(n6170), .C2(keyinput27), 
        .A(n6169), .ZN(n6178) );
  INV_X1 U7762 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n9797) );
  AOI22_X1 U7763 ( .A1(n9797), .A2(keyinput50), .B1(n6758), .B2(keyinput38), 
        .ZN(n6171) );
  OAI221_X1 U7764 ( .B1(n9797), .B2(keyinput50), .C1(n6758), .C2(keyinput38), 
        .A(n6171), .ZN(n6177) );
  INV_X1 U7765 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n6190) );
  INV_X1 U7766 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7546) );
  AOI22_X1 U7767 ( .A1(n6190), .A2(keyinput28), .B1(n7546), .B2(keyinput2), 
        .ZN(n6172) );
  OAI221_X1 U7768 ( .B1(n6190), .B2(keyinput28), .C1(n7546), .C2(keyinput2), 
        .A(n6172), .ZN(n6176) );
  XNOR2_X1 U7769 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput42), .ZN(n6174) );
  XNOR2_X1 U7770 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput57), .ZN(n6173) );
  NAND2_X1 U7771 ( .A1(n6174), .A2(n6173), .ZN(n6175) );
  NOR4_X1 U7772 ( .A1(n6178), .A2(n6177), .A3(n6176), .A4(n6175), .ZN(n6179)
         );
  NAND4_X1 U7773 ( .A1(n6182), .A2(n6181), .A3(n6180), .A4(n6179), .ZN(n6183)
         );
  NOR2_X1 U7774 ( .A1(n6184), .A2(n6183), .ZN(n6209) );
  NOR4_X1 U7775 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(P2_DATAO_REG_25__SCAN_IN), 
        .A3(P1_REG3_REG_19__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6207) );
  NOR2_X1 U7776 ( .A1(n9711), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6564) );
  INV_X1 U7777 ( .A(n6564), .ZN(n6189) );
  NAND4_X1 U7778 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_1__SCAN_IN), 
        .A3(n6186), .A4(n6185), .ZN(n6188) );
  NAND4_X1 U7779 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(SI_3_), .A3(n6758), .A4(
        n4535), .ZN(n6187) );
  NOR4_X1 U7780 ( .A1(n6190), .A2(n6189), .A3(n6188), .A4(n6187), .ZN(n6206)
         );
  NAND4_X1 U7781 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_DATAO_REG_16__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .A4(P2_REG1_REG_20__SCAN_IN), .ZN(n6194)
         );
  NAND4_X1 U7782 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_REG0_REG_19__SCAN_IN), .A4(P2_REG0_REG_23__SCAN_IN), .ZN(n6193) );
  NAND4_X1 U7783 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_REG0_REG_10__SCAN_IN), .A4(P2_REG0_REG_7__SCAN_IN), .ZN(n6192) );
  NAND4_X1 U7784 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .A3(
        P2_REG3_REG_13__SCAN_IN), .A4(P2_REG3_REG_12__SCAN_IN), .ZN(n6191) );
  NOR4_X1 U7785 ( .A1(n6194), .A2(n6193), .A3(n6192), .A4(n6191), .ZN(n6205)
         );
  NOR4_X1 U7786 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_REG0_REG_25__SCAN_IN), 
        .A3(P2_REG1_REG_22__SCAN_IN), .A4(P2_REG0_REG_30__SCAN_IN), .ZN(n6198)
         );
  NOR4_X1 U7787 ( .A1(P1_REG0_REG_6__SCAN_IN), .A2(P2_REG1_REG_12__SCAN_IN), 
        .A3(P2_REG1_REG_9__SCAN_IN), .A4(P2_REG0_REG_8__SCAN_IN), .ZN(n6197)
         );
  NOR4_X1 U7788 ( .A1(SI_23_), .A2(P1_REG2_REG_21__SCAN_IN), .A3(
        P1_REG2_REG_16__SCAN_IN), .A4(P2_WR_REG_SCAN_IN), .ZN(n6196) );
  INV_X1 U7789 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8359) );
  NOR4_X1 U7790 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG2_REG_24__SCAN_IN), 
        .A3(n6381), .A4(n8359), .ZN(n6195) );
  NAND4_X1 U7791 ( .A1(n6198), .A2(n6197), .A3(n6196), .A4(n6195), .ZN(n6203)
         );
  NAND4_X1 U7792 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_IR_REG_29__SCAN_IN), .A4(P1_REG0_REG_29__SCAN_IN), .ZN(n6202) );
  NAND4_X1 U7793 ( .A1(P1_D_REG_22__SCAN_IN), .A2(SI_24_), .A3(
        P1_REG3_REG_7__SCAN_IN), .A4(P1_REG3_REG_6__SCAN_IN), .ZN(n6201) );
  NAND3_X1 U7794 ( .A1(n9788), .A2(n9798), .A3(n9803), .ZN(n6422) );
  NAND4_X1 U7795 ( .A1(P1_REG1_REG_21__SCAN_IN), .A2(P1_REG1_REG_19__SCAN_IN), 
        .A3(P1_REG1_REG_18__SCAN_IN), .A4(P2_REG2_REG_18__SCAN_IN), .ZN(n6199)
         );
  OR4_X1 U7796 ( .A1(n7638), .A2(n5131), .A3(n6422), .A4(n6199), .ZN(n6200) );
  NOR4_X1 U7797 ( .A1(n6203), .A2(n6202), .A3(n6201), .A4(n6200), .ZN(n6204)
         );
  NAND4_X1 U7798 ( .A1(n6207), .A2(n6206), .A3(n6205), .A4(n6204), .ZN(n6208)
         );
  XNOR2_X1 U7799 ( .A(n6209), .B(n6208), .ZN(n6210) );
  XNOR2_X1 U7800 ( .A(n6211), .B(n6210), .ZN(P2_U3345) );
  INV_X1 U7801 ( .A(n6218), .ZN(n7666) );
  AND2_X4 U7802 ( .A1(n7666), .A2(n6224), .ZN(n6750) );
  NAND2_X1 U7803 ( .A1(n6750), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6222) );
  INV_X4 U7804 ( .A(n7931), .ZN(n8105) );
  NAND2_X1 U7805 ( .A1(n8105), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6221) );
  AND2_X2 U7806 ( .A1(n7666), .A2(n6219), .ZN(n6463) );
  NAND2_X1 U7807 ( .A1(n8106), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7808 ( .A1(n4638), .A2(P2_U3966), .ZN(n6223) );
  OAI21_X1 U7809 ( .B1(P2_U3966), .B2(n5491), .A(n6223), .ZN(P2_U3583) );
  NAND2_X1 U7810 ( .A1(n6462), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6228) );
  NAND2_X1 U7811 ( .A1(n7916), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6227) );
  NAND2_X1 U7812 ( .A1(n6750), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U7813 ( .A1(n6463), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6225) );
  NAND4_X2 U7814 ( .A1(n6228), .A2(n6227), .A3(n6226), .A4(n6225), .ZN(n6453)
         );
  NAND2_X1 U7815 ( .A1(n6453), .A2(P2_U3966), .ZN(n6229) );
  OAI21_X1 U7816 ( .B1(P2_U3966), .B2(n4534), .A(n6229), .ZN(P2_U3552) );
  INV_X1 U7817 ( .A(n7744), .ZN(n6235) );
  OAI222_X1 U7818 ( .A1(n7497), .A2(P1_U3084), .B1(n9552), .B2(n6235), .C1(
        n6230), .C2(n7705), .ZN(P1_U3338) );
  NAND2_X1 U7819 ( .A1(n6232), .A2(n6231), .ZN(n6233) );
  NAND2_X1 U7820 ( .A1(n6233), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6234) );
  XNOR2_X1 U7821 ( .A(n6234), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8330) );
  INV_X1 U7822 ( .A(n8330), .ZN(n8322) );
  OAI222_X1 U7823 ( .A1(n8830), .A2(n6236), .B1(n7667), .B2(n6235), .C1(
        P2_U3152), .C2(n8322), .ZN(P2_U3343) );
  NAND2_X1 U7824 ( .A1(n5674), .A2(n9004), .ZN(n6237) );
  OAI21_X1 U7825 ( .B1(n9004), .B2(n4535), .A(n6237), .ZN(P1_U3555) );
  NAND2_X1 U7826 ( .A1(n6238), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6239) );
  MUX2_X1 U7827 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6239), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6240) );
  INV_X1 U7828 ( .A(n6298), .ZN(n6246) );
  AND2_X1 U7829 ( .A1(n6240), .A2(n6246), .ZN(n8349) );
  INV_X1 U7830 ( .A(n8349), .ZN(n6242) );
  INV_X1 U7831 ( .A(n7736), .ZN(n6243) );
  OAI222_X1 U7832 ( .A1(P2_U3152), .A2(n6242), .B1(n7667), .B2(n6243), .C1(
        n6241), .C2(n8830), .ZN(P2_U3342) );
  INV_X1 U7833 ( .A(n7644), .ZN(n7503) );
  OAI222_X1 U7834 ( .A1(n7705), .A2(n6244), .B1(n9552), .B2(n6243), .C1(
        P1_U3084), .C2(n7503), .ZN(P1_U3337) );
  INV_X1 U7835 ( .A(n7764), .ZN(n6249) );
  AOI22_X1 U7836 ( .A1(n9015), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9549), .ZN(n6245) );
  OAI21_X1 U7837 ( .B1(n6249), .B2(n9552), .A(n6245), .ZN(P1_U3336) );
  NAND2_X1 U7838 ( .A1(n6246), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6247) );
  XNOR2_X1 U7839 ( .A(n6247), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8363) );
  INV_X1 U7840 ( .A(n8363), .ZN(n8356) );
  OAI222_X1 U7841 ( .A1(P2_U3152), .A2(n8356), .B1(n7667), .B2(n6249), .C1(
        n6248), .C2(n8830), .ZN(P2_U3341) );
  OAI21_X1 U7842 ( .B1(n6252), .B2(n6250), .A(n6251), .ZN(n6353) );
  INV_X1 U7843 ( .A(n6353), .ZN(n6259) );
  INV_X1 U7844 ( .A(n6870), .ZN(n6255) );
  NAND3_X1 U7845 ( .A1(n6256), .A2(n6255), .A3(n6254), .ZN(n8947) );
  OAI22_X1 U7846 ( .A1(n8977), .A2(n6704), .B1(n6698), .B2(n6374), .ZN(n6257)
         );
  AOI21_X1 U7847 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n8947), .A(n6257), .ZN(
        n6258) );
  OAI21_X1 U7848 ( .B1(n6259), .B2(n8991), .A(n6258), .ZN(P1_U3230) );
  INV_X1 U7849 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6268) );
  INV_X1 U7850 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6296) );
  OAI22_X1 U7851 ( .A1(n5667), .A2(n6343), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6296), .ZN(n6262) );
  NOR2_X1 U7852 ( .A1(n5667), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6261) );
  INV_X1 U7853 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6260) );
  OAI21_X1 U7854 ( .B1(n6261), .B2(n6356), .A(n6260), .ZN(n6355) );
  OAI211_X1 U7855 ( .C1(n6356), .C2(n6262), .A(n6355), .B(P1_STATE_REG_SCAN_IN), .ZN(n6263) );
  NOR2_X1 U7856 ( .A1(n6264), .A2(n6263), .ZN(n6266) );
  AND3_X1 U7857 ( .A1(n9623), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6296), .ZN(n6265) );
  AOI211_X1 U7858 ( .C1(P1_REG3_REG_0__SCAN_IN), .C2(P1_U3084), .A(n6266), .B(
        n6265), .ZN(n6267) );
  OAI21_X1 U7859 ( .B1(n9039), .B2(n6268), .A(n6267), .ZN(P1_U3241) );
  INV_X1 U7860 ( .A(n7780), .ZN(n6300) );
  AOI22_X1 U7861 ( .A1(n9026), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9549), .ZN(n6269) );
  OAI21_X1 U7862 ( .B1(n6300), .B2(n9552), .A(n6269), .ZN(P1_U3335) );
  INV_X1 U7863 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U7864 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6898) );
  MUX2_X1 U7865 ( .A(n6000), .B(P1_REG1_REG_3__SCAN_IN), .S(n6270), .Z(n6272)
         );
  NAND3_X1 U7866 ( .A1(n6272), .A2(n6387), .A3(n6271), .ZN(n6273) );
  NAND3_X1 U7867 ( .A1(n9623), .A2(n6274), .A3(n6273), .ZN(n6275) );
  OAI211_X1 U7868 ( .C1(n9029), .C2(n6276), .A(n6898), .B(n6275), .ZN(n6277)
         );
  INV_X1 U7869 ( .A(n6277), .ZN(n6282) );
  OAI211_X1 U7870 ( .C1(n6280), .C2(n6279), .A(n9616), .B(n6278), .ZN(n6281)
         );
  OAI211_X1 U7871 ( .C1(n6283), .C2(n9039), .A(n6282), .B(n6281), .ZN(P1_U3244) );
  OR2_X1 U7872 ( .A1(n9510), .A2(n6284), .ZN(n6288) );
  AND2_X1 U7873 ( .A1(n6286), .A2(n6285), .ZN(n6287) );
  NOR2_X1 U7874 ( .A1(n6870), .A2(n6661), .ZN(n6289) );
  NAND2_X1 U7875 ( .A1(n7003), .A2(n6881), .ZN(n6290) );
  OR2_X1 U7876 ( .A1(n6291), .A2(n6290), .ZN(n6294) );
  NAND2_X1 U7877 ( .A1(n9309), .A2(n9005), .ZN(n6293) );
  AND2_X1 U7878 ( .A1(n6294), .A2(n6293), .ZN(n6878) );
  OAI21_X1 U7879 ( .B1(n6704), .B2(n6881), .A(n6878), .ZN(n6664) );
  NAND2_X1 U7880 ( .A1(n6664), .A2(n9697), .ZN(n6295) );
  OAI21_X1 U7881 ( .B1(n9697), .B2(n6296), .A(n6295), .ZN(P1_U3523) );
  INV_X1 U7882 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U7883 ( .A1(n6298), .A2(n6297), .ZN(n6299) );
  XNOR2_X1 U7884 ( .A(n6379), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8379) );
  INV_X1 U7885 ( .A(n8379), .ZN(n8369) );
  OAI222_X1 U7886 ( .A1(n8830), .A2(n6301), .B1(n7667), .B2(n6300), .C1(
        P2_U3152), .C2(n8369), .ZN(P2_U3340) );
  AOI21_X1 U7887 ( .B1(n9695), .B2(n6303), .A(n6302), .ZN(n6305) );
  INV_X1 U7888 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9575) );
  AOI22_X1 U7889 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6400), .B1(n6404), .B2(
        n9575), .ZN(n6304) );
  NOR2_X1 U7890 ( .A1(n6305), .A2(n6304), .ZN(n6399) );
  AOI21_X1 U7891 ( .B1(n6305), .B2(n6304), .A(n6399), .ZN(n6315) );
  INV_X1 U7892 ( .A(n9039), .ZN(n9611) );
  NAND2_X1 U7893 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n6404), .ZN(n6306) );
  OAI21_X1 U7894 ( .B1(n6404), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6306), .ZN(
        n6310) );
  AOI21_X1 U7895 ( .B1(n6310), .B2(n6309), .A(n6403), .ZN(n6311) );
  NAND2_X1 U7896 ( .A1(n9616), .A2(n6311), .ZN(n6312) );
  NAND2_X1 U7897 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7657) );
  OAI211_X1 U7898 ( .C1(n9029), .C2(n6400), .A(n6312), .B(n7657), .ZN(n6313)
         );
  AOI21_X1 U7899 ( .B1(n9611), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n6313), .ZN(
        n6314) );
  OAI21_X1 U7900 ( .B1(n6315), .B2(n9030), .A(n6314), .ZN(P1_U3251) );
  INV_X1 U7901 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6328) );
  OAI21_X1 U7902 ( .B1(n6318), .B2(n6317), .A(n6316), .ZN(n6326) );
  AOI21_X1 U7903 ( .B1(n6321), .B2(n6320), .A(n6319), .ZN(n6324) );
  NAND2_X1 U7904 ( .A1(n9610), .A2(n6322), .ZN(n6323) );
  NAND2_X1 U7905 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7559) );
  OAI211_X1 U7906 ( .C1(n6324), .C2(n9030), .A(n6323), .B(n7559), .ZN(n6325)
         );
  AOI21_X1 U7907 ( .B1(n9616), .B2(n6326), .A(n6325), .ZN(n6327) );
  OAI21_X1 U7908 ( .B1(n6328), .B2(n9039), .A(n6327), .ZN(P1_U3249) );
  INV_X1 U7909 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6341) );
  OAI21_X1 U7910 ( .B1(n6331), .B2(n6330), .A(n6329), .ZN(n6339) );
  AOI21_X1 U7911 ( .B1(n6334), .B2(n6333), .A(n6332), .ZN(n6337) );
  NAND2_X1 U7912 ( .A1(n9610), .A2(n6335), .ZN(n6336) );
  NAND2_X1 U7913 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7436) );
  OAI211_X1 U7914 ( .C1(n6337), .C2(n9030), .A(n6336), .B(n7436), .ZN(n6338)
         );
  AOI21_X1 U7915 ( .B1(n9616), .B2(n6339), .A(n6338), .ZN(n6340) );
  OAI21_X1 U7916 ( .B1(n6341), .B2(n9039), .A(n6340), .ZN(P1_U3248) );
  OAI211_X1 U7917 ( .C1(n6344), .C2(n6343), .A(n9616), .B(n6342), .ZN(n6345)
         );
  OAI21_X1 U7918 ( .B1(n9029), .B2(n4927), .A(n6345), .ZN(n6351) );
  INV_X1 U7919 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6349) );
  OAI211_X1 U7920 ( .C1(n6347), .C2(n6346), .A(n9623), .B(n6384), .ZN(n6348)
         );
  OAI21_X1 U7921 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6349), .A(n6348), .ZN(n6350) );
  AOI211_X1 U7922 ( .C1(n9611), .C2(P1_ADDR_REG_1__SCAN_IN), .A(n6351), .B(
        n6350), .ZN(n6352) );
  INV_X1 U7923 ( .A(n6352), .ZN(P1_U3242) );
  MUX2_X1 U7924 ( .A(n6354), .B(n6353), .S(n5667), .Z(n6357) );
  OAI211_X1 U7925 ( .C1(n6357), .C2(n6356), .A(n9004), .B(n6355), .ZN(n6397)
         );
  NAND2_X1 U7926 ( .A1(n4343), .A2(n4273), .ZN(n6358) );
  NAND2_X1 U7927 ( .A1(n6359), .A2(n6358), .ZN(n6360) );
  NAND2_X1 U7928 ( .A1(n9616), .A2(n6360), .ZN(n6366) );
  OAI21_X1 U7929 ( .B1(n6363), .B2(n6362), .A(n6361), .ZN(n6364) );
  AND2_X1 U7930 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7035) );
  AOI21_X1 U7931 ( .B1(n9623), .B2(n6364), .A(n7035), .ZN(n6365) );
  OAI211_X1 U7932 ( .C1(n9029), .C2(n6367), .A(n6366), .B(n6365), .ZN(n6368)
         );
  AOI21_X1 U7933 ( .B1(n9611), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6368), .ZN(
        n6369) );
  NAND2_X1 U7934 ( .A1(n6397), .A2(n6369), .ZN(P1_U3245) );
  NAND2_X1 U7935 ( .A1(n6370), .A2(n6371), .ZN(n6372) );
  XNOR2_X1 U7936 ( .A(n6373), .B(n6372), .ZN(n6377) );
  INV_X1 U7937 ( .A(n8987), .ZN(n8946) );
  INV_X2 U7938 ( .A(n6374), .ZN(n8984) );
  AOI22_X1 U7939 ( .A1(n8946), .A2(n5674), .B1(n8984), .B2(n9003), .ZN(n6376)
         );
  AOI22_X1 U7940 ( .A1(n8989), .A2(n5683), .B1(n8947), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6375) );
  OAI211_X1 U7941 ( .C1(n6377), .C2(n8991), .A(n6376), .B(n6375), .ZN(P1_U3220) );
  INV_X1 U7942 ( .A(n7793), .ZN(n6382) );
  OAI222_X1 U7943 ( .A1(n8830), .A2(n6380), .B1(n7667), .B2(n6382), .C1(n8389), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U7944 ( .A1(P1_U3084), .A2(n9250), .B1(n9552), .B2(n6382), .C1(
        n6381), .C2(n7705), .ZN(P1_U3334) );
  INV_X1 U7945 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7391) );
  INV_X1 U7946 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6389) );
  MUX2_X1 U7947 ( .A(n5996), .B(P1_REG1_REG_2__SCAN_IN), .S(n6396), .Z(n6385)
         );
  NAND3_X1 U7948 ( .A1(n6385), .A2(n6384), .A3(n6383), .ZN(n6386) );
  NAND3_X1 U7949 ( .A1(n9623), .A2(n6387), .A3(n6386), .ZN(n6388) );
  OAI21_X1 U7950 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6389), .A(n6388), .ZN(n6395) );
  OAI211_X1 U7951 ( .C1(n6392), .C2(n6391), .A(n9616), .B(n6390), .ZN(n6393)
         );
  INV_X1 U7952 ( .A(n6393), .ZN(n6394) );
  AOI211_X1 U7953 ( .C1(n9610), .C2(n6396), .A(n6395), .B(n6394), .ZN(n6398)
         );
  OAI211_X1 U7954 ( .C1(n7391), .C2(n9039), .A(n6398), .B(n6397), .ZN(P1_U3243) );
  AOI21_X1 U7955 ( .B1(n9575), .B2(n6400), .A(n6399), .ZN(n6633) );
  INV_X1 U7956 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9605) );
  NOR2_X1 U7957 ( .A1(n9605), .A2(n6408), .ZN(n6632) );
  AOI21_X1 U7958 ( .B1(n9605), .B2(n6408), .A(n6632), .ZN(n6401) );
  XNOR2_X1 U7959 ( .A(n6633), .B(n6401), .ZN(n6412) );
  NOR2_X1 U7960 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6641), .ZN(n6402) );
  AOI21_X1 U7961 ( .B1(n6641), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6402), .ZN(
        n6406) );
  OAI21_X1 U7962 ( .B1(n6406), .B2(n6405), .A(n6640), .ZN(n6410) );
  NAND2_X1 U7963 ( .A1(n9611), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U7964 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7671) );
  OAI211_X1 U7965 ( .C1(n9029), .C2(n6408), .A(n6407), .B(n7671), .ZN(n6409)
         );
  AOI21_X1 U7966 ( .B1(n9616), .B2(n6410), .A(n6409), .ZN(n6411) );
  OAI21_X1 U7967 ( .B1(n6412), .B2(n9030), .A(n6411), .ZN(P1_U3252) );
  XNOR2_X1 U7968 ( .A(n7354), .B(P2_B_REG_SCAN_IN), .ZN(n6413) );
  NAND2_X1 U7969 ( .A1(n7469), .A2(n7569), .ZN(n9817) );
  OAI21_X1 U7970 ( .B1(P2_D_REG_1__SCAN_IN), .B2(n6433), .A(n9817), .ZN(n7157)
         );
  NAND2_X1 U7971 ( .A1(n6679), .A2(n6483), .ZN(n6419) );
  NAND2_X1 U7972 ( .A1(n6480), .A2(n6419), .ZN(n6671) );
  INV_X1 U7973 ( .A(n6671), .ZN(n7155) );
  AND2_X1 U7974 ( .A1(n6470), .A2(n6456), .ZN(n6420) );
  NAND4_X1 U7975 ( .A1(n7157), .A2(n7154), .A3(n7155), .A4(n6674), .ZN(n6432)
         );
  NOR4_X1 U7976 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(n6422), .ZN(n6431) );
  NOR4_X1 U7977 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n6423) );
  NAND3_X1 U7978 ( .A1(n6423), .A2(n9795), .A3(n9797), .ZN(n6429) );
  NOR4_X1 U7979 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6427) );
  NOR4_X1 U7980 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6426) );
  NOR4_X1 U7981 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n6425) );
  NOR4_X1 U7982 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6424) );
  NAND4_X1 U7983 ( .A1(n6427), .A2(n6426), .A3(n6425), .A4(n6424), .ZN(n6428)
         );
  NOR4_X1 U7984 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        n6429), .A4(n6428), .ZN(n6430) );
  NAND2_X1 U7985 ( .A1(n7354), .A2(n7569), .ZN(n9815) );
  INV_X1 U7986 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6434) );
  NAND2_X1 U7987 ( .A1(n9783), .A2(n6434), .ZN(n6435) );
  INV_X1 U7988 ( .A(n7153), .ZN(n6436) );
  INV_X2 U7989 ( .A(n9895), .ZN(n9872) );
  INV_X1 U7990 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6475) );
  NAND2_X1 U7991 ( .A1(n7916), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U7992 ( .A1(n6462), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U7993 ( .A1(n6463), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6438) );
  NAND2_X1 U7994 ( .A1(n6750), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6437) );
  INV_X1 U7995 ( .A(SI_0_), .ZN(n6444) );
  NOR2_X1 U7996 ( .A1(n6445), .A2(n6444), .ZN(n6446) );
  XNOR2_X1 U7997 ( .A(n6446), .B(n4535), .ZN(n8831) );
  AND2_X1 U7998 ( .A1(n6453), .A2(n9821), .ZN(n6680) );
  INV_X1 U7999 ( .A(n6680), .ZN(n6448) );
  NAND2_X1 U8000 ( .A1(n6447), .A2(n6448), .ZN(n6762) );
  OAI21_X1 U8001 ( .B1(n6447), .B2(n6448), .A(n6762), .ZN(n7171) );
  INV_X1 U8002 ( .A(n7171), .ZN(n6473) );
  NAND2_X1 U8003 ( .A1(n6449), .A2(n6421), .ZN(n7161) );
  NAND2_X1 U8004 ( .A1(n7161), .A2(n6470), .ZN(n6451) );
  AND2_X1 U8005 ( .A1(n6676), .A2(n8389), .ZN(n6450) );
  NAND2_X1 U8006 ( .A1(n6451), .A2(n6450), .ZN(n9757) );
  INV_X1 U8007 ( .A(n6453), .ZN(n9705) );
  NAND2_X1 U8008 ( .A1(n9705), .A2(n9821), .ZN(n6454) );
  INV_X1 U8009 ( .A(n8170), .ZN(n6458) );
  INV_X1 U8010 ( .A(n6454), .ZN(n6455) );
  NAND2_X1 U8011 ( .A1(n6447), .A2(n6455), .ZN(n6457) );
  OR2_X1 U8012 ( .A1(n6449), .A2(n6877), .ZN(n8117) );
  INV_X1 U8013 ( .A(n6470), .ZN(n8307) );
  OAI211_X1 U8014 ( .C1(n8162), .C2(n6458), .A(n6457), .B(n9769), .ZN(n6469)
         );
  INV_X1 U8015 ( .A(n6460), .ZN(n6461) );
  NAND2_X1 U8016 ( .A1(n6462), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U8017 ( .A1(n7916), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U8018 ( .A1(n6463), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U8019 ( .A1(n6483), .A2(n6460), .ZN(n8694) );
  AOI22_X1 U8020 ( .A1(n9762), .A2(n6453), .B1(n8318), .B2(n9764), .ZN(n6468)
         );
  NAND2_X1 U8021 ( .A1(n6469), .A2(n6468), .ZN(n7166) );
  INV_X1 U8022 ( .A(n7166), .ZN(n6472) );
  AOI21_X1 U8023 ( .B1(n9821), .B2(n6734), .A(n4554), .ZN(n7167) );
  AOI22_X1 U8024 ( .A1(n7167), .A2(n9836), .B1(n9835), .B2(n6734), .ZN(n6471)
         );
  OAI211_X1 U8025 ( .C1(n6473), .C2(n8796), .A(n6472), .B(n6471), .ZN(n6477)
         );
  NAND2_X1 U8026 ( .A1(n9872), .A2(n6477), .ZN(n6474) );
  OAI21_X1 U8027 ( .B1(n9872), .B2(n6475), .A(n6474), .ZN(P2_U3454) );
  INV_X1 U8028 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6479) );
  NAND2_X1 U8029 ( .A1(n4260), .A2(n6477), .ZN(n6478) );
  OAI21_X1 U8030 ( .B1(n4260), .B2(n6479), .A(n6478), .ZN(P2_U3521) );
  INV_X1 U8031 ( .A(n6480), .ZN(n6481) );
  NAND2_X1 U8032 ( .A1(n6481), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6482) );
  OAI211_X1 U8033 ( .C1(n9782), .C2(n6483), .A(n8309), .B(n6482), .ZN(n6514)
         );
  NAND2_X1 U8034 ( .A1(n6514), .A2(n6768), .ZN(n6484) );
  NAND2_X1 U8035 ( .A1(n6484), .A2(n8319), .ZN(n8384) );
  NOR2_X1 U8036 ( .A1(n7453), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6507) );
  NAND2_X1 U8037 ( .A1(n7313), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6504) );
  INV_X1 U8038 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6485) );
  MUX2_X1 U8039 ( .A(n6485), .B(P2_REG2_REG_10__SCAN_IN), .S(n7313), .Z(n6486)
         );
  INV_X1 U8040 ( .A(n6486), .ZN(n6555) );
  NAND2_X1 U8041 ( .A1(n7286), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6503) );
  INV_X1 U8042 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6487) );
  MUX2_X1 U8043 ( .A(n6487), .B(P2_REG2_REG_9__SCAN_IN), .S(n7286), .Z(n6488)
         );
  INV_X1 U8044 ( .A(n6488), .ZN(n6629) );
  INV_X1 U8045 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6502) );
  MUX2_X1 U8046 ( .A(n6502), .B(P2_REG2_REG_8__SCAN_IN), .S(n7112), .Z(n6588)
         );
  NAND2_X1 U8047 ( .A1(n6526), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6501) );
  INV_X1 U8048 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6489) );
  MUX2_X1 U8049 ( .A(n6489), .B(P2_REG2_REG_7__SCAN_IN), .S(n6526), .Z(n6490)
         );
  INV_X1 U8050 ( .A(n6490), .ZN(n6545) );
  NAND2_X1 U8051 ( .A1(n6524), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6500) );
  INV_X1 U8052 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6491) );
  MUX2_X1 U8053 ( .A(n6491), .B(P2_REG2_REG_6__SCAN_IN), .S(n6524), .Z(n6492)
         );
  INV_X1 U8054 ( .A(n6492), .ZN(n6608) );
  NAND2_X1 U8055 ( .A1(n6522), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6499) );
  INV_X1 U8056 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6493) );
  MUX2_X1 U8057 ( .A(n6493), .B(P2_REG2_REG_5__SCAN_IN), .S(n6522), .Z(n6494)
         );
  INV_X1 U8058 ( .A(n6494), .ZN(n6578) );
  NAND2_X1 U8059 ( .A1(n6520), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6498) );
  INV_X1 U8060 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6495) );
  MUX2_X1 U8061 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6495), .S(n6520), .Z(n6598)
         );
  NAND2_X1 U8062 ( .A1(n6518), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6497) );
  INV_X1 U8063 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6496) );
  MUX2_X1 U8064 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6496), .S(n6518), .Z(n6619)
         );
  INV_X1 U8065 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7237) );
  MUX2_X1 U8066 ( .A(n7237), .B(P2_REG2_REG_2__SCAN_IN), .S(n6728), .Z(n9562)
         );
  INV_X1 U8067 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7163) );
  MUX2_X1 U8068 ( .A(n7163), .B(P2_REG2_REG_1__SCAN_IN), .S(n6571), .Z(n6567)
         );
  NAND3_X1 U8069 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n6567), .ZN(n6566) );
  OAI21_X1 U8070 ( .B1(n6571), .B2(n7163), .A(n6566), .ZN(n9563) );
  NAND2_X1 U8071 ( .A1(n9562), .A2(n9563), .ZN(n9561) );
  OAI21_X1 U8072 ( .B1(n6728), .B2(n7237), .A(n9561), .ZN(n6618) );
  NAND2_X1 U8073 ( .A1(n6619), .A2(n6618), .ZN(n6617) );
  NAND2_X1 U8074 ( .A1(n6497), .A2(n6617), .ZN(n6599) );
  NAND2_X1 U8075 ( .A1(n6598), .A2(n6599), .ZN(n6597) );
  NAND2_X1 U8076 ( .A1(n6498), .A2(n6597), .ZN(n6579) );
  NAND2_X1 U8077 ( .A1(n6578), .A2(n6579), .ZN(n6577) );
  NAND2_X1 U8078 ( .A1(n6499), .A2(n6577), .ZN(n6609) );
  NAND2_X1 U8079 ( .A1(n6608), .A2(n6609), .ZN(n6607) );
  NAND2_X1 U8080 ( .A1(n6500), .A2(n6607), .ZN(n6546) );
  NAND2_X1 U8081 ( .A1(n6545), .A2(n6546), .ZN(n6544) );
  NAND2_X1 U8082 ( .A1(n6501), .A2(n6544), .ZN(n6589) );
  NAND2_X1 U8083 ( .A1(n6588), .A2(n6589), .ZN(n6587) );
  OAI21_X1 U8084 ( .B1(n7112), .B2(n6502), .A(n6587), .ZN(n6628) );
  NAND2_X1 U8085 ( .A1(n6629), .A2(n6628), .ZN(n6627) );
  NAND2_X1 U8086 ( .A1(n6503), .A2(n6627), .ZN(n6556) );
  NAND2_X1 U8087 ( .A1(n6555), .A2(n6556), .ZN(n6554) );
  NAND2_X1 U8088 ( .A1(n6504), .A2(n6554), .ZN(n6788) );
  INV_X1 U8089 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6505) );
  MUX2_X1 U8090 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n6505), .S(n7453), .Z(n6506)
         );
  INV_X1 U8091 ( .A(n6506), .ZN(n6787) );
  NOR2_X1 U8092 ( .A1(n6788), .A2(n6787), .ZN(n6786) );
  NOR2_X1 U8093 ( .A1(n6507), .A2(n6786), .ZN(n6512) );
  INV_X1 U8094 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6508) );
  MUX2_X1 U8095 ( .A(n6508), .B(P2_REG2_REG_12__SCAN_IN), .S(n7539), .Z(n6509)
         );
  INV_X1 U8096 ( .A(n6509), .ZN(n6511) );
  NOR2_X1 U8097 ( .A1(n6460), .A2(n8828), .ZN(n6510) );
  NAND2_X1 U8098 ( .A1(n6511), .A2(n6512), .ZN(n6797) );
  OAI211_X1 U8099 ( .C1(n6512), .C2(n6511), .A(n9714), .B(n6797), .ZN(n6538)
         );
  AND2_X1 U8100 ( .A1(n6768), .A2(n8828), .ZN(n6513) );
  INV_X1 U8101 ( .A(n6728), .ZN(n9559) );
  INV_X1 U8102 ( .A(n6571), .ZN(n6515) );
  NAND2_X1 U8103 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n6562) );
  INV_X1 U8104 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6516) );
  MUX2_X1 U8105 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6516), .S(n6728), .Z(n9556)
         );
  NOR2_X1 U8106 ( .A1(n9557), .A2(n9556), .ZN(n9555) );
  AOI21_X1 U8107 ( .B1(n9559), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9555), .ZN(
        n6614) );
  NAND2_X1 U8108 ( .A1(n6518), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6517) );
  OAI21_X1 U8109 ( .B1(n6518), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6517), .ZN(
        n6613) );
  NOR2_X1 U8110 ( .A1(n6614), .A2(n6613), .ZN(n6612) );
  AOI21_X1 U8111 ( .B1(n6518), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6612), .ZN(
        n6594) );
  NAND2_X1 U8112 ( .A1(n6520), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6519) );
  OAI21_X1 U8113 ( .B1(n6520), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6519), .ZN(
        n6593) );
  NOR2_X1 U8114 ( .A1(n6594), .A2(n6593), .ZN(n6592) );
  AOI21_X1 U8115 ( .B1(n6520), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6592), .ZN(
        n6574) );
  NAND2_X1 U8116 ( .A1(n6522), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6521) );
  OAI21_X1 U8117 ( .B1(n6522), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6521), .ZN(
        n6573) );
  NAND2_X1 U8118 ( .A1(n6524), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6523) );
  OAI21_X1 U8119 ( .B1(n6524), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6523), .ZN(
        n6603) );
  NAND2_X1 U8120 ( .A1(n6526), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6525) );
  OAI21_X1 U8121 ( .B1(n6526), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6525), .ZN(
        n6541) );
  NOR2_X1 U8122 ( .A1(n4288), .A2(n6541), .ZN(n6540) );
  INV_X1 U8123 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6527) );
  MUX2_X1 U8124 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6527), .S(n7112), .Z(n6583)
         );
  NAND2_X1 U8125 ( .A1(n7286), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6528) );
  OAI21_X1 U8126 ( .B1(n7286), .B2(P2_REG1_REG_9__SCAN_IN), .A(n6528), .ZN(
        n6623) );
  INV_X1 U8127 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6529) );
  MUX2_X1 U8128 ( .A(n6529), .B(P2_REG1_REG_10__SCAN_IN), .S(n7313), .Z(n6550)
         );
  NOR2_X1 U8129 ( .A1(n6551), .A2(n6550), .ZN(n6549) );
  AOI21_X1 U8130 ( .B1(n7313), .B2(P2_REG1_REG_10__SCAN_IN), .A(n6549), .ZN(
        n6791) );
  INV_X1 U8131 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6530) );
  MUX2_X1 U8132 ( .A(n6530), .B(P2_REG1_REG_11__SCAN_IN), .S(n7453), .Z(n6790)
         );
  NOR2_X1 U8133 ( .A1(n6791), .A2(n6790), .ZN(n6789) );
  MUX2_X1 U8134 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n9911), .S(n7539), .Z(n6531)
         );
  OAI21_X1 U8135 ( .B1(n6532), .B2(n6531), .A(n6804), .ZN(n6536) );
  NOR2_X1 U8136 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7546), .ZN(n6535) );
  INV_X1 U8137 ( .A(n9715), .ZN(n6808) );
  INV_X1 U8138 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6533) );
  NOR2_X1 U8139 ( .A1(n6808), .A2(n6533), .ZN(n6534) );
  AOI211_X1 U8140 ( .C1(n9713), .C2(n6536), .A(n6535), .B(n6534), .ZN(n6537)
         );
  OAI211_X1 U8141 ( .C1(n9717), .C2(n6539), .A(n6538), .B(n6537), .ZN(P2_U3257) );
  AND2_X1 U8142 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6543) );
  AOI211_X1 U8143 ( .C1(n4288), .C2(n6541), .A(n6540), .B(n9718), .ZN(n6542)
         );
  AOI211_X1 U8144 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n9715), .A(n6543), .B(
        n6542), .ZN(n6548) );
  OAI211_X1 U8145 ( .C1(n6546), .C2(n6545), .A(n9714), .B(n6544), .ZN(n6547)
         );
  OAI211_X1 U8146 ( .C1(n9717), .C2(n7134), .A(n6548), .B(n6547), .ZN(P2_U3252) );
  NAND2_X1 U8147 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7325) );
  INV_X1 U8148 ( .A(n7325), .ZN(n6553) );
  AOI211_X1 U8149 ( .C1(n6551), .C2(n6550), .A(n6549), .B(n9718), .ZN(n6552)
         );
  AOI211_X1 U8150 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n9715), .A(n6553), .B(
        n6552), .ZN(n6558) );
  OAI211_X1 U8151 ( .C1(n6556), .C2(n6555), .A(n9714), .B(n6554), .ZN(n6557)
         );
  OAI211_X1 U8152 ( .C1(n9717), .C2(n6559), .A(n6558), .B(n6557), .ZN(P2_U3255) );
  AOI211_X1 U8153 ( .C1(n6562), .C2(n6561), .A(n6560), .B(n9718), .ZN(n6563)
         );
  AOI211_X1 U8154 ( .C1(P2_ADDR_REG_1__SCAN_IN), .C2(n9715), .A(n6564), .B(
        n6563), .ZN(n6570) );
  INV_X1 U8155 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6565) );
  INV_X1 U8156 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7207) );
  NOR2_X1 U8157 ( .A1(n6565), .A2(n7207), .ZN(n6568) );
  OAI211_X1 U8158 ( .C1(n6568), .C2(n6567), .A(n9714), .B(n6566), .ZN(n6569)
         );
  OAI211_X1 U8159 ( .C1(n9717), .C2(n6571), .A(n6570), .B(n6569), .ZN(P2_U3246) );
  INV_X1 U8160 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6824) );
  NOR2_X1 U8161 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6824), .ZN(n6576) );
  AOI211_X1 U8162 ( .C1(n6574), .C2(n6573), .A(n6572), .B(n9718), .ZN(n6575)
         );
  AOI211_X1 U8163 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n9715), .A(n6576), .B(
        n6575), .ZN(n6581) );
  OAI211_X1 U8164 ( .C1(n6579), .C2(n6578), .A(n9714), .B(n6577), .ZN(n6580)
         );
  OAI211_X1 U8165 ( .C1(n9717), .C2(n6834), .A(n6581), .B(n6580), .ZN(P2_U3250) );
  NAND2_X1 U8166 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7121) );
  INV_X1 U8167 ( .A(n7121), .ZN(n6586) );
  AOI211_X1 U8168 ( .C1(n6584), .C2(n6583), .A(n6582), .B(n9718), .ZN(n6585)
         );
  AOI211_X1 U8169 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n9715), .A(n6586), .B(
        n6585), .ZN(n6591) );
  OAI211_X1 U8170 ( .C1(n6589), .C2(n6588), .A(n9714), .B(n6587), .ZN(n6590)
         );
  OAI211_X1 U8171 ( .C1(n9717), .C2(n7112), .A(n6591), .B(n6590), .ZN(P2_U3253) );
  AND2_X1 U8172 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6596) );
  AOI211_X1 U8173 ( .C1(n6594), .C2(n6593), .A(n6592), .B(n9718), .ZN(n6595)
         );
  AOI211_X1 U8174 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n9715), .A(n6596), .B(
        n6595), .ZN(n6601) );
  OAI211_X1 U8175 ( .C1(n6599), .C2(n6598), .A(n9714), .B(n6597), .ZN(n6600)
         );
  OAI211_X1 U8176 ( .C1(n9717), .C2(n6821), .A(n6601), .B(n6600), .ZN(P2_U3249) );
  NAND2_X1 U8177 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n6943) );
  INV_X1 U8178 ( .A(n6943), .ZN(n6606) );
  AOI211_X1 U8179 ( .C1(n6604), .C2(n6603), .A(n6602), .B(n9718), .ZN(n6605)
         );
  AOI211_X1 U8180 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n9715), .A(n6606), .B(
        n6605), .ZN(n6611) );
  OAI211_X1 U8181 ( .C1(n6609), .C2(n6608), .A(n9714), .B(n6607), .ZN(n6610)
         );
  OAI211_X1 U8182 ( .C1(n9717), .C2(n6930), .A(n6611), .B(n6610), .ZN(P2_U3251) );
  NOR2_X1 U8183 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6749), .ZN(n6616) );
  AOI211_X1 U8184 ( .C1(n6614), .C2(n6613), .A(n6612), .B(n9718), .ZN(n6615)
         );
  AOI211_X1 U8185 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n9715), .A(n6616), .B(
        n6615), .ZN(n6621) );
  OAI211_X1 U8186 ( .C1(n6619), .C2(n6618), .A(n9714), .B(n6617), .ZN(n6620)
         );
  OAI211_X1 U8187 ( .C1(n9717), .C2(n6767), .A(n6621), .B(n6620), .ZN(P2_U3248) );
  NAND2_X1 U8188 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7304) );
  INV_X1 U8189 ( .A(n7304), .ZN(n6626) );
  AOI211_X1 U8190 ( .C1(n6624), .C2(n6623), .A(n6622), .B(n9718), .ZN(n6625)
         );
  AOI211_X1 U8191 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n9715), .A(n6626), .B(
        n6625), .ZN(n6631) );
  OAI211_X1 U8192 ( .C1(n6629), .C2(n6628), .A(n9714), .B(n6627), .ZN(n6630)
         );
  OAI211_X1 U8193 ( .C1(n9717), .C2(n4449), .A(n6631), .B(n6630), .ZN(P2_U3254) );
  NAND2_X1 U8194 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8926) );
  XOR2_X1 U8195 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6954), .Z(n6635) );
  XOR2_X1 U8196 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6642), .Z(n6650) );
  OAI22_X1 U8197 ( .A1(n6633), .A2(n6632), .B1(n6641), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n6651) );
  NAND2_X1 U8198 ( .A1(n6650), .A2(n6651), .ZN(n6649) );
  OAI21_X1 U8199 ( .B1(n6642), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6649), .ZN(
        n6634) );
  NAND2_X1 U8200 ( .A1(n6635), .A2(n6634), .ZN(n6948) );
  OAI21_X1 U8201 ( .B1(n6635), .B2(n6634), .A(n6948), .ZN(n6636) );
  NAND2_X1 U8202 ( .A1(n9623), .A2(n6636), .ZN(n6637) );
  OAI211_X1 U8203 ( .C1(n9029), .C2(n6638), .A(n8926), .B(n6637), .ZN(n6647)
         );
  NAND2_X1 U8204 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6642), .ZN(n6639) );
  OAI21_X1 U8205 ( .B1(n6642), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6639), .ZN(
        n6655) );
  OAI21_X1 U8206 ( .B1(n6641), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6640), .ZN(
        n6656) );
  NOR2_X1 U8207 ( .A1(n6655), .A2(n6656), .ZN(n6654) );
  AOI21_X1 U8208 ( .B1(n6642), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6654), .ZN(
        n6645) );
  NAND2_X1 U8209 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n6954), .ZN(n6643) );
  OAI21_X1 U8210 ( .B1(n6954), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6643), .ZN(
        n6644) );
  NOR2_X1 U8211 ( .A1(n6645), .A2(n6644), .ZN(n6953) );
  AOI211_X1 U8212 ( .C1(n6645), .C2(n6644), .A(n6953), .B(n9017), .ZN(n6646)
         );
  AOI211_X1 U8213 ( .C1(P1_ADDR_REG_13__SCAN_IN), .C2(n9611), .A(n6647), .B(
        n6646), .ZN(n6648) );
  INV_X1 U8214 ( .A(n6648), .ZN(P1_U3254) );
  OAI21_X1 U8215 ( .B1(n6651), .B2(n6650), .A(n6649), .ZN(n6659) );
  NAND2_X1 U8216 ( .A1(n9611), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6652) );
  NAND2_X1 U8217 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8877) );
  OAI211_X1 U8218 ( .C1(n9029), .C2(n6653), .A(n6652), .B(n8877), .ZN(n6658)
         );
  AOI211_X1 U8219 ( .C1(n6656), .C2(n6655), .A(n6654), .B(n9017), .ZN(n6657)
         );
  AOI211_X1 U8220 ( .C1(n6659), .C2(n9623), .A(n6658), .B(n6657), .ZN(n6660)
         );
  INV_X1 U8221 ( .A(n6660), .ZN(P1_U3253) );
  INV_X1 U8222 ( .A(n6661), .ZN(n9533) );
  INV_X1 U8223 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U8224 ( .A1(n6664), .A2(n9530), .ZN(n6665) );
  OAI21_X1 U8225 ( .B1(n9530), .B2(n6666), .A(n6665), .ZN(P1_U3454) );
  OR2_X1 U8226 ( .A1(n7157), .A2(n7153), .ZN(n6667) );
  NOR2_X1 U8227 ( .A1(n7158), .A2(n6667), .ZN(n6669) );
  INV_X1 U8228 ( .A(n9782), .ZN(n8305) );
  INV_X1 U8229 ( .A(n6679), .ZN(n8304) );
  NAND2_X1 U8230 ( .A1(n6678), .A2(n8304), .ZN(n8071) );
  NOR2_X1 U8231 ( .A1(n8071), .A2(n8694), .ZN(n7986) );
  INV_X1 U8232 ( .A(n6669), .ZN(n6673) );
  INV_X1 U8233 ( .A(n6670), .ZN(n6672) );
  AOI211_X1 U8234 ( .C1(n6673), .C2(n6674), .A(n6672), .B(n6671), .ZN(n6941)
         );
  AND2_X1 U8235 ( .A1(n6941), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9712) );
  INV_X1 U8236 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7206) );
  OAI22_X1 U8237 ( .A1(n9703), .A2(n6668), .B1(n9712), .B2(n7206), .ZN(n6685)
         );
  NOR2_X1 U8238 ( .A1(n6449), .A2(n6729), .ZN(n7164) );
  NAND2_X1 U8239 ( .A1(n6678), .A2(n7164), .ZN(n6675) );
  INV_X1 U8240 ( .A(n9821), .ZN(n8160) );
  AND2_X1 U8241 ( .A1(n9887), .A2(n6676), .ZN(n6677) );
  NAND2_X1 U8242 ( .A1(n6680), .A2(n6739), .ZN(n6732) );
  NAND2_X1 U8243 ( .A1(n6453), .A2(n8118), .ZN(n6681) );
  NAND2_X1 U8244 ( .A1(n6681), .A2(n8160), .ZN(n6682) );
  NAND2_X1 U8245 ( .A1(n6732), .A2(n6682), .ZN(n6683) );
  OAI22_X1 U8246 ( .A1(n9701), .A2(n8160), .B1(n8085), .B2(n6683), .ZN(n6684)
         );
  OR2_X1 U8247 ( .A1(n6685), .A2(n6684), .ZN(P2_U3234) );
  INV_X1 U8248 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6697) );
  AOI21_X1 U8249 ( .B1(n6688), .B2(n6687), .A(n6686), .ZN(n6689) );
  NAND2_X1 U8250 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7378) );
  OAI21_X1 U8251 ( .B1(n9030), .B2(n6689), .A(n7378), .ZN(n6694) );
  AOI211_X1 U8252 ( .C1(n6692), .C2(n6691), .A(n6690), .B(n9017), .ZN(n6693)
         );
  AOI211_X1 U8253 ( .C1(n9610), .C2(n6695), .A(n6694), .B(n6693), .ZN(n6696)
         );
  OAI21_X1 U8254 ( .B1(n9039), .B2(n6697), .A(n6696), .ZN(P1_U3247) );
  INV_X1 U8255 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6723) );
  INV_X1 U8256 ( .A(n9510), .ZN(n9687) );
  NAND2_X1 U8257 ( .A1(n6698), .A2(n9664), .ZN(n6700) );
  NAND2_X1 U8258 ( .A1(n5674), .A2(n6883), .ZN(n6857) );
  NAND2_X1 U8259 ( .A1(n6702), .A2(n6701), .ZN(n6962) );
  OR2_X1 U8260 ( .A1(n6702), .A2(n6701), .ZN(n6703) );
  NAND2_X1 U8261 ( .A1(n6962), .A2(n6703), .ZN(n7083) );
  NAND3_X1 U8262 ( .A1(n9664), .A2(n6960), .A3(n6704), .ZN(n7047) );
  NAND2_X1 U8263 ( .A1(n9664), .A2(n6704), .ZN(n6705) );
  NAND2_X1 U8264 ( .A1(n8948), .A2(n6705), .ZN(n6706) );
  NAND2_X1 U8265 ( .A1(n7047), .A2(n6706), .ZN(n7079) );
  NAND2_X1 U8266 ( .A1(n9568), .A2(n8948), .ZN(n6708) );
  OAI21_X1 U8267 ( .B1(n7079), .B2(n9682), .A(n6708), .ZN(n6721) );
  INV_X1 U8268 ( .A(n9643), .ZN(n9376) );
  NAND2_X1 U8269 ( .A1(n7083), .A2(n9376), .ZN(n6720) );
  XNOR2_X1 U8270 ( .A(n6711), .B(n6710), .ZN(n6715) );
  NAND2_X1 U8271 ( .A1(n6712), .A2(n9207), .ZN(n6714) );
  OR2_X1 U8272 ( .A1(n5670), .A2(n6759), .ZN(n6713) );
  NAND2_X1 U8273 ( .A1(n6715), .A2(n9640), .ZN(n6719) );
  AOI22_X1 U8274 ( .A1(n9002), .A2(n9309), .B1(n9311), .B2(n9005), .ZN(n6718)
         );
  NAND3_X1 U8275 ( .A1(n6720), .A2(n6719), .A3(n6718), .ZN(n7080) );
  AOI211_X1 U8276 ( .C1(n9687), .C2(n7083), .A(n6721), .B(n7080), .ZN(n6887)
         );
  OR2_X1 U8277 ( .A1(n6887), .A2(n9688), .ZN(n6722) );
  OAI21_X1 U8278 ( .B1(n9530), .B2(n6723), .A(n6722), .ZN(P1_U3460) );
  OR2_X1 U8279 ( .A1(n6815), .A2(n6725), .ZN(n6726) );
  NAND3_X1 U8280 ( .A1(n6730), .A2(n6729), .A3(n6877), .ZN(n6731) );
  NAND2_X2 U8281 ( .A1(n7161), .A2(n6731), .ZN(n6912) );
  OR2_X1 U8282 ( .A1(n9821), .A2(n6912), .ZN(n6733) );
  XNOR2_X1 U8283 ( .A(n6734), .B(n6912), .ZN(n6735) );
  NAND2_X1 U8284 ( .A1(n8320), .A2(n6739), .ZN(n6736) );
  XNOR2_X1 U8285 ( .A(n6735), .B(n6736), .ZN(n9699) );
  INV_X1 U8286 ( .A(n6735), .ZN(n6737) );
  NAND2_X1 U8287 ( .A1(n6737), .A2(n6736), .ZN(n6738) );
  XNOR2_X1 U8288 ( .A(n6919), .B(n9827), .ZN(n6743) );
  INV_X1 U8289 ( .A(n6743), .ZN(n6741) );
  NAND2_X1 U8290 ( .A1(n8318), .A2(n6739), .ZN(n6742) );
  INV_X1 U8291 ( .A(n6742), .ZN(n6740) );
  NAND2_X1 U8292 ( .A1(n6743), .A2(n6742), .ZN(n6744) );
  NAND2_X1 U8293 ( .A1(n6746), .A2(n6745), .ZN(n6747) );
  NAND2_X1 U8294 ( .A1(n6904), .A2(n6747), .ZN(n6748) );
  OAI22_X1 U8295 ( .A1(n9701), .A2(n6763), .B1(n6748), .B2(n8085), .ZN(n6756)
         );
  NAND2_X1 U8296 ( .A1(n8105), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6754) );
  INV_X1 U8297 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6749) );
  NAND2_X1 U8298 ( .A1(n7141), .A2(n6749), .ZN(n6753) );
  NAND2_X1 U8299 ( .A1(n6750), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6752) );
  NAND2_X1 U8300 ( .A1(n6463), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6751) );
  NAND4_X2 U8301 ( .A1(n6754), .A2(n6753), .A3(n6752), .A4(n6751), .ZN(n8317)
         );
  INV_X1 U8302 ( .A(n8317), .ZN(n6839) );
  INV_X1 U8303 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7238) );
  OAI22_X1 U8304 ( .A1(n9703), .A2(n6839), .B1(n7238), .B2(n9712), .ZN(n6755)
         );
  AOI211_X1 U8305 ( .C1(n7985), .C2(n8320), .A(n6756), .B(n6755), .ZN(n6757)
         );
  INV_X1 U8306 ( .A(n6757), .ZN(P2_U3239) );
  INV_X1 U8307 ( .A(n7808), .ZN(n6991) );
  OAI222_X1 U8308 ( .A1(n6759), .A2(P1_U3084), .B1(n9552), .B2(n6991), .C1(
        n6758), .C2(n7705), .ZN(P1_U3333) );
  INV_X1 U8309 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6782) );
  INV_X1 U8310 ( .A(n9856), .ZN(n9878) );
  NAND2_X1 U8311 ( .A1(n6668), .A2(n6760), .ZN(n6761) );
  NAND2_X1 U8312 ( .A1(n6763), .A2(n8318), .ZN(n8173) );
  NAND2_X1 U8313 ( .A1(n7233), .A2(n8120), .ZN(n7232) );
  NAND2_X1 U8314 ( .A1(n9702), .A2(n6763), .ZN(n6764) );
  NAND2_X1 U8315 ( .A1(n7232), .A2(n6764), .ZN(n6769) );
  NAND2_X1 U8316 ( .A1(n6769), .A2(n6837), .ZN(n6814) );
  OR2_X1 U8317 ( .A1(n6769), .A2(n6837), .ZN(n6770) );
  NAND2_X1 U8318 ( .A1(n6814), .A2(n6770), .ZN(n7198) );
  AND2_X1 U8319 ( .A1(n7234), .A2(n7204), .ZN(n6771) );
  OR2_X1 U8320 ( .A1(n6771), .A2(n7261), .ZN(n7195) );
  OAI22_X1 U8321 ( .A1(n7195), .A2(n9889), .B1(n8147), .B2(n9887), .ZN(n6780)
         );
  NAND2_X1 U8322 ( .A1(n8162), .A2(n8170), .ZN(n7226) );
  NAND2_X1 U8323 ( .A1(n7228), .A2(n8171), .ZN(n6838) );
  XNOR2_X1 U8324 ( .A(n6838), .B(n6837), .ZN(n6779) );
  INV_X1 U8325 ( .A(n9757), .ZN(n7344) );
  NAND2_X1 U8326 ( .A1(n7198), .A2(n7344), .ZN(n6778) );
  NAND2_X1 U8327 ( .A1(n8105), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6776) );
  NAND2_X1 U8328 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6825) );
  OAI21_X1 U8329 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n6825), .ZN(n7265) );
  INV_X1 U8330 ( .A(n7265), .ZN(n6772) );
  NAND2_X1 U8331 ( .A1(n7141), .A2(n6772), .ZN(n6775) );
  NAND2_X1 U8332 ( .A1(n6750), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6774) );
  NAND2_X1 U8333 ( .A1(n6463), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6773) );
  NAND4_X1 U8334 ( .A1(n6776), .A2(n6775), .A3(n6774), .A4(n6773), .ZN(n8316)
         );
  AOI22_X1 U8335 ( .A1(n9762), .A2(n8318), .B1(n8316), .B2(n9764), .ZN(n6777)
         );
  OAI211_X1 U8336 ( .C1(n8690), .C2(n6779), .A(n6778), .B(n6777), .ZN(n7199)
         );
  AOI211_X1 U8337 ( .C1(n9878), .C2(n7198), .A(n6780), .B(n7199), .ZN(n6783)
         );
  OR2_X1 U8338 ( .A1(n6783), .A2(n9910), .ZN(n6781) );
  OAI21_X1 U8339 ( .B1(n4260), .B2(n6782), .A(n6781), .ZN(P2_U3523) );
  INV_X1 U8340 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6785) );
  OR2_X1 U8341 ( .A1(n6783), .A2(n9895), .ZN(n6784) );
  OAI21_X1 U8342 ( .B1(n9872), .B2(n6785), .A(n6784), .ZN(P2_U3460) );
  AOI21_X1 U8343 ( .B1(n6788), .B2(n6787), .A(n6786), .ZN(n6796) );
  INV_X1 U8344 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7463) );
  NOR2_X1 U8345 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7463), .ZN(n6793) );
  AOI211_X1 U8346 ( .C1(n6791), .C2(n6790), .A(n6789), .B(n9718), .ZN(n6792)
         );
  AOI211_X1 U8347 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n9715), .A(n6793), .B(
        n6792), .ZN(n6795) );
  INV_X1 U8348 ( .A(n9717), .ZN(n9560) );
  NAND2_X1 U8349 ( .A1(n9560), .A2(n7453), .ZN(n6794) );
  OAI211_X1 U8350 ( .C1(n6796), .C2(n9716), .A(n6795), .B(n6794), .ZN(P2_U3256) );
  NAND2_X1 U8351 ( .A1(n7539), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6798) );
  NAND2_X1 U8352 ( .A1(n6798), .A2(n6797), .ZN(n6801) );
  INV_X1 U8353 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6799) );
  INV_X1 U8354 ( .A(n7578), .ZN(n6802) );
  AOI22_X1 U8355 ( .A1(n7578), .A2(n6799), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n6802), .ZN(n6800) );
  NOR2_X1 U8356 ( .A1(n6801), .A2(n6800), .ZN(n6982) );
  AOI21_X1 U8357 ( .B1(n6801), .B2(n6800), .A(n6982), .ZN(n6812) );
  INV_X1 U8358 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6803) );
  AOI22_X1 U8359 ( .A1(n7578), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n6803), .B2(
        n6802), .ZN(n6806) );
  OAI21_X1 U8360 ( .B1(n6806), .B2(n6805), .A(n6978), .ZN(n6807) );
  NAND2_X1 U8361 ( .A1(n6807), .A2(n9713), .ZN(n6811) );
  OAI22_X1 U8362 ( .A1(n6808), .A2(n6185), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7582), .ZN(n6809) );
  AOI21_X1 U8363 ( .B1(n9560), .B2(n7578), .A(n6809), .ZN(n6810) );
  OAI211_X1 U8364 ( .C1(n6812), .C2(n9716), .A(n6811), .B(n6810), .ZN(P2_U3258) );
  INV_X1 U8365 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6852) );
  NAND2_X1 U8366 ( .A1(n6839), .A2(n8147), .ZN(n6813) );
  INV_X1 U8367 ( .A(n8316), .ZN(n7009) );
  OR2_X1 U8368 ( .A1(n6815), .A2(n6816), .ZN(n6820) );
  OR2_X1 U8369 ( .A1(n6817), .A2(n6818), .ZN(n6819) );
  OAI211_X1 U8370 ( .C1(n6768), .C2(n6821), .A(n6820), .B(n6819), .ZN(n9834)
         );
  NAND2_X1 U8371 ( .A1(n7009), .A2(n9834), .ZN(n8154) );
  NAND2_X1 U8372 ( .A1(n7260), .A2(n8121), .ZN(n7259) );
  NAND2_X1 U8373 ( .A1(n7009), .A2(n7021), .ZN(n6822) );
  NAND2_X1 U8374 ( .A1(n7259), .A2(n6822), .ZN(n6835) );
  NAND2_X1 U8375 ( .A1(n8105), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6830) );
  INV_X1 U8376 ( .A(n6825), .ZN(n6823) );
  NAND2_X1 U8377 ( .A1(n6823), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6843) );
  NAND2_X1 U8378 ( .A1(n6825), .A2(n6824), .ZN(n6826) );
  AND2_X1 U8379 ( .A1(n6843), .A2(n6826), .ZN(n8018) );
  NAND2_X1 U8380 ( .A1(n7141), .A2(n8018), .ZN(n6829) );
  NAND2_X1 U8381 ( .A1(n6750), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6828) );
  NAND2_X1 U8382 ( .A1(n6463), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6827) );
  NAND4_X1 U8383 ( .A1(n6830), .A2(n6829), .A3(n6828), .A4(n6827), .ZN(n8315)
         );
  INV_X1 U8384 ( .A(n8315), .ZN(n7182) );
  OR2_X1 U8385 ( .A1(n8111), .A2(n6832), .ZN(n6833) );
  NAND2_X1 U8386 ( .A1(n8155), .A2(n8150), .ZN(n8125) );
  NAND2_X1 U8387 ( .A1(n6835), .A2(n8125), .ZN(n7184) );
  OAI21_X1 U8388 ( .B1(n6835), .B2(n8125), .A(n7184), .ZN(n6836) );
  INV_X1 U8389 ( .A(n6836), .ZN(n7180) );
  INV_X1 U8390 ( .A(n6837), .ZN(n8165) );
  NAND2_X1 U8391 ( .A1(n6839), .A2(n7204), .ZN(n8153) );
  NAND2_X1 U8392 ( .A1(n7255), .A2(n8149), .ZN(n6840) );
  XNOR2_X1 U8393 ( .A(n6840), .B(n8125), .ZN(n6849) );
  NAND2_X1 U8394 ( .A1(n8105), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6848) );
  INV_X1 U8395 ( .A(n6843), .ZN(n6841) );
  NAND2_X1 U8396 ( .A1(n6841), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6935) );
  INV_X1 U8397 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6842) );
  NAND2_X1 U8398 ( .A1(n6843), .A2(n6842), .ZN(n6844) );
  AND2_X1 U8399 ( .A1(n6935), .A2(n6844), .ZN(n7186) );
  NAND2_X1 U8400 ( .A1(n7141), .A2(n7186), .ZN(n6847) );
  NAND2_X1 U8401 ( .A1(n6750), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6846) );
  NAND2_X1 U8402 ( .A1(n8106), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6845) );
  NAND4_X1 U8403 ( .A1(n6848), .A2(n6847), .A3(n6846), .A4(n6845), .ZN(n8314)
         );
  INV_X1 U8404 ( .A(n8314), .ZN(n8179) );
  OAI22_X1 U8405 ( .A1(n7009), .A2(n8692), .B1(n8179), .B2(n8694), .ZN(n8019)
         );
  AOI21_X1 U8406 ( .B1(n6849), .B2(n9769), .A(n8019), .ZN(n7177) );
  NAND2_X1 U8407 ( .A1(n7261), .A2(n7021), .ZN(n7262) );
  AOI211_X1 U8408 ( .C1(n8017), .C2(n7262), .A(n9889), .B(n4560), .ZN(n7176)
         );
  AOI21_X1 U8409 ( .B1(n9835), .B2(n8017), .A(n7176), .ZN(n6850) );
  OAI211_X1 U8410 ( .C1(n7180), .C2(n8796), .A(n7177), .B(n6850), .ZN(n6853)
         );
  NAND2_X1 U8411 ( .A1(n6853), .A2(n9872), .ZN(n6851) );
  OAI21_X1 U8412 ( .B1(n9872), .B2(n6852), .A(n6851), .ZN(P2_U3466) );
  INV_X1 U8413 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6855) );
  NAND2_X1 U8414 ( .A1(n6853), .A2(n4260), .ZN(n6854) );
  OAI21_X1 U8415 ( .B1(n4260), .B2(n6855), .A(n6854), .ZN(P2_U3525) );
  INV_X2 U8416 ( .A(n9245), .ZN(n9645) );
  XNOR2_X1 U8417 ( .A(n9664), .B(n6883), .ZN(n6856) );
  NAND2_X1 U8418 ( .A1(n9500), .A2(n6856), .ZN(n9662) );
  NOR2_X1 U8419 ( .A1(n9662), .A2(n9207), .ZN(n6867) );
  NAND2_X1 U8420 ( .A1(n9661), .A2(n9376), .ZN(n6866) );
  AOI22_X1 U8421 ( .A1(n9309), .A2(n9003), .B1(n9311), .B2(n5674), .ZN(n6865)
         );
  INV_X1 U8422 ( .A(n6858), .ZN(n6860) );
  NAND2_X1 U8423 ( .A1(n6860), .A2(n6859), .ZN(n6862) );
  NAND2_X1 U8424 ( .A1(n6862), .A2(n6861), .ZN(n6863) );
  NAND2_X1 U8425 ( .A1(n6863), .A2(n9640), .ZN(n6864) );
  NAND3_X1 U8426 ( .A1(n6866), .A2(n6865), .A3(n6864), .ZN(n9666) );
  AOI211_X1 U8427 ( .C1(n9645), .C2(P1_REG3_REG_1__SCAN_IN), .A(n6867), .B(
        n9666), .ZN(n6876) );
  OR2_X1 U8428 ( .A1(n6868), .A2(n9533), .ZN(n6869) );
  NAND2_X1 U8429 ( .A1(n9650), .A2(n6871), .ZN(n9585) );
  INV_X1 U8430 ( .A(n9585), .ZN(n9632) );
  NAND2_X2 U8431 ( .A1(n9650), .A2(n6872), .ZN(n9595) );
  OAI22_X1 U8432 ( .A1(n9595), .A2(n9664), .B1(n6873), .B2(n9650), .ZN(n6874)
         );
  AOI21_X1 U8433 ( .B1(n9632), .B2(n9661), .A(n6874), .ZN(n6875) );
  OAI21_X1 U8434 ( .B1(n6876), .B2(n9647), .A(n6875), .ZN(P1_U3290) );
  INV_X1 U8435 ( .A(n7826), .ZN(n7707) );
  OAI222_X1 U8436 ( .A1(n8830), .A2(n7827), .B1(P2_U3152), .B2(n6877), .C1(
        n7667), .C2(n7707), .ZN(P2_U3337) );
  INV_X1 U8437 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6886) );
  INV_X1 U8438 ( .A(n6878), .ZN(n6879) );
  AOI22_X1 U8439 ( .A1(n6879), .A2(n9650), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9645), .ZN(n6885) );
  NOR2_X1 U8440 ( .A1(n6881), .A2(n6880), .ZN(n6882) );
  NAND2_X1 U8441 ( .A1(n9650), .A2(n6882), .ZN(n9584) );
  OAI21_X1 U8442 ( .B1(n9631), .B2(n9254), .A(n6883), .ZN(n6884) );
  OAI211_X1 U8443 ( .C1(n6886), .C2(n9650), .A(n6885), .B(n6884), .ZN(P1_U3291) );
  OR2_X1 U8444 ( .A1(n6887), .A2(n9694), .ZN(n6888) );
  OAI21_X1 U8445 ( .B1(n9697), .B2(n5996), .A(n6888), .ZN(P1_U3525) );
  INV_X1 U8446 ( .A(n6890), .ZN(n6894) );
  INV_X1 U8447 ( .A(n6891), .ZN(n6893) );
  NOR3_X1 U8448 ( .A1(n6894), .A2(n6893), .A3(n6892), .ZN(n6897) );
  INV_X1 U8449 ( .A(n6895), .ZN(n6896) );
  OAI21_X1 U8450 ( .B1(n6897), .B2(n6896), .A(n8970), .ZN(n6902) );
  INV_X1 U8451 ( .A(n6898), .ZN(n6900) );
  OAI22_X1 U8452 ( .A1(n8977), .A2(n5706), .B1(n8987), .B2(n7043), .ZN(n6899)
         );
  AOI211_X1 U8453 ( .C1(n8984), .C2(n9001), .A(n6900), .B(n6899), .ZN(n6901)
         );
  OAI211_X1 U8454 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8906), .A(n6902), .B(
        n6901), .ZN(P1_U3216) );
  NAND2_X1 U8455 ( .A1(n6904), .A2(n6903), .ZN(n7013) );
  XNOR2_X1 U8456 ( .A(n6919), .B(n7204), .ZN(n6906) );
  NAND2_X1 U8457 ( .A1(n8317), .A2(n6739), .ZN(n6907) );
  NAND2_X1 U8458 ( .A1(n6906), .A2(n6907), .ZN(n6910) );
  INV_X1 U8459 ( .A(n6906), .ZN(n6909) );
  INV_X1 U8460 ( .A(n6907), .ZN(n6908) );
  NAND2_X1 U8461 ( .A1(n6909), .A2(n6908), .ZN(n6911) );
  XNOR2_X1 U8462 ( .A(n9834), .B(n6912), .ZN(n6914) );
  AND2_X1 U8463 ( .A1(n8316), .A2(n6739), .ZN(n6915) );
  XNOR2_X1 U8464 ( .A(n6914), .B(n6915), .ZN(n7020) );
  INV_X1 U8465 ( .A(n6914), .ZN(n6917) );
  INV_X1 U8466 ( .A(n6915), .ZN(n6916) );
  NAND2_X1 U8467 ( .A1(n6917), .A2(n6916), .ZN(n6918) );
  XNOR2_X1 U8468 ( .A(n6919), .B(n8017), .ZN(n6920) );
  NAND2_X1 U8469 ( .A1(n8315), .A2(n6739), .ZN(n6921) );
  NAND2_X1 U8470 ( .A1(n6920), .A2(n6921), .ZN(n6924) );
  INV_X1 U8471 ( .A(n6920), .ZN(n6923) );
  INV_X1 U8472 ( .A(n6921), .ZN(n6922) );
  NAND2_X1 U8473 ( .A1(n6923), .A2(n6922), .ZN(n6925) );
  AND2_X1 U8474 ( .A1(n6924), .A2(n6925), .ZN(n8021) );
  OR2_X1 U8475 ( .A1(n6815), .A2(n6926), .ZN(n6929) );
  OR2_X1 U8476 ( .A1(n8111), .A2(n6927), .ZN(n6928) );
  OAI211_X1 U8477 ( .C1(n6768), .C2(n6930), .A(n6929), .B(n6928), .ZN(n8178)
         );
  XNOR2_X1 U8478 ( .A(n8178), .B(n6912), .ZN(n7125) );
  NAND2_X1 U8479 ( .A1(n8314), .A2(n8118), .ZN(n7126) );
  XNOR2_X1 U8480 ( .A(n7125), .B(n7126), .ZN(n6931) );
  OAI21_X1 U8481 ( .B1(n6932), .B2(n6931), .A(n7129), .ZN(n6946) );
  NAND2_X1 U8482 ( .A1(n8105), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6940) );
  INV_X1 U8483 ( .A(n6935), .ZN(n6933) );
  NAND2_X1 U8484 ( .A1(n6933), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7118) );
  INV_X1 U8485 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6934) );
  NAND2_X1 U8486 ( .A1(n6935), .A2(n6934), .ZN(n6936) );
  AND2_X1 U8487 ( .A1(n7118), .A2(n6936), .ZN(n7712) );
  NAND2_X1 U8488 ( .A1(n7141), .A2(n7712), .ZN(n6939) );
  NAND2_X1 U8489 ( .A1(n6750), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6938) );
  NAND2_X1 U8490 ( .A1(n8106), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6937) );
  NAND4_X1 U8491 ( .A1(n6940), .A2(n6939), .A3(n6938), .A4(n6937), .ZN(n9763)
         );
  INV_X1 U8492 ( .A(n9763), .ZN(n7333) );
  OAI22_X1 U8493 ( .A1(n9703), .A2(n7333), .B1(n9844), .B2(n9701), .ZN(n6945)
         );
  NAND2_X1 U8494 ( .A1(n8073), .A2(n7186), .ZN(n6942) );
  OAI211_X1 U8495 ( .C1(n9704), .C2(n7182), .A(n6943), .B(n6942), .ZN(n6944)
         );
  AOI211_X1 U8496 ( .C1(n9709), .C2(n6946), .A(n6945), .B(n6944), .ZN(n6947)
         );
  INV_X1 U8497 ( .A(n6947), .ZN(P2_U3241) );
  NAND2_X1 U8498 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8836) );
  XNOR2_X1 U8499 ( .A(n7269), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n6950) );
  OAI21_X1 U8500 ( .B1(n6954), .B2(P1_REG1_REG_13__SCAN_IN), .A(n6948), .ZN(
        n6949) );
  NAND2_X1 U8501 ( .A1(n6950), .A2(n6949), .ZN(n7277) );
  OAI21_X1 U8502 ( .B1(n6950), .B2(n6949), .A(n7277), .ZN(n6951) );
  NAND2_X1 U8503 ( .A1(n9623), .A2(n6951), .ZN(n6952) );
  OAI211_X1 U8504 ( .C1(n9029), .C2(n7269), .A(n8836), .B(n6952), .ZN(n6958)
         );
  INV_X1 U8505 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6955) );
  AOI211_X1 U8506 ( .C1(n6956), .C2(n6955), .A(n7271), .B(n9017), .ZN(n6957)
         );
  AOI211_X1 U8507 ( .C1(P1_ADDR_REG_14__SCAN_IN), .C2(n9611), .A(n6958), .B(
        n6957), .ZN(n6959) );
  INV_X1 U8508 ( .A(n6959), .ZN(P1_U3255) );
  NAND2_X1 U8509 ( .A1(n7043), .A2(n6960), .ZN(n6961) );
  NAND2_X1 U8510 ( .A1(n6962), .A2(n6961), .ZN(n7042) );
  NAND2_X1 U8511 ( .A1(n7042), .A2(n7041), .ZN(n7040) );
  NAND2_X1 U8512 ( .A1(n7032), .A2(n5706), .ZN(n6963) );
  NAND2_X1 U8513 ( .A1(n7040), .A2(n6963), .ZN(n6965) );
  NAND2_X1 U8514 ( .A1(n6965), .A2(n6964), .ZN(n6999) );
  OAI21_X1 U8515 ( .B1(n6965), .B2(n6964), .A(n6999), .ZN(n7058) );
  OAI22_X1 U8516 ( .A1(n9638), .A2(n7032), .B1(n7379), .B2(n9635), .ZN(n6970)
         );
  XNOR2_X1 U8517 ( .A(n6967), .B(n6966), .ZN(n6968) );
  NOR2_X1 U8518 ( .A1(n6968), .A2(n9370), .ZN(n6969) );
  AOI211_X1 U8519 ( .C1(n9376), .C2(n7058), .A(n6970), .B(n6969), .ZN(n7062)
         );
  INV_X1 U8520 ( .A(n6971), .ZN(n7048) );
  NAND2_X1 U8521 ( .A1(n6971), .A2(n7033), .ZN(n6993) );
  INV_X1 U8522 ( .A(n6993), .ZN(n6972) );
  AOI21_X1 U8523 ( .B1(n7059), .B2(n7048), .A(n6972), .ZN(n7060) );
  NAND2_X1 U8524 ( .A1(n7060), .A2(n9631), .ZN(n6974) );
  AOI22_X1 U8525 ( .A1(n9647), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7027), .B2(
        n9645), .ZN(n6973) );
  OAI211_X1 U8526 ( .C1(n7033), .C2(n9595), .A(n6974), .B(n6973), .ZN(n6975)
         );
  AOI21_X1 U8527 ( .B1(n7058), .B2(n9632), .A(n6975), .ZN(n6976) );
  OAI21_X1 U8528 ( .B1(n7062), .B2(n9647), .A(n6976), .ZN(P1_U3287) );
  INV_X1 U8529 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6977) );
  AOI22_X1 U8530 ( .A1(n7726), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n6977), .B2(
        n7422), .ZN(n6980) );
  OAI21_X1 U8531 ( .B1(n7578), .B2(P2_REG1_REG_13__SCAN_IN), .A(n6978), .ZN(
        n6979) );
  NAND2_X1 U8532 ( .A1(n6980), .A2(n6979), .ZN(n7417) );
  OAI21_X1 U8533 ( .B1(n6980), .B2(n6979), .A(n7417), .ZN(n6989) );
  AND2_X1 U8534 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7942) );
  AOI21_X1 U8535 ( .B1(n9715), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n7942), .ZN(
        n6981) );
  OAI21_X1 U8536 ( .B1(n9717), .B2(n7422), .A(n6981), .ZN(n6988) );
  NOR2_X1 U8537 ( .A1(n7578), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6983) );
  NOR2_X1 U8538 ( .A1(n6983), .A2(n6982), .ZN(n6985) );
  INV_X1 U8539 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7421) );
  AOI22_X1 U8540 ( .A1(n7726), .A2(n7421), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7422), .ZN(n6984) );
  NOR2_X1 U8541 ( .A1(n6985), .A2(n6984), .ZN(n7420) );
  AOI21_X1 U8542 ( .B1(n6985), .B2(n6984), .A(n7420), .ZN(n6986) );
  NOR2_X1 U8543 ( .A1(n6986), .A2(n9716), .ZN(n6987) );
  AOI211_X1 U8544 ( .C1(n6989), .C2(n9713), .A(n6988), .B(n6987), .ZN(n6990)
         );
  INV_X1 U8545 ( .A(n6990), .ZN(P2_U3259) );
  OAI222_X1 U8546 ( .A1(n8830), .A2(n7809), .B1(P2_U3152), .B2(n6449), .C1(
        n7667), .C2(n6991), .ZN(P2_U3338) );
  OR2_X1 U8547 ( .A1(n6993), .A2(n7089), .ZN(n7365) );
  INV_X1 U8548 ( .A(n7365), .ZN(n6992) );
  AOI211_X1 U8549 ( .C1(n7089), .C2(n6993), .A(n9682), .B(n6992), .ZN(n7070)
         );
  INV_X1 U8550 ( .A(n7250), .ZN(n6994) );
  NOR2_X1 U8551 ( .A1(n9245), .A2(n6994), .ZN(n6997) );
  XOR2_X1 U8552 ( .A(n6995), .B(n7000), .Z(n6996) );
  OAI222_X1 U8553 ( .A1(n9638), .A2(n7246), .B1(n9635), .B2(n7438), .C1(n6996), 
        .C2(n9370), .ZN(n7069) );
  AOI211_X1 U8554 ( .C1(n7070), .C2(n9250), .A(n6997), .B(n7069), .ZN(n7008)
         );
  NAND2_X1 U8555 ( .A1(n7246), .A2(n7033), .ZN(n6998) );
  INV_X1 U8556 ( .A(n7000), .ZN(n7001) );
  OAI21_X1 U8557 ( .B1(n7002), .B2(n7001), .A(n7091), .ZN(n7072) );
  INV_X1 U8558 ( .A(n7072), .ZN(n7006) );
  INV_X1 U8559 ( .A(n9364), .ZN(n9323) );
  OAI22_X1 U8560 ( .A1(n9595), .A2(n7247), .B1(n4386), .B2(n9650), .ZN(n7005)
         );
  AOI21_X1 U8561 ( .B1(n7006), .B2(n9323), .A(n7005), .ZN(n7007) );
  OAI21_X1 U8562 ( .B1(n7008), .B2(n9647), .A(n7007), .ZN(P1_U3286) );
  OAI22_X1 U8563 ( .A1(n9703), .A2(n7009), .B1(n8147), .B2(n9701), .ZN(n7011)
         );
  OAI22_X1 U8564 ( .A1(n8080), .A2(P2_REG3_REG_3__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n6749), .ZN(n7010) );
  AOI211_X1 U8565 ( .C1(n7985), .C2(n8318), .A(n7011), .B(n7010), .ZN(n7016)
         );
  OAI211_X1 U8566 ( .C1(n7014), .C2(n7013), .A(n9709), .B(n7012), .ZN(n7015)
         );
  NAND2_X1 U8567 ( .A1(n7016), .A2(n7015), .ZN(P2_U3220) );
  INV_X1 U8568 ( .A(n7017), .ZN(n7018) );
  AOI21_X1 U8569 ( .B1(n7020), .B2(n7019), .A(n7018), .ZN(n7026) );
  OAI22_X1 U8570 ( .A1(n9703), .A2(n7182), .B1(n7021), .B2(n9701), .ZN(n7024)
         );
  INV_X1 U8571 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7022) );
  OAI22_X1 U8572 ( .A1(n8080), .A2(n7265), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7022), .ZN(n7023) );
  AOI211_X1 U8573 ( .C1(n7985), .C2(n8317), .A(n7024), .B(n7023), .ZN(n7025)
         );
  OAI21_X1 U8574 ( .B1(n7026), .B2(n8085), .A(n7025), .ZN(P2_U3232) );
  INV_X1 U8575 ( .A(n7027), .ZN(n7038) );
  OAI21_X1 U8576 ( .B1(n7030), .B2(n7029), .A(n7028), .ZN(n7031) );
  NAND2_X1 U8577 ( .A1(n7031), .A2(n8970), .ZN(n7037) );
  OAI22_X1 U8578 ( .A1(n8977), .A2(n7033), .B1(n8987), .B2(n7032), .ZN(n7034)
         );
  AOI211_X1 U8579 ( .C1(n8984), .C2(n9000), .A(n7035), .B(n7034), .ZN(n7036)
         );
  OAI211_X1 U8580 ( .C1(n8906), .C2(n7038), .A(n7037), .B(n7036), .ZN(P1_U3228) );
  XNOR2_X1 U8581 ( .A(n7039), .B(n7041), .ZN(n7046) );
  OAI21_X1 U8582 ( .B1(n7042), .B2(n7041), .A(n7040), .ZN(n9671) );
  OAI22_X1 U8583 ( .A1(n9638), .A2(n7043), .B1(n7246), .B2(n9635), .ZN(n7044)
         );
  AOI21_X1 U8584 ( .B1(n9671), .B2(n9376), .A(n7044), .ZN(n7045) );
  OAI21_X1 U8585 ( .B1(n9370), .B2(n7046), .A(n7045), .ZN(n9669) );
  INV_X1 U8586 ( .A(n9669), .ZN(n7056) );
  INV_X1 U8587 ( .A(n7047), .ZN(n7049) );
  OAI21_X1 U8588 ( .B1(n5706), .B2(n7049), .A(n7048), .ZN(n9668) );
  AOI22_X1 U8589 ( .A1(n9647), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9645), .B2(
        n7050), .ZN(n7053) );
  NAND2_X1 U8590 ( .A1(n9254), .A2(n7051), .ZN(n7052) );
  OAI211_X1 U8591 ( .C1(n9668), .C2(n9584), .A(n7053), .B(n7052), .ZN(n7054)
         );
  AOI21_X1 U8592 ( .B1(n9671), .B2(n9632), .A(n7054), .ZN(n7055) );
  OAI21_X1 U8593 ( .B1(n7056), .B2(n9647), .A(n7055), .ZN(P1_U3288) );
  INV_X1 U8594 ( .A(n7839), .ZN(n7668) );
  OAI222_X1 U8595 ( .A1(P1_U3084), .A2(n5678), .B1(n9552), .B2(n7668), .C1(
        n7057), .C2(n7705), .ZN(P1_U3331) );
  INV_X1 U8596 ( .A(n7058), .ZN(n7063) );
  AOI22_X1 U8597 ( .A1(n7060), .A2(n9500), .B1(n9568), .B2(n7059), .ZN(n7061)
         );
  OAI211_X1 U8598 ( .C1(n7063), .C2(n9510), .A(n7062), .B(n7061), .ZN(n7066)
         );
  NAND2_X1 U8599 ( .A1(n7066), .A2(n9697), .ZN(n7064) );
  OAI21_X1 U8600 ( .B1(n9697), .B2(n7065), .A(n7064), .ZN(P1_U3527) );
  INV_X1 U8601 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7068) );
  NAND2_X1 U8602 ( .A1(n7066), .A2(n9530), .ZN(n7067) );
  OAI21_X1 U8603 ( .B1(n9530), .B2(n7068), .A(n7067), .ZN(P1_U3466) );
  AOI211_X1 U8604 ( .C1(n9568), .C2(n7089), .A(n7070), .B(n7069), .ZN(n7071)
         );
  OAI21_X1 U8605 ( .B1(n9497), .B2(n7072), .A(n7071), .ZN(n7075) );
  NAND2_X1 U8606 ( .A1(n7075), .A2(n9697), .ZN(n7073) );
  OAI21_X1 U8607 ( .B1(n9697), .B2(n7074), .A(n7073), .ZN(P1_U3528) );
  INV_X1 U8608 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7077) );
  NAND2_X1 U8609 ( .A1(n7075), .A2(n9530), .ZN(n7076) );
  OAI21_X1 U8610 ( .B1(n9530), .B2(n7077), .A(n7076), .ZN(P1_U3469) );
  AOI22_X1 U8611 ( .A1(n9254), .A2(n8948), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9645), .ZN(n7078) );
  OAI21_X1 U8612 ( .B1(n9584), .B2(n7079), .A(n7078), .ZN(n7082) );
  MUX2_X1 U8613 ( .A(n7080), .B(P1_REG2_REG_2__SCAN_IN), .S(n9647), .Z(n7081)
         );
  AOI211_X1 U8614 ( .C1(n9632), .C2(n7083), .A(n7082), .B(n7081), .ZN(n7084)
         );
  INV_X1 U8615 ( .A(n7084), .ZN(P1_U3289) );
  NAND2_X1 U8616 ( .A1(n7086), .A2(n7085), .ZN(n7087) );
  XNOR2_X1 U8617 ( .A(n8998), .B(n9675), .ZN(n7094) );
  XNOR2_X1 U8618 ( .A(n7087), .B(n7094), .ZN(n7088) );
  AOI222_X1 U8619 ( .A1(n9640), .A2(n7088), .B1(n8997), .B2(n9309), .C1(n8999), 
        .C2(n9311), .ZN(n9674) );
  NAND2_X1 U8620 ( .A1(n9000), .A2(n7089), .ZN(n7090) );
  NAND2_X1 U8621 ( .A1(n7438), .A2(n7380), .ZN(n7093) );
  OAI21_X1 U8622 ( .B1(n7095), .B2(n7094), .A(n7476), .ZN(n9677) );
  OR2_X1 U8623 ( .A1(n7365), .A2(n7523), .ZN(n7363) );
  INV_X1 U8624 ( .A(n7484), .ZN(n7485) );
  AOI21_X1 U8625 ( .B1(n7363), .B2(n7098), .A(n9682), .ZN(n7096) );
  NAND2_X1 U8626 ( .A1(n7485), .A2(n7096), .ZN(n9673) );
  NOR2_X1 U8627 ( .A1(n7097), .A2(n9207), .ZN(n9406) );
  INV_X1 U8628 ( .A(n9406), .ZN(n7101) );
  AOI22_X1 U8629 ( .A1(n9647), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7442), .B2(
        n9645), .ZN(n7100) );
  NAND2_X1 U8630 ( .A1(n9254), .A2(n7098), .ZN(n7099) );
  OAI211_X1 U8631 ( .C1(n9673), .C2(n7101), .A(n7100), .B(n7099), .ZN(n7102)
         );
  AOI21_X1 U8632 ( .B1(n9677), .B2(n9323), .A(n7102), .ZN(n7103) );
  OAI21_X1 U8633 ( .B1(n9674), .B2(n9647), .A(n7103), .ZN(P1_U3284) );
  NAND2_X1 U8634 ( .A1(n8106), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7110) );
  NAND2_X1 U8635 ( .A1(n6750), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7109) );
  INV_X1 U8636 ( .A(n7120), .ZN(n7104) );
  NAND2_X1 U8637 ( .A1(n7104), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7319) );
  INV_X1 U8638 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7105) );
  NAND2_X1 U8639 ( .A1(n7120), .A2(n7105), .ZN(n7106) );
  AND2_X1 U8640 ( .A1(n7319), .A2(n7106), .ZN(n7303) );
  NAND2_X1 U8641 ( .A1(n7141), .A2(n7303), .ZN(n7108) );
  NAND2_X1 U8642 ( .A1(n8105), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7107) );
  NAND4_X1 U8643 ( .A1(n7110), .A2(n7109), .A3(n7108), .A4(n7107), .ZN(n9765)
         );
  INV_X1 U8644 ( .A(n9765), .ZN(n7336) );
  AND2_X1 U8645 ( .A1(n7111), .A2(n8110), .ZN(n7116) );
  NOR2_X1 U8646 ( .A1(n6768), .A2(n7112), .ZN(n7115) );
  NOR2_X1 U8647 ( .A1(n8111), .A2(n7113), .ZN(n7114) );
  OAI22_X1 U8648 ( .A1(n9703), .A2(n7336), .B1(n9858), .B2(n9701), .ZN(n7124)
         );
  NAND2_X1 U8649 ( .A1(n7118), .A2(n7117), .ZN(n7119) );
  AND2_X1 U8650 ( .A1(n7120), .A2(n7119), .ZN(n9774) );
  INV_X1 U8651 ( .A(n9774), .ZN(n7122) );
  OAI21_X1 U8652 ( .B1(n8080), .B2(n7122), .A(n7121), .ZN(n7123) );
  AOI211_X1 U8653 ( .C1(n7985), .C2(n9763), .A(n7124), .B(n7123), .ZN(n7149)
         );
  INV_X1 U8654 ( .A(n7125), .ZN(n7127) );
  NAND2_X1 U8655 ( .A1(n7127), .A2(n7126), .ZN(n7128) );
  OR2_X1 U8656 ( .A1(n7130), .A2(n6815), .ZN(n7133) );
  OR2_X1 U8657 ( .A1(n8111), .A2(n7131), .ZN(n7132) );
  OAI211_X1 U8658 ( .C1(n6768), .C2(n7134), .A(n7133), .B(n7132), .ZN(n7711)
         );
  XNOR2_X1 U8659 ( .A(n6919), .B(n7711), .ZN(n7135) );
  NAND2_X1 U8660 ( .A1(n9763), .A2(n8118), .ZN(n7136) );
  NAND2_X1 U8661 ( .A1(n7135), .A2(n7136), .ZN(n7139) );
  INV_X1 U8662 ( .A(n7135), .ZN(n7138) );
  INV_X1 U8663 ( .A(n7136), .ZN(n7137) );
  NAND2_X1 U8664 ( .A1(n7138), .A2(n7137), .ZN(n7140) );
  AND2_X1 U8665 ( .A1(n7139), .A2(n7140), .ZN(n7709) );
  XNOR2_X1 U8666 ( .A(n8185), .B(n6912), .ZN(n7295) );
  NAND2_X1 U8667 ( .A1(n8105), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7145) );
  NAND2_X1 U8668 ( .A1(n7901), .A2(n9774), .ZN(n7144) );
  NAND2_X1 U8669 ( .A1(n6750), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7143) );
  NAND2_X1 U8670 ( .A1(n8106), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7142) );
  NAND4_X1 U8671 ( .A1(n7145), .A2(n7144), .A3(n7143), .A4(n7142), .ZN(n8313)
         );
  NAND2_X1 U8672 ( .A1(n8313), .A2(n8118), .ZN(n7293) );
  XNOR2_X1 U8673 ( .A(n7295), .B(n7293), .ZN(n7146) );
  OAI211_X1 U8674 ( .C1(n7147), .C2(n7146), .A(n7297), .B(n9709), .ZN(n7148)
         );
  NAND2_X1 U8675 ( .A1(n7149), .A2(n7148), .ZN(P2_U3223) );
  INV_X1 U8676 ( .A(n7852), .ZN(n7152) );
  NAND2_X1 U8677 ( .A1(n9549), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7150) );
  OAI211_X1 U8678 ( .C1(n7152), .C2(n9552), .A(n7151), .B(n7150), .ZN(P1_U3330) );
  NAND3_X1 U8679 ( .A1(n7155), .A2(n7154), .A3(n7153), .ZN(n7156) );
  NOR2_X1 U8680 ( .A1(n7157), .A2(n7156), .ZN(n7160) );
  INV_X1 U8681 ( .A(n7158), .ZN(n7159) );
  NAND2_X1 U8682 ( .A1(n7160), .A2(n7159), .ZN(n7165) );
  OR2_X1 U8683 ( .A1(n7161), .A2(n8389), .ZN(n7196) );
  NAND2_X1 U8684 ( .A1(n9757), .A2(n7196), .ZN(n7162) );
  INV_X1 U8685 ( .A(n8703), .ZN(n8522) );
  OAI22_X1 U8686 ( .A1(n8613), .A2(n9711), .B1(n7163), .B2(n9779), .ZN(n7170)
         );
  AOI22_X1 U8687 ( .A1(n9733), .A2(n7167), .B1(n9779), .B2(n7166), .ZN(n7168)
         );
  OAI21_X1 U8688 ( .B1(n6760), .B2(n9777), .A(n7168), .ZN(n7169) );
  AOI211_X1 U8689 ( .C1(n8522), .C2(n7171), .A(n7170), .B(n7169), .ZN(n7172)
         );
  INV_X1 U8690 ( .A(n7172), .ZN(P2_U3295) );
  NAND2_X1 U8691 ( .A1(n7852), .A2(n8825), .ZN(n7173) );
  OAI211_X1 U8692 ( .C1(n7853), .C2(n8830), .A(n7173), .B(n8309), .ZN(P2_U3335) );
  NOR2_X1 U8693 ( .A1(n9775), .A2(n6456), .ZN(n8585) );
  INV_X1 U8694 ( .A(n8018), .ZN(n7174) );
  OAI22_X1 U8695 ( .A1(n9777), .A2(n7181), .B1(n8613), .B2(n7174), .ZN(n7175)
         );
  AOI21_X1 U8696 ( .B1(n8585), .B2(n7176), .A(n7175), .ZN(n7179) );
  MUX2_X1 U8697 ( .A(n7177), .B(n6493), .S(n9775), .Z(n7178) );
  OAI211_X1 U8698 ( .C1(n7180), .C2(n8703), .A(n7179), .B(n7178), .ZN(P2_U3291) );
  NAND2_X1 U8699 ( .A1(n7182), .A2(n7181), .ZN(n7183) );
  XNOR2_X1 U8700 ( .A(n8314), .B(n8178), .ZN(n8130) );
  XOR2_X1 U8701 ( .A(n7212), .B(n8130), .Z(n9848) );
  INV_X1 U8702 ( .A(n7214), .ZN(n7216) );
  AOI21_X1 U8703 ( .B1(n8178), .B2(n7185), .A(n7216), .ZN(n9843) );
  AOI22_X1 U8704 ( .A1(n9733), .A2(n9843), .B1(n7186), .B2(n9773), .ZN(n7187)
         );
  OAI21_X1 U8705 ( .B1(n9844), .B2(n9777), .A(n7187), .ZN(n7193) );
  AND2_X1 U8706 ( .A1(n8149), .A2(n8150), .ZN(n8145) );
  NAND2_X1 U8707 ( .A1(n7188), .A2(n8155), .ZN(n7218) );
  XNOR2_X1 U8708 ( .A(n7218), .B(n8130), .ZN(n7189) );
  NAND2_X1 U8709 ( .A1(n7189), .A2(n9769), .ZN(n7191) );
  AOI22_X1 U8710 ( .A1(n9762), .A2(n8315), .B1(n9763), .B2(n9764), .ZN(n7190)
         );
  NAND2_X1 U8711 ( .A1(n7191), .A2(n7190), .ZN(n9847) );
  MUX2_X1 U8712 ( .A(n9847), .B(P2_REG2_REG_6__SCAN_IN), .S(n9775), .Z(n7192)
         );
  AOI211_X1 U8713 ( .C1(n8522), .C2(n9848), .A(n7193), .B(n7192), .ZN(n7194)
         );
  INV_X1 U8714 ( .A(n7194), .ZN(P2_U3290) );
  OAI22_X1 U8715 ( .A1(n9754), .A2(n7195), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8613), .ZN(n7203) );
  INV_X1 U8716 ( .A(n7196), .ZN(n7197) );
  NAND2_X1 U8717 ( .A1(n9779), .A2(n7197), .ZN(n9755) );
  INV_X1 U8718 ( .A(n9755), .ZN(n9734) );
  NAND2_X1 U8719 ( .A1(n9734), .A2(n7198), .ZN(n7201) );
  NAND2_X1 U8720 ( .A1(n7199), .A2(n9779), .ZN(n7200) );
  OAI211_X1 U8721 ( .C1(n6496), .C2(n9779), .A(n7201), .B(n7200), .ZN(n7202)
         );
  AOI211_X1 U8722 ( .C1(n8698), .C2(n7204), .A(n7203), .B(n7202), .ZN(n7205)
         );
  INV_X1 U8723 ( .A(n7205), .ZN(P2_U3293) );
  XNOR2_X1 U8724 ( .A(n6453), .B(n9821), .ZN(n8126) );
  INV_X1 U8725 ( .A(n8126), .ZN(n9823) );
  AOI22_X1 U8726 ( .A1(n9823), .A2(n9769), .B1(n9764), .B2(n8320), .ZN(n9825)
         );
  OAI21_X1 U8727 ( .B1(n7206), .B2(n8613), .A(n9825), .ZN(n7209) );
  NOR2_X1 U8728 ( .A1(n9779), .A2(n7207), .ZN(n7208) );
  AOI21_X1 U8729 ( .B1(n9779), .B2(n7209), .A(n7208), .ZN(n7211) );
  OAI21_X1 U8730 ( .B1(n8698), .B2(n9733), .A(n9821), .ZN(n7210) );
  OAI211_X1 U8731 ( .C1(n8126), .C2(n8703), .A(n7211), .B(n7210), .ZN(P2_U3296) );
  NAND2_X1 U8732 ( .A1(n7212), .A2(n9844), .ZN(n7213) );
  NAND2_X1 U8733 ( .A1(n7333), .A2(n7711), .ZN(n8194) );
  NAND2_X1 U8734 ( .A1(n9850), .A2(n9763), .ZN(n8182) );
  NAND2_X1 U8735 ( .A1(n8194), .A2(n8182), .ZN(n7331) );
  XNOR2_X1 U8736 ( .A(n7332), .B(n7331), .ZN(n9854) );
  INV_X1 U8737 ( .A(n9854), .ZN(n7225) );
  INV_X1 U8738 ( .A(n9751), .ZN(n7215) );
  OAI21_X1 U8739 ( .B1(n9850), .B2(n7216), .A(n7215), .ZN(n9851) );
  INV_X1 U8740 ( .A(n7712), .ZN(n7217) );
  OAI22_X1 U8741 ( .A1(n9851), .A2(n9754), .B1(n7217), .B2(n8613), .ZN(n7223)
         );
  NOR2_X1 U8742 ( .A1(n9844), .A2(n8314), .ZN(n8156) );
  INV_X1 U8743 ( .A(n7331), .ZN(n8181) );
  OAI211_X1 U8744 ( .C1(n7219), .C2(n8181), .A(n7340), .B(n9769), .ZN(n7221)
         );
  AOI22_X1 U8745 ( .A1(n9764), .A2(n8313), .B1(n8314), .B2(n9762), .ZN(n7220)
         );
  NAND2_X1 U8746 ( .A1(n7221), .A2(n7220), .ZN(n9852) );
  MUX2_X1 U8747 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9852), .S(n9779), .Z(n7222)
         );
  AOI211_X1 U8748 ( .C1(n8698), .C2(n7711), .A(n7223), .B(n7222), .ZN(n7224)
         );
  OAI21_X1 U8749 ( .B1(n7225), .B2(n8703), .A(n7224), .ZN(P2_U3289) );
  NAND2_X1 U8750 ( .A1(n7226), .A2(n8120), .ZN(n7227) );
  NAND2_X1 U8751 ( .A1(n7228), .A2(n7227), .ZN(n7229) );
  NAND2_X1 U8752 ( .A1(n7229), .A2(n9769), .ZN(n7231) );
  AOI22_X1 U8753 ( .A1(n9762), .A2(n8320), .B1(n8317), .B2(n9764), .ZN(n7230)
         );
  AND2_X1 U8754 ( .A1(n7231), .A2(n7230), .ZN(n9830) );
  OAI21_X1 U8755 ( .B1(n7233), .B2(n8120), .A(n7232), .ZN(n9832) );
  AOI22_X1 U8756 ( .A1(n8522), .A2(n9832), .B1(n8698), .B2(n9827), .ZN(n7241)
         );
  INV_X1 U8757 ( .A(n7234), .ZN(n7235) );
  AOI21_X1 U8758 ( .B1(n9827), .B2(n7236), .A(n7235), .ZN(n9828) );
  OAI22_X1 U8759 ( .A1(n8613), .A2(n7238), .B1(n7237), .B2(n9779), .ZN(n7239)
         );
  AOI21_X1 U8760 ( .B1(n9733), .B2(n9828), .A(n7239), .ZN(n7240) );
  OAI211_X1 U8761 ( .C1(n9775), .C2(n9830), .A(n7241), .B(n7240), .ZN(P2_U3294) );
  NAND2_X1 U8762 ( .A1(n7243), .A2(n7242), .ZN(n7371) );
  OAI21_X1 U8763 ( .B1(n7243), .B2(n7242), .A(n7371), .ZN(n7244) );
  NOR2_X1 U8764 ( .A1(n7244), .A2(n7245), .ZN(n7374) );
  AOI21_X1 U8765 ( .B1(n7245), .B2(n7244), .A(n7374), .ZN(n7253) );
  NAND2_X1 U8766 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9626) );
  INV_X1 U8767 ( .A(n9626), .ZN(n7249) );
  OAI22_X1 U8768 ( .A1(n8977), .A2(n7247), .B1(n8987), .B2(n7246), .ZN(n7248)
         );
  AOI211_X1 U8769 ( .C1(n8984), .C2(n8999), .A(n7249), .B(n7248), .ZN(n7252)
         );
  NAND2_X1 U8770 ( .A1(n8982), .A2(n7250), .ZN(n7251) );
  OAI211_X1 U8771 ( .C1(n7253), .C2(n8991), .A(n7252), .B(n7251), .ZN(P1_U3225) );
  AOI21_X1 U8772 ( .B1(n7254), .B2(n8121), .A(n8690), .ZN(n7256) );
  NAND2_X1 U8773 ( .A1(n7256), .A2(n7255), .ZN(n7258) );
  AOI22_X1 U8774 ( .A1(n9762), .A2(n8317), .B1(n8315), .B2(n9764), .ZN(n7257)
         );
  AND2_X1 U8775 ( .A1(n7258), .A2(n7257), .ZN(n9839) );
  OAI21_X1 U8776 ( .B1(n7260), .B2(n8121), .A(n7259), .ZN(n9841) );
  AOI22_X1 U8777 ( .A1(n8522), .A2(n9841), .B1(n8698), .B2(n9834), .ZN(n7268)
         );
  INV_X1 U8778 ( .A(n7261), .ZN(n7264) );
  INV_X1 U8779 ( .A(n7262), .ZN(n7263) );
  AOI21_X1 U8780 ( .B1(n9834), .B2(n7264), .A(n7263), .ZN(n9837) );
  OAI22_X1 U8781 ( .A1(n8613), .A2(n7265), .B1(n6495), .B2(n9779), .ZN(n7266)
         );
  AOI21_X1 U8782 ( .B1(n9733), .B2(n9837), .A(n7266), .ZN(n7267) );
  OAI211_X1 U8783 ( .C1(n9775), .C2(n9839), .A(n7268), .B(n7267), .ZN(P2_U3292) );
  NOR2_X1 U8784 ( .A1(n7270), .A2(n7269), .ZN(n7272) );
  XNOR2_X1 U8785 ( .A(n7490), .B(n7497), .ZN(n7274) );
  INV_X1 U8786 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7273) );
  NOR2_X1 U8787 ( .A1(n7273), .A2(n7274), .ZN(n7491) );
  AOI211_X1 U8788 ( .C1(n7274), .C2(n7273), .A(n7491), .B(n9017), .ZN(n7275)
         );
  INV_X1 U8789 ( .A(n7275), .ZN(n7284) );
  NOR2_X1 U8790 ( .A1(n7276), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8983) );
  OAI21_X1 U8791 ( .B1(n7278), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7277), .ZN(
        n7496) );
  INV_X1 U8792 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7279) );
  NOR2_X1 U8793 ( .A1(n7279), .A2(n7280), .ZN(n7498) );
  AOI211_X1 U8794 ( .C1(n7280), .C2(n7279), .A(n7498), .B(n9030), .ZN(n7281)
         );
  AOI211_X1 U8795 ( .C1(n9610), .C2(n7282), .A(n8983), .B(n7281), .ZN(n7283)
         );
  OAI211_X1 U8796 ( .C1(n9039), .C2(n6093), .A(n7284), .B(n7283), .ZN(P1_U3256) );
  NAND2_X1 U8797 ( .A1(n7285), .A2(n8110), .ZN(n7288) );
  AOI22_X1 U8798 ( .A1(n7795), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7794), .B2(
        n7286), .ZN(n7287) );
  XNOR2_X1 U8799 ( .A(n9864), .B(n6919), .ZN(n7289) );
  NAND2_X1 U8800 ( .A1(n9765), .A2(n8118), .ZN(n7290) );
  NAND2_X1 U8801 ( .A1(n7289), .A2(n7290), .ZN(n7309) );
  INV_X1 U8802 ( .A(n7289), .ZN(n7292) );
  INV_X1 U8803 ( .A(n7290), .ZN(n7291) );
  NAND2_X1 U8804 ( .A1(n7292), .A2(n7291), .ZN(n7311) );
  NAND2_X1 U8805 ( .A1(n7309), .A2(n7311), .ZN(n7298) );
  INV_X1 U8806 ( .A(n7293), .ZN(n7294) );
  NAND2_X1 U8807 ( .A1(n7295), .A2(n7294), .ZN(n7296) );
  XOR2_X1 U8808 ( .A(n7298), .B(n7310), .Z(n7308) );
  NAND2_X1 U8809 ( .A1(n8105), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7302) );
  XNOR2_X1 U8810 ( .A(n7319), .B(P2_REG3_REG_10__SCAN_IN), .ZN(n9742) );
  NAND2_X1 U8811 ( .A1(n7901), .A2(n9742), .ZN(n7301) );
  NAND2_X1 U8812 ( .A1(n6750), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7300) );
  NAND2_X1 U8813 ( .A1(n8106), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7299) );
  NAND4_X1 U8814 ( .A1(n7302), .A2(n7301), .A3(n7300), .A4(n7299), .ZN(n8312)
         );
  AOI22_X1 U8815 ( .A1(n9864), .A2(n8083), .B1(n7986), .B2(n8312), .ZN(n7307)
         );
  INV_X1 U8816 ( .A(n7303), .ZN(n7346) );
  OAI21_X1 U8817 ( .B1(n8080), .B2(n7346), .A(n7304), .ZN(n7305) );
  AOI21_X1 U8818 ( .B1(n7985), .B2(n8313), .A(n7305), .ZN(n7306) );
  OAI211_X1 U8819 ( .C1(n7308), .C2(n8085), .A(n7307), .B(n7306), .ZN(P2_U3233) );
  NAND2_X1 U8820 ( .A1(n7310), .A2(n7309), .ZN(n7312) );
  NAND2_X1 U8821 ( .A1(n7312), .A2(n7311), .ZN(n7446) );
  AOI22_X1 U8822 ( .A1(n7795), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7794), .B2(
        n7313), .ZN(n7316) );
  NAND2_X1 U8823 ( .A1(n7314), .A2(n8110), .ZN(n7315) );
  NAND2_X1 U8824 ( .A1(n7316), .A2(n7315), .ZN(n7516) );
  XNOR2_X1 U8825 ( .A(n7516), .B(n6912), .ZN(n7449) );
  NAND2_X1 U8826 ( .A1(n8312), .A2(n8118), .ZN(n7447) );
  XNOR2_X1 U8827 ( .A(n7449), .B(n7447), .ZN(n7445) );
  XNOR2_X1 U8828 ( .A(n7446), .B(n7445), .ZN(n7330) );
  NAND2_X1 U8829 ( .A1(n8106), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7324) );
  INV_X1 U8830 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7317) );
  OAI21_X1 U8831 ( .B1(n7319), .B2(n7317), .A(n7463), .ZN(n7320) );
  NAND2_X1 U8832 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n7318) );
  AND2_X1 U8833 ( .A1(n7320), .A2(n7457), .ZN(n7517) );
  NAND2_X1 U8834 ( .A1(n7901), .A2(n7517), .ZN(n7323) );
  NAND2_X1 U8835 ( .A1(n6750), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7322) );
  NAND2_X1 U8836 ( .A1(n8105), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7321) );
  NAND4_X1 U8837 ( .A1(n7324), .A2(n7323), .A3(n7322), .A4(n7321), .ZN(n9735)
         );
  INV_X1 U8838 ( .A(n7516), .ZN(n9873) );
  OAI22_X1 U8839 ( .A1(n9703), .A2(n8691), .B1(n9873), .B2(n9701), .ZN(n7328)
         );
  INV_X1 U8840 ( .A(n9742), .ZN(n7326) );
  OAI21_X1 U8841 ( .B1(n8080), .B2(n7326), .A(n7325), .ZN(n7327) );
  AOI211_X1 U8842 ( .C1(n7985), .C2(n9765), .A(n7328), .B(n7327), .ZN(n7329)
         );
  OAI21_X1 U8843 ( .B1(n7330), .B2(n8085), .A(n7329), .ZN(P2_U3219) );
  NAND2_X1 U8844 ( .A1(n7333), .A2(n9850), .ZN(n7334) );
  XNOR2_X1 U8845 ( .A(n8185), .B(n8313), .ZN(n9749) );
  NAND2_X1 U8846 ( .A1(n8185), .A2(n8313), .ZN(n7335) );
  OR2_X1 U8847 ( .A1(n7336), .A2(n9864), .ZN(n8190) );
  NAND2_X1 U8848 ( .A1(n9864), .A2(n7336), .ZN(n8191) );
  NAND2_X1 U8849 ( .A1(n7338), .A2(n7512), .ZN(n7339) );
  NAND2_X1 U8850 ( .A1(n7508), .A2(n7339), .ZN(n9868) );
  INV_X1 U8851 ( .A(n9749), .ZN(n9758) );
  INV_X1 U8852 ( .A(n8313), .ZN(n8186) );
  NAND2_X1 U8853 ( .A1(n8186), .A2(n8185), .ZN(n8183) );
  XNOR2_X1 U8854 ( .A(n7513), .B(n7337), .ZN(n7342) );
  AOI22_X1 U8855 ( .A1(n9762), .A2(n8313), .B1(n8312), .B2(n9764), .ZN(n7341)
         );
  OAI21_X1 U8856 ( .B1(n7342), .B2(n8690), .A(n7341), .ZN(n7343) );
  AOI21_X1 U8857 ( .B1(n9868), .B2(n7344), .A(n7343), .ZN(n9870) );
  NAND2_X1 U8858 ( .A1(n9753), .A2(n9864), .ZN(n7345) );
  NAND2_X1 U8859 ( .A1(n9728), .A2(n7345), .ZN(n9866) );
  OAI22_X1 U8860 ( .A1(n9779), .A2(n6487), .B1(n7346), .B2(n8613), .ZN(n7347)
         );
  AOI21_X1 U8861 ( .B1(n8698), .B2(n9864), .A(n7347), .ZN(n7348) );
  OAI21_X1 U8862 ( .B1(n9754), .B2(n9866), .A(n7348), .ZN(n7349) );
  AOI21_X1 U8863 ( .B1(n9868), .B2(n9734), .A(n7349), .ZN(n7350) );
  OAI21_X1 U8864 ( .B1(n9870), .B2(n9775), .A(n7350), .ZN(P2_U3287) );
  INV_X1 U8865 ( .A(n7865), .ZN(n7353) );
  INV_X1 U8866 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7351) );
  OAI222_X1 U8867 ( .A1(n7352), .A2(P1_U3084), .B1(n9552), .B2(n7353), .C1(
        n7351), .C2(n7705), .ZN(P1_U3329) );
  INV_X1 U8868 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7866) );
  OAI222_X1 U8869 ( .A1(n7354), .A2(P2_U3152), .B1(n7667), .B2(n7353), .C1(
        n7866), .C2(n8830), .ZN(P2_U3334) );
  XOR2_X1 U8870 ( .A(n7355), .B(n7359), .Z(n7362) );
  OAI22_X1 U8871 ( .A1(n9638), .A2(n7379), .B1(n7563), .B2(n9635), .ZN(n7361)
         );
  INV_X1 U8872 ( .A(n7356), .ZN(n7357) );
  AOI21_X1 U8873 ( .B1(n7359), .B2(n7358), .A(n7357), .ZN(n7526) );
  NOR2_X1 U8874 ( .A1(n7526), .A2(n9643), .ZN(n7360) );
  AOI211_X1 U8875 ( .C1(n9640), .C2(n7362), .A(n7361), .B(n7360), .ZN(n7525)
         );
  INV_X1 U8876 ( .A(n7363), .ZN(n7364) );
  AOI211_X1 U8877 ( .C1(n7523), .C2(n7365), .A(n9682), .B(n7364), .ZN(n7522)
         );
  AOI22_X1 U8878 ( .A1(n9647), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7370), .B2(
        n9645), .ZN(n7366) );
  OAI21_X1 U8879 ( .B1(n7380), .B2(n9595), .A(n7366), .ZN(n7368) );
  NOR2_X1 U8880 ( .A1(n7526), .A2(n9585), .ZN(n7367) );
  AOI211_X1 U8881 ( .C1(n7522), .C2(n9406), .A(n7368), .B(n7367), .ZN(n7369)
         );
  OAI21_X1 U8882 ( .B1(n7525), .B2(n9647), .A(n7369), .ZN(P1_U3285) );
  INV_X1 U8883 ( .A(n7370), .ZN(n7385) );
  INV_X1 U8884 ( .A(n7371), .ZN(n7372) );
  NOR3_X1 U8885 ( .A1(n7374), .A2(n7373), .A3(n7372), .ZN(n7377) );
  INV_X1 U8886 ( .A(n7375), .ZN(n7376) );
  OAI21_X1 U8887 ( .B1(n7377), .B2(n7376), .A(n8970), .ZN(n7384) );
  INV_X1 U8888 ( .A(n7378), .ZN(n7382) );
  OAI22_X1 U8889 ( .A1(n8977), .A2(n7380), .B1(n8987), .B2(n7379), .ZN(n7381)
         );
  AOI211_X1 U8890 ( .C1(n8984), .C2(n8998), .A(n7382), .B(n7381), .ZN(n7383)
         );
  OAI211_X1 U8891 ( .C1(n8906), .C2(n7385), .A(n7384), .B(n7383), .ZN(P1_U3237) );
  INV_X1 U8892 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9948) );
  NOR2_X1 U8893 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7386) );
  AOI21_X1 U8894 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7386), .ZN(n9920) );
  NOR2_X1 U8895 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7387) );
  AOI21_X1 U8896 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7387), .ZN(n9923) );
  NOR2_X1 U8897 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n7388) );
  AOI21_X1 U8898 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n7388), .ZN(n9926) );
  NOR2_X1 U8899 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7389) );
  AOI21_X1 U8900 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7389), .ZN(n9929) );
  NOR2_X1 U8901 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7390) );
  AOI21_X1 U8902 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7390), .ZN(n9932) );
  NOR2_X1 U8903 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7397) );
  XNOR2_X1 U8904 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9960) );
  NAND2_X1 U8905 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7395) );
  XOR2_X1 U8906 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n9958) );
  NAND2_X1 U8907 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7393) );
  XNOR2_X1 U8908 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n7391), .ZN(n9956) );
  AOI21_X1 U8909 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9913) );
  INV_X1 U8910 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9917) );
  NAND3_X1 U8911 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9915) );
  OAI21_X1 U8912 ( .B1(n9913), .B2(n9917), .A(n9915), .ZN(n9955) );
  NAND2_X1 U8913 ( .A1(n9956), .A2(n9955), .ZN(n7392) );
  NAND2_X1 U8914 ( .A1(n7393), .A2(n7392), .ZN(n9957) );
  NAND2_X1 U8915 ( .A1(n9958), .A2(n9957), .ZN(n7394) );
  NAND2_X1 U8916 ( .A1(n7395), .A2(n7394), .ZN(n9959) );
  NOR2_X1 U8917 ( .A1(n9960), .A2(n9959), .ZN(n7396) );
  NOR2_X1 U8918 ( .A1(n7397), .A2(n7396), .ZN(n7398) );
  NOR2_X1 U8919 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7398), .ZN(n9944) );
  AND2_X1 U8920 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7398), .ZN(n9943) );
  NOR2_X1 U8921 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9943), .ZN(n7399) );
  NOR2_X1 U8922 ( .A1(n9944), .A2(n7399), .ZN(n7400) );
  NAND2_X1 U8923 ( .A1(n7400), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7402) );
  XOR2_X1 U8924 ( .A(n7400), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n9942) );
  NAND2_X1 U8925 ( .A1(n9942), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7401) );
  NAND2_X1 U8926 ( .A1(n7402), .A2(n7401), .ZN(n7403) );
  NAND2_X1 U8927 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7403), .ZN(n7405) );
  XOR2_X1 U8928 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7403), .Z(n9954) );
  NAND2_X1 U8929 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n9954), .ZN(n7404) );
  NAND2_X1 U8930 ( .A1(n7405), .A2(n7404), .ZN(n7406) );
  NAND2_X1 U8931 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7406), .ZN(n7408) );
  XOR2_X1 U8932 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7406), .Z(n9953) );
  NAND2_X1 U8933 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n9953), .ZN(n7407) );
  NAND2_X1 U8934 ( .A1(n7408), .A2(n7407), .ZN(n7409) );
  AND2_X1 U8935 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7409), .ZN(n7410) );
  XNOR2_X1 U8936 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7409), .ZN(n9951) );
  NOR2_X1 U8937 ( .A1(n9952), .A2(n9951), .ZN(n9950) );
  NAND2_X1 U8938 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7411) );
  OAI21_X1 U8939 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7411), .ZN(n9940) );
  NAND2_X1 U8940 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7412) );
  OAI21_X1 U8941 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7412), .ZN(n9937) );
  NOR2_X1 U8942 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7413) );
  AOI21_X1 U8943 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7413), .ZN(n9934) );
  NAND2_X1 U8944 ( .A1(n9935), .A2(n9934), .ZN(n9933) );
  NAND2_X1 U8945 ( .A1(n9932), .A2(n9931), .ZN(n9930) );
  NAND2_X1 U8946 ( .A1(n9929), .A2(n9928), .ZN(n9927) );
  OAI21_X1 U8947 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9927), .ZN(n9925) );
  NAND2_X1 U8948 ( .A1(n9926), .A2(n9925), .ZN(n9924) );
  OAI21_X1 U8949 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9924), .ZN(n9922) );
  NAND2_X1 U8950 ( .A1(n9923), .A2(n9922), .ZN(n9921) );
  OAI21_X1 U8951 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9921), .ZN(n9919) );
  NAND2_X1 U8952 ( .A1(n9920), .A2(n9919), .ZN(n9918) );
  OAI21_X1 U8953 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9918), .ZN(n9947) );
  NOR2_X1 U8954 ( .A1(n9948), .A2(n9947), .ZN(n7414) );
  NAND2_X1 U8955 ( .A1(n9948), .A2(n9947), .ZN(n9946) );
  OAI21_X1 U8956 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7414), .A(n9946), .ZN(
        n7416) );
  XNOR2_X1 U8957 ( .A(n9040), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7415) );
  XNOR2_X1 U8958 ( .A(n7416), .B(n7415), .ZN(ADD_1071_U4) );
  INV_X1 U8959 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7418) );
  AOI211_X1 U8960 ( .C1(n7419), .C2(n7418), .A(n8323), .B(n9718), .ZN(n7429)
         );
  AOI21_X1 U8961 ( .B1(n7422), .B2(n7421), .A(n7420), .ZN(n8329) );
  XNOR2_X1 U8962 ( .A(n8329), .B(n8330), .ZN(n7423) );
  NOR2_X1 U8963 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7423), .ZN(n8331) );
  AOI21_X1 U8964 ( .B1(n7423), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8331), .ZN(
        n7424) );
  NOR2_X1 U8965 ( .A1(n7424), .A2(n9716), .ZN(n7428) );
  INV_X1 U8966 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8078) );
  NOR2_X1 U8967 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8078), .ZN(n7425) );
  AOI21_X1 U8968 ( .B1(n9715), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7425), .ZN(
        n7426) );
  OAI21_X1 U8969 ( .B1(n9717), .B2(n8322), .A(n7426), .ZN(n7427) );
  OR3_X1 U8970 ( .A1(n7429), .A2(n7428), .A3(n7427), .ZN(P2_U3260) );
  INV_X1 U8971 ( .A(n7430), .ZN(n7435) );
  AOI21_X1 U8972 ( .B1(n7432), .B2(n7434), .A(n7431), .ZN(n7433) );
  AOI21_X1 U8973 ( .B1(n7435), .B2(n7434), .A(n7433), .ZN(n7444) );
  INV_X1 U8974 ( .A(n7436), .ZN(n7437) );
  AOI21_X1 U8975 ( .B1(n8984), .B2(n8997), .A(n7437), .ZN(n7440) );
  OR2_X1 U8976 ( .A1(n8987), .A2(n7438), .ZN(n7439) );
  OAI211_X1 U8977 ( .C1(n9675), .C2(n8977), .A(n7440), .B(n7439), .ZN(n7441)
         );
  AOI21_X1 U8978 ( .B1(n7442), .B2(n8982), .A(n7441), .ZN(n7443) );
  OAI21_X1 U8979 ( .B1(n7444), .B2(n8991), .A(n7443), .ZN(P1_U3211) );
  NAND2_X1 U8980 ( .A1(n7446), .A2(n7445), .ZN(n7451) );
  INV_X1 U8981 ( .A(n7447), .ZN(n7448) );
  NAND2_X1 U8982 ( .A1(n7449), .A2(n7448), .ZN(n7450) );
  NAND2_X1 U8983 ( .A1(n7451), .A2(n7450), .ZN(n7532) );
  NAND2_X1 U8984 ( .A1(n7452), .A2(n8110), .ZN(n7455) );
  AOI22_X1 U8985 ( .A1(n7795), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7794), .B2(
        n7453), .ZN(n7454) );
  NAND2_X1 U8986 ( .A1(n7455), .A2(n7454), .ZN(n8400) );
  XNOR2_X1 U8987 ( .A(n8400), .B(n6912), .ZN(n7535) );
  NAND2_X1 U8988 ( .A1(n9735), .A2(n8118), .ZN(n7533) );
  XNOR2_X1 U8989 ( .A(n7535), .B(n7533), .ZN(n7531) );
  XNOR2_X1 U8990 ( .A(n7532), .B(n7531), .ZN(n7468) );
  NAND2_X1 U8991 ( .A1(n8105), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7462) );
  INV_X1 U8992 ( .A(n7457), .ZN(n7456) );
  NAND2_X1 U8993 ( .A1(n7456), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7583) );
  NAND2_X1 U8994 ( .A1(n7457), .A2(n7546), .ZN(n7458) );
  AND2_X1 U8995 ( .A1(n7583), .A2(n7458), .ZN(n8696) );
  NAND2_X1 U8996 ( .A1(n7901), .A2(n8696), .ZN(n7461) );
  NAND2_X1 U8997 ( .A1(n6750), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7460) );
  NAND2_X1 U8998 ( .A1(n8106), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7459) );
  NAND4_X1 U8999 ( .A1(n7462), .A2(n7461), .A3(n7460), .A4(n7459), .ZN(n8403)
         );
  INV_X1 U9000 ( .A(n8400), .ZN(n9881) );
  OAI22_X1 U9001 ( .A1(n9703), .A2(n8669), .B1(n9881), .B2(n9701), .ZN(n7466)
         );
  INV_X1 U9002 ( .A(n7517), .ZN(n7464) );
  OAI22_X1 U9003 ( .A1(n8080), .A2(n7464), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7463), .ZN(n7465) );
  AOI211_X1 U9004 ( .C1(n7985), .C2(n8312), .A(n7466), .B(n7465), .ZN(n7467)
         );
  OAI21_X1 U9005 ( .B1(n7468), .B2(n8085), .A(n7467), .ZN(P2_U3238) );
  INV_X1 U9006 ( .A(n7880), .ZN(n7471) );
  OAI222_X1 U9007 ( .A1(n8830), .A2(n7881), .B1(n7667), .B2(n7471), .C1(n7469), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI222_X1 U9008 ( .A1(P1_U3084), .A2(n7472), .B1(n9552), .B2(n7471), .C1(
        n7470), .C2(n7705), .ZN(P1_U3328) );
  XNOR2_X1 U9009 ( .A(n7474), .B(n7478), .ZN(n7483) );
  OAI22_X1 U9010 ( .A1(n9638), .A2(n7563), .B1(n7661), .B2(n9635), .ZN(n7482)
         );
  NAND2_X1 U9011 ( .A1(n7563), .A2(n9675), .ZN(n7475) );
  NAND2_X1 U9012 ( .A1(n7479), .A2(n7478), .ZN(n7480) );
  NAND2_X1 U9013 ( .A1(n7477), .A2(n7480), .ZN(n7597) );
  NOR2_X1 U9014 ( .A1(n7597), .A2(n9643), .ZN(n7481) );
  AOI211_X1 U9015 ( .C1(n7483), .C2(n9640), .A(n7482), .B(n7481), .ZN(n7596)
         );
  AOI21_X1 U9016 ( .B1(n7603), .B2(n7485), .A(n4336), .ZN(n7594) );
  AOI22_X1 U9017 ( .A1(n9647), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7558), .B2(
        n9645), .ZN(n7486) );
  OAI21_X1 U9018 ( .B1(n7557), .B2(n9595), .A(n7486), .ZN(n7488) );
  NOR2_X1 U9019 ( .A1(n7597), .A2(n9585), .ZN(n7487) );
  AOI211_X1 U9020 ( .C1(n7594), .C2(n9631), .A(n7488), .B(n7487), .ZN(n7489)
         );
  OAI21_X1 U9021 ( .B1(n7596), .B2(n9647), .A(n7489), .ZN(P1_U3283) );
  NOR2_X1 U9022 ( .A1(n7490), .A2(n7497), .ZN(n7492) );
  NOR2_X1 U9023 ( .A1(n7492), .A2(n7491), .ZN(n7495) );
  NAND2_X1 U9024 ( .A1(n7644), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7493) );
  OAI21_X1 U9025 ( .B1(n7644), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7493), .ZN(
        n7494) );
  NOR2_X1 U9026 ( .A1(n7495), .A2(n7494), .ZN(n7643) );
  AOI211_X1 U9027 ( .C1(n7495), .C2(n7494), .A(n7643), .B(n9017), .ZN(n7506)
         );
  NOR2_X1 U9028 ( .A1(n7497), .A2(n7496), .ZN(n7499) );
  NOR2_X1 U9029 ( .A1(n7499), .A2(n7498), .ZN(n7501) );
  XNOR2_X1 U9030 ( .A(n7644), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7500) );
  NOR2_X1 U9031 ( .A1(n7501), .A2(n7500), .ZN(n7639) );
  AOI211_X1 U9032 ( .C1(n7501), .C2(n7500), .A(n7639), .B(n9030), .ZN(n7505)
         );
  NAND2_X1 U9033 ( .A1(n9611), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7502) );
  NAND2_X1 U9034 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8897) );
  OAI211_X1 U9035 ( .C1(n7503), .C2(n9029), .A(n7502), .B(n8897), .ZN(n7504)
         );
  OR3_X1 U9036 ( .A1(n7506), .A2(n7505), .A3(n7504), .ZN(P1_U3257) );
  OR2_X1 U9037 ( .A1(n9864), .A2(n9765), .ZN(n7507) );
  NAND2_X1 U9038 ( .A1(n9873), .A2(n8312), .ZN(n8197) );
  INV_X1 U9039 ( .A(n8312), .ZN(n7515) );
  NAND2_X1 U9040 ( .A1(n7515), .A2(n7516), .ZN(n8199) );
  NAND2_X1 U9041 ( .A1(n7516), .A2(n8312), .ZN(n7510) );
  OR2_X1 U9042 ( .A1(n8400), .A2(n8691), .ZN(n8204) );
  NAND2_X1 U9043 ( .A1(n8400), .A2(n8691), .ZN(n8208) );
  NAND2_X1 U9044 ( .A1(n8204), .A2(n8208), .ZN(n8132) );
  NAND2_X1 U9045 ( .A1(n7511), .A2(n8132), .ZN(n8402) );
  OAI21_X1 U9046 ( .B1(n7511), .B2(n8132), .A(n8402), .ZN(n9880) );
  INV_X1 U9047 ( .A(n8191), .ZN(n8189) );
  NAND2_X1 U9048 ( .A1(n9738), .A2(n9737), .ZN(n9736) );
  NAND2_X1 U9049 ( .A1(n9736), .A2(n8197), .ZN(n8088) );
  XOR2_X1 U9050 ( .A(n8132), .B(n8088), .Z(n7514) );
  OAI222_X1 U9051 ( .A1(n8694), .A2(n8669), .B1(n8692), .B2(n7515), .C1(n8690), 
        .C2(n7514), .ZN(n9883) );
  XNOR2_X1 U9052 ( .A(n9729), .B(n9881), .ZN(n9882) );
  AOI22_X1 U9053 ( .A1(n9775), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7517), .B2(
        n9773), .ZN(n7519) );
  NAND2_X1 U9054 ( .A1(n8698), .A2(n8400), .ZN(n7518) );
  OAI211_X1 U9055 ( .C1(n9882), .C2(n9754), .A(n7519), .B(n7518), .ZN(n7520)
         );
  AOI21_X1 U9056 ( .B1(n9883), .B2(n9779), .A(n7520), .ZN(n7521) );
  OAI21_X1 U9057 ( .B1(n8703), .B2(n9880), .A(n7521), .ZN(P2_U3285) );
  AOI21_X1 U9058 ( .B1(n9568), .B2(n7523), .A(n7522), .ZN(n7524) );
  OAI211_X1 U9059 ( .C1(n7526), .C2(n9510), .A(n7525), .B(n7524), .ZN(n7528)
         );
  NAND2_X1 U9060 ( .A1(n7528), .A2(n9697), .ZN(n7527) );
  OAI21_X1 U9061 ( .B1(n9697), .B2(n6005), .A(n7527), .ZN(P1_U3529) );
  NAND2_X1 U9062 ( .A1(n7528), .A2(n9530), .ZN(n7529) );
  OAI21_X1 U9063 ( .B1(n9530), .B2(n7530), .A(n7529), .ZN(P1_U3472) );
  NAND2_X1 U9064 ( .A1(n7532), .A2(n7531), .ZN(n7537) );
  INV_X1 U9065 ( .A(n7533), .ZN(n7534) );
  NAND2_X1 U9066 ( .A1(n7535), .A2(n7534), .ZN(n7536) );
  NAND2_X1 U9067 ( .A1(n7537), .A2(n7536), .ZN(n7571) );
  NAND2_X1 U9068 ( .A1(n7538), .A2(n8110), .ZN(n7541) );
  AOI22_X1 U9069 ( .A1(n7795), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7794), .B2(
        n7539), .ZN(n7540) );
  NAND2_X1 U9070 ( .A1(n7541), .A2(n7540), .ZN(n8697) );
  XNOR2_X1 U9071 ( .A(n8697), .B(n6912), .ZN(n7574) );
  NAND2_X1 U9072 ( .A1(n8403), .A2(n8118), .ZN(n7572) );
  XNOR2_X1 U9073 ( .A(n7574), .B(n7572), .ZN(n7570) );
  XNOR2_X1 U9074 ( .A(n7571), .B(n7570), .ZN(n7551) );
  NAND2_X1 U9075 ( .A1(n8106), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7545) );
  XNOR2_X1 U9076 ( .A(n7583), .B(P2_REG3_REG_13__SCAN_IN), .ZN(n8678) );
  NAND2_X1 U9077 ( .A1(n7901), .A2(n8678), .ZN(n7544) );
  NAND2_X1 U9078 ( .A1(n6750), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7543) );
  NAND2_X1 U9079 ( .A1(n8105), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7542) );
  NAND4_X1 U9080 ( .A1(n7545), .A2(n7544), .A3(n7543), .A4(n7542), .ZN(n8405)
         );
  OAI22_X1 U9081 ( .A1(n8691), .A2(n9704), .B1(n9703), .B2(n8693), .ZN(n7549)
         );
  INV_X1 U9082 ( .A(n8696), .ZN(n7547) );
  OAI22_X1 U9083 ( .A1(n8080), .A2(n7547), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7546), .ZN(n7548) );
  AOI211_X1 U9084 ( .C1(n8697), .C2(n8083), .A(n7549), .B(n7548), .ZN(n7550)
         );
  OAI21_X1 U9085 ( .B1(n7551), .B2(n8085), .A(n7550), .ZN(P2_U3226) );
  INV_X1 U9086 ( .A(n7894), .ZN(n7568) );
  AOI22_X1 U9087 ( .A1(n5916), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n9549), .ZN(n7552) );
  OAI21_X1 U9088 ( .B1(n7568), .B2(n9552), .A(n7552), .ZN(P1_U3327) );
  NAND2_X1 U9089 ( .A1(n7553), .A2(n7554), .ZN(n7556) );
  XNOR2_X1 U9090 ( .A(n7556), .B(n7555), .ZN(n7566) );
  NOR2_X1 U9091 ( .A1(n8977), .A2(n7557), .ZN(n7565) );
  NAND2_X1 U9092 ( .A1(n8982), .A2(n7558), .ZN(n7562) );
  INV_X1 U9093 ( .A(n7559), .ZN(n7560) );
  AOI21_X1 U9094 ( .B1(n8984), .B2(n8996), .A(n7560), .ZN(n7561) );
  OAI211_X1 U9095 ( .C1(n7563), .C2(n8987), .A(n7562), .B(n7561), .ZN(n7564)
         );
  AOI211_X1 U9096 ( .C1(n7566), .C2(n8970), .A(n7565), .B(n7564), .ZN(n7567)
         );
  INV_X1 U9097 ( .A(n7567), .ZN(P1_U3219) );
  OAI222_X1 U9098 ( .A1(n7569), .A2(P2_U3152), .B1(n7667), .B2(n7568), .C1(
        n7895), .C2(n8830), .ZN(P2_U3332) );
  NAND2_X1 U9099 ( .A1(n7571), .A2(n7570), .ZN(n7576) );
  INV_X1 U9100 ( .A(n7572), .ZN(n7573) );
  NAND2_X1 U9101 ( .A1(n7574), .A2(n7573), .ZN(n7575) );
  NAND2_X1 U9102 ( .A1(n7577), .A2(n8110), .ZN(n7580) );
  AOI22_X1 U9103 ( .A1(n7795), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7794), .B2(
        n7578), .ZN(n7579) );
  XNOR2_X1 U9104 ( .A(n8797), .B(n6912), .ZN(n7723) );
  NAND2_X1 U9105 ( .A1(n8405), .A2(n8118), .ZN(n7721) );
  XNOR2_X1 U9106 ( .A(n7723), .B(n7721), .ZN(n7719) );
  XNOR2_X1 U9107 ( .A(n7720), .B(n7719), .ZN(n7593) );
  NAND2_X1 U9108 ( .A1(n8106), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7588) );
  NAND2_X1 U9109 ( .A1(n6750), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7587) );
  INV_X1 U9110 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7581) );
  OAI21_X1 U9111 ( .B1(n7583), .B2(n7582), .A(n7581), .ZN(n7584) );
  AND2_X1 U9112 ( .A1(n7584), .A2(n7747), .ZN(n8654) );
  NAND2_X1 U9113 ( .A1(n7901), .A2(n8654), .ZN(n7586) );
  NAND2_X1 U9114 ( .A1(n8105), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7585) );
  NAND4_X1 U9115 ( .A1(n7588), .A2(n7587), .A3(n7586), .A4(n7585), .ZN(n8407)
         );
  OAI22_X1 U9116 ( .A1(n8669), .A2(n9704), .B1(n9703), .B2(n8668), .ZN(n7591)
         );
  INV_X1 U9117 ( .A(n8678), .ZN(n7589) );
  OAI22_X1 U9118 ( .A1(n8080), .A2(n7589), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7582), .ZN(n7590) );
  AOI211_X1 U9119 ( .C1(n8797), .C2(n8083), .A(n7591), .B(n7590), .ZN(n7592)
         );
  OAI21_X1 U9120 ( .B1(n7593), .B2(n8085), .A(n7592), .ZN(P2_U3236) );
  AOI22_X1 U9121 ( .A1(n7594), .A2(n9500), .B1(n9568), .B2(n7603), .ZN(n7595)
         );
  OAI211_X1 U9122 ( .C1(n9510), .C2(n7597), .A(n7596), .B(n7595), .ZN(n7600)
         );
  NAND2_X1 U9123 ( .A1(n7600), .A2(n9697), .ZN(n7598) );
  OAI21_X1 U9124 ( .B1(n9697), .B2(n7599), .A(n7598), .ZN(P1_U3531) );
  INV_X1 U9125 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7602) );
  NAND2_X1 U9126 ( .A1(n7600), .A2(n9530), .ZN(n7601) );
  OAI21_X1 U9127 ( .B1(n9530), .B2(n7602), .A(n7601), .ZN(P1_U3478) );
  NAND2_X1 U9128 ( .A1(n8997), .A2(n7603), .ZN(n7604) );
  NAND2_X1 U9129 ( .A1(n7605), .A2(n7604), .ZN(n9628) );
  AND2_X1 U9130 ( .A1(n8996), .A2(n7635), .ZN(n7606) );
  OAI22_X2 U9131 ( .A1(n9628), .A2(n7606), .B1(n8996), .B2(n7635), .ZN(n9053)
         );
  XOR2_X1 U9132 ( .A(n9053), .B(n9052), .Z(n9567) );
  AOI22_X1 U9133 ( .A1(n9056), .A2(n9309), .B1(n9311), .B2(n8996), .ZN(n7618)
         );
  NAND2_X1 U9134 ( .A1(n7611), .A2(n7610), .ZN(n9094) );
  INV_X1 U9135 ( .A(n7611), .ZN(n7614) );
  INV_X1 U9136 ( .A(n7612), .ZN(n7613) );
  OAI21_X1 U9137 ( .B1(n7614), .B2(n7613), .A(n9052), .ZN(n7615) );
  OAI211_X1 U9138 ( .C1(n7616), .C2(n9094), .A(n7615), .B(n9640), .ZN(n7617)
         );
  OAI211_X1 U9139 ( .C1(n9567), .C2(n9643), .A(n7618), .B(n7617), .ZN(n9571)
         );
  NAND2_X1 U9140 ( .A1(n9571), .A2(n9650), .ZN(n7626) );
  INV_X1 U9141 ( .A(n9629), .ZN(n7621) );
  INV_X1 U9142 ( .A(n9581), .ZN(n7620) );
  OAI211_X1 U9143 ( .C1(n9570), .C2(n7621), .A(n7620), .B(n9500), .ZN(n9569)
         );
  INV_X1 U9144 ( .A(n9569), .ZN(n7624) );
  AOI22_X1 U9145 ( .A1(n9647), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7656), .B2(
        n9645), .ZN(n7622) );
  OAI21_X1 U9146 ( .B1(n9570), .B2(n9595), .A(n7622), .ZN(n7623) );
  AOI21_X1 U9147 ( .B1(n7624), .B2(n9406), .A(n7623), .ZN(n7625) );
  OAI211_X1 U9148 ( .C1(n9567), .C2(n9585), .A(n7626), .B(n7625), .ZN(P1_U3281) );
  INV_X1 U9149 ( .A(n7628), .ZN(n7629) );
  AOI21_X1 U9150 ( .B1(n7630), .B2(n7627), .A(n7629), .ZN(n7637) );
  NAND2_X1 U9151 ( .A1(n8982), .A2(n9646), .ZN(n7633) );
  AOI21_X1 U9152 ( .B1(n8984), .B2(n8995), .A(n7631), .ZN(n7632) );
  OAI211_X1 U9153 ( .C1(n9637), .C2(n8987), .A(n7633), .B(n7632), .ZN(n7634)
         );
  AOI21_X1 U9154 ( .B1(n7635), .B2(n8989), .A(n7634), .ZN(n7636) );
  OAI21_X1 U9155 ( .B1(n7637), .B2(n8991), .A(n7636), .ZN(P1_U3229) );
  INV_X1 U9156 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7651) );
  NOR2_X1 U9157 ( .A1(n7638), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7680) );
  AOI21_X1 U9158 ( .B1(n7644), .B2(P1_REG1_REG_16__SCAN_IN), .A(n7639), .ZN(
        n7641) );
  XNOR2_X1 U9159 ( .A(n9015), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n7640) );
  NOR2_X1 U9160 ( .A1(n7641), .A2(n7640), .ZN(n9007) );
  AOI211_X1 U9161 ( .C1(n7641), .C2(n7640), .A(n9007), .B(n9030), .ZN(n7642)
         );
  AOI211_X1 U9162 ( .C1(n9015), .C2(n9610), .A(n7680), .B(n7642), .ZN(n7650)
         );
  AOI21_X1 U9163 ( .B1(n7644), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7643), .ZN(
        n7647) );
  NAND2_X1 U9164 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9015), .ZN(n7645) );
  OAI21_X1 U9165 ( .B1(n9015), .B2(P1_REG2_REG_17__SCAN_IN), .A(n7645), .ZN(
        n7646) );
  NOR2_X1 U9166 ( .A1(n7647), .A2(n7646), .ZN(n9014) );
  AOI211_X1 U9167 ( .C1(n7647), .C2(n7646), .A(n9014), .B(n9017), .ZN(n7648)
         );
  INV_X1 U9168 ( .A(n7648), .ZN(n7649) );
  OAI211_X1 U9169 ( .C1(n7651), .C2(n9039), .A(n7650), .B(n7649), .ZN(P1_U3258) );
  XNOR2_X1 U9170 ( .A(n7653), .B(n7652), .ZN(n7654) );
  XNOR2_X1 U9171 ( .A(n7655), .B(n7654), .ZN(n7664) );
  NOR2_X1 U9172 ( .A1(n8977), .A2(n9570), .ZN(n7663) );
  NAND2_X1 U9173 ( .A1(n8982), .A2(n7656), .ZN(n7660) );
  INV_X1 U9174 ( .A(n7657), .ZN(n7658) );
  AOI21_X1 U9175 ( .B1(n8984), .B2(n9056), .A(n7658), .ZN(n7659) );
  OAI211_X1 U9176 ( .C1(n7661), .C2(n8987), .A(n7660), .B(n7659), .ZN(n7662)
         );
  AOI211_X1 U9177 ( .C1(n7664), .C2(n8970), .A(n7663), .B(n7662), .ZN(n7665)
         );
  INV_X1 U9178 ( .A(n7665), .ZN(P1_U3215) );
  INV_X1 U9179 ( .A(n8101), .ZN(n9542) );
  OAI222_X1 U9180 ( .A1(n8830), .A2(n8102), .B1(n7667), .B2(n9542), .C1(n7666), 
        .C2(P2_U3152), .ZN(P2_U3328) );
  INV_X1 U9181 ( .A(n8097), .ZN(n9545) );
  INV_X1 U9182 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8098) );
  OAI222_X1 U9183 ( .A1(n7667), .A2(n9545), .B1(P2_U3152), .B2(n6219), .C1(
        n8098), .C2(n8830), .ZN(P2_U3329) );
  OAI222_X1 U9184 ( .A1(n8830), .A2(n7840), .B1(n7667), .B2(n7668), .C1(n6470), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  XNOR2_X1 U9185 ( .A(n7669), .B(n7670), .ZN(n7676) );
  INV_X1 U9186 ( .A(n9589), .ZN(n9058) );
  NAND2_X1 U9187 ( .A1(n8984), .A2(n9058), .ZN(n7672) );
  OAI211_X1 U9188 ( .C1(n8987), .C2(n9636), .A(n7672), .B(n7671), .ZN(n7673)
         );
  AOI21_X1 U9189 ( .B1(n9593), .B2(n8982), .A(n7673), .ZN(n7675) );
  NAND2_X1 U9190 ( .A1(n8989), .A2(n9055), .ZN(n7674) );
  OAI211_X1 U9191 ( .C1(n7676), .C2(n8991), .A(n7675), .B(n7674), .ZN(P1_U3234) );
  XNOR2_X1 U9192 ( .A(n7678), .B(n7677), .ZN(n7679) );
  XNOR2_X1 U9193 ( .A(n8953), .B(n7679), .ZN(n7685) );
  NAND2_X1 U9194 ( .A1(n8982), .A2(n9305), .ZN(n7682) );
  INV_X1 U9195 ( .A(n9275), .ZN(n9310) );
  AOI21_X1 U9196 ( .B1(n8984), .B2(n9310), .A(n7680), .ZN(n7681) );
  OAI211_X1 U9197 ( .C1(n9336), .C2(n8987), .A(n7682), .B(n7681), .ZN(n7683)
         );
  AOI21_X1 U9198 ( .B1(n9476), .B2(n8989), .A(n7683), .ZN(n7684) );
  OAI21_X1 U9199 ( .B1(n7685), .B2(n8991), .A(n7684), .ZN(P1_U3226) );
  NAND2_X1 U9200 ( .A1(n9423), .A2(n5743), .ZN(n7687) );
  NAND2_X1 U9201 ( .A1(n9090), .A2(n7689), .ZN(n7686) );
  NAND2_X1 U9202 ( .A1(n7687), .A2(n7686), .ZN(n7688) );
  XNOR2_X1 U9203 ( .A(n7688), .B(n5708), .ZN(n7692) );
  NAND2_X1 U9204 ( .A1(n9423), .A2(n7689), .ZN(n7690) );
  OAI21_X1 U9205 ( .B1(n9089), .B2(n5721), .A(n7690), .ZN(n7691) );
  XNOR2_X1 U9206 ( .A(n7692), .B(n7691), .ZN(n7693) );
  INV_X1 U9207 ( .A(n7693), .ZN(n7698) );
  NAND3_X1 U9208 ( .A1(n7698), .A2(n8970), .A3(n7697), .ZN(n7703) );
  NAND3_X1 U9209 ( .A1(n7704), .A2(n8970), .A3(n7693), .ZN(n7702) );
  AOI22_X1 U9210 ( .A1(n8993), .A2(n8984), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n7696) );
  INV_X1 U9211 ( .A(n7694), .ZN(n9146) );
  NAND2_X1 U9212 ( .A1(n8982), .A2(n9146), .ZN(n7695) );
  OAI211_X1 U9213 ( .C1(n9143), .C2(n8987), .A(n7696), .B(n7695), .ZN(n7700)
         );
  NOR3_X1 U9214 ( .A1(n7698), .A2(n8991), .A3(n7697), .ZN(n7699) );
  AOI211_X1 U9215 ( .C1(n9423), .C2(n8989), .A(n7700), .B(n7699), .ZN(n7701)
         );
  OAI211_X1 U9216 ( .C1(n7704), .C2(n7703), .A(n7702), .B(n7701), .ZN(P1_U3218) );
  INV_X1 U9217 ( .A(n7968), .ZN(n9548) );
  OAI222_X1 U9218 ( .A1(n8830), .A2(n7969), .B1(P2_U3152), .B2(n6460), .C1(
        n7667), .C2(n9548), .ZN(P2_U3330) );
  OAI222_X1 U9219 ( .A1(n5670), .A2(P1_U3084), .B1(n9552), .B2(n7707), .C1(
        n7706), .C2(n7705), .ZN(P1_U3332) );
  OAI211_X1 U9220 ( .C1(n7710), .C2(n7709), .A(n7708), .B(n9709), .ZN(n7716)
         );
  AOI22_X1 U9221 ( .A1(n7711), .A2(n8083), .B1(n7986), .B2(n8313), .ZN(n7715)
         );
  AOI22_X1 U9222 ( .A1(n8073), .A2(n7712), .B1(P2_REG3_REG_7__SCAN_IN), .B2(
        P2_U3152), .ZN(n7714) );
  NAND2_X1 U9223 ( .A1(n7985), .A2(n8314), .ZN(n7713) );
  NAND4_X1 U9224 ( .A1(n7716), .A2(n7715), .A3(n7714), .A4(n7713), .ZN(
        P2_U3215) );
  NAND2_X1 U9225 ( .A1(n8827), .A2(n8110), .ZN(n7718) );
  OR2_X1 U9226 ( .A1(n8111), .A2(n8829), .ZN(n7717) );
  INV_X1 U9227 ( .A(n8725), .ZN(n8460) );
  INV_X1 U9228 ( .A(n7721), .ZN(n7722) );
  NAND2_X1 U9229 ( .A1(n7723), .A2(n7722), .ZN(n7724) );
  NAND2_X1 U9230 ( .A1(n7725), .A2(n8110), .ZN(n7728) );
  AOI22_X1 U9231 ( .A1(n7795), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7794), .B2(
        n7726), .ZN(n7727) );
  XNOR2_X1 U9232 ( .A(n8791), .B(n6919), .ZN(n7729) );
  NAND2_X1 U9233 ( .A1(n8407), .A2(n8118), .ZN(n7730) );
  NAND2_X1 U9234 ( .A1(n7729), .A2(n7730), .ZN(n7735) );
  INV_X1 U9235 ( .A(n7729), .ZN(n7732) );
  INV_X1 U9236 ( .A(n7730), .ZN(n7731) );
  NAND2_X1 U9237 ( .A1(n7732), .A2(n7731), .ZN(n7733) );
  NAND2_X1 U9238 ( .A1(n7735), .A2(n7733), .ZN(n7940) );
  NAND2_X1 U9239 ( .A1(n7736), .A2(n8110), .ZN(n7738) );
  AOI22_X1 U9240 ( .A1(n7795), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7794), .B2(
        n8349), .ZN(n7737) );
  XNOR2_X1 U9241 ( .A(n8781), .B(n6919), .ZN(n7757) );
  NAND2_X1 U9242 ( .A1(n8105), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7743) );
  INV_X1 U9243 ( .A(n7747), .ZN(n7739) );
  NAND2_X1 U9244 ( .A1(n7739), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7767) );
  XNOR2_X1 U9245 ( .A(n7767), .B(P2_REG3_REG_16__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U9246 ( .A1(n7141), .A2(n8628), .ZN(n7742) );
  NAND2_X1 U9247 ( .A1(n6750), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7741) );
  NAND2_X1 U9248 ( .A1(n8106), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7740) );
  NAND4_X1 U9249 ( .A1(n7743), .A2(n7742), .A3(n7741), .A4(n7740), .ZN(n8411)
         );
  NAND2_X1 U9250 ( .A1(n8411), .A2(n8118), .ZN(n7758) );
  AND2_X1 U9251 ( .A1(n7757), .A2(n7758), .ZN(n7754) );
  NAND2_X1 U9252 ( .A1(n7744), .A2(n8110), .ZN(n7746) );
  AOI22_X1 U9253 ( .A1(n7795), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7794), .B2(
        n8330), .ZN(n7745) );
  XNOR2_X1 U9254 ( .A(n8786), .B(n6919), .ZN(n8007) );
  NAND2_X1 U9255 ( .A1(n8106), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7752) );
  NAND2_X1 U9256 ( .A1(n6750), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7751) );
  NAND2_X1 U9257 ( .A1(n7747), .A2(n8078), .ZN(n7748) );
  AND2_X1 U9258 ( .A1(n7767), .A2(n7748), .ZN(n8638) );
  NAND2_X1 U9259 ( .A1(n7901), .A2(n8638), .ZN(n7750) );
  NAND2_X1 U9260 ( .A1(n8105), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7749) );
  NAND4_X1 U9261 ( .A1(n7752), .A2(n7751), .A3(n7750), .A4(n7749), .ZN(n8409)
         );
  NAND2_X1 U9262 ( .A1(n8409), .A2(n8118), .ZN(n8076) );
  AND2_X1 U9263 ( .A1(n8007), .A2(n8076), .ZN(n7753) );
  INV_X1 U9264 ( .A(n7754), .ZN(n8009) );
  INV_X1 U9265 ( .A(n8076), .ZN(n7756) );
  INV_X1 U9266 ( .A(n8007), .ZN(n7755) );
  NAND3_X1 U9267 ( .A1(n8009), .A2(n7756), .A3(n7755), .ZN(n7761) );
  INV_X1 U9268 ( .A(n7757), .ZN(n7760) );
  INV_X1 U9269 ( .A(n7758), .ZN(n7759) );
  NAND2_X1 U9270 ( .A1(n7760), .A2(n7759), .ZN(n8008) );
  AND2_X1 U9271 ( .A1(n7761), .A2(n8008), .ZN(n7762) );
  NAND2_X1 U9272 ( .A1(n7764), .A2(n8110), .ZN(n7766) );
  AOI22_X1 U9273 ( .A1(n7795), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7794), .B2(
        n8363), .ZN(n7765) );
  XNOR2_X1 U9274 ( .A(n8778), .B(n6912), .ZN(n7777) );
  NAND2_X1 U9275 ( .A1(n8106), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7774) );
  NAND2_X1 U9276 ( .A1(n6750), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7773) );
  INV_X1 U9277 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8013) );
  INV_X1 U9278 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8347) );
  OAI21_X1 U9279 ( .B1(n7767), .B2(n8013), .A(n8347), .ZN(n7770) );
  INV_X1 U9280 ( .A(n7767), .ZN(n7769) );
  AND2_X1 U9281 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n7768) );
  NAND2_X1 U9282 ( .A1(n7769), .A2(n7768), .ZN(n7783) );
  AND2_X1 U9283 ( .A1(n7770), .A2(n7783), .ZN(n8028) );
  NAND2_X1 U9284 ( .A1(n7901), .A2(n8028), .ZN(n7772) );
  NAND2_X1 U9285 ( .A1(n8105), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7771) );
  NAND4_X1 U9286 ( .A1(n7774), .A2(n7773), .A3(n7772), .A4(n7771), .ZN(n8596)
         );
  NAND2_X1 U9287 ( .A1(n8596), .A2(n8118), .ZN(n7775) );
  XNOR2_X1 U9288 ( .A(n7777), .B(n7775), .ZN(n8026) );
  NAND2_X1 U9289 ( .A1(n8027), .A2(n8026), .ZN(n7779) );
  INV_X1 U9290 ( .A(n7775), .ZN(n7776) );
  NAND2_X1 U9291 ( .A1(n7777), .A2(n7776), .ZN(n7778) );
  NAND2_X1 U9292 ( .A1(n7779), .A2(n7778), .ZN(n8060) );
  NAND2_X1 U9293 ( .A1(n7780), .A2(n8110), .ZN(n7782) );
  AOI22_X1 U9294 ( .A1(n7795), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7794), .B2(
        n8379), .ZN(n7781) );
  XNOR2_X1 U9295 ( .A(n8771), .B(n6912), .ZN(n7791) );
  NAND2_X1 U9296 ( .A1(n8105), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7788) );
  NAND2_X1 U9297 ( .A1(n7783), .A2(n8359), .ZN(n7784) );
  AND2_X1 U9298 ( .A1(n7815), .A2(n7784), .ZN(n8590) );
  NAND2_X1 U9299 ( .A1(n7141), .A2(n8590), .ZN(n7787) );
  NAND2_X1 U9300 ( .A1(n6750), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7786) );
  NAND2_X1 U9301 ( .A1(n8106), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7785) );
  NAND4_X1 U9302 ( .A1(n7788), .A2(n7787), .A3(n7786), .A4(n7785), .ZN(n8580)
         );
  NAND2_X1 U9303 ( .A1(n8580), .A2(n8118), .ZN(n7789) );
  XNOR2_X1 U9304 ( .A(n7791), .B(n7789), .ZN(n8061) );
  INV_X1 U9305 ( .A(n7789), .ZN(n7790) );
  NAND2_X1 U9306 ( .A1(n7791), .A2(n7790), .ZN(n7792) );
  NAND2_X1 U9307 ( .A1(n7793), .A2(n8110), .ZN(n7797) );
  AOI22_X1 U9308 ( .A1(n7795), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6456), .B2(
        n7794), .ZN(n7796) );
  XNOR2_X1 U9309 ( .A(n8767), .B(n6919), .ZN(n7802) );
  NAND2_X1 U9310 ( .A1(n8105), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n7801) );
  XNOR2_X1 U9311 ( .A(n7815), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n8574) );
  NAND2_X1 U9312 ( .A1(n7901), .A2(n8574), .ZN(n7800) );
  NAND2_X1 U9313 ( .A1(n6750), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n7799) );
  NAND2_X1 U9314 ( .A1(n8106), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n7798) );
  NAND4_X1 U9315 ( .A1(n7801), .A2(n7800), .A3(n7799), .A4(n7798), .ZN(n8597)
         );
  NAND2_X1 U9316 ( .A1(n8597), .A2(n8118), .ZN(n7803) );
  NAND2_X1 U9317 ( .A1(n7802), .A2(n7803), .ZN(n7807) );
  INV_X1 U9318 ( .A(n7802), .ZN(n7805) );
  INV_X1 U9319 ( .A(n7803), .ZN(n7804) );
  NAND2_X1 U9320 ( .A1(n7805), .A2(n7804), .ZN(n7806) );
  NAND2_X1 U9321 ( .A1(n7807), .A2(n7806), .ZN(n7960) );
  NAND2_X1 U9322 ( .A1(n7808), .A2(n8110), .ZN(n7811) );
  OR2_X1 U9323 ( .A1(n8111), .A2(n7809), .ZN(n7810) );
  XNOR2_X1 U9324 ( .A(n8761), .B(n6919), .ZN(n7821) );
  NAND2_X1 U9325 ( .A1(n8105), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n7820) );
  INV_X1 U9326 ( .A(n7815), .ZN(n7813) );
  AND2_X1 U9327 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .ZN(n7812) );
  NAND2_X1 U9328 ( .A1(n7813), .A2(n7812), .ZN(n7830) );
  INV_X1 U9329 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7961) );
  INV_X1 U9330 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7814) );
  OAI21_X1 U9331 ( .B1(n7815), .B2(n7961), .A(n7814), .ZN(n7816) );
  AND2_X1 U9332 ( .A1(n7830), .A2(n7816), .ZN(n8559) );
  NAND2_X1 U9333 ( .A1(n7901), .A2(n8559), .ZN(n7819) );
  NAND2_X1 U9334 ( .A1(n6750), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n7818) );
  NAND2_X1 U9335 ( .A1(n8106), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n7817) );
  NAND4_X1 U9336 ( .A1(n7820), .A2(n7819), .A3(n7818), .A4(n7817), .ZN(n8581)
         );
  NAND2_X1 U9337 ( .A1(n8581), .A2(n8118), .ZN(n7822) );
  XNOR2_X1 U9338 ( .A(n7821), .B(n7822), .ZN(n8041) );
  INV_X1 U9339 ( .A(n7821), .ZN(n7824) );
  INV_X1 U9340 ( .A(n7822), .ZN(n7823) );
  NAND2_X1 U9341 ( .A1(n7824), .A2(n7823), .ZN(n7825) );
  NAND2_X1 U9342 ( .A1(n7826), .A2(n8110), .ZN(n7829) );
  OR2_X1 U9343 ( .A1(n8111), .A2(n7827), .ZN(n7828) );
  XNOR2_X1 U9344 ( .A(n8756), .B(n6912), .ZN(n7838) );
  NAND2_X1 U9345 ( .A1(n8106), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7835) );
  INV_X1 U9346 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7991) );
  NAND2_X1 U9347 ( .A1(n7830), .A2(n7991), .ZN(n7831) );
  AND2_X1 U9348 ( .A1(n7858), .A2(n7831), .ZN(n8544) );
  NAND2_X1 U9349 ( .A1(n7141), .A2(n8544), .ZN(n7834) );
  NAND2_X1 U9350 ( .A1(n6750), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n7833) );
  NAND2_X1 U9351 ( .A1(n8105), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7832) );
  NAND4_X1 U9352 ( .A1(n7835), .A2(n7834), .A3(n7833), .A4(n7832), .ZN(n8415)
         );
  NAND2_X1 U9353 ( .A1(n8415), .A2(n8118), .ZN(n7836) );
  XNOR2_X1 U9354 ( .A(n7838), .B(n7836), .ZN(n7990) );
  INV_X1 U9355 ( .A(n7836), .ZN(n7837) );
  NAND2_X1 U9356 ( .A1(n7839), .A2(n8110), .ZN(n7842) );
  OR2_X1 U9357 ( .A1(n8111), .A2(n7840), .ZN(n7841) );
  XOR2_X1 U9358 ( .A(n6912), .B(n8751), .Z(n7847) );
  XNOR2_X1 U9359 ( .A(n7848), .B(n7847), .ZN(n8052) );
  XNOR2_X1 U9360 ( .A(n7858), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U9361 ( .A1(n7141), .A2(n8528), .ZN(n7846) );
  NAND2_X1 U9362 ( .A1(n6750), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n7845) );
  NAND2_X1 U9363 ( .A1(n8105), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n7844) );
  NAND2_X1 U9364 ( .A1(n8106), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n7843) );
  NOR2_X1 U9365 ( .A1(n8416), .A2(n6905), .ZN(n8053) );
  NOR2_X1 U9366 ( .A1(n8052), .A2(n8053), .ZN(n8051) );
  INV_X1 U9367 ( .A(n7847), .ZN(n7850) );
  NAND2_X1 U9368 ( .A1(n7852), .A2(n8110), .ZN(n7855) );
  OR2_X1 U9369 ( .A1(n8111), .A2(n7853), .ZN(n7854) );
  XNOR2_X1 U9370 ( .A(n8745), .B(n6912), .ZN(n7864) );
  NAND2_X1 U9371 ( .A1(n8105), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n7863) );
  INV_X1 U9372 ( .A(n7858), .ZN(n7857) );
  AND2_X1 U9373 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n7856) );
  NAND2_X1 U9374 ( .A1(n7857), .A2(n7856), .ZN(n7870) );
  INV_X1 U9375 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8054) );
  INV_X1 U9376 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7951) );
  OAI21_X1 U9377 ( .B1(n7858), .B2(n8054), .A(n7951), .ZN(n7859) );
  AND2_X1 U9378 ( .A1(n7870), .A2(n7859), .ZN(n8515) );
  NAND2_X1 U9379 ( .A1(n7901), .A2(n8515), .ZN(n7862) );
  NAND2_X1 U9380 ( .A1(n6750), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n7861) );
  NAND2_X1 U9381 ( .A1(n8106), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n7860) );
  NAND4_X1 U9382 ( .A1(n7863), .A2(n7862), .A3(n7861), .A4(n7860), .ZN(n8501)
         );
  NAND2_X1 U9383 ( .A1(n8501), .A2(n8118), .ZN(n7949) );
  NAND2_X1 U9384 ( .A1(n7865), .A2(n8110), .ZN(n7868) );
  OR2_X1 U9385 ( .A1(n8111), .A2(n7866), .ZN(n7867) );
  XNOR2_X1 U9386 ( .A(n8740), .B(n6912), .ZN(n7876) );
  INV_X1 U9387 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8035) );
  NAND2_X1 U9388 ( .A1(n7870), .A2(n8035), .ZN(n7871) );
  AND2_X1 U9389 ( .A1(n7899), .A2(n7871), .ZN(n8496) );
  NAND2_X1 U9390 ( .A1(n8496), .A2(n7901), .ZN(n7875) );
  NAND2_X1 U9391 ( .A1(n8105), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n7874) );
  NAND2_X1 U9392 ( .A1(n6750), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n7873) );
  NAND2_X1 U9393 ( .A1(n6463), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n7872) );
  NAND4_X1 U9394 ( .A1(n7875), .A2(n7874), .A3(n7873), .A4(n7872), .ZN(n8511)
         );
  AND2_X1 U9395 ( .A1(n8511), .A2(n8118), .ZN(n8034) );
  NAND2_X1 U9396 ( .A1(n8033), .A2(n8034), .ZN(n7879) );
  NAND2_X1 U9397 ( .A1(n7877), .A2(n7876), .ZN(n7878) );
  NAND2_X1 U9398 ( .A1(n7879), .A2(n7878), .ZN(n7890) );
  NAND2_X1 U9399 ( .A1(n7880), .A2(n8110), .ZN(n7883) );
  OR2_X1 U9400 ( .A1(n8111), .A2(n7881), .ZN(n7882) );
  NAND2_X2 U9401 ( .A1(n7883), .A2(n7882), .ZN(n8737) );
  XNOR2_X1 U9402 ( .A(n8737), .B(n6912), .ZN(n7891) );
  NAND2_X1 U9403 ( .A1(n7890), .A2(n7891), .ZN(n7889) );
  INV_X1 U9404 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n7888) );
  NAND2_X1 U9405 ( .A1(n8105), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U9406 ( .A1(n8106), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n7884) );
  AND2_X1 U9407 ( .A1(n7885), .A2(n7884), .ZN(n7887) );
  XNOR2_X1 U9408 ( .A(n7899), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U9409 ( .A1(n8488), .A2(n7141), .ZN(n7886) );
  OAI211_X1 U9410 ( .C1(n7984), .C2(n7888), .A(n7887), .B(n7886), .ZN(n8502)
         );
  NAND2_X1 U9411 ( .A1(n8502), .A2(n8118), .ZN(n7998) );
  NAND2_X1 U9412 ( .A1(n7889), .A2(n7998), .ZN(n7893) );
  INV_X1 U9413 ( .A(n7890), .ZN(n7997) );
  INV_X1 U9414 ( .A(n7891), .ZN(n7999) );
  NAND2_X1 U9415 ( .A1(n7997), .A2(n7999), .ZN(n7892) );
  NAND2_X1 U9416 ( .A1(n7894), .A2(n8110), .ZN(n7897) );
  OR2_X1 U9417 ( .A1(n8111), .A2(n7895), .ZN(n7896) );
  NAND2_X2 U9418 ( .A1(n7897), .A2(n7896), .ZN(n8732) );
  XNOR2_X1 U9419 ( .A(n8732), .B(n6919), .ZN(n7908) );
  INV_X1 U9420 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n7906) );
  INV_X1 U9421 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8001) );
  INV_X1 U9422 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8070) );
  OAI21_X1 U9423 ( .B1(n7899), .B2(n8001), .A(n8070), .ZN(n7900) );
  NAND2_X1 U9424 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .ZN(n7898) );
  AND2_X1 U9425 ( .A1(n7900), .A2(n7914), .ZN(n8476) );
  NAND2_X1 U9426 ( .A1(n8476), .A2(n7901), .ZN(n7905) );
  NAND2_X1 U9427 ( .A1(n8105), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n7903) );
  NAND2_X1 U9428 ( .A1(n6463), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7902) );
  AND2_X1 U9429 ( .A1(n7903), .A2(n7902), .ZN(n7904) );
  OAI211_X1 U9430 ( .C1(n7984), .C2(n7906), .A(n7905), .B(n7904), .ZN(n8464)
         );
  NAND2_X1 U9431 ( .A1(n8464), .A2(n8118), .ZN(n7907) );
  NOR2_X1 U9432 ( .A1(n7908), .A2(n7907), .ZN(n7909) );
  AOI21_X1 U9433 ( .B1(n7908), .B2(n7907), .A(n7909), .ZN(n8068) );
  INV_X1 U9434 ( .A(n7909), .ZN(n7910) );
  XNOR2_X1 U9435 ( .A(n8725), .B(n6919), .ZN(n7921) );
  INV_X1 U9436 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n7919) );
  INV_X1 U9437 ( .A(n7914), .ZN(n7912) );
  NAND2_X1 U9438 ( .A1(n7912), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n7926) );
  INV_X1 U9439 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7913) );
  NAND2_X1 U9440 ( .A1(n7914), .A2(n7913), .ZN(n7915) );
  NAND2_X1 U9441 ( .A1(n7926), .A2(n7915), .ZN(n8457) );
  INV_X1 U9442 ( .A(n7141), .ZN(n7980) );
  OR2_X1 U9443 ( .A1(n8457), .A2(n7980), .ZN(n7918) );
  AOI22_X1 U9444 ( .A1(n8105), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n6463), .B2(
        P2_REG0_REG_27__SCAN_IN), .ZN(n7917) );
  OAI211_X1 U9445 ( .C1(n7984), .C2(n7919), .A(n7918), .B(n7917), .ZN(n8311)
         );
  NAND2_X1 U9446 ( .A1(n8311), .A2(n8118), .ZN(n7920) );
  NOR2_X1 U9447 ( .A1(n7921), .A2(n7920), .ZN(n7966) );
  AOI21_X1 U9448 ( .B1(n7921), .B2(n7920), .A(n7966), .ZN(n7922) );
  OAI211_X1 U9449 ( .C1(n7923), .C2(n7922), .A(n7967), .B(n9709), .ZN(n7938)
         );
  NOR2_X1 U9450 ( .A1(n8080), .A2(n8457), .ZN(n7936) );
  INV_X1 U9451 ( .A(n7926), .ZN(n7924) );
  NAND2_X1 U9452 ( .A1(n7924), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8431) );
  INV_X1 U9453 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7925) );
  NAND2_X1 U9454 ( .A1(n7926), .A2(n7925), .ZN(n7927) );
  NAND2_X1 U9455 ( .A1(n8431), .A2(n7927), .ZN(n7979) );
  OR2_X1 U9456 ( .A1(n7979), .A2(n7980), .ZN(n7934) );
  INV_X1 U9457 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U9458 ( .A1(n6750), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7929) );
  NAND2_X1 U9459 ( .A1(n6463), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7928) );
  OAI211_X1 U9460 ( .C1(n7931), .C2(n7930), .A(n7929), .B(n7928), .ZN(n7932)
         );
  INV_X1 U9461 ( .A(n7932), .ZN(n7933) );
  NAND2_X1 U9462 ( .A1(n7934), .A2(n7933), .ZN(n8463) );
  INV_X1 U9463 ( .A(n8464), .ZN(n8274) );
  OAI22_X1 U9464 ( .A1(n8420), .A2(n9703), .B1(n9704), .B2(n8274), .ZN(n7935)
         );
  AOI211_X1 U9465 ( .C1(P2_REG3_REG_27__SCAN_IN), .C2(P2_U3152), .A(n7936), 
        .B(n7935), .ZN(n7937) );
  OAI211_X1 U9466 ( .C1(n8460), .C2(n9701), .A(n7938), .B(n7937), .ZN(P2_U3216) );
  AOI21_X1 U9467 ( .B1(n7940), .B2(n7939), .A(n4333), .ZN(n7945) );
  OAI22_X1 U9468 ( .A1(n8660), .A2(n9703), .B1(n9704), .B2(n8693), .ZN(n7941)
         );
  AOI211_X1 U9469 ( .C1(n8073), .C2(n8654), .A(n7942), .B(n7941), .ZN(n7944)
         );
  NAND2_X1 U9470 ( .A1(n8083), .A2(n8791), .ZN(n7943) );
  OAI211_X1 U9471 ( .C1(n7945), .C2(n8085), .A(n7944), .B(n7943), .ZN(P2_U3217) );
  INV_X1 U9472 ( .A(n7946), .ZN(n7948) );
  NAND2_X1 U9473 ( .A1(n7948), .A2(n7947), .ZN(n7950) );
  XNOR2_X1 U9474 ( .A(n7950), .B(n7949), .ZN(n7956) );
  INV_X1 U9475 ( .A(n8515), .ZN(n7952) );
  OAI22_X1 U9476 ( .A1(n8080), .A2(n7952), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7951), .ZN(n7954) );
  INV_X1 U9477 ( .A(n8511), .ZN(n8256) );
  OAI22_X1 U9478 ( .A1(n8256), .A2(n9703), .B1(n9704), .B2(n8416), .ZN(n7953)
         );
  AOI211_X1 U9479 ( .C1(n8745), .C2(n8083), .A(n7954), .B(n7953), .ZN(n7955)
         );
  OAI21_X1 U9480 ( .B1(n7956), .B2(n8085), .A(n7955), .ZN(P2_U3218) );
  INV_X1 U9481 ( .A(n7958), .ZN(n7959) );
  AOI21_X1 U9482 ( .B1(n7957), .B2(n7960), .A(n7959), .ZN(n7965) );
  NOR2_X1 U9483 ( .A1(n7961), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8390) );
  INV_X1 U9484 ( .A(n8581), .ZN(n8092) );
  OAI22_X1 U9485 ( .A1(n8609), .A2(n9704), .B1(n9703), .B2(n8092), .ZN(n7962)
         );
  AOI211_X1 U9486 ( .C1(n8073), .C2(n8574), .A(n8390), .B(n7962), .ZN(n7964)
         );
  NAND2_X1 U9487 ( .A1(n8767), .A2(n8083), .ZN(n7963) );
  OAI211_X1 U9488 ( .C1(n7965), .C2(n8085), .A(n7964), .B(n7963), .ZN(P2_U3221) );
  NAND2_X1 U9489 ( .A1(n7968), .A2(n8110), .ZN(n7971) );
  OR2_X1 U9490 ( .A1(n8111), .A2(n7969), .ZN(n7970) );
  NAND2_X1 U9491 ( .A1(n8463), .A2(n8118), .ZN(n7972) );
  XNOR2_X1 U9492 ( .A(n7972), .B(n6912), .ZN(n7975) );
  NOR3_X1 U9493 ( .A1(n8448), .A2(n7975), .A3(n8083), .ZN(n7973) );
  AOI21_X1 U9494 ( .B1(n8448), .B2(n7975), .A(n7973), .ZN(n7978) );
  NAND3_X1 U9495 ( .A1(n8720), .A2(n9701), .A3(n7975), .ZN(n7974) );
  OAI21_X1 U9496 ( .B1(n8720), .B2(n7975), .A(n7974), .ZN(n7976) );
  OAI21_X1 U9497 ( .B1(n8448), .B2(n9701), .A(n8085), .ZN(n7977) );
  INV_X1 U9498 ( .A(n7979), .ZN(n8446) );
  AOI22_X1 U9499 ( .A1(n8073), .A2(n8446), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n7988) );
  INV_X1 U9500 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7983) );
  OR2_X1 U9501 ( .A1(n8431), .A2(n7980), .ZN(n7982) );
  AOI22_X1 U9502 ( .A1(n8105), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8106), .B2(
        P2_REG0_REG_29__SCAN_IN), .ZN(n7981) );
  OAI211_X1 U9503 ( .C1(n7984), .C2(n7983), .A(n7982), .B(n7981), .ZN(n8310)
         );
  AOI22_X1 U9504 ( .A1(n7986), .A2(n8310), .B1(n7985), .B2(n8311), .ZN(n7987)
         );
  XNOR2_X1 U9505 ( .A(n7989), .B(n7990), .ZN(n7996) );
  INV_X1 U9506 ( .A(n8544), .ZN(n7992) );
  OAI22_X1 U9507 ( .A1(n8080), .A2(n7992), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7991), .ZN(n7994) );
  OAI22_X1 U9508 ( .A1(n8416), .A2(n9703), .B1(n9704), .B2(n8092), .ZN(n7993)
         );
  AOI211_X1 U9509 ( .C1(n8756), .C2(n8083), .A(n7994), .B(n7993), .ZN(n7995)
         );
  OAI21_X1 U9510 ( .B1(n7996), .B2(n8085), .A(n7995), .ZN(P2_U3225) );
  XNOR2_X1 U9511 ( .A(n7999), .B(n7998), .ZN(n8000) );
  XNOR2_X1 U9512 ( .A(n7997), .B(n8000), .ZN(n8005) );
  AOI22_X1 U9513 ( .A1(n8464), .A2(n9764), .B1(n9762), .B2(n8511), .ZN(n8485)
         );
  OAI22_X1 U9514 ( .A1(n8071), .A2(n8485), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8001), .ZN(n8003) );
  INV_X1 U9515 ( .A(n8737), .ZN(n8491) );
  NOR2_X1 U9516 ( .A1(n8491), .A2(n9701), .ZN(n8002) );
  AOI211_X1 U9517 ( .C1(n8073), .C2(n8488), .A(n8003), .B(n8002), .ZN(n8004)
         );
  OAI21_X1 U9518 ( .B1(n8005), .B2(n8085), .A(n8004), .ZN(P2_U3227) );
  INV_X1 U9519 ( .A(n8781), .ZN(n8630) );
  XNOR2_X1 U9520 ( .A(n8006), .B(n8007), .ZN(n8077) );
  OAI22_X1 U9521 ( .A1(n8077), .A2(n8076), .B1(n8007), .B2(n8006), .ZN(n8011)
         );
  NAND2_X1 U9522 ( .A1(n8009), .A2(n8008), .ZN(n8010) );
  XNOR2_X1 U9523 ( .A(n8011), .B(n8010), .ZN(n8012) );
  NAND2_X1 U9524 ( .A1(n8012), .A2(n9709), .ZN(n8016) );
  NOR2_X1 U9525 ( .A1(n8013), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8328) );
  INV_X1 U9526 ( .A(n8596), .ZN(n8619) );
  OAI22_X1 U9527 ( .A1(n8660), .A2(n9704), .B1(n9703), .B2(n8619), .ZN(n8014)
         );
  AOI211_X1 U9528 ( .C1(n8073), .C2(n8628), .A(n8328), .B(n8014), .ZN(n8015)
         );
  OAI211_X1 U9529 ( .C1(n8630), .C2(n9701), .A(n8016), .B(n8015), .ZN(P2_U3228) );
  AOI22_X1 U9530 ( .A1(n8073), .A2(n8018), .B1(n8083), .B2(n8017), .ZN(n8025)
         );
  INV_X1 U9531 ( .A(n8071), .ZN(n8045) );
  AOI22_X1 U9532 ( .A1(n8045), .A2(n8019), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n8024) );
  OAI211_X1 U9533 ( .C1(n8022), .C2(n8021), .A(n8020), .B(n9709), .ZN(n8023)
         );
  NAND3_X1 U9534 ( .A1(n8025), .A2(n8024), .A3(n8023), .ZN(P2_U3229) );
  XNOR2_X1 U9535 ( .A(n8027), .B(n8026), .ZN(n8032) );
  OAI22_X1 U9536 ( .A1(n8644), .A2(n9704), .B1(n9703), .B2(n8609), .ZN(n8030)
         );
  INV_X1 U9537 ( .A(n8028), .ZN(n8612) );
  OAI22_X1 U9538 ( .A1(n8080), .A2(n8612), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8347), .ZN(n8029) );
  AOI211_X1 U9539 ( .C1(n8778), .C2(n8083), .A(n8030), .B(n8029), .ZN(n8031)
         );
  OAI21_X1 U9540 ( .B1(n8032), .B2(n8085), .A(n8031), .ZN(P2_U3230) );
  XNOR2_X1 U9541 ( .A(n8033), .B(n8034), .ZN(n8040) );
  INV_X1 U9542 ( .A(n8496), .ZN(n8036) );
  OAI22_X1 U9543 ( .A1(n8080), .A2(n8036), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8035), .ZN(n8038) );
  INV_X1 U9544 ( .A(n8502), .ZN(n8094) );
  OAI22_X1 U9545 ( .A1(n8537), .A2(n9704), .B1(n9703), .B2(n8094), .ZN(n8037)
         );
  AOI211_X1 U9546 ( .C1(n8740), .C2(n8083), .A(n8038), .B(n8037), .ZN(n8039)
         );
  OAI21_X1 U9547 ( .B1(n8040), .B2(n8085), .A(n8039), .ZN(P2_U3231) );
  XNOR2_X1 U9548 ( .A(n8042), .B(n8041), .ZN(n8050) );
  INV_X1 U9549 ( .A(n8559), .ZN(n8047) );
  NAND2_X1 U9550 ( .A1(n8597), .A2(n9762), .ZN(n8044) );
  NAND2_X1 U9551 ( .A1(n8415), .A2(n9764), .ZN(n8043) );
  NAND2_X1 U9552 ( .A1(n8044), .A2(n8043), .ZN(n8567) );
  AOI22_X1 U9553 ( .A1(n8045), .A2(n8567), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8046) );
  OAI21_X1 U9554 ( .B1(n8080), .B2(n8047), .A(n8046), .ZN(n8048) );
  AOI21_X1 U9555 ( .B1(n8761), .B2(n8083), .A(n8048), .ZN(n8049) );
  OAI21_X1 U9556 ( .B1(n8050), .B2(n8085), .A(n8049), .ZN(P2_U3235) );
  AOI21_X1 U9557 ( .B1(n8053), .B2(n8052), .A(n8051), .ZN(n8059) );
  INV_X1 U9558 ( .A(n8528), .ZN(n8055) );
  OAI22_X1 U9559 ( .A1(n8080), .A2(n8055), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8054), .ZN(n8057) );
  INV_X1 U9560 ( .A(n8415), .ZN(n8536) );
  OAI22_X1 U9561 ( .A1(n8537), .A2(n9703), .B1(n9704), .B2(n8536), .ZN(n8056)
         );
  AOI211_X1 U9562 ( .C1(n8751), .C2(n8083), .A(n8057), .B(n8056), .ZN(n8058)
         );
  OAI21_X1 U9563 ( .B1(n8059), .B2(n8085), .A(n8058), .ZN(P2_U3237) );
  XNOR2_X1 U9564 ( .A(n8060), .B(n8061), .ZN(n8066) );
  INV_X1 U9565 ( .A(n8597), .ZN(n8413) );
  OAI22_X1 U9566 ( .A1(n8619), .A2(n9704), .B1(n9703), .B2(n8413), .ZN(n8064)
         );
  INV_X1 U9567 ( .A(n8590), .ZN(n8062) );
  OAI22_X1 U9568 ( .A1(n8080), .A2(n8062), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8359), .ZN(n8063) );
  AOI211_X1 U9569 ( .C1(n8771), .C2(n8083), .A(n8064), .B(n8063), .ZN(n8065)
         );
  OAI21_X1 U9570 ( .B1(n8066), .B2(n8085), .A(n8065), .ZN(P2_U3240) );
  INV_X1 U9571 ( .A(n8732), .ZN(n8479) );
  OAI211_X1 U9572 ( .C1(n8069), .C2(n8068), .A(n8067), .B(n9709), .ZN(n8075)
         );
  AOI22_X1 U9573 ( .A1(n8311), .A2(n9764), .B1(n9762), .B2(n8502), .ZN(n8472)
         );
  OAI22_X1 U9574 ( .A1(n8071), .A2(n8472), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8070), .ZN(n8072) );
  AOI21_X1 U9575 ( .B1(n8073), .B2(n8476), .A(n8072), .ZN(n8074) );
  OAI211_X1 U9576 ( .C1(n8479), .C2(n9701), .A(n8075), .B(n8074), .ZN(P2_U3242) );
  XNOR2_X1 U9577 ( .A(n8077), .B(n8076), .ZN(n8086) );
  OAI22_X1 U9578 ( .A1(n8644), .A2(n9703), .B1(n9704), .B2(n8668), .ZN(n8082)
         );
  INV_X1 U9579 ( .A(n8638), .ZN(n8079) );
  OAI22_X1 U9580 ( .A1(n8080), .A2(n8079), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8078), .ZN(n8081) );
  AOI211_X1 U9581 ( .C1(n8786), .C2(n8083), .A(n8082), .B(n8081), .ZN(n8084)
         );
  OAI21_X1 U9582 ( .B1(n8086), .B2(n8085), .A(n8084), .ZN(P2_U3243) );
  INV_X1 U9583 ( .A(n8204), .ZN(n8087) );
  AOI21_X2 U9584 ( .B1(n8088), .B2(n8208), .A(n8087), .ZN(n8687) );
  NAND2_X1 U9585 ( .A1(n8697), .A2(n8669), .ZN(n8209) );
  INV_X1 U9586 ( .A(n8209), .ZN(n8203) );
  OR2_X1 U9587 ( .A1(n8697), .A2(n8669), .ZN(n8210) );
  OR2_X1 U9588 ( .A1(n8797), .A2(n8693), .ZN(n8216) );
  NAND2_X1 U9589 ( .A1(n8797), .A2(n8693), .ZN(n8215) );
  INV_X1 U9590 ( .A(n8670), .ZN(n8667) );
  OAI21_X1 U9591 ( .B1(n8666), .B2(n8667), .A(n8215), .ZN(n8658) );
  NAND2_X1 U9592 ( .A1(n8791), .A2(n8668), .ZN(n8219) );
  INV_X1 U9593 ( .A(n8653), .ZN(n8659) );
  INV_X1 U9594 ( .A(n8218), .ZN(n8089) );
  XNOR2_X1 U9595 ( .A(n8786), .B(n8660), .ZN(n8643) );
  INV_X1 U9596 ( .A(n8786), .ZN(n8640) );
  OR2_X1 U9597 ( .A1(n8781), .A2(n8644), .ZN(n8225) );
  NAND2_X1 U9598 ( .A1(n8781), .A2(n8644), .ZN(n8224) );
  OR2_X1 U9599 ( .A1(n8778), .A2(n8619), .ZN(n8091) );
  NAND2_X1 U9600 ( .A1(n8778), .A2(n8619), .ZN(n8229) );
  NAND2_X1 U9601 ( .A1(n8091), .A2(n8229), .ZN(n8603) );
  INV_X1 U9602 ( .A(n8603), .ZN(n8606) );
  INV_X1 U9603 ( .A(n8091), .ZN(n8227) );
  NOR2_X1 U9604 ( .A1(n8771), .A2(n8609), .ZN(n8233) );
  AND2_X1 U9605 ( .A1(n8771), .A2(n8609), .ZN(n8235) );
  NOR2_X1 U9606 ( .A1(n8233), .A2(n8235), .ZN(n8594) );
  NAND2_X1 U9607 ( .A1(n8595), .A2(n8594), .ZN(n8593) );
  INV_X1 U9608 ( .A(n8235), .ZN(n8243) );
  NAND2_X1 U9609 ( .A1(n8593), .A2(n8243), .ZN(n8578) );
  OR2_X1 U9610 ( .A1(n8767), .A2(n8413), .ZN(n8241) );
  NAND2_X1 U9611 ( .A1(n8767), .A2(n8413), .ZN(n8564) );
  NAND2_X1 U9612 ( .A1(n8761), .A2(n8092), .ZN(n8245) );
  NAND2_X1 U9613 ( .A1(n8247), .A2(n8245), .ZN(n8554) );
  INV_X1 U9614 ( .A(n8554), .ZN(n8563) );
  OR2_X1 U9615 ( .A1(n8756), .A2(n8536), .ZN(n8246) );
  NAND2_X1 U9616 ( .A1(n8756), .A2(n8536), .ZN(n8533) );
  NAND2_X1 U9617 ( .A1(n8751), .A2(n8416), .ZN(n8263) );
  NAND2_X1 U9618 ( .A1(n8238), .A2(n8263), .ZN(n8417) );
  INV_X1 U9619 ( .A(n8417), .ZN(n8532) );
  OR2_X1 U9620 ( .A1(n8745), .A2(n8537), .ZN(n8266) );
  NAND2_X1 U9621 ( .A1(n8745), .A2(n8537), .ZN(n8253) );
  NAND2_X1 U9622 ( .A1(n8266), .A2(n8253), .ZN(n8519) );
  INV_X1 U9623 ( .A(n8238), .ZN(n8508) );
  NOR2_X1 U9624 ( .A1(n8519), .A2(n8508), .ZN(n8255) );
  NAND2_X1 U9625 ( .A1(n8507), .A2(n8255), .ZN(n8509) );
  NAND2_X1 U9626 ( .A1(n8740), .A2(n8511), .ZN(n8093) );
  NAND2_X1 U9627 ( .A1(n8418), .A2(n8093), .ZN(n8500) );
  INV_X1 U9628 ( .A(n8500), .ZN(n8270) );
  NAND2_X1 U9629 ( .A1(n8737), .A2(n8094), .ZN(n8260) );
  NAND2_X1 U9630 ( .A1(n8732), .A2(n8274), .ZN(n8095) );
  INV_X1 U9631 ( .A(n8311), .ZN(n8440) );
  NOR2_X1 U9632 ( .A1(n8725), .A2(n8440), .ZN(n8281) );
  NAND2_X1 U9633 ( .A1(n8720), .A2(n8420), .ZN(n8096) );
  NOR2_X1 U9634 ( .A1(n8439), .A2(n8450), .ZN(n8438) );
  NAND2_X1 U9635 ( .A1(n8097), .A2(n8110), .ZN(n8100) );
  OR2_X1 U9636 ( .A1(n8111), .A2(n8098), .ZN(n8099) );
  NAND2_X1 U9637 ( .A1(n8100), .A2(n8099), .ZN(n8391) );
  INV_X1 U9638 ( .A(n8310), .ZN(n8441) );
  OR2_X1 U9639 ( .A1(n8391), .A2(n8441), .ZN(n8286) );
  NAND2_X1 U9640 ( .A1(n8391), .A2(n8441), .ZN(n8285) );
  NAND2_X1 U9641 ( .A1(n8101), .A2(n8110), .ZN(n8104) );
  OR2_X1 U9642 ( .A1(n8111), .A2(n8102), .ZN(n8103) );
  NAND2_X1 U9643 ( .A1(n8105), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U9644 ( .A1(n6750), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8108) );
  NAND2_X1 U9645 ( .A1(n8106), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8107) );
  NAND3_X1 U9646 ( .A1(n8109), .A2(n8108), .A3(n8107), .ZN(n8426) );
  INV_X1 U9647 ( .A(n8426), .ZN(n8114) );
  OR2_X1 U9648 ( .A1(n8396), .A2(n8114), .ZN(n8289) );
  NAND2_X1 U9649 ( .A1(n9534), .A2(n8110), .ZN(n8113) );
  OR2_X1 U9650 ( .A1(n8111), .A2(n8822), .ZN(n8112) );
  OR2_X1 U9651 ( .A1(n8705), .A2(n8115), .ZN(n8296) );
  NAND2_X1 U9652 ( .A1(n8396), .A2(n8114), .ZN(n8288) );
  NAND2_X1 U9653 ( .A1(n8296), .A2(n8288), .ZN(n8119) );
  XNOR2_X1 U9654 ( .A(n8116), .B(n8389), .ZN(n8303) );
  NAND2_X1 U9655 ( .A1(n8118), .A2(n8117), .ZN(n8302) );
  INV_X1 U9656 ( .A(n8119), .ZN(n8291) );
  AND2_X1 U9657 ( .A1(n4298), .A2(n8289), .ZN(n8290) );
  INV_X1 U9658 ( .A(n8547), .ZN(n8138) );
  NAND2_X1 U9659 ( .A1(n8225), .A2(n8224), .ZN(n8620) );
  NOR2_X1 U9660 ( .A1(n8120), .A2(n6449), .ZN(n8124) );
  INV_X1 U9661 ( .A(n8121), .ZN(n8123) );
  INV_X1 U9662 ( .A(n6447), .ZN(n8122) );
  NAND4_X1 U9663 ( .A1(n8124), .A2(n8123), .A3(n8122), .A4(n8165), .ZN(n8129)
         );
  INV_X1 U9664 ( .A(n8125), .ZN(n8127) );
  NAND2_X1 U9665 ( .A1(n8127), .A2(n8126), .ZN(n8128) );
  NOR2_X1 U9666 ( .A1(n8129), .A2(n8128), .ZN(n8131) );
  NAND4_X1 U9667 ( .A1(n8131), .A2(n8181), .A3(n9737), .A4(n8130), .ZN(n8133)
         );
  NOR4_X1 U9668 ( .A1(n8133), .A2(n9758), .A3(n7337), .A4(n8132), .ZN(n8134)
         );
  NAND4_X1 U9669 ( .A1(n8653), .A2(n8134), .A3(n8670), .A4(n8688), .ZN(n8135)
         );
  NOR4_X1 U9670 ( .A1(n8603), .A2(n8620), .A3(n8643), .A4(n8135), .ZN(n8136)
         );
  NAND4_X1 U9671 ( .A1(n8563), .A2(n8579), .A3(n8594), .A4(n8136), .ZN(n8137)
         );
  NOR4_X1 U9672 ( .A1(n8519), .A2(n8417), .A3(n8138), .A4(n8137), .ZN(n8139)
         );
  NAND3_X1 U9673 ( .A1(n8483), .A2(n8139), .A3(n8500), .ZN(n8140) );
  NOR4_X1 U9674 ( .A1(n8450), .A2(n8461), .A3(n8471), .A4(n8140), .ZN(n8141)
         );
  NAND4_X1 U9675 ( .A1(n8291), .A2(n8290), .A3(n8421), .A4(n8141), .ZN(n8142)
         );
  XNOR2_X1 U9676 ( .A(n8142), .B(n8389), .ZN(n8143) );
  INV_X1 U9677 ( .A(n6449), .ZN(n8297) );
  OAI22_X1 U9678 ( .A1(n8143), .A2(n6421), .B1(n8297), .B2(n6730), .ZN(n8301)
         );
  INV_X1 U9679 ( .A(n6730), .ZN(n8144) );
  NOR2_X1 U9680 ( .A1(n8144), .A2(n9822), .ZN(n8300) );
  INV_X1 U9681 ( .A(n8295), .ZN(n8280) );
  AOI21_X1 U9682 ( .B1(n8440), .B2(n8725), .A(n8450), .ZN(n8277) );
  AND2_X1 U9683 ( .A1(n8155), .A2(n8154), .ZN(n8146) );
  MUX2_X1 U9684 ( .A(n8146), .B(n8145), .S(n8295), .Z(n8166) );
  NAND2_X1 U9685 ( .A1(n8147), .A2(n8317), .ZN(n8148) );
  NAND2_X1 U9686 ( .A1(n8149), .A2(n8148), .ZN(n8152) );
  NAND2_X1 U9687 ( .A1(n9844), .A2(n8314), .ZN(n8176) );
  NAND2_X1 U9688 ( .A1(n8150), .A2(n8176), .ZN(n8151) );
  AOI21_X1 U9689 ( .B1(n8166), .B2(n8152), .A(n8151), .ZN(n8177) );
  NAND2_X1 U9690 ( .A1(n8154), .A2(n8153), .ZN(n8159) );
  INV_X1 U9691 ( .A(n8155), .ZN(n8157) );
  OR2_X1 U9692 ( .A1(n8157), .A2(n8156), .ZN(n8158) );
  AOI21_X1 U9693 ( .B1(n8166), .B2(n8159), .A(n8158), .ZN(n8168) );
  NAND2_X1 U9694 ( .A1(n8160), .A2(n6453), .ZN(n8169) );
  AND2_X1 U9695 ( .A1(n8169), .A2(n6421), .ZN(n8161) );
  OAI211_X1 U9696 ( .C1(n8162), .C2(n8161), .A(n8173), .B(n8170), .ZN(n8163)
         );
  NAND3_X1 U9697 ( .A1(n8163), .A2(n8171), .A3(n8295), .ZN(n8164) );
  NAND3_X1 U9698 ( .A1(n8166), .A2(n8165), .A3(n8164), .ZN(n8167) );
  NAND2_X1 U9699 ( .A1(n8170), .A2(n8169), .ZN(n8172) );
  NAND3_X1 U9700 ( .A1(n8172), .A2(n8171), .A3(n6452), .ZN(n8174) );
  NAND3_X1 U9701 ( .A1(n8174), .A2(n8280), .A3(n8173), .ZN(n8175) );
  NAND3_X1 U9702 ( .A1(n8179), .A2(n8280), .A3(n8178), .ZN(n8180) );
  NAND3_X1 U9703 ( .A1(n8196), .A2(n9749), .A3(n8182), .ZN(n8184) );
  NAND2_X1 U9704 ( .A1(n8184), .A2(n8183), .ZN(n8188) );
  OAI21_X1 U9705 ( .B1(n8186), .B2(n8185), .A(n8190), .ZN(n8187) );
  NAND2_X1 U9706 ( .A1(n9737), .A2(n8190), .ZN(n8193) );
  NAND2_X1 U9707 ( .A1(n8191), .A2(n8199), .ZN(n8192) );
  MUX2_X1 U9708 ( .A(n8193), .B(n8192), .S(n8295), .Z(n8202) );
  INV_X1 U9709 ( .A(n8202), .ZN(n8195) );
  NAND4_X1 U9710 ( .A1(n8196), .A2(n8195), .A3(n9749), .A4(n8194), .ZN(n8198)
         );
  NAND3_X1 U9711 ( .A1(n8198), .A2(n8204), .A3(n8197), .ZN(n8201) );
  NAND2_X1 U9712 ( .A1(n8208), .A2(n8199), .ZN(n8200) );
  INV_X1 U9713 ( .A(n8210), .ZN(n8205) );
  NOR2_X1 U9714 ( .A1(n8206), .A2(n8205), .ZN(n8214) );
  INV_X1 U9715 ( .A(n8207), .ZN(n8212) );
  NAND2_X1 U9716 ( .A1(n8209), .A2(n8208), .ZN(n8211) );
  OAI21_X1 U9717 ( .B1(n8212), .B2(n8211), .A(n8210), .ZN(n8213) );
  MUX2_X1 U9718 ( .A(n8216), .B(n8215), .S(n8295), .Z(n8217) );
  MUX2_X1 U9719 ( .A(n8219), .B(n8218), .S(n8295), .Z(n8220) );
  NAND2_X1 U9720 ( .A1(n8409), .A2(n8280), .ZN(n8222) );
  NAND2_X1 U9721 ( .A1(n8660), .A2(n8295), .ZN(n8221) );
  MUX2_X1 U9722 ( .A(n8222), .B(n8221), .S(n8786), .Z(n8223) );
  MUX2_X1 U9723 ( .A(n8225), .B(n8224), .S(n8295), .Z(n8226) );
  NAND2_X1 U9724 ( .A1(n8606), .A2(n8226), .ZN(n8231) );
  NOR2_X1 U9725 ( .A1(n8233), .A2(n8227), .ZN(n8228) );
  MUX2_X1 U9726 ( .A(n8229), .B(n8228), .S(n8295), .Z(n8230) );
  OAI21_X1 U9727 ( .B1(n8232), .B2(n8231), .A(n8230), .ZN(n8244) );
  INV_X1 U9728 ( .A(n8233), .ZN(n8234) );
  OAI211_X1 U9729 ( .C1(n8244), .C2(n8235), .A(n8241), .B(n8234), .ZN(n8237)
         );
  INV_X1 U9730 ( .A(n8247), .ZN(n8236) );
  AOI21_X1 U9731 ( .B1(n8237), .B2(n8564), .A(n8236), .ZN(n8240) );
  NAND2_X1 U9732 ( .A1(n8533), .A2(n8245), .ZN(n8239) );
  OAI211_X1 U9733 ( .C1(n8240), .C2(n8239), .A(n8238), .B(n8246), .ZN(n8252)
         );
  INV_X1 U9734 ( .A(n8241), .ZN(n8242) );
  AOI21_X1 U9735 ( .B1(n8244), .B2(n8243), .A(n8242), .ZN(n8249) );
  NAND2_X1 U9736 ( .A1(n8245), .A2(n8564), .ZN(n8248) );
  OAI211_X1 U9737 ( .C1(n8249), .C2(n8248), .A(n8247), .B(n8246), .ZN(n8250)
         );
  NAND3_X1 U9738 ( .A1(n8250), .A2(n8263), .A3(n8533), .ZN(n8251) );
  MUX2_X1 U9739 ( .A(n8252), .B(n8251), .S(n8295), .Z(n8265) );
  INV_X1 U9740 ( .A(n8253), .ZN(n8254) );
  AOI21_X1 U9741 ( .B1(n8265), .B2(n8255), .A(n8254), .ZN(n8261) );
  NAND2_X1 U9742 ( .A1(n8511), .A2(n8295), .ZN(n8258) );
  NAND2_X1 U9743 ( .A1(n8256), .A2(n8280), .ZN(n8257) );
  MUX2_X1 U9744 ( .A(n8258), .B(n8257), .S(n8740), .Z(n8259) );
  NAND2_X1 U9745 ( .A1(n8483), .A2(n8259), .ZN(n8268) );
  INV_X1 U9746 ( .A(n8471), .ZN(n8469) );
  OAI211_X1 U9747 ( .C1(n8261), .C2(n8268), .A(n8469), .B(n8260), .ZN(n8262)
         );
  INV_X1 U9748 ( .A(n8519), .ZN(n8264) );
  NAND3_X1 U9749 ( .A1(n8265), .A2(n8264), .A3(n8263), .ZN(n8267) );
  AOI21_X1 U9750 ( .B1(n8267), .B2(n8266), .A(n8295), .ZN(n8271) );
  INV_X1 U9751 ( .A(n8268), .ZN(n8269) );
  AOI21_X1 U9752 ( .B1(n8273), .B2(n8272), .A(n8295), .ZN(n8276) );
  NAND3_X1 U9753 ( .A1(n8732), .A2(n8274), .A3(n8280), .ZN(n8275) );
  NAND2_X1 U9754 ( .A1(n8278), .A2(n8279), .ZN(n8284) );
  INV_X1 U9755 ( .A(n8279), .ZN(n8423) );
  OAI21_X1 U9756 ( .B1(n8423), .B2(n8281), .A(n8280), .ZN(n8283) );
  NOR3_X1 U9757 ( .A1(n8448), .A2(n8463), .A3(n8295), .ZN(n8282) );
  INV_X1 U9758 ( .A(n8421), .ZN(n8422) );
  AOI211_X1 U9759 ( .C1(n8284), .C2(n8283), .A(n8282), .B(n8422), .ZN(n8294)
         );
  MUX2_X1 U9760 ( .A(n8286), .B(n8285), .S(n8295), .Z(n8287) );
  NAND3_X1 U9761 ( .A1(n8289), .A2(n8288), .A3(n8287), .ZN(n8293) );
  MUX2_X1 U9762 ( .A(n8291), .B(n8290), .S(n8295), .Z(n8292) );
  OAI21_X1 U9763 ( .B1(n8294), .B2(n8293), .A(n8292), .ZN(n8299) );
  MUX2_X1 U9764 ( .A(n4298), .B(n8296), .S(n8295), .Z(n8298) );
  INV_X1 U9765 ( .A(n8828), .ZN(n8392) );
  NAND4_X1 U9766 ( .A1(n8305), .A2(n8392), .A3(n8304), .A4(n9762), .ZN(n8306)
         );
  OAI211_X1 U9767 ( .C1(n8307), .C2(n8309), .A(n8306), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8308) );
  MUX2_X1 U9768 ( .A(n8426), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8319), .Z(
        P2_U3582) );
  MUX2_X1 U9769 ( .A(n8310), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8319), .Z(
        P2_U3581) );
  MUX2_X1 U9770 ( .A(n8463), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8319), .Z(
        P2_U3580) );
  MUX2_X1 U9771 ( .A(n8311), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8319), .Z(
        P2_U3579) );
  MUX2_X1 U9772 ( .A(n8464), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8319), .Z(
        P2_U3578) );
  MUX2_X1 U9773 ( .A(n8502), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8319), .Z(
        P2_U3577) );
  MUX2_X1 U9774 ( .A(n8511), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8319), .Z(
        P2_U3576) );
  MUX2_X1 U9775 ( .A(n8501), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8319), .Z(
        P2_U3575) );
  INV_X1 U9776 ( .A(n8416), .ZN(n8549) );
  MUX2_X1 U9777 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8549), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9778 ( .A(n8415), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8319), .Z(
        P2_U3573) );
  MUX2_X1 U9779 ( .A(n8581), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8319), .Z(
        P2_U3572) );
  MUX2_X1 U9780 ( .A(n8597), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8319), .Z(
        P2_U3571) );
  MUX2_X1 U9781 ( .A(n8580), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8319), .Z(
        P2_U3570) );
  MUX2_X1 U9782 ( .A(n8596), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8319), .Z(
        P2_U3569) );
  MUX2_X1 U9783 ( .A(n8411), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8319), .Z(
        P2_U3568) );
  MUX2_X1 U9784 ( .A(n8409), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8319), .Z(
        P2_U3567) );
  MUX2_X1 U9785 ( .A(n8407), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8319), .Z(
        P2_U3566) );
  MUX2_X1 U9786 ( .A(n8405), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8319), .Z(
        P2_U3565) );
  MUX2_X1 U9787 ( .A(n8403), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8319), .Z(
        P2_U3564) );
  MUX2_X1 U9788 ( .A(n9735), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8319), .Z(
        P2_U3563) );
  MUX2_X1 U9789 ( .A(n8312), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8319), .Z(
        P2_U3562) );
  MUX2_X1 U9790 ( .A(n9765), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8319), .Z(
        P2_U3561) );
  MUX2_X1 U9791 ( .A(n8313), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8319), .Z(
        P2_U3560) );
  MUX2_X1 U9792 ( .A(n9763), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8319), .Z(
        P2_U3559) );
  MUX2_X1 U9793 ( .A(n8314), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8319), .Z(
        P2_U3558) );
  MUX2_X1 U9794 ( .A(n8315), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8319), .Z(
        P2_U3557) );
  MUX2_X1 U9795 ( .A(n8316), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8319), .Z(
        P2_U3556) );
  MUX2_X1 U9796 ( .A(n8317), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8319), .Z(
        P2_U3555) );
  MUX2_X1 U9797 ( .A(n8318), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8319), .Z(
        P2_U3554) );
  MUX2_X1 U9798 ( .A(n8320), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8319), .Z(
        P2_U3553) );
  NOR2_X1 U9799 ( .A1(n8322), .A2(n8321), .ZN(n8324) );
  XOR2_X1 U9800 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8349), .Z(n8325) );
  NAND2_X1 U9801 ( .A1(n8325), .A2(n8326), .ZN(n8348) );
  OAI21_X1 U9802 ( .B1(n8326), .B2(n8325), .A(n8348), .ZN(n8327) );
  NAND2_X1 U9803 ( .A1(n8327), .A2(n9713), .ZN(n8340) );
  AOI21_X1 U9804 ( .B1(n9715), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8328), .ZN(
        n8339) );
  NOR2_X1 U9805 ( .A1(n8330), .A2(n8329), .ZN(n8332) );
  NOR2_X1 U9806 ( .A1(n8332), .A2(n8331), .ZN(n8336) );
  INV_X1 U9807 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8333) );
  MUX2_X1 U9808 ( .A(n8333), .B(P2_REG2_REG_16__SCAN_IN), .S(n8349), .Z(n8334)
         );
  INV_X1 U9809 ( .A(n8334), .ZN(n8335) );
  NAND2_X1 U9810 ( .A1(n8335), .A2(n8336), .ZN(n8341) );
  OAI211_X1 U9811 ( .C1(n8336), .C2(n8335), .A(n9714), .B(n8341), .ZN(n8338)
         );
  NAND2_X1 U9812 ( .A1(n9560), .A2(n8349), .ZN(n8337) );
  NAND4_X1 U9813 ( .A1(n8340), .A2(n8339), .A3(n8338), .A4(n8337), .ZN(
        P2_U3261) );
  NAND2_X1 U9814 ( .A1(n8349), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8342) );
  NAND2_X1 U9815 ( .A1(n8342), .A2(n8341), .ZN(n8346) );
  INV_X1 U9816 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8344) );
  NAND2_X1 U9817 ( .A1(n8363), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8358) );
  INV_X1 U9818 ( .A(n8358), .ZN(n8343) );
  AOI21_X1 U9819 ( .B1(n8344), .B2(n8356), .A(n8343), .ZN(n8345) );
  NAND2_X1 U9820 ( .A1(n8345), .A2(n8346), .ZN(n8357) );
  OAI211_X1 U9821 ( .C1(n8346), .C2(n8345), .A(n9714), .B(n8357), .ZN(n8355)
         );
  NOR2_X1 U9822 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8347), .ZN(n8353) );
  OAI21_X1 U9823 ( .B1(n8349), .B2(P2_REG1_REG_16__SCAN_IN), .A(n8348), .ZN(
        n8351) );
  XNOR2_X1 U9824 ( .A(n8363), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8350) );
  NOR2_X1 U9825 ( .A1(n8350), .A2(n8351), .ZN(n8362) );
  AOI211_X1 U9826 ( .C1(n8351), .C2(n8350), .A(n8362), .B(n9718), .ZN(n8352)
         );
  AOI211_X1 U9827 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n9715), .A(n8353), .B(
        n8352), .ZN(n8354) );
  OAI211_X1 U9828 ( .C1(n9717), .C2(n8356), .A(n8355), .B(n8354), .ZN(P2_U3262) );
  NAND2_X1 U9829 ( .A1(n8358), .A2(n8357), .ZN(n8380) );
  XNOR2_X1 U9830 ( .A(n8380), .B(n8379), .ZN(n8377) );
  XOR2_X1 U9831 ( .A(P2_REG2_REG_18__SCAN_IN), .B(n8377), .Z(n8372) );
  NOR2_X1 U9832 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8359), .ZN(n8360) );
  AOI21_X1 U9833 ( .B1(n9715), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8360), .ZN(
        n8368) );
  INV_X1 U9834 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8361) );
  XNOR2_X1 U9835 ( .A(n8379), .B(n8361), .ZN(n8365) );
  NAND2_X1 U9836 ( .A1(n8365), .A2(n8364), .ZN(n8374) );
  OAI21_X1 U9837 ( .B1(n8365), .B2(n8364), .A(n8374), .ZN(n8366) );
  NAND2_X1 U9838 ( .A1(n9713), .A2(n8366), .ZN(n8367) );
  OAI211_X1 U9839 ( .C1(n9717), .C2(n8369), .A(n8368), .B(n8367), .ZN(n8370)
         );
  INV_X1 U9840 ( .A(n8370), .ZN(n8371) );
  OAI21_X1 U9841 ( .B1(n8372), .B2(n9716), .A(n8371), .ZN(P2_U3263) );
  OR2_X1 U9842 ( .A1(n8379), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8373) );
  NAND2_X1 U9843 ( .A1(n8374), .A2(n8373), .ZN(n8376) );
  INV_X1 U9844 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8375) );
  XNOR2_X1 U9845 ( .A(n8376), .B(n8375), .ZN(n8387) );
  INV_X1 U9846 ( .A(n8387), .ZN(n8386) );
  INV_X1 U9847 ( .A(n8377), .ZN(n8378) );
  NAND2_X1 U9848 ( .A1(n8378), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U9849 ( .A1(n8380), .A2(n8379), .ZN(n8381) );
  NAND2_X1 U9850 ( .A1(n8382), .A2(n8381), .ZN(n8383) );
  XNOR2_X1 U9851 ( .A(n8383), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8388) );
  NAND3_X1 U9852 ( .A1(n8388), .A2(n8392), .A3(n8384), .ZN(n8385) );
  INV_X1 U9853 ( .A(n8697), .ZN(n9888) );
  NOR2_X1 U9854 ( .A1(n4274), .A2(n8791), .ZN(n8635) );
  NAND2_X1 U9855 ( .A1(n8636), .A2(n8630), .ZN(n8625) );
  OR2_X2 U9856 ( .A1(n8625), .A2(n8778), .ZN(n8610) );
  OR2_X2 U9857 ( .A1(n8610), .A2(n8771), .ZN(n8588) );
  INV_X1 U9858 ( .A(n8761), .ZN(n8561) );
  NAND2_X1 U9859 ( .A1(n8573), .A2(n8561), .ZN(n8556) );
  OR2_X2 U9860 ( .A1(n8556), .A2(n8756), .ZN(n8527) );
  INV_X1 U9861 ( .A(n8740), .ZN(n8498) );
  OR2_X2 U9862 ( .A1(n8487), .A2(n8732), .ZN(n8474) );
  XOR2_X1 U9863 ( .A(n8705), .B(n8395), .Z(n8707) );
  AOI21_X1 U9864 ( .B1(n8392), .B2(P2_B_REG_SCAN_IN), .A(n8694), .ZN(n8427) );
  NAND2_X1 U9865 ( .A1(n8427), .A2(n4638), .ZN(n8710) );
  NOR2_X1 U9866 ( .A1(n9775), .A2(n8710), .ZN(n8397) );
  AOI21_X1 U9867 ( .B1(P2_REG2_REG_31__SCAN_IN), .B2(n9775), .A(n8397), .ZN(
        n8394) );
  NAND2_X1 U9868 ( .A1(n8705), .A2(n8698), .ZN(n8393) );
  OAI211_X1 U9869 ( .C1(n8707), .C2(n9754), .A(n8394), .B(n8393), .ZN(P2_U3265) );
  INV_X1 U9870 ( .A(n8396), .ZN(n8712) );
  INV_X1 U9871 ( .A(n8395), .ZN(n8709) );
  NAND2_X1 U9872 ( .A1(n8430), .A2(n8396), .ZN(n8708) );
  NAND3_X1 U9873 ( .A1(n8709), .A2(n9733), .A3(n8708), .ZN(n8399) );
  AOI21_X1 U9874 ( .B1(n9775), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8397), .ZN(
        n8398) );
  OAI211_X1 U9875 ( .C1(n8712), .C2(n9777), .A(n8399), .B(n8398), .ZN(P2_U3266) );
  NAND2_X1 U9876 ( .A1(n8400), .A2(n9735), .ZN(n8401) );
  OR2_X1 U9877 ( .A1(n8697), .A2(n8403), .ZN(n8404) );
  NAND2_X1 U9878 ( .A1(n8797), .A2(n8405), .ZN(n8406) );
  OR2_X1 U9879 ( .A1(n8791), .A2(n8407), .ZN(n8408) );
  NOR2_X1 U9880 ( .A1(n8786), .A2(n8409), .ZN(n8410) );
  AOI21_X2 U9881 ( .B1(n8634), .B2(n8643), .A(n8410), .ZN(n8621) );
  INV_X1 U9882 ( .A(n8771), .ZN(n8592) );
  INV_X1 U9883 ( .A(n8767), .ZN(n8576) );
  INV_X1 U9884 ( .A(n8756), .ZN(n8546) );
  NAND2_X1 U9885 ( .A1(n8543), .A2(n4835), .ZN(n8414) );
  INV_X1 U9886 ( .A(n8751), .ZN(n8530) );
  NAND2_X1 U9887 ( .A1(n8520), .A2(n8519), .ZN(n8521) );
  INV_X1 U9888 ( .A(n8713), .ZN(n8437) );
  OAI21_X1 U9889 ( .B1(n8438), .B2(n8423), .A(n8422), .ZN(n8425) );
  AND2_X1 U9890 ( .A1(n8425), .A2(n8424), .ZN(n8429) );
  AOI22_X1 U9891 ( .A1(n8463), .A2(n9762), .B1(n8427), .B2(n8426), .ZN(n8428)
         );
  OAI21_X1 U9892 ( .B1(n8429), .B2(n8690), .A(n8428), .ZN(n8717) );
  OAI21_X1 U9893 ( .B1(n8444), .B2(n8714), .A(n8430), .ZN(n8715) );
  NOR2_X1 U9894 ( .A1(n8715), .A2(n9754), .ZN(n8435) );
  INV_X1 U9895 ( .A(n8431), .ZN(n8432) );
  AOI22_X1 U9896 ( .A1(n9775), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8432), .B2(
        n9773), .ZN(n8433) );
  OAI21_X1 U9897 ( .B1(n8714), .B2(n9777), .A(n8433), .ZN(n8434) );
  AOI211_X1 U9898 ( .C1(n8717), .C2(n9779), .A(n8435), .B(n8434), .ZN(n8436)
         );
  OAI21_X1 U9899 ( .B1(n8437), .B2(n8703), .A(n8436), .ZN(P2_U3267) );
  AOI211_X1 U9900 ( .C1(n8439), .C2(n8450), .A(n8690), .B(n8438), .ZN(n8443)
         );
  OAI22_X1 U9901 ( .A1(n8441), .A2(n8694), .B1(n8440), .B2(n8692), .ZN(n8442)
         );
  NOR2_X1 U9902 ( .A1(n8443), .A2(n8442), .ZN(n8723) );
  INV_X1 U9903 ( .A(n8456), .ZN(n8445) );
  AOI21_X1 U9904 ( .B1(n8720), .B2(n8445), .A(n8444), .ZN(n8721) );
  AOI22_X1 U9905 ( .A1(n9775), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8446), .B2(
        n9773), .ZN(n8447) );
  OAI21_X1 U9906 ( .B1(n8448), .B2(n9777), .A(n8447), .ZN(n8449) );
  AOI21_X1 U9907 ( .B1(n8721), .B2(n9733), .A(n8449), .ZN(n8453) );
  INV_X1 U9908 ( .A(n8450), .ZN(n8451) );
  OR2_X1 U9909 ( .A1(n8724), .A2(n8703), .ZN(n8452) );
  OAI211_X1 U9910 ( .C1(n8723), .C2(n9775), .A(n8453), .B(n8452), .ZN(P2_U3268) );
  XNOR2_X1 U9911 ( .A(n8454), .B(n8455), .ZN(n8729) );
  AOI21_X1 U9912 ( .B1(n8725), .B2(n8474), .A(n8456), .ZN(n8726) );
  INV_X1 U9913 ( .A(n8457), .ZN(n8458) );
  AOI22_X1 U9914 ( .A1(n9775), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8458), .B2(
        n9773), .ZN(n8459) );
  OAI21_X1 U9915 ( .B1(n8460), .B2(n9777), .A(n8459), .ZN(n8467) );
  XNOR2_X1 U9916 ( .A(n8462), .B(n8461), .ZN(n8465) );
  AOI222_X1 U9917 ( .A1(n9769), .A2(n8465), .B1(n8464), .B2(n9762), .C1(n8463), 
        .C2(n9764), .ZN(n8728) );
  NOR2_X1 U9918 ( .A1(n8728), .A2(n9775), .ZN(n8466) );
  AOI211_X1 U9919 ( .C1(n9733), .C2(n8726), .A(n8467), .B(n8466), .ZN(n8468)
         );
  OAI21_X1 U9920 ( .B1(n8729), .B2(n8703), .A(n8468), .ZN(P2_U3269) );
  XNOR2_X1 U9921 ( .A(n8470), .B(n8469), .ZN(n8734) );
  OAI21_X1 U9922 ( .B1(n8473), .B2(n8690), .A(n8472), .ZN(n8730) );
  INV_X1 U9923 ( .A(n8474), .ZN(n8475) );
  AOI211_X1 U9924 ( .C1(n8732), .C2(n8487), .A(n9889), .B(n8475), .ZN(n8731)
         );
  NAND2_X1 U9925 ( .A1(n8731), .A2(n8585), .ZN(n8478) );
  AOI22_X1 U9926 ( .A1(n9775), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8476), .B2(
        n9773), .ZN(n8477) );
  OAI211_X1 U9927 ( .C1(n8479), .C2(n9777), .A(n8478), .B(n8477), .ZN(n8480)
         );
  AOI21_X1 U9928 ( .B1(n8730), .B2(n9779), .A(n8480), .ZN(n8481) );
  OAI21_X1 U9929 ( .B1(n8734), .B2(n8703), .A(n8481), .ZN(P2_U3270) );
  XOR2_X1 U9930 ( .A(n8483), .B(n8482), .Z(n8739) );
  XNOR2_X1 U9931 ( .A(n8484), .B(n8483), .ZN(n8486) );
  OAI21_X1 U9932 ( .B1(n8486), .B2(n8690), .A(n8485), .ZN(n8735) );
  AOI211_X1 U9933 ( .C1(n8737), .C2(n4271), .A(n9889), .B(n4555), .ZN(n8736)
         );
  NAND2_X1 U9934 ( .A1(n8736), .A2(n8585), .ZN(n8490) );
  AOI22_X1 U9935 ( .A1(n9775), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8488), .B2(
        n9773), .ZN(n8489) );
  OAI211_X1 U9936 ( .C1(n8491), .C2(n9777), .A(n8490), .B(n8489), .ZN(n8492)
         );
  AOI21_X1 U9937 ( .B1(n8735), .B2(n9779), .A(n8492), .ZN(n8493) );
  OAI21_X1 U9938 ( .B1(n8739), .B2(n8703), .A(n8493), .ZN(P2_U3271) );
  AOI21_X1 U9939 ( .B1(n8495), .B2(n8500), .A(n8494), .ZN(n8744) );
  XNOR2_X1 U9940 ( .A(n8513), .B(n8740), .ZN(n8741) );
  AOI22_X1 U9941 ( .A1(n9775), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8496), .B2(
        n9773), .ZN(n8497) );
  OAI21_X1 U9942 ( .B1(n8498), .B2(n9777), .A(n8497), .ZN(n8505) );
  XNOR2_X1 U9943 ( .A(n8499), .B(n8500), .ZN(n8503) );
  AOI222_X1 U9944 ( .A1(n9769), .A2(n8503), .B1(n8502), .B2(n9764), .C1(n8501), 
        .C2(n9762), .ZN(n8743) );
  NOR2_X1 U9945 ( .A1(n8743), .A2(n9775), .ZN(n8504) );
  AOI211_X1 U9946 ( .C1(n8741), .C2(n9733), .A(n8505), .B(n8504), .ZN(n8506)
         );
  OAI21_X1 U9947 ( .B1(n8744), .B2(n8703), .A(n8506), .ZN(P2_U3272) );
  INV_X1 U9948 ( .A(n8507), .ZN(n8535) );
  OAI21_X1 U9949 ( .B1(n8535), .B2(n8508), .A(n8519), .ZN(n8510) );
  NAND2_X1 U9950 ( .A1(n8510), .A2(n8509), .ZN(n8512) );
  AOI222_X1 U9951 ( .A1(n9769), .A2(n8512), .B1(n8549), .B2(n9762), .C1(n8511), 
        .C2(n9764), .ZN(n8750) );
  INV_X1 U9952 ( .A(n8526), .ZN(n8514) );
  AOI21_X1 U9953 ( .B1(n8745), .B2(n8514), .A(n8513), .ZN(n8746) );
  AOI22_X1 U9954 ( .A1(n9775), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8515), .B2(
        n9773), .ZN(n8516) );
  OAI21_X1 U9955 ( .B1(n8517), .B2(n9777), .A(n8516), .ZN(n8518) );
  AOI21_X1 U9956 ( .B1(n8746), .B2(n9733), .A(n8518), .ZN(n8524) );
  OR2_X1 U9957 ( .A1(n8520), .A2(n8519), .ZN(n8747) );
  NAND3_X1 U9958 ( .A1(n8747), .A2(n8521), .A3(n8522), .ZN(n8523) );
  OAI211_X1 U9959 ( .C1(n8750), .C2(n9775), .A(n8524), .B(n8523), .ZN(P2_U3273) );
  XNOR2_X1 U9960 ( .A(n8525), .B(n8532), .ZN(n8755) );
  AOI21_X1 U9961 ( .B1(n8751), .B2(n8527), .A(n8526), .ZN(n8752) );
  AOI22_X1 U9962 ( .A1(n9775), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8528), .B2(
        n9773), .ZN(n8529) );
  OAI21_X1 U9963 ( .B1(n8530), .B2(n9777), .A(n8529), .ZN(n8541) );
  AOI21_X1 U9964 ( .B1(n8531), .B2(n8533), .A(n8532), .ZN(n8534) );
  NOR3_X1 U9965 ( .A1(n8535), .A2(n8534), .A3(n8690), .ZN(n8539) );
  OAI22_X1 U9966 ( .A1(n8537), .A2(n8694), .B1(n8536), .B2(n8692), .ZN(n8538)
         );
  NOR2_X1 U9967 ( .A1(n8539), .A2(n8538), .ZN(n8754) );
  NOR2_X1 U9968 ( .A1(n8754), .A2(n9775), .ZN(n8540) );
  AOI211_X1 U9969 ( .C1(n8752), .C2(n9733), .A(n8541), .B(n8540), .ZN(n8542)
         );
  OAI21_X1 U9970 ( .B1(n8755), .B2(n8703), .A(n8542), .ZN(P2_U3274) );
  XNOR2_X1 U9971 ( .A(n8543), .B(n8547), .ZN(n8760) );
  XNOR2_X1 U9972 ( .A(n8556), .B(n8546), .ZN(n8757) );
  AOI22_X1 U9973 ( .A1(n9775), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8544), .B2(
        n9773), .ZN(n8545) );
  OAI21_X1 U9974 ( .B1(n8546), .B2(n9777), .A(n8545), .ZN(n8552) );
  OAI21_X1 U9975 ( .B1(n8548), .B2(n8547), .A(n8531), .ZN(n8550) );
  AOI222_X1 U9976 ( .A1(n9769), .A2(n8550), .B1(n8581), .B2(n9762), .C1(n8549), 
        .C2(n9764), .ZN(n8759) );
  NOR2_X1 U9977 ( .A1(n8759), .A2(n9775), .ZN(n8551) );
  AOI211_X1 U9978 ( .C1(n8757), .C2(n9733), .A(n8552), .B(n8551), .ZN(n8553)
         );
  OAI21_X1 U9979 ( .B1(n8703), .B2(n8760), .A(n8553), .ZN(P2_U3275) );
  XNOR2_X1 U9980 ( .A(n8555), .B(n8554), .ZN(n8765) );
  INV_X1 U9981 ( .A(n8573), .ZN(n8558) );
  INV_X1 U9982 ( .A(n8556), .ZN(n8557) );
  AOI21_X1 U9983 ( .B1(n8761), .B2(n8558), .A(n8557), .ZN(n8762) );
  AOI22_X1 U9984 ( .A1(n9775), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8559), .B2(
        n9773), .ZN(n8560) );
  OAI21_X1 U9985 ( .B1(n8561), .B2(n9777), .A(n8560), .ZN(n8570) );
  INV_X1 U9986 ( .A(n8562), .ZN(n8566) );
  AOI21_X1 U9987 ( .B1(n8577), .B2(n8564), .A(n8563), .ZN(n8565) );
  NOR3_X1 U9988 ( .A1(n8566), .A2(n8565), .A3(n8690), .ZN(n8568) );
  NOR2_X1 U9989 ( .A1(n8568), .A2(n8567), .ZN(n8764) );
  NOR2_X1 U9990 ( .A1(n8764), .A2(n9775), .ZN(n8569) );
  AOI211_X1 U9991 ( .C1(n8762), .C2(n9733), .A(n8570), .B(n8569), .ZN(n8571)
         );
  OAI21_X1 U9992 ( .B1(n8703), .B2(n8765), .A(n8571), .ZN(P2_U3276) );
  XNOR2_X1 U9993 ( .A(n8572), .B(n8579), .ZN(n8770) );
  AOI211_X1 U9994 ( .C1(n8767), .C2(n8588), .A(n9889), .B(n8573), .ZN(n8766)
         );
  AOI22_X1 U9995 ( .A1(n9775), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8574), .B2(
        n9773), .ZN(n8575) );
  OAI21_X1 U9996 ( .B1(n8576), .B2(n9777), .A(n8575), .ZN(n8584) );
  OAI21_X1 U9997 ( .B1(n8579), .B2(n8578), .A(n8577), .ZN(n8582) );
  AOI222_X1 U9998 ( .A1(n9769), .A2(n8582), .B1(n8581), .B2(n9764), .C1(n8580), 
        .C2(n9762), .ZN(n8769) );
  NOR2_X1 U9999 ( .A1(n8769), .A2(n9775), .ZN(n8583) );
  AOI211_X1 U10000 ( .C1(n8766), .C2(n8585), .A(n8584), .B(n8583), .ZN(n8586)
         );
  OAI21_X1 U10001 ( .B1(n8703), .B2(n8770), .A(n8586), .ZN(P2_U3277) );
  XNOR2_X1 U10002 ( .A(n8587), .B(n8594), .ZN(n8775) );
  INV_X1 U10003 ( .A(n8588), .ZN(n8589) );
  AOI21_X1 U10004 ( .B1(n8771), .B2(n8610), .A(n8589), .ZN(n8772) );
  AOI22_X1 U10005 ( .A1(n9775), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8590), .B2(
        n9773), .ZN(n8591) );
  OAI21_X1 U10006 ( .B1(n8592), .B2(n9777), .A(n8591), .ZN(n8600) );
  OAI21_X1 U10007 ( .B1(n8595), .B2(n8594), .A(n8593), .ZN(n8598) );
  AOI222_X1 U10008 ( .A1(n9769), .A2(n8598), .B1(n8597), .B2(n9764), .C1(n8596), .C2(n9762), .ZN(n8774) );
  NOR2_X1 U10009 ( .A1(n8774), .A2(n9775), .ZN(n8599) );
  AOI211_X1 U10010 ( .C1(n8772), .C2(n9733), .A(n8600), .B(n8599), .ZN(n8601)
         );
  OAI21_X1 U10011 ( .B1(n8775), .B2(n8703), .A(n8601), .ZN(P2_U3278) );
  OAI21_X1 U10012 ( .B1(n8604), .B2(n8603), .A(n8602), .ZN(n8605) );
  INV_X1 U10013 ( .A(n8605), .ZN(n8780) );
  XNOR2_X1 U10014 ( .A(n8607), .B(n8606), .ZN(n8608) );
  OAI222_X1 U10015 ( .A1(n8694), .A2(n8609), .B1(n8692), .B2(n8644), .C1(n8608), .C2(n8690), .ZN(n8776) );
  INV_X1 U10016 ( .A(n8610), .ZN(n8611) );
  AOI211_X1 U10017 ( .C1(n8778), .C2(n8625), .A(n9889), .B(n8611), .ZN(n8777)
         );
  INV_X1 U10018 ( .A(n8777), .ZN(n8614) );
  OAI22_X1 U10019 ( .A1(n8614), .A2(n6456), .B1(n8613), .B2(n8612), .ZN(n8615)
         );
  OAI21_X1 U10020 ( .B1(n8776), .B2(n8615), .A(n9779), .ZN(n8617) );
  AOI22_X1 U10021 ( .A1(n8778), .A2(n8698), .B1(n9775), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n8616) );
  OAI211_X1 U10022 ( .C1(n8780), .C2(n8703), .A(n8617), .B(n8616), .ZN(
        P2_U3279) );
  XOR2_X1 U10023 ( .A(n8620), .B(n8618), .Z(n8624) );
  OAI22_X1 U10024 ( .A1(n8660), .A2(n8692), .B1(n8619), .B2(n8694), .ZN(n8623)
         );
  XNOR2_X1 U10025 ( .A(n8621), .B(n8620), .ZN(n8785) );
  NOR2_X1 U10026 ( .A1(n8785), .A2(n9757), .ZN(n8622) );
  AOI211_X1 U10027 ( .C1(n8624), .C2(n9769), .A(n8623), .B(n8622), .ZN(n8784)
         );
  INV_X1 U10028 ( .A(n8636), .ZN(n8627) );
  INV_X1 U10029 ( .A(n8625), .ZN(n8626) );
  AOI21_X1 U10030 ( .B1(n8781), .B2(n8627), .A(n8626), .ZN(n8782) );
  AOI22_X1 U10031 ( .A1(n9775), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8628), .B2(
        n9773), .ZN(n8629) );
  OAI21_X1 U10032 ( .B1(n8630), .B2(n9777), .A(n8629), .ZN(n8632) );
  NOR2_X1 U10033 ( .A1(n8785), .A2(n9755), .ZN(n8631) );
  AOI211_X1 U10034 ( .C1(n8782), .C2(n9733), .A(n8632), .B(n8631), .ZN(n8633)
         );
  OAI21_X1 U10035 ( .B1(n8784), .B2(n9775), .A(n8633), .ZN(P2_U3280) );
  XNOR2_X1 U10036 ( .A(n8634), .B(n4628), .ZN(n8790) );
  INV_X1 U10037 ( .A(n8635), .ZN(n8637) );
  AOI21_X1 U10038 ( .B1(n8786), .B2(n8637), .A(n8636), .ZN(n8787) );
  AOI22_X1 U10039 ( .A1(n9775), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8638), .B2(
        n9773), .ZN(n8639) );
  OAI21_X1 U10040 ( .B1(n8640), .B2(n9777), .A(n8639), .ZN(n8648) );
  AOI211_X1 U10041 ( .C1(n8643), .C2(n8642), .A(n8690), .B(n8641), .ZN(n8646)
         );
  OAI22_X1 U10042 ( .A1(n8644), .A2(n8694), .B1(n8668), .B2(n8692), .ZN(n8645)
         );
  NOR2_X1 U10043 ( .A1(n8646), .A2(n8645), .ZN(n8789) );
  NOR2_X1 U10044 ( .A1(n8789), .A2(n9775), .ZN(n8647) );
  AOI211_X1 U10045 ( .C1(n8787), .C2(n9733), .A(n8648), .B(n8647), .ZN(n8649)
         );
  OAI21_X1 U10046 ( .B1(n8703), .B2(n8790), .A(n8649), .ZN(P2_U3281) );
  INV_X1 U10047 ( .A(n8650), .ZN(n8651) );
  AOI21_X1 U10048 ( .B1(n8653), .B2(n8652), .A(n8651), .ZN(n8795) );
  INV_X1 U10049 ( .A(n4274), .ZN(n8677) );
  XNOR2_X1 U10050 ( .A(n8677), .B(n8791), .ZN(n8792) );
  INV_X1 U10051 ( .A(n8791), .ZN(n8656) );
  AOI22_X1 U10052 ( .A1(n9775), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8654), .B2(
        n9773), .ZN(n8655) );
  OAI21_X1 U10053 ( .B1(n8656), .B2(n9777), .A(n8655), .ZN(n8664) );
  AOI211_X1 U10054 ( .C1(n8659), .C2(n8658), .A(n8690), .B(n8657), .ZN(n8662)
         );
  OAI22_X1 U10055 ( .A1(n8660), .A2(n8694), .B1(n8693), .B2(n8692), .ZN(n8661)
         );
  NOR2_X1 U10056 ( .A1(n8662), .A2(n8661), .ZN(n8794) );
  NOR2_X1 U10057 ( .A1(n8794), .A2(n9775), .ZN(n8663) );
  AOI211_X1 U10058 ( .C1(n8792), .C2(n9733), .A(n8664), .B(n8663), .ZN(n8665)
         );
  OAI21_X1 U10059 ( .B1(n8795), .B2(n8703), .A(n8665), .ZN(P2_U3282) );
  XNOR2_X1 U10060 ( .A(n8666), .B(n8667), .ZN(n8676) );
  OAI22_X1 U10061 ( .A1(n8669), .A2(n8692), .B1(n8668), .B2(n8694), .ZN(n8675)
         );
  NAND2_X1 U10062 ( .A1(n8671), .A2(n8670), .ZN(n8672) );
  NAND2_X1 U10063 ( .A1(n8673), .A2(n8672), .ZN(n8801) );
  NOR2_X1 U10064 ( .A1(n8801), .A2(n9757), .ZN(n8674) );
  AOI211_X1 U10065 ( .C1(n9769), .C2(n8676), .A(n8675), .B(n8674), .ZN(n8800)
         );
  AOI21_X1 U10066 ( .B1(n8797), .B2(n4337), .A(n8677), .ZN(n8798) );
  INV_X1 U10067 ( .A(n8797), .ZN(n8680) );
  AOI22_X1 U10068 ( .A1(n9775), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8678), .B2(
        n9773), .ZN(n8679) );
  OAI21_X1 U10069 ( .B1(n8680), .B2(n9777), .A(n8679), .ZN(n8682) );
  NOR2_X1 U10070 ( .A1(n8801), .A2(n9755), .ZN(n8681) );
  AOI211_X1 U10071 ( .C1(n8798), .C2(n9733), .A(n8682), .B(n8681), .ZN(n8683)
         );
  OAI21_X1 U10072 ( .B1(n8800), .B2(n9775), .A(n8683), .ZN(P2_U3283) );
  INV_X1 U10073 ( .A(n8688), .ZN(n8685) );
  OAI21_X1 U10074 ( .B1(n8686), .B2(n8685), .A(n8684), .ZN(n9893) );
  INV_X1 U10075 ( .A(n9893), .ZN(n8704) );
  XOR2_X1 U10076 ( .A(n8688), .B(n8687), .Z(n8689) );
  OAI222_X1 U10077 ( .A1(n8694), .A2(n8693), .B1(n8692), .B2(n8691), .C1(n8690), .C2(n8689), .ZN(n9891) );
  OAI21_X1 U10078 ( .B1(n8695), .B2(n9888), .A(n4337), .ZN(n9890) );
  AOI22_X1 U10079 ( .A1(n9775), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n8696), .B2(
        n9773), .ZN(n8700) );
  NAND2_X1 U10080 ( .A1(n8698), .A2(n8697), .ZN(n8699) );
  OAI211_X1 U10081 ( .C1(n9890), .C2(n9754), .A(n8700), .B(n8699), .ZN(n8701)
         );
  AOI21_X1 U10082 ( .B1(n9891), .B2(n9779), .A(n8701), .ZN(n8702) );
  OAI21_X1 U10083 ( .B1(n8704), .B2(n8703), .A(n8702), .ZN(P2_U3284) );
  NAND2_X1 U10084 ( .A1(n8705), .A2(n9835), .ZN(n8706) );
  OAI211_X1 U10085 ( .C1(n8707), .C2(n9889), .A(n8706), .B(n8710), .ZN(n8802)
         );
  MUX2_X1 U10086 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8802), .S(n4260), .Z(
        P2_U3551) );
  NAND3_X1 U10087 ( .A1(n8709), .A2(n9836), .A3(n8708), .ZN(n8711) );
  OAI211_X1 U10088 ( .C1(n8712), .C2(n9887), .A(n8711), .B(n8710), .ZN(n8803)
         );
  MUX2_X1 U10089 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8803), .S(n4260), .Z(
        P2_U3550) );
  NAND2_X1 U10090 ( .A1(n8713), .A2(n9894), .ZN(n8719) );
  OAI22_X1 U10091 ( .A1(n8715), .A2(n9889), .B1(n8714), .B2(n9887), .ZN(n8716)
         );
  NOR2_X1 U10092 ( .A1(n8717), .A2(n8716), .ZN(n8718) );
  NAND2_X1 U10093 ( .A1(n8719), .A2(n8718), .ZN(n8804) );
  MUX2_X1 U10094 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8804), .S(n4260), .Z(
        P2_U3549) );
  AOI22_X1 U10095 ( .A1(n8721), .A2(n9836), .B1(n9835), .B2(n8720), .ZN(n8722)
         );
  AOI22_X1 U10096 ( .A1(n8726), .A2(n9836), .B1(n9835), .B2(n8725), .ZN(n8727)
         );
  OAI211_X1 U10097 ( .C1(n8729), .C2(n8796), .A(n8728), .B(n8727), .ZN(n8806)
         );
  MUX2_X1 U10098 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8806), .S(n4260), .Z(
        P2_U3547) );
  OAI21_X1 U10099 ( .B1(n8734), .B2(n8796), .A(n8733), .ZN(n8807) );
  MUX2_X1 U10100 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8807), .S(n4260), .Z(
        P2_U3546) );
  AOI211_X1 U10101 ( .C1(n9835), .C2(n8737), .A(n8736), .B(n8735), .ZN(n8738)
         );
  OAI21_X1 U10102 ( .B1(n8739), .B2(n8796), .A(n8738), .ZN(n8808) );
  MUX2_X1 U10103 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8808), .S(n4260), .Z(
        P2_U3545) );
  AOI22_X1 U10104 ( .A1(n8741), .A2(n9836), .B1(n9835), .B2(n8740), .ZN(n8742)
         );
  OAI211_X1 U10105 ( .C1(n8744), .C2(n8796), .A(n8743), .B(n8742), .ZN(n8809)
         );
  MUX2_X1 U10106 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8809), .S(n4260), .Z(
        P2_U3544) );
  AOI22_X1 U10107 ( .A1(n8746), .A2(n9836), .B1(n9835), .B2(n8745), .ZN(n8749)
         );
  NAND3_X1 U10108 ( .A1(n8747), .A2(n8521), .A3(n9894), .ZN(n8748) );
  NAND3_X1 U10109 ( .A1(n8750), .A2(n8749), .A3(n8748), .ZN(n8810) );
  MUX2_X1 U10110 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8810), .S(n4260), .Z(
        P2_U3543) );
  AOI22_X1 U10111 ( .A1(n8752), .A2(n9836), .B1(n9835), .B2(n8751), .ZN(n8753)
         );
  OAI211_X1 U10112 ( .C1(n8755), .C2(n8796), .A(n8754), .B(n8753), .ZN(n8811)
         );
  MUX2_X1 U10113 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8811), .S(n4260), .Z(
        P2_U3542) );
  AOI22_X1 U10114 ( .A1(n8757), .A2(n9836), .B1(n9835), .B2(n8756), .ZN(n8758)
         );
  OAI211_X1 U10115 ( .C1(n8796), .C2(n8760), .A(n8759), .B(n8758), .ZN(n8812)
         );
  MUX2_X1 U10116 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8812), .S(n4260), .Z(
        P2_U3541) );
  AOI22_X1 U10117 ( .A1(n8762), .A2(n9836), .B1(n9835), .B2(n8761), .ZN(n8763)
         );
  OAI211_X1 U10118 ( .C1(n8796), .C2(n8765), .A(n8764), .B(n8763), .ZN(n8813)
         );
  MUX2_X1 U10119 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8813), .S(n4260), .Z(
        P2_U3540) );
  AOI21_X1 U10120 ( .B1(n9835), .B2(n8767), .A(n8766), .ZN(n8768) );
  OAI211_X1 U10121 ( .C1(n8796), .C2(n8770), .A(n8769), .B(n8768), .ZN(n8814)
         );
  MUX2_X1 U10122 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8814), .S(n4260), .Z(
        P2_U3539) );
  AOI22_X1 U10123 ( .A1(n8772), .A2(n9836), .B1(n9835), .B2(n8771), .ZN(n8773)
         );
  OAI211_X1 U10124 ( .C1(n8796), .C2(n8775), .A(n8774), .B(n8773), .ZN(n8815)
         );
  MUX2_X1 U10125 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8815), .S(n4260), .Z(
        P2_U3538) );
  AOI211_X1 U10126 ( .C1(n9835), .C2(n8778), .A(n8777), .B(n8776), .ZN(n8779)
         );
  OAI21_X1 U10127 ( .B1(n8796), .B2(n8780), .A(n8779), .ZN(n8816) );
  MUX2_X1 U10128 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8816), .S(n4260), .Z(
        P2_U3537) );
  AOI22_X1 U10129 ( .A1(n8782), .A2(n9836), .B1(n9835), .B2(n8781), .ZN(n8783)
         );
  OAI211_X1 U10130 ( .C1(n8785), .C2(n9856), .A(n8784), .B(n8783), .ZN(n8817)
         );
  MUX2_X1 U10131 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8817), .S(n4260), .Z(
        P2_U3536) );
  AOI22_X1 U10132 ( .A1(n8787), .A2(n9836), .B1(n9835), .B2(n8786), .ZN(n8788)
         );
  OAI211_X1 U10133 ( .C1(n8796), .C2(n8790), .A(n8789), .B(n8788), .ZN(n8818)
         );
  MUX2_X1 U10134 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8818), .S(n4260), .Z(
        P2_U3535) );
  AOI22_X1 U10135 ( .A1(n8792), .A2(n9836), .B1(n9835), .B2(n8791), .ZN(n8793)
         );
  OAI211_X1 U10136 ( .C1(n8796), .C2(n8795), .A(n8794), .B(n8793), .ZN(n8819)
         );
  MUX2_X1 U10137 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8819), .S(n4260), .Z(
        P2_U3534) );
  AOI22_X1 U10138 ( .A1(n8798), .A2(n9836), .B1(n9835), .B2(n8797), .ZN(n8799)
         );
  OAI211_X1 U10139 ( .C1(n9856), .C2(n8801), .A(n8800), .B(n8799), .ZN(n8820)
         );
  MUX2_X1 U10140 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8820), .S(n4260), .Z(
        P2_U3533) );
  MUX2_X1 U10141 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8802), .S(n9872), .Z(
        P2_U3519) );
  MUX2_X1 U10142 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8803), .S(n9872), .Z(
        P2_U3518) );
  MUX2_X1 U10143 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8804), .S(n9872), .Z(
        P2_U3517) );
  MUX2_X1 U10144 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8805), .S(n9872), .Z(
        P2_U3516) );
  MUX2_X1 U10145 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8806), .S(n9872), .Z(
        P2_U3515) );
  MUX2_X1 U10146 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8807), .S(n9872), .Z(
        P2_U3514) );
  MUX2_X1 U10147 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8808), .S(n9872), .Z(
        P2_U3513) );
  MUX2_X1 U10148 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8809), .S(n9872), .Z(
        P2_U3512) );
  MUX2_X1 U10149 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8810), .S(n9872), .Z(
        P2_U3511) );
  MUX2_X1 U10150 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8811), .S(n9872), .Z(
        P2_U3510) );
  MUX2_X1 U10151 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8812), .S(n9872), .Z(
        P2_U3509) );
  MUX2_X1 U10152 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8813), .S(n9872), .Z(
        P2_U3508) );
  MUX2_X1 U10153 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8814), .S(n9872), .Z(
        P2_U3507) );
  MUX2_X1 U10154 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8815), .S(n9872), .Z(
        P2_U3505) );
  MUX2_X1 U10155 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8816), .S(n9872), .Z(
        P2_U3502) );
  MUX2_X1 U10156 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8817), .S(n9872), .Z(
        P2_U3499) );
  MUX2_X1 U10157 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8818), .S(n9872), .Z(
        P2_U3496) );
  MUX2_X1 U10158 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8819), .S(n9872), .Z(
        P2_U3493) );
  MUX2_X1 U10159 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8820), .S(n9872), .Z(
        P2_U3490) );
  INV_X1 U10160 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8821) );
  NAND3_X1 U10161 ( .A1(n8821), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8823) );
  OAI22_X1 U10162 ( .A1(n6216), .A2(n8823), .B1(n8822), .B2(n8830), .ZN(n8824)
         );
  AOI21_X1 U10163 ( .B1(n9534), .B2(n8825), .A(n8824), .ZN(n8826) );
  INV_X1 U10164 ( .A(n8826), .ZN(P2_U3327) );
  INV_X1 U10165 ( .A(n8827), .ZN(n9553) );
  OAI222_X1 U10166 ( .A1(n8830), .A2(n8829), .B1(n7667), .B2(n9553), .C1(n8828), .C2(P2_U3152), .ZN(P2_U3331) );
  MUX2_X1 U10167 ( .A(n8831), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XOR2_X1 U10168 ( .A(n8833), .B(n8832), .Z(n8834) );
  XNOR2_X1 U10169 ( .A(n8835), .B(n8834), .ZN(n8841) );
  NAND2_X1 U10170 ( .A1(n8984), .A2(n8994), .ZN(n8837) );
  OAI211_X1 U10171 ( .C1(n8987), .C2(n9390), .A(n8837), .B(n8836), .ZN(n8839)
         );
  INV_X1 U10172 ( .A(n9495), .ZN(n9361) );
  NOR2_X1 U10173 ( .A1(n9361), .A2(n8977), .ZN(n8838) );
  AOI211_X1 U10174 ( .C1(n9358), .C2(n8982), .A(n8839), .B(n8838), .ZN(n8840)
         );
  OAI21_X1 U10175 ( .B1(n8841), .B2(n8991), .A(n8840), .ZN(P1_U3213) );
  INV_X1 U10176 ( .A(n8842), .ZN(n8844) );
  NAND2_X1 U10177 ( .A1(n8844), .A2(n8843), .ZN(n8846) );
  XNOR2_X1 U10178 ( .A(n8846), .B(n8845), .ZN(n8853) );
  INV_X1 U10179 ( .A(n8847), .ZN(n9222) );
  NAND2_X1 U10180 ( .A1(n8984), .A2(n9192), .ZN(n8849) );
  NAND2_X1 U10181 ( .A1(P1_U3084), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8848) );
  OAI211_X1 U10182 ( .C1(n8987), .C2(n9248), .A(n8849), .B(n8848), .ZN(n8850)
         );
  AOI21_X1 U10183 ( .B1(n9222), .B2(n8982), .A(n8850), .ZN(n8852) );
  NAND2_X1 U10184 ( .A1(n9447), .A2(n8989), .ZN(n8851) );
  OAI211_X1 U10185 ( .C1(n8853), .C2(n8991), .A(n8852), .B(n8851), .ZN(
        P1_U3214) );
  INV_X1 U10186 ( .A(n8854), .ZN(n8856) );
  NOR2_X1 U10187 ( .A1(n8856), .A2(n8855), .ZN(n8857) );
  XNOR2_X1 U10188 ( .A(n8858), .B(n8857), .ZN(n8864) );
  NAND2_X1 U10189 ( .A1(n8982), .A2(n9279), .ZN(n8861) );
  NOR2_X1 U10190 ( .A1(n8859), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9037) );
  AOI21_X1 U10191 ( .B1(n8984), .B2(n9073), .A(n9037), .ZN(n8860) );
  OAI211_X1 U10192 ( .C1(n9275), .C2(n8987), .A(n8861), .B(n8860), .ZN(n8862)
         );
  AOI21_X1 U10193 ( .B1(n9468), .B2(n8989), .A(n8862), .ZN(n8863) );
  OAI21_X1 U10194 ( .B1(n8864), .B2(n8991), .A(n8863), .ZN(P1_U3217) );
  NAND2_X1 U10195 ( .A1(n8866), .A2(n8865), .ZN(n8867) );
  XNOR2_X1 U10196 ( .A(n4283), .B(n8867), .ZN(n8872) );
  NAND2_X1 U10197 ( .A1(n8982), .A2(n9243), .ZN(n8869) );
  AOI22_X1 U10198 ( .A1(n8984), .A2(n9075), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8868) );
  OAI211_X1 U10199 ( .C1(n9274), .C2(n8987), .A(n8869), .B(n8868), .ZN(n8870)
         );
  AOI21_X1 U10200 ( .B1(n9458), .B2(n8989), .A(n8870), .ZN(n8871) );
  OAI21_X1 U10201 ( .B1(n8872), .B2(n8991), .A(n8871), .ZN(P1_U3221) );
  NAND2_X1 U10202 ( .A1(n8875), .A2(n8874), .ZN(n8876) );
  XNOR2_X1 U10203 ( .A(n8873), .B(n8876), .ZN(n8883) );
  INV_X1 U10204 ( .A(n9506), .ZN(n9403) );
  NOR2_X1 U10205 ( .A1(n8977), .A2(n9403), .ZN(n8882) );
  NAND2_X1 U10206 ( .A1(n8982), .A2(n9401), .ZN(n8880) );
  INV_X1 U10207 ( .A(n8877), .ZN(n8878) );
  AOI21_X1 U10208 ( .B1(n8984), .B2(n9061), .A(n8878), .ZN(n8879) );
  OAI211_X1 U10209 ( .C1(n9391), .C2(n8987), .A(n8880), .B(n8879), .ZN(n8881)
         );
  AOI211_X1 U10210 ( .C1(n8883), .C2(n8970), .A(n8882), .B(n8881), .ZN(n8884)
         );
  INV_X1 U10211 ( .A(n8884), .ZN(P1_U3222) );
  AOI21_X1 U10212 ( .B1(n8886), .B2(n8885), .A(n8968), .ZN(n8891) );
  AOI22_X1 U10213 ( .A1(n9193), .A2(n8984), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8888) );
  NAND2_X1 U10214 ( .A1(n8982), .A2(n9187), .ZN(n8887) );
  OAI211_X1 U10215 ( .C1(n9218), .C2(n8987), .A(n8888), .B(n8887), .ZN(n8889)
         );
  AOI21_X1 U10216 ( .B1(n9435), .B2(n8989), .A(n8889), .ZN(n8890) );
  OAI21_X1 U10217 ( .B1(n8891), .B2(n8991), .A(n8890), .ZN(P1_U3223) );
  INV_X1 U10218 ( .A(n8893), .ZN(n8895) );
  NOR2_X1 U10219 ( .A1(n8895), .A2(n8894), .ZN(n8896) );
  XNOR2_X1 U10220 ( .A(n8892), .B(n8896), .ZN(n8902) );
  NAND2_X1 U10221 ( .A1(n8984), .A2(n9296), .ZN(n8898) );
  OAI211_X1 U10222 ( .C1(n8987), .C2(n9355), .A(n8898), .B(n8897), .ZN(n8900)
         );
  NOR2_X1 U10223 ( .A1(n4445), .A2(n8977), .ZN(n8899) );
  AOI211_X1 U10224 ( .C1(n9326), .C2(n8982), .A(n8900), .B(n8899), .ZN(n8901)
         );
  OAI21_X1 U10225 ( .B1(n8902), .B2(n8991), .A(n8901), .ZN(P1_U3224) );
  AOI21_X1 U10226 ( .B1(n8905), .B2(n8904), .A(n8903), .ZN(n8911) );
  NOR2_X1 U10227 ( .A1(n8906), .A2(n9206), .ZN(n8909) );
  AOI22_X1 U10228 ( .A1(n9177), .A2(n8984), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8907) );
  OAI21_X1 U10229 ( .B1(n9203), .B2(n8987), .A(n8907), .ZN(n8908) );
  AOI211_X1 U10230 ( .C1(n9442), .C2(n8989), .A(n8909), .B(n8908), .ZN(n8910)
         );
  OAI21_X1 U10231 ( .B1(n8911), .B2(n8991), .A(n8910), .ZN(P1_U3227) );
  INV_X1 U10232 ( .A(n9463), .ZN(n9267) );
  OAI21_X1 U10233 ( .B1(n5865), .B2(n8915), .A(n8914), .ZN(n8916) );
  OAI211_X1 U10234 ( .C1(n8917), .C2(n5865), .A(n8970), .B(n8916), .ZN(n8921)
         );
  INV_X1 U10235 ( .A(n9262), .ZN(n9234) );
  AOI22_X1 U10236 ( .A1(n8984), .A2(n9234), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8918) );
  OAI21_X1 U10237 ( .B1(n9263), .B2(n8987), .A(n8918), .ZN(n8919) );
  AOI21_X1 U10238 ( .B1(n9264), .B2(n8982), .A(n8919), .ZN(n8920) );
  OAI211_X1 U10239 ( .C1(n9267), .C2(n8977), .A(n8921), .B(n8920), .ZN(
        P1_U3231) );
  XNOR2_X1 U10240 ( .A(n8924), .B(n8923), .ZN(n8925) );
  XNOR2_X1 U10241 ( .A(n8922), .B(n8925), .ZN(n8932) );
  INV_X1 U10242 ( .A(n9499), .ZN(n9380) );
  NOR2_X1 U10243 ( .A1(n9380), .A2(n8977), .ZN(n8931) );
  NAND2_X1 U10244 ( .A1(n8982), .A2(n9378), .ZN(n8929) );
  INV_X1 U10245 ( .A(n9373), .ZN(n9064) );
  INV_X1 U10246 ( .A(n8926), .ZN(n8927) );
  AOI21_X1 U10247 ( .B1(n8984), .B2(n9064), .A(n8927), .ZN(n8928) );
  OAI211_X1 U10248 ( .C1(n9589), .C2(n8987), .A(n8929), .B(n8928), .ZN(n8930)
         );
  AOI211_X1 U10249 ( .C1(n8932), .C2(n8970), .A(n8931), .B(n8930), .ZN(n8933)
         );
  INV_X1 U10250 ( .A(n8933), .ZN(P1_U3232) );
  XNOR2_X1 U10251 ( .A(n8936), .B(n8935), .ZN(n8937) );
  XNOR2_X1 U10252 ( .A(n8934), .B(n8937), .ZN(n8942) );
  NAND2_X1 U10253 ( .A1(n8982), .A2(n9230), .ZN(n8939) );
  AOI22_X1 U10254 ( .A1(n8984), .A2(n9235), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8938) );
  OAI211_X1 U10255 ( .C1(n9262), .C2(n8987), .A(n8939), .B(n8938), .ZN(n8940)
         );
  AOI21_X1 U10256 ( .B1(n9450), .B2(n8989), .A(n8940), .ZN(n8941) );
  OAI21_X1 U10257 ( .B1(n8942), .B2(n8991), .A(n8941), .ZN(P1_U3233) );
  OAI21_X1 U10258 ( .B1(n8943), .B2(n8944), .A(n6890), .ZN(n8945) );
  NAND2_X1 U10259 ( .A1(n8945), .A2(n8970), .ZN(n8951) );
  AOI22_X1 U10260 ( .A1(n8946), .A2(n9005), .B1(n8984), .B2(n9002), .ZN(n8950)
         );
  AOI22_X1 U10261 ( .A1(n8989), .A2(n8948), .B1(n8947), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n8949) );
  NAND3_X1 U10262 ( .A1(n8951), .A2(n8950), .A3(n8949), .ZN(P1_U3235) );
  OR2_X1 U10263 ( .A1(n8953), .A2(n8952), .ZN(n8955) );
  NAND2_X1 U10264 ( .A1(n8955), .A2(n8954), .ZN(n8957) );
  NAND2_X1 U10265 ( .A1(n8957), .A2(n8956), .ZN(n8958) );
  XOR2_X1 U10266 ( .A(n8959), .B(n8958), .Z(n8964) );
  NAND2_X1 U10267 ( .A1(n8982), .A2(n9289), .ZN(n8961) );
  AOI22_X1 U10268 ( .A1(n8984), .A2(n9297), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3084), .ZN(n8960) );
  OAI211_X1 U10269 ( .C1(n9068), .C2(n8987), .A(n8961), .B(n8960), .ZN(n8962)
         );
  AOI21_X1 U10270 ( .B1(n9471), .B2(n8989), .A(n8962), .ZN(n8963) );
  OAI21_X1 U10271 ( .B1(n8964), .B2(n8991), .A(n8963), .ZN(P1_U3236) );
  INV_X1 U10272 ( .A(n8965), .ZN(n8971) );
  OAI21_X1 U10273 ( .B1(n8968), .B2(n8967), .A(n8966), .ZN(n8969) );
  NAND3_X1 U10274 ( .A1(n8971), .A2(n8970), .A3(n8969), .ZN(n8976) );
  INV_X1 U10275 ( .A(n8972), .ZN(n9170) );
  AOI22_X1 U10276 ( .A1(n9178), .A2(n8984), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8973) );
  OAI21_X1 U10277 ( .B1(n9204), .B2(n8987), .A(n8973), .ZN(n8974) );
  AOI21_X1 U10278 ( .B1(n9170), .B2(n8982), .A(n8974), .ZN(n8975) );
  OAI211_X1 U10279 ( .C1(n9172), .C2(n8977), .A(n8976), .B(n8975), .ZN(
        P1_U3238) );
  XNOR2_X1 U10280 ( .A(n8979), .B(n8978), .ZN(n8980) );
  XNOR2_X1 U10281 ( .A(n8981), .B(n8980), .ZN(n8992) );
  NAND2_X1 U10282 ( .A1(n8982), .A2(n9343), .ZN(n8986) );
  INV_X1 U10283 ( .A(n9336), .ZN(n9312) );
  AOI21_X1 U10284 ( .B1(n8984), .B2(n9312), .A(n8983), .ZN(n8985) );
  OAI211_X1 U10285 ( .C1(n9373), .C2(n8987), .A(n8986), .B(n8985), .ZN(n8988)
         );
  AOI21_X1 U10286 ( .B1(n9487), .B2(n8989), .A(n8988), .ZN(n8990) );
  OAI21_X1 U10287 ( .B1(n8992), .B2(n8991), .A(n8990), .ZN(P1_U3239) );
  MUX2_X1 U10288 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9045), .S(n9004), .Z(
        P1_U3586) );
  MUX2_X1 U10289 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9121), .S(n9004), .Z(
        P1_U3585) );
  MUX2_X1 U10290 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n8993), .S(n9004), .Z(
        P1_U3584) );
  MUX2_X1 U10291 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9090), .S(n9004), .Z(
        P1_U3583) );
  MUX2_X1 U10292 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9178), .S(n9004), .Z(
        P1_U3582) );
  MUX2_X1 U10293 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9193), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10294 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9177), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10295 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9192), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10296 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9235), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10297 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9075), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10298 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9234), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10299 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9073), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10300 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9297), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10301 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9310), .S(n9004), .Z(
        P1_U3573) );
  MUX2_X1 U10302 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9296), .S(n9004), .Z(
        P1_U3572) );
  MUX2_X1 U10303 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9312), .S(n9004), .Z(
        P1_U3571) );
  MUX2_X1 U10304 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n8994), .S(n9004), .Z(
        P1_U3570) );
  MUX2_X1 U10305 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9064), .S(n9004), .Z(
        P1_U3569) );
  MUX2_X1 U10306 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9061), .S(n9004), .Z(
        P1_U3568) );
  MUX2_X1 U10307 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9058), .S(n9004), .Z(
        P1_U3567) );
  MUX2_X1 U10308 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9056), .S(n9004), .Z(
        P1_U3566) );
  MUX2_X1 U10309 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n8995), .S(n9004), .Z(
        P1_U3565) );
  MUX2_X1 U10310 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n8996), .S(n9004), .Z(
        P1_U3564) );
  MUX2_X1 U10311 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n8997), .S(n9004), .Z(
        P1_U3563) );
  MUX2_X1 U10312 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8998), .S(n9004), .Z(
        P1_U3562) );
  MUX2_X1 U10313 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8999), .S(n9004), .Z(
        P1_U3561) );
  MUX2_X1 U10314 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9000), .S(n9004), .Z(
        P1_U3560) );
  MUX2_X1 U10315 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9001), .S(n9004), .Z(
        P1_U3559) );
  MUX2_X1 U10316 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9002), .S(n9004), .Z(
        P1_U3558) );
  MUX2_X1 U10317 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9003), .S(n9004), .Z(
        P1_U3557) );
  MUX2_X1 U10318 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9005), .S(n9004), .Z(
        P1_U3556) );
  INV_X1 U10319 ( .A(n9026), .ZN(n9013) );
  NAND2_X1 U10320 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3084), .ZN(n9012) );
  XOR2_X1 U10321 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9026), .Z(n9009) );
  AOI21_X1 U10322 ( .B1(n9015), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9007), .ZN(
        n9008) );
  NAND2_X1 U10323 ( .A1(n9009), .A2(n9008), .ZN(n9025) );
  OAI21_X1 U10324 ( .B1(n9009), .B2(n9008), .A(n9025), .ZN(n9010) );
  NAND2_X1 U10325 ( .A1(n9623), .A2(n9010), .ZN(n9011) );
  OAI211_X1 U10326 ( .C1(n9029), .C2(n9013), .A(n9012), .B(n9011), .ZN(n9021)
         );
  AOI21_X1 U10327 ( .B1(n9015), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9014), .ZN(
        n9019) );
  NAND2_X1 U10328 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n9026), .ZN(n9016) );
  OAI21_X1 U10329 ( .B1(n9026), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9016), .ZN(
        n9018) );
  NOR2_X1 U10330 ( .A1(n9019), .A2(n9018), .ZN(n9023) );
  AOI211_X1 U10331 ( .C1(n9019), .C2(n9018), .A(n9023), .B(n9017), .ZN(n9020)
         );
  AOI211_X1 U10332 ( .C1(P1_ADDR_REG_18__SCAN_IN), .C2(n9611), .A(n9021), .B(
        n9020), .ZN(n9022) );
  INV_X1 U10333 ( .A(n9022), .ZN(P1_U3259) );
  AOI21_X1 U10334 ( .B1(n9026), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9023), .ZN(
        n9024) );
  INV_X1 U10335 ( .A(n9035), .ZN(n9033) );
  OAI21_X1 U10336 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9026), .A(n9025), .ZN(
        n9028) );
  XOR2_X1 U10337 ( .A(n9028), .B(n9027), .Z(n9034) );
  OAI21_X1 U10338 ( .B1(n9034), .B2(n9030), .A(n9029), .ZN(n9031) );
  AOI21_X1 U10339 ( .B1(n9033), .B2(n9032), .A(n9031), .ZN(n9036) );
  INV_X1 U10340 ( .A(n9037), .ZN(n9038) );
  INV_X1 U10341 ( .A(n9487), .ZN(n9345) );
  INV_X1 U10342 ( .A(n9471), .ZN(n9291) );
  INV_X1 U10343 ( .A(n9468), .ZN(n9282) );
  NAND2_X1 U10344 ( .A1(n9229), .A2(n9225), .ZN(n9219) );
  NAND2_X1 U10345 ( .A1(n9205), .A2(n9189), .ZN(n9184) );
  NAND2_X1 U10346 ( .A1(n9169), .A2(n9165), .ZN(n9159) );
  NOR2_X1 U10347 ( .A1(n9125), .A2(n9410), .ZN(n9042) );
  XNOR2_X1 U10348 ( .A(n9042), .B(n9046), .ZN(n9409) );
  AND2_X1 U10349 ( .A1(n9043), .A2(P1_B_REG_SCAN_IN), .ZN(n9044) );
  NOR2_X1 U10350 ( .A1(n9635), .A2(n9044), .ZN(n9122) );
  NAND2_X1 U10351 ( .A1(n9122), .A2(n9045), .ZN(n9412) );
  NOR2_X1 U10352 ( .A1(n9647), .A2(n9412), .ZN(n9049) );
  NOR2_X1 U10353 ( .A1(n9046), .A2(n9595), .ZN(n9047) );
  AOI211_X1 U10354 ( .C1(n9647), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9049), .B(
        n9047), .ZN(n9048) );
  OAI21_X1 U10355 ( .B1(n9409), .B2(n9584), .A(n9048), .ZN(P1_U3261) );
  XNOR2_X1 U10356 ( .A(n9125), .B(n9410), .ZN(n9413) );
  AOI21_X1 U10357 ( .B1(n9647), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9049), .ZN(
        n9051) );
  NAND2_X1 U10358 ( .A1(n9410), .A2(n9254), .ZN(n9050) );
  OAI211_X1 U10359 ( .C1(n9413), .C2(n9584), .A(n9051), .B(n9050), .ZN(
        P1_U3262) );
  NAND2_X1 U10360 ( .A1(n9636), .A2(n9570), .ZN(n9054) );
  NAND2_X1 U10361 ( .A1(n9056), .A2(n9055), .ZN(n9057) );
  NAND2_X1 U10362 ( .A1(n9577), .A2(n9057), .ZN(n9393) );
  NAND2_X1 U10363 ( .A1(n9393), .A2(n9392), .ZN(n9395) );
  NAND2_X1 U10364 ( .A1(n9506), .A2(n9058), .ZN(n9059) );
  NAND2_X1 U10365 ( .A1(n9395), .A2(n9059), .ZN(n9365) );
  OR2_X1 U10366 ( .A1(n9499), .A2(n9061), .ZN(n9060) );
  NAND2_X1 U10367 ( .A1(n9365), .A2(n9060), .ZN(n9063) );
  NAND2_X1 U10368 ( .A1(n9499), .A2(n9061), .ZN(n9062) );
  OR2_X1 U10369 ( .A1(n9495), .A2(n9064), .ZN(n9065) );
  NAND2_X1 U10370 ( .A1(n9320), .A2(n9319), .ZN(n9321) );
  OAI21_X1 U10371 ( .B1(n9336), .B2(n4445), .A(n9321), .ZN(n9303) );
  NAND2_X1 U10372 ( .A1(n9069), .A2(n9068), .ZN(n9070) );
  NAND2_X1 U10373 ( .A1(n9303), .A2(n9070), .ZN(n9071) );
  NOR2_X1 U10374 ( .A1(n9468), .A2(n9297), .ZN(n9072) );
  NAND2_X1 U10375 ( .A1(n9253), .A2(n4831), .ZN(n9228) );
  OR2_X1 U10376 ( .A1(n9450), .A2(n9075), .ZN(n9076) );
  NAND2_X1 U10377 ( .A1(n9228), .A2(n9076), .ZN(n9077) );
  NAND2_X1 U10378 ( .A1(n9077), .A2(n4832), .ZN(n9212) );
  NAND2_X1 U10379 ( .A1(n9225), .A2(n9203), .ZN(n9079) );
  AOI21_X2 U10380 ( .B1(n9212), .B2(n9079), .A(n9078), .ZN(n9198) );
  OAI21_X1 U10381 ( .B1(n9218), .B2(n9080), .A(n9198), .ZN(n9082) );
  NAND2_X1 U10382 ( .A1(n9080), .A2(n9218), .ZN(n9081) );
  AOI21_X2 U10383 ( .B1(n9183), .B2(n9190), .A(n9083), .ZN(n9168) );
  NAND2_X1 U10384 ( .A1(n9172), .A2(n9158), .ZN(n9085) );
  NOR2_X1 U10385 ( .A1(n9172), .A2(n9158), .ZN(n9084) );
  NAND2_X1 U10386 ( .A1(n9165), .A2(n9143), .ZN(n9087) );
  INV_X1 U10387 ( .A(n9423), .ZN(n9149) );
  NAND2_X1 U10388 ( .A1(n9423), .A2(n9090), .ZN(n9091) );
  XNOR2_X1 U10389 ( .A(n9092), .B(n9120), .ZN(n9414) );
  INV_X1 U10390 ( .A(n9414), .ZN(n9133) );
  INV_X1 U10391 ( .A(n9098), .ZN(n9099) );
  NAND2_X1 U10392 ( .A1(n9233), .A2(n9110), .ZN(n9214) );
  INV_X1 U10393 ( .A(n9113), .ZN(n9114) );
  NAND3_X1 U10394 ( .A1(n9138), .A2(n9139), .A3(n9140), .ZN(n9137) );
  NAND2_X1 U10395 ( .A1(n9137), .A2(n9118), .ZN(n9119) );
  XOR2_X1 U10396 ( .A(n9120), .B(n9119), .Z(n9124) );
  AOI22_X1 U10397 ( .A1(n9090), .A2(n9311), .B1(n9122), .B2(n9121), .ZN(n9123)
         );
  OAI21_X1 U10398 ( .B1(n9124), .B2(n9370), .A(n9123), .ZN(n9416) );
  NOR2_X1 U10399 ( .A1(n9415), .A2(n9584), .ZN(n9131) );
  INV_X1 U10400 ( .A(n9126), .ZN(n9127) );
  AOI22_X1 U10401 ( .A1(n9127), .A2(n9645), .B1(n9647), .B2(
        P1_REG2_REG_29__SCAN_IN), .ZN(n9128) );
  OAI21_X1 U10402 ( .B1(n9129), .B2(n9595), .A(n9128), .ZN(n9130) );
  AOI211_X1 U10403 ( .C1(n9416), .C2(n9650), .A(n9131), .B(n9130), .ZN(n9132)
         );
  OAI21_X1 U10404 ( .B1(n9133), .B2(n9364), .A(n9132), .ZN(P1_U3355) );
  NAND2_X1 U10405 ( .A1(n9134), .A2(n9139), .ZN(n9135) );
  INV_X1 U10406 ( .A(n9420), .ZN(n9152) );
  INV_X1 U10407 ( .A(n9137), .ZN(n9142) );
  AOI21_X1 U10408 ( .B1(n9138), .B2(n9140), .A(n9139), .ZN(n9141) );
  AOI211_X1 U10409 ( .C1(n9423), .C2(n9159), .A(n9682), .B(n9145), .ZN(n9422)
         );
  NAND2_X1 U10410 ( .A1(n9422), .A2(n9406), .ZN(n9148) );
  AOI22_X1 U10411 ( .A1(n9146), .A2(n9645), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9647), .ZN(n9147) );
  OAI211_X1 U10412 ( .C1(n9149), .C2(n9595), .A(n9148), .B(n9147), .ZN(n9150)
         );
  AOI21_X1 U10413 ( .B1(n9421), .B2(n9650), .A(n9150), .ZN(n9151) );
  OAI21_X1 U10414 ( .B1(n9152), .B2(n9364), .A(n9151), .ZN(P1_U3263) );
  XNOR2_X1 U10415 ( .A(n9153), .B(n9154), .ZN(n9429) );
  OAI211_X1 U10416 ( .C1(n9155), .C2(n9154), .A(n9138), .B(n9640), .ZN(n9157)
         );
  NAND2_X1 U10417 ( .A1(n9090), .A2(n9309), .ZN(n9156) );
  OAI211_X1 U10418 ( .C1(n9158), .C2(n9638), .A(n9157), .B(n9156), .ZN(n9425)
         );
  INV_X1 U10419 ( .A(n9169), .ZN(n9161) );
  INV_X1 U10420 ( .A(n9159), .ZN(n9160) );
  AOI211_X1 U10421 ( .C1(n9427), .C2(n9161), .A(n9682), .B(n9160), .ZN(n9426)
         );
  NAND2_X1 U10422 ( .A1(n9426), .A2(n9406), .ZN(n9164) );
  AOI22_X1 U10423 ( .A1(n9647), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9162), .B2(
        n9645), .ZN(n9163) );
  OAI211_X1 U10424 ( .C1(n9165), .C2(n9595), .A(n9164), .B(n9163), .ZN(n9166)
         );
  AOI21_X1 U10425 ( .B1(n9425), .B2(n9650), .A(n9166), .ZN(n9167) );
  OAI21_X1 U10426 ( .B1(n9429), .B2(n9364), .A(n9167), .ZN(P1_U3264) );
  XNOR2_X1 U10427 ( .A(n9168), .B(n9175), .ZN(n9434) );
  AOI21_X1 U10428 ( .B1(n9430), .B2(n9184), .A(n9169), .ZN(n9431) );
  AOI22_X1 U10429 ( .A1(n9647), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9170), .B2(
        n9645), .ZN(n9171) );
  OAI21_X1 U10430 ( .B1(n9172), .B2(n9595), .A(n9171), .ZN(n9181) );
  NAND2_X1 U10431 ( .A1(n9174), .A2(n9173), .ZN(n9176) );
  XNOR2_X1 U10432 ( .A(n9176), .B(n9175), .ZN(n9179) );
  AOI222_X1 U10433 ( .A1(n9640), .A2(n9179), .B1(n9178), .B2(n9309), .C1(n9177), .C2(n9311), .ZN(n9433) );
  NOR2_X1 U10434 ( .A1(n9433), .A2(n9647), .ZN(n9180) );
  AOI211_X1 U10435 ( .C1(n9431), .C2(n9631), .A(n9181), .B(n9180), .ZN(n9182)
         );
  OAI21_X1 U10436 ( .B1(n9434), .B2(n9364), .A(n9182), .ZN(P1_U3265) );
  XOR2_X1 U10437 ( .A(n9190), .B(n9183), .Z(n9439) );
  INV_X1 U10438 ( .A(n9205), .ZN(n9186) );
  INV_X1 U10439 ( .A(n9184), .ZN(n9185) );
  AOI21_X1 U10440 ( .B1(n9435), .B2(n9186), .A(n9185), .ZN(n9436) );
  AOI22_X1 U10441 ( .A1(n9647), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9187), .B2(
        n9645), .ZN(n9188) );
  OAI21_X1 U10442 ( .B1(n9189), .B2(n9595), .A(n9188), .ZN(n9196) );
  XNOR2_X1 U10443 ( .A(n9191), .B(n9190), .ZN(n9194) );
  AOI222_X1 U10444 ( .A1(n9640), .A2(n9194), .B1(n9193), .B2(n9309), .C1(n9192), .C2(n9311), .ZN(n9438) );
  NOR2_X1 U10445 ( .A1(n9438), .A2(n9647), .ZN(n9195) );
  AOI211_X1 U10446 ( .C1(n9436), .C2(n9631), .A(n9196), .B(n9195), .ZN(n9197)
         );
  OAI21_X1 U10447 ( .B1(n9439), .B2(n9364), .A(n9197), .ZN(P1_U3266) );
  XOR2_X1 U10448 ( .A(n9200), .B(n9198), .Z(n9444) );
  AOI22_X1 U10449 ( .A1(n9442), .A2(n9254), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9647), .ZN(n9211) );
  AOI21_X1 U10450 ( .B1(n9201), .B2(n9200), .A(n9199), .ZN(n9202) );
  OAI222_X1 U10451 ( .A1(n9635), .A2(n9204), .B1(n9638), .B2(n9203), .C1(n9370), .C2(n9202), .ZN(n9440) );
  AOI211_X1 U10452 ( .C1(n9442), .C2(n9219), .A(n9682), .B(n9205), .ZN(n9441)
         );
  INV_X1 U10453 ( .A(n9441), .ZN(n9208) );
  OAI22_X1 U10454 ( .A1(n9208), .A2(n9207), .B1(n9245), .B2(n9206), .ZN(n9209)
         );
  OAI21_X1 U10455 ( .B1(n9440), .B2(n9209), .A(n9650), .ZN(n9210) );
  OAI211_X1 U10456 ( .C1(n9444), .C2(n9364), .A(n9211), .B(n9210), .ZN(
        P1_U3267) );
  XNOR2_X1 U10457 ( .A(n9212), .B(n9216), .ZN(n9449) );
  NAND2_X1 U10458 ( .A1(n9214), .A2(n9213), .ZN(n9215) );
  XOR2_X1 U10459 ( .A(n9216), .B(n9215), .Z(n9217) );
  OAI222_X1 U10460 ( .A1(n9638), .A2(n9248), .B1(n9635), .B2(n9218), .C1(n9370), .C2(n9217), .ZN(n9445) );
  INV_X1 U10461 ( .A(n9229), .ZN(n9221) );
  INV_X1 U10462 ( .A(n9219), .ZN(n9220) );
  AOI211_X1 U10463 ( .C1(n9447), .C2(n9221), .A(n9682), .B(n9220), .ZN(n9446)
         );
  NAND2_X1 U10464 ( .A1(n9446), .A2(n9406), .ZN(n9224) );
  AOI22_X1 U10465 ( .A1(n9647), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9222), .B2(
        n9645), .ZN(n9223) );
  OAI211_X1 U10466 ( .C1(n9225), .C2(n9595), .A(n9224), .B(n9223), .ZN(n9226)
         );
  AOI21_X1 U10467 ( .B1(n9445), .B2(n9650), .A(n9226), .ZN(n9227) );
  OAI21_X1 U10468 ( .B1(n9449), .B2(n9364), .A(n9227), .ZN(P1_U3268) );
  XNOR2_X1 U10469 ( .A(n9228), .B(n9232), .ZN(n9454) );
  AOI21_X1 U10470 ( .B1(n9450), .B2(n9241), .A(n9229), .ZN(n9451) );
  AOI22_X1 U10471 ( .A1(n9647), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9230), .B2(
        n9645), .ZN(n9231) );
  OAI21_X1 U10472 ( .B1(n4439), .B2(n9595), .A(n9231), .ZN(n9238) );
  XNOR2_X1 U10473 ( .A(n9233), .B(n9232), .ZN(n9236) );
  AOI222_X1 U10474 ( .A1(n9640), .A2(n9236), .B1(n9235), .B2(n9309), .C1(n9234), .C2(n9311), .ZN(n9453) );
  NOR2_X1 U10475 ( .A1(n9453), .A2(n9647), .ZN(n9237) );
  AOI211_X1 U10476 ( .C1(n9451), .C2(n9631), .A(n9238), .B(n9237), .ZN(n9239)
         );
  OAI21_X1 U10477 ( .B1(n9454), .B2(n9364), .A(n9239), .ZN(P1_U3269) );
  INV_X1 U10478 ( .A(n9241), .ZN(n9242) );
  AOI211_X1 U10479 ( .C1(n9458), .C2(n4443), .A(n9682), .B(n9242), .ZN(n9457)
         );
  INV_X1 U10480 ( .A(n9243), .ZN(n9244) );
  NOR2_X1 U10481 ( .A1(n9245), .A2(n9244), .ZN(n9249) );
  XNOR2_X1 U10482 ( .A(n9246), .B(n9251), .ZN(n9247) );
  OAI222_X1 U10483 ( .A1(n9635), .A2(n9248), .B1(n9638), .B2(n9274), .C1(n9247), .C2(n9370), .ZN(n9456) );
  AOI211_X1 U10484 ( .C1(n9457), .C2(n9250), .A(n9249), .B(n9456), .ZN(n9257)
         );
  OR2_X1 U10485 ( .A1(n9252), .A2(n9251), .ZN(n9455) );
  NAND3_X1 U10486 ( .A1(n9455), .A2(n9253), .A3(n9323), .ZN(n9256) );
  AOI22_X1 U10487 ( .A1(n9458), .A2(n9254), .B1(n9647), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9255) );
  OAI211_X1 U10488 ( .C1(n9647), .C2(n9257), .A(n9256), .B(n9255), .ZN(
        P1_U3270) );
  XNOR2_X1 U10489 ( .A(n9258), .B(n9259), .ZN(n9465) );
  XNOR2_X1 U10490 ( .A(n9260), .B(n4586), .ZN(n9261) );
  OAI222_X1 U10491 ( .A1(n9638), .A2(n9263), .B1(n9635), .B2(n9262), .C1(n9261), .C2(n9370), .ZN(n9461) );
  AOI211_X1 U10492 ( .C1(n9463), .C2(n9276), .A(n9682), .B(n9240), .ZN(n9462)
         );
  NAND2_X1 U10493 ( .A1(n9462), .A2(n9406), .ZN(n9266) );
  AOI22_X1 U10494 ( .A1(n9647), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9264), .B2(
        n9645), .ZN(n9265) );
  OAI211_X1 U10495 ( .C1(n9267), .C2(n9595), .A(n9266), .B(n9265), .ZN(n9268)
         );
  AOI21_X1 U10496 ( .B1(n9461), .B2(n9650), .A(n9268), .ZN(n9269) );
  OAI21_X1 U10497 ( .B1(n9465), .B2(n9364), .A(n9269), .ZN(P1_U3271) );
  XNOR2_X1 U10498 ( .A(n9270), .B(n9272), .ZN(n9470) );
  XOR2_X1 U10499 ( .A(n9272), .B(n9271), .Z(n9273) );
  OAI222_X1 U10500 ( .A1(n9638), .A2(n9275), .B1(n9635), .B2(n9274), .C1(n9273), .C2(n9370), .ZN(n9466) );
  INV_X1 U10501 ( .A(n9287), .ZN(n9278) );
  INV_X1 U10502 ( .A(n9276), .ZN(n9277) );
  AOI211_X1 U10503 ( .C1(n9468), .C2(n9278), .A(n9682), .B(n9277), .ZN(n9467)
         );
  NAND2_X1 U10504 ( .A1(n9467), .A2(n9406), .ZN(n9281) );
  AOI22_X1 U10505 ( .A1(n9647), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9279), .B2(
        n9645), .ZN(n9280) );
  OAI211_X1 U10506 ( .C1(n9282), .C2(n9595), .A(n9281), .B(n9280), .ZN(n9283)
         );
  AOI21_X1 U10507 ( .B1(n9466), .B2(n9650), .A(n9283), .ZN(n9284) );
  OAI21_X1 U10508 ( .B1(n9470), .B2(n9364), .A(n9284), .ZN(P1_U3272) );
  XNOR2_X1 U10509 ( .A(n9285), .B(n9286), .ZN(n9475) );
  INV_X1 U10510 ( .A(n9304), .ZN(n9288) );
  AOI21_X1 U10511 ( .B1(n9471), .B2(n9288), .A(n9287), .ZN(n9472) );
  AOI22_X1 U10512 ( .A1(n9647), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9289), .B2(
        n9645), .ZN(n9290) );
  OAI21_X1 U10513 ( .B1(n9291), .B2(n9595), .A(n9290), .ZN(n9300) );
  INV_X1 U10514 ( .A(n9292), .ZN(n9293) );
  NOR2_X1 U10515 ( .A1(n4289), .A2(n9293), .ZN(n9295) );
  XNOR2_X1 U10516 ( .A(n9295), .B(n9294), .ZN(n9298) );
  AOI222_X1 U10517 ( .A1(n9640), .A2(n9298), .B1(n9297), .B2(n9309), .C1(n9296), .C2(n9311), .ZN(n9474) );
  NOR2_X1 U10518 ( .A1(n9474), .A2(n9647), .ZN(n9299) );
  AOI211_X1 U10519 ( .C1(n9472), .C2(n9631), .A(n9300), .B(n9299), .ZN(n9301)
         );
  OAI21_X1 U10520 ( .B1(n9364), .B2(n9475), .A(n9301), .ZN(P1_U3273) );
  XNOR2_X1 U10521 ( .A(n9303), .B(n9302), .ZN(n9480) );
  AOI21_X1 U10522 ( .B1(n9476), .B2(n9324), .A(n9304), .ZN(n9477) );
  AOI22_X1 U10523 ( .A1(n9647), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9305), .B2(
        n9645), .ZN(n9306) );
  OAI21_X1 U10524 ( .B1(n9069), .B2(n9595), .A(n9306), .ZN(n9315) );
  XNOR2_X1 U10525 ( .A(n9307), .B(n9308), .ZN(n9313) );
  AOI222_X1 U10526 ( .A1(n9640), .A2(n9313), .B1(n9312), .B2(n9311), .C1(n9310), .C2(n9309), .ZN(n9479) );
  NOR2_X1 U10527 ( .A1(n9479), .A2(n9647), .ZN(n9314) );
  AOI211_X1 U10528 ( .C1(n9477), .C2(n9631), .A(n9315), .B(n9314), .ZN(n9316)
         );
  OAI21_X1 U10529 ( .B1(n9364), .B2(n9480), .A(n9316), .ZN(P1_U3274) );
  XOR2_X1 U10530 ( .A(n9319), .B(n9317), .Z(n9318) );
  OAI222_X1 U10531 ( .A1(n9638), .A2(n9355), .B1(n9635), .B2(n9068), .C1(n9318), .C2(n9370), .ZN(n9481) );
  INV_X1 U10532 ( .A(n9481), .ZN(n9331) );
  OR2_X1 U10533 ( .A1(n9320), .A2(n9319), .ZN(n9484) );
  NAND3_X1 U10534 ( .A1(n9484), .A2(n9322), .A3(n9323), .ZN(n9330) );
  INV_X1 U10535 ( .A(n9324), .ZN(n9325) );
  AOI211_X1 U10536 ( .C1(n9483), .C2(n9342), .A(n9682), .B(n9325), .ZN(n9482)
         );
  AOI22_X1 U10537 ( .A1(n9647), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9326), .B2(
        n9645), .ZN(n9327) );
  OAI21_X1 U10538 ( .B1(n4445), .B2(n9595), .A(n9327), .ZN(n9328) );
  AOI21_X1 U10539 ( .B1(n9482), .B2(n9406), .A(n9328), .ZN(n9329) );
  OAI211_X1 U10540 ( .C1(n9647), .C2(n9331), .A(n9330), .B(n9329), .ZN(
        P1_U3275) );
  XNOR2_X1 U10541 ( .A(n9332), .B(n4367), .ZN(n9333) );
  INV_X1 U10542 ( .A(n9333), .ZN(n9490) );
  NAND2_X1 U10543 ( .A1(n9333), .A2(n9376), .ZN(n9340) );
  XNOR2_X1 U10544 ( .A(n9335), .B(n9334), .ZN(n9338) );
  OAI22_X1 U10545 ( .A1(n9638), .A2(n9373), .B1(n9336), .B2(n9635), .ZN(n9337)
         );
  AOI21_X1 U10546 ( .B1(n9338), .B2(n9640), .A(n9337), .ZN(n9339) );
  NAND2_X1 U10547 ( .A1(n9340), .A2(n9339), .ZN(n9492) );
  NAND2_X1 U10548 ( .A1(n9492), .A2(n9650), .ZN(n9348) );
  OR2_X1 U10549 ( .A1(n9356), .A2(n9345), .ZN(n9341) );
  AND2_X1 U10550 ( .A1(n9342), .A2(n9341), .ZN(n9488) );
  AOI22_X1 U10551 ( .A1(n9647), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9343), .B2(
        n9645), .ZN(n9344) );
  OAI21_X1 U10552 ( .B1(n9345), .B2(n9595), .A(n9344), .ZN(n9346) );
  AOI21_X1 U10553 ( .B1(n9488), .B2(n9631), .A(n9346), .ZN(n9347) );
  OAI211_X1 U10554 ( .C1(n9490), .C2(n9585), .A(n9348), .B(n9347), .ZN(
        P1_U3276) );
  INV_X1 U10555 ( .A(n9349), .ZN(n9350) );
  AOI21_X1 U10556 ( .B1(n9352), .B2(n9351), .A(n9350), .ZN(n9498) );
  XNOR2_X1 U10557 ( .A(n9353), .B(n9352), .ZN(n9354) );
  OAI222_X1 U10558 ( .A1(n9638), .A2(n9390), .B1(n9635), .B2(n9355), .C1(n9354), .C2(n9370), .ZN(n9493) );
  INV_X1 U10559 ( .A(n9377), .ZN(n9357) );
  AOI211_X1 U10560 ( .C1(n9495), .C2(n9357), .A(n9682), .B(n9356), .ZN(n9494)
         );
  NAND2_X1 U10561 ( .A1(n9494), .A2(n9406), .ZN(n9360) );
  AOI22_X1 U10562 ( .A1(n9647), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9358), .B2(
        n9645), .ZN(n9359) );
  OAI211_X1 U10563 ( .C1(n9361), .C2(n9595), .A(n9360), .B(n9359), .ZN(n9362)
         );
  AOI21_X1 U10564 ( .B1(n9493), .B2(n9650), .A(n9362), .ZN(n9363) );
  OAI21_X1 U10565 ( .B1(n9498), .B2(n9364), .A(n9363), .ZN(P1_U3277) );
  XNOR2_X1 U10566 ( .A(n9367), .B(n9366), .ZN(n9381) );
  NAND2_X1 U10567 ( .A1(n9369), .A2(n9368), .ZN(n9371) );
  AOI21_X1 U10568 ( .B1(n9372), .B2(n9371), .A(n9370), .ZN(n9375) );
  OAI22_X1 U10569 ( .A1(n9638), .A2(n9589), .B1(n9373), .B2(n9635), .ZN(n9374)
         );
  AOI211_X1 U10570 ( .C1(n9381), .C2(n9376), .A(n9375), .B(n9374), .ZN(n9503)
         );
  AOI21_X1 U10571 ( .B1(n9499), .B2(n9399), .A(n9377), .ZN(n9501) );
  AOI22_X1 U10572 ( .A1(n9647), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9378), .B2(
        n9645), .ZN(n9379) );
  OAI21_X1 U10573 ( .B1(n9380), .B2(n9595), .A(n9379), .ZN(n9383) );
  INV_X1 U10574 ( .A(n9381), .ZN(n9504) );
  NOR2_X1 U10575 ( .A1(n9504), .A2(n9585), .ZN(n9382) );
  AOI211_X1 U10576 ( .C1(n9501), .C2(n9631), .A(n9383), .B(n9382), .ZN(n9384)
         );
  OAI21_X1 U10577 ( .B1(n9647), .B2(n9503), .A(n9384), .ZN(P1_U3278) );
  INV_X1 U10578 ( .A(n9385), .ZN(n9386) );
  AOI21_X1 U10579 ( .B1(n9588), .B2(n9387), .A(n9386), .ZN(n9389) );
  XNOR2_X1 U10580 ( .A(n9389), .B(n9388), .ZN(n9398) );
  OAI22_X1 U10581 ( .A1(n9638), .A2(n9391), .B1(n9390), .B2(n9635), .ZN(n9397)
         );
  OR2_X1 U10582 ( .A1(n9393), .A2(n9392), .ZN(n9394) );
  NAND2_X1 U10583 ( .A1(n9395), .A2(n9394), .ZN(n9509) );
  NOR2_X1 U10584 ( .A1(n9509), .A2(n9643), .ZN(n9396) );
  AOI211_X1 U10585 ( .C1(n9640), .C2(n9398), .A(n9397), .B(n9396), .ZN(n9508)
         );
  INV_X1 U10586 ( .A(n9399), .ZN(n9400) );
  AOI211_X1 U10587 ( .C1(n9506), .C2(n9583), .A(n9682), .B(n9400), .ZN(n9505)
         );
  AOI22_X1 U10588 ( .A1(n9647), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9401), .B2(
        n9645), .ZN(n9402) );
  OAI21_X1 U10589 ( .B1(n9403), .B2(n9595), .A(n9402), .ZN(n9405) );
  NOR2_X1 U10590 ( .A1(n9509), .A2(n9585), .ZN(n9404) );
  AOI211_X1 U10591 ( .C1(n9505), .C2(n9406), .A(n9405), .B(n9404), .ZN(n9407)
         );
  OAI21_X1 U10592 ( .B1(n9508), .B2(n9647), .A(n9407), .ZN(P1_U3279) );
  NAND2_X1 U10593 ( .A1(n4651), .A2(n9568), .ZN(n9408) );
  OAI211_X1 U10594 ( .C1(n9409), .C2(n9682), .A(n9408), .B(n9412), .ZN(n9511)
         );
  MUX2_X1 U10595 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9511), .S(n9697), .Z(
        P1_U3554) );
  NAND2_X1 U10596 ( .A1(n9410), .A2(n9568), .ZN(n9411) );
  OAI211_X1 U10597 ( .C1(n9413), .C2(n9682), .A(n9412), .B(n9411), .ZN(n9512)
         );
  MUX2_X1 U10598 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9512), .S(n9697), .Z(
        P1_U3553) );
  NAND2_X1 U10599 ( .A1(n9414), .A2(n9678), .ZN(n9419) );
  NAND2_X1 U10600 ( .A1(n9419), .A2(n9418), .ZN(n9513) );
  MUX2_X1 U10601 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9513), .S(n9697), .Z(
        P1_U3552) );
  NAND2_X1 U10602 ( .A1(n9420), .A2(n9678), .ZN(n9424) );
  MUX2_X1 U10603 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9514), .S(n9697), .Z(
        P1_U3551) );
  AOI211_X1 U10604 ( .C1(n9568), .C2(n9427), .A(n9426), .B(n9425), .ZN(n9428)
         );
  OAI21_X1 U10605 ( .B1(n9429), .B2(n9497), .A(n9428), .ZN(n9515) );
  MUX2_X1 U10606 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9515), .S(n9697), .Z(
        P1_U3550) );
  AOI22_X1 U10607 ( .A1(n9431), .A2(n9500), .B1(n9568), .B2(n9430), .ZN(n9432)
         );
  OAI211_X1 U10608 ( .C1(n9434), .C2(n9497), .A(n9433), .B(n9432), .ZN(n9516)
         );
  MUX2_X1 U10609 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9516), .S(n9697), .Z(
        P1_U3549) );
  AOI22_X1 U10610 ( .A1(n9436), .A2(n9500), .B1(n9568), .B2(n9435), .ZN(n9437)
         );
  OAI211_X1 U10611 ( .C1(n9439), .C2(n9497), .A(n9438), .B(n9437), .ZN(n9517)
         );
  MUX2_X1 U10612 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9517), .S(n9697), .Z(
        P1_U3548) );
  AOI211_X1 U10613 ( .C1(n9568), .C2(n9442), .A(n9441), .B(n9440), .ZN(n9443)
         );
  OAI21_X1 U10614 ( .B1(n9444), .B2(n9497), .A(n9443), .ZN(n9518) );
  MUX2_X1 U10615 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9518), .S(n9697), .Z(
        P1_U3547) );
  AOI211_X1 U10616 ( .C1(n9568), .C2(n9447), .A(n9446), .B(n9445), .ZN(n9448)
         );
  OAI21_X1 U10617 ( .B1(n9449), .B2(n9497), .A(n9448), .ZN(n9519) );
  MUX2_X1 U10618 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9519), .S(n9697), .Z(
        P1_U3546) );
  AOI22_X1 U10619 ( .A1(n9451), .A2(n9500), .B1(n9568), .B2(n9450), .ZN(n9452)
         );
  OAI211_X1 U10620 ( .C1(n9454), .C2(n9497), .A(n9453), .B(n9452), .ZN(n9520)
         );
  MUX2_X1 U10621 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9520), .S(n9697), .Z(
        P1_U3545) );
  NAND3_X1 U10622 ( .A1(n9455), .A2(n9253), .A3(n9678), .ZN(n9460) );
  AOI211_X1 U10623 ( .C1(n9568), .C2(n9458), .A(n9457), .B(n9456), .ZN(n9459)
         );
  NAND2_X1 U10624 ( .A1(n9460), .A2(n9459), .ZN(n9521) );
  MUX2_X1 U10625 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9521), .S(n9697), .Z(
        P1_U3544) );
  AOI211_X1 U10626 ( .C1(n9568), .C2(n9463), .A(n9462), .B(n9461), .ZN(n9464)
         );
  OAI21_X1 U10627 ( .B1(n9465), .B2(n9497), .A(n9464), .ZN(n9522) );
  MUX2_X1 U10628 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9522), .S(n9697), .Z(
        P1_U3543) );
  AOI211_X1 U10629 ( .C1(n9568), .C2(n9468), .A(n9467), .B(n9466), .ZN(n9469)
         );
  OAI21_X1 U10630 ( .B1(n9470), .B2(n9497), .A(n9469), .ZN(n9523) );
  MUX2_X1 U10631 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9523), .S(n9697), .Z(
        P1_U3542) );
  AOI22_X1 U10632 ( .A1(n9472), .A2(n9500), .B1(n9568), .B2(n9471), .ZN(n9473)
         );
  OAI211_X1 U10633 ( .C1(n9475), .C2(n9497), .A(n9474), .B(n9473), .ZN(n9524)
         );
  MUX2_X1 U10634 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9524), .S(n9697), .Z(
        P1_U3541) );
  AOI22_X1 U10635 ( .A1(n9477), .A2(n9500), .B1(n9568), .B2(n9476), .ZN(n9478)
         );
  OAI211_X1 U10636 ( .C1(n9480), .C2(n9497), .A(n9479), .B(n9478), .ZN(n9525)
         );
  MUX2_X1 U10637 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9525), .S(n9697), .Z(
        P1_U3540) );
  AOI211_X1 U10638 ( .C1(n9568), .C2(n9483), .A(n9482), .B(n9481), .ZN(n9486)
         );
  NAND3_X1 U10639 ( .A1(n9484), .A2(n9322), .A3(n9678), .ZN(n9485) );
  NAND2_X1 U10640 ( .A1(n9486), .A2(n9485), .ZN(n9526) );
  MUX2_X1 U10641 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9526), .S(n9697), .Z(
        P1_U3539) );
  AOI22_X1 U10642 ( .A1(n9488), .A2(n9500), .B1(n9568), .B2(n9487), .ZN(n9489)
         );
  OAI21_X1 U10643 ( .B1(n9490), .B2(n9510), .A(n9489), .ZN(n9491) );
  MUX2_X1 U10644 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9527), .S(n9697), .Z(
        P1_U3538) );
  AOI211_X1 U10645 ( .C1(n9568), .C2(n9495), .A(n9494), .B(n9493), .ZN(n9496)
         );
  OAI21_X1 U10646 ( .B1(n9498), .B2(n9497), .A(n9496), .ZN(n9528) );
  MUX2_X1 U10647 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9528), .S(n9697), .Z(
        P1_U3537) );
  AOI22_X1 U10648 ( .A1(n9501), .A2(n9500), .B1(n9568), .B2(n9499), .ZN(n9502)
         );
  OAI211_X1 U10649 ( .C1(n9510), .C2(n9504), .A(n9503), .B(n9502), .ZN(n9529)
         );
  MUX2_X1 U10650 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9529), .S(n9697), .Z(
        P1_U3536) );
  AOI21_X1 U10651 ( .B1(n9568), .B2(n9506), .A(n9505), .ZN(n9507) );
  OAI211_X1 U10652 ( .C1(n9510), .C2(n9509), .A(n9508), .B(n9507), .ZN(n9531)
         );
  MUX2_X1 U10653 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9531), .S(n9697), .Z(
        P1_U3535) );
  MUX2_X1 U10654 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9511), .S(n9530), .Z(
        P1_U3522) );
  MUX2_X1 U10655 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9512), .S(n9530), .Z(
        P1_U3521) );
  MUX2_X1 U10656 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9513), .S(n9530), .Z(
        P1_U3520) );
  MUX2_X1 U10657 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9514), .S(n9530), .Z(
        P1_U3519) );
  MUX2_X1 U10658 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9515), .S(n9530), .Z(
        P1_U3518) );
  MUX2_X1 U10659 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9516), .S(n9530), .Z(
        P1_U3517) );
  MUX2_X1 U10660 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9517), .S(n9530), .Z(
        P1_U3516) );
  MUX2_X1 U10661 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9518), .S(n9530), .Z(
        P1_U3515) );
  MUX2_X1 U10662 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9519), .S(n9530), .Z(
        P1_U3514) );
  MUX2_X1 U10663 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9520), .S(n9530), .Z(
        P1_U3513) );
  MUX2_X1 U10664 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9521), .S(n9530), .Z(
        P1_U3512) );
  MUX2_X1 U10665 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9522), .S(n9530), .Z(
        P1_U3511) );
  MUX2_X1 U10666 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9523), .S(n9530), .Z(
        P1_U3510) );
  MUX2_X1 U10667 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9524), .S(n9530), .Z(
        P1_U3508) );
  MUX2_X1 U10668 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9525), .S(n9530), .Z(
        P1_U3505) );
  MUX2_X1 U10669 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9526), .S(n9530), .Z(
        P1_U3502) );
  MUX2_X1 U10670 ( .A(n9527), .B(P1_REG0_REG_15__SCAN_IN), .S(n9688), .Z(
        P1_U3499) );
  MUX2_X1 U10671 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9528), .S(n9530), .Z(
        P1_U3496) );
  MUX2_X1 U10672 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9529), .S(n9530), .Z(
        P1_U3493) );
  MUX2_X1 U10673 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9531), .S(n9530), .Z(
        P1_U3490) );
  MUX2_X1 U10674 ( .A(P1_D_REG_1__SCAN_IN), .B(n9532), .S(n9654), .Z(P1_U3441)
         );
  MUX2_X1 U10675 ( .A(P1_D_REG_0__SCAN_IN), .B(n9533), .S(n9654), .Z(P1_U3440)
         );
  INV_X1 U10676 ( .A(n9534), .ZN(n9539) );
  NOR4_X1 U10677 ( .A1(n9536), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9535), .ZN(n9537) );
  AOI21_X1 U10678 ( .B1(n9549), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9537), .ZN(
        n9538) );
  OAI21_X1 U10679 ( .B1(n9539), .B2(n9552), .A(n9538), .ZN(P1_U3322) );
  AOI22_X1 U10680 ( .A1(n9540), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9549), .ZN(n9541) );
  OAI21_X1 U10681 ( .B1(n9542), .B2(n9552), .A(n9541), .ZN(P1_U3323) );
  AOI22_X1 U10682 ( .A1(n9543), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9549), .ZN(n9544) );
  OAI21_X1 U10683 ( .B1(n9545), .B2(n9552), .A(n9544), .ZN(P1_U3324) );
  AOI21_X1 U10684 ( .B1(n9549), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n9546), .ZN(
        n9547) );
  OAI21_X1 U10685 ( .B1(n9548), .B2(n9552), .A(n9547), .ZN(P1_U3325) );
  NAND2_X1 U10686 ( .A1(n9549), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9550) );
  OAI211_X1 U10687 ( .C1(n9553), .C2(n9552), .A(n9551), .B(n9550), .ZN(
        P1_U3326) );
  MUX2_X1 U10688 ( .A(n9554), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10689 ( .A1(n9715), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9566) );
  AOI211_X1 U10690 ( .C1(n9557), .C2(n9556), .A(n9555), .B(n9718), .ZN(n9558)
         );
  AOI21_X1 U10691 ( .B1(n9560), .B2(n9559), .A(n9558), .ZN(n9565) );
  OAI211_X1 U10692 ( .C1(n9563), .C2(n9562), .A(n9714), .B(n9561), .ZN(n9564)
         );
  NAND3_X1 U10693 ( .A1(n9566), .A2(n9565), .A3(n9564), .ZN(P2_U3247) );
  INV_X1 U10694 ( .A(n9567), .ZN(n9573) );
  OAI21_X1 U10695 ( .B1(n9570), .B2(n9680), .A(n9569), .ZN(n9572) );
  AOI211_X1 U10696 ( .C1(n9687), .C2(n9573), .A(n9572), .B(n9571), .ZN(n9576)
         );
  INV_X1 U10697 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9574) );
  AOI22_X1 U10698 ( .A1(n9530), .A2(n9576), .B1(n9574), .B2(n9688), .ZN(
        P1_U3484) );
  AOI22_X1 U10699 ( .A1(n9697), .A2(n9576), .B1(n9575), .B2(n9694), .ZN(
        P1_U3533) );
  NAND2_X1 U10700 ( .A1(n9578), .A2(n9579), .ZN(n9580) );
  NAND2_X1 U10701 ( .A1(n9577), .A2(n9580), .ZN(n9599) );
  OR2_X1 U10702 ( .A1(n9581), .A2(n9600), .ZN(n9582) );
  NAND2_X1 U10703 ( .A1(n9583), .A2(n9582), .ZN(n9601) );
  OAI22_X1 U10704 ( .A1(n9599), .A2(n9585), .B1(n9584), .B2(n9601), .ZN(n9586)
         );
  INV_X1 U10705 ( .A(n9586), .ZN(n9598) );
  XNOR2_X1 U10706 ( .A(n9588), .B(n9587), .ZN(n9591) );
  OAI22_X1 U10707 ( .A1(n9638), .A2(n9636), .B1(n9589), .B2(n9635), .ZN(n9590)
         );
  AOI21_X1 U10708 ( .B1(n9591), .B2(n9640), .A(n9590), .ZN(n9592) );
  OAI21_X1 U10709 ( .B1(n9599), .B2(n9643), .A(n9592), .ZN(n9602) );
  AOI22_X1 U10710 ( .A1(n9647), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9593), .B2(
        n9645), .ZN(n9594) );
  OAI21_X1 U10711 ( .B1(n9600), .B2(n9595), .A(n9594), .ZN(n9596) );
  AOI21_X1 U10712 ( .B1(n9602), .B2(n9650), .A(n9596), .ZN(n9597) );
  NAND2_X1 U10713 ( .A1(n9598), .A2(n9597), .ZN(P1_U3280) );
  INV_X1 U10714 ( .A(n9599), .ZN(n9604) );
  OAI22_X1 U10715 ( .A1(n9601), .A2(n9682), .B1(n9600), .B2(n9680), .ZN(n9603)
         );
  AOI211_X1 U10716 ( .C1(n9687), .C2(n9604), .A(n9603), .B(n9602), .ZN(n9607)
         );
  AOI22_X1 U10717 ( .A1(n9697), .A2(n9607), .B1(n9605), .B2(n9694), .ZN(
        P1_U3534) );
  INV_X1 U10718 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9606) );
  AOI22_X1 U10719 ( .A1(n9530), .A2(n9607), .B1(n9606), .B2(n9688), .ZN(
        P1_U3487) );
  XOR2_X1 U10720 ( .A(n9608), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  XNOR2_X1 U10721 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  AOI22_X1 U10722 ( .A1(n9611), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n9610), .B2(
        n9609), .ZN(n9627) );
  INV_X1 U10723 ( .A(n9612), .ZN(n9618) );
  NOR3_X1 U10724 ( .A1(n9615), .A2(n9614), .A3(n9613), .ZN(n9617) );
  OAI21_X1 U10725 ( .B1(n9618), .B2(n9617), .A(n9616), .ZN(n9625) );
  NAND2_X1 U10726 ( .A1(n9620), .A2(n9619), .ZN(n9621) );
  NAND3_X1 U10727 ( .A1(n9623), .A2(n9622), .A3(n9621), .ZN(n9624) );
  NAND4_X1 U10728 ( .A1(n9627), .A2(n9626), .A3(n9625), .A4(n9624), .ZN(
        P1_U3246) );
  XNOR2_X1 U10729 ( .A(n9628), .B(n9633), .ZN(n9644) );
  INV_X1 U10730 ( .A(n9644), .ZN(n9686) );
  OAI21_X1 U10731 ( .B1(n4336), .B2(n9681), .A(n9629), .ZN(n9683) );
  INV_X1 U10732 ( .A(n9683), .ZN(n9630) );
  AOI22_X1 U10733 ( .A1(n9686), .A2(n9632), .B1(n9631), .B2(n9630), .ZN(n9652)
         );
  XNOR2_X1 U10734 ( .A(n9634), .B(n9633), .ZN(n9641) );
  OAI22_X1 U10735 ( .A1(n9638), .A2(n9637), .B1(n9636), .B2(n9635), .ZN(n9639)
         );
  AOI21_X1 U10736 ( .B1(n9641), .B2(n9640), .A(n9639), .ZN(n9642) );
  OAI21_X1 U10737 ( .B1(n9644), .B2(n9643), .A(n9642), .ZN(n9684) );
  AOI22_X1 U10738 ( .A1(n9647), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n9646), .B2(
        n9645), .ZN(n9648) );
  OAI21_X1 U10739 ( .B1(n9681), .B2(n9595), .A(n9648), .ZN(n9649) );
  AOI21_X1 U10740 ( .B1(n9684), .B2(n9650), .A(n9649), .ZN(n9651) );
  NAND2_X1 U10741 ( .A1(n9652), .A2(n9651), .ZN(P1_U3282) );
  AND2_X1 U10742 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9660), .ZN(P1_U3292) );
  NOR2_X1 U10743 ( .A1(n9659), .A2(n9655), .ZN(P1_U3293) );
  AND2_X1 U10744 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9660), .ZN(P1_U3294) );
  AND2_X1 U10745 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9660), .ZN(P1_U3295) );
  NOR2_X1 U10746 ( .A1(n9659), .A2(n9656), .ZN(P1_U3296) );
  AND2_X1 U10747 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9660), .ZN(P1_U3297) );
  AND2_X1 U10748 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9660), .ZN(P1_U3298) );
  AND2_X1 U10749 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9660), .ZN(P1_U3299) );
  AND2_X1 U10750 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9660), .ZN(P1_U3300) );
  NOR2_X1 U10751 ( .A1(n9659), .A2(n9657), .ZN(P1_U3301) );
  AND2_X1 U10752 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9660), .ZN(P1_U3302) );
  AND2_X1 U10753 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9660), .ZN(P1_U3303) );
  AND2_X1 U10754 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9660), .ZN(P1_U3304) );
  AND2_X1 U10755 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9660), .ZN(P1_U3305) );
  AND2_X1 U10756 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9660), .ZN(P1_U3306) );
  AND2_X1 U10757 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9660), .ZN(P1_U3307) );
  AND2_X1 U10758 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9660), .ZN(P1_U3308) );
  AND2_X1 U10759 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9660), .ZN(P1_U3309) );
  AND2_X1 U10760 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9660), .ZN(P1_U3310) );
  AND2_X1 U10761 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9660), .ZN(P1_U3311) );
  AND2_X1 U10762 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9660), .ZN(P1_U3312) );
  AND2_X1 U10763 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9660), .ZN(P1_U3313) );
  AND2_X1 U10764 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9660), .ZN(P1_U3314) );
  AND2_X1 U10765 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9660), .ZN(P1_U3315) );
  AND2_X1 U10766 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9660), .ZN(P1_U3316) );
  AND2_X1 U10767 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9660), .ZN(P1_U3317) );
  AND2_X1 U10768 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9660), .ZN(P1_U3318) );
  NOR2_X1 U10769 ( .A1(n9659), .A2(n9658), .ZN(P1_U3319) );
  AND2_X1 U10770 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9660), .ZN(P1_U3320) );
  AND2_X1 U10771 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9660), .ZN(P1_U3321) );
  NAND2_X1 U10772 ( .A1(n9661), .A2(n9687), .ZN(n9663) );
  OAI211_X1 U10773 ( .C1(n9664), .C2(n9680), .A(n9663), .B(n9662), .ZN(n9665)
         );
  NOR2_X1 U10774 ( .A1(n9666), .A2(n9665), .ZN(n9690) );
  INV_X1 U10775 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9667) );
  AOI22_X1 U10776 ( .A1(n9530), .A2(n9690), .B1(n9667), .B2(n9688), .ZN(
        P1_U3457) );
  OAI22_X1 U10777 ( .A1(n9668), .A2(n9682), .B1(n5706), .B2(n9680), .ZN(n9670)
         );
  AOI211_X1 U10778 ( .C1(n9687), .C2(n9671), .A(n9670), .B(n9669), .ZN(n9691)
         );
  INV_X1 U10779 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9672) );
  AOI22_X1 U10780 ( .A1(n9530), .A2(n9691), .B1(n9672), .B2(n9688), .ZN(
        P1_U3463) );
  OAI211_X1 U10781 ( .C1(n9675), .C2(n9680), .A(n9674), .B(n9673), .ZN(n9676)
         );
  AOI21_X1 U10782 ( .B1(n9678), .B2(n9677), .A(n9676), .ZN(n9693) );
  INV_X1 U10783 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9679) );
  AOI22_X1 U10784 ( .A1(n9530), .A2(n9693), .B1(n9679), .B2(n9688), .ZN(
        P1_U3475) );
  OAI22_X1 U10785 ( .A1(n9683), .A2(n9682), .B1(n9681), .B2(n9680), .ZN(n9685)
         );
  AOI211_X1 U10786 ( .C1(n9687), .C2(n9686), .A(n9685), .B(n9684), .ZN(n9696)
         );
  INV_X1 U10787 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9689) );
  AOI22_X1 U10788 ( .A1(n9530), .A2(n9696), .B1(n9689), .B2(n9688), .ZN(
        P1_U3481) );
  AOI22_X1 U10789 ( .A1(n9697), .A2(n9690), .B1(n5997), .B2(n9694), .ZN(
        P1_U3524) );
  AOI22_X1 U10790 ( .A1(n9697), .A2(n9691), .B1(n6000), .B2(n9694), .ZN(
        P1_U3526) );
  AOI22_X1 U10791 ( .A1(n9697), .A2(n9693), .B1(n9692), .B2(n9694), .ZN(
        P1_U3530) );
  AOI22_X1 U10792 ( .A1(n9697), .A2(n9696), .B1(n9695), .B2(n9694), .ZN(
        P1_U3532) );
  OAI21_X1 U10793 ( .B1(n9700), .B2(n9699), .A(n9698), .ZN(n9708) );
  NOR2_X1 U10794 ( .A1(n9701), .A2(n6760), .ZN(n9707) );
  OAI22_X1 U10795 ( .A1(n9705), .A2(n9704), .B1(n9703), .B2(n9702), .ZN(n9706)
         );
  AOI211_X1 U10796 ( .C1(n9709), .C2(n9708), .A(n9707), .B(n9706), .ZN(n9710)
         );
  OAI21_X1 U10797 ( .B1(n9712), .B2(n9711), .A(n9710), .ZN(P2_U3224) );
  AOI22_X1 U10798 ( .A1(n9714), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9713), .ZN(n9723) );
  AOI22_X1 U10799 ( .A1(n9715), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9722) );
  NOR2_X1 U10800 ( .A1(n9716), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9720) );
  OAI21_X1 U10801 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n9718), .A(n9717), .ZN(
        n9719) );
  OAI21_X1 U10802 ( .B1(n9720), .B2(n9719), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9721) );
  OAI211_X1 U10803 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9723), .A(n9722), .B(
        n9721), .ZN(P2_U3245) );
  NAND2_X1 U10804 ( .A1(n9725), .A2(n9737), .ZN(n9726) );
  NAND2_X1 U10805 ( .A1(n9727), .A2(n9726), .ZN(n9741) );
  INV_X1 U10806 ( .A(n9741), .ZN(n9877) );
  INV_X1 U10807 ( .A(n9728), .ZN(n9731) );
  INV_X1 U10808 ( .A(n9729), .ZN(n9730) );
  OAI21_X1 U10809 ( .B1(n9873), .B2(n9731), .A(n9730), .ZN(n9874) );
  INV_X1 U10810 ( .A(n9874), .ZN(n9732) );
  AOI22_X1 U10811 ( .A1(n9877), .A2(n9734), .B1(n9733), .B2(n9732), .ZN(n9746)
         );
  AOI22_X1 U10812 ( .A1(n9762), .A2(n9765), .B1(n9735), .B2(n9764), .ZN(n9740)
         );
  OAI211_X1 U10813 ( .C1(n9738), .C2(n9737), .A(n9736), .B(n9769), .ZN(n9739)
         );
  OAI211_X1 U10814 ( .C1(n9741), .C2(n9757), .A(n9740), .B(n9739), .ZN(n9875)
         );
  AOI22_X1 U10815 ( .A1(n9775), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n9742), .B2(
        n9773), .ZN(n9743) );
  OAI21_X1 U10816 ( .B1(n9873), .B2(n9777), .A(n9743), .ZN(n9744) );
  AOI21_X1 U10817 ( .B1(n9875), .B2(n9779), .A(n9744), .ZN(n9745) );
  NAND2_X1 U10818 ( .A1(n9746), .A2(n9745), .ZN(P2_U3286) );
  NAND2_X1 U10819 ( .A1(n9748), .A2(n9749), .ZN(n9750) );
  NAND2_X1 U10820 ( .A1(n9747), .A2(n9750), .ZN(n9857) );
  OR2_X1 U10821 ( .A1(n9751), .A2(n9858), .ZN(n9752) );
  NAND2_X1 U10822 ( .A1(n9753), .A2(n9752), .ZN(n9859) );
  OAI22_X1 U10823 ( .A1(n9857), .A2(n9755), .B1(n9754), .B2(n9859), .ZN(n9756)
         );
  INV_X1 U10824 ( .A(n9756), .ZN(n9781) );
  OR2_X1 U10825 ( .A1(n9857), .A2(n9757), .ZN(n9772) );
  NAND2_X1 U10826 ( .A1(n9759), .A2(n9758), .ZN(n9760) );
  NAND2_X1 U10827 ( .A1(n9761), .A2(n9760), .ZN(n9770) );
  NAND2_X1 U10828 ( .A1(n9763), .A2(n9762), .ZN(n9767) );
  NAND2_X1 U10829 ( .A1(n9765), .A2(n9764), .ZN(n9766) );
  NAND2_X1 U10830 ( .A1(n9767), .A2(n9766), .ZN(n9768) );
  AOI21_X1 U10831 ( .B1(n9770), .B2(n9769), .A(n9768), .ZN(n9771) );
  NAND2_X1 U10832 ( .A1(n9772), .A2(n9771), .ZN(n9862) );
  AOI22_X1 U10833 ( .A1(n9775), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n9774), .B2(
        n9773), .ZN(n9776) );
  OAI21_X1 U10834 ( .B1(n9858), .B2(n9777), .A(n9776), .ZN(n9778) );
  AOI21_X1 U10835 ( .B1(n9862), .B2(n9779), .A(n9778), .ZN(n9780) );
  NAND2_X1 U10836 ( .A1(n9781), .A2(n9780), .ZN(P2_U3288) );
  INV_X1 U10837 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n9784) );
  NOR2_X1 U10838 ( .A1(n9819), .A2(n9784), .ZN(P2_U3297) );
  INV_X1 U10839 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n9785) );
  NOR2_X1 U10840 ( .A1(n9819), .A2(n9785), .ZN(P2_U3298) );
  INV_X1 U10841 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n9786) );
  NOR2_X1 U10842 ( .A1(n9819), .A2(n9786), .ZN(P2_U3299) );
  INV_X1 U10843 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n9787) );
  NOR2_X1 U10844 ( .A1(n9819), .A2(n9787), .ZN(P2_U3300) );
  NOR2_X1 U10845 ( .A1(n9819), .A2(n9788), .ZN(P2_U3301) );
  INV_X1 U10846 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n9789) );
  NOR2_X1 U10847 ( .A1(n9799), .A2(n9789), .ZN(P2_U3302) );
  INV_X1 U10848 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9790) );
  NOR2_X1 U10849 ( .A1(n9799), .A2(n9790), .ZN(P2_U3303) );
  INV_X1 U10850 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n9791) );
  NOR2_X1 U10851 ( .A1(n9799), .A2(n9791), .ZN(P2_U3304) );
  INV_X1 U10852 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n9792) );
  NOR2_X1 U10853 ( .A1(n9799), .A2(n9792), .ZN(P2_U3305) );
  INV_X1 U10854 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n9793) );
  NOR2_X1 U10855 ( .A1(n9799), .A2(n9793), .ZN(P2_U3306) );
  NOR2_X1 U10856 ( .A1(n9799), .A2(n9794), .ZN(P2_U3307) );
  NOR2_X1 U10857 ( .A1(n9799), .A2(n9795), .ZN(P2_U3308) );
  INV_X1 U10858 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n9796) );
  NOR2_X1 U10859 ( .A1(n9799), .A2(n9796), .ZN(P2_U3309) );
  NOR2_X1 U10860 ( .A1(n9799), .A2(n9797), .ZN(P2_U3310) );
  NOR2_X1 U10861 ( .A1(n9799), .A2(n9798), .ZN(P2_U3311) );
  INV_X1 U10862 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9800) );
  NOR2_X1 U10863 ( .A1(n9819), .A2(n9800), .ZN(P2_U3312) );
  INV_X1 U10864 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n9801) );
  NOR2_X1 U10865 ( .A1(n9819), .A2(n9801), .ZN(P2_U3313) );
  INV_X1 U10866 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n9802) );
  NOR2_X1 U10867 ( .A1(n9819), .A2(n9802), .ZN(P2_U3314) );
  NOR2_X1 U10868 ( .A1(n9819), .A2(n9803), .ZN(P2_U3315) );
  NOR2_X1 U10869 ( .A1(n9819), .A2(n9804), .ZN(P2_U3316) );
  INV_X1 U10870 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n9805) );
  NOR2_X1 U10871 ( .A1(n9819), .A2(n9805), .ZN(P2_U3317) );
  INV_X1 U10872 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n9806) );
  NOR2_X1 U10873 ( .A1(n9819), .A2(n9806), .ZN(P2_U3318) );
  INV_X1 U10874 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n9807) );
  NOR2_X1 U10875 ( .A1(n9819), .A2(n9807), .ZN(P2_U3319) );
  INV_X1 U10876 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n9808) );
  NOR2_X1 U10877 ( .A1(n9819), .A2(n9808), .ZN(P2_U3320) );
  INV_X1 U10878 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n9809) );
  NOR2_X1 U10879 ( .A1(n9819), .A2(n9809), .ZN(P2_U3321) );
  INV_X1 U10880 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n9810) );
  NOR2_X1 U10881 ( .A1(n9819), .A2(n9810), .ZN(P2_U3322) );
  INV_X1 U10882 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n9811) );
  NOR2_X1 U10883 ( .A1(n9819), .A2(n9811), .ZN(P2_U3323) );
  INV_X1 U10884 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n9812) );
  NOR2_X1 U10885 ( .A1(n9819), .A2(n9812), .ZN(P2_U3324) );
  INV_X1 U10886 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n9813) );
  NOR2_X1 U10887 ( .A1(n9819), .A2(n9813), .ZN(P2_U3325) );
  INV_X1 U10888 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9814) );
  NOR2_X1 U10889 ( .A1(n9819), .A2(n9814), .ZN(P2_U3326) );
  OAI22_X1 U10890 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n9819), .B1(n9818), .B2(
        n9815), .ZN(n9816) );
  INV_X1 U10891 ( .A(n9816), .ZN(P2_U3437) );
  OAI22_X1 U10892 ( .A1(P2_D_REG_1__SCAN_IN), .A2(n9819), .B1(n9818), .B2(
        n9817), .ZN(n9820) );
  INV_X1 U10893 ( .A(n9820), .ZN(P2_U3438) );
  AOI22_X1 U10894 ( .A1(n9823), .A2(n9894), .B1(n9822), .B2(n9821), .ZN(n9824)
         );
  AND2_X1 U10895 ( .A1(n9825), .A2(n9824), .ZN(n9898) );
  INV_X1 U10896 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9826) );
  AOI22_X1 U10897 ( .A1(n9872), .A2(n9898), .B1(n9826), .B2(n9895), .ZN(
        P2_U3451) );
  AOI22_X1 U10898 ( .A1(n9828), .A2(n9836), .B1(n9835), .B2(n9827), .ZN(n9829)
         );
  NAND2_X1 U10899 ( .A1(n9830), .A2(n9829), .ZN(n9831) );
  AOI21_X1 U10900 ( .B1(n9894), .B2(n9832), .A(n9831), .ZN(n9899) );
  INV_X1 U10901 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9833) );
  AOI22_X1 U10902 ( .A1(n9872), .A2(n9899), .B1(n9833), .B2(n9895), .ZN(
        P2_U3457) );
  AOI22_X1 U10903 ( .A1(n9837), .A2(n9836), .B1(n9835), .B2(n9834), .ZN(n9838)
         );
  NAND2_X1 U10904 ( .A1(n9839), .A2(n9838), .ZN(n9840) );
  AOI21_X1 U10905 ( .B1(n9894), .B2(n9841), .A(n9840), .ZN(n9901) );
  INV_X1 U10906 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9842) );
  AOI22_X1 U10907 ( .A1(n9872), .A2(n9901), .B1(n9842), .B2(n9895), .ZN(
        P2_U3463) );
  INV_X1 U10908 ( .A(n9843), .ZN(n9845) );
  OAI22_X1 U10909 ( .A1(n9845), .A2(n9889), .B1(n9844), .B2(n9887), .ZN(n9846)
         );
  AOI211_X1 U10910 ( .C1(n9848), .C2(n9894), .A(n9847), .B(n9846), .ZN(n9903)
         );
  INV_X1 U10911 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9849) );
  AOI22_X1 U10912 ( .A1(n9872), .A2(n9903), .B1(n9849), .B2(n9895), .ZN(
        P2_U3469) );
  OAI22_X1 U10913 ( .A1(n9851), .A2(n9889), .B1(n9850), .B2(n9887), .ZN(n9853)
         );
  AOI211_X1 U10914 ( .C1(n9854), .C2(n9894), .A(n9853), .B(n9852), .ZN(n9905)
         );
  AOI22_X1 U10915 ( .A1(n9872), .A2(n9905), .B1(n9855), .B2(n9895), .ZN(
        P2_U3472) );
  NOR2_X1 U10916 ( .A1(n9857), .A2(n9856), .ZN(n9861) );
  OAI22_X1 U10917 ( .A1(n9859), .A2(n9889), .B1(n9858), .B2(n9887), .ZN(n9860)
         );
  NOR3_X1 U10918 ( .A1(n9862), .A2(n9861), .A3(n9860), .ZN(n9906) );
  AOI22_X1 U10919 ( .A1(n9872), .A2(n9906), .B1(n9863), .B2(n9895), .ZN(
        P2_U3475) );
  INV_X1 U10920 ( .A(n9864), .ZN(n9865) );
  OAI22_X1 U10921 ( .A1(n9866), .A2(n9889), .B1(n9865), .B2(n9887), .ZN(n9867)
         );
  AOI21_X1 U10922 ( .B1(n9868), .B2(n9878), .A(n9867), .ZN(n9869) );
  AND2_X1 U10923 ( .A1(n9870), .A2(n9869), .ZN(n9907) );
  INV_X1 U10924 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9871) );
  AOI22_X1 U10925 ( .A1(n9872), .A2(n9907), .B1(n9871), .B2(n9895), .ZN(
        P2_U3478) );
  OAI22_X1 U10926 ( .A1(n9874), .A2(n9889), .B1(n9873), .B2(n9887), .ZN(n9876)
         );
  AOI211_X1 U10927 ( .C1(n9878), .C2(n9877), .A(n9876), .B(n9875), .ZN(n9908)
         );
  AOI22_X1 U10928 ( .A1(n9872), .A2(n9908), .B1(n9879), .B2(n9895), .ZN(
        P2_U3481) );
  INV_X1 U10929 ( .A(n9880), .ZN(n9885) );
  OAI22_X1 U10930 ( .A1(n9882), .A2(n9889), .B1(n9881), .B2(n9887), .ZN(n9884)
         );
  AOI211_X1 U10931 ( .C1(n9885), .C2(n9894), .A(n9884), .B(n9883), .ZN(n9909)
         );
  INV_X1 U10932 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9886) );
  AOI22_X1 U10933 ( .A1(n9872), .A2(n9909), .B1(n9886), .B2(n9895), .ZN(
        P2_U3484) );
  OAI22_X1 U10934 ( .A1(n9890), .A2(n9889), .B1(n9888), .B2(n9887), .ZN(n9892)
         );
  AOI211_X1 U10935 ( .C1(n9894), .C2(n9893), .A(n9892), .B(n9891), .ZN(n9912)
         );
  INV_X1 U10936 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9896) );
  AOI22_X1 U10937 ( .A1(n9872), .A2(n9912), .B1(n9896), .B2(n9895), .ZN(
        P2_U3487) );
  INV_X1 U10938 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9897) );
  AOI22_X1 U10939 ( .A1(n4260), .A2(n9898), .B1(n9897), .B2(n9910), .ZN(
        P2_U3520) );
  AOI22_X1 U10940 ( .A1(n4260), .A2(n9899), .B1(n6516), .B2(n9910), .ZN(
        P2_U3522) );
  INV_X1 U10941 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9900) );
  AOI22_X1 U10942 ( .A1(n4260), .A2(n9901), .B1(n9900), .B2(n9910), .ZN(
        P2_U3524) );
  INV_X1 U10943 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9902) );
  AOI22_X1 U10944 ( .A1(n4260), .A2(n9903), .B1(n9902), .B2(n9910), .ZN(
        P2_U3526) );
  INV_X1 U10945 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9904) );
  AOI22_X1 U10946 ( .A1(n4260), .A2(n9905), .B1(n9904), .B2(n9910), .ZN(
        P2_U3527) );
  AOI22_X1 U10947 ( .A1(n4260), .A2(n9906), .B1(n6527), .B2(n9910), .ZN(
        P2_U3528) );
  AOI22_X1 U10948 ( .A1(n4260), .A2(n9907), .B1(n4448), .B2(n9910), .ZN(
        P2_U3529) );
  AOI22_X1 U10949 ( .A1(n4260), .A2(n9908), .B1(n6529), .B2(n9910), .ZN(
        P2_U3530) );
  AOI22_X1 U10950 ( .A1(n4260), .A2(n9909), .B1(n6530), .B2(n9910), .ZN(
        P2_U3531) );
  AOI22_X1 U10951 ( .A1(n4260), .A2(n9912), .B1(n9911), .B2(n9910), .ZN(
        P2_U3532) );
  INV_X1 U10952 ( .A(n9913), .ZN(n9914) );
  NAND2_X1 U10953 ( .A1(n9915), .A2(n9914), .ZN(n9916) );
  XOR2_X1 U10954 ( .A(n9917), .B(n9916), .Z(ADD_1071_U5) );
  XOR2_X1 U10955 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U10956 ( .B1(n9920), .B2(n9919), .A(n9918), .ZN(ADD_1071_U56) );
  OAI21_X1 U10957 ( .B1(n9923), .B2(n9922), .A(n9921), .ZN(ADD_1071_U57) );
  OAI21_X1 U10958 ( .B1(n9926), .B2(n9925), .A(n9924), .ZN(ADD_1071_U58) );
  OAI21_X1 U10959 ( .B1(n9929), .B2(n9928), .A(n9927), .ZN(ADD_1071_U59) );
  OAI21_X1 U10960 ( .B1(n9932), .B2(n9931), .A(n9930), .ZN(ADD_1071_U60) );
  OAI21_X1 U10961 ( .B1(n9935), .B2(n9934), .A(n9933), .ZN(ADD_1071_U61) );
  AOI21_X1 U10962 ( .B1(n9938), .B2(n9937), .A(n9936), .ZN(ADD_1071_U62) );
  AOI21_X1 U10963 ( .B1(n9941), .B2(n9940), .A(n9939), .ZN(ADD_1071_U63) );
  XOR2_X1 U10964 ( .A(n9942), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U10965 ( .A1(n9944), .A2(n9943), .ZN(n9945) );
  XOR2_X1 U10966 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n9945), .Z(ADD_1071_U51) );
  OAI21_X1 U10967 ( .B1(n9948), .B2(n9947), .A(n9946), .ZN(n9949) );
  XNOR2_X1 U10968 ( .A(n9949), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U10969 ( .B1(n9952), .B2(n9951), .A(n9950), .ZN(ADD_1071_U47) );
  XOR2_X1 U10970 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n9953), .Z(ADD_1071_U48) );
  XOR2_X1 U10971 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n9954), .Z(ADD_1071_U49) );
  XOR2_X1 U10972 ( .A(n9956), .B(n9955), .Z(ADD_1071_U54) );
  XOR2_X1 U10973 ( .A(n9958), .B(n9957), .Z(ADD_1071_U53) );
  XNOR2_X1 U10974 ( .A(n9960), .B(n9959), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4767 ( .A(n6463), .Z(n8106) );
  CLKBUF_X1 U4768 ( .A(n7141), .Z(n7901) );
  CLKBUF_X2 U4779 ( .A(n5746), .Z(n5900) );
endmodule

