

module b21_C_gen_AntiSAT_k_128_9 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, 
        keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, 
        keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, 
        keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, 
        keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, 
        keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, 
        keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, 
        keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, 
        keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, 
        keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, 
        keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, 
        keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, 
        keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117;

  INV_X1 U4815 ( .A(n5022), .ZN(n8840) );
  CLKBUF_X2 U4816 ( .A(n5634), .Z(n5215) );
  CLKBUF_X2 U4817 ( .A(n5013), .Z(n5685) );
  INV_X1 U4819 ( .A(n4964), .ZN(n8835) );
  NAND2_X1 U4820 ( .A1(n9508), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4916) );
  CLKBUF_X1 U4821 ( .A(n7796), .Z(n4310) );
  OAI21_X1 U4822 ( .B1(n6492), .B2(n6468), .A(n8440), .ZN(n7796) );
  NOR2_X2 U4823 ( .A1(n5719), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n4865) );
  INV_X1 U4824 ( .A(n5606), .ZN(n8625) );
  XNOR2_X1 U4825 ( .A(n6500), .B(n8969), .ZN(n6501) );
  INV_X2 U4826 ( .A(n8539), .ZN(n10050) );
  INV_X1 U4827 ( .A(n7157), .ZN(n10009) );
  INV_X1 U4828 ( .A(n5010), .ZN(n5477) );
  NAND2_X1 U4829 ( .A1(n6211), .A2(n5676), .ZN(n4949) );
  INV_X1 U4830 ( .A(n7246), .ZN(n9949) );
  OAI211_X2 U4831 ( .C1(n5864), .C2(n6243), .A(n5776), .B(n5775), .ZN(n7217)
         );
  AOI211_X1 U4832 ( .C1(n9935), .C2(n9429), .A(n9428), .B(n9427), .ZN(n9430)
         );
  NAND2_X1 U4833 ( .A1(n7692), .A2(n7693), .ZN(n7691) );
  AND2_X1 U4834 ( .A1(n8718), .A2(n4449), .ZN(n8645) );
  NAND3_X1 U4835 ( .A1(n4864), .A2(n4865), .A3(n4355), .ZN(n4311) );
  XNOR2_X2 U4836 ( .A(n4919), .B(n4918), .ZN(n4922) );
  XNOR2_X2 U4837 ( .A(n4916), .B(P1_IR_REG_30__SCAN_IN), .ZN(n4920) );
  OAI22_X2 U4838 ( .A1(n7768), .A2(n7767), .B1(n7632), .B2(n7631), .ZN(n7726)
         );
  OAI211_X2 U4839 ( .C1(n8837), .C2(n6257), .A(n5086), .B(n5085), .ZN(n7139)
         );
  NAND3_X2 U4840 ( .A1(n5646), .A2(n5641), .A3(n5643), .ZN(n4934) );
  NAND3_X2 U4841 ( .A1(n5863), .A2(n5862), .A3(n4430), .ZN(n6937) );
  OAI222_X1 U4842 ( .A1(n7689), .A2(n6263), .B1(n9512), .B2(n6262), .C1(
        P1_U3084), .C2(n6261), .ZN(P1_U3346) );
  OAI222_X1 U4843 ( .A1(n7365), .A2(n6260), .B1(n8597), .B2(n6262), .C1(n7694), 
        .C2(n6709), .ZN(P2_U3351) );
  XNOR2_X2 U4844 ( .A(n4892), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5663) );
  AND2_X1 U4845 ( .A1(n6485), .A2(n6542), .ZN(n6489) );
  INV_X1 U4846 ( .A(n5800), .ZN(n5779) );
  NAND2_X1 U4847 ( .A1(n6480), .A2(n4742), .ZN(n6546) );
  NAND2_X4 U4848 ( .A1(n8591), .A2(n5733), .ZN(n5801) );
  NAND2_X1 U4849 ( .A1(n6605), .A2(n6609), .ZN(n6603) );
  INV_X1 U4850 ( .A(n4934), .ZN(n6199) );
  INV_X2 U4851 ( .A(n7833), .ZN(n8152) );
  OR2_X1 U4853 ( .A1(n8678), .A2(n4368), .ZN(n4790) );
  AOI21_X1 U4854 ( .B1(n5490), .B2(n4524), .A(n4797), .ZN(n5537) );
  NAND2_X1 U4855 ( .A1(n4440), .A2(n4442), .ZN(n5490) );
  OAI21_X1 U4856 ( .B1(n8892), .B2(n8891), .A(n9002), .ZN(n8893) );
  NOR2_X1 U4857 ( .A1(n8857), .A2(n8856), .ZN(n8892) );
  MUX2_X1 U4858 ( .A(n8847), .B(n8846), .S(n8850), .Z(n8857) );
  AOI21_X1 U4859 ( .B1(n5415), .B2(n4521), .A(n4518), .ZN(n4517) );
  NAND2_X1 U4860 ( .A1(n8668), .A2(n5392), .ZN(n5415) );
  NAND2_X1 U4861 ( .A1(n8659), .A2(n5367), .ZN(n8669) );
  NAND2_X1 U4862 ( .A1(n4726), .A2(n4727), .ZN(n7755) );
  INV_X1 U4863 ( .A(n7475), .ZN(n5280) );
  OR2_X1 U4864 ( .A1(n4324), .A2(n8479), .ZN(n8236) );
  NAND2_X1 U4865 ( .A1(n7369), .A2(n5223), .ZN(n7502) );
  NAND2_X1 U4866 ( .A1(n7491), .A2(n7490), .ZN(n7535) );
  NAND3_X1 U4867 ( .A1(n4814), .A2(n5174), .A3(n7092), .ZN(n7222) );
  NAND2_X1 U4868 ( .A1(n7091), .A2(n7093), .ZN(n4814) );
  NAND2_X1 U4869 ( .A1(n5146), .A2(n5145), .ZN(n7092) );
  NAND2_X1 U4870 ( .A1(n5401), .A2(n5400), .ZN(n9468) );
  NAND2_X1 U4871 ( .A1(n5762), .A2(n5761), .ZN(n8449) );
  NAND2_X1 U4872 ( .A1(n5923), .A2(n5922), .ZN(n10046) );
  OR2_X1 U4873 ( .A1(n7240), .A2(n7294), .ZN(n7290) );
  INV_X2 U4874 ( .A(n8438), .ZN(n8406) );
  NAND2_X1 U4875 ( .A1(n6489), .A2(n6488), .ZN(n6543) );
  OAI21_X1 U4876 ( .B1(n6421), .B2(n4817), .A(n6424), .ZN(n4816) );
  AND3_X1 U4877 ( .A1(n4937), .A2(n4936), .A3(n4935), .ZN(n6367) );
  NOR2_X1 U4878 ( .A1(n9806), .A2(n7018), .ZN(n9787) );
  AND4_X1 U4879 ( .A1(n5794), .A2(n5793), .A3(n5792), .A4(n5791), .ZN(n6772)
         );
  NAND2_X1 U4880 ( .A1(n4613), .A2(n4925), .ZN(n9028) );
  NOR2_X1 U4881 ( .A1(n4338), .A2(n4612), .ZN(n4613) );
  INV_X2 U4882 ( .A(n6546), .ZN(n7650) );
  CLKBUF_X3 U4883 ( .A(n6546), .Z(n7666) );
  INV_X1 U4884 ( .A(n7056), .ZN(n9927) );
  INV_X2 U4885 ( .A(n5864), .ZN(n7828) );
  AND2_X2 U4886 ( .A1(n4951), .A2(n4326), .ZN(n8969) );
  INV_X2 U4888 ( .A(n6603), .ZN(n5993) );
  NAND2_X1 U4889 ( .A1(n7688), .A2(n7587), .ZN(n5010) );
  AND2_X2 U4890 ( .A1(n5729), .A2(n5728), .ZN(n8595) );
  XNOR2_X1 U4891 ( .A(n6131), .B(n6130), .ZN(n8020) );
  NAND2_X1 U4892 ( .A1(n4949), .A2(n7824), .ZN(n5022) );
  OR2_X1 U4893 ( .A1(n5727), .A2(n4847), .ZN(n5728) );
  XNOR2_X1 U4894 ( .A(n6126), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8019) );
  NAND2_X1 U4895 ( .A1(n4848), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5724) );
  XNOR2_X1 U4896 ( .A(n6128), .B(n6127), .ZN(n7833) );
  XNOR2_X1 U4897 ( .A(n4888), .B(n4897), .ZN(n6866) );
  XNOR2_X1 U4898 ( .A(n4903), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5646) );
  OAI21_X1 U4899 ( .B1(n4889), .B2(n4531), .A(n4532), .ZN(n4892) );
  AND2_X1 U4900 ( .A1(n4403), .A2(n4900), .ZN(n4402) );
  AND2_X1 U4901 ( .A1(n5053), .A2(n4879), .ZN(n4403) );
  AND2_X1 U4902 ( .A1(n4882), .A2(n4822), .ZN(n4821) );
  AND3_X1 U4903 ( .A1(n4516), .A2(n4881), .A3(n4880), .ZN(n4882) );
  AND3_X1 U4904 ( .A1(n6114), .A2(n6127), .A3(n4592), .ZN(n5713) );
  NOR2_X1 U4905 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4880) );
  NOR2_X1 U4906 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4516) );
  NOR2_X1 U4907 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4881) );
  NOR2_X1 U4908 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5795) );
  INV_X1 U4909 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6114) );
  NOR2_X1 U4910 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5019) );
  INV_X4 U4911 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U4912 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9731) );
  XNOR2_X1 U4913 ( .A(n4931), .B(P1_IR_REG_28__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U4914 ( .A1(n4920), .A2(n4922), .ZN(n4313) );
  NOR2_X2 U4915 ( .A1(n7317), .A2(n8559), .ZN(n7355) );
  INV_X1 U4916 ( .A(n8595), .ZN(n5733) );
  NAND2_X1 U4917 ( .A1(n4922), .A2(n7587), .ZN(n5013) );
  AND2_X1 U4918 ( .A1(n7688), .A2(n4920), .ZN(n4987) );
  INV_X1 U4919 ( .A(n5057), .ZN(n5427) );
  INV_X1 U4920 ( .A(n8837), .ZN(n5426) );
  INV_X1 U4921 ( .A(n7734), .ZN(n4739) );
  NAND2_X1 U4922 ( .A1(n4419), .A2(n4325), .ZN(n4418) );
  INV_X1 U4923 ( .A(n6066), .ZN(n4834) );
  OR2_X1 U4924 ( .A1(n8476), .A2(n8245), .ZN(n7980) );
  NOR2_X1 U4925 ( .A1(n8279), .A2(n4844), .ZN(n4843) );
  INV_X1 U4926 ( .A(n6025), .ZN(n4844) );
  NOR2_X1 U4927 ( .A1(n4691), .A2(n4688), .ZN(n4687) );
  INV_X1 U4928 ( .A(n7934), .ZN(n4688) );
  INV_X1 U4929 ( .A(n4692), .ZN(n4691) );
  OR2_X1 U4930 ( .A1(n8521), .A2(n8369), .ZN(n7947) );
  AOI21_X1 U4931 ( .B1(n4679), .B2(n4681), .A(n4678), .ZN(n4677) );
  INV_X1 U4932 ( .A(n4684), .ZN(n4679) );
  INV_X1 U4933 ( .A(n7928), .ZN(n4678) );
  NAND2_X1 U4934 ( .A1(n8027), .A2(n8152), .ZN(n8017) );
  NAND2_X1 U4935 ( .A1(n5737), .A2(n5722), .ZN(n5739) );
  AND2_X1 U4936 ( .A1(n4355), .A2(n5721), .ZN(n4605) );
  INV_X1 U4937 ( .A(n5860), .ZN(n4864) );
  AND2_X1 U4938 ( .A1(n5966), .A2(n4743), .ZN(n6125) );
  AND2_X1 U4939 ( .A1(n4744), .A2(n4361), .ZN(n4743) );
  INV_X1 U4940 ( .A(n5964), .ZN(n5966) );
  NOR2_X2 U4941 ( .A1(n4858), .A2(n5807), .ZN(n5835) );
  OR2_X1 U4942 ( .A1(n4860), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n4858) );
  AND2_X1 U4943 ( .A1(n5555), .A2(n5554), .ZN(n5557) );
  AND2_X1 U4944 ( .A1(n7569), .A2(n4806), .ZN(n4809) );
  OR2_X1 U4945 ( .A1(n9421), .A2(n9192), .ZN(n9150) );
  NOR2_X1 U4946 ( .A1(n9381), .A2(n8902), .ZN(n4631) );
  AND2_X1 U4947 ( .A1(n4655), .A2(n4413), .ZN(n4412) );
  OR2_X1 U4948 ( .A1(n4663), .A2(n4414), .ZN(n4413) );
  AND2_X1 U4949 ( .A1(n4660), .A2(n4315), .ZN(n4655) );
  AND2_X1 U4950 ( .A1(n8872), .A2(n6516), .ZN(n4407) );
  OR2_X1 U4951 ( .A1(n6409), .A2(n6408), .ZN(n6943) );
  OR2_X1 U4952 ( .A1(n7583), .A2(n7582), .ZN(n7584) );
  OAI21_X1 U4953 ( .B1(n5589), .B2(n5588), .A(n5587), .ZN(n5614) );
  NAND2_X1 U4954 ( .A1(n4755), .A2(n4373), .ZN(n4474) );
  AND2_X1 U4955 ( .A1(n5538), .A2(n4479), .ZN(n4478) );
  NOR2_X1 U4956 ( .A1(n5493), .A2(n4762), .ZN(n4761) );
  INV_X1 U4957 ( .A(n5471), .ZN(n4762) );
  INV_X1 U4958 ( .A(n5447), .ZN(n4480) );
  AND2_X1 U4959 ( .A1(n5471), .A2(n5452), .ZN(n5469) );
  OAI21_X1 U4960 ( .B1(n5315), .B2(n5314), .A(n5317), .ZN(n5340) );
  INV_X1 U4961 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4822) );
  AND2_X1 U4962 ( .A1(n5287), .A2(n5263), .ZN(n5285) );
  INV_X1 U4963 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4879) );
  OAI21_X1 U4964 ( .B1(n4456), .B2(n4453), .A(n4451), .ZN(n5198) );
  NOR2_X1 U4965 ( .A1(n4341), .A2(n4452), .ZN(n4451) );
  INV_X1 U4966 ( .A(n5178), .ZN(n4452) );
  OR2_X1 U4967 ( .A1(n7735), .A2(n4739), .ZN(n4738) );
  NAND2_X1 U4968 ( .A1(n7735), .A2(n4739), .ZN(n4737) );
  OAI21_X1 U4969 ( .B1(n4397), .B2(n8016), .A(n8015), .ZN(n8021) );
  AOI21_X1 U4970 ( .B1(n8009), .B2(n8008), .A(n4398), .ZN(n4397) );
  OR3_X1 U4971 ( .A1(n7368), .A2(n6133), .A3(n6135), .ZN(n6599) );
  AND2_X1 U4972 ( .A1(n4832), .A2(n4420), .ZN(n4419) );
  OR2_X1 U4973 ( .A1(n4325), .A2(n8224), .ZN(n4420) );
  INV_X1 U4974 ( .A(n4833), .ZN(n4832) );
  OAI21_X1 U4975 ( .B1(n8208), .B2(n4834), .A(n8194), .ZN(n4833) );
  OR2_X1 U4976 ( .A1(n8256), .A2(n4705), .ZN(n4702) );
  OR2_X1 U4977 ( .A1(n4707), .A2(n8224), .ZN(n4705) );
  OR2_X1 U4978 ( .A1(n8256), .A2(n4707), .ZN(n4706) );
  OR2_X1 U4979 ( .A1(n8493), .A2(n8257), .ZN(n8254) );
  NAND2_X1 U4980 ( .A1(n4825), .A2(n4823), .ZN(n8302) );
  NAND2_X1 U4981 ( .A1(n8332), .A2(n4826), .ZN(n4825) );
  NAND2_X1 U4982 ( .A1(n4588), .A2(n4317), .ZN(n7916) );
  AND4_X1 U4983 ( .A1(n5832), .A2(n5831), .A3(n5830), .A4(n5829), .ZN(n7166)
         );
  NAND2_X1 U4984 ( .A1(n6603), .A2(n8835), .ZN(n5864) );
  AND2_X1 U4985 ( .A1(n6603), .A2(n7824), .ZN(n5821) );
  NAND2_X1 U4986 ( .A1(n6139), .A2(n6138), .ZN(n6141) );
  OR2_X1 U4987 ( .A1(n8686), .A2(n4445), .ZN(n4440) );
  NAND2_X1 U4988 ( .A1(n4521), .A2(n4520), .ZN(n4519) );
  INV_X1 U4989 ( .A(n4533), .ZN(n4531) );
  AOI21_X1 U4990 ( .B1(n4533), .B2(n9507), .A(n9507), .ZN(n4532) );
  AOI21_X1 U4991 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_20__SCAN_IN), .ZN(n4533) );
  INV_X1 U4992 ( .A(n9170), .ZN(n9130) );
  AND2_X1 U4993 ( .A1(n5629), .A2(n5628), .ZN(n9210) );
  AOI21_X1 U4994 ( .B1(n9246), .B2(n9118), .A(n9117), .ZN(n9233) );
  OR2_X1 U4995 ( .A1(n9346), .A2(n9112), .ZN(n4652) );
  OR2_X1 U4996 ( .A1(n9818), .A2(n9375), .ZN(n4873) );
  OR2_X1 U4997 ( .A1(n9393), .A2(n9107), .ZN(n9108) );
  AND2_X1 U4998 ( .A1(n8914), .A2(n8913), .ZN(n8870) );
  AND4_X1 U4999 ( .A1(n5018), .A2(n5017), .A3(n5016), .A4(n5015), .ZN(n7045)
         );
  INV_X1 U5000 ( .A(n9772), .ZN(n9798) );
  OR2_X1 U5001 ( .A1(n6412), .A2(n6507), .ZN(n9796) );
  NAND2_X1 U5002 ( .A1(n5429), .A2(n5428), .ZN(n9462) );
  OR2_X1 U5003 ( .A1(n8850), .A2(n9002), .ZN(n9824) );
  XNOR2_X1 U5004 ( .A(n6096), .B(n6095), .ZN(n8616) );
  INV_X1 U5005 ( .A(n4751), .ZN(n6096) );
  AOI21_X1 U5006 ( .B1(n6077), .B2(n6076), .A(n4754), .ZN(n4751) );
  XNOR2_X1 U5007 ( .A(n5614), .B(n5613), .ZN(n7510) );
  NAND2_X1 U5008 ( .A1(n4963), .A2(n4962), .ZN(n5001) );
  MUX2_X1 U5009 ( .A(n7921), .B(n7920), .S(n8012), .Z(n7922) );
  MUX2_X1 U5010 ( .A(n7970), .B(n7969), .S(n8012), .Z(n7971) );
  AND2_X1 U5011 ( .A1(n7972), .A2(n8012), .ZN(n4578) );
  NOR2_X1 U5012 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4894) );
  NOR2_X1 U5013 ( .A1(n6171), .A2(n4682), .ZN(n4681) );
  OR2_X1 U5014 ( .A1(n8524), .A2(n8533), .ZN(n4602) );
  NAND2_X1 U5015 ( .A1(n4773), .A2(n5419), .ZN(n4772) );
  NAND2_X1 U5016 ( .A1(n7002), .A2(n4555), .ZN(n4554) );
  OR2_X1 U5017 ( .A1(n8455), .A2(n4611), .ZN(n4610) );
  OR2_X1 U5018 ( .A1(n8459), .A2(n8464), .ZN(n4611) );
  OR2_X1 U5019 ( .A1(n8459), .A2(n8196), .ZN(n7994) );
  NAND2_X1 U5020 ( .A1(n7974), .A2(n7976), .ZN(n4707) );
  NAND2_X1 U5021 ( .A1(n8276), .A2(n4561), .ZN(n4609) );
  OR2_X1 U5022 ( .A1(n8521), .A2(n4602), .ZN(n4601) );
  NOR2_X1 U5023 ( .A1(n6172), .A2(n4693), .ZN(n4692) );
  INV_X1 U5024 ( .A(n7940), .ZN(n4693) );
  OR2_X1 U5025 ( .A1(n8538), .A2(n8431), .ZN(n7934) );
  OR2_X1 U5026 ( .A1(n8533), .A2(n8413), .ZN(n7940) );
  NOR2_X1 U5027 ( .A1(n7854), .A2(n4856), .ZN(n4855) );
  INV_X1 U5028 ( .A(n5918), .ZN(n4856) );
  INV_X1 U5029 ( .A(n4681), .ZN(n4680) );
  NOR2_X1 U5030 ( .A1(n6170), .A2(n4685), .ZN(n4684) );
  INV_X1 U5031 ( .A(n7916), .ZN(n4685) );
  AND2_X1 U5032 ( .A1(n7907), .A2(n7915), .ZN(n7849) );
  NOR2_X1 U5033 ( .A1(n7896), .A2(n4383), .ZN(n4837) );
  NAND2_X1 U5034 ( .A1(n8046), .A2(n10019), .ZN(n7890) );
  OR2_X1 U5035 ( .A1(n5801), .A2(n6637), .ZN(n5802) );
  NAND2_X1 U5036 ( .A1(n8047), .A2(n10014), .ZN(n7889) );
  NAND2_X1 U5037 ( .A1(n7165), .A2(n6777), .ZN(n7882) );
  INV_X1 U5038 ( .A(n8020), .ZN(n7841) );
  NOR2_X1 U5039 ( .A1(n8236), .A2(n8476), .ZN(n8227) );
  NOR2_X1 U5040 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n4744) );
  NOR2_X1 U5041 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4746) );
  INV_X1 U5042 ( .A(n5807), .ZN(n4859) );
  INV_X1 U5043 ( .A(n5041), .ZN(n4813) );
  INV_X1 U5044 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4918) );
  INV_X1 U5045 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4893) );
  NOR2_X1 U5046 ( .A1(n7435), .A2(n7434), .ZN(n9043) );
  NAND2_X1 U5047 ( .A1(n4625), .A2(n9236), .ZN(n4624) );
  OR2_X1 U5048 ( .A1(n9434), .A2(n9238), .ZN(n8946) );
  AND2_X1 U5049 ( .A1(n9272), .A2(n9114), .ZN(n9143) );
  NAND2_X1 U5050 ( .A1(n4668), .A2(n9115), .ZN(n4667) );
  OR2_X1 U5051 ( .A1(n9449), .A2(n9114), .ZN(n9115) );
  OR2_X1 U5052 ( .A1(n9444), .A2(n9265), .ZN(n9145) );
  AOI21_X1 U5053 ( .B1(n4645), .B2(n4646), .A(n4347), .ZN(n4644) );
  INV_X1 U5054 ( .A(n4650), .ZN(n4645) );
  NAND2_X1 U5055 ( .A1(n4653), .A2(n9112), .ZN(n4648) );
  OR2_X1 U5056 ( .A1(n9486), .A2(n9779), .ZN(n4505) );
  NAND2_X1 U5057 ( .A1(n4504), .A2(n9818), .ZN(n4503) );
  INV_X1 U5058 ( .A(n4505), .ZN(n4504) );
  INV_X1 U5059 ( .A(n7520), .ZN(n4414) );
  AND2_X1 U5060 ( .A1(n4867), .A2(n7519), .ZN(n4663) );
  NAND2_X1 U5061 ( .A1(n9795), .A2(n8768), .ZN(n7553) );
  NAND2_X1 U5062 ( .A1(n4320), .A2(n7113), .ZN(n4633) );
  NAND2_X1 U5063 ( .A1(n5662), .A2(n9001), .ZN(n6497) );
  NAND2_X1 U5064 ( .A1(n4633), .A2(n4632), .ZN(n9795) );
  AND2_X1 U5065 ( .A1(n8898), .A2(n8897), .ZN(n4632) );
  AND2_X1 U5066 ( .A1(n4405), .A2(n4404), .ZN(n7039) );
  INV_X1 U5067 ( .A(n6804), .ZN(n4406) );
  OAI21_X1 U5068 ( .B1(n4750), .B2(n4753), .A(n4749), .ZN(n7583) );
  AOI21_X1 U5069 ( .B1(n4752), .B2(n4754), .A(n4386), .ZN(n4749) );
  NAND2_X1 U5070 ( .A1(n5616), .A2(n5615), .ZN(n6077) );
  NAND2_X1 U5071 ( .A1(n5614), .A2(n5613), .ZN(n5616) );
  NAND2_X1 U5072 ( .A1(n5567), .A2(n5566), .ZN(n5589) );
  NOR2_X1 U5073 ( .A1(n4476), .A2(n4377), .ZN(n4473) );
  AND2_X1 U5074 ( .A1(n5538), .A2(n4477), .ZN(n4476) );
  INV_X1 U5075 ( .A(n5515), .ZN(n4477) );
  NAND2_X1 U5076 ( .A1(n5449), .A2(n5448), .ZN(n5470) );
  NAND2_X1 U5077 ( .A1(n4459), .A2(n4460), .ZN(n5315) );
  AOI21_X1 U5078 ( .B1(n4463), .B2(n5225), .A(n4461), .ZN(n4460) );
  AND2_X1 U5079 ( .A1(n5178), .A2(n5153), .ZN(n5176) );
  NAND2_X1 U5080 ( .A1(n4929), .A2(n4928), .ZN(n4964) );
  NAND2_X1 U5081 ( .A1(n9730), .A2(n4926), .ZN(n4929) );
  NAND2_X1 U5082 ( .A1(n9731), .A2(n4927), .ZN(n4928) );
  INV_X1 U5083 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4926) );
  INV_X1 U5084 ( .A(n6912), .ZN(n4723) );
  INV_X1 U5085 ( .A(n6796), .ZN(n4720) );
  INV_X1 U5086 ( .A(n6910), .ZN(n4724) );
  INV_X1 U5087 ( .A(n7604), .ZN(n4730) );
  OR2_X1 U5088 ( .A1(n7611), .A2(n4729), .ZN(n4728) );
  NAND2_X1 U5089 ( .A1(n7702), .A2(n7604), .ZN(n4729) );
  AND2_X1 U5090 ( .A1(n7396), .A2(n7393), .ZN(n4717) );
  INV_X1 U5091 ( .A(n4737), .ZN(n4736) );
  AND2_X1 U5092 ( .A1(n7791), .A2(n4734), .ZN(n4733) );
  NAND2_X1 U5093 ( .A1(n4735), .A2(n4737), .ZN(n4734) );
  NAND2_X1 U5094 ( .A1(n6113), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6124) );
  AND2_X1 U5095 ( .A1(n5730), .A2(n8595), .ZN(n5798) );
  AND4_X1 U5096 ( .A1(n5859), .A2(n5858), .A3(n5857), .A4(n5856), .ZN(n6914)
         );
  NOR2_X1 U5097 ( .A1(n6644), .A2(n4329), .ZN(n6632) );
  OR2_X1 U5098 ( .A1(n6632), .A2(n6631), .ZN(n4541) );
  OR2_X1 U5099 ( .A1(n8056), .A2(n8057), .ZN(n4539) );
  AND2_X1 U5100 ( .A1(n4539), .A2(n4538), .ZN(n8070) );
  NAND2_X1 U5101 ( .A1(n8054), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4538) );
  OR2_X1 U5102 ( .A1(n8070), .A2(n8071), .ZN(n4537) );
  AND2_X1 U5103 ( .A1(n8090), .A2(n7006), .ZN(n4550) );
  INV_X1 U5104 ( .A(n7006), .ZN(n4547) );
  NOR2_X1 U5105 ( .A1(n4554), .A2(n8100), .ZN(n4553) );
  NAND2_X1 U5106 ( .A1(n5740), .A2(n5739), .ZN(n6605) );
  MUX2_X1 U5107 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5738), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n5740) );
  NOR2_X1 U5108 ( .A1(n8211), .A2(n4610), .ZN(n8165) );
  NOR2_X1 U5109 ( .A1(n4877), .A2(n8459), .ZN(n8173) );
  INV_X1 U5110 ( .A(n6056), .ZN(n4831) );
  NAND2_X1 U5111 ( .A1(n4702), .A2(n4700), .ZN(n4458) );
  AND2_X1 U5112 ( .A1(n4703), .A2(n4701), .ZN(n4700) );
  INV_X1 U5113 ( .A(n4704), .ZN(n4703) );
  OAI21_X1 U5114 ( .B1(n8224), .B2(n6178), .A(n7980), .ZN(n4704) );
  NAND2_X1 U5115 ( .A1(n8220), .A2(n6056), .ZN(n8204) );
  NAND2_X1 U5116 ( .A1(n8204), .A2(n8208), .ZN(n8203) );
  AND2_X1 U5117 ( .A1(n6055), .A2(n6054), .ZN(n8245) );
  OAI21_X1 U5118 ( .B1(n8284), .B2(n8269), .A(n8264), .ZN(n8235) );
  AND2_X1 U5119 ( .A1(n8252), .A2(n6177), .ZN(n8256) );
  AOI21_X1 U5120 ( .B1(n4843), .B2(n4425), .A(n4344), .ZN(n4424) );
  INV_X1 U5121 ( .A(n6024), .ZN(n4425) );
  OR2_X1 U5122 ( .A1(n8290), .A2(n4426), .ZN(n4423) );
  INV_X1 U5123 ( .A(n4843), .ZN(n4426) );
  NAND2_X1 U5124 ( .A1(n4423), .A2(n4421), .ZN(n8264) );
  NOR2_X1 U5125 ( .A1(n4422), .A2(n8261), .ZN(n4421) );
  INV_X1 U5126 ( .A(n4424), .ZN(n4422) );
  OR2_X1 U5127 ( .A1(n8319), .A2(n8510), .ZN(n8306) );
  AOI21_X1 U5128 ( .B1(n4829), .B2(n4827), .A(n4342), .ZN(n4826) );
  INV_X1 U5129 ( .A(n5991), .ZN(n4827) );
  AND2_X1 U5130 ( .A1(n8317), .A2(n4333), .ZN(n4829) );
  AND2_X1 U5131 ( .A1(n6173), .A2(n7947), .ZN(n8340) );
  NAND2_X1 U5132 ( .A1(n8349), .A2(n5979), .ZN(n8332) );
  AND2_X1 U5133 ( .A1(n7947), .A2(n7948), .ZN(n8352) );
  AND2_X1 U5134 ( .A1(n8383), .A2(n5949), .ZN(n8366) );
  NAND2_X1 U5135 ( .A1(n8366), .A2(n8367), .ZN(n8365) );
  OAI21_X1 U5136 ( .B1(n5919), .B2(n4853), .A(n4849), .ZN(n5934) );
  AND2_X1 U5137 ( .A1(n4334), .A2(n4850), .ZN(n4849) );
  OR2_X1 U5138 ( .A1(n10046), .A2(n8040), .ZN(n4857) );
  NAND2_X1 U5139 ( .A1(n5919), .A2(n4855), .ZN(n4854) );
  NAND2_X1 U5140 ( .A1(n4854), .A2(n4852), .ZN(n8426) );
  NAND2_X1 U5141 ( .A1(n6169), .A2(n4684), .ZN(n4683) );
  AND2_X1 U5142 ( .A1(n7928), .A2(n7926), .ZN(n7854) );
  AOI21_X1 U5143 ( .B1(n4862), .B2(n7901), .A(n4356), .ZN(n4434) );
  NAND2_X1 U5144 ( .A1(n7256), .A2(n4862), .ZN(n7309) );
  AND4_X1 U5145 ( .A1(n5888), .A2(n5887), .A3(n5886), .A4(n5885), .ZN(n7349)
         );
  AND4_X1 U5146 ( .A1(n5917), .A2(n5916), .A3(n5915), .A4(n5914), .ZN(n7467)
         );
  AND4_X1 U5147 ( .A1(n5873), .A2(n5872), .A3(n5871), .A4(n5870), .ZN(n7313)
         );
  NAND2_X1 U5148 ( .A1(n4433), .A2(n5878), .ZN(n7256) );
  OR2_X1 U5149 ( .A1(n7027), .A2(n6937), .ZN(n7260) );
  OR2_X1 U5150 ( .A1(n5850), .A2(n4841), .ZN(n4840) );
  AND2_X1 U5151 ( .A1(n7899), .A2(n7898), .ZN(n7896) );
  OR2_X1 U5152 ( .A1(n7153), .A2(n6777), .ZN(n7171) );
  NAND2_X1 U5153 ( .A1(n6490), .A2(n6605), .ZN(n8430) );
  NOR2_X1 U5154 ( .A1(n7217), .A2(n10001), .ZN(n7154) );
  OR3_X1 U5155 ( .A1(n6153), .A2(n6465), .A3(n6152), .ZN(n6193) );
  OR2_X1 U5156 ( .A1(n6479), .A2(n7841), .ZN(n6936) );
  AND2_X1 U5157 ( .A1(n4672), .A2(n4670), .ZN(n8457) );
  AOI21_X1 U5158 ( .B1(n8032), .B2(n8341), .A(n4671), .ZN(n4670) );
  NAND2_X1 U5159 ( .A1(n6181), .A2(n8434), .ZN(n4672) );
  NOR2_X1 U5160 ( .A1(n6187), .A2(n6186), .ZN(n4671) );
  AND2_X1 U5161 ( .A1(n6136), .A2(n7511), .ZN(n9992) );
  NAND2_X1 U5162 ( .A1(n5739), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5727) );
  NAND2_X1 U5163 ( .A1(n5743), .A2(n5742), .ZN(n6609) );
  MUX2_X1 U5164 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5741), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5743) );
  NAND2_X1 U5165 ( .A1(n4435), .A2(n4436), .ZN(n8601) );
  AND2_X1 U5166 ( .A1(n4437), .A2(n4794), .ZN(n4436) );
  AOI21_X1 U5167 ( .B1(n4795), .B2(n4439), .A(n4371), .ZN(n4794) );
  NAND2_X1 U5168 ( .A1(n6456), .A2(n4986), .ZN(n6533) );
  NOR2_X1 U5169 ( .A1(n5417), .A2(n8706), .ZN(n4520) );
  OAI211_X1 U5170 ( .C1(n4809), .C2(n4807), .A(n4345), .B(n4803), .ZN(n8659)
         );
  INV_X1 U5171 ( .A(n8730), .ZN(n4807) );
  NAND2_X1 U5172 ( .A1(n8669), .A2(n8670), .ZN(n8668) );
  NAND2_X1 U5173 ( .A1(n6533), .A2(n6534), .ZN(n6584) );
  NAND2_X1 U5174 ( .A1(n5634), .A2(n9028), .ZN(n4939) );
  AND2_X1 U5175 ( .A1(n8610), .A2(n4522), .ZN(n4521) );
  OR2_X1 U5176 ( .A1(n5416), .A2(n4523), .ZN(n4522) );
  INV_X1 U5177 ( .A(n5239), .ZN(n5237) );
  NOR2_X1 U5178 ( .A1(n4801), .A2(n4800), .ZN(n4799) );
  INV_X1 U5179 ( .A(n5490), .ZN(n4801) );
  NAND2_X1 U5180 ( .A1(n5415), .A2(n5416), .ZN(n8704) );
  NAND2_X1 U5181 ( .A1(n5296), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5327) );
  INV_X1 U5182 ( .A(n5298), .ZN(n5296) );
  NAND2_X1 U5183 ( .A1(n4515), .A2(n9005), .ZN(n4514) );
  INV_X1 U5184 ( .A(n4952), .ZN(n4513) );
  OAI22_X1 U5185 ( .A1(n4313), .A2(n6325), .B1(n5013), .B2(n4954), .ZN(n4783)
         );
  NOR2_X2 U5186 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4966) );
  OR2_X1 U5187 ( .A1(n5157), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5202) );
  NOR2_X1 U5188 ( .A1(n6578), .A2(n6577), .ZN(n6846) );
  OR2_X1 U5189 ( .A1(n6851), .A2(n6850), .ZN(n4485) );
  XNOR2_X1 U5190 ( .A(n9043), .B(n9049), .ZN(n7436) );
  AOI21_X1 U5191 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n9083), .A(n9077), .ZN(
        n9915) );
  NAND2_X1 U5192 ( .A1(n8829), .A2(n8828), .ZN(n9099) );
  XNOR2_X1 U5193 ( .A(n9412), .B(n9012), .ZN(n9152) );
  NAND2_X1 U5194 ( .A1(n5574), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5596) );
  INV_X1 U5195 ( .A(n5576), .ZN(n5574) );
  AOI21_X1 U5196 ( .B1(n9219), .B2(n9222), .A(n9123), .ZN(n9205) );
  NOR2_X1 U5197 ( .A1(n9434), .A2(n9014), .ZN(n9123) );
  AND2_X1 U5198 ( .A1(n5603), .A2(n5602), .ZN(n9224) );
  OAI21_X1 U5199 ( .B1(n9248), .B2(n9247), .A(n9145), .ZN(n9235) );
  NOR2_X1 U5200 ( .A1(n9235), .A2(n9236), .ZN(n9234) );
  AOI21_X1 U5201 ( .B1(n9278), .B2(n9144), .A(n9143), .ZN(n9248) );
  OR2_X1 U5202 ( .A1(n5455), .A2(n8690), .ZN(n5475) );
  INV_X1 U5203 ( .A(n9114), .ZN(n9285) );
  NAND2_X1 U5204 ( .A1(n9279), .A2(n4399), .ZN(n9278) );
  AND2_X1 U5205 ( .A1(n9280), .A2(n9303), .ZN(n4399) );
  NAND2_X1 U5206 ( .A1(n9301), .A2(n9142), .ZN(n9279) );
  OAI22_X1 U5207 ( .A1(n9293), .A2(n9113), .B1(n9323), .B2(n9457), .ZN(n9275)
         );
  AND2_X1 U5208 ( .A1(n8865), .A2(n9261), .ZN(n9280) );
  AND3_X1 U5209 ( .A1(n5481), .A2(n5480), .A3(n5479), .ZN(n9306) );
  OR2_X1 U5210 ( .A1(n9457), .A2(n9284), .ZN(n9303) );
  AND2_X1 U5211 ( .A1(n8934), .A2(n8933), .ZN(n9320) );
  NAND2_X1 U5212 ( .A1(n9351), .A2(n9376), .ZN(n4653) );
  NOR2_X1 U5213 ( .A1(n9335), .A2(n4651), .ZN(n4650) );
  INV_X1 U5214 ( .A(n4653), .ZN(n4651) );
  AND2_X1 U5215 ( .A1(n8866), .A2(n9139), .ZN(n9335) );
  OR2_X1 U5216 ( .A1(n5379), .A2(n8672), .ZN(n5404) );
  NAND2_X1 U5217 ( .A1(n4629), .A2(n4627), .ZN(n9357) );
  NAND2_X1 U5218 ( .A1(n9136), .A2(n4628), .ZN(n4627) );
  NAND2_X1 U5219 ( .A1(n8923), .A2(n9137), .ZN(n4628) );
  NAND2_X1 U5220 ( .A1(n9111), .A2(n9110), .ZN(n9346) );
  NAND2_X1 U5221 ( .A1(n9481), .A2(n9385), .ZN(n9110) );
  NAND2_X1 U5222 ( .A1(n9134), .A2(n4631), .ZN(n4630) );
  AND2_X1 U5223 ( .A1(n7555), .A2(n8767), .ZN(n4868) );
  NOR2_X1 U5224 ( .A1(n4661), .A2(n7551), .ZN(n4660) );
  INV_X1 U5225 ( .A(n8879), .ZN(n4661) );
  INV_X1 U5226 ( .A(n4658), .ZN(n4657) );
  OAI22_X1 U5227 ( .A1(n7551), .A2(n4659), .B1(n8771), .B2(n9825), .ZN(n4658)
         );
  INV_X1 U5228 ( .A(n7549), .ZN(n4659) );
  NOR2_X1 U5229 ( .A1(n9760), .A2(n9779), .ZN(n9761) );
  NAND2_X1 U5230 ( .A1(n4411), .A2(n7520), .ZN(n7550) );
  NAND2_X1 U5231 ( .A1(n4664), .A2(n4663), .ZN(n4411) );
  OR2_X1 U5232 ( .A1(n5186), .A2(n6393), .ZN(n5209) );
  NAND2_X1 U5233 ( .A1(n5097), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U5234 ( .A1(n5121), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5162) );
  INV_X1 U5235 ( .A(n5122), .ZN(n5121) );
  NAND2_X1 U5236 ( .A1(n7125), .A2(n7106), .ZN(n7239) );
  NAND2_X1 U5237 ( .A1(n8914), .A2(n4615), .ZN(n4614) );
  INV_X1 U5238 ( .A(n8912), .ZN(n4615) );
  NAND2_X1 U5239 ( .A1(n6806), .A2(n8867), .ZN(n6954) );
  AND2_X1 U5240 ( .A1(n6504), .A2(n6503), .ZN(n9802) );
  NAND2_X1 U5241 ( .A1(n6517), .A2(n4407), .ZN(n4641) );
  XNOR2_X1 U5242 ( .A(n9026), .B(n9403), .ZN(n8872) );
  AND2_X1 U5243 ( .A1(n4512), .A2(n4511), .ZN(n9414) );
  NAND2_X1 U5244 ( .A1(n7117), .A2(n9824), .ZN(n9967) );
  NAND2_X1 U5245 ( .A1(n4617), .A2(n8912), .ZN(n7111) );
  NOR2_X1 U5246 ( .A1(n6943), .A2(n6410), .ZN(n6416) );
  AND2_X1 U5247 ( .A1(n4821), .A2(n4669), .ZN(n4401) );
  AND2_X1 U5248 ( .A1(n4819), .A2(n4901), .ZN(n4669) );
  AND2_X1 U5249 ( .A1(n4366), .A2(n4902), .ZN(n4819) );
  NAND2_X1 U5250 ( .A1(n4913), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4933) );
  AOI21_X1 U5251 ( .B1(n4761), .B2(n4759), .A(n4376), .ZN(n4758) );
  INV_X1 U5252 ( .A(n5469), .ZN(n4759) );
  INV_X1 U5253 ( .A(n5516), .ZN(n4479) );
  NOR2_X1 U5254 ( .A1(n4760), .A2(n4757), .ZN(n4756) );
  INV_X1 U5255 ( .A(n5448), .ZN(n4757) );
  INV_X1 U5256 ( .A(n4761), .ZN(n4760) );
  NAND2_X1 U5257 ( .A1(n4481), .A2(n4770), .ZN(n5446) );
  NAND2_X1 U5258 ( .A1(n4470), .A2(n5259), .ZN(n5286) );
  NAND2_X1 U5259 ( .A1(n4471), .A2(n4462), .ZN(n4470) );
  INV_X1 U5260 ( .A(n4464), .ZN(n4462) );
  NAND2_X1 U5261 ( .A1(n4471), .A2(n5228), .ZN(n5258) );
  XNOR2_X1 U5262 ( .A(n5177), .B(n5176), .ZN(n6273) );
  OAI21_X1 U5263 ( .B1(n4453), .B2(n4454), .A(n5149), .ZN(n5177) );
  NAND2_X1 U5264 ( .A1(n4568), .A2(n4457), .ZN(n4454) );
  NAND2_X1 U5265 ( .A1(n5083), .A2(n5082), .ZN(n5107) );
  NAND2_X1 U5266 ( .A1(n5027), .A2(n5026), .ZN(n5059) );
  XNOR2_X1 U5267 ( .A(n4961), .B(n4946), .ZN(n4960) );
  NAND2_X1 U5268 ( .A1(n5745), .A2(n5744), .ZN(n8484) );
  AND4_X1 U5269 ( .A1(n5767), .A2(n5766), .A3(n5765), .A4(n5764), .ZN(n8414)
         );
  AND3_X1 U5270 ( .A1(n6044), .A2(n6043), .A3(n6042), .ZN(n8258) );
  NAND2_X1 U5271 ( .A1(n6038), .A2(n6037), .ZN(n8479) );
  NOR2_X1 U5272 ( .A1(n6790), .A2(n4741), .ZN(n4740) );
  NAND2_X1 U5273 ( .A1(n6795), .A2(n6796), .ZN(n6857) );
  INV_X1 U5274 ( .A(n7810), .ZN(n7789) );
  AND2_X1 U5275 ( .A1(n6560), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7794) );
  AND2_X1 U5276 ( .A1(n6599), .A2(n10000), .ZN(n9994) );
  AND2_X1 U5277 ( .A1(n8020), .A2(n7833), .ZN(n8024) );
  NAND2_X1 U5278 ( .A1(n4591), .A2(n4590), .ZN(n4589) );
  OR2_X1 U5279 ( .A1(n8018), .A2(n8019), .ZN(n4590) );
  OAI21_X1 U5280 ( .B1(n8021), .B2(n8022), .A(n8020), .ZN(n4591) );
  XNOR2_X1 U5281 ( .A(n6124), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8027) );
  INV_X1 U5282 ( .A(n7467), .ZN(n8041) );
  NAND2_X1 U5283 ( .A1(n7830), .A2(n7829), .ZN(n9749) );
  XNOR2_X1 U5284 ( .A(n4314), .B(n9749), .ZN(n9747) );
  XNOR2_X1 U5285 ( .A(n6111), .B(n6110), .ZN(n8458) );
  OR2_X1 U5286 ( .A1(n8459), .A2(n8032), .ZN(n6094) );
  AND2_X1 U5287 ( .A1(n6085), .A2(n6061), .ZN(n8214) );
  AND2_X1 U5288 ( .A1(n5722), .A2(n4847), .ZN(n4846) );
  INV_X1 U5289 ( .A(n4795), .ZN(n4524) );
  NAND2_X1 U5290 ( .A1(n8619), .A2(n8618), .ZN(n9421) );
  NOR2_X1 U5291 ( .A1(n5638), .A2(n5637), .ZN(n4449) );
  XNOR2_X1 U5292 ( .A(n4956), .B(n5031), .ZN(n6424) );
  OAI21_X1 U5293 ( .B1(n8969), .B2(n4952), .A(n4955), .ZN(n4956) );
  NAND2_X1 U5294 ( .A1(n4441), .A2(n8688), .ZN(n8646) );
  NAND2_X1 U5295 ( .A1(n8686), .A2(n8687), .ZN(n4441) );
  INV_X1 U5296 ( .A(n9299), .ZN(n9457) );
  NAND2_X1 U5297 ( .A1(n6364), .A2(n5667), .ZN(n8726) );
  AND2_X1 U5298 ( .A1(n5664), .A2(n9961), .ZN(n8717) );
  NAND2_X1 U5299 ( .A1(n5325), .A2(n5324), .ZN(n9393) );
  AND2_X1 U5300 ( .A1(n6231), .A2(n6507), .ZN(n9921) );
  OAI21_X1 U5301 ( .B1(n9088), .B2(n9087), .A(n4497), .ZN(n4496) );
  AOI21_X1 U5302 ( .B1(n9089), .B2(n9920), .A(n9912), .ZN(n4497) );
  NAND2_X1 U5303 ( .A1(n4638), .A2(n4637), .ZN(n9419) );
  INV_X1 U5304 ( .A(n9178), .ZN(n4637) );
  NAND2_X1 U5305 ( .A1(n4640), .A2(n4639), .ZN(n4638) );
  AND2_X1 U5306 ( .A1(n9172), .A2(n9173), .ZN(n9418) );
  AND2_X1 U5307 ( .A1(n5595), .A2(n5594), .ZN(n9216) );
  AND2_X1 U5308 ( .A1(n5523), .A2(n5522), .ZN(n9257) );
  NOR2_X1 U5309 ( .A1(n7912), .A2(n7911), .ZN(n7919) );
  AND2_X1 U5310 ( .A1(n7928), .A2(n7924), .ZN(n4582) );
  NOR2_X1 U5311 ( .A1(n6171), .A2(n8012), .ZN(n4580) );
  NAND2_X1 U5312 ( .A1(n4585), .A2(n4584), .ZN(n4583) );
  NOR2_X1 U5313 ( .A1(n6171), .A2(n4682), .ZN(n4586) );
  AND2_X1 U5314 ( .A1(n8352), .A2(n7946), .ZN(n4395) );
  AOI21_X1 U5315 ( .B1(n7957), .B2(n7956), .A(n6174), .ZN(n4562) );
  AND2_X1 U5316 ( .A1(n7965), .A2(n7966), .ZN(n4394) );
  NAND2_X1 U5317 ( .A1(n4577), .A2(n4576), .ZN(n4575) );
  NAND2_X1 U5318 ( .A1(n4354), .A2(n8000), .ZN(n4576) );
  OAI21_X1 U5319 ( .B1(n7971), .B2(n4578), .A(n8261), .ZN(n4577) );
  INV_X1 U5320 ( .A(n8224), .ZN(n4572) );
  NAND2_X1 U5321 ( .A1(n7979), .A2(n8012), .ZN(n4571) );
  AOI21_X1 U5322 ( .B1(n4574), .B2(n4573), .A(n4570), .ZN(n7989) );
  NAND2_X1 U5323 ( .A1(n7977), .A2(n8012), .ZN(n4573) );
  NAND2_X1 U5324 ( .A1(n4572), .A2(n4571), .ZN(n4570) );
  NAND2_X1 U5325 ( .A1(n4575), .A2(n7978), .ZN(n4574) );
  OR2_X1 U5326 ( .A1(n8455), .A2(n7672), .ZN(n8004) );
  NAND2_X1 U5327 ( .A1(n4328), .A2(n4748), .ZN(n8851) );
  INV_X1 U5328 ( .A(n9743), .ZN(n4748) );
  OR2_X1 U5329 ( .A1(n9422), .A2(n9210), .ZN(n8945) );
  NOR2_X1 U5330 ( .A1(n9421), .A2(n9422), .ZN(n4510) );
  OR2_X1 U5331 ( .A1(n4509), .A2(n9449), .ZN(n4508) );
  NAND2_X1 U5332 ( .A1(n9290), .A2(n9257), .ZN(n4509) );
  INV_X1 U5333 ( .A(SI_30_), .ZN(n4779) );
  INV_X1 U5334 ( .A(n5540), .ZN(n4774) );
  INV_X1 U5335 ( .A(n5564), .ZN(n4776) );
  NOR2_X1 U5336 ( .A1(n4899), .A2(n4898), .ZN(n4900) );
  NAND2_X1 U5337 ( .A1(n5344), .A2(n5343), .ZN(n5370) );
  NAND2_X1 U5338 ( .A1(n5318), .A2(n9602), .ZN(n5341) );
  INV_X1 U5339 ( .A(n5285), .ZN(n4469) );
  INV_X1 U5340 ( .A(n4466), .ZN(n4461) );
  AOI21_X1 U5341 ( .B1(n5285), .B2(n4468), .A(n4467), .ZN(n4466) );
  INV_X1 U5342 ( .A(n5259), .ZN(n4468) );
  INV_X1 U5343 ( .A(n5287), .ZN(n4467) );
  INV_X1 U5344 ( .A(n5149), .ZN(n4455) );
  INV_X1 U5345 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4927) );
  INV_X1 U5346 ( .A(SI_9_), .ZN(n9705) );
  INV_X1 U5347 ( .A(n4738), .ZN(n4735) );
  NAND2_X1 U5348 ( .A1(n8006), .A2(n7837), .ZN(n4398) );
  OR2_X1 U5349 ( .A1(n5801), .A2(n6619), .ZN(n5772) );
  NAND2_X1 U5350 ( .A1(n8004), .A2(n8005), .ZN(n7996) );
  AOI21_X1 U5351 ( .B1(n4696), .B2(n4695), .A(n4350), .ZN(n4694) );
  INV_X1 U5352 ( .A(n6175), .ZN(n4695) );
  OR2_X1 U5353 ( .A1(n5971), .A2(n9661), .ZN(n5985) );
  OR2_X1 U5354 ( .A1(n5941), .A2(n5701), .ZN(n5957) );
  NAND2_X1 U5355 ( .A1(n4852), .A2(n4851), .ZN(n4850) );
  INV_X1 U5356 ( .A(n4855), .ZN(n4851) );
  AND2_X1 U5357 ( .A1(n7934), .A2(n7935), .ZN(n7932) );
  INV_X1 U5358 ( .A(n10046), .ZN(n4596) );
  NOR2_X1 U5359 ( .A1(n8555), .A2(n7386), .ZN(n4597) );
  NOR2_X1 U5360 ( .A1(n5878), .A2(n4708), .ZN(n4712) );
  INV_X1 U5361 ( .A(n7899), .ZN(n4708) );
  NAND2_X1 U5362 ( .A1(n8048), .A2(n10009), .ZN(n7869) );
  NAND2_X1 U5363 ( .A1(n7183), .A2(n10001), .ZN(n6435) );
  NOR2_X1 U5364 ( .A1(n8402), .A2(n4602), .ZN(n8377) );
  AND2_X1 U5365 ( .A1(n6599), .A2(n6132), .ZN(n6471) );
  INV_X1 U5366 ( .A(n7384), .ZN(n6135) );
  INV_X1 U5367 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4606) );
  INV_X1 U5368 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5720) );
  INV_X1 U5369 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6138) );
  OR2_X1 U5370 ( .A1(n5908), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5920) );
  NAND2_X1 U5371 ( .A1(n5835), .A2(n5709), .ZN(n5860) );
  INV_X1 U5372 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5708) );
  INV_X1 U5373 ( .A(n4529), .ZN(n4528) );
  OAI21_X1 U5374 ( .B1(n4530), .B2(n4323), .A(n5311), .ZN(n4529) );
  AND2_X1 U5375 ( .A1(n8647), .A2(n4443), .ZN(n4442) );
  NAND2_X1 U5376 ( .A1(n8688), .A2(n4444), .ZN(n4443) );
  INV_X1 U5377 ( .A(n8687), .ZN(n4444) );
  NAND2_X1 U5378 ( .A1(n4438), .A2(n4445), .ZN(n4437) );
  OR2_X1 U5379 ( .A1(n5338), .A2(n8730), .ZN(n4804) );
  AND2_X1 U5380 ( .A1(n4526), .A2(n8661), .ZN(n4525) );
  NAND2_X1 U5381 ( .A1(n4331), .A2(n4530), .ZN(n4526) );
  INV_X1 U5382 ( .A(n8851), .ZN(n8959) );
  OR2_X1 U5383 ( .A1(n9099), .A2(n8859), .ZN(n8993) );
  AND2_X1 U5384 ( .A1(n4485), .A2(n4484), .ZN(n7433) );
  NAND2_X1 U5385 ( .A1(n7199), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4484) );
  NOR2_X1 U5386 ( .A1(n9176), .A2(n9175), .ZN(n9174) );
  AND2_X1 U5387 ( .A1(n8945), .A2(n8949), .ZN(n9128) );
  OR2_X1 U5388 ( .A1(n9454), .A2(n9306), .ZN(n8865) );
  AND2_X1 U5389 ( .A1(n8919), .A2(n8918), .ZN(n4634) );
  INV_X1 U5390 ( .A(n7238), .ZN(n8874) );
  NAND2_X1 U5391 ( .A1(n9949), .A2(n9021), .ZN(n8974) );
  NOR2_X1 U5392 ( .A1(n8911), .A2(n4619), .ZN(n4618) );
  NAND2_X1 U5393 ( .A1(n9211), .A2(n4510), .ZN(n9179) );
  NOR3_X1 U5394 ( .A1(n9294), .A2(n9449), .A3(n9454), .ZN(n9266) );
  NOR2_X1 U5395 ( .A1(n9294), .A2(n9454), .ZN(n9286) );
  NAND2_X1 U5396 ( .A1(n4515), .A2(n9161), .ZN(n8850) );
  INV_X1 U5397 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4820) );
  NAND2_X1 U5398 ( .A1(n7822), .A2(n4779), .ZN(n4778) );
  INV_X1 U5399 ( .A(n6078), .ZN(n4754) );
  AND2_X1 U5400 ( .A1(n5615), .A2(n5593), .ZN(n5613) );
  NAND2_X1 U5401 ( .A1(n5371), .A2(n4482), .ZN(n4481) );
  NOR2_X1 U5402 ( .A1(n4772), .A2(n4483), .ZN(n4482) );
  INV_X1 U5403 ( .A(n5370), .ZN(n4483) );
  INV_X1 U5404 ( .A(n4771), .ZN(n4770) );
  OAI21_X1 U5405 ( .B1(n4772), .B2(n5395), .A(n5422), .ZN(n4771) );
  AND2_X1 U5406 ( .A1(n4883), .A2(n4893), .ZN(n4447) );
  NOR2_X1 U5407 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4883) );
  OAI21_X1 U5408 ( .B1(n5340), .B2(n5339), .A(n5341), .ZN(n5369) );
  INV_X1 U5409 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U5410 ( .A1(n5230), .A2(n9652), .ZN(n5259) );
  NAND2_X1 U5411 ( .A1(n4465), .A2(n5228), .ZN(n4464) );
  INV_X1 U5412 ( .A(n5257), .ZN(n4465) );
  OR2_X1 U5413 ( .A1(n5226), .A2(n5225), .ZN(n4471) );
  INV_X1 U5414 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5154) );
  INV_X1 U5415 ( .A(n5148), .ZN(n4457) );
  AND2_X1 U5416 ( .A1(n5129), .A2(n5106), .ZN(n4567) );
  AOI21_X1 U5417 ( .B1(n4569), .B2(n5129), .A(n4346), .ZN(n4568) );
  INV_X1 U5418 ( .A(n5109), .ZN(n4569) );
  INV_X1 U5419 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4878) );
  INV_X1 U5420 ( .A(SI_21_), .ZN(n9646) );
  NAND2_X1 U5421 ( .A1(n4731), .A2(n7603), .ZN(n7699) );
  INV_X1 U5422 ( .A(n7701), .ZN(n4731) );
  OR2_X1 U5423 ( .A1(n7395), .A2(n7394), .ZN(n4718) );
  AND2_X1 U5424 ( .A1(n7675), .A2(n7671), .ZN(n7693) );
  INV_X1 U5425 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5880) );
  NAND2_X1 U5426 ( .A1(n7621), .A2(n4747), .ZN(n7718) );
  AND2_X1 U5427 ( .A1(n7627), .A2(n7620), .ZN(n4747) );
  INV_X1 U5428 ( .A(n7720), .ZN(n7627) );
  OR2_X1 U5429 ( .A1(n5897), .A2(n9604), .ZN(n5925) );
  INV_X1 U5430 ( .A(n6556), .ZN(n4741) );
  NAND2_X1 U5431 ( .A1(n7699), .A2(n7604), .ZN(n7743) );
  OR2_X1 U5432 ( .A1(n6470), .A2(n6466), .ZN(n6492) );
  NAND2_X1 U5433 ( .A1(n8068), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4536) );
  NOR2_X1 U5434 ( .A1(n8082), .A2(n4543), .ZN(n6738) );
  AND2_X1 U5435 ( .A1(n8081), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4543) );
  NOR2_X1 U5436 ( .A1(n6738), .A2(n6737), .ZN(n6828) );
  NOR2_X1 U5437 ( .A1(n6828), .A2(n4542), .ZN(n6830) );
  AND2_X1 U5438 ( .A1(n6829), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4542) );
  NAND2_X1 U5439 ( .A1(n6830), .A2(n6831), .ZN(n6900) );
  NOR2_X1 U5440 ( .A1(n8127), .A2(n4389), .ZN(n8131) );
  INV_X1 U5441 ( .A(n6598), .ZN(n6490) );
  NAND2_X1 U5442 ( .A1(n8131), .A2(n8130), .ZN(n8144) );
  NAND2_X1 U5443 ( .A1(n8198), .A2(n7992), .ZN(n8179) );
  NAND2_X1 U5444 ( .A1(n4418), .A2(n6075), .ZN(n4417) );
  NAND2_X1 U5445 ( .A1(n8193), .A2(n7987), .ZN(n8198) );
  AND2_X1 U5446 ( .A1(n4458), .A2(n7985), .ZN(n8193) );
  OR2_X1 U5447 ( .A1(n8174), .A2(n6087), .ZN(n6093) );
  OR2_X1 U5448 ( .A1(n8211), .A2(n8464), .ZN(n4877) );
  OR2_X1 U5449 ( .A1(n6060), .A2(n6059), .ZN(n6085) );
  NAND2_X1 U5450 ( .A1(n8221), .A2(n8224), .ZN(n8220) );
  CLKBUF_X1 U5451 ( .A(n8252), .Z(n8253) );
  OR2_X1 U5452 ( .A1(n4609), .A2(n8484), .ZN(n4608) );
  OR2_X1 U5453 ( .A1(n6028), .A2(n9606), .ZN(n6030) );
  NAND2_X1 U5454 ( .A1(n4561), .A2(n4560), .ZN(n7966) );
  NAND2_X1 U5455 ( .A1(n8324), .A2(n6175), .ZN(n4699) );
  NAND2_X1 U5456 ( .A1(n4699), .A2(n4696), .ZN(n8296) );
  NOR3_X1 U5457 ( .A1(n8306), .A2(n8499), .A3(n8504), .ZN(n8291) );
  NOR2_X1 U5458 ( .A1(n8306), .A2(n8504), .ZN(n8305) );
  INV_X1 U5459 ( .A(n4829), .ZN(n4828) );
  NOR2_X1 U5460 ( .A1(n8402), .A2(n4601), .ZN(n8356) );
  NOR2_X1 U5461 ( .A1(n4601), .A2(n8514), .ZN(n4600) );
  AND2_X1 U5462 ( .A1(n7956), .A2(n7955), .ZN(n8339) );
  AOI21_X1 U5463 ( .B1(n4692), .B2(n8391), .A(n4690), .ZN(n4689) );
  INV_X1 U5464 ( .A(n7944), .ZN(n4690) );
  NAND2_X1 U5465 ( .A1(n8395), .A2(n7940), .ZN(n8368) );
  NAND2_X1 U5466 ( .A1(n8390), .A2(n7937), .ZN(n8395) );
  NAND2_X1 U5467 ( .A1(n8416), .A2(n7934), .ZN(n8390) );
  NAND2_X1 U5468 ( .A1(n4676), .A2(n4674), .ZN(n8412) );
  AND2_X1 U5469 ( .A1(n4675), .A2(n7930), .ZN(n4674) );
  AND2_X1 U5470 ( .A1(n7355), .A2(n4593), .ZN(n8445) );
  NOR2_X1 U5471 ( .A1(n8449), .A2(n4595), .ZN(n4593) );
  AND4_X1 U5472 ( .A1(n5932), .A2(n5931), .A3(n5930), .A4(n5929), .ZN(n8432)
         );
  NAND2_X1 U5473 ( .A1(n4673), .A2(n4677), .ZN(n8429) );
  OR2_X1 U5474 ( .A1(n6169), .A2(n4680), .ZN(n4673) );
  NAND2_X1 U5475 ( .A1(n7355), .A2(n4597), .ZN(n7460) );
  NAND2_X1 U5476 ( .A1(n7355), .A2(n10039), .ZN(n7357) );
  AND2_X1 U5477 ( .A1(n7256), .A2(n5879), .ZN(n7310) );
  NAND2_X1 U5478 ( .A1(n4837), .A2(n4840), .ZN(n4835) );
  OR2_X1 U5479 ( .A1(n7260), .A2(n7263), .ZN(n7317) );
  NAND2_X1 U5480 ( .A1(n4713), .A2(n7899), .ZN(n7253) );
  OAI21_X1 U5481 ( .B1(n7278), .B2(n6164), .A(n7883), .ZN(n7023) );
  NOR2_X1 U5482 ( .A1(n7171), .A2(n7176), .ZN(n7273) );
  AND2_X1 U5483 ( .A1(n7273), .A2(n10019), .ZN(n7271) );
  AND4_X1 U5484 ( .A1(n5805), .A2(n5804), .A3(n5803), .A4(n5802), .ZN(n7165)
         );
  NAND2_X1 U5485 ( .A1(n7889), .A2(n7881), .ZN(n7840) );
  NAND2_X1 U5486 ( .A1(n5779), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5791) );
  AND4_X1 U5487 ( .A1(n5820), .A2(n5819), .A3(n5818), .A4(n5817), .ZN(n6771)
         );
  INV_X1 U5488 ( .A(n8430), .ZN(n8343) );
  NAND2_X1 U5489 ( .A1(n7159), .A2(n7839), .ZN(n7158) );
  OR2_X1 U5490 ( .A1(n10050), .A2(n7833), .ZN(n6469) );
  OR2_X1 U5491 ( .A1(n6262), .A2(n5864), .ZN(n4430) );
  INV_X1 U5492 ( .A(n7176), .ZN(n10014) );
  OAI211_X1 U5493 ( .C1(n5864), .C2(n6249), .A(n5811), .B(n5810), .ZN(n6777)
         );
  AND2_X1 U5494 ( .A1(n9992), .A2(n9995), .ZN(n6137) );
  INV_X1 U5495 ( .A(n7511), .ZN(n6133) );
  INV_X1 U5496 ( .A(n5742), .ZN(n5737) );
  OR2_X1 U5497 ( .A1(n6125), .A2(n8588), .ZN(n6126) );
  INV_X1 U5498 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U5499 ( .A1(n6112), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6128) );
  AND2_X1 U5500 ( .A1(n5835), .A2(n4358), .ZN(n5951) );
  INV_X1 U5501 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5952) );
  OR2_X1 U5502 ( .A1(n5904), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U5503 ( .A1(n5836), .A2(n4746), .ZN(n5746) );
  CLKBUF_X1 U5504 ( .A(n5835), .Z(n5836) );
  NAND2_X1 U5505 ( .A1(n5708), .A2(n4861), .ZN(n4860) );
  INV_X1 U5506 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4861) );
  NAND2_X1 U5507 ( .A1(n4448), .A2(n4528), .ZN(n7569) );
  NAND2_X1 U5508 ( .A1(n7475), .A2(n7473), .ZN(n4448) );
  NAND2_X1 U5509 ( .A1(n4798), .A2(n5489), .ZN(n4795) );
  NAND2_X1 U5510 ( .A1(n8697), .A2(n5514), .ZN(n4798) );
  AND2_X1 U5511 ( .A1(n5612), .A2(n5611), .ZN(n5637) );
  NAND2_X1 U5512 ( .A1(n5207), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5239) );
  INV_X1 U5513 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5161) );
  NAND2_X1 U5514 ( .A1(n5606), .A2(n9028), .ZN(n4937) );
  INV_X1 U5515 ( .A(n5432), .ZN(n5430) );
  INV_X1 U5516 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5268) );
  OR2_X1 U5517 ( .A1(n5269), .A2(n5268), .ZN(n5298) );
  NAND2_X1 U5518 ( .A1(n4813), .A2(n5069), .ZN(n4811) );
  NAND2_X1 U5519 ( .A1(n4792), .A2(n4793), .ZN(n4789) );
  NAND2_X1 U5520 ( .A1(n4792), .A2(n5562), .ZN(n4788) );
  OR2_X1 U5521 ( .A1(n8894), .A2(n8890), .ZN(n4767) );
  AND4_X1 U5522 ( .A1(n5244), .A2(n5243), .A3(n5242), .A4(n5241), .ZN(n9797)
         );
  NAND2_X1 U5523 ( .A1(n6380), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4486) );
  NOR2_X1 U5524 ( .A1(n6356), .A2(n4330), .ZN(n6355) );
  AOI21_X1 U5525 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n6359), .A(n6355), .ZN(
        n9855) );
  NOR2_X1 U5526 ( .A1(n9886), .A2(n4488), .ZN(n6334) );
  NOR2_X1 U5527 ( .A1(n6257), .A2(n7134), .ZN(n4488) );
  NAND2_X1 U5528 ( .A1(n6334), .A2(n6335), .ZN(n6333) );
  AOI21_X1 U5529 ( .B1(n6400), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6394), .ZN(
        n6397) );
  NOR2_X1 U5530 ( .A1(n6573), .A2(n4493), .ZN(n9030) );
  AND2_X1 U5531 ( .A1(n6574), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4493) );
  NAND2_X1 U5532 ( .A1(n9030), .A2(n9031), .ZN(n9029) );
  NAND2_X1 U5533 ( .A1(n9029), .A2(n4492), .ZN(n6578) );
  OR2_X1 U5534 ( .A1(n6575), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4492) );
  AND2_X1 U5535 ( .A1(n5264), .A2(n4893), .ZN(n5289) );
  XNOR2_X1 U5536 ( .A(n7433), .B(n7432), .ZN(n7201) );
  NOR2_X1 U5537 ( .A1(n7201), .A2(n7200), .ZN(n7434) );
  NOR2_X1 U5538 ( .A1(n7436), .A2(n9391), .ZN(n9044) );
  INV_X1 U5539 ( .A(n9174), .ZN(n4640) );
  OAI21_X1 U5540 ( .B1(n9235), .B2(n4623), .A(n4620), .ZN(n9190) );
  AOI21_X1 U5541 ( .B1(n4622), .B2(n9146), .A(n4621), .ZN(n4620) );
  INV_X1 U5542 ( .A(n9147), .ZN(n4621) );
  NOR2_X1 U5543 ( .A1(n9190), .A2(n9191), .ZN(n9189) );
  AND2_X1 U5544 ( .A1(n5689), .A2(n5688), .ZN(n9192) );
  NAND2_X1 U5545 ( .A1(n9127), .A2(n9126), .ZN(n9188) );
  NAND2_X1 U5546 ( .A1(n9439), .A2(n9120), .ZN(n9119) );
  NAND2_X1 U5547 ( .A1(n8946), .A2(n8861), .ZN(n9222) );
  INV_X1 U5548 ( .A(n4666), .ZN(n4665) );
  OAI21_X1 U5549 ( .B1(n4667), .B2(n4872), .A(n4871), .ZN(n4666) );
  AND2_X1 U5550 ( .A1(n5533), .A2(n5532), .ZN(n9265) );
  OR2_X1 U5551 ( .A1(n5475), .A2(n5474), .ZN(n5502) );
  NAND2_X1 U5552 ( .A1(n4408), .A2(n4642), .ZN(n9293) );
  AOI21_X1 U5553 ( .B1(n4644), .B2(n4647), .A(n4353), .ZN(n4642) );
  NAND2_X1 U5554 ( .A1(n9346), .A2(n4644), .ZN(n4408) );
  AND2_X1 U5555 ( .A1(n9303), .A2(n9142), .ZN(n9300) );
  OAI21_X1 U5556 ( .B1(n9330), .B2(n9140), .A(n9139), .ZN(n9321) );
  NOR2_X2 U5557 ( .A1(n9349), .A2(n9468), .ZN(n9338) );
  INV_X1 U5558 ( .A(n5353), .ZN(n5351) );
  OR2_X1 U5559 ( .A1(n5327), .A2(n5326), .ZN(n5353) );
  NOR2_X1 U5560 ( .A1(n4503), .A2(n9481), .ZN(n4501) );
  NOR2_X1 U5561 ( .A1(n9760), .A2(n4505), .ZN(n9388) );
  NAND2_X1 U5562 ( .A1(n4357), .A2(n4315), .ZN(n4654) );
  NAND2_X1 U5563 ( .A1(n4412), .A2(n4414), .ZN(n4409) );
  NAND2_X1 U5564 ( .A1(n4664), .A2(n4412), .ZN(n4410) );
  INV_X1 U5565 ( .A(n7556), .ZN(n7557) );
  OR2_X1 U5566 ( .A1(n5162), .A2(n5161), .ZN(n5186) );
  NAND2_X1 U5567 ( .A1(n4633), .A2(n8898), .ZN(n7513) );
  AND2_X1 U5568 ( .A1(n7338), .A2(n7372), .ZN(n9783) );
  NAND2_X1 U5569 ( .A1(n7113), .A2(n4634), .ZN(n7329) );
  AND2_X1 U5570 ( .A1(n8762), .A2(n8759), .ZN(n8876) );
  AND2_X1 U5571 ( .A1(n7108), .A2(n7107), .ZN(n4662) );
  AND2_X1 U5572 ( .A1(n8919), .A2(n8758), .ZN(n8875) );
  NAND2_X1 U5573 ( .A1(n7113), .A2(n8918), .ZN(n7284) );
  NOR2_X1 U5574 ( .A1(n7135), .A2(n7139), .ZN(n7241) );
  NAND2_X1 U5575 ( .A1(n9949), .A2(n7241), .ZN(n7240) );
  AND4_X1 U5576 ( .A1(n5128), .A2(n5127), .A3(n5126), .A4(n5125), .ZN(n7287)
         );
  NAND2_X1 U5577 ( .A1(n7239), .A2(n7238), .ZN(n7237) );
  INV_X1 U5578 ( .A(n7127), .ZN(n7105) );
  AND2_X1 U5579 ( .A1(n8915), .A2(n8967), .ZN(n7127) );
  NAND2_X1 U5580 ( .A1(n4498), .A2(n6968), .ZN(n7135) );
  AND4_X1 U5581 ( .A1(n4993), .A2(n4992), .A3(n4991), .A4(n4990), .ZN(n6807)
         );
  NAND2_X1 U5582 ( .A1(n7044), .A2(n8910), .ZN(n6959) );
  AND4_X1 U5583 ( .A1(n5051), .A2(n5050), .A3(n5049), .A4(n5048), .ZN(n7129)
         );
  NOR2_X1 U5584 ( .A1(n6525), .A2(n6810), .ZN(n7051) );
  AND2_X1 U5585 ( .A1(n8890), .A2(n6507), .ZN(n9772) );
  AND2_X1 U5586 ( .A1(n9028), .A2(n7019), .ZN(n6502) );
  OR2_X1 U5587 ( .A1(n5022), .A2(n6243), .ZN(n4951) );
  NAND2_X1 U5588 ( .A1(n4949), .A2(n4336), .ZN(n4499) );
  AND2_X1 U5589 ( .A1(n6499), .A2(n6498), .ZN(n7117) );
  INV_X1 U5590 ( .A(n9216), .ZN(n9429) );
  INV_X1 U5591 ( .A(n9393), .ZN(n9818) );
  NAND2_X1 U5592 ( .A1(n5185), .A2(n5184), .ZN(n9735) );
  OR2_X1 U5593 ( .A1(n7017), .A2(n9002), .ZN(n9963) );
  NAND2_X1 U5594 ( .A1(n4641), .A2(n6804), .ZN(n7041) );
  INV_X1 U5595 ( .A(n9935), .ZN(n9961) );
  AND2_X1 U5596 ( .A1(n6413), .A2(n7016), .ZN(n9935) );
  NAND2_X1 U5597 ( .A1(n4515), .A2(n6948), .ZN(n7017) );
  OAI211_X1 U5598 ( .C1(P1_B_REG_SCAN_IN), .C2(n7364), .A(n5646), .B(n5642), 
        .ZN(n9504) );
  XNOR2_X1 U5599 ( .A(n7823), .B(n7586), .ZN(n8826) );
  NAND2_X1 U5600 ( .A1(n4912), .A2(n4870), .ZN(n4919) );
  XNOR2_X1 U5601 ( .A(n7583), .B(n6100), .ZN(n8841) );
  XNOR2_X1 U5602 ( .A(n6077), .B(n6076), .ZN(n7543) );
  AND2_X1 U5603 ( .A1(n4909), .A2(n4335), .ZN(n5643) );
  INV_X1 U5604 ( .A(n4476), .ZN(n4472) );
  NAND2_X1 U5605 ( .A1(n4763), .A2(n5471), .ZN(n5494) );
  NAND2_X1 U5606 ( .A1(n5470), .A2(n5469), .ZN(n4763) );
  XNOR2_X1 U5607 ( .A(n5198), .B(n5197), .ZN(n6278) );
  NAND2_X1 U5608 ( .A1(n4429), .A2(n5061), .ZN(n5080) );
  XNOR2_X1 U5609 ( .A(n5081), .B(n9649), .ZN(n5079) );
  NAND2_X1 U5610 ( .A1(n5004), .A2(n5003), .ZN(n5024) );
  OR2_X1 U5611 ( .A1(n4966), .A2(n9507), .ZN(n4995) );
  AOI21_X1 U5612 ( .B1(n9881), .B2(n9527), .A(n10111), .ZN(n9528) );
  NAND2_X1 U5613 ( .A1(n5753), .A2(n5752), .ZN(n8538) );
  NAND2_X1 U5614 ( .A1(n4718), .A2(n7393), .ZN(n7397) );
  NAND2_X1 U5615 ( .A1(n7621), .A2(n7620), .ZN(n7721) );
  NAND2_X1 U5616 ( .A1(n5995), .A2(n5994), .ZN(n8510) );
  NAND2_X1 U5617 ( .A1(n6080), .A2(n6079), .ZN(n8459) );
  INV_X1 U5618 ( .A(n4722), .ZN(n4721) );
  AOI21_X1 U5619 ( .B1(n4720), .B2(n4722), .A(n4352), .ZN(n4719) );
  AND2_X1 U5620 ( .A1(n4723), .A2(n6856), .ZN(n4722) );
  AND4_X1 U5621 ( .A1(n5977), .A2(n5976), .A3(n5975), .A4(n5974), .ZN(n8369)
         );
  AND4_X1 U5622 ( .A1(n5962), .A2(n5961), .A3(n5960), .A4(n5959), .ZN(n8393)
         );
  AND2_X1 U5623 ( .A1(n4728), .A2(n7610), .ZN(n4727) );
  NAND2_X1 U5624 ( .A1(n5894), .A2(n5893), .ZN(n8559) );
  NAND2_X1 U5625 ( .A1(n4716), .A2(n4714), .ZN(n7406) );
  AOI21_X1 U5626 ( .B1(n4717), .B2(n7394), .A(n4715), .ZN(n4714) );
  INV_X1 U5627 ( .A(n7404), .ZN(n4715) );
  AND4_X1 U5628 ( .A1(n6004), .A2(n6003), .A3(n6002), .A4(n6001), .ZN(n7785)
         );
  INV_X1 U5629 ( .A(n7793), .ZN(n7803) );
  NAND2_X1 U5630 ( .A1(n6058), .A2(n6057), .ZN(n8471) );
  NAND2_X1 U5631 ( .A1(n4732), .A2(n4737), .ZN(n7792) );
  NAND2_X1 U5632 ( .A1(n7737), .A2(n4738), .ZN(n4732) );
  AND4_X1 U5633 ( .A1(n5759), .A2(n5758), .A3(n5757), .A4(n5756), .ZN(n8431)
         );
  INV_X1 U5634 ( .A(n7795), .ZN(n7806) );
  NAND2_X1 U5635 ( .A1(n5938), .A2(n5937), .ZN(n8533) );
  INV_X1 U5636 ( .A(n7785), .ZN(n8344) );
  INV_X1 U5637 ( .A(n7313), .ZN(n8043) );
  INV_X1 U5638 ( .A(n6772), .ZN(n8048) );
  INV_X1 U5639 ( .A(n4541), .ZN(n6678) );
  NOR2_X1 U5640 ( .A1(n6681), .A2(n6680), .ZN(n6695) );
  AND2_X1 U5641 ( .A1(n4541), .A2(n4540), .ZN(n6681) );
  NAND2_X1 U5642 ( .A1(n6683), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4540) );
  INV_X1 U5643 ( .A(n4539), .ZN(n8055) );
  INV_X1 U5644 ( .A(n4537), .ZN(n8069) );
  AOI21_X1 U5645 ( .B1(n4551), .B2(n4547), .A(n4553), .ZN(n4546) );
  AND2_X1 U5646 ( .A1(n6615), .A2(n6605), .ZN(n8150) );
  XNOR2_X1 U5647 ( .A(n4544), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8146) );
  NAND2_X1 U5648 ( .A1(n8144), .A2(n4545), .ZN(n4544) );
  OR2_X1 U5649 ( .A1(n8145), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4545) );
  AND2_X1 U5650 ( .A1(n6617), .A2(n6616), .ZN(n9986) );
  OAI21_X1 U5651 ( .B1(n8221), .B2(n4325), .A(n4419), .ZN(n8186) );
  NAND2_X1 U5652 ( .A1(n8203), .A2(n6066), .ZN(n8187) );
  INV_X1 U5653 ( .A(n8440), .ZN(n8404) );
  NAND2_X1 U5654 ( .A1(n4702), .A2(n4703), .ZN(n8207) );
  INV_X1 U5655 ( .A(n4458), .ZN(n8206) );
  NAND2_X1 U5656 ( .A1(n6046), .A2(n6045), .ZN(n8476) );
  AND2_X1 U5657 ( .A1(n4706), .A2(n6178), .ZN(n8223) );
  AND2_X1 U5658 ( .A1(n8264), .A2(n8263), .ZN(n8489) );
  NAND2_X1 U5659 ( .A1(n4423), .A2(n4424), .ZN(n8262) );
  NAND2_X1 U5660 ( .A1(n6027), .A2(n6026), .ZN(n8493) );
  NAND2_X1 U5661 ( .A1(n4845), .A2(n6025), .ZN(n8273) );
  NAND2_X1 U5662 ( .A1(n8290), .A2(n6024), .ZN(n4845) );
  NAND2_X1 U5663 ( .A1(n4830), .A2(n4829), .ZN(n8316) );
  AND2_X1 U5664 ( .A1(n4830), .A2(n4333), .ZN(n8318) );
  NAND2_X1 U5665 ( .A1(n8332), .A2(n5991), .ZN(n4830) );
  NAND2_X1 U5666 ( .A1(n8365), .A2(n5963), .ZN(n8351) );
  NAND2_X1 U5667 ( .A1(n4854), .A2(n4857), .ZN(n8424) );
  NAND2_X1 U5668 ( .A1(n4683), .A2(n7925), .ZN(n7466) );
  NAND2_X1 U5669 ( .A1(n5919), .A2(n5918), .ZN(n7459) );
  NAND2_X1 U5670 ( .A1(n6169), .A2(n7916), .ZN(n7302) );
  AND2_X1 U5671 ( .A1(n7309), .A2(n5896), .ZN(n7346) );
  INV_X1 U5672 ( .A(n4838), .ZN(n6931) );
  AOI21_X1 U5673 ( .B1(n4842), .B2(n4839), .A(n4383), .ZN(n4838) );
  INV_X1 U5674 ( .A(n4840), .ZN(n4839) );
  NAND2_X1 U5675 ( .A1(n4842), .A2(n5840), .ZN(n7022) );
  NAND2_X1 U5676 ( .A1(n8438), .A2(n6467), .ZN(n8408) );
  NOR2_X1 U5677 ( .A1(n6193), .A2(n8152), .ZN(n7324) );
  OAI211_X1 U5678 ( .C1(n5864), .C2(n6246), .A(n5797), .B(n5796), .ZN(n7157)
         );
  NAND2_X1 U5679 ( .A1(n9994), .A2(n6154), .ZN(n8440) );
  INV_X1 U5680 ( .A(n6469), .ZN(n6154) );
  NAND2_X1 U5681 ( .A1(n5821), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5776) );
  AND2_X1 U5682 ( .A1(n7324), .A2(n8539), .ZN(n8420) );
  AND2_X2 U5683 ( .A1(n6445), .A2(n6465), .ZN(n10069) );
  AOI211_X1 U5684 ( .C1(n10045), .C2(n9749), .A(n9753), .B(n9748), .ZN(n9756)
         );
  AOI211_X1 U5685 ( .C1(n10045), .C2(n9754), .A(n9753), .B(n9752), .ZN(n9757)
         );
  OAI21_X1 U5686 ( .B1(n8458), .B2(n10028), .A(n4318), .ZN(n8563) );
  AND2_X1 U5687 ( .A1(n6557), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10000) );
  NOR2_X1 U5688 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5726) );
  NAND2_X1 U5689 ( .A1(n6141), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6117) );
  INV_X1 U5690 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7038) );
  INV_X1 U5691 ( .A(n8027), .ZN(n7036) );
  INV_X1 U5692 ( .A(n8019), .ZN(n7815) );
  INV_X1 U5693 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6868) );
  INV_X1 U5694 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6747) );
  INV_X1 U5695 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6346) );
  INV_X1 U5696 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6295) );
  INV_X1 U5697 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6269) );
  XNOR2_X1 U5698 ( .A(n4556), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6635) );
  NAND2_X1 U5699 ( .A1(n4557), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4556) );
  INV_X1 U5700 ( .A(n5795), .ZN(n4557) );
  AND4_X1 U5701 ( .A1(n5077), .A2(n5076), .A3(n5075), .A4(n5074), .ZN(n7233)
         );
  OAI211_X1 U5702 ( .C1(n8837), .C2(n6261), .A(n5112), .B(n5111), .ZN(n7246)
         );
  INV_X1 U5703 ( .A(n9257), .ZN(n9444) );
  OAI21_X1 U5704 ( .B1(n5415), .B2(n4520), .A(n4521), .ZN(n8609) );
  NAND2_X1 U5705 ( .A1(n8704), .A2(n8706), .ZN(n4810) );
  AND3_X1 U5706 ( .A1(n5461), .A2(n5460), .A3(n5459), .ZN(n9284) );
  NAND2_X1 U5707 ( .A1(n4450), .A2(n4790), .ZN(n8715) );
  INV_X1 U5708 ( .A(n4786), .ZN(n4785) );
  NAND2_X1 U5709 ( .A1(n4784), .A2(n4793), .ZN(n4791) );
  OAI21_X1 U5710 ( .B1(n8679), .B2(n8677), .A(n5561), .ZN(n4786) );
  NAND2_X1 U5711 ( .A1(n5573), .A2(n5572), .ZN(n9434) );
  AND2_X1 U5712 ( .A1(n4808), .A2(n8727), .ZN(n8660) );
  AND4_X1 U5713 ( .A1(n5359), .A2(n5358), .A3(n5357), .A4(n5356), .ZN(n9359)
         );
  NAND2_X1 U5714 ( .A1(n5037), .A2(n6584), .ZN(n6585) );
  NAND2_X1 U5715 ( .A1(n4814), .A2(n7092), .ZN(n7224) );
  NAND2_X1 U5716 ( .A1(n4519), .A2(n5445), .ZN(n4518) );
  NAND2_X1 U5717 ( .A1(n4799), .A2(n4796), .ZN(n8696) );
  AND4_X1 U5718 ( .A1(n5192), .A2(n5191), .A3(n5190), .A4(n5189), .ZN(n9799)
         );
  NAND2_X1 U5719 ( .A1(n4816), .A2(n4815), .ZN(n6457) );
  NAND2_X1 U5720 ( .A1(n6421), .A2(n4817), .ZN(n4815) );
  INV_X1 U5721 ( .A(n6422), .ZN(n4817) );
  AND2_X1 U5722 ( .A1(n4985), .A2(n4986), .ZN(n6458) );
  AND4_X1 U5723 ( .A1(n5104), .A2(n5103), .A3(n5102), .A4(n5101), .ZN(n7128)
         );
  INV_X1 U5724 ( .A(n8723), .ZN(n8736) );
  INV_X1 U5725 ( .A(n8717), .ZN(n8740) );
  NAND2_X1 U5726 ( .A1(n4886), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4887) );
  INV_X1 U5727 ( .A(n9192), .ZN(n9157) );
  INV_X1 U5728 ( .A(n9265), .ZN(n9116) );
  NAND2_X1 U5729 ( .A1(n5509), .A2(n5508), .ZN(n9114) );
  INV_X1 U5730 ( .A(n7129), .ZN(n9023) );
  INV_X1 U5731 ( .A(n6807), .ZN(n9025) );
  NAND3_X1 U5732 ( .A1(n4976), .A2(n4975), .A3(n4974), .ZN(n9026) );
  NAND2_X1 U5733 ( .A1(n4987), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4780) );
  NAND2_X1 U5734 ( .A1(n4953), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4781) );
  NAND2_X1 U5735 ( .A1(n6389), .A2(n6388), .ZN(n6387) );
  AND2_X1 U5736 ( .A1(n4966), .A2(n5019), .ZN(n5020) );
  NAND2_X1 U5737 ( .A1(n6333), .A2(n4487), .ZN(n9896) );
  OR2_X1 U5738 ( .A1(n6337), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4487) );
  NAND2_X1 U5739 ( .A1(n9896), .A2(n9897), .ZN(n9895) );
  INV_X1 U5740 ( .A(n4485), .ZN(n7198) );
  NAND2_X1 U5741 ( .A1(n4491), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4490) );
  NAND2_X1 U5742 ( .A1(n9045), .A2(n4491), .ZN(n4489) );
  INV_X1 U5743 ( .A(n9047), .ZN(n4491) );
  AND2_X1 U5744 ( .A1(n6231), .A2(n4312), .ZN(n9912) );
  NAND2_X1 U5745 ( .A1(n8838), .A2(n8837), .ZN(n9743) );
  MUX2_X1 U5746 ( .A(n8836), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8835), .Z(n8838) );
  INV_X1 U5747 ( .A(n9099), .ZN(n9814) );
  AND2_X1 U5748 ( .A1(n5679), .A2(n5597), .ZN(n9213) );
  NOR2_X1 U5749 ( .A1(n4327), .A2(n9206), .ZN(n9208) );
  NAND2_X1 U5750 ( .A1(n4370), .A2(n4872), .ZN(n9260) );
  AND2_X1 U5751 ( .A1(n5454), .A2(n5453), .ZN(n9299) );
  NAND2_X1 U5752 ( .A1(n9346), .A2(n4650), .ZN(n4643) );
  NAND2_X1 U5753 ( .A1(n4652), .A2(n4653), .ZN(n9336) );
  AND2_X1 U5754 ( .A1(n4630), .A2(n8923), .ZN(n9373) );
  NAND2_X1 U5755 ( .A1(n9792), .A2(n6967), .ZN(n9404) );
  NAND2_X1 U5756 ( .A1(n4656), .A2(n4657), .ZN(n9103) );
  NAND2_X1 U5757 ( .A1(n7550), .A2(n4660), .ZN(n4656) );
  NAND2_X1 U5758 ( .A1(n5267), .A2(n5266), .ZN(n9779) );
  NAND2_X1 U5759 ( .A1(n5236), .A2(n5235), .ZN(n7548) );
  NAND2_X1 U5760 ( .A1(n5205), .A2(n5204), .ZN(n9809) );
  NAND2_X1 U5761 ( .A1(n5160), .A2(n5159), .ZN(n7335) );
  OR3_X1 U5762 ( .A1(n5138), .A2(n5137), .A3(n5136), .ZN(n7294) );
  NAND2_X1 U5763 ( .A1(n6954), .A2(n6953), .ZN(n6956) );
  NOR2_X1 U5764 ( .A1(n9415), .A2(n4869), .ZN(n9416) );
  OR2_X1 U5765 ( .A1(n9414), .A2(n9413), .ZN(n4869) );
  INV_X1 U5766 ( .A(n9419), .ZN(n4636) );
  AOI21_X1 U5767 ( .B1(n9418), .B2(n9967), .A(n4415), .ZN(n4635) );
  OR2_X1 U5768 ( .A1(n9420), .A2(n4378), .ZN(n4415) );
  AND2_X2 U5769 ( .A1(n6416), .A2(n6411), .ZN(n9971) );
  INV_X1 U5770 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4932) );
  INV_X1 U5771 ( .A(n5641), .ZN(n7364) );
  INV_X1 U5772 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7210) );
  XNOR2_X1 U5773 ( .A(n5539), .B(n5538), .ZN(n7207) );
  NAND2_X1 U5774 ( .A1(n4475), .A2(n5515), .ZN(n5539) );
  INV_X1 U5775 ( .A(n5663), .ZN(n6948) );
  INV_X1 U5776 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6865) );
  NAND2_X1 U5777 ( .A1(n4535), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4888) );
  INV_X1 U5778 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6745) );
  AND2_X1 U5779 ( .A1(n5376), .A2(n5398), .ZN(n9083) );
  INV_X1 U5780 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6371) );
  INV_X1 U5781 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6275) );
  INV_X1 U5782 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6272) );
  XNOR2_X1 U5783 ( .A(n4431), .B(n5129), .ZN(n6262) );
  NAND2_X1 U5784 ( .A1(n4432), .A2(n5109), .ZN(n4431) );
  NAND2_X1 U5785 ( .A1(n5107), .A2(n5106), .ZN(n4432) );
  XNOR2_X1 U5786 ( .A(n4948), .B(n4947), .ZN(n6242) );
  NOR2_X1 U5787 ( .A1(n9538), .A2(n10099), .ZN(n10098) );
  AOI21_X1 U5788 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10096), .ZN(n10095) );
  NOR2_X1 U5789 ( .A1(n10095), .A2(n10094), .ZN(n10093) );
  AOI21_X1 U5790 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10093), .ZN(n10092) );
  AND2_X1 U5791 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9730) );
  INV_X1 U5792 ( .A(SI_8_), .ZN(n9727) );
  CLKBUF_X1 U5793 ( .A(n7694), .Z(P2_U3152) );
  NAND2_X1 U5794 ( .A1(n6857), .A2(n6856), .ZN(n6913) );
  AOI21_X1 U5795 ( .B1(n4589), .B2(n8023), .A(n4319), .ZN(n8030) );
  OAI21_X1 U5796 ( .B1(n9201), .B2(n8726), .A(n5693), .ZN(n5694) );
  OAI21_X1 U5797 ( .B1(n9090), .B2(n9161), .A(n4494), .ZN(P1_U3260) );
  AOI21_X1 U5798 ( .B1(n4496), .B2(n9161), .A(n4495), .ZN(n4494) );
  OAI21_X1 U5799 ( .B1(n9925), .B2(n9092), .A(n9091), .ZN(n4495) );
  XNOR2_X1 U5800 ( .A(n4887), .B(P1_IR_REG_22__SCAN_IN), .ZN(n5662) );
  INV_X1 U5801 ( .A(n5821), .ZN(n5877) );
  OR3_X1 U5802 ( .A1(n8211), .A2(n4610), .A3(n9754), .ZN(n4314) );
  INV_X1 U5803 ( .A(n6936), .ZN(n6478) );
  INV_X1 U5804 ( .A(n9376), .ZN(n9332) );
  AND4_X1 U5805 ( .A1(n5385), .A2(n5384), .A3(n5383), .A4(n5382), .ZN(n9376)
         );
  NAND2_X1 U5806 ( .A1(n4859), .A2(n5708), .ZN(n5806) );
  AND2_X1 U5807 ( .A1(n6178), .A2(n7978), .ZN(n7974) );
  INV_X1 U5808 ( .A(n4797), .ZN(n4439) );
  OR2_X1 U5809 ( .A1(n9486), .A2(n9770), .ZN(n4315) );
  OR2_X1 U5810 ( .A1(n5415), .A2(n5416), .ZN(n4316) );
  AND2_X1 U5811 ( .A1(n4587), .A2(n5906), .ZN(n4317) );
  INV_X1 U5812 ( .A(n4647), .ZN(n4646) );
  OAI21_X1 U5813 ( .B1(n9335), .B2(n4648), .A(n4348), .ZN(n4647) );
  INV_X1 U5814 ( .A(n7901), .ZN(n5878) );
  AND2_X1 U5815 ( .A1(n7905), .A2(n7904), .ZN(n7901) );
  AND2_X1 U5816 ( .A1(n8457), .A2(n8456), .ZN(n4318) );
  INV_X1 U5817 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5965) );
  NOR2_X1 U5818 ( .A1(n7835), .A2(n4390), .ZN(n4319) );
  AND2_X1 U5819 ( .A1(n8920), .A2(n4634), .ZN(n4320) );
  OAI21_X1 U5820 ( .B1(n8679), .B2(n4789), .A(n4788), .ZN(n4787) );
  INV_X1 U5821 ( .A(n4787), .ZN(n4450) );
  INV_X1 U5822 ( .A(n8289), .ZN(n4698) );
  AND2_X1 U5823 ( .A1(n5308), .A2(n7473), .ZN(n4321) );
  NAND2_X1 U5824 ( .A1(n7959), .A2(n8309), .ZN(n4322) );
  INV_X1 U5825 ( .A(n4863), .ZN(n4862) );
  NAND2_X1 U5826 ( .A1(n5895), .A2(n5879), .ZN(n4863) );
  AND4_X1 U5827 ( .A1(n6014), .A2(n6013), .A3(n6012), .A4(n6011), .ZN(n7729)
         );
  INV_X1 U5828 ( .A(n7729), .ZN(n4560) );
  NAND2_X1 U5829 ( .A1(n6068), .A2(n6067), .ZN(n8464) );
  NAND2_X1 U5830 ( .A1(n4400), .A2(n4882), .ZN(n5233) );
  AND2_X1 U5831 ( .A1(n6093), .A2(n6092), .ZN(n8196) );
  INV_X1 U5832 ( .A(n7165), .ZN(n6674) );
  INV_X1 U5833 ( .A(n5012), .ZN(n5623) );
  NAND2_X2 U5834 ( .A1(n4920), .A2(n4922), .ZN(n5012) );
  NAND2_X1 U5835 ( .A1(n5281), .A2(n5282), .ZN(n4323) );
  NAND2_X4 U5836 ( .A1(n5730), .A2(n5733), .ZN(n5800) );
  NAND2_X1 U5837 ( .A1(n6017), .A2(n6016), .ZN(n8499) );
  OR3_X1 U5838 ( .A1(n8306), .A2(n4608), .A3(n8499), .ZN(n4324) );
  OR2_X1 U5839 ( .A1(n4834), .A2(n4831), .ZN(n4325) );
  AND2_X1 U5840 ( .A1(n4950), .A2(n4499), .ZN(n4326) );
  AND2_X1 U5841 ( .A1(n8254), .A2(n7960), .ZN(n8279) );
  NOR2_X1 U5842 ( .A1(n9234), .A2(n9146), .ZN(n4327) );
  OR2_X1 U5843 ( .A1(n9486), .A2(n9105), .ZN(n9133) );
  OR2_X1 U5844 ( .A1(n9481), .A2(n9359), .ZN(n9136) );
  NAND2_X1 U5845 ( .A1(n8993), .A2(n9096), .ZN(n4328) );
  INV_X1 U5846 ( .A(n7925), .ZN(n4682) );
  AND2_X1 U5847 ( .A1(n6650), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4329) );
  INV_X1 U5848 ( .A(n9449), .ZN(n9272) );
  NAND2_X1 U5849 ( .A1(n5499), .A2(n5498), .ZN(n9449) );
  OR2_X1 U5850 ( .A1(n8479), .A2(n8258), .ZN(n6178) );
  AND2_X1 U5851 ( .A1(n6387), .A2(n4486), .ZN(n4330) );
  INV_X1 U5852 ( .A(n8208), .ZN(n4701) );
  AND2_X1 U5853 ( .A1(n4528), .A2(n5338), .ZN(n4331) );
  OR2_X1 U5854 ( .A1(n8027), .A2(n8019), .ZN(n6479) );
  NAND3_X1 U5855 ( .A1(n4864), .A2(n4865), .A3(n4605), .ZN(n5742) );
  NAND2_X1 U5856 ( .A1(n4588), .A2(n5906), .ZN(n7386) );
  AND3_X1 U5857 ( .A1(n4966), .A2(n5019), .A3(n4878), .ZN(n5053) );
  NAND2_X1 U5858 ( .A1(n5295), .A2(n5294), .ZN(n9486) );
  AND2_X1 U5859 ( .A1(n4537), .A2(n4536), .ZN(n4332) );
  OR2_X1 U5860 ( .A1(n8514), .A2(n8327), .ZN(n4333) );
  NOR2_X1 U5861 ( .A1(n7932), .A2(n5768), .ZN(n4334) );
  INV_X1 U5862 ( .A(n8653), .ZN(n4792) );
  INV_X1 U5863 ( .A(n9146), .ZN(n4625) );
  OR2_X1 U5864 ( .A1(n4906), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4335) );
  NOR3_X1 U5865 ( .A1(n9294), .A2(n4508), .A3(n9439), .ZN(n4506) );
  AND2_X1 U5866 ( .A1(n8835), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4336) );
  INV_X1 U5867 ( .A(n7473), .ZN(n4530) );
  AND2_X1 U5868 ( .A1(n4900), .A2(n4901), .ZN(n4337) );
  INV_X1 U5869 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8588) );
  NOR2_X1 U5870 ( .A1(n5010), .A2(n4921), .ZN(n4338) );
  AND2_X1 U5871 ( .A1(n5978), .A2(n5963), .ZN(n4339) );
  NAND2_X1 U5872 ( .A1(n7814), .A2(n7813), .ZN(n9754) );
  AND2_X1 U5873 ( .A1(n4699), .A2(n7966), .ZN(n4340) );
  NAND2_X1 U5874 ( .A1(n5982), .A2(n5981), .ZN(n8514) );
  INV_X1 U5875 ( .A(n4507), .ZN(n9251) );
  NOR2_X1 U5876 ( .A1(n9294), .A2(n4508), .ZN(n4507) );
  NAND2_X1 U5877 ( .A1(n5795), .A2(n5707), .ZN(n5807) );
  AND2_X1 U5878 ( .A1(n5176), .A2(n4455), .ZN(n4341) );
  INV_X1 U5879 ( .A(n8706), .ZN(n4523) );
  AND2_X1 U5880 ( .A1(n8510), .A2(n8344), .ZN(n4342) );
  AND2_X1 U5881 ( .A1(n4791), .A2(n4785), .ZN(n4343) );
  INV_X1 U5882 ( .A(n9005), .ZN(n7016) );
  AND2_X1 U5883 ( .A1(n6866), .A2(n9001), .ZN(n9005) );
  INV_X1 U5884 ( .A(n5489), .ZN(n4800) );
  OR2_X1 U5885 ( .A1(n4889), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n4535) );
  NOR2_X1 U5886 ( .A1(n8493), .A2(n8297), .ZN(n4344) );
  INV_X1 U5887 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5709) );
  AND2_X1 U5888 ( .A1(n7973), .A2(n7976), .ZN(n8261) );
  AND2_X1 U5889 ( .A1(n4527), .A2(n4525), .ZN(n4345) );
  INV_X1 U5890 ( .A(n4595), .ZN(n4594) );
  NAND2_X1 U5891 ( .A1(n4597), .A2(n4596), .ZN(n4595) );
  AND2_X1 U5892 ( .A1(n5130), .A2(SI_7_), .ZN(n4346) );
  NOR2_X1 U5893 ( .A1(n9462), .A2(n9333), .ZN(n4347) );
  NAND2_X1 U5894 ( .A1(n9468), .A2(n9322), .ZN(n4348) );
  INV_X1 U5895 ( .A(n4853), .ZN(n4852) );
  NAND2_X1 U5896 ( .A1(n8428), .A2(n4857), .ZN(n4853) );
  AND2_X1 U5897 ( .A1(n6794), .A2(n6793), .ZN(n4349) );
  OR2_X1 U5898 ( .A1(n6036), .A2(n6176), .ZN(n4350) );
  INV_X1 U5899 ( .A(n4623), .ZN(n4622) );
  NAND2_X1 U5900 ( .A1(n4626), .A2(n4624), .ZN(n4623) );
  AND2_X1 U5901 ( .A1(n7929), .A2(n7930), .ZN(n8423) );
  AND2_X1 U5902 ( .A1(n5264), .A2(n4337), .ZN(n4351) );
  AND2_X1 U5903 ( .A1(n4725), .A2(n4724), .ZN(n4352) );
  NOR2_X1 U5904 ( .A1(n9319), .A2(n9305), .ZN(n4353) );
  NAND2_X1 U5905 ( .A1(n7974), .A2(n7973), .ZN(n4354) );
  INV_X1 U5906 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4897) );
  AND2_X1 U5907 ( .A1(n5720), .A2(n4606), .ZN(n4355) );
  NAND2_X1 U5908 ( .A1(n7347), .A2(n5896), .ZN(n4356) );
  AND2_X1 U5909 ( .A1(n8753), .A2(n8759), .ZN(n8920) );
  AND3_X1 U5910 ( .A1(n4969), .A2(n4968), .A3(n4967), .ZN(n9403) );
  NAND2_X1 U5911 ( .A1(n9106), .A2(n4657), .ZN(n4357) );
  INV_X1 U5912 ( .A(n8303), .ZN(n4824) );
  INV_X1 U5913 ( .A(n9351), .ZN(n9476) );
  AND2_X1 U5914 ( .A1(n5378), .A2(n5377), .ZN(n9351) );
  AND2_X1 U5915 ( .A1(n4746), .A2(n4745), .ZN(n4358) );
  NAND2_X1 U5916 ( .A1(n5970), .A2(n5969), .ZN(n8521) );
  AND2_X1 U5917 ( .A1(n8423), .A2(n4677), .ZN(n4359) );
  NOR2_X1 U5918 ( .A1(n7611), .A2(n4730), .ZN(n4360) );
  AND2_X1 U5919 ( .A1(n6127), .A2(n6130), .ZN(n4361) );
  NOR2_X1 U5920 ( .A1(n5807), .A2(n4860), .ZN(n5833) );
  OAI21_X1 U5921 ( .B1(n9188), .B2(n9128), .A(n9129), .ZN(n9170) );
  NAND2_X1 U5922 ( .A1(n6102), .A2(n6101), .ZN(n8455) );
  OR2_X1 U5923 ( .A1(n4799), .A2(n4796), .ZN(n4362) );
  AND2_X1 U5924 ( .A1(n9136), .A2(n4631), .ZN(n4363) );
  NOR2_X1 U5925 ( .A1(n4469), .A2(n4464), .ZN(n4463) );
  OR2_X1 U5926 ( .A1(n9735), .A2(n9799), .ZN(n8897) );
  AND2_X1 U5927 ( .A1(n4447), .A2(n4446), .ZN(n4364) );
  AND2_X1 U5928 ( .A1(n7105), .A2(n7103), .ZN(n4365) );
  AND2_X1 U5929 ( .A1(n4910), .A2(n4820), .ZN(n4366) );
  AND2_X1 U5930 ( .A1(n4810), .A2(n4316), .ZN(n4367) );
  AND2_X1 U5931 ( .A1(n4442), .A2(n4439), .ZN(n4438) );
  INV_X1 U5932 ( .A(n4697), .ZN(n4696) );
  NAND2_X1 U5933 ( .A1(n4698), .A2(n7966), .ZN(n4697) );
  OR2_X1 U5934 ( .A1(n8653), .A2(n8677), .ZN(n4368) );
  INV_X1 U5935 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4592) );
  NOR2_X1 U5936 ( .A1(n8713), .A2(n8714), .ZN(n4369) );
  INV_X1 U5937 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4446) );
  INV_X1 U5938 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4534) );
  INV_X1 U5939 ( .A(n5798), .ZN(n6107) );
  INV_X1 U5940 ( .A(n5010), .ZN(n4953) );
  AND4_X1 U5941 ( .A1(n5903), .A2(n5902), .A3(n5901), .A4(n5900), .ZN(n7387)
         );
  INV_X1 U5942 ( .A(n7387), .ZN(n4587) );
  INV_X1 U5943 ( .A(n5514), .ZN(n4796) );
  AND2_X1 U5944 ( .A1(n5552), .A2(n5551), .ZN(n9250) );
  INV_X1 U5945 ( .A(n9250), .ZN(n9120) );
  NAND2_X1 U5946 ( .A1(n5966), .A2(n5965), .ZN(n5992) );
  INV_X1 U5947 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n4428) );
  AOI21_X1 U5948 ( .B1(n7550), .B2(n8879), .A(n7549), .ZN(n9758) );
  NAND2_X1 U5949 ( .A1(n4664), .A2(n7519), .ZN(n9782) );
  OR2_X1 U5950 ( .A1(n9275), .A2(n9280), .ZN(n4370) );
  XOR2_X1 U5951 ( .A(n5534), .B(n6950), .Z(n4371) );
  AND2_X1 U5952 ( .A1(n4643), .A2(n4646), .ZN(n4372) );
  NAND2_X1 U5953 ( .A1(n5473), .A2(n5472), .ZN(n9454) );
  NAND2_X1 U5954 ( .A1(n8844), .A2(n8843), .ZN(n9412) );
  INV_X1 U5955 ( .A(n9148), .ZN(n4626) );
  AND2_X1 U5956 ( .A1(n4758), .A2(n4478), .ZN(n4373) );
  OR2_X1 U5957 ( .A1(n4503), .A2(n9760), .ZN(n4374) );
  INV_X1 U5958 ( .A(n4607), .ZN(n8494) );
  NOR3_X1 U5959 ( .A1(n8306), .A2(n8499), .A3(n4609), .ZN(n4607) );
  NOR2_X1 U5960 ( .A1(n9044), .A2(n9045), .ZN(n4375) );
  INV_X1 U5961 ( .A(n8210), .ZN(n8180) );
  AND2_X1 U5962 ( .A1(n6074), .A2(n6073), .ZN(n8210) );
  AND2_X1 U5963 ( .A1(n9150), .A2(n8950), .ZN(n9171) );
  INV_X1 U5964 ( .A(n9422), .ZN(n9201) );
  NAND2_X1 U5965 ( .A1(n5622), .A2(n5621), .ZN(n9422) );
  AND2_X1 U5966 ( .A1(n5935), .A2(n5751), .ZN(n7419) );
  INV_X1 U5967 ( .A(n8677), .ZN(n4793) );
  NOR2_X1 U5968 ( .A1(n8402), .A2(n8533), .ZN(n4604) );
  NAND2_X1 U5969 ( .A1(n8365), .A2(n4339), .ZN(n8349) );
  INV_X1 U5970 ( .A(n8688), .ZN(n4445) );
  AND2_X1 U5971 ( .A1(n5264), .A2(n4364), .ZN(n5372) );
  AND2_X1 U5972 ( .A1(n5492), .A2(SI_21_), .ZN(n4376) );
  OR2_X1 U5973 ( .A1(n4776), .A2(n4774), .ZN(n4377) );
  NOR2_X1 U5974 ( .A1(n8697), .A2(n5514), .ZN(n4797) );
  INV_X1 U5975 ( .A(n4649), .ZN(n9473) );
  NAND2_X1 U5976 ( .A1(n4652), .A2(n4650), .ZN(n4649) );
  INV_X1 U5977 ( .A(n4400), .ZN(n5052) );
  AND2_X1 U5978 ( .A1(n9421), .A2(n9935), .ZN(n4378) );
  AND2_X1 U5979 ( .A1(n4758), .A2(n4479), .ZN(n4379) );
  AND2_X1 U5980 ( .A1(n4510), .A2(n9166), .ZN(n4380) );
  INV_X1 U5981 ( .A(n9243), .ZN(n9439) );
  AND2_X1 U5982 ( .A1(n5543), .A2(n5542), .ZN(n9243) );
  AND2_X1 U5983 ( .A1(n4770), .A2(n4480), .ZN(n4381) );
  INV_X1 U5984 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4847) );
  INV_X1 U5985 ( .A(n4552), .ZN(n4551) );
  NAND2_X1 U5986 ( .A1(n7270), .A2(n7838), .ZN(n4842) );
  NAND2_X1 U5987 ( .A1(n5350), .A2(n5349), .ZN(n9481) );
  INV_X1 U5988 ( .A(n9481), .ZN(n4502) );
  AND2_X1 U5989 ( .A1(n6585), .A2(n5041), .ZN(n4382) );
  INV_X1 U5990 ( .A(n8910), .ZN(n4619) );
  NAND2_X1 U5991 ( .A1(n6755), .A2(n6556), .ZN(n6789) );
  AND2_X1 U5992 ( .A1(n8045), .A2(n10024), .ZN(n4383) );
  NAND2_X1 U5993 ( .A1(n5956), .A2(n5955), .ZN(n8524) );
  INV_X1 U5994 ( .A(n8524), .ZN(n4603) );
  AND2_X1 U5995 ( .A1(n4864), .A2(n4865), .ZN(n4384) );
  NAND2_X1 U5996 ( .A1(n6006), .A2(n6005), .ZN(n8504) );
  INV_X1 U5997 ( .A(n8504), .ZN(n4561) );
  NAND2_X1 U5998 ( .A1(n7237), .A2(n7107), .ZN(n7109) );
  NAND2_X1 U5999 ( .A1(n7237), .A2(n4662), .ZN(n7296) );
  AND2_X1 U6000 ( .A1(n4718), .A2(n4717), .ZN(n4385) );
  AND2_X1 U6001 ( .A1(n6099), .A2(n6098), .ZN(n4386) );
  INV_X1 U6002 ( .A(n4753), .ZN(n4752) );
  OAI21_X1 U6003 ( .B1(n6076), .B2(n4754), .A(n6095), .ZN(n4753) );
  NAND2_X1 U6004 ( .A1(n7355), .A2(n4594), .ZN(n4598) );
  AND2_X1 U6005 ( .A1(n7104), .A2(n7103), .ZN(n4387) );
  NAND2_X1 U6006 ( .A1(n4402), .A2(n4821), .ZN(n4388) );
  XNOR2_X1 U6007 ( .A(n4933), .B(n4932), .ZN(n6211) );
  CLKBUF_X1 U6008 ( .A(n5777), .Z(n6673) );
  NAND2_X1 U6009 ( .A1(n6457), .A2(n6458), .ZN(n6456) );
  NAND2_X1 U6010 ( .A1(n6367), .A2(n6366), .ZN(n6365) );
  AND2_X1 U6011 ( .A1(n8128), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4389) );
  INV_X1 U6012 ( .A(n4498), .ZN(n6962) );
  NOR2_X1 U6013 ( .A1(n7053), .A2(n6816), .ZN(n4498) );
  AND2_X1 U6014 ( .A1(n10050), .A2(n7836), .ZN(n4390) );
  INV_X1 U6015 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n4555) );
  AND2_X1 U6016 ( .A1(n6517), .A2(n6516), .ZN(n4391) );
  OR2_X1 U6017 ( .A1(n7822), .A2(n4779), .ZN(n4392) );
  XNOR2_X1 U6018 ( .A(n4919), .B(P1_IR_REG_29__SCAN_IN), .ZN(n7688) );
  INV_X1 U6019 ( .A(n4848), .ZN(n5725) );
  NAND2_X1 U6020 ( .A1(n5737), .A2(n4846), .ZN(n4848) );
  INV_X1 U6021 ( .A(n9001), .ZN(n9161) );
  INV_X1 U6022 ( .A(n8012), .ZN(n8000) );
  MUX2_X1 U6023 ( .A(n7910), .B(n7909), .S(n8012), .Z(n7912) );
  OR2_X2 U6024 ( .A1(n8027), .A2(n7864), .ZN(n8012) );
  AOI21_X1 U6025 ( .B1(n4393), .B2(n8280), .A(n7968), .ZN(n7969) );
  NAND2_X1 U6026 ( .A1(n7967), .A2(n4394), .ZN(n4393) );
  NAND2_X1 U6027 ( .A1(n4396), .A2(n4395), .ZN(n7954) );
  NAND3_X1 U6028 ( .A1(n7943), .A2(n7941), .A3(n7942), .ZN(n4396) );
  NAND2_X2 U6029 ( .A1(n4868), .A2(n7557), .ZN(n9134) );
  NAND2_X2 U6030 ( .A1(n7655), .A2(n7654), .ZN(n7762) );
  NAND2_X2 U6031 ( .A1(n7597), .A2(n7596), .ZN(n7701) );
  AOI21_X2 U6032 ( .B1(n6755), .B2(n4740), .A(n4349), .ZN(n6795) );
  CLKBUF_X1 U6033 ( .A(n4403), .Z(n4400) );
  NAND2_X1 U6034 ( .A1(n4402), .A2(n4401), .ZN(n4913) );
  NAND3_X1 U6035 ( .A1(n4400), .A2(n4821), .A3(n4447), .ZN(n5347) );
  AND2_X1 U6036 ( .A1(n4403), .A2(n4821), .ZN(n5264) );
  NAND3_X1 U6037 ( .A1(n6517), .A2(n4407), .A3(n7040), .ZN(n4405) );
  NAND2_X1 U6038 ( .A1(n7040), .A2(n4406), .ZN(n4404) );
  NAND3_X1 U6039 ( .A1(n4410), .A2(n4654), .A3(n4409), .ZN(n9380) );
  NAND2_X1 U6040 ( .A1(n4365), .A2(n7104), .ZN(n7125) );
  AOI21_X1 U6041 ( .B1(n8221), .B2(n4419), .A(n4417), .ZN(n4416) );
  INV_X1 U6042 ( .A(n4416), .ZN(n8171) );
  INV_X4 U6043 ( .A(n8835), .ZN(n7824) );
  NAND2_X1 U6044 ( .A1(n5080), .A2(n5079), .ZN(n5083) );
  OAI21_X1 U6045 ( .B1(n8835), .B2(n4428), .A(n4427), .ZN(n5081) );
  NAND2_X1 U6046 ( .A1(n8835), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n4427) );
  NAND2_X1 U6047 ( .A1(n5059), .A2(n5058), .ZN(n4429) );
  INV_X1 U6048 ( .A(n7254), .ZN(n4433) );
  OAI21_X1 U6049 ( .B1(n4433), .B2(n4863), .A(n4434), .ZN(n7345) );
  NAND2_X1 U6050 ( .A1(n8686), .A2(n4438), .ZN(n4435) );
  NAND2_X2 U6051 ( .A1(n7447), .A2(n5256), .ZN(n7475) );
  INV_X2 U6052 ( .A(n5634), .ZN(n5605) );
  NAND2_X1 U6053 ( .A1(n6810), .A2(n5634), .ZN(n4980) );
  AND2_X4 U6054 ( .A1(n4934), .A2(n4940), .ZN(n5634) );
  AND2_X2 U6055 ( .A1(n6866), .A2(n5663), .ZN(n4940) );
  NAND3_X1 U6056 ( .A1(n4450), .A2(n4790), .A3(n4369), .ZN(n8718) );
  INV_X1 U6057 ( .A(n4566), .ZN(n4453) );
  NAND3_X1 U6058 ( .A1(n4568), .A2(n5176), .A3(n4457), .ZN(n4456) );
  NAND2_X1 U6059 ( .A1(n4566), .A2(n4568), .ZN(n5147) );
  NAND2_X1 U6060 ( .A1(n5226), .A2(n4463), .ZN(n4459) );
  NAND2_X1 U6061 ( .A1(n4755), .A2(n4379), .ZN(n4475) );
  AND2_X1 U6062 ( .A1(n4474), .A2(n4472), .ZN(n4775) );
  NAND2_X1 U6063 ( .A1(n4474), .A2(n4473), .ZN(n5567) );
  NAND2_X1 U6064 ( .A1(n4755), .A2(n4758), .ZN(n5517) );
  NAND2_X1 U6065 ( .A1(n4481), .A2(n4381), .ZN(n5449) );
  NAND2_X1 U6066 ( .A1(n5371), .A2(n5370), .ZN(n5397) );
  OAI21_X1 U6067 ( .B1(n7436), .B2(n4490), .A(n4489), .ZN(n9067) );
  NAND2_X2 U6068 ( .A1(n4949), .A2(n8835), .ZN(n5057) );
  INV_X1 U6069 ( .A(n9760), .ZN(n4500) );
  NAND2_X1 U6070 ( .A1(n4501), .A2(n4500), .ZN(n9365) );
  INV_X1 U6071 ( .A(n4506), .ZN(n9239) );
  NAND2_X1 U6072 ( .A1(n9211), .A2(n4380), .ZN(n4511) );
  NAND2_X1 U6073 ( .A1(n9211), .A2(n9201), .ZN(n9195) );
  INV_X1 U6074 ( .A(n4511), .ZN(n9160) );
  AOI21_X1 U6075 ( .B1(n9179), .B2(n9412), .A(n9963), .ZN(n4512) );
  AND2_X4 U6076 ( .A1(n4514), .A2(n4513), .ZN(n5606) );
  OR2_X4 U6077 ( .A1(n4940), .A2(n6199), .ZN(n4952) );
  INV_X1 U6078 ( .A(n5662), .ZN(n4515) );
  INV_X1 U6079 ( .A(n4517), .ZN(n8686) );
  NAND2_X1 U6080 ( .A1(n5280), .A2(n4331), .ZN(n4527) );
  NAND2_X1 U6081 ( .A1(n5280), .A2(n4323), .ZN(n4818) );
  NAND2_X1 U6082 ( .A1(n7005), .A2(n7006), .ZN(n7416) );
  NAND3_X1 U6083 ( .A1(n4549), .A2(n4548), .A3(n4546), .ZN(n7418) );
  NAND2_X1 U6084 ( .A1(n7005), .A2(n4550), .ZN(n4548) );
  OR2_X1 U6085 ( .A1(n7005), .A2(n4552), .ZN(n4549) );
  NAND2_X1 U6086 ( .A1(n7416), .A2(n4554), .ZN(n8089) );
  NOR2_X1 U6087 ( .A1(n7417), .A2(n7418), .ZN(n8091) );
  NAND2_X1 U6088 ( .A1(n4554), .A2(n8100), .ZN(n4552) );
  MUX2_X1 U6089 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n8835), .Z(n5025) );
  MUX2_X1 U6090 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8835), .Z(n5060) );
  NAND2_X1 U6091 ( .A1(n4563), .A2(n4558), .ZN(n7967) );
  OAI21_X1 U6092 ( .B1(n4562), .B2(n4559), .A(n8000), .ZN(n4558) );
  NAND2_X1 U6093 ( .A1(n7966), .A2(n7958), .ZN(n4559) );
  OAI21_X1 U6094 ( .B1(n4564), .B2(n4322), .A(n8012), .ZN(n4563) );
  AOI21_X1 U6095 ( .B1(n7957), .B2(n7955), .A(n4565), .ZN(n4564) );
  INV_X1 U6096 ( .A(n7958), .ZN(n4565) );
  NAND2_X1 U6097 ( .A1(n4567), .A2(n5107), .ZN(n4566) );
  NAND3_X1 U6098 ( .A1(n4583), .A2(n4579), .A3(n8423), .ZN(n7933) );
  NAND2_X1 U6099 ( .A1(n4581), .A2(n4580), .ZN(n4579) );
  NAND2_X1 U6100 ( .A1(n7927), .A2(n4582), .ZN(n4581) );
  AND2_X1 U6101 ( .A1(n7928), .A2(n8012), .ZN(n4584) );
  NAND2_X1 U6102 ( .A1(n7927), .A2(n4586), .ZN(n4585) );
  NAND2_X1 U6103 ( .A1(n6278), .A2(n7828), .ZN(n4588) );
  INV_X1 U6104 ( .A(n4598), .ZN(n8443) );
  INV_X1 U6105 ( .A(n8402), .ZN(n4599) );
  NAND2_X1 U6106 ( .A1(n4600), .A2(n4599), .ZN(n8319) );
  INV_X1 U6107 ( .A(n4604), .ZN(n8386) );
  NAND3_X1 U6108 ( .A1(n4864), .A2(n4865), .A3(n5720), .ZN(n6118) );
  NAND2_X1 U6109 ( .A1(n4924), .A2(n4923), .ZN(n4612) );
  NAND3_X1 U6110 ( .A1(n7044), .A2(n8914), .A3(n4618), .ZN(n4616) );
  NAND2_X1 U6111 ( .A1(n7044), .A2(n4618), .ZN(n4617) );
  NAND3_X1 U6112 ( .A1(n4616), .A2(n4614), .A3(n8913), .ZN(n7126) );
  NAND2_X1 U6113 ( .A1(n9134), .A2(n4363), .ZN(n4629) );
  NAND2_X1 U6114 ( .A1(n9134), .A2(n9133), .ZN(n9382) );
  INV_X1 U6115 ( .A(n4630), .ZN(n9384) );
  NAND2_X1 U6116 ( .A1(n4636), .A2(n4635), .ZN(n9490) );
  AOI21_X1 U6117 ( .B1(n9176), .B2(n9175), .A(n9802), .ZN(n4639) );
  OR2_X1 U6118 ( .A1(n5042), .A2(n4917), .ZN(n4925) );
  NAND2_X1 U6119 ( .A1(n6521), .A2(n6520), .ZN(n6809) );
  NAND2_X1 U6120 ( .A1(n7554), .A2(n8776), .ZN(n9767) );
  INV_X1 U6121 ( .A(n7040), .ZN(n8868) );
  NOR2_X1 U6122 ( .A1(n9189), .A2(n9149), .ZN(n9176) );
  NOR2_X1 U6123 ( .A1(n9357), .A2(n9138), .ZN(n9330) );
  NOR2_X2 U6124 ( .A1(n9028), .A2(n6509), .ZN(n6505) );
  AOI21_X1 U6125 ( .B1(n9321), .B2(n9320), .A(n9141), .ZN(n9301) );
  NOR2_X2 U6126 ( .A1(n7290), .A2(n7335), .ZN(n7338) );
  OAI21_X1 U6127 ( .B1(n8872), .B2(n4391), .A(n4641), .ZN(n9407) );
  NAND2_X1 U6128 ( .A1(n7518), .A2(n8878), .ZN(n4664) );
  OAI21_X1 U6129 ( .B1(n9275), .B2(n4667), .A(n4665), .ZN(n9246) );
  NAND2_X1 U6130 ( .A1(n9280), .A2(n4872), .ZN(n4668) );
  NAND3_X1 U6131 ( .A1(n6954), .A2(n6953), .A3(n6955), .ZN(n7104) );
  INV_X2 U6132 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U6133 ( .A1(n6169), .A2(n4359), .ZN(n4676) );
  NAND3_X1 U6134 ( .A1(n8423), .A2(n4677), .A3(n4680), .ZN(n4675) );
  NAND2_X1 U6135 ( .A1(n8416), .A2(n4687), .ZN(n4686) );
  NAND2_X1 U6136 ( .A1(n4686), .A2(n4689), .ZN(n8353) );
  OAI21_X1 U6137 ( .B1(n8324), .B2(n4697), .A(n4694), .ZN(n8252) );
  INV_X1 U6138 ( .A(n4706), .ZN(n8242) );
  NAND2_X1 U6139 ( .A1(n4709), .A2(n4712), .ZN(n4710) );
  INV_X1 U6140 ( .A(n6166), .ZN(n4709) );
  OAI211_X1 U6141 ( .C1(n6932), .C2(n4711), .A(n7905), .B(n4710), .ZN(n6167)
         );
  INV_X1 U6142 ( .A(n4712), .ZN(n4711) );
  NAND2_X1 U6143 ( .A1(n4713), .A2(n4712), .ZN(n7251) );
  NAND2_X1 U6144 ( .A1(n6932), .A2(n6166), .ZN(n4713) );
  NAND2_X1 U6145 ( .A1(n7395), .A2(n4717), .ZN(n4716) );
  OAI21_X2 U6146 ( .B1(n6795), .B2(n4721), .A(n4719), .ZN(n6973) );
  NAND2_X1 U6147 ( .A1(n6973), .A2(n6972), .ZN(n6978) );
  INV_X1 U6148 ( .A(n6911), .ZN(n4725) );
  NAND2_X1 U6149 ( .A1(n7701), .A2(n4360), .ZN(n4726) );
  OAI21_X2 U6150 ( .B1(n7737), .B2(n4736), .A(n4733), .ZN(n7790) );
  NAND2_X2 U6151 ( .A1(n6555), .A2(n6554), .ZN(n6755) );
  NAND3_X1 U6152 ( .A1(n7815), .A2(n6479), .A3(n8017), .ZN(n4742) );
  NAND2_X1 U6153 ( .A1(n5966), .A2(n4744), .ZN(n6112) );
  INV_X1 U6154 ( .A(n5950), .ZN(n4745) );
  NAND2_X1 U6155 ( .A1(n5951), .A2(n5952), .ZN(n5964) );
  NAND2_X1 U6156 ( .A1(n7718), .A2(n7628), .ZN(n7768) );
  INV_X1 U6157 ( .A(n6077), .ZN(n4750) );
  NAND2_X1 U6158 ( .A1(n5449), .A2(n4756), .ZN(n4755) );
  NAND2_X1 U6159 ( .A1(n4764), .A2(n9006), .ZN(n4768) );
  NAND3_X1 U6160 ( .A1(n4766), .A2(n4769), .A3(n4765), .ZN(n4764) );
  OAI211_X1 U6161 ( .C1(n8892), .C2(n8894), .A(n4767), .B(n9161), .ZN(n4765)
         );
  INV_X1 U6162 ( .A(n8893), .ZN(n4766) );
  NAND2_X1 U6163 ( .A1(n4768), .A2(n9011), .ZN(P1_U3240) );
  NAND2_X1 U6164 ( .A1(n4874), .A2(n9001), .ZN(n4769) );
  OAI21_X1 U6165 ( .B1(n5397), .B2(n5396), .A(n5395), .ZN(n5420) );
  NAND2_X1 U6166 ( .A1(n5396), .A2(n5395), .ZN(n4773) );
  NAND2_X1 U6167 ( .A1(n4775), .A2(n5540), .ZN(n5563) );
  NAND2_X1 U6168 ( .A1(n7584), .A2(n7585), .ZN(n7823) );
  NAND2_X1 U6169 ( .A1(n4777), .A2(n4778), .ZN(n7827) );
  NAND3_X1 U6170 ( .A1(n7584), .A2(n7585), .A3(n4392), .ZN(n4777) );
  NAND3_X2 U6171 ( .A1(n4782), .A2(n4781), .A3(n4780), .ZN(n6500) );
  INV_X1 U6172 ( .A(n4783), .ZN(n4782) );
  INV_X1 U6173 ( .A(n8678), .ZN(n4784) );
  AOI21_X1 U6174 ( .B1(n8679), .B2(n8678), .A(n8677), .ZN(n8681) );
  INV_X1 U6175 ( .A(n5312), .ZN(n4805) );
  NAND2_X1 U6176 ( .A1(n4802), .A2(n5338), .ZN(n8727) );
  NAND2_X1 U6177 ( .A1(n5312), .A2(n7569), .ZN(n4802) );
  NAND2_X1 U6178 ( .A1(n4805), .A2(n4804), .ZN(n4803) );
  INV_X1 U6179 ( .A(n5338), .ZN(n4806) );
  NAND2_X1 U6180 ( .A1(n8728), .A2(n8730), .ZN(n4808) );
  NAND2_X1 U6181 ( .A1(n4809), .A2(n5312), .ZN(n8728) );
  NAND3_X1 U6182 ( .A1(n4812), .A2(n5095), .A3(n4811), .ZN(n6873) );
  NAND3_X1 U6183 ( .A1(n6584), .A2(n5037), .A3(n5069), .ZN(n4812) );
  NAND2_X1 U6184 ( .A1(n4818), .A2(n4321), .ZN(n7568) );
  NAND2_X1 U6185 ( .A1(n4351), .A2(n4902), .ZN(n4906) );
  OAI21_X1 U6186 ( .B1(n8332), .B2(n4828), .A(n4826), .ZN(n8304) );
  AOI21_X1 U6187 ( .B1(n4826), .B2(n4828), .A(n4824), .ZN(n4823) );
  NAND3_X1 U6188 ( .A1(n4836), .A2(n5865), .A3(n4835), .ZN(n7254) );
  NAND3_X1 U6189 ( .A1(n7270), .A2(n4837), .A3(n7838), .ZN(n4836) );
  INV_X1 U6190 ( .A(n5840), .ZN(n4841) );
  OR2_X1 U6191 ( .A1(n8855), .A2(n8858), .ZN(n8856) );
  OAI21_X2 U6192 ( .B1(n7126), .B2(n7112), .A(n8915), .ZN(n8964) );
  NOR3_X1 U6193 ( .A1(n6196), .A2(n6195), .A3(n6194), .ZN(n6197) );
  OR2_X1 U6194 ( .A1(n8629), .A2(n4313), .ZN(n5689) );
  INV_X1 U6195 ( .A(n4931), .ZN(n4912) );
  NAND2_X1 U6196 ( .A1(n4933), .A2(n4911), .ZN(n4931) );
  INV_X1 U6197 ( .A(n9346), .ZN(n9348) );
  NAND2_X1 U6198 ( .A1(n6436), .A2(n5790), .ZN(n7159) );
  OR2_X1 U6199 ( .A1(n8458), .A2(n8422), .ZN(n6198) );
  OR2_X1 U6200 ( .A1(n4934), .A2(n6309), .ZN(n4866) );
  OR2_X1 U6201 ( .A1(n9809), .A2(n9017), .ZN(n4867) );
  INV_X1 U6202 ( .A(n8352), .ZN(n5978) );
  INV_X1 U6203 ( .A(n9486), .ZN(n9104) );
  AND2_X1 U6204 ( .A1(n5583), .A2(n5582), .ZN(n9238) );
  INV_X1 U6205 ( .A(n7996), .ZN(n6110) );
  NAND2_X1 U6206 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n4870) );
  AND2_X1 U6207 ( .A1(n6490), .A2(n6616), .ZN(n8341) );
  OR2_X1 U6208 ( .A1(n9285), .A2(n9272), .ZN(n4871) );
  OR2_X1 U6209 ( .A1(n9290), .A2(n9306), .ZN(n4872) );
  AND2_X1 U6210 ( .A1(n8961), .A2(n8960), .ZN(n4874) );
  AND2_X1 U6211 ( .A1(n5779), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n4875) );
  INV_X1 U6212 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9507) );
  NOR2_X1 U6213 ( .A1(n5813), .A2(n6160), .ZN(n4876) );
  AOI21_X1 U6214 ( .B1(n8214), .B2(n5815), .A(n6065), .ZN(n8226) );
  NAND2_X1 U6215 ( .A1(n8017), .A2(n7836), .ZN(n8434) );
  INV_X1 U6216 ( .A(n8870), .ZN(n6955) );
  INV_X1 U6217 ( .A(n7849), .ZN(n5895) );
  AND2_X2 U6218 ( .A1(n7242), .A2(n9789), .ZN(n9806) );
  INV_X1 U6219 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4896) );
  INV_X1 U6220 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5707) );
  AOI21_X1 U6221 ( .B1(n8179), .B2(n7861), .A(n6179), .ZN(n6180) );
  INV_X1 U6222 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5722) );
  INV_X1 U6223 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4910) );
  INV_X1 U6224 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4901) );
  OR2_X1 U6225 ( .A1(n5997), .A2(n5996), .ZN(n6007) );
  NAND2_X1 U6226 ( .A1(n5700), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5941) );
  INV_X1 U6227 ( .A(n7839), .ZN(n6159) );
  NAND2_X1 U6228 ( .A1(n7184), .A2(n7865), .ZN(n7871) );
  NAND2_X1 U6229 ( .A1(n6124), .A2(n6114), .ZN(n6115) );
  INV_X1 U6230 ( .A(n5526), .ZN(n5524) );
  INV_X1 U6231 ( .A(n5502), .ZN(n5500) );
  INV_X1 U6232 ( .A(n5404), .ZN(n5402) );
  INV_X1 U6233 ( .A(n5209), .ZN(n5207) );
  AND2_X1 U6234 ( .A1(n9412), .A2(n9935), .ZN(n9413) );
  INV_X1 U6235 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4902) );
  INV_X1 U6236 ( .A(SI_22_), .ZN(n9580) );
  INV_X1 U6237 ( .A(n5418), .ZN(n5419) );
  INV_X1 U6238 ( .A(SI_10_), .ZN(n9651) );
  INV_X1 U6239 ( .A(n7702), .ZN(n7603) );
  INV_X1 U6240 ( .A(n7398), .ZN(n7396) );
  OR2_X1 U6241 ( .A1(n6030), .A2(n7712), .ZN(n6040) );
  AND2_X1 U6242 ( .A1(n5841), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U6243 ( .A1(n5781), .A2(n5780), .ZN(n5782) );
  INV_X1 U6244 ( .A(n6643), .ZN(n6683) );
  OR2_X1 U6245 ( .A1(n8476), .A2(n8034), .ZN(n6056) );
  NAND2_X1 U6246 ( .A1(n6115), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U6247 ( .A1(n5524), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5545) );
  INV_X1 U6248 ( .A(n5143), .ZN(n5146) );
  INV_X1 U6249 ( .A(n5416), .ZN(n5417) );
  NAND2_X1 U6250 ( .A1(n5500), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U6251 ( .A1(n5430), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5455) );
  INV_X1 U6252 ( .A(n9152), .ZN(n9153) );
  NAND2_X1 U6253 ( .A1(n5402), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U6254 ( .A1(n5351), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6255 ( .A1(n5237), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5269) );
  NOR2_X1 U6256 ( .A1(n9351), .A2(n9376), .ZN(n9112) );
  INV_X1 U6257 ( .A(n6866), .ZN(n9002) );
  INV_X1 U6258 ( .A(SI_17_), .ZN(n9618) );
  NAND2_X1 U6259 ( .A1(n5261), .A2(n9634), .ZN(n5287) );
  NAND2_X1 U6260 ( .A1(n7657), .A2(n7656), .ZN(n7658) );
  AND3_X1 U6261 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5841) );
  OR2_X1 U6262 ( .A1(n5881), .A2(n5880), .ZN(n5897) );
  INV_X1 U6263 ( .A(n7794), .ZN(n7805) );
  INV_X1 U6264 ( .A(n5800), .ZN(n6104) );
  INV_X1 U6265 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9604) );
  INV_X1 U6266 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9661) );
  NAND2_X1 U6267 ( .A1(n7980), .A2(n7981), .ZN(n8224) );
  OR2_X1 U6268 ( .A1(n6603), .A2(n5774), .ZN(n5775) );
  INV_X1 U6269 ( .A(n8434), .ZN(n8410) );
  OR2_X1 U6270 ( .A1(n5545), .A2(n5544), .ZN(n5576) );
  OR2_X1 U6271 ( .A1(n5596), .A2(n8719), .ZN(n5679) );
  OR2_X1 U6272 ( .A1(n9226), .A2(n4313), .ZN(n5583) );
  INV_X1 U6273 ( .A(n5013), .ZN(n5478) );
  INV_X1 U6274 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6393) );
  AND2_X1 U6275 ( .A1(n9444), .A2(n9116), .ZN(n9117) );
  INV_X1 U6276 ( .A(n9333), .ZN(n9305) );
  XNOR2_X1 U6277 ( .A(n7827), .B(n7826), .ZN(n8836) );
  AND2_X1 U6278 ( .A1(n6078), .A2(n5620), .ZN(n6076) );
  AND2_X1 U6279 ( .A1(n5540), .A2(n5521), .ZN(n5538) );
  AND2_X1 U6280 ( .A1(n5370), .A2(n5346), .ZN(n5368) );
  AND2_X1 U6281 ( .A1(n5199), .A2(n5182), .ZN(n5197) );
  NOR2_X1 U6282 ( .A1(n10117), .A2(n10116), .ZN(n9525) );
  NAND2_X1 U6283 ( .A1(n6543), .A2(n6542), .ZN(n6672) );
  NOR2_X1 U6284 ( .A1(n7409), .A2(n8430), .ZN(n7793) );
  AND4_X1 U6285 ( .A1(n6035), .A2(n6034), .A3(n6033), .A4(n6032), .ZN(n8257)
         );
  AND4_X1 U6286 ( .A1(n5948), .A2(n5947), .A3(n5946), .A4(n5945), .ZN(n8413)
         );
  INV_X1 U6287 ( .A(n9981), .ZN(n9983) );
  AND2_X1 U6288 ( .A1(n6610), .A2(n6609), .ZN(n9981) );
  INV_X1 U6289 ( .A(n7974), .ZN(n8243) );
  INV_X1 U6290 ( .A(n7932), .ZN(n8411) );
  NAND2_X1 U6291 ( .A1(n7345), .A2(n5907), .ZN(n7300) );
  AND2_X1 U6292 ( .A1(n7897), .A2(n7894), .ZN(n7843) );
  INV_X1 U6293 ( .A(n8408), .ZN(n8450) );
  NOR2_X1 U6294 ( .A1(n9996), .A2(n6137), .ZN(n6465) );
  AND2_X1 U6295 ( .A1(n8427), .A2(n10031), .ZN(n10028) );
  AND2_X1 U6296 ( .A1(n7256), .A2(n7255), .ZN(n10036) );
  INV_X1 U6297 ( .A(n10028), .ZN(n10052) );
  NOR2_X1 U6298 ( .A1(n6432), .A2(n6431), .ZN(n6445) );
  AND2_X1 U6299 ( .A1(n6120), .A2(n4311), .ZN(n7511) );
  AND2_X1 U6300 ( .A1(n6202), .A2(n6232), .ZN(n6216) );
  INV_X1 U6301 ( .A(n8732), .ZN(n8708) );
  INV_X1 U6302 ( .A(n8720), .ZN(n8734) );
  OR2_X1 U6303 ( .A1(n5057), .A2(n6247), .ZN(n4968) );
  NAND2_X1 U6304 ( .A1(n5673), .A2(n6364), .ZN(n8723) );
  INV_X1 U6305 ( .A(n8726), .ZN(n8738) );
  AND4_X1 U6306 ( .A1(n5409), .A2(n5408), .A3(n5407), .A4(n5406), .ZN(n9360)
         );
  INV_X1 U6307 ( .A(n9921), .ZN(n9885) );
  AND2_X1 U6308 ( .A1(n6216), .A2(n6215), .ZN(n9920) );
  INV_X1 U6309 ( .A(n9128), .ZN(n9191) );
  INV_X1 U6310 ( .A(n9802), .ZN(n9768) );
  OR2_X1 U6311 ( .A1(n9824), .A2(n6949), .ZN(n9789) );
  INV_X1 U6312 ( .A(n9404), .ZN(n9810) );
  AND2_X1 U6313 ( .A1(n5647), .A2(n9506), .ZN(n6945) );
  INV_X1 U6314 ( .A(n9963), .ZN(n9816) );
  INV_X1 U6315 ( .A(n9967), .ZN(n9932) );
  INV_X1 U6316 ( .A(n7117), .ZN(n9805) );
  INV_X1 U6317 ( .A(n6945), .ZN(n6411) );
  AND2_X1 U6318 ( .A1(n5293), .A2(n5321), .ZN(n7439) );
  AND2_X1 U6319 ( .A1(n5158), .A2(n5202), .ZN(n6400) );
  INV_X1 U6320 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9520) );
  NOR2_X1 U6321 ( .A1(n9526), .A2(n9525), .ZN(n10112) );
  INV_X1 U6322 ( .A(n8157), .ZN(n9987) );
  INV_X1 U6323 ( .A(n7217), .ZN(n6496) );
  OR2_X1 U6324 ( .A1(n6492), .A2(n6491), .ZN(n7810) );
  INV_X1 U6325 ( .A(n8196), .ZN(n8032) );
  AND3_X1 U6326 ( .A1(n5736), .A2(n5735), .A3(n5734), .ZN(n8284) );
  INV_X1 U6327 ( .A(n8432), .ZN(n8040) );
  INV_X1 U6328 ( .A(n8150), .ZN(n9982) );
  INV_X1 U6329 ( .A(n9986), .ZN(n8138) );
  NAND2_X1 U6330 ( .A1(n6298), .A2(n6297), .ZN(n8157) );
  NAND2_X1 U6331 ( .A1(n8438), .A2(n6156), .ZN(n8422) );
  INV_X1 U6332 ( .A(n10069), .ZN(n10067) );
  INV_X1 U6333 ( .A(n10055), .ZN(n10054) );
  AND2_X2 U6334 ( .A1(n6445), .A2(n6433), .ZN(n10055) );
  NAND2_X1 U6335 ( .A1(n9994), .A2(n9993), .ZN(n9997) );
  XNOR2_X1 U6336 ( .A(n6117), .B(n6116), .ZN(n7368) );
  INV_X1 U6337 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6373) );
  INV_X1 U6338 ( .A(P2_STATE_REG_SCAN_IN), .ZN(n7694) );
  INV_X1 U6339 ( .A(n8594), .ZN(n7365) );
  INV_X1 U6340 ( .A(n9462), .ZN(n9319) );
  INV_X1 U6341 ( .A(n9224), .ZN(n9125) );
  INV_X1 U6342 ( .A(n9360), .ZN(n9322) );
  INV_X1 U6343 ( .A(n7287), .ZN(n9020) );
  INV_X1 U6344 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9866) );
  OR2_X1 U6345 ( .A1(P1_U3083), .A2(n6233), .ZN(n9925) );
  NAND2_X1 U6346 ( .A1(n9792), .A2(n6952), .ZN(n9398) );
  INV_X1 U6347 ( .A(n9980), .ZN(n9978) );
  AND2_X2 U6348 ( .A1(n6416), .A2(n6945), .ZN(n9980) );
  AND2_X1 U6349 ( .A1(n9830), .A2(n9829), .ZN(n9847) );
  AND2_X1 U6350 ( .A1(n9841), .A2(n9840), .ZN(n9851) );
  INV_X1 U6351 ( .A(n9971), .ZN(n9969) );
  AND2_X1 U6352 ( .A1(n4934), .A2(n5660), .ZN(n9505) );
  INV_X1 U6353 ( .A(n4920), .ZN(n7587) );
  INV_X1 U6354 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7431) );
  INV_X1 U6355 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7035) );
  INV_X1 U6356 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6455) );
  INV_X1 U6357 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6280) );
  NOR2_X1 U6358 ( .A1(n10101), .A2(n10100), .ZN(n10099) );
  NOR2_X1 U6359 ( .A1(n10098), .A2(n10097), .ZN(n10096) );
  INV_X1 U6360 ( .A(n8049), .ZN(P2_U3966) );
  NAND2_X1 U6361 ( .A1(n6198), .A2(n6197), .ZN(P2_U3267) );
  INV_X1 U6362 ( .A(n9027), .ZN(P1_U4006) );
  NOR2_X1 U6363 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4884) );
  NAND2_X1 U6364 ( .A1(n5372), .A2(n4884), .ZN(n4889) );
  INV_X1 U6365 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4885) );
  NAND2_X1 U6366 ( .A1(n4892), .A2(n4885), .ZN(n4886) );
  NAND2_X1 U6367 ( .A1(n4889), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4890) );
  MUX2_X1 U6368 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4890), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n4891) );
  NAND2_X1 U6369 ( .A1(n4891), .A2(n4535), .ZN(n9001) );
  NOR2_X1 U6370 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4895) );
  NAND4_X1 U6371 ( .A1(n4895), .A2(n4894), .A3(n4893), .A4(n5291), .ZN(n4899)
         );
  NAND4_X1 U6372 ( .A1(n4897), .A2(n4534), .A3(n4446), .A4(n4896), .ZN(n4898)
         );
  NAND2_X1 U6373 ( .A1(n4335), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4903) );
  INV_X1 U6374 ( .A(n4351), .ZN(n4904) );
  NAND2_X1 U6375 ( .A1(n4904), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4905) );
  MUX2_X1 U6376 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4905), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n4907) );
  AND2_X1 U6377 ( .A1(n4907), .A2(n4906), .ZN(n5641) );
  NAND2_X1 U6378 ( .A1(n4906), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4908) );
  MUX2_X1 U6379 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4908), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n4909) );
  NAND2_X1 U6380 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n4911) );
  INV_X1 U6381 ( .A(n4913), .ZN(n4915) );
  NOR3_X1 U6382 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .A3(
        P1_IR_REG_29__SCAN_IN), .ZN(n4914) );
  NAND2_X1 U6383 ( .A1(n4915), .A2(n4914), .ZN(n9508) );
  INV_X1 U6384 ( .A(n4987), .ZN(n5042) );
  INV_X1 U6385 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n4917) );
  INV_X1 U6386 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7014) );
  OR2_X1 U6387 ( .A1(n5012), .A2(n7014), .ZN(n4924) );
  INV_X1 U6388 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n4921) );
  NAND2_X1 U6389 ( .A1(n5478), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4923) );
  NAND2_X1 U6390 ( .A1(n7824), .A2(SI_0_), .ZN(n4930) );
  XNOR2_X1 U6391 ( .A(n4930), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9514) );
  MUX2_X1 U6392 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9514), .S(n8837), .Z(n7019) );
  NAND2_X1 U6393 ( .A1(n7019), .A2(n5634), .ZN(n4936) );
  NAND2_X1 U6394 ( .A1(n6199), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n4935) );
  INV_X4 U6395 ( .A(n4952), .ZN(n8620) );
  NAND2_X1 U6396 ( .A1(n7019), .A2(n8620), .ZN(n4938) );
  INV_X1 U6397 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6309) );
  NAND3_X1 U6398 ( .A1(n4939), .A2(n4938), .A3(n4866), .ZN(n6366) );
  INV_X1 U6399 ( .A(n6366), .ZN(n4941) );
  INV_X1 U6400 ( .A(n4940), .ZN(n5674) );
  NAND2_X4 U6401 ( .A1(n5674), .A2(n6497), .ZN(n6950) );
  NAND2_X1 U6402 ( .A1(n4941), .A2(n6950), .ZN(n4942) );
  NAND2_X1 U6403 ( .A1(n6365), .A2(n4942), .ZN(n6421) );
  INV_X1 U6404 ( .A(n4964), .ZN(n4944) );
  AND2_X1 U6405 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4943) );
  NAND2_X1 U6406 ( .A1(n4944), .A2(n4943), .ZN(n5788) );
  NAND3_X1 U6407 ( .A1(n4964), .A2(SI_0_), .A3(P2_DATAO_REG_0__SCAN_IN), .ZN(
        n4945) );
  NAND2_X1 U6408 ( .A1(n5788), .A2(n4945), .ZN(n4961) );
  INV_X1 U6409 ( .A(SI_1_), .ZN(n4946) );
  MUX2_X1 U6410 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4964), .Z(n4959) );
  XNOR2_X1 U6411 ( .A(n4960), .B(n4959), .ZN(n6243) );
  INV_X1 U6412 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4948) );
  NAND2_X1 U6413 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4947) );
  OR2_X1 U6414 ( .A1(n4949), .A2(n6242), .ZN(n4950) );
  INV_X1 U6415 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n4954) );
  INV_X1 U6416 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U6417 ( .A1(n6500), .A2(n5634), .ZN(n4955) );
  INV_X2 U6418 ( .A(n6950), .ZN(n5031) );
  OR2_X1 U6419 ( .A1(n8969), .A2(n5605), .ZN(n4958) );
  NAND2_X1 U6420 ( .A1(n5606), .A2(n6500), .ZN(n4957) );
  NAND2_X1 U6421 ( .A1(n4958), .A2(n4957), .ZN(n6422) );
  NAND2_X1 U6422 ( .A1(n4960), .A2(n4959), .ZN(n4963) );
  NAND2_X1 U6423 ( .A1(n4961), .A2(SI_1_), .ZN(n4962) );
  MUX2_X1 U6424 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4964), .Z(n5002) );
  INV_X1 U6425 ( .A(SI_2_), .ZN(n4965) );
  XNOR2_X1 U6426 ( .A(n5002), .B(n4965), .ZN(n5000) );
  XNOR2_X1 U6427 ( .A(n5001), .B(n5000), .ZN(n6246) );
  OR2_X1 U6428 ( .A1(n5022), .A2(n6246), .ZN(n4969) );
  INV_X1 U6429 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6247) );
  INV_X1 U6430 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4994) );
  XNOR2_X1 U6431 ( .A(n4995), .B(n4994), .ZN(n6245) );
  OR2_X1 U6432 ( .A1(n8837), .A2(n6245), .ZN(n4967) );
  INV_X1 U6433 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n4971) );
  NAND2_X1 U6434 ( .A1(n4987), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4970) );
  OAI21_X1 U6435 ( .B1(n5010), .B2(n4971), .A(n4970), .ZN(n4972) );
  INV_X1 U6436 ( .A(n4972), .ZN(n4976) );
  INV_X1 U6437 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n4973) );
  OR2_X1 U6438 ( .A1(n5013), .A2(n4973), .ZN(n4975) );
  INV_X1 U6439 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9402) );
  OR2_X1 U6440 ( .A1(n5012), .A2(n9402), .ZN(n4974) );
  NAND2_X1 U6441 ( .A1(n9026), .A2(n5634), .ZN(n4977) );
  OAI21_X1 U6442 ( .B1(n9403), .B2(n4952), .A(n4977), .ZN(n4978) );
  XNOR2_X1 U6443 ( .A(n4978), .B(n5031), .ZN(n4981) );
  NAND2_X1 U6444 ( .A1(n5606), .A2(n9026), .ZN(n4979) );
  AND2_X1 U6445 ( .A1(n4980), .A2(n4979), .ZN(n4982) );
  NAND2_X1 U6446 ( .A1(n4981), .A2(n4982), .ZN(n4986) );
  INV_X1 U6447 ( .A(n4981), .ZN(n4984) );
  INV_X1 U6448 ( .A(n4982), .ZN(n4983) );
  NAND2_X1 U6449 ( .A1(n4984), .A2(n4983), .ZN(n4985) );
  NAND2_X1 U6450 ( .A1(n8830), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4993) );
  OR2_X1 U6451 ( .A1(n5012), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n4992) );
  INV_X1 U6452 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n4988) );
  OR2_X1 U6453 ( .A1(n5013), .A2(n4988), .ZN(n4991) );
  INV_X1 U6454 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n4989) );
  OR2_X1 U6455 ( .A1(n5010), .A2(n4989), .ZN(n4990) );
  NAND2_X1 U6456 ( .A1(n4995), .A2(n4994), .ZN(n4996) );
  NAND2_X1 U6457 ( .A1(n4996), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4998) );
  INV_X1 U6458 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4997) );
  XNOR2_X1 U6459 ( .A(n4998), .B(n4997), .ZN(n6248) );
  INV_X1 U6460 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6250) );
  OR2_X1 U6461 ( .A1(n5057), .A2(n6250), .ZN(n5006) );
  INV_X1 U6462 ( .A(SI_3_), .ZN(n4999) );
  XNOR2_X1 U6463 ( .A(n5025), .B(n4999), .ZN(n5023) );
  NAND2_X1 U6464 ( .A1(n5001), .A2(n5000), .ZN(n5004) );
  NAND2_X1 U6465 ( .A1(n5002), .A2(SI_2_), .ZN(n5003) );
  XNOR2_X1 U6466 ( .A(n5023), .B(n5024), .ZN(n6249) );
  OR2_X1 U6467 ( .A1(n5022), .A2(n6249), .ZN(n5005) );
  OAI211_X1 U6468 ( .C1(n8837), .C2(n6248), .A(n5006), .B(n5005), .ZN(n7056)
         );
  NAND2_X1 U6469 ( .A1(n7056), .A2(n8620), .ZN(n5007) );
  OAI21_X1 U6470 ( .B1(n6807), .B2(n5605), .A(n5007), .ZN(n5008) );
  XNOR2_X1 U6471 ( .A(n5008), .B(n5031), .ZN(n5034) );
  NAND2_X1 U6472 ( .A1(n7056), .A2(n5215), .ZN(n5009) );
  OAI21_X1 U6473 ( .B1(n6807), .B2(n8625), .A(n5009), .ZN(n5035) );
  XNOR2_X1 U6474 ( .A(n5034), .B(n5035), .ZN(n6534) );
  NAND2_X1 U6475 ( .A1(n8830), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5018) );
  INV_X1 U6476 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5011) );
  OR2_X1 U6477 ( .A1(n5010), .A2(n5011), .ZN(n5017) );
  XNOR2_X1 U6478 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7061) );
  OR2_X1 U6479 ( .A1(n5012), .A2(n7061), .ZN(n5016) );
  INV_X1 U6480 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5014) );
  OR2_X1 U6481 ( .A1(n5685), .A2(n5014), .ZN(n5015) );
  OR2_X1 U6482 ( .A1(n5020), .A2(n9507), .ZN(n5021) );
  XNOR2_X1 U6483 ( .A(n5021), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9863) );
  INV_X1 U6484 ( .A(n9863), .ZN(n6251) );
  INV_X1 U6485 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6253) );
  OR2_X1 U6486 ( .A1(n5057), .A2(n6253), .ZN(n5029) );
  NAND2_X1 U6487 ( .A1(n5024), .A2(n5023), .ZN(n5027) );
  NAND2_X1 U6488 ( .A1(n5025), .A2(SI_3_), .ZN(n5026) );
  INV_X1 U6489 ( .A(SI_4_), .ZN(n9674) );
  XNOR2_X1 U6490 ( .A(n5060), .B(n9674), .ZN(n5058) );
  XNOR2_X1 U6491 ( .A(n5059), .B(n5058), .ZN(n6252) );
  OR2_X1 U6492 ( .A1(n5022), .A2(n6252), .ZN(n5028) );
  OAI211_X1 U6493 ( .C1(n8837), .C2(n6251), .A(n5029), .B(n5028), .ZN(n6816)
         );
  NAND2_X1 U6494 ( .A1(n6816), .A2(n8620), .ZN(n5030) );
  OAI21_X1 U6495 ( .B1(n7045), .B2(n5605), .A(n5030), .ZN(n5032) );
  XNOR2_X1 U6496 ( .A(n5032), .B(n5031), .ZN(n5038) );
  NAND2_X1 U6497 ( .A1(n6816), .A2(n5215), .ZN(n5033) );
  OAI21_X1 U6498 ( .B1(n7045), .B2(n8625), .A(n5033), .ZN(n5039) );
  XNOR2_X1 U6499 ( .A(n5038), .B(n5039), .ZN(n6586) );
  INV_X1 U6500 ( .A(n5034), .ZN(n5036) );
  OR2_X1 U6501 ( .A1(n5036), .A2(n5035), .ZN(n6583) );
  AND2_X1 U6502 ( .A1(n6586), .A2(n6583), .ZN(n5037) );
  INV_X1 U6503 ( .A(n5038), .ZN(n5040) );
  NAND2_X1 U6504 ( .A1(n5040), .A2(n5039), .ZN(n5041) );
  NAND2_X1 U6505 ( .A1(n5477), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5051) );
  INV_X1 U6506 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5043) );
  OR2_X1 U6507 ( .A1(n5042), .A2(n5043), .ZN(n5050) );
  NAND3_X1 U6508 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5072) );
  INV_X1 U6509 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5045) );
  NAND2_X1 U6510 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5044) );
  NAND2_X1 U6511 ( .A1(n5045), .A2(n5044), .ZN(n5046) );
  NAND2_X1 U6512 ( .A1(n5072), .A2(n5046), .ZN(n6964) );
  OR2_X1 U6513 ( .A1(n5012), .A2(n6964), .ZN(n5049) );
  INV_X1 U6514 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5047) );
  OR2_X1 U6515 ( .A1(n5685), .A2(n5047), .ZN(n5048) );
  NOR2_X1 U6516 ( .A1(n5053), .A2(n9507), .ZN(n5054) );
  MUX2_X1 U6517 ( .A(n9507), .B(n5054), .S(P1_IR_REG_5__SCAN_IN), .Z(n5055) );
  INV_X1 U6518 ( .A(n5055), .ZN(n5056) );
  AND2_X1 U6519 ( .A1(n5052), .A2(n5056), .ZN(n9867) );
  INV_X1 U6520 ( .A(n9867), .ZN(n6254) );
  OR2_X1 U6521 ( .A1(n5057), .A2(n4428), .ZN(n5063) );
  NAND2_X1 U6522 ( .A1(n5060), .A2(SI_4_), .ZN(n5061) );
  INV_X1 U6523 ( .A(SI_5_), .ZN(n9649) );
  XNOR2_X1 U6524 ( .A(n5080), .B(n5079), .ZN(n6255) );
  OR2_X1 U6525 ( .A1(n5022), .A2(n6255), .ZN(n5062) );
  OAI211_X1 U6526 ( .C1(n8837), .C2(n6254), .A(n5063), .B(n5062), .ZN(n9934)
         );
  NAND2_X1 U6527 ( .A1(n9934), .A2(n8620), .ZN(n5064) );
  OAI21_X1 U6528 ( .B1(n7129), .B2(n5605), .A(n5064), .ZN(n5065) );
  XNOR2_X1 U6529 ( .A(n5065), .B(n5031), .ZN(n6885) );
  OR2_X1 U6530 ( .A1(n7129), .A2(n8625), .ZN(n5067) );
  NAND2_X1 U6531 ( .A1(n9934), .A2(n5215), .ZN(n5066) );
  NAND2_X1 U6532 ( .A1(n5067), .A2(n5066), .ZN(n6887) );
  INV_X1 U6533 ( .A(n6887), .ZN(n5068) );
  NAND2_X1 U6534 ( .A1(n6885), .A2(n5068), .ZN(n5069) );
  NAND2_X1 U6535 ( .A1(n5477), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5077) );
  INV_X1 U6536 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7134) );
  OR2_X1 U6537 ( .A1(n5042), .A2(n7134), .ZN(n5076) );
  INV_X1 U6538 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5070) );
  OR2_X1 U6539 ( .A1(n5685), .A2(n5070), .ZN(n5075) );
  INV_X1 U6540 ( .A(n5072), .ZN(n5071) );
  NAND2_X1 U6541 ( .A1(n5071), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5099) );
  INV_X1 U6542 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6926) );
  NAND2_X1 U6543 ( .A1(n5072), .A2(n6926), .ZN(n5073) );
  NAND2_X1 U6544 ( .A1(n5099), .A2(n5073), .ZN(n7133) );
  OR2_X1 U6545 ( .A1(n5012), .A2(n7133), .ZN(n5074) );
  NAND2_X1 U6546 ( .A1(n5052), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5078) );
  XNOR2_X1 U6547 ( .A(n5078), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9892) );
  INV_X1 U6548 ( .A(n9892), .ZN(n6257) );
  NAND2_X1 U6549 ( .A1(n5081), .A2(SI_5_), .ZN(n5082) );
  MUX2_X1 U6550 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7824), .Z(n5108) );
  INV_X1 U6551 ( .A(SI_6_), .ZN(n5084) );
  XNOR2_X1 U6552 ( .A(n5108), .B(n5084), .ZN(n5106) );
  XNOR2_X1 U6553 ( .A(n5107), .B(n5106), .ZN(n6258) );
  OR2_X1 U6554 ( .A1(n5022), .A2(n6258), .ZN(n5086) );
  INV_X1 U6555 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6259) );
  OR2_X1 U6556 ( .A1(n5057), .A2(n6259), .ZN(n5085) );
  NAND2_X1 U6557 ( .A1(n7139), .A2(n8620), .ZN(n5087) );
  OAI21_X1 U6558 ( .B1(n7233), .B2(n5605), .A(n5087), .ZN(n5088) );
  XNOR2_X1 U6559 ( .A(n5088), .B(n6950), .ZN(n5091) );
  NAND2_X1 U6560 ( .A1(n7139), .A2(n5215), .ZN(n5089) );
  OAI21_X1 U6561 ( .B1(n7233), .B2(n8625), .A(n5089), .ZN(n5090) );
  OR2_X1 U6562 ( .A1(n5091), .A2(n5090), .ZN(n6874) );
  NAND2_X1 U6563 ( .A1(n5091), .A2(n5090), .ZN(n5092) );
  NAND2_X1 U6564 ( .A1(n6874), .A2(n5092), .ZN(n6919) );
  INV_X1 U6565 ( .A(n6885), .ZN(n5093) );
  AND2_X1 U6566 ( .A1(n5093), .A2(n6887), .ZN(n5094) );
  NOR2_X1 U6567 ( .A1(n6919), .A2(n5094), .ZN(n5095) );
  NAND2_X1 U6568 ( .A1(n6873), .A2(n6874), .ZN(n5119) );
  NAND2_X1 U6569 ( .A1(n5477), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5104) );
  INV_X1 U6570 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7244) );
  OR2_X1 U6571 ( .A1(n5042), .A2(n7244), .ZN(n5103) );
  INV_X1 U6572 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5096) );
  OR2_X1 U6573 ( .A1(n5685), .A2(n5096), .ZN(n5102) );
  INV_X1 U6574 ( .A(n5099), .ZN(n5097) );
  INV_X1 U6575 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5098) );
  NAND2_X1 U6576 ( .A1(n5099), .A2(n5098), .ZN(n5100) );
  NAND2_X1 U6577 ( .A1(n5122), .A2(n5100), .ZN(n7243) );
  OR2_X1 U6578 ( .A1(n5012), .A2(n7243), .ZN(n5101) );
  OR2_X1 U6579 ( .A1(n5052), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5134) );
  NAND2_X1 U6580 ( .A1(n5134), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5105) );
  XNOR2_X1 U6581 ( .A(n5105), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6337) );
  INV_X1 U6582 ( .A(n6337), .ZN(n6261) );
  INV_X1 U6583 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6263) );
  OR2_X1 U6584 ( .A1(n5057), .A2(n6263), .ZN(n5112) );
  NAND2_X1 U6585 ( .A1(n5108), .A2(SI_6_), .ZN(n5109) );
  MUX2_X1 U6586 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7824), .Z(n5130) );
  INV_X1 U6587 ( .A(SI_7_), .ZN(n5110) );
  XNOR2_X1 U6588 ( .A(n5130), .B(n5110), .ZN(n5129) );
  OR2_X1 U6589 ( .A1(n5022), .A2(n6262), .ZN(n5111) );
  NAND2_X1 U6590 ( .A1(n7246), .A2(n8620), .ZN(n5113) );
  OAI21_X1 U6591 ( .B1(n7128), .B2(n5605), .A(n5113), .ZN(n5114) );
  XNOR2_X1 U6592 ( .A(n5114), .B(n6950), .ZN(n5117) );
  NAND2_X1 U6593 ( .A1(n7246), .A2(n5215), .ZN(n5115) );
  OAI21_X1 U6594 ( .B1(n7128), .B2(n8625), .A(n5115), .ZN(n5116) );
  OR2_X1 U6595 ( .A1(n5117), .A2(n5116), .ZN(n5120) );
  NAND2_X1 U6596 ( .A1(n5117), .A2(n5116), .ZN(n5118) );
  AND2_X1 U6597 ( .A1(n5120), .A2(n5118), .ZN(n6875) );
  NAND2_X1 U6598 ( .A1(n5119), .A2(n6875), .ZN(n6877) );
  NAND2_X1 U6599 ( .A1(n6877), .A2(n5120), .ZN(n5143) );
  NAND2_X1 U6600 ( .A1(n5478), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5128) );
  INV_X1 U6601 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7119) );
  OR2_X1 U6602 ( .A1(n5042), .A2(n7119), .ZN(n5127) );
  INV_X1 U6603 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7095) );
  NAND2_X1 U6604 ( .A1(n5122), .A2(n7095), .ZN(n5123) );
  NAND2_X1 U6605 ( .A1(n5162), .A2(n5123), .ZN(n7118) );
  OR2_X1 U6606 ( .A1(n5012), .A2(n7118), .ZN(n5126) );
  INV_X1 U6607 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5124) );
  OR2_X1 U6608 ( .A1(n5010), .A2(n5124), .ZN(n5125) );
  OR2_X1 U6609 ( .A1(n7287), .A2(n8625), .ZN(n5140) );
  MUX2_X1 U6610 ( .A(n6269), .B(n6272), .S(n7824), .Z(n5131) );
  NAND2_X1 U6611 ( .A1(n5131), .A2(n9727), .ZN(n5149) );
  INV_X1 U6612 ( .A(n5131), .ZN(n5132) );
  NAND2_X1 U6613 ( .A1(n5132), .A2(SI_8_), .ZN(n5133) );
  NAND2_X1 U6614 ( .A1(n5149), .A2(n5133), .ZN(n5148) );
  XNOR2_X1 U6615 ( .A(n5147), .B(n5148), .ZN(n6267) );
  AND2_X1 U6616 ( .A1(n8840), .A2(n6267), .ZN(n5138) );
  NOR2_X1 U6617 ( .A1(n5134), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5155) );
  OR2_X1 U6618 ( .A1(n5155), .A2(n9507), .ZN(n5135) );
  XNOR2_X1 U6619 ( .A(n5135), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9905) );
  INV_X1 U6620 ( .A(n9905), .ZN(n6270) );
  NOR2_X1 U6621 ( .A1(n8837), .A2(n6270), .ZN(n5137) );
  NOR2_X1 U6622 ( .A1(n5057), .A2(n6272), .ZN(n5136) );
  NAND2_X1 U6623 ( .A1(n7294), .A2(n5215), .ZN(n5139) );
  AND2_X1 U6624 ( .A1(n5140), .A2(n5139), .ZN(n5144) );
  NAND2_X1 U6625 ( .A1(n5143), .A2(n5144), .ZN(n7091) );
  NAND2_X1 U6626 ( .A1(n7294), .A2(n8620), .ZN(n5141) );
  OAI21_X1 U6627 ( .B1(n7287), .B2(n5605), .A(n5141), .ZN(n5142) );
  XNOR2_X1 U6628 ( .A(n5142), .B(n6950), .ZN(n7093) );
  INV_X1 U6629 ( .A(n5144), .ZN(n5145) );
  INV_X1 U6630 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5150) );
  MUX2_X1 U6631 ( .A(n5150), .B(n6275), .S(n7824), .Z(n5151) );
  NAND2_X1 U6632 ( .A1(n5151), .A2(n9705), .ZN(n5178) );
  INV_X1 U6633 ( .A(n5151), .ZN(n5152) );
  NAND2_X1 U6634 ( .A1(n5152), .A2(SI_9_), .ZN(n5153) );
  NAND2_X1 U6635 ( .A1(n6273), .A2(n8840), .ZN(n5160) );
  NAND2_X1 U6636 ( .A1(n5155), .A2(n5154), .ZN(n5157) );
  NAND2_X1 U6637 ( .A1(n5157), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5156) );
  MUX2_X1 U6638 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5156), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n5158) );
  AOI22_X1 U6639 ( .A1(n5427), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5426), .B2(
        n6400), .ZN(n5159) );
  NAND2_X1 U6640 ( .A1(n7335), .A2(n8620), .ZN(n5169) );
  NAND2_X1 U6641 ( .A1(n8830), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6642 ( .A1(n5477), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6643 ( .A1(n5162), .A2(n5161), .ZN(n5163) );
  NAND2_X1 U6644 ( .A1(n5186), .A2(n5163), .ZN(n7288) );
  OR2_X1 U6645 ( .A1(n4313), .A2(n7288), .ZN(n5165) );
  INV_X1 U6646 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6217) );
  OR2_X1 U6647 ( .A1(n5685), .A2(n6217), .ZN(n5164) );
  NAND4_X1 U6648 ( .A1(n5167), .A2(n5166), .A3(n5165), .A4(n5164), .ZN(n9019)
         );
  NAND2_X1 U6649 ( .A1(n9019), .A2(n5215), .ZN(n5168) );
  NAND2_X1 U6650 ( .A1(n5169), .A2(n5168), .ZN(n5170) );
  XNOR2_X1 U6651 ( .A(n5170), .B(n5031), .ZN(n5172) );
  AOI22_X1 U6652 ( .A1(n7335), .A2(n5634), .B1(n5606), .B2(n9019), .ZN(n5171)
         );
  NAND2_X1 U6653 ( .A1(n5172), .A2(n5171), .ZN(n5175) );
  OR2_X1 U6654 ( .A1(n5172), .A2(n5171), .ZN(n5173) );
  NAND2_X1 U6655 ( .A1(n5175), .A2(n5173), .ZN(n7225) );
  INV_X1 U6656 ( .A(n7225), .ZN(n5174) );
  NAND2_X1 U6657 ( .A1(n7222), .A2(n5175), .ZN(n7370) );
  INV_X1 U6658 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5179) );
  MUX2_X1 U6659 ( .A(n5179), .B(n6280), .S(n7824), .Z(n5180) );
  NAND2_X1 U6660 ( .A1(n5180), .A2(n9651), .ZN(n5199) );
  INV_X1 U6661 ( .A(n5180), .ZN(n5181) );
  NAND2_X1 U6662 ( .A1(n5181), .A2(SI_10_), .ZN(n5182) );
  NAND2_X1 U6663 ( .A1(n6278), .A2(n8840), .ZN(n5185) );
  NAND2_X1 U6664 ( .A1(n5202), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5183) );
  XNOR2_X1 U6665 ( .A(n5183), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6574) );
  AOI22_X1 U6666 ( .A1(n5427), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5426), .B2(
        n6574), .ZN(n5184) );
  NAND2_X1 U6667 ( .A1(n9735), .A2(n8620), .ZN(n5194) );
  NAND2_X1 U6668 ( .A1(n5477), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5192) );
  INV_X1 U6669 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7340) );
  OR2_X1 U6670 ( .A1(n5042), .A2(n7340), .ZN(n5191) );
  NAND2_X1 U6671 ( .A1(n5186), .A2(n6393), .ZN(n5187) );
  NAND2_X1 U6672 ( .A1(n5209), .A2(n5187), .ZN(n7374) );
  OR2_X1 U6673 ( .A1(n5012), .A2(n7374), .ZN(n5190) );
  INV_X1 U6674 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5188) );
  OR2_X1 U6675 ( .A1(n5685), .A2(n5188), .ZN(n5189) );
  INV_X1 U6676 ( .A(n9799), .ZN(n9018) );
  NAND2_X1 U6677 ( .A1(n9018), .A2(n5215), .ZN(n5193) );
  NAND2_X1 U6678 ( .A1(n5194), .A2(n5193), .ZN(n5195) );
  XNOR2_X1 U6679 ( .A(n5195), .B(n6950), .ZN(n5220) );
  NOR2_X1 U6680 ( .A1(n9799), .A2(n8625), .ZN(n5196) );
  AOI21_X1 U6681 ( .B1(n9735), .B2(n5634), .A(n5196), .ZN(n5221) );
  XNOR2_X1 U6682 ( .A(n5220), .B(n5221), .ZN(n7371) );
  NAND2_X1 U6683 ( .A1(n7370), .A2(n7371), .ZN(n7369) );
  NAND2_X1 U6684 ( .A1(n5198), .A2(n5197), .ZN(n5200) );
  NAND2_X1 U6685 ( .A1(n5200), .A2(n5199), .ZN(n5226) );
  MUX2_X1 U6686 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n7824), .Z(n5227) );
  INV_X1 U6687 ( .A(SI_11_), .ZN(n5201) );
  XNOR2_X1 U6688 ( .A(n5227), .B(n5201), .ZN(n5224) );
  XNOR2_X1 U6689 ( .A(n5226), .B(n5224), .ZN(n6282) );
  NAND2_X1 U6690 ( .A1(n6282), .A2(n8840), .ZN(n5205) );
  OAI21_X1 U6691 ( .B1(n5202), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5203) );
  XNOR2_X1 U6692 ( .A(n5203), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6575) );
  AOI22_X1 U6693 ( .A1(n5427), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5426), .B2(
        n6575), .ZN(n5204) );
  NAND2_X1 U6694 ( .A1(n9809), .A2(n8620), .ZN(n5217) );
  INV_X1 U6695 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9791) );
  OR2_X1 U6696 ( .A1(n5042), .A2(n9791), .ZN(n5214) );
  NAND2_X1 U6697 ( .A1(n5477), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5213) );
  INV_X1 U6698 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5206) );
  OR2_X1 U6699 ( .A1(n5685), .A2(n5206), .ZN(n5212) );
  INV_X1 U6700 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5208) );
  NAND2_X1 U6701 ( .A1(n5209), .A2(n5208), .ZN(n5210) );
  NAND2_X1 U6702 ( .A1(n5239), .A2(n5210), .ZN(n9790) );
  OR2_X1 U6703 ( .A1(n5012), .A2(n9790), .ZN(n5211) );
  NAND4_X1 U6704 ( .A1(n5214), .A2(n5213), .A3(n5212), .A4(n5211), .ZN(n9017)
         );
  NAND2_X1 U6705 ( .A1(n9017), .A2(n5215), .ZN(n5216) );
  NAND2_X1 U6706 ( .A1(n5217), .A2(n5216), .ZN(n5218) );
  XNOR2_X1 U6707 ( .A(n5218), .B(n6950), .ZN(n5251) );
  AND2_X1 U6708 ( .A1(n5606), .A2(n9017), .ZN(n5219) );
  AOI21_X1 U6709 ( .B1(n9809), .B2(n5634), .A(n5219), .ZN(n5249) );
  XNOR2_X1 U6710 ( .A(n5251), .B(n5249), .ZN(n7503) );
  INV_X1 U6711 ( .A(n5220), .ZN(n5222) );
  NAND2_X1 U6712 ( .A1(n5222), .A2(n5221), .ZN(n7504) );
  AND2_X1 U6713 ( .A1(n7503), .A2(n7504), .ZN(n5223) );
  INV_X1 U6714 ( .A(n5224), .ZN(n5225) );
  NAND2_X1 U6715 ( .A1(n5227), .A2(SI_11_), .ZN(n5228) );
  INV_X1 U6716 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5229) );
  MUX2_X1 U6717 ( .A(n6295), .B(n5229), .S(n7824), .Z(n5230) );
  INV_X1 U6718 ( .A(n5230), .ZN(n5231) );
  NAND2_X1 U6719 ( .A1(n5231), .A2(SI_12_), .ZN(n5232) );
  NAND2_X1 U6720 ( .A1(n5259), .A2(n5232), .ZN(n5257) );
  XNOR2_X1 U6721 ( .A(n5258), .B(n5257), .ZN(n6286) );
  NAND2_X1 U6722 ( .A1(n6286), .A2(n8840), .ZN(n5236) );
  NAND2_X1 U6723 ( .A1(n5233), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5234) );
  XNOR2_X1 U6724 ( .A(n5234), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6847) );
  AOI22_X1 U6725 ( .A1(n5427), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5426), .B2(
        n6847), .ZN(n5235) );
  NAND2_X1 U6726 ( .A1(n7548), .A2(n8620), .ZN(n5246) );
  NAND2_X1 U6727 ( .A1(n5477), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5244) );
  INV_X1 U6728 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7523) );
  OR2_X1 U6729 ( .A1(n5042), .A2(n7523), .ZN(n5243) );
  INV_X1 U6730 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U6731 ( .A1(n5239), .A2(n5238), .ZN(n5240) );
  NAND2_X1 U6732 ( .A1(n5269), .A2(n5240), .ZN(n7522) );
  OR2_X1 U6733 ( .A1(n4313), .A2(n7522), .ZN(n5242) );
  INV_X1 U6734 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6567) );
  OR2_X1 U6735 ( .A1(n5685), .A2(n6567), .ZN(n5241) );
  INV_X1 U6736 ( .A(n9797), .ZN(n9773) );
  NAND2_X1 U6737 ( .A1(n9773), .A2(n5215), .ZN(n5245) );
  NAND2_X1 U6738 ( .A1(n5246), .A2(n5245), .ZN(n5247) );
  XNOR2_X1 U6739 ( .A(n5247), .B(n6950), .ZN(n5253) );
  NOR2_X1 U6740 ( .A1(n9797), .A2(n8625), .ZN(n5248) );
  AOI21_X1 U6741 ( .B1(n7548), .B2(n5634), .A(n5248), .ZN(n5254) );
  XNOR2_X1 U6742 ( .A(n5253), .B(n5254), .ZN(n7448) );
  INV_X1 U6743 ( .A(n5249), .ZN(n5250) );
  NAND2_X1 U6744 ( .A1(n5251), .A2(n5250), .ZN(n7449) );
  AND2_X1 U6745 ( .A1(n7448), .A2(n7449), .ZN(n5252) );
  NAND2_X1 U6746 ( .A1(n7502), .A2(n5252), .ZN(n7447) );
  INV_X1 U6747 ( .A(n5253), .ZN(n5255) );
  NAND2_X1 U6748 ( .A1(n5255), .A2(n5254), .ZN(n5256) );
  INV_X1 U6749 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5260) );
  MUX2_X1 U6750 ( .A(n6346), .B(n5260), .S(n7824), .Z(n5261) );
  INV_X1 U6751 ( .A(n5261), .ZN(n5262) );
  NAND2_X1 U6752 ( .A1(n5262), .A2(SI_13_), .ZN(n5263) );
  XNOR2_X1 U6753 ( .A(n5286), .B(n5285), .ZN(n6304) );
  NAND2_X1 U6754 ( .A1(n6304), .A2(n8840), .ZN(n5267) );
  OR2_X1 U6755 ( .A1(n5264), .A2(n9507), .ZN(n5265) );
  XNOR2_X1 U6756 ( .A(n5265), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7199) );
  AOI22_X1 U6757 ( .A1(n5427), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5426), .B2(
        n7199), .ZN(n5266) );
  NAND2_X1 U6758 ( .A1(n9779), .A2(n8620), .ZN(n5277) );
  NAND2_X1 U6759 ( .A1(n5477), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5275) );
  INV_X1 U6760 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6848) );
  OR2_X1 U6761 ( .A1(n5042), .A2(n6848), .ZN(n5274) );
  NAND2_X1 U6762 ( .A1(n5269), .A2(n5268), .ZN(n5270) );
  NAND2_X1 U6763 ( .A1(n5298), .A2(n5270), .ZN(n9765) );
  OR2_X1 U6764 ( .A1(n5012), .A2(n9765), .ZN(n5273) );
  INV_X1 U6765 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n5271) );
  OR2_X1 U6766 ( .A1(n5685), .A2(n5271), .ZN(n5272) );
  NAND4_X1 U6767 ( .A1(n5275), .A2(n5274), .A3(n5273), .A4(n5272), .ZN(n9016)
         );
  NAND2_X1 U6768 ( .A1(n9016), .A2(n5215), .ZN(n5276) );
  NAND2_X1 U6769 ( .A1(n5277), .A2(n5276), .ZN(n5278) );
  XNOR2_X1 U6770 ( .A(n5278), .B(n5031), .ZN(n5281) );
  AND2_X1 U6771 ( .A1(n5606), .A2(n9016), .ZN(n5279) );
  AOI21_X1 U6772 ( .B1(n9779), .B2(n5634), .A(n5279), .ZN(n5282) );
  INV_X1 U6773 ( .A(n5281), .ZN(n5284) );
  INV_X1 U6774 ( .A(n5282), .ZN(n5283) );
  NAND2_X1 U6775 ( .A1(n5284), .A2(n5283), .ZN(n7473) );
  MUX2_X1 U6776 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7824), .Z(n5316) );
  INV_X1 U6777 ( .A(SI_14_), .ZN(n5288) );
  XNOR2_X1 U6778 ( .A(n5316), .B(n5288), .ZN(n5313) );
  XNOR2_X1 U6779 ( .A(n5315), .B(n5313), .ZN(n6347) );
  NAND2_X1 U6780 ( .A1(n6347), .A2(n8840), .ZN(n5295) );
  OR2_X1 U6781 ( .A1(n5289), .A2(n9507), .ZN(n5292) );
  INV_X1 U6782 ( .A(n5292), .ZN(n5290) );
  NAND2_X1 U6783 ( .A1(n5290), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6784 ( .A1(n5292), .A2(n5291), .ZN(n5321) );
  AOI22_X1 U6785 ( .A1(n5427), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5426), .B2(
        n7439), .ZN(n5294) );
  NAND2_X1 U6786 ( .A1(n9486), .A2(n8620), .ZN(n5306) );
  NAND2_X1 U6787 ( .A1(n5477), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U6788 ( .A1(n8830), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5303) );
  INV_X1 U6789 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5297) );
  NAND2_X1 U6790 ( .A1(n5298), .A2(n5297), .ZN(n5299) );
  NAND2_X1 U6791 ( .A1(n5327), .A2(n5299), .ZN(n7576) );
  OR2_X1 U6792 ( .A1(n4313), .A2(n7576), .ZN(n5302) );
  INV_X1 U6793 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5300) );
  OR2_X1 U6794 ( .A1(n5685), .A2(n5300), .ZN(n5301) );
  NAND4_X1 U6795 ( .A1(n5304), .A2(n5303), .A3(n5302), .A4(n5301), .ZN(n9770)
         );
  NAND2_X1 U6796 ( .A1(n9770), .A2(n5215), .ZN(n5305) );
  NAND2_X1 U6797 ( .A1(n5306), .A2(n5305), .ZN(n5307) );
  XNOR2_X1 U6798 ( .A(n5307), .B(n6950), .ZN(n5311) );
  INV_X1 U6799 ( .A(n5311), .ZN(n5308) );
  NAND2_X1 U6800 ( .A1(n9486), .A2(n5215), .ZN(n5310) );
  NAND2_X1 U6801 ( .A1(n5606), .A2(n9770), .ZN(n5309) );
  NAND2_X1 U6802 ( .A1(n5310), .A2(n5309), .ZN(n7571) );
  NAND2_X1 U6803 ( .A1(n7568), .A2(n7571), .ZN(n5312) );
  INV_X1 U6804 ( .A(n5313), .ZN(n5314) );
  NAND2_X1 U6805 ( .A1(n5316), .A2(SI_14_), .ZN(n5317) );
  MUX2_X1 U6806 ( .A(n6373), .B(n6371), .S(n7824), .Z(n5318) );
  INV_X1 U6807 ( .A(n5318), .ZN(n5319) );
  NAND2_X1 U6808 ( .A1(n5319), .A2(SI_15_), .ZN(n5320) );
  NAND2_X1 U6809 ( .A1(n5341), .A2(n5320), .ZN(n5339) );
  XNOR2_X1 U6810 ( .A(n5340), .B(n5339), .ZN(n6370) );
  NAND2_X1 U6811 ( .A1(n6370), .A2(n8840), .ZN(n5325) );
  NAND2_X1 U6812 ( .A1(n5321), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5323) );
  INV_X1 U6813 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5322) );
  XNOR2_X1 U6814 ( .A(n5323), .B(n5322), .ZN(n9049) );
  INV_X1 U6815 ( .A(n9049), .ZN(n7443) );
  AOI22_X1 U6816 ( .A1(n5427), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5426), .B2(
        n7443), .ZN(n5324) );
  NAND2_X1 U6817 ( .A1(n9393), .A2(n8620), .ZN(n5334) );
  NAND2_X1 U6818 ( .A1(n5477), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U6819 ( .A1(n5478), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5331) );
  INV_X1 U6820 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6821 ( .A1(n5327), .A2(n5326), .ZN(n5328) );
  NAND2_X1 U6822 ( .A1(n5353), .A2(n5328), .ZN(n9390) );
  OR2_X1 U6823 ( .A1(n5012), .A2(n9390), .ZN(n5330) );
  INV_X1 U6824 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9391) );
  OR2_X1 U6825 ( .A1(n5042), .A2(n9391), .ZN(n5329) );
  NAND4_X1 U6826 ( .A1(n5332), .A2(n5331), .A3(n5330), .A4(n5329), .ZN(n9107)
         );
  NAND2_X1 U6827 ( .A1(n9107), .A2(n5215), .ZN(n5333) );
  NAND2_X1 U6828 ( .A1(n5334), .A2(n5333), .ZN(n5335) );
  XNOR2_X1 U6829 ( .A(n5335), .B(n6950), .ZN(n5338) );
  NAND2_X1 U6830 ( .A1(n9393), .A2(n5215), .ZN(n5337) );
  NAND2_X1 U6831 ( .A1(n5606), .A2(n9107), .ZN(n5336) );
  NAND2_X1 U6832 ( .A1(n5337), .A2(n5336), .ZN(n8730) );
  INV_X1 U6833 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5342) );
  MUX2_X1 U6834 ( .A(n5342), .B(n6455), .S(n7824), .Z(n5344) );
  INV_X1 U6835 ( .A(SI_16_), .ZN(n5343) );
  INV_X1 U6836 ( .A(n5344), .ZN(n5345) );
  NAND2_X1 U6837 ( .A1(n5345), .A2(SI_16_), .ZN(n5346) );
  XNOR2_X1 U6838 ( .A(n5369), .B(n5368), .ZN(n6419) );
  NAND2_X1 U6839 ( .A1(n6419), .A2(n8840), .ZN(n5350) );
  NAND2_X1 U6840 ( .A1(n5347), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5348) );
  XNOR2_X1 U6841 ( .A(n5348), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9068) );
  AOI22_X1 U6842 ( .A1(n5427), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5426), .B2(
        n9068), .ZN(n5349) );
  NAND2_X1 U6843 ( .A1(n9481), .A2(n8620), .ZN(n5361) );
  NAND2_X1 U6844 ( .A1(n5477), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5359) );
  INV_X1 U6845 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9368) );
  OR2_X1 U6846 ( .A1(n5042), .A2(n9368), .ZN(n5358) );
  INV_X1 U6847 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U6848 ( .A1(n5353), .A2(n5352), .ZN(n5354) );
  NAND2_X1 U6849 ( .A1(n5379), .A2(n5354), .ZN(n9367) );
  OR2_X1 U6850 ( .A1(n4313), .A2(n9367), .ZN(n5357) );
  INV_X1 U6851 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n5355) );
  OR2_X1 U6852 ( .A1(n5685), .A2(n5355), .ZN(n5356) );
  INV_X1 U6853 ( .A(n9359), .ZN(n9385) );
  NAND2_X1 U6854 ( .A1(n9385), .A2(n5215), .ZN(n5360) );
  NAND2_X1 U6855 ( .A1(n5361), .A2(n5360), .ZN(n5362) );
  XNOR2_X1 U6856 ( .A(n5362), .B(n6950), .ZN(n5364) );
  NOR2_X1 U6857 ( .A1(n9359), .A2(n8625), .ZN(n5363) );
  AOI21_X1 U6858 ( .B1(n9481), .B2(n5634), .A(n5363), .ZN(n5365) );
  XNOR2_X1 U6859 ( .A(n5364), .B(n5365), .ZN(n8661) );
  INV_X1 U6860 ( .A(n5364), .ZN(n5366) );
  NAND2_X1 U6861 ( .A1(n5366), .A2(n5365), .ZN(n5367) );
  NAND2_X1 U6862 ( .A1(n5369), .A2(n5368), .ZN(n5371) );
  MUX2_X1 U6863 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n7824), .Z(n5394) );
  XNOR2_X1 U6864 ( .A(n5394), .B(n9618), .ZN(n5393) );
  XNOR2_X1 U6865 ( .A(n5397), .B(n5393), .ZN(n6450) );
  NAND2_X1 U6866 ( .A1(n6450), .A2(n8840), .ZN(n5378) );
  INV_X1 U6867 ( .A(n5372), .ZN(n5373) );
  NAND2_X1 U6868 ( .A1(n5373), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5375) );
  INV_X1 U6869 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5374) );
  OR2_X1 U6870 ( .A1(n5375), .A2(n5374), .ZN(n5376) );
  NAND2_X1 U6871 ( .A1(n5375), .A2(n5374), .ZN(n5398) );
  AOI22_X1 U6872 ( .A1(n5427), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5426), .B2(
        n9083), .ZN(n5377) );
  NAND2_X1 U6873 ( .A1(n4953), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5385) );
  INV_X1 U6874 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9069) );
  OR2_X1 U6875 ( .A1(n5042), .A2(n9069), .ZN(n5384) );
  INV_X1 U6876 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8672) );
  NAND2_X1 U6877 ( .A1(n5379), .A2(n8672), .ZN(n5380) );
  NAND2_X1 U6878 ( .A1(n5404), .A2(n5380), .ZN(n9352) );
  OR2_X1 U6879 ( .A1(n5012), .A2(n9352), .ZN(n5383) );
  INV_X1 U6880 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n5381) );
  OR2_X1 U6881 ( .A1(n5685), .A2(n5381), .ZN(n5382) );
  OAI22_X1 U6882 ( .A1(n9351), .A2(n4952), .B1(n9376), .B2(n5605), .ZN(n5386)
         );
  XNOR2_X1 U6883 ( .A(n5386), .B(n5031), .ZN(n5391) );
  OR2_X1 U6884 ( .A1(n9351), .A2(n5605), .ZN(n5388) );
  NAND2_X1 U6885 ( .A1(n9332), .A2(n5606), .ZN(n5387) );
  NAND2_X1 U6886 ( .A1(n5388), .A2(n5387), .ZN(n5389) );
  XNOR2_X1 U6887 ( .A(n5391), .B(n5389), .ZN(n8670) );
  INV_X1 U6888 ( .A(n5389), .ZN(n5390) );
  NAND2_X1 U6889 ( .A1(n5391), .A2(n5390), .ZN(n5392) );
  INV_X1 U6890 ( .A(n5393), .ZN(n5396) );
  NAND2_X1 U6891 ( .A1(n5394), .A2(SI_17_), .ZN(n5395) );
  MUX2_X1 U6892 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7824), .Z(n5421) );
  XNOR2_X1 U6893 ( .A(n5421), .B(SI_18_), .ZN(n5418) );
  XNOR2_X1 U6894 ( .A(n5420), .B(n5418), .ZN(n6594) );
  NAND2_X1 U6895 ( .A1(n6594), .A2(n8840), .ZN(n5401) );
  NAND2_X1 U6896 ( .A1(n5398), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5399) );
  XNOR2_X1 U6897 ( .A(n5399), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9911) );
  AOI22_X1 U6898 ( .A1(n5427), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5426), .B2(
        n9911), .ZN(n5400) );
  NAND2_X1 U6899 ( .A1(n9468), .A2(n8620), .ZN(n5411) );
  NAND2_X1 U6900 ( .A1(n5477), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5409) );
  INV_X1 U6901 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9341) );
  OR2_X1 U6902 ( .A1(n5042), .A2(n9341), .ZN(n5408) );
  INV_X1 U6903 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U6904 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  NAND2_X1 U6905 ( .A1(n5432), .A2(n5405), .ZN(n9340) );
  OR2_X1 U6906 ( .A1(n4313), .A2(n9340), .ZN(n5407) );
  INV_X1 U6907 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9081) );
  OR2_X1 U6908 ( .A1(n5685), .A2(n9081), .ZN(n5406) );
  NAND2_X1 U6909 ( .A1(n9322), .A2(n5215), .ZN(n5410) );
  NAND2_X1 U6910 ( .A1(n5411), .A2(n5410), .ZN(n5412) );
  XNOR2_X1 U6911 ( .A(n5412), .B(n5031), .ZN(n5416) );
  NAND2_X1 U6912 ( .A1(n9468), .A2(n5215), .ZN(n5414) );
  NAND2_X1 U6913 ( .A1(n9322), .A2(n5606), .ZN(n5413) );
  NAND2_X1 U6914 ( .A1(n5414), .A2(n5413), .ZN(n8706) );
  NAND2_X1 U6915 ( .A1(n5421), .A2(SI_18_), .ZN(n5422) );
  MUX2_X1 U6916 ( .A(n6747), .B(n6745), .S(n7824), .Z(n5423) );
  NAND2_X1 U6917 ( .A1(n5423), .A2(n9614), .ZN(n5448) );
  INV_X1 U6918 ( .A(n5423), .ZN(n5424) );
  NAND2_X1 U6919 ( .A1(n5424), .A2(SI_19_), .ZN(n5425) );
  NAND2_X1 U6920 ( .A1(n5448), .A2(n5425), .ZN(n5447) );
  XNOR2_X1 U6921 ( .A(n5446), .B(n5447), .ZN(n6744) );
  NAND2_X1 U6922 ( .A1(n6744), .A2(n8840), .ZN(n5429) );
  AOI22_X1 U6923 ( .A1(n5427), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9161), .B2(
        n5426), .ZN(n5428) );
  NAND2_X1 U6924 ( .A1(n9462), .A2(n8620), .ZN(n5439) );
  INV_X1 U6925 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6926 ( .A1(n5432), .A2(n5431), .ZN(n5433) );
  NAND2_X1 U6927 ( .A1(n5455), .A2(n5433), .ZN(n9315) );
  OR2_X1 U6928 ( .A1(n9315), .A2(n5012), .ZN(n5437) );
  NAND2_X1 U6929 ( .A1(n8830), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U6930 ( .A1(n5477), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5435) );
  INV_X1 U6931 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9084) );
  OR2_X1 U6932 ( .A1(n5685), .A2(n9084), .ZN(n5434) );
  NAND4_X1 U6933 ( .A1(n5437), .A2(n5436), .A3(n5435), .A4(n5434), .ZN(n9333)
         );
  NAND2_X1 U6934 ( .A1(n9333), .A2(n5215), .ZN(n5438) );
  NAND2_X1 U6935 ( .A1(n5439), .A2(n5438), .ZN(n5440) );
  XNOR2_X1 U6936 ( .A(n5440), .B(n6950), .ZN(n5442) );
  AND2_X1 U6937 ( .A1(n5606), .A2(n9333), .ZN(n5441) );
  AOI21_X1 U6938 ( .B1(n9462), .B2(n5634), .A(n5441), .ZN(n5443) );
  XNOR2_X1 U6939 ( .A(n5442), .B(n5443), .ZN(n8610) );
  INV_X1 U6940 ( .A(n5442), .ZN(n5444) );
  NAND2_X1 U6941 ( .A1(n5444), .A2(n5443), .ZN(n5445) );
  MUX2_X1 U6942 ( .A(n6868), .B(n6865), .S(n7824), .Z(n5450) );
  INV_X1 U6943 ( .A(SI_20_), .ZN(n9643) );
  NAND2_X1 U6944 ( .A1(n5450), .A2(n9643), .ZN(n5471) );
  INV_X1 U6945 ( .A(n5450), .ZN(n5451) );
  NAND2_X1 U6946 ( .A1(n5451), .A2(SI_20_), .ZN(n5452) );
  XNOR2_X1 U6947 ( .A(n5470), .B(n5469), .ZN(n6864) );
  NAND2_X1 U6948 ( .A1(n6864), .A2(n8840), .ZN(n5454) );
  OR2_X1 U6949 ( .A1(n5057), .A2(n6865), .ZN(n5453) );
  INV_X1 U6950 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8690) );
  NAND2_X1 U6951 ( .A1(n5455), .A2(n8690), .ZN(n5456) );
  NAND2_X1 U6952 ( .A1(n5475), .A2(n5456), .ZN(n9296) );
  OR2_X1 U6953 ( .A1(n9296), .A2(n4313), .ZN(n5461) );
  NAND2_X1 U6954 ( .A1(n8830), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U6955 ( .A1(n5478), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5457) );
  AND2_X1 U6956 ( .A1(n5458), .A2(n5457), .ZN(n5460) );
  NAND2_X1 U6957 ( .A1(n5477), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5459) );
  OAI22_X1 U6958 ( .A1(n9299), .A2(n4952), .B1(n9284), .B2(n5605), .ZN(n5462)
         );
  XNOR2_X1 U6959 ( .A(n5462), .B(n6950), .ZN(n5465) );
  OR2_X1 U6960 ( .A1(n9299), .A2(n5605), .ZN(n5464) );
  INV_X1 U6961 ( .A(n9284), .ZN(n9323) );
  NAND2_X1 U6962 ( .A1(n9323), .A2(n5606), .ZN(n5463) );
  NAND2_X1 U6963 ( .A1(n5464), .A2(n5463), .ZN(n5466) );
  NAND2_X1 U6964 ( .A1(n5465), .A2(n5466), .ZN(n8687) );
  INV_X1 U6965 ( .A(n5465), .ZN(n5468) );
  INV_X1 U6966 ( .A(n5466), .ZN(n5467) );
  NAND2_X1 U6967 ( .A1(n5468), .A2(n5467), .ZN(n8688) );
  MUX2_X1 U6968 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7824), .Z(n5492) );
  XNOR2_X1 U6969 ( .A(n5492), .B(n9646), .ZN(n5491) );
  XNOR2_X1 U6970 ( .A(n5494), .B(n5491), .ZN(n6869) );
  NAND2_X1 U6971 ( .A1(n6869), .A2(n8840), .ZN(n5473) );
  INV_X1 U6972 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6870) );
  OR2_X1 U6973 ( .A1(n5057), .A2(n6870), .ZN(n5472) );
  NAND2_X1 U6974 ( .A1(n9454), .A2(n8620), .ZN(n5483) );
  INV_X1 U6975 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U6976 ( .A1(n5475), .A2(n5474), .ZN(n5476) );
  AND2_X1 U6977 ( .A1(n5502), .A2(n5476), .ZN(n9287) );
  NAND2_X1 U6978 ( .A1(n9287), .A2(n5623), .ZN(n5481) );
  AOI22_X1 U6979 ( .A1(n8830), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n5477), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U6980 ( .A1(n5478), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5479) );
  INV_X1 U6981 ( .A(n9306), .ZN(n9015) );
  NAND2_X1 U6982 ( .A1(n9015), .A2(n5215), .ZN(n5482) );
  NAND2_X1 U6983 ( .A1(n5483), .A2(n5482), .ZN(n5484) );
  XNOR2_X1 U6984 ( .A(n5484), .B(n6950), .ZN(n5486) );
  NOR2_X1 U6985 ( .A1(n9306), .A2(n8625), .ZN(n5485) );
  AOI21_X1 U6986 ( .B1(n9454), .B2(n5634), .A(n5485), .ZN(n5487) );
  XNOR2_X1 U6987 ( .A(n5486), .B(n5487), .ZN(n8647) );
  INV_X1 U6988 ( .A(n5486), .ZN(n5488) );
  NAND2_X1 U6989 ( .A1(n5488), .A2(n5487), .ZN(n5489) );
  INV_X1 U6990 ( .A(n5491), .ZN(n5493) );
  MUX2_X1 U6991 ( .A(n7038), .B(n7035), .S(n7824), .Z(n5495) );
  NAND2_X1 U6992 ( .A1(n5495), .A2(n9580), .ZN(n5515) );
  INV_X1 U6993 ( .A(n5495), .ZN(n5496) );
  NAND2_X1 U6994 ( .A1(n5496), .A2(SI_22_), .ZN(n5497) );
  NAND2_X1 U6995 ( .A1(n5515), .A2(n5497), .ZN(n5516) );
  XNOR2_X1 U6996 ( .A(n5517), .B(n5516), .ZN(n7034) );
  NAND2_X1 U6997 ( .A1(n7034), .A2(n8840), .ZN(n5499) );
  OR2_X1 U6998 ( .A1(n5057), .A2(n7035), .ZN(n5498) );
  INV_X1 U6999 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U7000 ( .A1(n5502), .A2(n5501), .ZN(n5503) );
  NAND2_X1 U7001 ( .A1(n5526), .A2(n5503), .ZN(n9268) );
  OR2_X1 U7002 ( .A1(n9268), .A2(n5012), .ZN(n5509) );
  INV_X1 U7003 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U7004 ( .A1(n8830), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U7005 ( .A1(n5477), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5504) );
  OAI211_X1 U7006 ( .C1(n5506), .C2(n5685), .A(n5505), .B(n5504), .ZN(n5507)
         );
  INV_X1 U7007 ( .A(n5507), .ZN(n5508) );
  AND2_X1 U7008 ( .A1(n5606), .A2(n9114), .ZN(n5510) );
  AOI21_X1 U7009 ( .B1(n9449), .B2(n5634), .A(n5510), .ZN(n5514) );
  NAND2_X1 U7010 ( .A1(n9449), .A2(n8620), .ZN(n5512) );
  NAND2_X1 U7011 ( .A1(n9114), .A2(n5215), .ZN(n5511) );
  NAND2_X1 U7012 ( .A1(n5512), .A2(n5511), .ZN(n5513) );
  XNOR2_X1 U7013 ( .A(n5513), .B(n5031), .ZN(n8697) );
  INV_X1 U7014 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5518) );
  MUX2_X1 U7015 ( .A(n5518), .B(n7210), .S(n7824), .Z(n5519) );
  INV_X1 U7016 ( .A(SI_23_), .ZN(n9591) );
  NAND2_X1 U7017 ( .A1(n5519), .A2(n9591), .ZN(n5540) );
  INV_X1 U7018 ( .A(n5519), .ZN(n5520) );
  NAND2_X1 U7019 ( .A1(n5520), .A2(SI_23_), .ZN(n5521) );
  NAND2_X1 U7020 ( .A1(n7207), .A2(n8840), .ZN(n5523) );
  OR2_X1 U7021 ( .A1(n5057), .A2(n7210), .ZN(n5522) );
  INV_X1 U7022 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U7023 ( .A1(n5526), .A2(n5525), .ZN(n5527) );
  NAND2_X1 U7024 ( .A1(n5545), .A2(n5527), .ZN(n9253) );
  OR2_X1 U7025 ( .A1(n9253), .A2(n5012), .ZN(n5533) );
  INV_X1 U7026 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U7027 ( .A1(n5477), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U7028 ( .A1(n8830), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5528) );
  OAI211_X1 U7029 ( .C1(n5530), .C2(n5685), .A(n5529), .B(n5528), .ZN(n5531)
         );
  INV_X1 U7030 ( .A(n5531), .ZN(n5532) );
  OAI22_X1 U7031 ( .A1(n9257), .A2(n4952), .B1(n9265), .B2(n5605), .ZN(n5534)
         );
  OR2_X1 U7032 ( .A1(n9257), .A2(n5605), .ZN(n5536) );
  NAND2_X1 U7033 ( .A1(n9116), .A2(n5606), .ZN(n5535) );
  AND2_X1 U7034 ( .A1(n5536), .A2(n5535), .ZN(n8600) );
  NAND2_X1 U7035 ( .A1(n8601), .A2(n8600), .ZN(n8679) );
  NAND2_X1 U7036 ( .A1(n5537), .A2(n4371), .ZN(n8678) );
  MUX2_X1 U7037 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n7824), .Z(n5565) );
  INV_X1 U7038 ( .A(SI_24_), .ZN(n5541) );
  XNOR2_X1 U7039 ( .A(n5565), .B(n5541), .ZN(n5564) );
  XNOR2_X1 U7040 ( .A(n5563), .B(n5564), .ZN(n7362) );
  NAND2_X1 U7041 ( .A1(n7362), .A2(n8840), .ZN(n5543) );
  INV_X1 U7042 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7363) );
  OR2_X1 U7043 ( .A1(n5057), .A2(n7363), .ZN(n5542) );
  INV_X1 U7044 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7045 ( .A1(n5545), .A2(n5544), .ZN(n5546) );
  AND2_X1 U7046 ( .A1(n5576), .A2(n5546), .ZN(n9240) );
  NAND2_X1 U7047 ( .A1(n9240), .A2(n5623), .ZN(n5552) );
  INV_X1 U7048 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U7049 ( .A1(n8830), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U7050 ( .A1(n5477), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5547) );
  OAI211_X1 U7051 ( .C1(n5549), .C2(n5685), .A(n5548), .B(n5547), .ZN(n5550)
         );
  INV_X1 U7052 ( .A(n5550), .ZN(n5551) );
  OAI22_X1 U7053 ( .A1(n9243), .A2(n4952), .B1(n9250), .B2(n5605), .ZN(n5553)
         );
  XNOR2_X1 U7054 ( .A(n5553), .B(n5031), .ZN(n5556) );
  OR2_X1 U7055 ( .A1(n9243), .A2(n5605), .ZN(n5555) );
  NAND2_X1 U7056 ( .A1(n9120), .A2(n5606), .ZN(n5554) );
  NAND2_X1 U7057 ( .A1(n5556), .A2(n5557), .ZN(n5561) );
  INV_X1 U7058 ( .A(n5556), .ZN(n5559) );
  INV_X1 U7059 ( .A(n5557), .ZN(n5558) );
  NAND2_X1 U7060 ( .A1(n5559), .A2(n5558), .ZN(n5560) );
  NAND2_X1 U7061 ( .A1(n5561), .A2(n5560), .ZN(n8677) );
  INV_X1 U7062 ( .A(n5561), .ZN(n5562) );
  NAND2_X1 U7063 ( .A1(n5565), .A2(SI_24_), .ZN(n5566) );
  INV_X1 U7064 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n5568) );
  MUX2_X1 U7065 ( .A(n5568), .B(n7431), .S(n7824), .Z(n5569) );
  INV_X1 U7066 ( .A(SI_25_), .ZN(n9663) );
  NAND2_X1 U7067 ( .A1(n5569), .A2(n9663), .ZN(n5587) );
  INV_X1 U7068 ( .A(n5569), .ZN(n5570) );
  NAND2_X1 U7069 ( .A1(n5570), .A2(SI_25_), .ZN(n5571) );
  NAND2_X1 U7070 ( .A1(n5587), .A2(n5571), .ZN(n5588) );
  XNOR2_X1 U7071 ( .A(n5589), .B(n5588), .ZN(n7383) );
  NAND2_X1 U7072 ( .A1(n7383), .A2(n8840), .ZN(n5573) );
  OR2_X1 U7073 ( .A1(n5057), .A2(n7431), .ZN(n5572) );
  NAND2_X1 U7074 ( .A1(n9434), .A2(n8620), .ZN(n5585) );
  INV_X1 U7075 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U7076 ( .A1(n5576), .A2(n5575), .ZN(n5577) );
  NAND2_X1 U7077 ( .A1(n5596), .A2(n5577), .ZN(n9226) );
  INV_X1 U7078 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U7079 ( .A1(n5477), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U7080 ( .A1(n8830), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5578) );
  OAI211_X1 U7081 ( .C1(n5580), .C2(n5685), .A(n5579), .B(n5578), .ZN(n5581)
         );
  INV_X1 U7082 ( .A(n5581), .ZN(n5582) );
  INV_X1 U7083 ( .A(n9238), .ZN(n9014) );
  NAND2_X1 U7084 ( .A1(n9014), .A2(n5215), .ZN(n5584) );
  NAND2_X1 U7085 ( .A1(n5585), .A2(n5584), .ZN(n5586) );
  XNOR2_X1 U7086 ( .A(n5586), .B(n6950), .ZN(n5610) );
  INV_X1 U7087 ( .A(n9434), .ZN(n9230) );
  OAI22_X1 U7088 ( .A1(n9230), .A2(n5605), .B1(n9238), .B2(n8625), .ZN(n5609)
         );
  XNOR2_X1 U7089 ( .A(n5610), .B(n5609), .ZN(n8653) );
  INV_X1 U7090 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5590) );
  INV_X1 U7091 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7531) );
  MUX2_X1 U7092 ( .A(n5590), .B(n7531), .S(n7824), .Z(n5591) );
  INV_X1 U7093 ( .A(SI_26_), .ZN(n9593) );
  NAND2_X1 U7094 ( .A1(n5591), .A2(n9593), .ZN(n5615) );
  INV_X1 U7095 ( .A(n5591), .ZN(n5592) );
  NAND2_X1 U7096 ( .A1(n5592), .A2(SI_26_), .ZN(n5593) );
  NAND2_X1 U7097 ( .A1(n7510), .A2(n8840), .ZN(n5595) );
  OR2_X1 U7098 ( .A1(n5057), .A2(n7531), .ZN(n5594) );
  INV_X1 U7099 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8719) );
  NAND2_X1 U7100 ( .A1(n5596), .A2(n8719), .ZN(n5597) );
  NAND2_X1 U7101 ( .A1(n9213), .A2(n5623), .ZN(n5603) );
  INV_X1 U7102 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7103 ( .A1(n5477), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U7104 ( .A1(n8830), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5598) );
  OAI211_X1 U7105 ( .C1(n5600), .C2(n5685), .A(n5599), .B(n5598), .ZN(n5601)
         );
  INV_X1 U7106 ( .A(n5601), .ZN(n5602) );
  OAI22_X1 U7107 ( .A1(n9216), .A2(n4952), .B1(n9224), .B2(n5605), .ZN(n5604)
         );
  XNOR2_X1 U7108 ( .A(n5604), .B(n6950), .ZN(n5612) );
  OR2_X1 U7109 ( .A1(n9216), .A2(n5605), .ZN(n5608) );
  NAND2_X1 U7110 ( .A1(n9125), .A2(n5606), .ZN(n5607) );
  NAND2_X1 U7111 ( .A1(n5608), .A2(n5607), .ZN(n5611) );
  XNOR2_X1 U7112 ( .A(n5612), .B(n5611), .ZN(n8713) );
  NOR2_X1 U7113 ( .A1(n5610), .A2(n5609), .ZN(n8714) );
  INV_X1 U7114 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5617) );
  INV_X1 U7115 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7546) );
  MUX2_X1 U7116 ( .A(n5617), .B(n7546), .S(n7824), .Z(n5618) );
  INV_X1 U7117 ( .A(SI_27_), .ZN(n9645) );
  NAND2_X1 U7118 ( .A1(n5618), .A2(n9645), .ZN(n6078) );
  INV_X1 U7119 ( .A(n5618), .ZN(n5619) );
  NAND2_X1 U7120 ( .A1(n5619), .A2(SI_27_), .ZN(n5620) );
  NAND2_X1 U7121 ( .A1(n7543), .A2(n8840), .ZN(n5622) );
  OR2_X1 U7122 ( .A1(n5057), .A2(n7546), .ZN(n5621) );
  NAND2_X1 U7123 ( .A1(n9422), .A2(n8620), .ZN(n5631) );
  XNOR2_X1 U7124 ( .A(n5679), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9198) );
  NAND2_X1 U7125 ( .A1(n9198), .A2(n5623), .ZN(n5629) );
  INV_X1 U7126 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U7127 ( .A1(n8830), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7128 ( .A1(n5477), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5624) );
  OAI211_X1 U7129 ( .C1(n5685), .C2(n5626), .A(n5625), .B(n5624), .ZN(n5627)
         );
  INV_X1 U7130 ( .A(n5627), .ZN(n5628) );
  INV_X1 U7131 ( .A(n9210), .ZN(n9013) );
  NAND2_X1 U7132 ( .A1(n9013), .A2(n5215), .ZN(n5630) );
  NAND2_X1 U7133 ( .A1(n5631), .A2(n5630), .ZN(n5632) );
  XNOR2_X1 U7134 ( .A(n5632), .B(n5031), .ZN(n5636) );
  NOR2_X1 U7135 ( .A1(n9210), .A2(n8625), .ZN(n5633) );
  AOI21_X1 U7136 ( .B1(n9422), .B2(n5634), .A(n5633), .ZN(n5635) );
  NAND2_X1 U7137 ( .A1(n5636), .A2(n5635), .ZN(n8638) );
  OAI21_X1 U7138 ( .B1(n5636), .B2(n5635), .A(n8638), .ZN(n5638) );
  INV_X1 U7139 ( .A(n5637), .ZN(n5640) );
  INV_X1 U7140 ( .A(n5638), .ZN(n5639) );
  AOI21_X1 U7141 ( .B1(n8718), .B2(n5640), .A(n5639), .ZN(n5665) );
  INV_X1 U7142 ( .A(n5643), .ZN(n7429) );
  NAND3_X1 U7143 ( .A1(n7429), .A2(P1_B_REG_SCAN_IN), .A3(n7364), .ZN(n5642)
         );
  OAI22_X1 U7144 ( .A1(n9504), .A2(P1_D_REG_1__SCAN_IN), .B1(n5646), .B2(n5643), .ZN(n6944) );
  INV_X1 U7145 ( .A(n6944), .ZN(n6264) );
  INV_X1 U7146 ( .A(n9504), .ZN(n5645) );
  INV_X1 U7147 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U7148 ( .A1(n5645), .A2(n5644), .ZN(n5647) );
  INV_X1 U7149 ( .A(n5646), .ZN(n7532) );
  NAND2_X1 U7150 ( .A1(n7532), .A2(n7364), .ZN(n9506) );
  NOR4_X1 U7151 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5656) );
  NOR4_X1 U7152 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5655) );
  OR4_X1 U7153 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5653) );
  NOR4_X1 U7154 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5651) );
  NOR4_X1 U7155 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5650) );
  NOR4_X1 U7156 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5649) );
  NOR4_X1 U7157 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5648) );
  NAND4_X1 U7158 ( .A1(n5651), .A2(n5650), .A3(n5649), .A4(n5648), .ZN(n5652)
         );
  NOR4_X1 U7159 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5653), .A4(n5652), .ZN(n5654) );
  AND3_X1 U7160 ( .A1(n5656), .A2(n5655), .A3(n5654), .ZN(n5657) );
  NOR2_X1 U7161 ( .A1(n9504), .A2(n5657), .ZN(n6408) );
  INV_X1 U7162 ( .A(n6408), .ZN(n5658) );
  NAND3_X1 U7163 ( .A1(n6264), .A2(n6945), .A3(n5658), .ZN(n5669) );
  NAND2_X1 U7164 ( .A1(n4388), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5659) );
  XNOR2_X1 U7165 ( .A(n5659), .B(n4901), .ZN(n6201) );
  AND2_X1 U7166 ( .A1(n6201), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5660) );
  INV_X1 U7167 ( .A(n9505), .ZN(n5661) );
  OR2_X1 U7168 ( .A1(n5669), .A2(n5661), .ZN(n5675) );
  NAND2_X1 U7169 ( .A1(n5662), .A2(n5663), .ZN(n6412) );
  INV_X1 U7170 ( .A(n6412), .ZN(n8890) );
  NOR2_X1 U7171 ( .A1(n5675), .A2(n8890), .ZN(n5664) );
  INV_X1 U7172 ( .A(n7017), .ZN(n6413) );
  OAI21_X1 U7173 ( .B1(n8645), .B2(n5665), .A(n8717), .ZN(n5696) );
  AND2_X1 U7174 ( .A1(n5669), .A2(n9505), .ZN(n5666) );
  NOR2_X1 U7175 ( .A1(n7017), .A2(n6866), .ZN(n6967) );
  NAND2_X1 U7176 ( .A1(n5666), .A2(n6967), .ZN(n6364) );
  OR2_X1 U7177 ( .A1(n6412), .A2(n9005), .ZN(n5668) );
  NAND2_X1 U7178 ( .A1(n5668), .A2(n9505), .ZN(n6409) );
  NOR2_X1 U7179 ( .A1(n9961), .A2(n6409), .ZN(n5667) );
  AND3_X1 U7180 ( .A1(n5668), .A2(n4934), .A3(n6201), .ZN(n5671) );
  INV_X1 U7181 ( .A(n5669), .ZN(n5670) );
  OR2_X1 U7182 ( .A1(n9935), .A2(n5670), .ZN(n6362) );
  NAND2_X1 U7183 ( .A1(n5671), .A2(n6362), .ZN(n5672) );
  NAND2_X1 U7184 ( .A1(n5672), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5673) );
  OR2_X1 U7185 ( .A1(n6497), .A2(n5674), .ZN(n6951) );
  NOR2_X1 U7186 ( .A1(n5675), .A2(n6951), .ZN(n5690) );
  INV_X1 U7187 ( .A(n4312), .ZN(n6507) );
  NAND2_X1 U7188 ( .A1(n5690), .A2(n6507), .ZN(n8732) );
  INV_X1 U7189 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5678) );
  OAI22_X1 U7190 ( .A1(n9224), .A2(n8732), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5678), .ZN(n5692) );
  INV_X1 U7191 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5677) );
  OAI21_X1 U7192 ( .B1(n5679), .B2(n5678), .A(n5677), .ZN(n5682) );
  INV_X1 U7193 ( .A(n5679), .ZN(n5681) );
  AND2_X1 U7194 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5680) );
  NAND2_X1 U7195 ( .A1(n5681), .A2(n5680), .ZN(n9162) );
  NAND2_X1 U7196 ( .A1(n5682), .A2(n9162), .ZN(n8629) );
  INV_X1 U7197 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U7198 ( .A1(n8830), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U7199 ( .A1(n5477), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5683) );
  OAI211_X1 U7200 ( .C1(n5686), .C2(n5685), .A(n5684), .B(n5683), .ZN(n5687)
         );
  INV_X1 U7201 ( .A(n5687), .ZN(n5688) );
  NAND2_X1 U7202 ( .A1(n5690), .A2(n4312), .ZN(n8720) );
  NOR2_X1 U7203 ( .A1(n9192), .A2(n8720), .ZN(n5691) );
  AOI211_X1 U7204 ( .C1(n9198), .C2(n8723), .A(n5692), .B(n5691), .ZN(n5693)
         );
  INV_X1 U7205 ( .A(n5694), .ZN(n5695) );
  NAND2_X1 U7206 ( .A1(n5696), .A2(n5695), .ZN(P1_U3212) );
  NAND2_X1 U7207 ( .A1(n5851), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5866) );
  INV_X1 U7208 ( .A(n5866), .ZN(n5697) );
  NAND2_X1 U7209 ( .A1(n5697), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5881) );
  INV_X1 U7210 ( .A(n5925), .ZN(n5699) );
  AND2_X1 U7211 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n5698) );
  NAND2_X1 U7212 ( .A1(n5699), .A2(n5698), .ZN(n5927) );
  INV_X1 U7213 ( .A(n5927), .ZN(n5700) );
  NAND2_X1 U7214 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n5701) );
  INV_X1 U7215 ( .A(n5957), .ZN(n5702) );
  NAND2_X1 U7216 ( .A1(n5702), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5971) );
  INV_X1 U7217 ( .A(n5985), .ZN(n5703) );
  NAND2_X1 U7218 ( .A1(n5703), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5997) );
  INV_X1 U7219 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5996) );
  INV_X1 U7220 ( .A(n6007), .ZN(n5704) );
  NAND2_X1 U7221 ( .A1(n5704), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6018) );
  INV_X1 U7222 ( .A(n6018), .ZN(n5705) );
  NAND2_X1 U7223 ( .A1(n5705), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6028) );
  INV_X1 U7224 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9606) );
  INV_X1 U7225 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7712) );
  NAND2_X1 U7226 ( .A1(n6030), .A2(n7712), .ZN(n5706) );
  AND2_X1 U7227 ( .A1(n6040), .A2(n5706), .ZN(n8267) );
  NOR2_X1 U7228 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5712) );
  NOR2_X1 U7229 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5711) );
  NOR2_X1 U7230 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5710) );
  NAND4_X1 U7231 ( .A1(n5713), .A2(n5712), .A3(n5711), .A4(n5710), .ZN(n5718)
         );
  NOR2_X1 U7232 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5717) );
  NOR2_X1 U7233 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5716) );
  NOR2_X1 U7234 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5715) );
  NOR2_X1 U7235 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5714) );
  NAND4_X1 U7236 ( .A1(n5717), .A2(n5716), .A3(n5715), .A4(n5714), .ZN(n5950)
         );
  OR2_X2 U7237 ( .A1(n5718), .A2(n5950), .ZN(n5719) );
  INV_X1 U7238 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5721) );
  INV_X1 U7239 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5723) );
  XNOR2_X2 U7240 ( .A(n5724), .B(n5723), .ZN(n5730) );
  INV_X2 U7241 ( .A(n5730), .ZN(n8591) );
  NOR2_X1 U7242 ( .A1(n5725), .A2(n5726), .ZN(n5729) );
  AND2_X4 U7243 ( .A1(n8591), .A2(n8595), .ZN(n5815) );
  NAND2_X1 U7244 ( .A1(n8267), .A2(n5815), .ZN(n5736) );
  NAND2_X1 U7245 ( .A1(n6104), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5732) );
  NAND2_X1 U7246 ( .A1(n6182), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5731) );
  AND2_X1 U7247 ( .A1(n5732), .A2(n5731), .ZN(n5735) );
  INV_X2 U7248 ( .A(n5801), .ZN(n5778) );
  NAND2_X1 U7249 ( .A1(n5778), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5734) );
  NAND2_X1 U7250 ( .A1(n5742), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U7251 ( .A1(n4311), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5741) );
  NAND2_X1 U7252 ( .A1(n7207), .A2(n7828), .ZN(n5745) );
  INV_X2 U7253 ( .A(n5877), .ZN(n7812) );
  NAND2_X1 U7254 ( .A1(n7812), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5744) );
  INV_X1 U7255 ( .A(n8484), .ZN(n8269) );
  NAND2_X1 U7256 ( .A1(n6347), .A2(n7828), .ZN(n5753) );
  NOR2_X1 U7257 ( .A1(n5746), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5889) );
  INV_X1 U7258 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U7259 ( .A1(n5889), .A2(n5890), .ZN(n5904) );
  OAI21_X1 U7260 ( .B1(n5920), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5760) );
  INV_X1 U7261 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5747) );
  NAND2_X1 U7262 ( .A1(n5760), .A2(n5747), .ZN(n5748) );
  NAND2_X1 U7263 ( .A1(n5748), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5750) );
  INV_X1 U7264 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5749) );
  NAND2_X1 U7265 ( .A1(n5750), .A2(n5749), .ZN(n5935) );
  OR2_X1 U7266 ( .A1(n5750), .A2(n5749), .ZN(n5751) );
  AOI22_X1 U7267 ( .A1(n7812), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5993), .B2(
        n7419), .ZN(n5752) );
  INV_X2 U7268 ( .A(n6107), .ZN(n6182) );
  NAND2_X1 U7269 ( .A1(n6182), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5759) );
  XNOR2_X1 U7270 ( .A(n5941), .B(P2_REG3_REG_14__SCAN_IN), .ZN(n8405) );
  NAND2_X1 U7271 ( .A1(n5815), .A2(n8405), .ZN(n5758) );
  INV_X1 U7272 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n5754) );
  OR2_X1 U7273 ( .A1(n5800), .A2(n5754), .ZN(n5757) );
  INV_X1 U7274 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5755) );
  OR2_X1 U7275 ( .A1(n5801), .A2(n5755), .ZN(n5756) );
  NAND2_X1 U7276 ( .A1(n8538), .A2(n8431), .ZN(n7935) );
  NAND2_X1 U7277 ( .A1(n6304), .A2(n7828), .ZN(n5762) );
  XNOR2_X1 U7278 ( .A(n5760), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7004) );
  AOI22_X1 U7279 ( .A1(n7812), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5993), .B2(
        n7004), .ZN(n5761) );
  NAND2_X1 U7280 ( .A1(n6182), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5767) );
  INV_X1 U7281 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9633) );
  NAND2_X1 U7282 ( .A1(n5927), .A2(n9633), .ZN(n5763) );
  AND2_X1 U7283 ( .A1(n5941), .A2(n5763), .ZN(n8439) );
  NAND2_X1 U7284 ( .A1(n5815), .A2(n8439), .ZN(n5766) );
  INV_X1 U7285 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8583) );
  OR2_X1 U7286 ( .A1(n5800), .A2(n8583), .ZN(n5765) );
  INV_X1 U7287 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8442) );
  OR2_X1 U7288 ( .A1(n5801), .A2(n8442), .ZN(n5764) );
  INV_X1 U7289 ( .A(n8414), .ZN(n8039) );
  NAND2_X1 U7290 ( .A1(n8449), .A2(n8039), .ZN(n8400) );
  INV_X1 U7291 ( .A(n8400), .ZN(n5768) );
  INV_X1 U7292 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6619) );
  NAND2_X1 U7293 ( .A1(n5779), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5771) );
  NAND2_X1 U7294 ( .A1(n5798), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U7295 ( .A1(n5815), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5769) );
  NAND4_X1 U7296 ( .A1(n5772), .A2(n5771), .A3(n5770), .A4(n5769), .ZN(n5777)
         );
  INV_X1 U7297 ( .A(n5777), .ZN(n5789) );
  NAND2_X1 U7298 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5773) );
  XNOR2_X1 U7299 ( .A(n5773), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6618) );
  INV_X1 U7300 ( .A(n6618), .ZN(n5774) );
  NAND2_X1 U7301 ( .A1(n5789), .A2(n7217), .ZN(n7865) );
  NAND2_X1 U7302 ( .A1(n6673), .A2(n6496), .ZN(n6158) );
  NAND2_X1 U7303 ( .A1(n7865), .A2(n6158), .ZN(n6434) );
  NAND2_X1 U7304 ( .A1(n5778), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5784) );
  NAND2_X1 U7305 ( .A1(n5798), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5781) );
  NAND2_X1 U7306 ( .A1(n5815), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5780) );
  NOR2_X1 U7307 ( .A1(n4875), .A2(n5782), .ZN(n5783) );
  NAND2_X1 U7308 ( .A1(n5784), .A2(n5783), .ZN(n7183) );
  INV_X1 U7309 ( .A(SI_0_), .ZN(n5786) );
  INV_X1 U7310 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5785) );
  OAI21_X1 U7311 ( .B1(n7824), .B2(n5786), .A(n5785), .ZN(n5787) );
  AND2_X1 U7312 ( .A1(n5788), .A2(n5787), .ZN(n8599) );
  MUX2_X1 U7313 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8599), .S(n6603), .Z(n10001)
         );
  NAND2_X1 U7314 ( .A1(n6434), .A2(n6435), .ZN(n6436) );
  NAND2_X1 U7315 ( .A1(n5789), .A2(n6496), .ZN(n5790) );
  NAND2_X1 U7316 ( .A1(n5798), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7317 ( .A1(n5815), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5793) );
  INV_X1 U7318 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6620) );
  OR2_X1 U7319 ( .A1(n5801), .A2(n6620), .ZN(n5792) );
  NAND2_X1 U7320 ( .A1(n5821), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5797) );
  NAND2_X1 U7321 ( .A1(n5993), .A2(n6635), .ZN(n5796) );
  NAND2_X1 U7322 ( .A1(n6772), .A2(n7157), .ZN(n7872) );
  NAND2_X1 U7323 ( .A1(n7869), .A2(n7872), .ZN(n7839) );
  NAND2_X1 U7324 ( .A1(n6772), .A2(n10009), .ZN(n6766) );
  NAND2_X1 U7325 ( .A1(n5798), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5805) );
  INV_X1 U7326 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6752) );
  NAND2_X1 U7327 ( .A1(n5815), .A2(n6752), .ZN(n5804) );
  INV_X1 U7328 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5799) );
  OR2_X1 U7329 ( .A1(n5800), .A2(n5799), .ZN(n5803) );
  INV_X1 U7330 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6637) );
  NAND2_X1 U7331 ( .A1(n5821), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U7332 ( .A1(n5807), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5808) );
  MUX2_X1 U7333 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5808), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5809) );
  AND2_X1 U7334 ( .A1(n5806), .A2(n5809), .ZN(n6636) );
  NAND2_X1 U7335 ( .A1(n5993), .A2(n6636), .ZN(n5810) );
  INV_X1 U7336 ( .A(n6777), .ZN(n7086) );
  NAND2_X1 U7337 ( .A1(n7165), .A2(n7086), .ZN(n5812) );
  AND2_X1 U7338 ( .A1(n6766), .A2(n5812), .ZN(n5814) );
  INV_X1 U7339 ( .A(n5812), .ZN(n5813) );
  NAND2_X1 U7340 ( .A1(n6674), .A2(n7086), .ZN(n7888) );
  NAND2_X1 U7341 ( .A1(n7888), .A2(n7882), .ZN(n6160) );
  AOI21_X1 U7342 ( .B1(n7158), .B2(n5814), .A(n4876), .ZN(n7177) );
  NAND2_X1 U7343 ( .A1(n6182), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5820) );
  XNOR2_X1 U7344 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7170) );
  INV_X1 U7345 ( .A(n7170), .ZN(n6763) );
  NAND2_X1 U7346 ( .A1(n5815), .A2(n6763), .ZN(n5819) );
  INV_X1 U7347 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5816) );
  OR2_X1 U7348 ( .A1(n5800), .A2(n5816), .ZN(n5818) );
  INV_X1 U7349 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6639) );
  OR2_X1 U7350 ( .A1(n5801), .A2(n6639), .ZN(n5817) );
  INV_X1 U7351 ( .A(n6771), .ZN(n8047) );
  NAND2_X1 U7352 ( .A1(n5821), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U7353 ( .A1(n5806), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5822) );
  XNOR2_X1 U7354 ( .A(n5822), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6650) );
  NAND2_X1 U7355 ( .A1(n5993), .A2(n6650), .ZN(n5823) );
  OAI211_X1 U7356 ( .C1(n5864), .C2(n6252), .A(n5824), .B(n5823), .ZN(n7176)
         );
  NAND2_X1 U7357 ( .A1(n6771), .A2(n7176), .ZN(n7881) );
  NAND2_X1 U7358 ( .A1(n7177), .A2(n7840), .ZN(n7178) );
  NAND2_X1 U7359 ( .A1(n6771), .A2(n10014), .ZN(n5825) );
  NAND2_X1 U7360 ( .A1(n7178), .A2(n5825), .ZN(n7270) );
  NAND2_X1 U7361 ( .A1(n6182), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5832) );
  AOI21_X1 U7362 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5826) );
  NOR2_X1 U7363 ( .A1(n5826), .A2(n5841), .ZN(n7274) );
  NAND2_X1 U7364 ( .A1(n5815), .A2(n7274), .ZN(n5831) );
  INV_X1 U7365 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5827) );
  OR2_X1 U7366 ( .A1(n5800), .A2(n5827), .ZN(n5830) );
  INV_X1 U7367 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5828) );
  OR2_X1 U7368 ( .A1(n5801), .A2(n5828), .ZN(n5829) );
  NAND2_X1 U7369 ( .A1(n7812), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5839) );
  NOR2_X1 U7370 ( .A1(n5833), .A2(n8588), .ZN(n5834) );
  MUX2_X1 U7371 ( .A(n8588), .B(n5834), .S(P2_IR_REG_5__SCAN_IN), .Z(n5837) );
  OR2_X1 U7372 ( .A1(n5837), .A2(n5836), .ZN(n6643) );
  NAND2_X1 U7373 ( .A1(n5993), .A2(n6683), .ZN(n5838) );
  OAI211_X1 U7374 ( .C1(n5864), .C2(n6255), .A(n5839), .B(n5838), .ZN(n7275)
         );
  NAND2_X1 U7375 ( .A1(n7166), .A2(n7275), .ZN(n7883) );
  INV_X1 U7376 ( .A(n7166), .ZN(n8046) );
  INV_X1 U7377 ( .A(n7275), .ZN(n10019) );
  NAND2_X1 U7378 ( .A1(n7883), .A2(n7890), .ZN(n7838) );
  NAND2_X1 U7379 ( .A1(n7166), .A2(n10019), .ZN(n5840) );
  NAND2_X1 U7380 ( .A1(n6182), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5846) );
  INV_X1 U7381 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7025) );
  OR2_X1 U7382 ( .A1(n5801), .A2(n7025), .ZN(n5845) );
  NOR2_X1 U7383 ( .A1(n5841), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5842) );
  NOR2_X1 U7384 ( .A1(n5851), .A2(n5842), .ZN(n7028) );
  NAND2_X1 U7385 ( .A1(n5815), .A2(n7028), .ZN(n5844) );
  NAND2_X1 U7386 ( .A1(n6104), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5843) );
  NAND4_X1 U7387 ( .A1(n5846), .A2(n5845), .A3(n5844), .A4(n5843), .ZN(n8045)
         );
  NAND2_X1 U7388 ( .A1(n7812), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5849) );
  OR2_X1 U7389 ( .A1(n5836), .A2(n8588), .ZN(n5847) );
  XNOR2_X1 U7390 ( .A(n5847), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6701) );
  NAND2_X1 U7391 ( .A1(n5993), .A2(n6701), .ZN(n5848) );
  OAI211_X1 U7392 ( .C1(n5864), .C2(n6258), .A(n5849), .B(n5848), .ZN(n10024)
         );
  NOR2_X1 U7393 ( .A1(n8045), .A2(n10024), .ZN(n5850) );
  NAND2_X1 U7394 ( .A1(n6182), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5859) );
  INV_X1 U7395 ( .A(n5851), .ZN(n5853) );
  INV_X1 U7396 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U7397 ( .A1(n5853), .A2(n5852), .ZN(n5854) );
  NAND2_X1 U7398 ( .A1(n5866), .A2(n5854), .ZN(n6990) );
  INV_X1 U7399 ( .A(n6990), .ZN(n6861) );
  NAND2_X1 U7400 ( .A1(n5815), .A2(n6861), .ZN(n5858) );
  INV_X1 U7401 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6704) );
  OR2_X1 U7402 ( .A1(n5801), .A2(n6704), .ZN(n5857) );
  INV_X1 U7403 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5855) );
  OR2_X1 U7404 ( .A1(n5800), .A2(n5855), .ZN(n5856) );
  NAND2_X1 U7405 ( .A1(n7812), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U7406 ( .A1(n5860), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5861) );
  XNOR2_X1 U7407 ( .A(n5861), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6732) );
  NAND2_X1 U7408 ( .A1(n5993), .A2(n6732), .ZN(n5862) );
  NAND2_X1 U7409 ( .A1(n6914), .A2(n6937), .ZN(n7898) );
  INV_X1 U7410 ( .A(n6914), .ZN(n8044) );
  INV_X1 U7411 ( .A(n6937), .ZN(n6991) );
  NAND2_X1 U7412 ( .A1(n8044), .A2(n6991), .ZN(n7899) );
  NAND2_X1 U7413 ( .A1(n6914), .A2(n6991), .ZN(n5865) );
  NAND2_X1 U7414 ( .A1(n6182), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5873) );
  INV_X1 U7415 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9659) );
  NAND2_X1 U7416 ( .A1(n5866), .A2(n9659), .ZN(n5867) );
  AND2_X1 U7417 ( .A1(n5881), .A2(n5867), .ZN(n7262) );
  NAND2_X1 U7418 ( .A1(n5815), .A2(n7262), .ZN(n5872) );
  INV_X1 U7419 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n5868) );
  OR2_X1 U7420 ( .A1(n5801), .A2(n5868), .ZN(n5871) );
  INV_X1 U7421 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5869) );
  OR2_X1 U7422 ( .A1(n5800), .A2(n5869), .ZN(n5870) );
  NAND2_X1 U7423 ( .A1(n7828), .A2(n6267), .ZN(n5876) );
  NAND2_X1 U7424 ( .A1(n5746), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5874) );
  XNOR2_X1 U7425 ( .A(n5874), .B(P2_IR_REG_8__SCAN_IN), .ZN(n8054) );
  NAND2_X1 U7426 ( .A1(n5993), .A2(n8054), .ZN(n5875) );
  OAI211_X1 U7427 ( .C1(n5877), .C2(n6269), .A(n5876), .B(n5875), .ZN(n7263)
         );
  NAND2_X1 U7428 ( .A1(n7313), .A2(n7263), .ZN(n7905) );
  INV_X1 U7429 ( .A(n7263), .ZN(n10032) );
  NAND2_X1 U7430 ( .A1(n8043), .A2(n10032), .ZN(n7904) );
  NAND2_X1 U7431 ( .A1(n8043), .A2(n7263), .ZN(n5879) );
  NAND2_X1 U7432 ( .A1(n6182), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U7433 ( .A1(n5881), .A2(n5880), .ZN(n5882) );
  AND2_X1 U7434 ( .A1(n5897), .A2(n5882), .ZN(n7318) );
  NAND2_X1 U7435 ( .A1(n5815), .A2(n7318), .ZN(n5887) );
  INV_X1 U7436 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5883) );
  OR2_X1 U7437 ( .A1(n5800), .A2(n5883), .ZN(n5886) );
  INV_X1 U7438 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5884) );
  OR2_X1 U7439 ( .A1(n5801), .A2(n5884), .ZN(n5885) );
  NAND2_X1 U7440 ( .A1(n6273), .A2(n7828), .ZN(n5894) );
  OR2_X1 U7441 ( .A1(n5889), .A2(n8588), .ZN(n5891) );
  MUX2_X1 U7442 ( .A(n5891), .B(P2_IR_REG_31__SCAN_IN), .S(n5890), .Z(n5892)
         );
  AND2_X1 U7443 ( .A1(n5892), .A2(n5904), .ZN(n8068) );
  AOI22_X1 U7444 ( .A1(n7812), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5993), .B2(
        n8068), .ZN(n5893) );
  NAND2_X1 U7445 ( .A1(n7349), .A2(n8559), .ZN(n7907) );
  INV_X1 U7446 ( .A(n8559), .ZN(n7320) );
  INV_X1 U7447 ( .A(n7349), .ZN(n8042) );
  NAND2_X1 U7448 ( .A1(n7320), .A2(n8042), .ZN(n7915) );
  NAND2_X1 U7449 ( .A1(n7349), .A2(n7320), .ZN(n5896) );
  NAND2_X1 U7450 ( .A1(n6182), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U7451 ( .A1(n5897), .A2(n9604), .ZN(n5898) );
  AND2_X1 U7452 ( .A1(n5925), .A2(n5898), .ZN(n7399) );
  NAND2_X1 U7453 ( .A1(n5815), .A2(n7399), .ZN(n5902) );
  INV_X1 U7454 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5899) );
  OR2_X1 U7455 ( .A1(n5800), .A2(n5899), .ZN(n5901) );
  INV_X1 U7456 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7354) );
  OR2_X1 U7457 ( .A1(n5801), .A2(n7354), .ZN(n5900) );
  NAND2_X1 U7458 ( .A1(n5904), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5905) );
  XNOR2_X1 U7459 ( .A(n5905), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8081) );
  AOI22_X1 U7460 ( .A1(n7812), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5993), .B2(
        n8081), .ZN(n5906) );
  NAND2_X1 U7461 ( .A1(n7386), .A2(n7387), .ZN(n7914) );
  NAND2_X1 U7462 ( .A1(n7916), .A2(n7914), .ZN(n7347) );
  NAND2_X1 U7463 ( .A1(n7386), .A2(n4587), .ZN(n5907) );
  NAND2_X1 U7464 ( .A1(n6282), .A2(n7828), .ZN(n5911) );
  NAND2_X1 U7465 ( .A1(n5908), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5909) );
  XNOR2_X1 U7466 ( .A(n5909), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6829) );
  AOI22_X1 U7467 ( .A1(n7812), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5993), .B2(
        n6829), .ZN(n5910) );
  NAND2_X1 U7468 ( .A1(n5911), .A2(n5910), .ZN(n8555) );
  NAND2_X1 U7469 ( .A1(n6182), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5917) );
  XNOR2_X1 U7470 ( .A(n5925), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n7411) );
  NAND2_X1 U7471 ( .A1(n5815), .A2(n7411), .ZN(n5916) );
  INV_X1 U7472 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5912) );
  OR2_X1 U7473 ( .A1(n5800), .A2(n5912), .ZN(n5915) );
  INV_X1 U7474 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5913) );
  OR2_X1 U7475 ( .A1(n5801), .A2(n5913), .ZN(n5914) );
  OR2_X1 U7476 ( .A1(n8555), .A2(n7467), .ZN(n7924) );
  NAND2_X1 U7477 ( .A1(n8555), .A2(n7467), .ZN(n7925) );
  NAND2_X1 U7478 ( .A1(n7924), .A2(n7925), .ZN(n7301) );
  NAND2_X1 U7479 ( .A1(n7300), .A2(n7301), .ZN(n5919) );
  NAND2_X1 U7480 ( .A1(n8555), .A2(n8041), .ZN(n5918) );
  NAND2_X1 U7481 ( .A1(n6286), .A2(n7828), .ZN(n5923) );
  NAND2_X1 U7482 ( .A1(n5920), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5921) );
  XNOR2_X1 U7483 ( .A(n5921), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6901) );
  AOI22_X1 U7484 ( .A1(n7812), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5993), .B2(
        n6901), .ZN(n5922) );
  NAND2_X1 U7485 ( .A1(n6182), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5932) );
  INV_X1 U7486 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7407) );
  INV_X1 U7487 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5924) );
  OAI21_X1 U7488 ( .B1(n5925), .B2(n7407), .A(n5924), .ZN(n5926) );
  AND2_X1 U7489 ( .A1(n5927), .A2(n5926), .ZN(n7493) );
  NAND2_X1 U7490 ( .A1(n5815), .A2(n7493), .ZN(n5931) );
  INV_X1 U7491 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7463) );
  OR2_X1 U7492 ( .A1(n5801), .A2(n7463), .ZN(n5930) );
  INV_X1 U7493 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5928) );
  OR2_X1 U7494 ( .A1(n5800), .A2(n5928), .ZN(n5929) );
  OR2_X1 U7495 ( .A1(n10046), .A2(n8432), .ZN(n7928) );
  NAND2_X1 U7496 ( .A1(n10046), .A2(n8432), .ZN(n7926) );
  OR2_X1 U7497 ( .A1(n8449), .A2(n8414), .ZN(n7929) );
  NAND2_X1 U7498 ( .A1(n8449), .A2(n8414), .ZN(n7930) );
  INV_X1 U7499 ( .A(n8431), .ZN(n8038) );
  OR2_X1 U7500 ( .A1(n8538), .A2(n8038), .ZN(n5933) );
  NAND2_X1 U7501 ( .A1(n5934), .A2(n5933), .ZN(n8384) );
  NAND2_X1 U7502 ( .A1(n6370), .A2(n7828), .ZN(n5938) );
  NAND2_X1 U7503 ( .A1(n5935), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5936) );
  XNOR2_X1 U7504 ( .A(n5936), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8100) );
  AOI22_X1 U7505 ( .A1(n8100), .A2(n5993), .B1(n7812), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U7506 ( .A1(n6182), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5948) );
  INV_X1 U7507 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5940) );
  INV_X1 U7508 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5939) );
  OAI21_X1 U7509 ( .B1(n5941), .B2(n5940), .A(n5939), .ZN(n5942) );
  AND2_X1 U7510 ( .A1(n5942), .A2(n5957), .ZN(n8387) );
  NAND2_X1 U7511 ( .A1(n5815), .A2(n8387), .ZN(n5947) );
  INV_X1 U7512 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n5943) );
  OR2_X1 U7513 ( .A1(n5801), .A2(n5943), .ZN(n5946) );
  INV_X1 U7514 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n5944) );
  OR2_X1 U7515 ( .A1(n5800), .A2(n5944), .ZN(n5945) );
  NAND2_X1 U7516 ( .A1(n8533), .A2(n8413), .ZN(n7939) );
  NAND2_X1 U7517 ( .A1(n7940), .A2(n7939), .ZN(n8391) );
  NAND2_X1 U7518 ( .A1(n8384), .A2(n8391), .ZN(n8383) );
  INV_X1 U7519 ( .A(n8413), .ZN(n8037) );
  OR2_X1 U7520 ( .A1(n8533), .A2(n8037), .ZN(n5949) );
  NAND2_X1 U7521 ( .A1(n6419), .A2(n7828), .ZN(n5956) );
  OR2_X1 U7522 ( .A1(n5951), .A2(n8588), .ZN(n5953) );
  MUX2_X1 U7523 ( .A(n5953), .B(P2_IR_REG_31__SCAN_IN), .S(n5952), .Z(n5954)
         );
  AND2_X1 U7524 ( .A1(n5964), .A2(n5954), .ZN(n8116) );
  AOI22_X1 U7525 ( .A1(n7812), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5993), .B2(
        n8116), .ZN(n5955) );
  NAND2_X1 U7526 ( .A1(n6182), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5962) );
  INV_X1 U7527 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9582) );
  NAND2_X1 U7528 ( .A1(n5957), .A2(n9582), .ZN(n5958) );
  AND2_X1 U7529 ( .A1(n5971), .A2(n5958), .ZN(n8374) );
  NAND2_X1 U7530 ( .A1(n5815), .A2(n8374), .ZN(n5961) );
  INV_X1 U7531 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8579) );
  OR2_X1 U7532 ( .A1(n5800), .A2(n8579), .ZN(n5960) );
  INV_X1 U7533 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8376) );
  OR2_X1 U7534 ( .A1(n5801), .A2(n8376), .ZN(n5959) );
  OR2_X1 U7535 ( .A1(n8524), .A2(n8393), .ZN(n7945) );
  NAND2_X1 U7536 ( .A1(n8524), .A2(n8393), .ZN(n7944) );
  NAND2_X1 U7537 ( .A1(n7945), .A2(n7944), .ZN(n8367) );
  INV_X1 U7538 ( .A(n8393), .ZN(n8036) );
  NAND2_X1 U7539 ( .A1(n8524), .A2(n8036), .ZN(n5963) );
  NAND2_X1 U7540 ( .A1(n6450), .A2(n7828), .ZN(n5970) );
  NAND2_X1 U7541 ( .A1(n5964), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5967) );
  MUX2_X1 U7542 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5967), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5968) );
  AND2_X1 U7543 ( .A1(n5992), .A2(n5968), .ZN(n8128) );
  AOI22_X1 U7544 ( .A1(n7812), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5993), .B2(
        n8128), .ZN(n5969) );
  NAND2_X1 U7545 ( .A1(n6182), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U7546 ( .A1(n5971), .A2(n9661), .ZN(n5972) );
  AND2_X1 U7547 ( .A1(n5985), .A2(n5972), .ZN(n8359) );
  NAND2_X1 U7548 ( .A1(n5815), .A2(n8359), .ZN(n5976) );
  INV_X1 U7549 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8111) );
  OR2_X1 U7550 ( .A1(n5801), .A2(n8111), .ZN(n5975) );
  INV_X1 U7551 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n5973) );
  OR2_X1 U7552 ( .A1(n5800), .A2(n5973), .ZN(n5974) );
  NAND2_X1 U7553 ( .A1(n8521), .A2(n8369), .ZN(n7948) );
  INV_X1 U7554 ( .A(n8369), .ZN(n8342) );
  OR2_X1 U7555 ( .A1(n8521), .A2(n8342), .ZN(n5979) );
  NAND2_X1 U7556 ( .A1(n6594), .A2(n7828), .ZN(n5982) );
  NAND2_X1 U7557 ( .A1(n5992), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5980) );
  XNOR2_X1 U7558 ( .A(n5980), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8145) );
  AOI22_X1 U7559 ( .A1(n7812), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5993), .B2(
        n8145), .ZN(n5981) );
  NAND2_X1 U7560 ( .A1(n6104), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5990) );
  INV_X1 U7561 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5983) );
  OR2_X1 U7562 ( .A1(n5801), .A2(n5983), .ZN(n5989) );
  NAND2_X1 U7563 ( .A1(n6182), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5988) );
  INV_X1 U7564 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7565 ( .A1(n5985), .A2(n5984), .ZN(n5986) );
  AND2_X1 U7566 ( .A1(n5997), .A2(n5986), .ZN(n8335) );
  NAND2_X1 U7567 ( .A1(n5815), .A2(n8335), .ZN(n5987) );
  NAND4_X1 U7568 ( .A1(n5990), .A2(n5989), .A3(n5988), .A4(n5987), .ZN(n8327)
         );
  NAND2_X1 U7569 ( .A1(n8514), .A2(n8327), .ZN(n5991) );
  NAND2_X1 U7570 ( .A1(n6744), .A2(n7828), .ZN(n5995) );
  AOI22_X1 U7571 ( .A1(n7812), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8152), .B2(
        n5993), .ZN(n5994) );
  NAND2_X1 U7572 ( .A1(n6182), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U7573 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  AND2_X1 U7574 ( .A1(n6007), .A2(n5998), .ZN(n8321) );
  NAND2_X1 U7575 ( .A1(n5815), .A2(n8321), .ZN(n6003) );
  INV_X1 U7576 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n5999) );
  OR2_X1 U7577 ( .A1(n5800), .A2(n5999), .ZN(n6002) );
  INV_X1 U7578 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6000) );
  OR2_X1 U7579 ( .A1(n5801), .A2(n6000), .ZN(n6001) );
  OR2_X1 U7580 ( .A1(n8510), .A2(n7785), .ZN(n7958) );
  NAND2_X1 U7581 ( .A1(n8510), .A2(n7785), .ZN(n8309) );
  NAND2_X1 U7582 ( .A1(n7958), .A2(n8309), .ZN(n8317) );
  NAND2_X1 U7583 ( .A1(n6864), .A2(n7828), .ZN(n6006) );
  NAND2_X1 U7584 ( .A1(n7812), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U7585 ( .A1(n6182), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6014) );
  INV_X1 U7586 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9642) );
  NAND2_X1 U7587 ( .A1(n6007), .A2(n9642), .ZN(n6008) );
  AND2_X1 U7588 ( .A1(n6018), .A2(n6008), .ZN(n8307) );
  NAND2_X1 U7589 ( .A1(n5815), .A2(n8307), .ZN(n6013) );
  INV_X1 U7590 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n6009) );
  OR2_X1 U7591 ( .A1(n5801), .A2(n6009), .ZN(n6012) );
  INV_X1 U7592 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n6010) );
  OR2_X1 U7593 ( .A1(n5800), .A2(n6010), .ZN(n6011) );
  NAND2_X1 U7594 ( .A1(n8504), .A2(n7729), .ZN(n7959) );
  NAND2_X1 U7595 ( .A1(n7966), .A2(n7959), .ZN(n8303) );
  NAND2_X1 U7596 ( .A1(n8504), .A2(n4560), .ZN(n6015) );
  NAND2_X1 U7597 ( .A1(n8302), .A2(n6015), .ZN(n8290) );
  NAND2_X1 U7598 ( .A1(n6869), .A2(n7828), .ZN(n6017) );
  NAND2_X1 U7599 ( .A1(n7812), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7600 ( .A1(n6104), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7601 ( .A1(n6182), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6022) );
  INV_X1 U7602 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9648) );
  NAND2_X1 U7603 ( .A1(n6018), .A2(n9648), .ZN(n6019) );
  AND2_X1 U7604 ( .A1(n6028), .A2(n6019), .ZN(n8293) );
  NAND2_X1 U7605 ( .A1(n5815), .A2(n8293), .ZN(n6021) );
  NAND2_X1 U7606 ( .A1(n5778), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6020) );
  NAND4_X1 U7607 ( .A1(n6023), .A2(n6022), .A3(n6021), .A4(n6020), .ZN(n8311)
         );
  OR2_X1 U7608 ( .A1(n8499), .A2(n8311), .ZN(n6024) );
  NAND2_X1 U7609 ( .A1(n8499), .A2(n8311), .ZN(n6025) );
  NAND2_X1 U7610 ( .A1(n7034), .A2(n7828), .ZN(n6027) );
  NAND2_X1 U7611 ( .A1(n7812), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U7612 ( .A1(n6182), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6035) );
  INV_X1 U7613 ( .A(n5815), .ZN(n6087) );
  NAND2_X1 U7614 ( .A1(n6028), .A2(n9606), .ZN(n6029) );
  NAND2_X1 U7615 ( .A1(n6030), .A2(n6029), .ZN(n8274) );
  OR2_X1 U7616 ( .A1(n6087), .A2(n8274), .ZN(n6034) );
  INV_X1 U7617 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n6031) );
  OR2_X1 U7618 ( .A1(n5800), .A2(n6031), .ZN(n6033) );
  INV_X1 U7619 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8275) );
  OR2_X1 U7620 ( .A1(n5801), .A2(n8275), .ZN(n6032) );
  NAND2_X1 U7621 ( .A1(n8493), .A2(n8257), .ZN(n7960) );
  INV_X1 U7622 ( .A(n8279), .ZN(n6036) );
  INV_X1 U7623 ( .A(n8257), .ZN(n8297) );
  OR2_X1 U7624 ( .A1(n8484), .A2(n8284), .ZN(n7973) );
  NAND2_X1 U7625 ( .A1(n8484), .A2(n8284), .ZN(n7976) );
  NAND2_X1 U7626 ( .A1(n7362), .A2(n7828), .ZN(n6038) );
  NAND2_X1 U7627 ( .A1(n7812), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6037) );
  INV_X1 U7628 ( .A(n6040), .ZN(n6039) );
  NAND2_X1 U7629 ( .A1(n6039), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6048) );
  INV_X1 U7630 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9673) );
  NAND2_X1 U7631 ( .A1(n6040), .A2(n9673), .ZN(n6041) );
  NAND2_X1 U7632 ( .A1(n6048), .A2(n6041), .ZN(n8238) );
  OR2_X1 U7633 ( .A1(n8238), .A2(n6087), .ZN(n6044) );
  AOI22_X1 U7634 ( .A1(n6104), .A2(P2_REG0_REG_24__SCAN_IN), .B1(n6182), .B2(
        P2_REG1_REG_24__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7635 ( .A1(n5778), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U7636 ( .A1(n8479), .A2(n8258), .ZN(n7978) );
  INV_X1 U7637 ( .A(n8258), .ZN(n8035) );
  OAI22_X1 U7638 ( .A1(n8235), .A2(n7974), .B1(n8035), .B2(n8479), .ZN(n8221)
         );
  NAND2_X1 U7639 ( .A1(n7383), .A2(n7828), .ZN(n6046) );
  NAND2_X1 U7640 ( .A1(n7812), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6045) );
  INV_X1 U7641 ( .A(n6048), .ZN(n6047) );
  NAND2_X1 U7642 ( .A1(n6047), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6060) );
  INV_X1 U7643 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U7644 ( .A1(n6048), .A2(n7738), .ZN(n6049) );
  NAND2_X1 U7645 ( .A1(n6060), .A2(n6049), .ZN(n8228) );
  OR2_X1 U7646 ( .A1(n8228), .A2(n6087), .ZN(n6055) );
  INV_X1 U7647 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7648 ( .A1(n5778), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7649 ( .A1(n6182), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6050) );
  OAI211_X1 U7650 ( .C1(n5800), .C2(n6052), .A(n6051), .B(n6050), .ZN(n6053)
         );
  INV_X1 U7651 ( .A(n6053), .ZN(n6054) );
  NAND2_X1 U7652 ( .A1(n8476), .A2(n8245), .ZN(n7981) );
  INV_X1 U7653 ( .A(n8245), .ZN(n8034) );
  NAND2_X1 U7654 ( .A1(n7510), .A2(n7828), .ZN(n6058) );
  NAND2_X1 U7655 ( .A1(n7812), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6057) );
  INV_X1 U7656 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7657 ( .A1(n6060), .A2(n6059), .ZN(n6061) );
  INV_X1 U7658 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7659 ( .A1(n5778), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7660 ( .A1(n6182), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6062) );
  OAI211_X1 U7661 ( .C1(n5800), .C2(n6064), .A(n6063), .B(n6062), .ZN(n6065)
         );
  OR2_X1 U7662 ( .A1(n8471), .A2(n8226), .ZN(n7984) );
  NAND2_X1 U7663 ( .A1(n8471), .A2(n8226), .ZN(n7985) );
  NAND2_X1 U7664 ( .A1(n7984), .A2(n7985), .ZN(n8208) );
  INV_X1 U7665 ( .A(n8226), .ZN(n8033) );
  NAND2_X1 U7666 ( .A1(n8217), .A2(n8226), .ZN(n6066) );
  NAND2_X1 U7667 ( .A1(n7543), .A2(n7828), .ZN(n6068) );
  NAND2_X1 U7668 ( .A1(n7812), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6067) );
  XNOR2_X1 U7669 ( .A(n6085), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8190) );
  NAND2_X1 U7670 ( .A1(n8190), .A2(n5815), .ZN(n6074) );
  INV_X1 U7671 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7672 ( .A1(n5778), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7673 ( .A1(n6182), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6069) );
  OAI211_X1 U7674 ( .C1(n5800), .C2(n6071), .A(n6070), .B(n6069), .ZN(n6072)
         );
  INV_X1 U7675 ( .A(n6072), .ZN(n6073) );
  XNOR2_X1 U7676 ( .A(n8464), .B(n8210), .ZN(n8194) );
  NAND2_X1 U7677 ( .A1(n8192), .A2(n8210), .ZN(n6075) );
  MUX2_X1 U7678 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7824), .Z(n6097) );
  INV_X1 U7679 ( .A(SI_28_), .ZN(n6098) );
  XNOR2_X1 U7680 ( .A(n6097), .B(n6098), .ZN(n6095) );
  NAND2_X1 U7681 ( .A1(n8616), .A2(n7828), .ZN(n6080) );
  NAND2_X1 U7682 ( .A1(n7812), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6079) );
  INV_X1 U7683 ( .A(n6085), .ZN(n6082) );
  AND2_X1 U7684 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6081) );
  NAND2_X1 U7685 ( .A1(n6082), .A2(n6081), .ZN(n6103) );
  INV_X1 U7686 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6084) );
  INV_X1 U7687 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6083) );
  OAI21_X1 U7688 ( .B1(n6085), .B2(n6084), .A(n6083), .ZN(n6086) );
  NAND2_X1 U7689 ( .A1(n6103), .A2(n6086), .ZN(n8174) );
  INV_X1 U7690 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7691 ( .A1(n5778), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7692 ( .A1(n5798), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6088) );
  OAI211_X1 U7693 ( .C1(n5800), .C2(n6090), .A(n6089), .B(n6088), .ZN(n6091)
         );
  INV_X1 U7694 ( .A(n6091), .ZN(n6092) );
  NAND2_X1 U7695 ( .A1(n8459), .A2(n8196), .ZN(n7998) );
  NAND2_X1 U7696 ( .A1(n7994), .A2(n7998), .ZN(n8178) );
  NAND2_X1 U7697 ( .A1(n8171), .A2(n8178), .ZN(n8170) );
  NAND2_X1 U7698 ( .A1(n8170), .A2(n6094), .ZN(n6111) );
  INV_X1 U7699 ( .A(n6097), .ZN(n6099) );
  MUX2_X1 U7700 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n7824), .Z(n7580) );
  INV_X1 U7701 ( .A(SI_29_), .ZN(n7582) );
  XNOR2_X1 U7702 ( .A(n7580), .B(n7582), .ZN(n6100) );
  NAND2_X1 U7703 ( .A1(n8841), .A2(n7828), .ZN(n6102) );
  NAND2_X1 U7704 ( .A1(n7812), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6101) );
  INV_X1 U7705 ( .A(n6103), .ZN(n6189) );
  INV_X1 U7706 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7707 ( .A1(n6104), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U7708 ( .A1(n5778), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6105) );
  OAI211_X1 U7709 ( .C1(n6108), .C2(n6107), .A(n6106), .B(n6105), .ZN(n6109)
         );
  AOI21_X1 U7710 ( .B1(n6189), .B2(n5815), .A(n6109), .ZN(n7672) );
  NAND2_X1 U7711 ( .A1(n8455), .A2(n7672), .ZN(n8005) );
  NAND2_X1 U7712 ( .A1(n6125), .A2(n4592), .ZN(n6113) );
  INV_X1 U7713 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U7714 ( .A1(n6118), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6119) );
  MUX2_X1 U7715 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6119), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6120) );
  NOR2_X1 U7716 ( .A1(n4384), .A2(n8588), .ZN(n6121) );
  MUX2_X1 U7717 ( .A(n8588), .B(n6121), .S(P2_IR_REG_25__SCAN_IN), .Z(n6122)
         );
  INV_X1 U7718 ( .A(n6122), .ZN(n6123) );
  AND2_X1 U7719 ( .A1(n6118), .A2(n6123), .ZN(n7384) );
  NAND2_X1 U7720 ( .A1(n8027), .A2(n8019), .ZN(n6598) );
  NAND2_X1 U7721 ( .A1(n6128), .A2(n6127), .ZN(n6129) );
  NAND2_X1 U7722 ( .A1(n6129), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6131) );
  OR2_X1 U7723 ( .A1(n6598), .A2(n8024), .ZN(n6132) );
  INV_X1 U7724 ( .A(n6471), .ZN(n6153) );
  AND2_X1 U7725 ( .A1(n7368), .A2(n6133), .ZN(n9996) );
  XNOR2_X1 U7726 ( .A(n7368), .B(P2_B_REG_SCAN_IN), .ZN(n6134) );
  NAND2_X1 U7727 ( .A1(n6135), .A2(n6134), .ZN(n6136) );
  INV_X1 U7728 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9995) );
  OR2_X1 U7729 ( .A1(n6139), .A2(n6138), .ZN(n6140) );
  NAND2_X1 U7730 ( .A1(n6141), .A2(n6140), .ZN(n6557) );
  INV_X1 U7731 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9998) );
  NOR2_X1 U7732 ( .A1(n7384), .A2(n7511), .ZN(n9999) );
  AOI21_X1 U7733 ( .B1(n9992), .B2(n9998), .A(n9999), .ZN(n6431) );
  NOR4_X1 U7734 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6145) );
  NOR4_X1 U7735 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6144) );
  NOR4_X1 U7736 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6143) );
  NOR4_X1 U7737 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6142) );
  NAND4_X1 U7738 ( .A1(n6145), .A2(n6144), .A3(n6143), .A4(n6142), .ZN(n6151)
         );
  NOR2_X1 U7739 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n6149) );
  NOR4_X1 U7740 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6148) );
  NOR4_X1 U7741 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6147) );
  NOR4_X1 U7742 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6146) );
  NAND4_X1 U7743 ( .A1(n6149), .A2(n6148), .A3(n6147), .A4(n6146), .ZN(n6150)
         );
  OAI21_X1 U7744 ( .B1(n6151), .B2(n6150), .A(n9992), .ZN(n6430) );
  AND2_X1 U7745 ( .A1(n6431), .A2(n6430), .ZN(n6464) );
  NAND2_X1 U7746 ( .A1(n10000), .A2(n6464), .ZN(n6152) );
  NAND2_X2 U7747 ( .A1(n6193), .A2(n8440), .ZN(n8438) );
  NAND2_X1 U7748 ( .A1(n8019), .A2(n8020), .ZN(n6480) );
  NAND2_X1 U7749 ( .A1(n7036), .A2(n6480), .ZN(n6155) );
  NAND3_X1 U7750 ( .A1(n6598), .A2(n6155), .A3(n7833), .ZN(n8427) );
  OR2_X1 U7751 ( .A1(n6480), .A2(n7833), .ZN(n7080) );
  NAND2_X1 U7752 ( .A1(n8427), .A2(n7080), .ZN(n6156) );
  INV_X1 U7753 ( .A(n7183), .ZN(n6157) );
  NAND2_X1 U7754 ( .A1(n6157), .A2(n10001), .ZN(n7184) );
  NAND3_X1 U7755 ( .A1(n6159), .A2(n7871), .A3(n6158), .ZN(n7149) );
  NAND2_X1 U7756 ( .A1(n7149), .A2(n7872), .ZN(n6770) );
  INV_X1 U7757 ( .A(n6160), .ZN(n7879) );
  NAND2_X1 U7758 ( .A1(n6770), .A2(n7879), .ZN(n6769) );
  INV_X1 U7759 ( .A(n7882), .ZN(n6161) );
  NOR2_X1 U7760 ( .A1(n7840), .A2(n6161), .ZN(n6162) );
  NAND2_X1 U7761 ( .A1(n6769), .A2(n6162), .ZN(n6163) );
  NAND2_X1 U7762 ( .A1(n6163), .A2(n7889), .ZN(n7278) );
  INV_X1 U7763 ( .A(n7890), .ZN(n6164) );
  INV_X1 U7764 ( .A(n8045), .ZN(n6858) );
  NAND2_X1 U7765 ( .A1(n6858), .A2(n10024), .ZN(n7897) );
  INV_X1 U7766 ( .A(n10024), .ZN(n7030) );
  NAND2_X1 U7767 ( .A1(n8045), .A2(n7030), .ZN(n7894) );
  NAND2_X1 U7768 ( .A1(n7023), .A2(n7843), .ZN(n6932) );
  INV_X1 U7769 ( .A(n7896), .ZN(n7847) );
  INV_X1 U7770 ( .A(n7897), .ZN(n6165) );
  NOR2_X1 U7771 ( .A1(n7847), .A2(n6165), .ZN(n6166) );
  NAND2_X1 U7772 ( .A1(n6167), .A2(n7849), .ZN(n7311) );
  INV_X1 U7773 ( .A(n7907), .ZN(n7909) );
  NOR2_X1 U7774 ( .A1(n7347), .A2(n7909), .ZN(n6168) );
  NAND2_X1 U7775 ( .A1(n7311), .A2(n6168), .ZN(n6169) );
  INV_X1 U7776 ( .A(n7924), .ZN(n6170) );
  INV_X1 U7777 ( .A(n7926), .ZN(n6171) );
  INV_X1 U7778 ( .A(n8423), .ZN(n8428) );
  OR2_X2 U7779 ( .A1(n8412), .A2(n8411), .ZN(n8416) );
  INV_X1 U7780 ( .A(n8391), .ZN(n7937) );
  INV_X1 U7781 ( .A(n7945), .ZN(n6172) );
  OR2_X1 U7782 ( .A1(n8353), .A2(n5978), .ZN(n6173) );
  INV_X1 U7783 ( .A(n8327), .ZN(n8355) );
  OR2_X1 U7784 ( .A1(n8514), .A2(n8355), .ZN(n7956) );
  NAND2_X1 U7785 ( .A1(n8514), .A2(n8355), .ZN(n7955) );
  NAND2_X1 U7786 ( .A1(n8340), .A2(n8339), .ZN(n8338) );
  NAND2_X1 U7787 ( .A1(n8338), .A2(n7955), .ZN(n8325) );
  INV_X1 U7788 ( .A(n8317), .ZN(n8326) );
  NAND2_X1 U7789 ( .A1(n8325), .A2(n8326), .ZN(n8324) );
  INV_X1 U7790 ( .A(n8309), .ZN(n6174) );
  NOR2_X1 U7791 ( .A1(n8303), .A2(n6174), .ZN(n6175) );
  INV_X1 U7792 ( .A(n8311), .ZN(n8283) );
  OR2_X1 U7793 ( .A1(n8499), .A2(n8283), .ZN(n7965) );
  NAND2_X1 U7794 ( .A1(n8499), .A2(n8283), .ZN(n8280) );
  NAND2_X1 U7795 ( .A1(n7965), .A2(n8280), .ZN(n8289) );
  INV_X1 U7796 ( .A(n8280), .ZN(n6176) );
  INV_X1 U7797 ( .A(n8261), .ZN(n7975) );
  INV_X1 U7798 ( .A(n8254), .ZN(n7968) );
  NOR2_X1 U7799 ( .A1(n7975), .A2(n7968), .ZN(n6177) );
  INV_X1 U7800 ( .A(n7976), .ZN(n8244) );
  INV_X1 U7801 ( .A(n6178), .ZN(n7979) );
  INV_X1 U7802 ( .A(n8194), .ZN(n7987) );
  INV_X1 U7803 ( .A(n8464), .ZN(n8192) );
  NAND2_X1 U7804 ( .A1(n8192), .A2(n8180), .ZN(n7992) );
  INV_X1 U7805 ( .A(n8178), .ZN(n7861) );
  INV_X1 U7806 ( .A(n7994), .ZN(n6179) );
  NAND2_X1 U7807 ( .A1(n6180), .A2(n6110), .ZN(n7820) );
  OAI21_X1 U7808 ( .B1(n6110), .B2(n6180), .A(n7820), .ZN(n6181) );
  NAND2_X1 U7809 ( .A1(n8019), .A2(n7841), .ZN(n7836) );
  INV_X1 U7810 ( .A(n6605), .ZN(n6616) );
  INV_X1 U7811 ( .A(n8341), .ZN(n6188) );
  INV_X1 U7812 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U7813 ( .A1(n6182), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7814 ( .A1(n5778), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6183) );
  OAI211_X1 U7815 ( .C1(n5800), .C2(n6185), .A(n6184), .B(n6183), .ZN(n8031)
         );
  INV_X1 U7816 ( .A(n8031), .ZN(n6187) );
  INV_X1 U7817 ( .A(n6609), .ZN(n8025) );
  AOI21_X1 U7818 ( .B1(n8025), .B2(P2_B_REG_SCAN_IN), .A(n8430), .ZN(n8160) );
  INV_X1 U7819 ( .A(n8160), .ZN(n6186) );
  NOR2_X1 U7820 ( .A1(n8457), .A2(n8406), .ZN(n6196) );
  INV_X1 U7821 ( .A(n8455), .ZN(n6191) );
  NOR2_X1 U7822 ( .A1(n6479), .A2(n8020), .ZN(n6467) );
  AOI22_X1 U7823 ( .A1(n8406), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n6189), .B2(
        n8404), .ZN(n6190) );
  OAI21_X1 U7824 ( .B1(n6191), .B2(n8408), .A(n6190), .ZN(n6195) );
  NAND2_X1 U7825 ( .A1(n7154), .A2(n10009), .ZN(n7153) );
  NAND2_X1 U7826 ( .A1(n7271), .A2(n7030), .ZN(n7027) );
  INV_X1 U7827 ( .A(n7386), .ZN(n10039) );
  INV_X1 U7828 ( .A(n8449), .ZN(n8544) );
  INV_X1 U7829 ( .A(n8538), .ZN(n8409) );
  NAND2_X1 U7830 ( .A1(n8445), .A2(n8409), .ZN(n8402) );
  INV_X1 U7831 ( .A(n8521), .ZN(n8362) );
  INV_X1 U7832 ( .A(n8514), .ZN(n8337) );
  INV_X1 U7833 ( .A(n8499), .ZN(n8295) );
  INV_X1 U7834 ( .A(n8493), .ZN(n8276) );
  INV_X1 U7835 ( .A(n8471), .ZN(n8217) );
  NAND2_X1 U7836 ( .A1(n8227), .A2(n8217), .ZN(n8211) );
  INV_X1 U7837 ( .A(n8173), .ZN(n6192) );
  AOI211_X1 U7838 ( .C1(n8455), .C2(n6192), .A(n10050), .B(n8165), .ZN(n8454)
         );
  AND2_X1 U7839 ( .A1(n8454), .A2(n7324), .ZN(n6194) );
  NAND2_X1 U7840 ( .A1(n6199), .A2(n6201), .ZN(n6232) );
  OR2_X2 U7841 ( .A1(n6232), .A2(P1_U3084), .ZN(n9027) );
  INV_X1 U7842 ( .A(n6599), .ZN(n6200) );
  NAND2_X2 U7843 ( .A1(n6200), .A2(n10000), .ZN(n8049) );
  INV_X1 U7844 ( .A(n6201), .ZN(n7208) );
  OR2_X1 U7845 ( .A1(n6412), .A2(n7208), .ZN(n6202) );
  NAND2_X1 U7846 ( .A1(n6216), .A2(n8837), .ZN(n6315) );
  NAND2_X1 U7847 ( .A1(n6315), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AND2_X1 U7848 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7227) );
  NOR2_X1 U7849 ( .A1(n9905), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6203) );
  AOI21_X1 U7850 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9905), .A(n6203), .ZN(
        n9897) );
  NOR2_X1 U7851 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6337), .ZN(n6204) );
  AOI21_X1 U7852 ( .B1(n6337), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6204), .ZN(
        n6335) );
  NOR2_X1 U7853 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9867), .ZN(n6205) );
  AOI21_X1 U7854 ( .B1(n9867), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6205), .ZN(
        n9876) );
  INV_X1 U7855 ( .A(n6248), .ZN(n6359) );
  INV_X1 U7856 ( .A(n6245), .ZN(n6380) );
  INV_X1 U7857 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6206) );
  MUX2_X1 U7858 ( .A(n6206), .B(P1_REG2_REG_2__SCAN_IN), .S(n6245), .Z(n6389)
         );
  INV_X1 U7859 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7072) );
  MUX2_X1 U7860 ( .A(n7072), .B(P1_REG2_REG_1__SCAN_IN), .S(n6242), .Z(n6329)
         );
  AND2_X1 U7861 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6374) );
  NAND2_X1 U7862 ( .A1(n6329), .A2(n6374), .ZN(n6328) );
  INV_X1 U7863 ( .A(n6242), .ZN(n6327) );
  NAND2_X1 U7864 ( .A1(n6327), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7865 ( .A1(n6328), .A2(n6207), .ZN(n6388) );
  XOR2_X1 U7866 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6248), .Z(n6356) );
  NOR2_X1 U7867 ( .A1(n9863), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6208) );
  AOI21_X1 U7868 ( .B1(n9863), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6208), .ZN(
        n9854) );
  NAND2_X1 U7869 ( .A1(n9855), .A2(n9854), .ZN(n9853) );
  OAI21_X1 U7870 ( .B1(n9863), .B2(P1_REG2_REG_4__SCAN_IN), .A(n9853), .ZN(
        n9877) );
  NAND2_X1 U7871 ( .A1(n9876), .A2(n9877), .ZN(n9875) );
  OAI21_X1 U7872 ( .B1(n9867), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9875), .ZN(
        n9888) );
  NAND2_X1 U7873 ( .A1(n9892), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6209) );
  OAI21_X1 U7874 ( .B1(n9892), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6209), .ZN(
        n9887) );
  NOR2_X1 U7875 ( .A1(n9888), .A2(n9887), .ZN(n9886) );
  OAI21_X1 U7876 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9905), .A(n9895), .ZN(
        n6214) );
  NAND2_X1 U7877 ( .A1(n6400), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6210) );
  OAI21_X1 U7878 ( .B1(n6400), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6210), .ZN(
        n6213) );
  NOR2_X1 U7879 ( .A1(n6213), .A2(n6214), .ZN(n6394) );
  NOR2_X1 U7880 ( .A1(n6211), .A2(P1_U3084), .ZN(n6212) );
  NAND2_X1 U7881 ( .A1(n6216), .A2(n6212), .ZN(n9087) );
  INV_X1 U7882 ( .A(n9087), .ZN(n6231) );
  AOI211_X1 U7883 ( .C1(n6214), .C2(n6213), .A(n6394), .B(n9885), .ZN(n6236)
         );
  INV_X1 U7884 ( .A(n6211), .ZN(n9094) );
  OR2_X1 U7885 ( .A1(n9094), .A2(n4312), .ZN(n6377) );
  NOR2_X1 U7886 ( .A1(n6377), .A2(P1_U3084), .ZN(n6215) );
  MUX2_X1 U7887 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n6217), .S(n6400), .Z(n6229)
         );
  NAND2_X1 U7888 ( .A1(n9905), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6218) );
  OAI21_X1 U7889 ( .B1(n9905), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6218), .ZN(
        n9900) );
  NOR2_X1 U7890 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6337), .ZN(n6219) );
  AOI21_X1 U7891 ( .B1(n6337), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6219), .ZN(
        n6340) );
  OR2_X1 U7892 ( .A1(n9867), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6221) );
  NAND2_X1 U7893 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9867), .ZN(n6220) );
  NAND2_X1 U7894 ( .A1(n6221), .A2(n6220), .ZN(n9869) );
  MUX2_X1 U7895 ( .A(n4973), .B(P1_REG1_REG_2__SCAN_IN), .S(n6245), .Z(n6383)
         );
  MUX2_X1 U7896 ( .A(n4954), .B(P1_REG1_REG_1__SCAN_IN), .S(n6242), .Z(n6323)
         );
  AND2_X1 U7897 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6322) );
  NAND2_X1 U7898 ( .A1(n6323), .A2(n6322), .ZN(n6321) );
  NAND2_X1 U7899 ( .A1(n6327), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6222) );
  NAND2_X1 U7900 ( .A1(n6321), .A2(n6222), .ZN(n6382) );
  NAND2_X1 U7901 ( .A1(n6383), .A2(n6382), .ZN(n6381) );
  NAND2_X1 U7902 ( .A1(n6380), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U7903 ( .A1(n6381), .A2(n6223), .ZN(n6352) );
  XNOR2_X1 U7904 ( .A(n6248), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n6353) );
  NAND2_X1 U7905 ( .A1(n6352), .A2(n6353), .ZN(n6351) );
  NAND2_X1 U7906 ( .A1(n6359), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6224) );
  AND2_X1 U7907 ( .A1(n6351), .A2(n6224), .ZN(n9857) );
  NOR2_X1 U7908 ( .A1(n9863), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6225) );
  AOI21_X1 U7909 ( .B1(n9863), .B2(P1_REG1_REG_4__SCAN_IN), .A(n6225), .ZN(
        n9858) );
  NAND2_X1 U7910 ( .A1(n9857), .A2(n9858), .ZN(n9856) );
  INV_X1 U7911 ( .A(n6225), .ZN(n6226) );
  NAND2_X1 U7912 ( .A1(n9856), .A2(n6226), .ZN(n9870) );
  NOR2_X1 U7913 ( .A1(n9869), .A2(n9870), .ZN(n9868) );
  AOI21_X1 U7914 ( .B1(n9867), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9868), .ZN(
        n9884) );
  NOR2_X1 U7915 ( .A1(n9892), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6227) );
  AOI21_X1 U7916 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n9892), .A(n6227), .ZN(
        n9883) );
  NAND2_X1 U7917 ( .A1(n9884), .A2(n9883), .ZN(n9882) );
  OAI21_X1 U7918 ( .B1(n9892), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9882), .ZN(
        n6339) );
  NAND2_X1 U7919 ( .A1(n6340), .A2(n6339), .ZN(n6338) );
  OAI21_X1 U7920 ( .B1(n6337), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6338), .ZN(
        n9901) );
  NOR2_X1 U7921 ( .A1(n9900), .A2(n9901), .ZN(n9899) );
  AOI21_X1 U7922 ( .B1(n9905), .B2(P1_REG1_REG_8__SCAN_IN), .A(n9899), .ZN(
        n6228) );
  NAND2_X1 U7923 ( .A1(n6228), .A2(n6229), .ZN(n6399) );
  OAI21_X1 U7924 ( .B1(n6229), .B2(n6228), .A(n6399), .ZN(n6230) );
  AND2_X1 U7925 ( .A1(n9920), .A2(n6230), .ZN(n6235) );
  INV_X1 U7926 ( .A(n9912), .ZN(n9057) );
  INV_X1 U7927 ( .A(n6400), .ZN(n6276) );
  INV_X1 U7928 ( .A(n6232), .ZN(n6233) );
  INV_X1 U7929 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10100) );
  OAI22_X1 U7930 ( .A1(n9057), .A2(n6276), .B1(n9925), .B2(n10100), .ZN(n6234)
         );
  OR4_X1 U7931 ( .A1(n7227), .A2(n6236), .A3(n6235), .A4(n6234), .ZN(P1_U3250)
         );
  XNOR2_X1 U7932 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OR2_X1 U7933 ( .A1(n7824), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7545) );
  AND2_X1 U7934 ( .A1(n7824), .A2(P2_U3152), .ZN(n8594) );
  AOI22_X1 U7935 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n8594), .B1(n6635), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6237) );
  OAI21_X1 U7936 ( .B1(n6246), .B2(n7545), .A(n6237), .ZN(P2_U3356) );
  INV_X1 U7937 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6238) );
  CLKBUF_X1 U7938 ( .A(n7545), .Z(n8597) );
  INV_X1 U7939 ( .A(n6636), .ZN(n6670) );
  OAI222_X1 U7940 ( .A1(n7365), .A2(n6238), .B1(n8597), .B2(n6249), .C1(n7694), 
        .C2(n6670), .ZN(P2_U3355) );
  INV_X1 U7941 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6239) );
  OAI222_X1 U7942 ( .A1(n7365), .A2(n6239), .B1(n8597), .B2(n6255), .C1(n7694), 
        .C2(n6643), .ZN(P2_U3353) );
  INV_X1 U7943 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6240) );
  OAI222_X1 U7944 ( .A1(n7365), .A2(n6240), .B1(n8597), .B2(n6243), .C1(n7694), 
        .C2(n5774), .ZN(P2_U3357) );
  INV_X1 U7945 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6241) );
  INV_X1 U7946 ( .A(n6650), .ZN(n6657) );
  OAI222_X1 U7947 ( .A1(n7365), .A2(n6241), .B1(n8597), .B2(n6252), .C1(n7694), 
        .C2(n6657), .ZN(P2_U3354) );
  OR2_X2 U7948 ( .A1(n7824), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7689) );
  INV_X1 U7949 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6244) );
  AND2_X1 U7950 ( .A1(n7824), .A2(P1_U3084), .ZN(n7206) );
  INV_X2 U7951 ( .A(n7206), .ZN(n9512) );
  OAI222_X1 U7952 ( .A1(n7689), .A2(n6244), .B1(n9512), .B2(n6243), .C1(
        P1_U3084), .C2(n6242), .ZN(P1_U3352) );
  OAI222_X1 U7953 ( .A1(n7689), .A2(n6247), .B1(n9512), .B2(n6246), .C1(
        P1_U3084), .C2(n6245), .ZN(P1_U3351) );
  OAI222_X1 U7954 ( .A1(n7689), .A2(n6250), .B1(n9512), .B2(n6249), .C1(
        P1_U3084), .C2(n6248), .ZN(P1_U3350) );
  OAI222_X1 U7955 ( .A1(n7689), .A2(n6253), .B1(n9512), .B2(n6252), .C1(
        P1_U3084), .C2(n6251), .ZN(P1_U3349) );
  OAI222_X1 U7956 ( .A1(n7689), .A2(n4428), .B1(n9512), .B2(n6255), .C1(
        P1_U3084), .C2(n6254), .ZN(P1_U3348) );
  INV_X1 U7957 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6256) );
  INV_X1 U7958 ( .A(n6701), .ZN(n6694) );
  OAI222_X1 U7959 ( .A1(n7365), .A2(n6256), .B1(n8597), .B2(n6258), .C1(n7694), 
        .C2(n6694), .ZN(P2_U3352) );
  OAI222_X1 U7960 ( .A1(n7689), .A2(n6259), .B1(n9512), .B2(n6258), .C1(
        P1_U3084), .C2(n6257), .ZN(P1_U3347) );
  INV_X1 U7961 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6260) );
  INV_X1 U7962 ( .A(n6732), .ZN(n6709) );
  INV_X1 U7963 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U7964 ( .A1(n6264), .A2(n9505), .ZN(n6265) );
  OAI21_X1 U7965 ( .B1(n9505), .B2(n6266), .A(n6265), .ZN(P1_U3441) );
  INV_X1 U7966 ( .A(n6267), .ZN(n6271) );
  INV_X1 U7967 ( .A(n8054), .ZN(n6268) );
  OAI222_X1 U7968 ( .A1(n7365), .A2(n6269), .B1(n8597), .B2(n6271), .C1(n7694), 
        .C2(n6268), .ZN(P2_U3350) );
  OAI222_X1 U7969 ( .A1(n7689), .A2(n6272), .B1(n9512), .B2(n6271), .C1(
        P1_U3084), .C2(n6270), .ZN(P1_U3345) );
  INV_X1 U7970 ( .A(n6273), .ZN(n6277) );
  AOI22_X1 U7971 ( .A1(n8068), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n8594), .ZN(n6274) );
  OAI21_X1 U7972 ( .B1(n6277), .B2(n8597), .A(n6274), .ZN(P2_U3349) );
  OAI222_X1 U7973 ( .A1(n9512), .A2(n6277), .B1(n6276), .B2(P1_U3084), .C1(
        n6275), .C2(n7689), .ZN(P1_U3344) );
  INV_X1 U7974 ( .A(n6278), .ZN(n6281) );
  AOI22_X1 U7975 ( .A1(n8081), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n8594), .ZN(n6279) );
  OAI21_X1 U7976 ( .B1(n6281), .B2(n8597), .A(n6279), .ZN(P2_U3348) );
  INV_X1 U7977 ( .A(n6574), .ZN(n6401) );
  OAI222_X1 U7978 ( .A1(n9512), .A2(n6281), .B1(n6401), .B2(P1_U3084), .C1(
        n6280), .C2(n7689), .ZN(P1_U3343) );
  INV_X1 U7979 ( .A(n6282), .ZN(n6285) );
  AOI22_X1 U7980 ( .A1(n6829), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n8594), .ZN(n6283) );
  OAI21_X1 U7981 ( .B1(n6285), .B2(n8597), .A(n6283), .ZN(P2_U3347) );
  INV_X1 U7982 ( .A(n6575), .ZN(n9037) );
  INV_X1 U7983 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6284) );
  OAI222_X1 U7984 ( .A1(n9512), .A2(n6285), .B1(n9037), .B2(P1_U3084), .C1(
        n6284), .C2(n7689), .ZN(P1_U3342) );
  INV_X1 U7985 ( .A(n6286), .ZN(n6294) );
  INV_X1 U7986 ( .A(n7689), .ZN(n9510) );
  AOI22_X1 U7987 ( .A1(n6847), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9510), .ZN(n6287) );
  OAI21_X1 U7988 ( .B1(n6294), .B2(n9512), .A(n6287), .ZN(P1_U3341) );
  INV_X1 U7989 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6293) );
  INV_X1 U7990 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U7991 ( .A1(n8830), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6290) );
  INV_X1 U7992 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6288) );
  OR2_X1 U7993 ( .A1(n5010), .A2(n6288), .ZN(n6289) );
  OAI211_X1 U7994 ( .C1(n5685), .C2(n6291), .A(n6290), .B(n6289), .ZN(n9096)
         );
  NAND2_X1 U7995 ( .A1(n9096), .A2(P1_U4006), .ZN(n6292) );
  OAI21_X1 U7996 ( .B1(P1_U4006), .B2(n6293), .A(n6292), .ZN(P1_U3586) );
  INV_X1 U7997 ( .A(n6901), .ZN(n6838) );
  OAI222_X1 U7998 ( .A1(n7365), .A2(n6295), .B1(n8597), .B2(n6294), .C1(
        P2_U3152), .C2(n6838), .ZN(P2_U3346) );
  NAND2_X1 U7999 ( .A1(n9994), .A2(n6490), .ZN(n6296) );
  NAND2_X1 U8000 ( .A1(n6296), .A2(n6603), .ZN(n6298) );
  OR2_X1 U8001 ( .A1(n6557), .A2(P2_U3152), .ZN(n8029) );
  INV_X1 U8002 ( .A(n8029), .ZN(n7144) );
  OR2_X1 U8003 ( .A1(n9994), .A2(n7144), .ZN(n6297) );
  NOR2_X1 U8004 ( .A1(n9987), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8005 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6303) );
  INV_X1 U8006 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U8007 ( .A1(n5798), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6300) );
  INV_X1 U8008 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8161) );
  OR2_X1 U8009 ( .A1(n5801), .A2(n8161), .ZN(n6299) );
  OAI211_X1 U8010 ( .C1(n5800), .C2(n6301), .A(n6300), .B(n6299), .ZN(n8159)
         );
  NAND2_X1 U8011 ( .A1(n8159), .A2(P2_U3966), .ZN(n6302) );
  OAI21_X1 U8012 ( .B1(n6303), .B2(P2_U3966), .A(n6302), .ZN(P2_U3583) );
  INV_X1 U8013 ( .A(n6304), .ZN(n6345) );
  AOI22_X1 U8014 ( .A1(n7199), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9510), .ZN(n6305) );
  OAI21_X1 U8015 ( .B1(n6345), .B2(n9512), .A(n6305), .ZN(P1_U3340) );
  INV_X1 U8016 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6307) );
  NAND2_X1 U8017 ( .A1(n7183), .A2(P2_U3966), .ZN(n6306) );
  OAI21_X1 U8018 ( .B1(n6307), .B2(P2_U3966), .A(n6306), .ZN(P2_U3552) );
  INV_X1 U8019 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6320) );
  OR2_X1 U8020 ( .A1(n4312), .A2(n4917), .ZN(n6308) );
  NAND2_X1 U8021 ( .A1(n6377), .A2(n6308), .ZN(n6312) );
  OR2_X1 U8022 ( .A1(n6312), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6375) );
  NAND2_X1 U8023 ( .A1(n6211), .A2(n6309), .ZN(n6310) );
  INV_X1 U8024 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6316) );
  NAND2_X1 U8025 ( .A1(n6310), .A2(n6316), .ZN(n6311) );
  NAND2_X1 U8026 ( .A1(n6312), .A2(n6311), .ZN(n6313) );
  NAND3_X1 U8027 ( .A1(n6375), .A2(P1_STATE_REG_SCAN_IN), .A3(n6313), .ZN(
        n6314) );
  NOR2_X1 U8028 ( .A1(n6315), .A2(n6314), .ZN(n6318) );
  INV_X1 U8029 ( .A(n9920), .ZN(n9898) );
  NOR3_X1 U8030 ( .A1(n9898), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n6316), .ZN(
        n6317) );
  AOI211_X1 U8031 ( .C1(P1_REG3_REG_0__SCAN_IN), .C2(P1_U3084), .A(n6318), .B(
        n6317), .ZN(n6319) );
  OAI21_X1 U8032 ( .B1(n9925), .B2(n6320), .A(n6319), .ZN(P1_U3241) );
  INV_X1 U8033 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6332) );
  OAI211_X1 U8034 ( .C1(n6323), .C2(n6322), .A(n9920), .B(n6321), .ZN(n6324)
         );
  OAI21_X1 U8035 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6325), .A(n6324), .ZN(n6326) );
  AOI21_X1 U8036 ( .B1(n6327), .B2(n9912), .A(n6326), .ZN(n6331) );
  OAI211_X1 U8037 ( .C1(n6329), .C2(n6374), .A(n9921), .B(n6328), .ZN(n6330)
         );
  OAI211_X1 U8038 ( .C1(n6332), .C2(n9925), .A(n6331), .B(n6330), .ZN(P1_U3242) );
  INV_X1 U8039 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6344) );
  OAI21_X1 U8040 ( .B1(n6335), .B2(n6334), .A(n6333), .ZN(n6336) );
  AOI22_X1 U8041 ( .A1(n6337), .A2(n9912), .B1(n9921), .B2(n6336), .ZN(n6343)
         );
  OAI21_X1 U8042 ( .B1(n6340), .B2(n6339), .A(n6338), .ZN(n6341) );
  AND2_X1 U8043 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6880) );
  AOI21_X1 U8044 ( .B1(n9920), .B2(n6341), .A(n6880), .ZN(n6342) );
  OAI211_X1 U8045 ( .C1(n9925), .C2(n6344), .A(n6343), .B(n6342), .ZN(P1_U3248) );
  INV_X1 U8046 ( .A(n7004), .ZN(n6999) );
  OAI222_X1 U8047 ( .A1(n7365), .A2(n6346), .B1(n8597), .B2(n6345), .C1(n6999), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8048 ( .A(n6347), .ZN(n6349) );
  INV_X1 U8049 ( .A(n7439), .ZN(n7432) );
  INV_X1 U8050 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6348) );
  OAI222_X1 U8051 ( .A1(n9512), .A2(n6349), .B1(n7432), .B2(P1_U3084), .C1(
        n6348), .C2(n7689), .ZN(P1_U3339) );
  INV_X1 U8052 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6350) );
  INV_X1 U8053 ( .A(n7419), .ZN(n7002) );
  OAI222_X1 U8054 ( .A1(n7365), .A2(n6350), .B1(n8597), .B2(n6349), .C1(n7002), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8055 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6361) );
  OAI211_X1 U8056 ( .C1(n6353), .C2(n6352), .A(n9920), .B(n6351), .ZN(n6354)
         );
  NAND2_X1 U8057 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U8058 ( .A1(n6354), .A2(n6536), .ZN(n6358) );
  AOI211_X1 U8059 ( .C1(n4330), .C2(n6356), .A(n6355), .B(n9885), .ZN(n6357)
         );
  AOI211_X1 U8060 ( .C1(n9912), .C2(n6359), .A(n6358), .B(n6357), .ZN(n6360)
         );
  OAI21_X1 U8061 ( .B1(n6361), .B2(n9925), .A(n6360), .ZN(P1_U3244) );
  INV_X1 U8062 ( .A(n7019), .ZN(n6509) );
  INV_X1 U8063 ( .A(n6409), .ZN(n6363) );
  NAND3_X1 U8064 ( .A1(n6364), .A2(n6363), .A3(n6362), .ZN(n6461) );
  AOI22_X1 U8065 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n6461), .B1(n8734), .B2(
        n6500), .ZN(n6369) );
  OAI21_X1 U8066 ( .B1(n6367), .B2(n6366), .A(n6365), .ZN(n6378) );
  NAND2_X1 U8067 ( .A1(n6378), .A2(n8717), .ZN(n6368) );
  OAI211_X1 U8068 ( .C1(n8726), .C2(n6509), .A(n6369), .B(n6368), .ZN(P1_U3230) );
  INV_X1 U8069 ( .A(n6370), .ZN(n6372) );
  OAI222_X1 U8070 ( .A1(n7689), .A2(n6371), .B1(n9512), .B2(n6372), .C1(
        P1_U3084), .C2(n9049), .ZN(P1_U3338) );
  INV_X1 U8071 ( .A(n8100), .ZN(n8090) );
  OAI222_X1 U8072 ( .A1(n7365), .A2(n6373), .B1(n7545), .B2(n6372), .C1(
        P2_U3152), .C2(n8090), .ZN(P2_U3343) );
  NOR2_X1 U8073 ( .A1(n4312), .A2(n6211), .ZN(n9007) );
  AOI21_X1 U8074 ( .B1(n9007), .B2(n6374), .A(n9027), .ZN(n6376) );
  OAI211_X1 U8075 ( .C1(n6378), .C2(n6377), .A(n6376), .B(n6375), .ZN(n6379)
         );
  INV_X1 U8076 ( .A(n6379), .ZN(n9861) );
  NAND2_X1 U8077 ( .A1(n9912), .A2(n6380), .ZN(n6385) );
  OAI211_X1 U8078 ( .C1(n6383), .C2(n6382), .A(n9920), .B(n6381), .ZN(n6384)
         );
  OAI211_X1 U8079 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9402), .A(n6385), .B(n6384), .ZN(n6386) );
  INV_X1 U8080 ( .A(n6386), .ZN(n6391) );
  OAI211_X1 U8081 ( .C1(n6389), .C2(n6388), .A(n9921), .B(n6387), .ZN(n6390)
         );
  OAI211_X1 U8082 ( .C1(n9520), .C2(n9925), .A(n6391), .B(n6390), .ZN(n6392)
         );
  OR2_X1 U8083 ( .A1(n9861), .A2(n6392), .ZN(P1_U3243) );
  INV_X1 U8084 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6407) );
  NOR2_X1 U8085 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6393), .ZN(n7373) );
  NAND2_X1 U8086 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n6574), .ZN(n6395) );
  OAI21_X1 U8087 ( .B1(n6574), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6395), .ZN(
        n6396) );
  NOR2_X1 U8088 ( .A1(n6397), .A2(n6396), .ZN(n6573) );
  AOI211_X1 U8089 ( .C1(n6397), .C2(n6396), .A(n6573), .B(n9885), .ZN(n6398)
         );
  AOI211_X1 U8090 ( .C1(n9912), .C2(n6574), .A(n7373), .B(n6398), .ZN(n6406)
         );
  OAI21_X1 U8091 ( .B1(n6400), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6399), .ZN(
        n6403) );
  AOI22_X1 U8092 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6574), .B1(n6401), .B2(
        n5188), .ZN(n6402) );
  NAND2_X1 U8093 ( .A1(n6402), .A2(n6403), .ZN(n6566) );
  OAI21_X1 U8094 ( .B1(n6403), .B2(n6402), .A(n6566), .ZN(n6404) );
  NAND2_X1 U8095 ( .A1(n6404), .A2(n9920), .ZN(n6405) );
  OAI211_X1 U8096 ( .C1(n9925), .C2(n6407), .A(n6406), .B(n6405), .ZN(P1_U3251) );
  OAI21_X1 U8097 ( .B1(n9824), .B2(n5663), .A(n6944), .ZN(n6410) );
  INV_X1 U8098 ( .A(n9796), .ZN(n9771) );
  AND2_X1 U8099 ( .A1(n6509), .A2(n9028), .ZN(n8965) );
  NOR2_X1 U8100 ( .A1(n6505), .A2(n8965), .ZN(n8871) );
  INV_X1 U8101 ( .A(n6951), .ZN(n9008) );
  NOR3_X1 U8102 ( .A1(n8871), .A2(n9008), .A3(n6413), .ZN(n6414) );
  AOI21_X1 U8103 ( .B1(n9771), .B2(n6500), .A(n6414), .ZN(n7013) );
  OAI21_X1 U8104 ( .B1(n6509), .B2(n7017), .A(n7013), .ZN(n6417) );
  NAND2_X1 U8105 ( .A1(n6417), .A2(n9971), .ZN(n6415) );
  OAI21_X1 U8106 ( .B1(n9971), .B2(n4921), .A(n6415), .ZN(P1_U3454) );
  NAND2_X1 U8107 ( .A1(n6417), .A2(n9980), .ZN(n6418) );
  OAI21_X1 U8108 ( .B1(n9980), .B2(n6309), .A(n6418), .ZN(P1_U3523) );
  INV_X1 U8109 ( .A(n6419), .ZN(n6454) );
  AOI22_X1 U8110 ( .A1(n8116), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8594), .ZN(n6420) );
  OAI21_X1 U8111 ( .B1(n6454), .B2(n8597), .A(n6420), .ZN(P2_U3342) );
  XNOR2_X1 U8112 ( .A(n6421), .B(n6422), .ZN(n6423) );
  XOR2_X1 U8113 ( .A(n6424), .B(n6423), .Z(n6429) );
  NOR2_X1 U8114 ( .A1(n8726), .A2(n8969), .ZN(n6427) );
  INV_X1 U8115 ( .A(n9026), .ZN(n7046) );
  INV_X1 U8116 ( .A(n9028), .ZN(n6425) );
  OAI22_X1 U8117 ( .A1(n7046), .A2(n8720), .B1(n8732), .B2(n6425), .ZN(n6426)
         );
  AOI211_X1 U8118 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n6461), .A(n6427), .B(
        n6426), .ZN(n6428) );
  OAI21_X1 U8119 ( .B1(n6429), .B2(n8740), .A(n6428), .ZN(P1_U3220) );
  NAND4_X1 U8120 ( .A1(n6430), .A2(n6471), .A3(n10000), .A4(n6469), .ZN(n6432)
         );
  INV_X1 U8121 ( .A(n6465), .ZN(n6433) );
  INV_X1 U8122 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6444) );
  INV_X1 U8123 ( .A(n6434), .ZN(n6438) );
  INV_X1 U8124 ( .A(n6435), .ZN(n6487) );
  INV_X1 U8125 ( .A(n6436), .ZN(n6437) );
  AOI21_X1 U8126 ( .B1(n6438), .B2(n6487), .A(n6437), .ZN(n7221) );
  AND2_X1 U8127 ( .A1(n8020), .A2(n8152), .ZN(n6439) );
  NAND2_X1 U8128 ( .A1(n7036), .A2(n6439), .ZN(n10031) );
  INV_X1 U8129 ( .A(n6158), .ZN(n7147) );
  INV_X1 U8130 ( .A(n7184), .ZN(n7685) );
  AOI21_X1 U8131 ( .B1(n6434), .B2(n7685), .A(n8410), .ZN(n6440) );
  OAI21_X1 U8132 ( .B1(n7147), .B2(n7871), .A(n6440), .ZN(n6441) );
  AOI22_X1 U8133 ( .A1(n8048), .A2(n8343), .B1(n8341), .B2(n7183), .ZN(n6475)
         );
  AND2_X1 U8134 ( .A1(n6441), .A2(n6475), .ZN(n7216) );
  INV_X1 U8135 ( .A(n6479), .ZN(n10002) );
  INV_X1 U8136 ( .A(n8024), .ZN(n6474) );
  AND2_X2 U8137 ( .A1(n10002), .A2(n6474), .ZN(n10045) );
  AOI211_X1 U8138 ( .C1(n10001), .C2(n7217), .A(n10050), .B(n7154), .ZN(n7211)
         );
  AOI21_X1 U8139 ( .B1(n10045), .B2(n7217), .A(n7211), .ZN(n6442) );
  OAI211_X1 U8140 ( .C1(n7221), .C2(n10028), .A(n7216), .B(n6442), .ZN(n6446)
         );
  NAND2_X1 U8141 ( .A1(n10055), .A2(n6446), .ZN(n6443) );
  OAI21_X1 U8142 ( .B1(n10055), .B2(n6444), .A(n6443), .ZN(P2_U3454) );
  INV_X1 U8143 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6448) );
  NAND2_X1 U8144 ( .A1(n10069), .A2(n6446), .ZN(n6447) );
  OAI21_X1 U8145 ( .B1(n10069), .B2(n6448), .A(n6447), .ZN(P2_U3521) );
  NAND2_X1 U8146 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n8049), .ZN(n6449) );
  OAI21_X1 U8147 ( .B1(n8284), .B2(n8049), .A(n6449), .ZN(P2_U3575) );
  INV_X1 U8148 ( .A(n6450), .ZN(n6453) );
  AOI22_X1 U8149 ( .A1(n8128), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n8594), .ZN(n6451) );
  OAI21_X1 U8150 ( .B1(n6453), .B2(n8597), .A(n6451), .ZN(P2_U3341) );
  AOI22_X1 U8151 ( .A1(n9083), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9510), .ZN(n6452) );
  OAI21_X1 U8152 ( .B1(n6453), .B2(n9512), .A(n6452), .ZN(P1_U3336) );
  INV_X1 U8153 ( .A(n9068), .ZN(n9056) );
  OAI222_X1 U8154 ( .A1(n7689), .A2(n6455), .B1(n9056), .B2(P1_U3084), .C1(
        n9512), .C2(n6454), .ZN(P1_U3337) );
  OAI21_X1 U8155 ( .B1(n6458), .B2(n6457), .A(n6456), .ZN(n6459) );
  NAND2_X1 U8156 ( .A1(n6459), .A2(n8717), .ZN(n6463) );
  INV_X1 U8157 ( .A(n6500), .ZN(n6519) );
  OAI22_X1 U8158 ( .A1(n6519), .A2(n8732), .B1(n8720), .B2(n6807), .ZN(n6460)
         );
  AOI21_X1 U8159 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n6461), .A(n6460), .ZN(
        n6462) );
  OAI211_X1 U8160 ( .C1(n9403), .C2(n8726), .A(n6463), .B(n6462), .ZN(P1_U3235) );
  NAND2_X1 U8161 ( .A1(n6465), .A2(n6464), .ZN(n6470) );
  INV_X1 U8162 ( .A(n9994), .ZN(n6466) );
  INV_X1 U8163 ( .A(n6467), .ZN(n6468) );
  INV_X1 U8164 ( .A(n4310), .ZN(n7414) );
  NAND2_X1 U8165 ( .A1(n6470), .A2(n6469), .ZN(n6472) );
  NAND2_X1 U8166 ( .A1(n6472), .A2(n6471), .ZN(n6559) );
  INV_X1 U8167 ( .A(n6559), .ZN(n6473) );
  NAND2_X1 U8168 ( .A1(n6473), .A2(n10000), .ZN(n7682) );
  OR2_X1 U8169 ( .A1(n6492), .A2(n6474), .ZN(n7409) );
  INV_X1 U8170 ( .A(n7409), .ZN(n6477) );
  INV_X1 U8171 ( .A(n6475), .ZN(n6476) );
  AOI22_X1 U8172 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(n7682), .B1(n6477), .B2(
        n6476), .ZN(n6495) );
  NOR2_X1 U8173 ( .A1(n5789), .A2(n6478), .ZN(n6481) );
  XNOR2_X1 U8174 ( .A(n7217), .B(n6546), .ZN(n6482) );
  NAND2_X1 U8175 ( .A1(n6481), .A2(n6482), .ZN(n6485) );
  INV_X1 U8176 ( .A(n6481), .ZN(n6484) );
  INV_X1 U8177 ( .A(n6482), .ZN(n6483) );
  NAND2_X1 U8178 ( .A1(n6484), .A2(n6483), .ZN(n6542) );
  NOR2_X1 U8179 ( .A1(n10001), .A2(n6546), .ZN(n6486) );
  AOI21_X1 U8180 ( .B1(n6487), .B2(n6936), .A(n6486), .ZN(n6488) );
  OAI21_X1 U8181 ( .B1(n6489), .B2(n6488), .A(n6543), .ZN(n6493) );
  OR2_X1 U8182 ( .A1(n10045), .A2(n6490), .ZN(n6491) );
  NAND2_X1 U8183 ( .A1(n6493), .A2(n7789), .ZN(n6494) );
  OAI211_X1 U8184 ( .C1(n6496), .C2(n7414), .A(n6495), .B(n6494), .ZN(P2_U3224) );
  OR2_X1 U8185 ( .A1(n6497), .A2(n4940), .ZN(n6499) );
  NAND3_X1 U8186 ( .A1(n4515), .A2(n5663), .A3(n9005), .ZN(n6498) );
  NAND2_X1 U8187 ( .A1(n6502), .A2(n6501), .ZN(n6517) );
  OAI21_X1 U8188 ( .B1(n6501), .B2(n6502), .A(n6517), .ZN(n7070) );
  NAND2_X1 U8189 ( .A1(n5662), .A2(n9161), .ZN(n6504) );
  NAND2_X1 U8190 ( .A1(n5663), .A2(n9002), .ZN(n6503) );
  INV_X1 U8191 ( .A(n6501), .ZN(n6506) );
  NAND2_X1 U8192 ( .A1(n6506), .A2(n6505), .ZN(n6521) );
  OAI21_X1 U8193 ( .B1(n6506), .B2(n6505), .A(n6521), .ZN(n6508) );
  AOI222_X1 U8194 ( .A1(n9768), .A2(n6508), .B1(n9028), .B2(n9772), .C1(n9026), 
        .C2(n9771), .ZN(n7075) );
  INV_X1 U8195 ( .A(n8969), .ZN(n6518) );
  OR2_X1 U8196 ( .A1(n6509), .A2(n8969), .ZN(n6510) );
  OR2_X1 U8197 ( .A1(n6518), .A2(n7019), .ZN(n6525) );
  AND3_X1 U8198 ( .A1(n6510), .A2(n9816), .A3(n6525), .ZN(n7073) );
  AOI21_X1 U8199 ( .B1(n9935), .B2(n6518), .A(n7073), .ZN(n6511) );
  OAI211_X1 U8200 ( .C1(n9932), .C2(n7070), .A(n7075), .B(n6511), .ZN(n6513)
         );
  NAND2_X1 U8201 ( .A1(n6513), .A2(n9980), .ZN(n6512) );
  OAI21_X1 U8202 ( .B1(n9980), .B2(n4954), .A(n6512), .ZN(P1_U3524) );
  INV_X1 U8203 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6515) );
  NAND2_X1 U8204 ( .A1(n6513), .A2(n9971), .ZN(n6514) );
  OAI21_X1 U8205 ( .B1(n9971), .B2(n6515), .A(n6514), .ZN(P1_U3457) );
  NAND2_X1 U8206 ( .A1(n6500), .A2(n6518), .ZN(n6516) );
  INV_X1 U8207 ( .A(n9407), .ZN(n6529) );
  NAND2_X1 U8208 ( .A1(n6519), .A2(n6518), .ZN(n6520) );
  XNOR2_X1 U8209 ( .A(n8872), .B(n6809), .ZN(n6524) );
  NAND2_X1 U8210 ( .A1(n9407), .A2(n9805), .ZN(n6523) );
  AOI22_X1 U8211 ( .A1(n9025), .A2(n9771), .B1(n9772), .B2(n6500), .ZN(n6522)
         );
  OAI211_X1 U8212 ( .C1(n9802), .C2(n6524), .A(n6523), .B(n6522), .ZN(n9400)
         );
  INV_X1 U8213 ( .A(n9400), .ZN(n6528) );
  INV_X1 U8214 ( .A(n9403), .ZN(n6810) );
  AND2_X1 U8215 ( .A1(n6810), .A2(n6525), .ZN(n6526) );
  NOR2_X1 U8216 ( .A1(n7051), .A2(n6526), .ZN(n9406) );
  AOI22_X1 U8217 ( .A1(n9406), .A2(n9816), .B1(n9935), .B2(n6810), .ZN(n6527)
         );
  OAI211_X1 U8218 ( .C1(n6529), .C2(n9824), .A(n6528), .B(n6527), .ZN(n6531)
         );
  NAND2_X1 U8219 ( .A1(n6531), .A2(n9971), .ZN(n6530) );
  OAI21_X1 U8220 ( .B1(n9971), .B2(n4971), .A(n6530), .ZN(P1_U3460) );
  NAND2_X1 U8221 ( .A1(n6531), .A2(n9980), .ZN(n6532) );
  OAI21_X1 U8222 ( .B1(n9980), .B2(n4973), .A(n6532), .ZN(P1_U3525) );
  OAI21_X1 U8223 ( .B1(n6534), .B2(n6533), .A(n6584), .ZN(n6535) );
  NAND2_X1 U8224 ( .A1(n6535), .A2(n8717), .ZN(n6541) );
  NOR2_X1 U8225 ( .A1(n8726), .A2(n9927), .ZN(n6539) );
  OR2_X1 U8226 ( .A1(n8732), .A2(n7046), .ZN(n6537) );
  OAI211_X1 U8227 ( .C1(n8720), .C2(n7045), .A(n6537), .B(n6536), .ZN(n6538)
         );
  NOR2_X1 U8228 ( .A1(n6539), .A2(n6538), .ZN(n6540) );
  OAI211_X1 U8229 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8736), .A(n6541), .B(
        n6540), .ZN(P1_U3216) );
  OR2_X1 U8230 ( .A1(n6772), .A2(n6478), .ZN(n6544) );
  XNOR2_X1 U8231 ( .A(n7157), .B(n7650), .ZN(n6545) );
  XNOR2_X1 U8232 ( .A(n6544), .B(n6545), .ZN(n6671) );
  OAI22_X2 U8233 ( .A1(n6672), .A2(n6671), .B1(n6545), .B2(n6544), .ZN(n6749)
         );
  OR2_X1 U8234 ( .A1(n7165), .A2(n6478), .ZN(n6547) );
  XNOR2_X1 U8235 ( .A(n6777), .B(n7666), .ZN(n6548) );
  XNOR2_X1 U8236 ( .A(n6547), .B(n6548), .ZN(n6748) );
  NAND2_X1 U8237 ( .A1(n6749), .A2(n6748), .ZN(n6551) );
  INV_X1 U8238 ( .A(n6547), .ZN(n6549) );
  NAND2_X1 U8239 ( .A1(n6549), .A2(n6548), .ZN(n6550) );
  NAND2_X1 U8240 ( .A1(n6551), .A2(n6550), .ZN(n6758) );
  INV_X1 U8241 ( .A(n6758), .ZN(n6555) );
  OR2_X1 U8242 ( .A1(n6771), .A2(n8539), .ZN(n6553) );
  XNOR2_X1 U8243 ( .A(n7176), .B(n7650), .ZN(n6552) );
  NAND2_X1 U8244 ( .A1(n6553), .A2(n6552), .ZN(n6556) );
  OAI21_X1 U8245 ( .B1(n6553), .B2(n6552), .A(n6556), .ZN(n6757) );
  INV_X1 U8246 ( .A(n6757), .ZN(n6554) );
  OR2_X1 U8247 ( .A1(n7166), .A2(n8539), .ZN(n6791) );
  XNOR2_X1 U8248 ( .A(n7275), .B(n7650), .ZN(n6792) );
  XNOR2_X1 U8249 ( .A(n6791), .B(n6792), .ZN(n6790) );
  XNOR2_X1 U8250 ( .A(n6789), .B(n6790), .ZN(n6565) );
  INV_X1 U8251 ( .A(n6557), .ZN(n6558) );
  OR2_X1 U8252 ( .A1(n6559), .A2(n6558), .ZN(n6560) );
  AOI22_X1 U8253 ( .A1(n8047), .A2(n8341), .B1(n8343), .B2(n8045), .ZN(n7279)
         );
  INV_X1 U8254 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6561) );
  OAI22_X1 U8255 ( .A1(n7409), .A2(n7279), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6561), .ZN(n6563) );
  NOR2_X1 U8256 ( .A1(n7414), .A2(n10019), .ZN(n6562) );
  AOI211_X1 U8257 ( .C1(n7794), .C2(n7274), .A(n6563), .B(n6562), .ZN(n6564)
         );
  OAI21_X1 U8258 ( .B1(n6565), .B2(n7810), .A(n6564), .ZN(P2_U3229) );
  AOI22_X1 U8259 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n6575), .B1(n9037), .B2(
        n5206), .ZN(n9035) );
  OAI21_X1 U8260 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n6574), .A(n6566), .ZN(
        n9034) );
  NAND2_X1 U8261 ( .A1(n9035), .A2(n9034), .ZN(n9033) );
  OAI21_X1 U8262 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6575), .A(n9033), .ZN(
        n6569) );
  MUX2_X1 U8263 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6567), .S(n6847), .Z(n6568)
         );
  NAND2_X1 U8264 ( .A1(n6568), .A2(n6569), .ZN(n6840) );
  OAI21_X1 U8265 ( .B1(n6569), .B2(n6568), .A(n6840), .ZN(n6581) );
  INV_X1 U8266 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6571) );
  NAND2_X1 U8267 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7452) );
  NAND2_X1 U8268 ( .A1(n9912), .A2(n6847), .ZN(n6570) );
  OAI211_X1 U8269 ( .C1(n9925), .C2(n6571), .A(n7452), .B(n6570), .ZN(n6580)
         );
  NOR2_X1 U8270 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6575), .ZN(n6572) );
  AOI21_X1 U8271 ( .B1(n6575), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6572), .ZN(
        n9031) );
  NAND2_X1 U8272 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6847), .ZN(n6576) );
  OAI21_X1 U8273 ( .B1(n6847), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6576), .ZN(
        n6577) );
  AOI211_X1 U8274 ( .C1(n6578), .C2(n6577), .A(n6846), .B(n9885), .ZN(n6579)
         );
  AOI211_X1 U8275 ( .C1(n9920), .C2(n6581), .A(n6580), .B(n6579), .ZN(n6582)
         );
  INV_X1 U8276 ( .A(n6582), .ZN(P1_U3253) );
  AND2_X1 U8277 ( .A1(n6584), .A2(n6583), .ZN(n6587) );
  OAI211_X1 U8278 ( .C1(n6587), .C2(n6586), .A(n8717), .B(n6585), .ZN(n6593)
         );
  INV_X1 U8279 ( .A(n6816), .ZN(n7060) );
  NOR2_X1 U8280 ( .A1(n8726), .A2(n7060), .ZN(n6591) );
  OR2_X1 U8281 ( .A1(n8732), .A2(n6807), .ZN(n6589) );
  AND2_X1 U8282 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9862) );
  INV_X1 U8283 ( .A(n9862), .ZN(n6588) );
  OAI211_X1 U8284 ( .C1(n8720), .C2(n7129), .A(n6589), .B(n6588), .ZN(n6590)
         );
  NOR2_X1 U8285 ( .A1(n6591), .A2(n6590), .ZN(n6592) );
  OAI211_X1 U8286 ( .C1(n8736), .C2(n7061), .A(n6593), .B(n6592), .ZN(P1_U3228) );
  INV_X1 U8287 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6595) );
  INV_X1 U8288 ( .A(n6594), .ZN(n6596) );
  INV_X1 U8289 ( .A(n8145), .ZN(n8134) );
  OAI222_X1 U8290 ( .A1(n7365), .A2(n6595), .B1(n7545), .B2(n6596), .C1(n7694), 
        .C2(n8134), .ZN(P2_U3340) );
  INV_X1 U8291 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6597) );
  INV_X1 U8292 ( .A(n9911), .ZN(n9080) );
  OAI222_X1 U8293 ( .A1(n7689), .A2(n6597), .B1(n9512), .B2(n6596), .C1(
        P1_U3084), .C2(n9080), .ZN(P1_U3335) );
  NAND2_X1 U8294 ( .A1(n9994), .A2(n6598), .ZN(n6602) );
  NAND2_X1 U8295 ( .A1(n6616), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7567) );
  OAI21_X1 U8296 ( .B1(n6599), .B2(n7567), .A(n8029), .ZN(n6600) );
  INV_X1 U8297 ( .A(n6600), .ZN(n6601) );
  NAND2_X1 U8298 ( .A1(n6602), .A2(n6601), .ZN(n6604) );
  NAND2_X1 U8299 ( .A1(n6604), .A2(n6603), .ZN(n6608) );
  NAND2_X1 U8300 ( .A1(n6608), .A2(n8049), .ZN(n6615) );
  INV_X1 U8301 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6606) );
  INV_X1 U8302 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7152) );
  OAI22_X1 U8303 ( .A1(n8157), .A2(n6606), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7152), .ZN(n6614) );
  MUX2_X1 U8304 ( .A(n6448), .B(P2_REG1_REG_1__SCAN_IN), .S(n6618), .Z(n6711)
         );
  INV_X1 U8305 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10056) );
  INV_X1 U8306 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9990) );
  NOR3_X1 U8307 ( .A1(n6711), .A2(n10056), .A3(n9990), .ZN(n6710) );
  AOI21_X1 U8308 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(n6618), .A(n6710), .ZN(
        n6612) );
  INV_X1 U8309 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6607) );
  MUX2_X1 U8310 ( .A(n6607), .B(P2_REG1_REG_2__SCAN_IN), .S(n6635), .Z(n6611)
         );
  NOR2_X1 U8311 ( .A1(n6612), .A2(n6611), .ZN(n6629) );
  INV_X1 U8312 ( .A(n6608), .ZN(n6610) );
  AOI211_X1 U8313 ( .C1(n6612), .C2(n6611), .A(n6629), .B(n9983), .ZN(n6613)
         );
  AOI211_X1 U8314 ( .C1(n8150), .C2(n6635), .A(n6614), .B(n6613), .ZN(n6628)
         );
  NAND2_X1 U8315 ( .A1(n6615), .A2(n8025), .ZN(n8147) );
  INV_X1 U8316 ( .A(n8147), .ZN(n6617) );
  MUX2_X1 U8317 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6619), .S(n6618), .Z(n6716)
         );
  NAND3_X1 U8318 ( .A1(n6716), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_REG2_REG_0__SCAN_IN), .ZN(n6715) );
  INV_X1 U8319 ( .A(n6715), .ZN(n6622) );
  NOR2_X1 U8320 ( .A1(n5774), .A2(n6619), .ZN(n6623) );
  MUX2_X1 U8321 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6620), .S(n6635), .Z(n6621)
         );
  OAI21_X1 U8322 ( .B1(n6622), .B2(n6623), .A(n6621), .ZN(n6665) );
  MUX2_X1 U8323 ( .A(n6620), .B(P2_REG2_REG_2__SCAN_IN), .S(n6635), .Z(n6625)
         );
  INV_X1 U8324 ( .A(n6623), .ZN(n6624) );
  NAND3_X1 U8325 ( .A1(n6625), .A2(n6715), .A3(n6624), .ZN(n6626) );
  NAND3_X1 U8326 ( .A1(n9986), .A2(n6665), .A3(n6626), .ZN(n6627) );
  NAND2_X1 U8327 ( .A1(n6628), .A2(n6627), .ZN(P2_U3247) );
  NOR2_X1 U8328 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6561), .ZN(n6634) );
  AOI21_X1 U8329 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n6635), .A(n6629), .ZN(
        n6660) );
  XNOR2_X1 U8330 ( .A(n6636), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n6659) );
  NOR2_X1 U8331 ( .A1(n6660), .A2(n6659), .ZN(n6658) );
  AOI21_X1 U8332 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n6636), .A(n6658), .ZN(
        n6646) );
  XNOR2_X1 U8333 ( .A(n6650), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n6645) );
  NOR2_X1 U8334 ( .A1(n6646), .A2(n6645), .ZN(n6644) );
  NAND2_X1 U8335 ( .A1(n6683), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6630) );
  OAI21_X1 U8336 ( .B1(n6683), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6630), .ZN(
        n6631) );
  AOI211_X1 U8337 ( .C1(n6632), .C2(n6631), .A(n6678), .B(n9983), .ZN(n6633)
         );
  AOI211_X1 U8338 ( .C1(n9987), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n6634), .B(
        n6633), .ZN(n6642) );
  NAND2_X1 U8339 ( .A1(n6635), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6664) );
  MUX2_X1 U8340 ( .A(n6637), .B(P2_REG2_REG_3__SCAN_IN), .S(n6636), .Z(n6663)
         );
  AOI21_X1 U8341 ( .B1(n6665), .B2(n6664), .A(n6663), .ZN(n6648) );
  NOR2_X1 U8342 ( .A1(n6670), .A2(n6637), .ZN(n6649) );
  MUX2_X1 U8343 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6639), .S(n6650), .Z(n6638)
         );
  OAI21_X1 U8344 ( .B1(n6648), .B2(n6649), .A(n6638), .ZN(n6654) );
  OAI21_X1 U8345 ( .B1(n6639), .B2(n6657), .A(n6654), .ZN(n6686) );
  MUX2_X1 U8346 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n5828), .S(n6643), .Z(n6684)
         );
  XNOR2_X1 U8347 ( .A(n6686), .B(n6684), .ZN(n6640) );
  NAND2_X1 U8348 ( .A1(n9986), .A2(n6640), .ZN(n6641) );
  OAI211_X1 U8349 ( .C1(n9982), .C2(n6643), .A(n6642), .B(n6641), .ZN(P2_U3250) );
  INV_X1 U8350 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9671) );
  NOR2_X1 U8351 ( .A1(n9671), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6759) );
  AOI211_X1 U8352 ( .C1(n6646), .C2(n6645), .A(n6644), .B(n9983), .ZN(n6647)
         );
  AOI211_X1 U8353 ( .C1(n9987), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6759), .B(
        n6647), .ZN(n6656) );
  INV_X1 U8354 ( .A(n6648), .ZN(n6667) );
  INV_X1 U8355 ( .A(n6649), .ZN(n6652) );
  MUX2_X1 U8356 ( .A(n6639), .B(P2_REG2_REG_4__SCAN_IN), .S(n6650), .Z(n6651)
         );
  NAND3_X1 U8357 ( .A1(n6667), .A2(n6652), .A3(n6651), .ZN(n6653) );
  NAND3_X1 U8358 ( .A1(n9986), .A2(n6654), .A3(n6653), .ZN(n6655) );
  OAI211_X1 U8359 ( .C1(n9982), .C2(n6657), .A(n6656), .B(n6655), .ZN(P2_U3249) );
  NOR2_X1 U8360 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6752), .ZN(n6662) );
  AOI211_X1 U8361 ( .C1(n6660), .C2(n6659), .A(n6658), .B(n9983), .ZN(n6661)
         );
  AOI211_X1 U8362 ( .C1(n9987), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6662), .B(
        n6661), .ZN(n6669) );
  NAND3_X1 U8363 ( .A1(n6665), .A2(n6664), .A3(n6663), .ZN(n6666) );
  NAND3_X1 U8364 ( .A1(n9986), .A2(n6667), .A3(n6666), .ZN(n6668) );
  OAI211_X1 U8365 ( .C1(n9982), .C2(n6670), .A(n6669), .B(n6668), .ZN(P2_U3248) );
  XNOR2_X1 U8366 ( .A(n6672), .B(n6671), .ZN(n6677) );
  NOR2_X2 U8367 ( .A1(n7409), .A2(n6188), .ZN(n7795) );
  AOI22_X1 U8368 ( .A1(n7795), .A2(n6673), .B1(n7793), .B2(n6674), .ZN(n6676)
         );
  AOI22_X1 U8369 ( .A1(n7157), .A2(n4310), .B1(n7682), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n6675) );
  OAI211_X1 U8370 ( .C1(n6677), .C2(n7810), .A(n6676), .B(n6675), .ZN(P2_U3239) );
  INV_X1 U8371 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9694) );
  NOR2_X1 U8372 ( .A1(n9694), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6797) );
  NAND2_X1 U8373 ( .A1(n6701), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6679) );
  OAI21_X1 U8374 ( .B1(n6701), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6679), .ZN(
        n6680) );
  AOI211_X1 U8375 ( .C1(n6681), .C2(n6680), .A(n6695), .B(n9983), .ZN(n6682)
         );
  AOI211_X1 U8376 ( .C1(n9987), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n6797), .B(
        n6682), .ZN(n6693) );
  NAND2_X1 U8377 ( .A1(n6683), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6688) );
  INV_X1 U8378 ( .A(n6684), .ZN(n6685) );
  NAND2_X1 U8379 ( .A1(n6686), .A2(n6685), .ZN(n6687) );
  NAND2_X1 U8380 ( .A1(n6688), .A2(n6687), .ZN(n6691) );
  MUX2_X1 U8381 ( .A(n7025), .B(P2_REG2_REG_6__SCAN_IN), .S(n6701), .Z(n6689)
         );
  INV_X1 U8382 ( .A(n6689), .ZN(n6690) );
  NAND2_X1 U8383 ( .A1(n6690), .A2(n6691), .ZN(n6702) );
  OAI211_X1 U8384 ( .C1(n6691), .C2(n6690), .A(n9986), .B(n6702), .ZN(n6692)
         );
  OAI211_X1 U8385 ( .C1(n9982), .C2(n6694), .A(n6693), .B(n6692), .ZN(P2_U3251) );
  NOR2_X1 U8386 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5852), .ZN(n6700) );
  AOI21_X1 U8387 ( .B1(n6701), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6695), .ZN(
        n6698) );
  NAND2_X1 U8388 ( .A1(n6732), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6696) );
  OAI21_X1 U8389 ( .B1(n6732), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6696), .ZN(
        n6697) );
  NOR2_X1 U8390 ( .A1(n6698), .A2(n6697), .ZN(n6731) );
  AOI211_X1 U8391 ( .C1(n6698), .C2(n6697), .A(n6731), .B(n9983), .ZN(n6699)
         );
  AOI211_X1 U8392 ( .C1(n9987), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n6700), .B(
        n6699), .ZN(n6708) );
  NAND2_X1 U8393 ( .A1(n6701), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6703) );
  NAND2_X1 U8394 ( .A1(n6703), .A2(n6702), .ZN(n6706) );
  MUX2_X1 U8395 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6704), .S(n6732), .Z(n6705)
         );
  NAND2_X1 U8396 ( .A1(n6705), .A2(n6706), .ZN(n6723) );
  OAI211_X1 U8397 ( .C1(n6706), .C2(n6705), .A(n9986), .B(n6723), .ZN(n6707)
         );
  OAI211_X1 U8398 ( .C1(n9982), .C2(n6709), .A(n6708), .B(n6707), .ZN(P2_U3252) );
  INV_X1 U8399 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10074) );
  NOR2_X1 U8400 ( .A1(n8157), .A2(n10074), .ZN(n6714) );
  NAND2_X1 U8401 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n6712) );
  AOI211_X1 U8402 ( .C1(n6712), .C2(n6711), .A(n6710), .B(n9983), .ZN(n6713)
         );
  AOI211_X1 U8403 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(P2_U3152), .A(n6714), .B(
        n6713), .ZN(n6719) );
  AND2_X1 U8404 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n6717) );
  OAI211_X1 U8405 ( .C1(n6717), .C2(n6716), .A(n9986), .B(n6715), .ZN(n6718)
         );
  OAI211_X1 U8406 ( .C1(n9982), .C2(n5774), .A(n6719), .B(n6718), .ZN(P2_U3246) );
  NAND2_X1 U8407 ( .A1(n8081), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6727) );
  MUX2_X1 U8408 ( .A(n7354), .B(P2_REG2_REG_10__SCAN_IN), .S(n8081), .Z(n6720)
         );
  INV_X1 U8409 ( .A(n6720), .ZN(n8078) );
  NAND2_X1 U8410 ( .A1(n8068), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6726) );
  MUX2_X1 U8411 ( .A(n5884), .B(P2_REG2_REG_9__SCAN_IN), .S(n8068), .Z(n6721)
         );
  INV_X1 U8412 ( .A(n6721), .ZN(n8064) );
  NAND2_X1 U8413 ( .A1(n8054), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6725) );
  MUX2_X1 U8414 ( .A(n5868), .B(P2_REG2_REG_8__SCAN_IN), .S(n8054), .Z(n6722)
         );
  INV_X1 U8415 ( .A(n6722), .ZN(n8051) );
  NAND2_X1 U8416 ( .A1(n6732), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6724) );
  NAND2_X1 U8417 ( .A1(n6724), .A2(n6723), .ZN(n8052) );
  NAND2_X1 U8418 ( .A1(n8051), .A2(n8052), .ZN(n8050) );
  NAND2_X1 U8419 ( .A1(n6725), .A2(n8050), .ZN(n8065) );
  NAND2_X1 U8420 ( .A1(n8064), .A2(n8065), .ZN(n8063) );
  NAND2_X1 U8421 ( .A1(n6726), .A2(n8063), .ZN(n8079) );
  NAND2_X1 U8422 ( .A1(n8078), .A2(n8079), .ZN(n8077) );
  NAND2_X1 U8423 ( .A1(n6727), .A2(n8077), .ZN(n6730) );
  MUX2_X1 U8424 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n5913), .S(n6829), .Z(n6728)
         );
  INV_X1 U8425 ( .A(n6728), .ZN(n6729) );
  NOR2_X1 U8426 ( .A1(n6730), .A2(n6729), .ZN(n6822) );
  AOI21_X1 U8427 ( .B1(n6730), .B2(n6729), .A(n6822), .ZN(n6743) );
  NOR2_X1 U8428 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7407), .ZN(n6740) );
  AOI21_X1 U8429 ( .B1(n6732), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6731), .ZN(
        n8056) );
  INV_X1 U8430 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6733) );
  MUX2_X1 U8431 ( .A(n6733), .B(P2_REG1_REG_8__SCAN_IN), .S(n8054), .Z(n8057)
         );
  INV_X1 U8432 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6734) );
  MUX2_X1 U8433 ( .A(n6734), .B(P2_REG1_REG_9__SCAN_IN), .S(n8068), .Z(n8071)
         );
  INV_X1 U8434 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6735) );
  MUX2_X1 U8435 ( .A(n6735), .B(P2_REG1_REG_10__SCAN_IN), .S(n8081), .Z(n8083)
         );
  NOR2_X1 U8436 ( .A1(n4332), .A2(n8083), .ZN(n8082) );
  INV_X1 U8437 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6736) );
  MUX2_X1 U8438 ( .A(n6736), .B(P2_REG1_REG_11__SCAN_IN), .S(n6829), .Z(n6737)
         );
  AOI211_X1 U8439 ( .C1(n6738), .C2(n6737), .A(n6828), .B(n9983), .ZN(n6739)
         );
  AOI211_X1 U8440 ( .C1(n9987), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n6740), .B(
        n6739), .ZN(n6742) );
  NAND2_X1 U8441 ( .A1(n8150), .A2(n6829), .ZN(n6741) );
  OAI211_X1 U8442 ( .C1(n6743), .C2(n8138), .A(n6742), .B(n6741), .ZN(P2_U3256) );
  INV_X1 U8443 ( .A(n6744), .ZN(n6746) );
  OAI222_X1 U8444 ( .A1(n7689), .A2(n6745), .B1(n9512), .B2(n6746), .C1(n9001), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  OAI222_X1 U8445 ( .A1(n7365), .A2(n6747), .B1(n7545), .B2(n6746), .C1(n7694), 
        .C2(n7833), .ZN(P2_U3339) );
  XNOR2_X1 U8446 ( .A(n6749), .B(n6748), .ZN(n6754) );
  OAI22_X1 U8447 ( .A1(n7414), .A2(n7086), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6752), .ZN(n6751) );
  OAI22_X1 U8448 ( .A1(n6772), .A2(n7806), .B1(n7803), .B2(n6771), .ZN(n6750)
         );
  AOI211_X1 U8449 ( .C1(n7794), .C2(n6752), .A(n6751), .B(n6750), .ZN(n6753)
         );
  OAI21_X1 U8450 ( .B1(n7810), .B2(n6754), .A(n6753), .ZN(P2_U3220) );
  INV_X1 U8451 ( .A(n6755), .ZN(n6756) );
  AOI21_X1 U8452 ( .B1(n6758), .B2(n6757), .A(n6756), .ZN(n6765) );
  INV_X1 U8453 ( .A(n6759), .ZN(n6760) );
  OAI21_X1 U8454 ( .B1(n7414), .B2(n10014), .A(n6760), .ZN(n6762) );
  OAI22_X1 U8455 ( .A1(n7166), .A2(n7803), .B1(n7806), .B2(n7165), .ZN(n6761)
         );
  AOI211_X1 U8456 ( .C1(n6763), .C2(n7794), .A(n6762), .B(n6761), .ZN(n6764)
         );
  OAI21_X1 U8457 ( .B1(n6765), .B2(n7810), .A(n6764), .ZN(P2_U3232) );
  INV_X1 U8458 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6781) );
  NAND2_X1 U8459 ( .A1(n7158), .A2(n6766), .ZN(n6768) );
  NAND2_X1 U8460 ( .A1(n6768), .A2(n6160), .ZN(n6767) );
  OAI21_X1 U8461 ( .B1(n6768), .B2(n6160), .A(n6767), .ZN(n7088) );
  INV_X1 U8462 ( .A(n7088), .ZN(n6779) );
  OAI21_X1 U8463 ( .B1(n7879), .B2(n6770), .A(n6769), .ZN(n6775) );
  OAI22_X1 U8464 ( .A1(n6772), .A2(n6188), .B1(n6771), .B2(n8430), .ZN(n6774)
         );
  NOR2_X1 U8465 ( .A1(n6779), .A2(n8427), .ZN(n6773) );
  AOI211_X1 U8466 ( .C1(n8434), .C2(n6775), .A(n6774), .B(n6773), .ZN(n7090)
         );
  AOI21_X1 U8467 ( .B1(n7153), .B2(n6777), .A(n10050), .ZN(n6776) );
  AND2_X1 U8468 ( .A1(n6776), .A2(n7171), .ZN(n7084) );
  AOI21_X1 U8469 ( .B1(n10045), .B2(n6777), .A(n7084), .ZN(n6778) );
  OAI211_X1 U8470 ( .C1(n6779), .C2(n10031), .A(n7090), .B(n6778), .ZN(n6782)
         );
  NAND2_X1 U8471 ( .A1(n6782), .A2(n10069), .ZN(n6780) );
  OAI21_X1 U8472 ( .B1(n10069), .B2(n6781), .A(n6780), .ZN(P2_U3523) );
  NAND2_X1 U8473 ( .A1(n6782), .A2(n10055), .ZN(n6783) );
  OAI21_X1 U8474 ( .B1(n10055), .B2(n5799), .A(n6783), .ZN(P2_U3460) );
  AND2_X1 U8475 ( .A1(n8045), .A2(n10050), .ZN(n6784) );
  XNOR2_X1 U8476 ( .A(n10024), .B(n7666), .ZN(n6785) );
  NAND2_X1 U8477 ( .A1(n6784), .A2(n6785), .ZN(n6788) );
  INV_X1 U8478 ( .A(n6784), .ZN(n6787) );
  INV_X1 U8479 ( .A(n6785), .ZN(n6786) );
  NAND2_X1 U8480 ( .A1(n6787), .A2(n6786), .ZN(n6856) );
  AND2_X1 U8481 ( .A1(n6788), .A2(n6856), .ZN(n6796) );
  INV_X1 U8482 ( .A(n6791), .ZN(n6794) );
  INV_X1 U8483 ( .A(n6792), .ZN(n6793) );
  OAI21_X1 U8484 ( .B1(n6796), .B2(n6795), .A(n6857), .ZN(n6802) );
  OAI22_X1 U8485 ( .A1(n7166), .A2(n7806), .B1(n7803), .B2(n6914), .ZN(n6801)
         );
  INV_X1 U8486 ( .A(n6797), .ZN(n6799) );
  NAND2_X1 U8487 ( .A1(n7794), .A2(n7028), .ZN(n6798) );
  OAI211_X1 U8488 ( .C1(n7414), .C2(n7030), .A(n6799), .B(n6798), .ZN(n6800)
         );
  AOI211_X1 U8489 ( .C1(n6802), .C2(n7789), .A(n6801), .B(n6800), .ZN(n6803)
         );
  INV_X1 U8490 ( .A(n6803), .ZN(P2_U3241) );
  NAND2_X1 U8491 ( .A1(n7046), .A2(n9403), .ZN(n6804) );
  NAND2_X1 U8492 ( .A1(n6807), .A2(n7056), .ZN(n8910) );
  NAND2_X1 U8493 ( .A1(n9927), .A2(n9025), .ZN(n8973) );
  NAND2_X1 U8494 ( .A1(n8910), .A2(n8973), .ZN(n7040) );
  NAND2_X1 U8495 ( .A1(n6807), .A2(n9927), .ZN(n6805) );
  NAND2_X1 U8496 ( .A1(n7039), .A2(n6805), .ZN(n6806) );
  NAND2_X1 U8497 ( .A1(n7045), .A2(n6816), .ZN(n6958) );
  INV_X1 U8498 ( .A(n7045), .ZN(n9024) );
  NAND2_X1 U8499 ( .A1(n7060), .A2(n9024), .ZN(n8912) );
  NAND2_X1 U8500 ( .A1(n6958), .A2(n8912), .ZN(n8867) );
  OAI21_X1 U8501 ( .B1(n6806), .B2(n8867), .A(n6954), .ZN(n7066) );
  INV_X1 U8502 ( .A(n7066), .ZN(n6818) );
  OAI22_X1 U8503 ( .A1(n6807), .A2(n9798), .B1(n7129), .B2(n9796), .ZN(n6815)
         );
  INV_X1 U8504 ( .A(n8872), .ZN(n6808) );
  NAND2_X1 U8505 ( .A1(n6809), .A2(n6808), .ZN(n6812) );
  NAND2_X1 U8506 ( .A1(n7046), .A2(n6810), .ZN(n6811) );
  NAND2_X1 U8507 ( .A1(n6812), .A2(n6811), .ZN(n7043) );
  NAND2_X1 U8508 ( .A1(n7043), .A2(n8868), .ZN(n7044) );
  XNOR2_X1 U8509 ( .A(n6959), .B(n8867), .ZN(n6813) );
  NOR2_X1 U8510 ( .A1(n6813), .A2(n9802), .ZN(n6814) );
  AOI211_X1 U8511 ( .C1(n9805), .C2(n7066), .A(n6815), .B(n6814), .ZN(n7069)
         );
  NAND2_X1 U8512 ( .A1(n7051), .A2(n9927), .ZN(n7053) );
  AOI21_X1 U8513 ( .B1(n6816), .B2(n7053), .A(n4498), .ZN(n7065) );
  AOI22_X1 U8514 ( .A1(n7065), .A2(n9816), .B1(n9935), .B2(n6816), .ZN(n6817)
         );
  OAI211_X1 U8515 ( .C1(n6818), .C2(n9824), .A(n7069), .B(n6817), .ZN(n6820)
         );
  NAND2_X1 U8516 ( .A1(n6820), .A2(n9980), .ZN(n6819) );
  OAI21_X1 U8517 ( .B1(n9980), .B2(n5014), .A(n6819), .ZN(P1_U3527) );
  NAND2_X1 U8518 ( .A1(n6820), .A2(n9971), .ZN(n6821) );
  OAI21_X1 U8519 ( .B1(n9971), .B2(n5011), .A(n6821), .ZN(P1_U3466) );
  NOR2_X1 U8520 ( .A1(n6829), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6823) );
  NOR2_X1 U8521 ( .A1(n6823), .A2(n6822), .ZN(n6826) );
  MUX2_X1 U8522 ( .A(n7463), .B(P2_REG2_REG_12__SCAN_IN), .S(n6901), .Z(n6824)
         );
  INV_X1 U8523 ( .A(n6824), .ZN(n6825) );
  NAND2_X1 U8524 ( .A1(n6825), .A2(n6826), .ZN(n6896) );
  OAI211_X1 U8525 ( .C1(n6826), .C2(n6825), .A(n9986), .B(n6896), .ZN(n6837)
         );
  INV_X1 U8526 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6827) );
  MUX2_X1 U8527 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6827), .S(n6901), .Z(n6831)
         );
  OAI21_X1 U8528 ( .B1(n6831), .B2(n6830), .A(n6900), .ZN(n6835) );
  NAND2_X1 U8529 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7494) );
  INV_X1 U8530 ( .A(n7494), .ZN(n6834) );
  INV_X1 U8531 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6832) );
  NOR2_X1 U8532 ( .A1(n8157), .A2(n6832), .ZN(n6833) );
  AOI211_X1 U8533 ( .C1(n9981), .C2(n6835), .A(n6834), .B(n6833), .ZN(n6836)
         );
  OAI211_X1 U8534 ( .C1(n9982), .C2(n6838), .A(n6837), .B(n6836), .ZN(P2_U3257) );
  INV_X1 U8535 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6855) );
  OR2_X1 U8536 ( .A1(n7199), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7193) );
  NAND2_X1 U8537 ( .A1(n7199), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6839) );
  AND2_X1 U8538 ( .A1(n7193), .A2(n6839), .ZN(n6843) );
  OR2_X1 U8539 ( .A1(n6847), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6841) );
  NAND2_X1 U8540 ( .A1(n6841), .A2(n6840), .ZN(n6842) );
  NAND2_X1 U8541 ( .A1(n6843), .A2(n6842), .ZN(n7192) );
  OAI21_X1 U8542 ( .B1(n6843), .B2(n6842), .A(n7192), .ZN(n6844) );
  NAND2_X1 U8543 ( .A1(n9920), .A2(n6844), .ZN(n6845) );
  NAND2_X1 U8544 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7476) );
  NAND2_X1 U8545 ( .A1(n6845), .A2(n7476), .ZN(n6853) );
  AOI21_X1 U8546 ( .B1(n6847), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6846), .ZN(
        n6851) );
  NOR2_X1 U8547 ( .A1(n7199), .A2(n6848), .ZN(n6849) );
  AOI21_X1 U8548 ( .B1(n7199), .B2(n6848), .A(n6849), .ZN(n6850) );
  AOI211_X1 U8549 ( .C1(n6851), .C2(n6850), .A(n7198), .B(n9885), .ZN(n6852)
         );
  AOI211_X1 U8550 ( .C1(n9912), .C2(n7199), .A(n6853), .B(n6852), .ZN(n6854)
         );
  OAI21_X1 U8551 ( .B1(n9925), .B2(n6855), .A(n6854), .ZN(P1_U3254) );
  OR2_X1 U8552 ( .A1(n6914), .A2(n8539), .ZN(n6910) );
  XNOR2_X1 U8553 ( .A(n6937), .B(n7650), .ZN(n6911) );
  XNOR2_X1 U8554 ( .A(n6910), .B(n6911), .ZN(n6912) );
  XNOR2_X1 U8555 ( .A(n6913), .B(n6912), .ZN(n6863) );
  OAI22_X1 U8556 ( .A1(n7414), .A2(n6991), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5852), .ZN(n6860) );
  OAI22_X1 U8557 ( .A1(n6858), .A2(n7806), .B1(n7803), .B2(n7313), .ZN(n6859)
         );
  AOI211_X1 U8558 ( .C1(n6861), .C2(n7794), .A(n6860), .B(n6859), .ZN(n6862)
         );
  OAI21_X1 U8559 ( .B1(n6863), .B2(n7810), .A(n6862), .ZN(P2_U3215) );
  INV_X1 U8560 ( .A(n6864), .ZN(n6867) );
  OAI222_X1 U8561 ( .A1(n9512), .A2(n6867), .B1(P1_U3084), .B2(n6866), .C1(
        n6865), .C2(n7689), .ZN(P1_U3333) );
  OAI222_X1 U8562 ( .A1(n7365), .A2(n6868), .B1(n7545), .B2(n6867), .C1(n8020), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  INV_X1 U8563 ( .A(n6869), .ZN(n6871) );
  OAI222_X1 U8564 ( .A1(n9512), .A2(n6871), .B1(P1_U3084), .B2(n6948), .C1(
        n6870), .C2(n7689), .ZN(P1_U3332) );
  INV_X1 U8565 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6872) );
  OAI222_X1 U8566 ( .A1(n7365), .A2(n6872), .B1(n7545), .B2(n6871), .C1(n7815), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  INV_X1 U8567 ( .A(n6873), .ZN(n6924) );
  INV_X1 U8568 ( .A(n6874), .ZN(n6876) );
  NOR3_X1 U8569 ( .A1(n6924), .A2(n6876), .A3(n6875), .ZN(n6879) );
  INV_X1 U8570 ( .A(n6877), .ZN(n6878) );
  OAI21_X1 U8571 ( .B1(n6879), .B2(n6878), .A(n8717), .ZN(n6884) );
  AOI21_X1 U8572 ( .B1(n8734), .B2(n9020), .A(n6880), .ZN(n6881) );
  OAI21_X1 U8573 ( .B1(n7233), .B2(n8732), .A(n6881), .ZN(n6882) );
  AOI21_X1 U8574 ( .B1(n8738), .B2(n7246), .A(n6882), .ZN(n6883) );
  OAI211_X1 U8575 ( .C1(n8736), .C2(n7243), .A(n6884), .B(n6883), .ZN(P1_U3211) );
  NAND2_X1 U8576 ( .A1(n4382), .A2(n6885), .ZN(n6920) );
  OAI21_X1 U8577 ( .B1(n4382), .B2(n6885), .A(n6920), .ZN(n6886) );
  NOR2_X1 U8578 ( .A1(n6886), .A2(n6887), .ZN(n6923) );
  AOI21_X1 U8579 ( .B1(n6887), .B2(n6886), .A(n6923), .ZN(n6895) );
  INV_X1 U8580 ( .A(n9934), .ZN(n6968) );
  NOR2_X1 U8581 ( .A1(n8726), .A2(n6968), .ZN(n6891) );
  OR2_X1 U8582 ( .A1(n8732), .A2(n7045), .ZN(n6889) );
  AND2_X1 U8583 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9871) );
  INV_X1 U8584 ( .A(n9871), .ZN(n6888) );
  OAI211_X1 U8585 ( .C1(n8720), .C2(n7233), .A(n6889), .B(n6888), .ZN(n6890)
         );
  NOR2_X1 U8586 ( .A1(n6891), .A2(n6890), .ZN(n6894) );
  INV_X1 U8587 ( .A(n6964), .ZN(n6892) );
  NAND2_X1 U8588 ( .A1(n8723), .A2(n6892), .ZN(n6893) );
  OAI211_X1 U8589 ( .C1(n6895), .C2(n8740), .A(n6894), .B(n6893), .ZN(P1_U3225) );
  NAND2_X1 U8590 ( .A1(n6901), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6897) );
  NAND2_X1 U8591 ( .A1(n6897), .A2(n6896), .ZN(n6899) );
  AOI22_X1 U8592 ( .A1(n7004), .A2(n8442), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n6999), .ZN(n6898) );
  NOR2_X1 U8593 ( .A1(n6899), .A2(n6898), .ZN(n6998) );
  AOI21_X1 U8594 ( .B1(n6899), .B2(n6898), .A(n6998), .ZN(n6909) );
  INV_X1 U8595 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8551) );
  AOI22_X1 U8596 ( .A1(n7004), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n8551), .B2(
        n6999), .ZN(n6903) );
  OAI21_X1 U8597 ( .B1(n6901), .B2(P2_REG1_REG_12__SCAN_IN), .A(n6900), .ZN(
        n6902) );
  NAND2_X1 U8598 ( .A1(n6903), .A2(n6902), .ZN(n7003) );
  OAI21_X1 U8599 ( .B1(n6903), .B2(n6902), .A(n7003), .ZN(n6904) );
  NAND2_X1 U8600 ( .A1(n6904), .A2(n9981), .ZN(n6908) );
  INV_X1 U8601 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6905) );
  NAND2_X1 U8602 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7538) );
  OAI21_X1 U8603 ( .B1(n8157), .B2(n6905), .A(n7538), .ZN(n6906) );
  AOI21_X1 U8604 ( .B1(n8150), .B2(n7004), .A(n6906), .ZN(n6907) );
  OAI211_X1 U8605 ( .C1(n6909), .C2(n8138), .A(n6908), .B(n6907), .ZN(P2_U3258) );
  OR2_X1 U8606 ( .A1(n7313), .A2(n6478), .ZN(n6974) );
  XNOR2_X1 U8607 ( .A(n7263), .B(n7666), .ZN(n6975) );
  XNOR2_X1 U8608 ( .A(n6974), .B(n6975), .ZN(n6972) );
  XNOR2_X1 U8609 ( .A(n6973), .B(n6972), .ZN(n6918) );
  OAI22_X1 U8610 ( .A1(n7414), .A2(n10032), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9659), .ZN(n6916) );
  OAI22_X1 U8611 ( .A1(n6914), .A2(n7806), .B1(n7803), .B2(n7349), .ZN(n6915)
         );
  AOI211_X1 U8612 ( .C1(n7262), .C2(n7794), .A(n6916), .B(n6915), .ZN(n6917)
         );
  OAI21_X1 U8613 ( .B1(n6918), .B2(n7810), .A(n6917), .ZN(P2_U3223) );
  INV_X1 U8614 ( .A(n6919), .ZN(n6922) );
  INV_X1 U8615 ( .A(n6920), .ZN(n6921) );
  NOR3_X1 U8616 ( .A1(n6923), .A2(n6922), .A3(n6921), .ZN(n6925) );
  OAI21_X1 U8617 ( .B1(n6925), .B2(n6924), .A(n8717), .ZN(n6930) );
  NOR2_X1 U8618 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6926), .ZN(n9890) );
  AOI21_X1 U8619 ( .B1(n8708), .B2(n9023), .A(n9890), .ZN(n6927) );
  OAI21_X1 U8620 ( .B1(n7128), .B2(n8720), .A(n6927), .ZN(n6928) );
  AOI21_X1 U8621 ( .B1(n8738), .B2(n7139), .A(n6928), .ZN(n6929) );
  OAI211_X1 U8622 ( .C1(n8736), .C2(n7133), .A(n6930), .B(n6929), .ZN(P1_U3237) );
  XNOR2_X1 U8623 ( .A(n6931), .B(n7847), .ZN(n6997) );
  NAND2_X1 U8624 ( .A1(n6932), .A2(n7897), .ZN(n6933) );
  XNOR2_X1 U8625 ( .A(n6933), .B(n7896), .ZN(n6934) );
  AOI222_X1 U8626 ( .A1(n8434), .A2(n6934), .B1(n8043), .B2(n8343), .C1(n8045), 
        .C2(n8341), .ZN(n6989) );
  INV_X1 U8627 ( .A(n7260), .ZN(n6935) );
  AOI21_X1 U8628 ( .B1(n6937), .B2(n7027), .A(n6935), .ZN(n6994) );
  INV_X2 U8629 ( .A(n6936), .ZN(n8539) );
  AOI22_X1 U8630 ( .A1(n6994), .A2(n8539), .B1(n10045), .B2(n6937), .ZN(n6938)
         );
  OAI211_X1 U8631 ( .C1(n10028), .C2(n6997), .A(n6989), .B(n6938), .ZN(n6940)
         );
  NAND2_X1 U8632 ( .A1(n6940), .A2(n10055), .ZN(n6939) );
  OAI21_X1 U8633 ( .B1(n10055), .B2(n5855), .A(n6939), .ZN(P2_U3472) );
  INV_X1 U8634 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6942) );
  NAND2_X1 U8635 ( .A1(n6940), .A2(n10069), .ZN(n6941) );
  OAI21_X1 U8636 ( .B1(n10069), .B2(n6942), .A(n6941), .ZN(P2_U3527) );
  INV_X1 U8637 ( .A(n6943), .ZN(n6947) );
  NOR2_X1 U8638 ( .A1(n6945), .A2(n6944), .ZN(n6946) );
  NAND2_X1 U8639 ( .A1(n6947), .A2(n6946), .ZN(n7242) );
  NAND2_X1 U8640 ( .A1(n6948), .A2(n9505), .ZN(n6949) );
  AND2_X1 U8641 ( .A1(n6951), .A2(n6950), .ZN(n6952) );
  NAND2_X1 U8642 ( .A1(n7045), .A2(n7060), .ZN(n6953) );
  NAND2_X1 U8643 ( .A1(n7129), .A2(n9934), .ZN(n8914) );
  NAND2_X1 U8644 ( .A1(n6968), .A2(n9023), .ZN(n8913) );
  NAND2_X1 U8645 ( .A1(n6956), .A2(n8870), .ZN(n6957) );
  NAND2_X1 U8646 ( .A1(n7104), .A2(n6957), .ZN(n9933) );
  INV_X1 U8647 ( .A(n6958), .ZN(n8911) );
  XNOR2_X1 U8648 ( .A(n7111), .B(n6955), .ZN(n6961) );
  OAI22_X1 U8649 ( .A1(n7045), .A2(n9798), .B1(n7233), .B2(n9796), .ZN(n6960)
         );
  AOI21_X1 U8650 ( .B1(n6961), .B2(n9768), .A(n6960), .ZN(n9939) );
  INV_X1 U8651 ( .A(n9939), .ZN(n6966) );
  AOI21_X1 U8652 ( .B1(n6962), .B2(n9934), .A(n9963), .ZN(n6963) );
  NAND2_X1 U8653 ( .A1(n6963), .A2(n7135), .ZN(n9937) );
  OAI22_X1 U8654 ( .A1(n9937), .A2(n9161), .B1(n9789), .B2(n6964), .ZN(n6965)
         );
  OAI21_X1 U8655 ( .B1(n6966), .B2(n6965), .A(n9792), .ZN(n6971) );
  INV_X2 U8656 ( .A(n9806), .ZN(n9792) );
  OAI22_X1 U8657 ( .A1(n9792), .A2(n5043), .B1(n9404), .B2(n6968), .ZN(n6969)
         );
  INV_X1 U8658 ( .A(n6969), .ZN(n6970) );
  OAI211_X1 U8659 ( .C1(n9398), .C2(n9933), .A(n6971), .B(n6970), .ZN(P1_U3286) );
  INV_X1 U8660 ( .A(n6974), .ZN(n6976) );
  NAND2_X1 U8661 ( .A1(n6976), .A2(n6975), .ZN(n6977) );
  NAND2_X1 U8662 ( .A1(n6978), .A2(n6977), .ZN(n7395) );
  NOR2_X1 U8663 ( .A1(n7349), .A2(n8539), .ZN(n6979) );
  XNOR2_X1 U8664 ( .A(n8559), .B(n7666), .ZN(n6980) );
  AND2_X1 U8665 ( .A1(n6979), .A2(n6980), .ZN(n7394) );
  INV_X1 U8666 ( .A(n6979), .ZN(n6982) );
  INV_X1 U8667 ( .A(n6980), .ZN(n6981) );
  NAND2_X1 U8668 ( .A1(n6982), .A2(n6981), .ZN(n7393) );
  INV_X1 U8669 ( .A(n7393), .ZN(n6983) );
  NOR2_X1 U8670 ( .A1(n7394), .A2(n6983), .ZN(n6984) );
  XNOR2_X1 U8671 ( .A(n7395), .B(n6984), .ZN(n6988) );
  AOI22_X1 U8672 ( .A1(n7795), .A2(n8043), .B1(n7794), .B2(n7318), .ZN(n6987)
         );
  NAND2_X1 U8673 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8066) );
  OAI21_X1 U8674 ( .B1(n7803), .B2(n7387), .A(n8066), .ZN(n6985) );
  AOI21_X1 U8675 ( .B1(n8559), .B2(n4310), .A(n6985), .ZN(n6986) );
  OAI211_X1 U8676 ( .C1(n6988), .C2(n7810), .A(n6987), .B(n6986), .ZN(P2_U3233) );
  OR2_X1 U8677 ( .A1(n6989), .A2(n8406), .ZN(n6996) );
  OAI22_X1 U8678 ( .A1(n8440), .A2(n6990), .B1(n6704), .B2(n8438), .ZN(n6993)
         );
  NOR2_X1 U8679 ( .A1(n8408), .A2(n6991), .ZN(n6992) );
  AOI211_X1 U8680 ( .C1(n6994), .C2(n8420), .A(n6993), .B(n6992), .ZN(n6995)
         );
  OAI211_X1 U8681 ( .C1(n6997), .C2(n8422), .A(n6996), .B(n6995), .ZN(P2_U3289) );
  AOI21_X1 U8682 ( .B1(n6999), .B2(n8442), .A(n6998), .ZN(n7001) );
  AOI22_X1 U8683 ( .A1(n7419), .A2(n5755), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7002), .ZN(n7000) );
  NOR2_X1 U8684 ( .A1(n7001), .A2(n7000), .ZN(n7420) );
  AOI21_X1 U8685 ( .B1(n7001), .B2(n7000), .A(n7420), .ZN(n7012) );
  AOI22_X1 U8686 ( .A1(n7419), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n4555), .B2(
        n7002), .ZN(n7006) );
  OAI21_X1 U8687 ( .B1(n7004), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7003), .ZN(
        n7005) );
  OAI21_X1 U8688 ( .B1(n7006), .B2(n7005), .A(n7416), .ZN(n7007) );
  NAND2_X1 U8689 ( .A1(n7007), .A2(n9981), .ZN(n7011) );
  INV_X1 U8690 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7008) );
  NAND2_X1 U8691 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7703) );
  OAI21_X1 U8692 ( .B1(n8157), .B2(n7008), .A(n7703), .ZN(n7009) );
  AOI21_X1 U8693 ( .B1(n8150), .B2(n7419), .A(n7009), .ZN(n7010) );
  OAI211_X1 U8694 ( .C1(n7012), .C2(n8138), .A(n7011), .B(n7010), .ZN(P2_U3259) );
  OAI21_X1 U8695 ( .B1(n7014), .B2(n9789), .A(n7013), .ZN(n7015) );
  NAND2_X1 U8696 ( .A1(n7015), .A2(n9792), .ZN(n7021) );
  OR2_X1 U8697 ( .A1(n7017), .A2(n7016), .ZN(n7018) );
  OAI21_X1 U8698 ( .B1(n9787), .B2(n9810), .A(n7019), .ZN(n7020) );
  OAI211_X1 U8699 ( .C1(n4917), .C2(n9792), .A(n7021), .B(n7020), .ZN(P1_U3291) );
  XNOR2_X1 U8700 ( .A(n7022), .B(n7843), .ZN(n10027) );
  OAI21_X1 U8701 ( .B1(n7843), .B2(n7023), .A(n6932), .ZN(n7024) );
  AOI222_X1 U8702 ( .A1(n8434), .A2(n7024), .B1(n8044), .B2(n8343), .C1(n8046), 
        .C2(n8341), .ZN(n10026) );
  MUX2_X1 U8703 ( .A(n7025), .B(n10026), .S(n8438), .Z(n7033) );
  OR2_X1 U8704 ( .A1(n7271), .A2(n7030), .ZN(n7026) );
  AND3_X1 U8705 ( .A1(n7027), .A2(n7026), .A3(n6478), .ZN(n10023) );
  INV_X1 U8706 ( .A(n7028), .ZN(n7029) );
  OAI22_X1 U8707 ( .A1(n8408), .A2(n7030), .B1(n8440), .B2(n7029), .ZN(n7031)
         );
  AOI21_X1 U8708 ( .B1(n10023), .B2(n7324), .A(n7031), .ZN(n7032) );
  OAI211_X1 U8709 ( .C1(n10027), .C2(n8422), .A(n7033), .B(n7032), .ZN(
        P2_U3290) );
  INV_X1 U8710 ( .A(n7034), .ZN(n7037) );
  OAI222_X1 U8711 ( .A1(n7689), .A2(n7035), .B1(n9512), .B2(n7037), .C1(n4515), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  OAI222_X1 U8712 ( .A1(n7365), .A2(n7038), .B1(n8597), .B2(n7037), .C1(n7694), 
        .C2(n7036), .ZN(P2_U3336) );
  OAI21_X1 U8713 ( .B1(n7041), .B2(n7040), .A(n7039), .ZN(n9931) );
  INV_X1 U8714 ( .A(n9931), .ZN(n7059) );
  NAND2_X1 U8715 ( .A1(n4940), .A2(n9161), .ZN(n7042) );
  NOR2_X1 U8716 ( .A1(n9806), .A2(n7042), .ZN(n9788) );
  INV_X1 U8717 ( .A(n9788), .ZN(n7142) );
  OAI21_X1 U8718 ( .B1(n8868), .B2(n7043), .A(n7044), .ZN(n7048) );
  OAI22_X1 U8719 ( .A1(n7046), .A2(n9798), .B1(n7045), .B2(n9796), .ZN(n7047)
         );
  AOI21_X1 U8720 ( .B1(n7048), .B2(n9768), .A(n7047), .ZN(n7049) );
  OAI21_X1 U8721 ( .B1(n7059), .B2(n7117), .A(n7049), .ZN(n9929) );
  NAND2_X1 U8722 ( .A1(n9929), .A2(n9792), .ZN(n7058) );
  NAND2_X1 U8723 ( .A1(n9806), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7050) );
  OAI21_X1 U8724 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(n9789), .A(n7050), .ZN(
        n7055) );
  INV_X1 U8725 ( .A(n9787), .ZN(n9395) );
  OR2_X1 U8726 ( .A1(n7051), .A2(n9927), .ZN(n7052) );
  NAND2_X1 U8727 ( .A1(n7053), .A2(n7052), .ZN(n9928) );
  NOR2_X1 U8728 ( .A1(n9395), .A2(n9928), .ZN(n7054) );
  AOI211_X1 U8729 ( .C1(n9810), .C2(n7056), .A(n7055), .B(n7054), .ZN(n7057)
         );
  OAI211_X1 U8730 ( .C1(n7059), .C2(n7142), .A(n7058), .B(n7057), .ZN(P1_U3288) );
  NOR2_X1 U8731 ( .A1(n9404), .A2(n7060), .ZN(n7064) );
  INV_X1 U8732 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7062) );
  OAI22_X1 U8733 ( .A1(n9792), .A2(n7062), .B1(n7061), .B2(n9789), .ZN(n7063)
         );
  AOI211_X1 U8734 ( .C1(n7065), .C2(n9787), .A(n7064), .B(n7063), .ZN(n7068)
         );
  NAND2_X1 U8735 ( .A1(n7066), .A2(n9788), .ZN(n7067) );
  OAI211_X1 U8736 ( .C1(n7069), .C2(n9806), .A(n7068), .B(n7067), .ZN(P1_U3287) );
  INV_X1 U8737 ( .A(n7070), .ZN(n7078) );
  NOR2_X1 U8738 ( .A1(n9806), .A2(n7117), .ZN(n7071) );
  OR2_X1 U8739 ( .A1(n9788), .A2(n7071), .ZN(n7521) );
  OAI22_X1 U8740 ( .A1(n9792), .A2(n7072), .B1(n9404), .B2(n8969), .ZN(n7077)
         );
  INV_X1 U8741 ( .A(n9789), .ZN(n9316) );
  AOI22_X1 U8742 ( .A1(n7073), .A2(n9001), .B1(n9316), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7074) );
  AOI21_X1 U8743 ( .B1(n7075), .B2(n7074), .A(n9806), .ZN(n7076) );
  AOI211_X1 U8744 ( .C1(n7078), .C2(n7521), .A(n7077), .B(n7076), .ZN(n7079)
         );
  INV_X1 U8745 ( .A(n7079), .ZN(P1_U3290) );
  INV_X1 U8746 ( .A(n7080), .ZN(n7081) );
  NAND2_X1 U8747 ( .A1(n8438), .A2(n7081), .ZN(n8453) );
  INV_X1 U8748 ( .A(n8453), .ZN(n7267) );
  NOR2_X1 U8749 ( .A1(n8440), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7083) );
  NOR2_X1 U8750 ( .A1(n8438), .A2(n6637), .ZN(n7082) );
  AOI211_X1 U8751 ( .C1(n7084), .C2(n7324), .A(n7083), .B(n7082), .ZN(n7085)
         );
  OAI21_X1 U8752 ( .B1(n7086), .B2(n8408), .A(n7085), .ZN(n7087) );
  AOI21_X1 U8753 ( .B1(n7267), .B2(n7088), .A(n7087), .ZN(n7089) );
  OAI21_X1 U8754 ( .B1(n7090), .B2(n8406), .A(n7089), .ZN(P2_U3293) );
  NAND2_X1 U8755 ( .A1(n7092), .A2(n7091), .ZN(n7094) );
  XNOR2_X1 U8756 ( .A(n7094), .B(n7093), .ZN(n7101) );
  INV_X1 U8757 ( .A(n7294), .ZN(n9955) );
  NOR2_X1 U8758 ( .A1(n8726), .A2(n9955), .ZN(n7100) );
  INV_X1 U8759 ( .A(n9019), .ZN(n7378) );
  INV_X1 U8760 ( .A(n7128), .ZN(n9021) );
  NOR2_X1 U8761 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7095), .ZN(n9903) );
  AOI21_X1 U8762 ( .B1(n8708), .B2(n9021), .A(n9903), .ZN(n7098) );
  INV_X1 U8763 ( .A(n7118), .ZN(n7096) );
  NAND2_X1 U8764 ( .A1(n8723), .A2(n7096), .ZN(n7097) );
  OAI211_X1 U8765 ( .C1(n7378), .C2(n8720), .A(n7098), .B(n7097), .ZN(n7099)
         );
  AOI211_X1 U8766 ( .C1(n7101), .C2(n8717), .A(n7100), .B(n7099), .ZN(n7102)
         );
  INV_X1 U8767 ( .A(n7102), .ZN(P1_U3219) );
  NAND2_X1 U8768 ( .A1(n9023), .A2(n9934), .ZN(n7103) );
  NAND2_X1 U8769 ( .A1(n7233), .A2(n7139), .ZN(n8915) );
  INV_X1 U8770 ( .A(n7139), .ZN(n9942) );
  INV_X1 U8771 ( .A(n7233), .ZN(n9022) );
  NAND2_X1 U8772 ( .A1(n9942), .A2(n9022), .ZN(n8967) );
  NAND2_X1 U8773 ( .A1(n7233), .A2(n9942), .ZN(n7106) );
  NAND2_X1 U8774 ( .A1(n7128), .A2(n7246), .ZN(n8918) );
  NAND2_X1 U8775 ( .A1(n8918), .A2(n8974), .ZN(n7238) );
  NAND2_X1 U8776 ( .A1(n7128), .A2(n9949), .ZN(n7107) );
  NAND2_X1 U8777 ( .A1(n7287), .A2(n7294), .ZN(n8919) );
  NAND2_X1 U8778 ( .A1(n9955), .A2(n9020), .ZN(n8758) );
  INV_X1 U8779 ( .A(n8875), .ZN(n7108) );
  NAND2_X1 U8780 ( .A1(n7109), .A2(n8875), .ZN(n7110) );
  NAND2_X1 U8781 ( .A1(n7296), .A2(n7110), .ZN(n9954) );
  INV_X1 U8782 ( .A(n8967), .ZN(n7112) );
  NAND2_X1 U8783 ( .A1(n8964), .A2(n8874), .ZN(n7113) );
  XNOR2_X1 U8784 ( .A(n7284), .B(n8875), .ZN(n7115) );
  OAI22_X1 U8785 ( .A1(n7128), .A2(n9798), .B1(n7378), .B2(n9796), .ZN(n7114)
         );
  AOI21_X1 U8786 ( .B1(n7115), .B2(n9768), .A(n7114), .ZN(n7116) );
  OAI21_X1 U8787 ( .B1(n9954), .B2(n7117), .A(n7116), .ZN(n9957) );
  NAND2_X1 U8788 ( .A1(n9957), .A2(n9792), .ZN(n7124) );
  OAI22_X1 U8789 ( .A1(n9792), .A2(n7119), .B1(n7118), .B2(n9789), .ZN(n7122)
         );
  NAND2_X1 U8790 ( .A1(n7240), .A2(n7294), .ZN(n7120) );
  NAND2_X1 U8791 ( .A1(n7290), .A2(n7120), .ZN(n9956) );
  NOR2_X1 U8792 ( .A1(n9956), .A2(n9395), .ZN(n7121) );
  AOI211_X1 U8793 ( .C1(n9810), .C2(n7294), .A(n7122), .B(n7121), .ZN(n7123)
         );
  OAI211_X1 U8794 ( .C1(n9954), .C2(n7142), .A(n7124), .B(n7123), .ZN(P1_U3283) );
  OAI21_X1 U8795 ( .B1(n4387), .B2(n7105), .A(n7125), .ZN(n9946) );
  INV_X1 U8796 ( .A(n9946), .ZN(n7143) );
  XNOR2_X1 U8797 ( .A(n7126), .B(n7127), .ZN(n7132) );
  OAI22_X1 U8798 ( .A1(n7129), .A2(n9798), .B1(n7128), .B2(n9796), .ZN(n7130)
         );
  AOI21_X1 U8799 ( .B1(n9946), .B2(n9805), .A(n7130), .ZN(n7131) );
  OAI21_X1 U8800 ( .B1(n9802), .B2(n7132), .A(n7131), .ZN(n9944) );
  NAND2_X1 U8801 ( .A1(n9944), .A2(n9792), .ZN(n7141) );
  OAI22_X1 U8802 ( .A1(n9792), .A2(n7134), .B1(n7133), .B2(n9789), .ZN(n7138)
         );
  AND2_X1 U8803 ( .A1(n7135), .A2(n7139), .ZN(n7136) );
  OR2_X1 U8804 ( .A1(n7136), .A2(n7241), .ZN(n9943) );
  NOR2_X1 U8805 ( .A1(n9943), .A2(n9395), .ZN(n7137) );
  AOI211_X1 U8806 ( .C1(n9810), .C2(n7139), .A(n7138), .B(n7137), .ZN(n7140)
         );
  OAI211_X1 U8807 ( .C1(n7143), .C2(n7142), .A(n7141), .B(n7140), .ZN(P1_U3285) );
  INV_X1 U8808 ( .A(n7207), .ZN(n7146) );
  AOI21_X1 U8809 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8594), .A(n7144), .ZN(
        n7145) );
  OAI21_X1 U8810 ( .B1(n7146), .B2(n7545), .A(n7145), .ZN(P2_U3335) );
  INV_X1 U8811 ( .A(n7871), .ZN(n7148) );
  OAI21_X1 U8812 ( .B1(n7148), .B2(n7147), .A(n7839), .ZN(n7150) );
  NAND2_X1 U8813 ( .A1(n7150), .A2(n7149), .ZN(n7151) );
  AOI222_X1 U8814 ( .A1(n8434), .A2(n7151), .B1(n6674), .B2(n8343), .C1(n6673), 
        .C2(n8341), .ZN(n10008) );
  OAI22_X1 U8815 ( .A1(n8440), .A2(n7152), .B1(n6620), .B2(n8438), .ZN(n7156)
         );
  INV_X1 U8816 ( .A(n7324), .ZN(n7213) );
  OAI211_X1 U8817 ( .C1(n7154), .C2(n10009), .A(n7153), .B(n8539), .ZN(n10007)
         );
  NOR2_X1 U8818 ( .A1(n7213), .A2(n10007), .ZN(n7155) );
  AOI211_X1 U8819 ( .C1(n8450), .C2(n7157), .A(n7156), .B(n7155), .ZN(n7161)
         );
  OAI21_X1 U8820 ( .B1(n7159), .B2(n7839), .A(n7158), .ZN(n10011) );
  INV_X1 U8821 ( .A(n8422), .ZN(n8265) );
  NAND2_X1 U8822 ( .A1(n10011), .A2(n8265), .ZN(n7160) );
  OAI211_X1 U8823 ( .C1(n10008), .C2(n8406), .A(n7161), .B(n7160), .ZN(
        P2_U3294) );
  NAND2_X1 U8824 ( .A1(n6769), .A2(n7882), .ZN(n7163) );
  INV_X1 U8825 ( .A(n7840), .ZN(n7162) );
  XNOR2_X1 U8826 ( .A(n7163), .B(n7162), .ZN(n7164) );
  NAND2_X1 U8827 ( .A1(n7164), .A2(n8434), .ZN(n7169) );
  OAI22_X1 U8828 ( .A1(n7166), .A2(n8430), .B1(n7165), .B2(n6188), .ZN(n7167)
         );
  INV_X1 U8829 ( .A(n7167), .ZN(n7168) );
  NAND2_X1 U8830 ( .A1(n7169), .A2(n7168), .ZN(n10015) );
  INV_X1 U8831 ( .A(n10015), .ZN(n7181) );
  OAI22_X1 U8832 ( .A1(n8440), .A2(n7170), .B1(n6639), .B2(n8438), .ZN(n7175)
         );
  INV_X1 U8833 ( .A(n7171), .ZN(n7173) );
  INV_X1 U8834 ( .A(n7273), .ZN(n7172) );
  OAI211_X1 U8835 ( .C1(n10014), .C2(n7173), .A(n7172), .B(n8539), .ZN(n10013)
         );
  NOR2_X1 U8836 ( .A1(n10013), .A2(n7213), .ZN(n7174) );
  AOI211_X1 U8837 ( .C1(n8450), .C2(n7176), .A(n7175), .B(n7174), .ZN(n7180)
         );
  OAI21_X1 U8838 ( .B1(n7177), .B2(n7840), .A(n7178), .ZN(n10017) );
  NAND2_X1 U8839 ( .A1(n10017), .A2(n8265), .ZN(n7179) );
  OAI211_X1 U8840 ( .C1(n7181), .C2(n8406), .A(n7180), .B(n7179), .ZN(P2_U3292) );
  INV_X1 U8841 ( .A(n10001), .ZN(n7182) );
  NAND2_X1 U8842 ( .A1(n7183), .A2(n7182), .ZN(n7868) );
  NAND2_X1 U8843 ( .A1(n7184), .A2(n7868), .ZN(n10003) );
  INV_X1 U8844 ( .A(n10003), .ZN(n7189) );
  AOI22_X1 U8845 ( .A1(n10003), .A2(n8434), .B1(n8343), .B2(n6673), .ZN(n10005) );
  NAND2_X1 U8846 ( .A1(n8404), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7185) );
  AOI21_X1 U8847 ( .B1(n10005), .B2(n7185), .A(n8406), .ZN(n7186) );
  AOI21_X1 U8848 ( .B1(n8406), .B2(P2_REG2_REG_0__SCAN_IN), .A(n7186), .ZN(
        n7188) );
  OAI21_X1 U8849 ( .B1(n8420), .B2(n8450), .A(n10001), .ZN(n7187) );
  OAI211_X1 U8850 ( .C1(n7189), .C2(n8422), .A(n7188), .B(n7187), .ZN(P2_U3296) );
  INV_X1 U8851 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7205) );
  OR2_X1 U8852 ( .A1(n7439), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7191) );
  NAND2_X1 U8853 ( .A1(n7439), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7190) );
  AND2_X1 U8854 ( .A1(n7191), .A2(n7190), .ZN(n7195) );
  NAND2_X1 U8855 ( .A1(n7193), .A2(n7192), .ZN(n7194) );
  NAND2_X1 U8856 ( .A1(n7195), .A2(n7194), .ZN(n7438) );
  OAI21_X1 U8857 ( .B1(n7195), .B2(n7194), .A(n7438), .ZN(n7196) );
  NAND2_X1 U8858 ( .A1(n9920), .A2(n7196), .ZN(n7197) );
  NAND2_X1 U8859 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7572) );
  NAND2_X1 U8860 ( .A1(n7197), .A2(n7572), .ZN(n7203) );
  INV_X1 U8861 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7200) );
  AOI211_X1 U8862 ( .C1(n7201), .C2(n7200), .A(n7434), .B(n9885), .ZN(n7202)
         );
  AOI211_X1 U8863 ( .C1(n9912), .C2(n7439), .A(n7203), .B(n7202), .ZN(n7204)
         );
  OAI21_X1 U8864 ( .B1(n9925), .B2(n7205), .A(n7204), .ZN(P1_U3255) );
  NAND2_X1 U8865 ( .A1(n7207), .A2(n7206), .ZN(n7209) );
  NAND2_X1 U8866 ( .A1(n7208), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9010) );
  OAI211_X1 U8867 ( .C1(n7210), .C2(n7689), .A(n7209), .B(n9010), .ZN(P1_U3330) );
  INV_X1 U8868 ( .A(n7211), .ZN(n7214) );
  INV_X1 U8869 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7212) );
  OAI22_X1 U8870 ( .A1(n7214), .A2(n7213), .B1(n7212), .B2(n8440), .ZN(n7215)
         );
  AOI21_X1 U8871 ( .B1(n8406), .B2(P2_REG2_REG_1__SCAN_IN), .A(n7215), .ZN(
        n7220) );
  INV_X1 U8872 ( .A(n7216), .ZN(n7218) );
  AOI22_X1 U8873 ( .A1(n7218), .A2(n8438), .B1(n8450), .B2(n7217), .ZN(n7219)
         );
  OAI211_X1 U8874 ( .C1(n7221), .C2(n8422), .A(n7220), .B(n7219), .ZN(P2_U3295) );
  INV_X1 U8875 ( .A(n7222), .ZN(n7223) );
  AOI21_X1 U8876 ( .B1(n7225), .B2(n7224), .A(n7223), .ZN(n7231) );
  NOR2_X1 U8877 ( .A1(n8732), .A2(n7287), .ZN(n7226) );
  AOI211_X1 U8878 ( .C1(n8734), .C2(n9018), .A(n7227), .B(n7226), .ZN(n7228)
         );
  OAI21_X1 U8879 ( .B1(n8736), .B2(n7288), .A(n7228), .ZN(n7229) );
  AOI21_X1 U8880 ( .B1(n8738), .B2(n7335), .A(n7229), .ZN(n7230) );
  OAI21_X1 U8881 ( .B1(n7231), .B2(n8740), .A(n7230), .ZN(P1_U3229) );
  XNOR2_X1 U8882 ( .A(n8964), .B(n8874), .ZN(n7232) );
  NAND2_X1 U8883 ( .A1(n7232), .A2(n9768), .ZN(n7236) );
  OAI22_X1 U8884 ( .A1(n7233), .A2(n9798), .B1(n7287), .B2(n9796), .ZN(n7234)
         );
  INV_X1 U8885 ( .A(n7234), .ZN(n7235) );
  NAND2_X1 U8886 ( .A1(n7236), .A2(n7235), .ZN(n9950) );
  INV_X1 U8887 ( .A(n9950), .ZN(n7250) );
  OAI21_X1 U8888 ( .B1(n7239), .B2(n7238), .A(n7237), .ZN(n9952) );
  INV_X1 U8889 ( .A(n9398), .ZN(n9337) );
  OAI211_X1 U8890 ( .C1(n7241), .C2(n9949), .A(n7240), .B(n9816), .ZN(n9948)
         );
  NOR2_X1 U8891 ( .A1(n7242), .A2(n9161), .ZN(n9371) );
  INV_X1 U8892 ( .A(n9371), .ZN(n7525) );
  OAI22_X1 U8893 ( .A1(n9792), .A2(n7244), .B1(n7243), .B2(n9789), .ZN(n7245)
         );
  AOI21_X1 U8894 ( .B1(n9810), .B2(n7246), .A(n7245), .ZN(n7247) );
  OAI21_X1 U8895 ( .B1(n9948), .B2(n7525), .A(n7247), .ZN(n7248) );
  AOI21_X1 U8896 ( .B1(n9952), .B2(n9337), .A(n7248), .ZN(n7249) );
  OAI21_X1 U8897 ( .B1(n9806), .B2(n7250), .A(n7249), .ZN(P1_U3284) );
  INV_X1 U8898 ( .A(n7251), .ZN(n7252) );
  AOI21_X1 U8899 ( .B1(n5878), .B2(n7253), .A(n7252), .ZN(n7259) );
  NAND2_X1 U8900 ( .A1(n7254), .A2(n7901), .ZN(n7255) );
  INV_X1 U8901 ( .A(n8427), .ZN(n7316) );
  NAND2_X1 U8902 ( .A1(n10036), .A2(n7316), .ZN(n7258) );
  AOI22_X1 U8903 ( .A1(n8341), .A2(n8044), .B1(n8042), .B2(n8343), .ZN(n7257)
         );
  OAI211_X1 U8904 ( .C1(n8410), .C2(n7259), .A(n7258), .B(n7257), .ZN(n10034)
         );
  INV_X1 U8905 ( .A(n10034), .ZN(n7269) );
  NAND2_X1 U8906 ( .A1(n7260), .A2(n7263), .ZN(n7261) );
  NAND2_X1 U8907 ( .A1(n7317), .A2(n7261), .ZN(n10033) );
  INV_X1 U8908 ( .A(n8420), .ZN(n8446) );
  AOI22_X1 U8909 ( .A1(n8406), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n7262), .B2(
        n8404), .ZN(n7265) );
  NAND2_X1 U8910 ( .A1(n8450), .A2(n7263), .ZN(n7264) );
  OAI211_X1 U8911 ( .C1(n10033), .C2(n8446), .A(n7265), .B(n7264), .ZN(n7266)
         );
  AOI21_X1 U8912 ( .B1(n10036), .B2(n7267), .A(n7266), .ZN(n7268) );
  OAI21_X1 U8913 ( .B1(n7269), .B2(n8406), .A(n7268), .ZN(P2_U3288) );
  XNOR2_X1 U8914 ( .A(n7270), .B(n7838), .ZN(n10022) );
  INV_X1 U8915 ( .A(n7271), .ZN(n7272) );
  OAI211_X1 U8916 ( .C1(n10019), .C2(n7273), .A(n7272), .B(n8539), .ZN(n10018)
         );
  AND2_X1 U8917 ( .A1(n8438), .A2(n7833), .ZN(n8358) );
  INV_X1 U8918 ( .A(n8358), .ZN(n7277) );
  AOI22_X1 U8919 ( .A1(n8450), .A2(n7275), .B1(n8404), .B2(n7274), .ZN(n7276)
         );
  OAI21_X1 U8920 ( .B1(n10018), .B2(n7277), .A(n7276), .ZN(n7282) );
  XOR2_X1 U8921 ( .A(n7278), .B(n7838), .Z(n7280) );
  OAI21_X1 U8922 ( .B1(n7280), .B2(n8410), .A(n7279), .ZN(n10020) );
  MUX2_X1 U8923 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10020), .S(n8438), .Z(n7281)
         );
  AOI211_X1 U8924 ( .C1(n8265), .C2(n10022), .A(n7282), .B(n7281), .ZN(n7283)
         );
  INV_X1 U8925 ( .A(n7283), .ZN(P2_U3291) );
  NAND2_X1 U8926 ( .A1(n7329), .A2(n8758), .ZN(n7285) );
  OR2_X1 U8927 ( .A1(n7378), .A2(n7335), .ZN(n8762) );
  NAND2_X1 U8928 ( .A1(n7335), .A2(n7378), .ZN(n8759) );
  XNOR2_X1 U8929 ( .A(n7285), .B(n8876), .ZN(n7286) );
  OAI222_X1 U8930 ( .A1(n9796), .A2(n9799), .B1(n9798), .B2(n7287), .C1(n9802), 
        .C2(n7286), .ZN(n9965) );
  INV_X1 U8931 ( .A(n9965), .ZN(n7299) );
  INV_X1 U8932 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7289) );
  OAI22_X1 U8933 ( .A1(n9792), .A2(n7289), .B1(n7288), .B2(n9789), .ZN(n7293)
         );
  INV_X1 U8934 ( .A(n7335), .ZN(n9962) );
  INV_X1 U8935 ( .A(n7290), .ZN(n7291) );
  INV_X1 U8936 ( .A(n7338), .ZN(n7339) );
  OAI21_X1 U8937 ( .B1(n9962), .B2(n7291), .A(n7339), .ZN(n9964) );
  NOR2_X1 U8938 ( .A1(n9964), .A2(n9395), .ZN(n7292) );
  AOI211_X1 U8939 ( .C1(n9810), .C2(n7335), .A(n7293), .B(n7292), .ZN(n7298)
         );
  NAND2_X1 U8940 ( .A1(n7294), .A2(n9020), .ZN(n7295) );
  NAND2_X1 U8941 ( .A1(n7296), .A2(n7295), .ZN(n7337) );
  XNOR2_X1 U8942 ( .A(n7337), .B(n8876), .ZN(n9968) );
  NAND2_X1 U8943 ( .A1(n9968), .A2(n7521), .ZN(n7297) );
  OAI211_X1 U8944 ( .C1(n7299), .C2(n9806), .A(n7298), .B(n7297), .ZN(P1_U3282) );
  XNOR2_X1 U8945 ( .A(n7300), .B(n7301), .ZN(n8557) );
  INV_X1 U8946 ( .A(n7301), .ZN(n7851) );
  XNOR2_X1 U8947 ( .A(n7302), .B(n7851), .ZN(n7303) );
  AOI22_X1 U8948 ( .A1(n8341), .A2(n4587), .B1(n8040), .B2(n8343), .ZN(n7408)
         );
  OAI21_X1 U8949 ( .B1(n7303), .B2(n8410), .A(n7408), .ZN(n8553) );
  INV_X1 U8950 ( .A(n8555), .ZN(n7415) );
  INV_X1 U8951 ( .A(n7460), .ZN(n7304) );
  AOI211_X1 U8952 ( .C1(n8555), .C2(n7357), .A(n10050), .B(n7304), .ZN(n8554)
         );
  NAND2_X1 U8953 ( .A1(n8554), .A2(n7324), .ZN(n7306) );
  AOI22_X1 U8954 ( .A1(n8406), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7411), .B2(
        n8404), .ZN(n7305) );
  OAI211_X1 U8955 ( .C1(n7415), .C2(n8408), .A(n7306), .B(n7305), .ZN(n7307)
         );
  AOI21_X1 U8956 ( .B1(n8438), .B2(n8553), .A(n7307), .ZN(n7308) );
  OAI21_X1 U8957 ( .B1(n8557), .B2(n8422), .A(n7308), .ZN(P2_U3285) );
  OAI21_X1 U8958 ( .B1(n7310), .B2(n5895), .A(n7309), .ZN(n7321) );
  NAND3_X1 U8959 ( .A1(n7251), .A2(n5895), .A3(n7905), .ZN(n7312) );
  AOI21_X1 U8960 ( .B1(n7311), .B2(n7312), .A(n8410), .ZN(n7315) );
  OAI22_X1 U8961 ( .A1(n7313), .A2(n6188), .B1(n7387), .B2(n8430), .ZN(n7314)
         );
  AOI211_X1 U8962 ( .C1(n7321), .C2(n7316), .A(n7315), .B(n7314), .ZN(n8561)
         );
  AOI211_X1 U8963 ( .C1(n8559), .C2(n7317), .A(n10050), .B(n7355), .ZN(n8558)
         );
  AOI22_X1 U8964 ( .A1(n8406), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7318), .B2(
        n8404), .ZN(n7319) );
  OAI21_X1 U8965 ( .B1(n7320), .B2(n8408), .A(n7319), .ZN(n7323) );
  INV_X1 U8966 ( .A(n7321), .ZN(n8562) );
  NOR2_X1 U8967 ( .A1(n8562), .A2(n8453), .ZN(n7322) );
  AOI211_X1 U8968 ( .C1(n8558), .C2(n7324), .A(n7323), .B(n7322), .ZN(n7325)
         );
  OAI21_X1 U8969 ( .B1(n8406), .B2(n8561), .A(n7325), .ZN(P2_U3287) );
  NAND2_X1 U8970 ( .A1(n9735), .A2(n9799), .ZN(n8753) );
  NAND2_X1 U8971 ( .A1(n8897), .A2(n8753), .ZN(n8878) );
  INV_X1 U8972 ( .A(n8878), .ZN(n7332) );
  NAND2_X1 U8973 ( .A1(n8762), .A2(n8758), .ZN(n7328) );
  INV_X1 U8974 ( .A(n7328), .ZN(n7327) );
  INV_X1 U8975 ( .A(n8759), .ZN(n7326) );
  AOI21_X1 U8976 ( .B1(n7329), .B2(n7327), .A(n7326), .ZN(n7331) );
  NAND2_X1 U8977 ( .A1(n8920), .A2(n7328), .ZN(n8898) );
  NAND2_X1 U8978 ( .A1(n7513), .A2(n8897), .ZN(n7330) );
  OAI211_X1 U8979 ( .C1(n7332), .C2(n7331), .A(n7330), .B(n9768), .ZN(n7334)
         );
  AOI22_X1 U8980 ( .A1(n9771), .A2(n9017), .B1(n9019), .B2(n9772), .ZN(n7333)
         );
  AND2_X1 U8981 ( .A1(n7334), .A2(n7333), .ZN(n9737) );
  AND2_X1 U8982 ( .A1(n7335), .A2(n9019), .ZN(n7336) );
  OAI22_X1 U8983 ( .A1(n7337), .A2(n7336), .B1(n7335), .B2(n9019), .ZN(n7518)
         );
  XOR2_X1 U8984 ( .A(n7518), .B(n8878), .Z(n9738) );
  INV_X1 U8985 ( .A(n9738), .ZN(n9740) );
  NAND2_X1 U8986 ( .A1(n9740), .A2(n7521), .ZN(n7344) );
  INV_X1 U8987 ( .A(n9735), .ZN(n7372) );
  AOI211_X1 U8988 ( .C1(n9735), .C2(n7339), .A(n9963), .B(n9783), .ZN(n9734)
         );
  NOR2_X1 U8989 ( .A1(n9404), .A2(n7372), .ZN(n7342) );
  OAI22_X1 U8990 ( .A1(n9792), .A2(n7340), .B1(n7374), .B2(n9789), .ZN(n7341)
         );
  AOI211_X1 U8991 ( .C1(n9734), .C2(n9371), .A(n7342), .B(n7341), .ZN(n7343)
         );
  OAI211_X1 U8992 ( .C1(n9806), .C2(n9737), .A(n7344), .B(n7343), .ZN(P1_U3281) );
  OAI21_X1 U8993 ( .B1(n7346), .B2(n7347), .A(n7345), .ZN(n10037) );
  NAND2_X1 U8994 ( .A1(n7311), .A2(n7907), .ZN(n7348) );
  INV_X1 U8995 ( .A(n7347), .ZN(n7850) );
  XNOR2_X1 U8996 ( .A(n7348), .B(n7850), .ZN(n7351) );
  OAI22_X1 U8997 ( .A1(n7349), .A2(n6188), .B1(n7467), .B2(n8430), .ZN(n7350)
         );
  AOI21_X1 U8998 ( .B1(n7351), .B2(n8434), .A(n7350), .ZN(n7352) );
  OAI21_X1 U8999 ( .B1(n10037), .B2(n8427), .A(n7352), .ZN(n10041) );
  NAND2_X1 U9000 ( .A1(n10041), .A2(n8438), .ZN(n7361) );
  INV_X1 U9001 ( .A(n7399), .ZN(n7353) );
  OAI22_X1 U9002 ( .A1(n8438), .A2(n7354), .B1(n7353), .B2(n8440), .ZN(n7359)
         );
  OR2_X1 U9003 ( .A1(n7355), .A2(n10039), .ZN(n7356) );
  NAND2_X1 U9004 ( .A1(n7357), .A2(n7356), .ZN(n10040) );
  NOR2_X1 U9005 ( .A1(n10040), .A2(n8446), .ZN(n7358) );
  AOI211_X1 U9006 ( .C1(n8450), .C2(n7386), .A(n7359), .B(n7358), .ZN(n7360)
         );
  OAI211_X1 U9007 ( .C1(n10037), .C2(n8453), .A(n7361), .B(n7360), .ZN(
        P2_U3286) );
  INV_X1 U9008 ( .A(n7362), .ZN(n7367) );
  OAI222_X1 U9009 ( .A1(n9512), .A2(n7367), .B1(P1_U3084), .B2(n7364), .C1(
        n7363), .C2(n7689), .ZN(P1_U3329) );
  INV_X1 U9010 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7366) );
  OAI222_X1 U9011 ( .A1(n7694), .A2(n7368), .B1(n8597), .B2(n7367), .C1(n7366), 
        .C2(n7365), .ZN(P2_U3334) );
  OAI21_X1 U9012 ( .B1(n7371), .B2(n7370), .A(n7369), .ZN(n7381) );
  NOR2_X1 U9013 ( .A1(n7372), .A2(n8726), .ZN(n7380) );
  AOI21_X1 U9014 ( .B1(n8734), .B2(n9017), .A(n7373), .ZN(n7377) );
  INV_X1 U9015 ( .A(n7374), .ZN(n7375) );
  NAND2_X1 U9016 ( .A1(n8723), .A2(n7375), .ZN(n7376) );
  OAI211_X1 U9017 ( .C1(n7378), .C2(n8732), .A(n7377), .B(n7376), .ZN(n7379)
         );
  AOI211_X1 U9018 ( .C1(n7381), .C2(n8717), .A(n7380), .B(n7379), .ZN(n7382)
         );
  INV_X1 U9019 ( .A(n7382), .ZN(P1_U3215) );
  INV_X1 U9020 ( .A(n7383), .ZN(n7430) );
  AOI22_X1 U9021 ( .A1(n7384), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n8594), .ZN(n7385) );
  OAI21_X1 U9022 ( .B1(n7430), .B2(n7545), .A(n7385), .ZN(P2_U3333) );
  XNOR2_X1 U9023 ( .A(n7386), .B(n7666), .ZN(n7388) );
  NOR2_X1 U9024 ( .A1(n7387), .A2(n8539), .ZN(n7389) );
  NAND2_X1 U9025 ( .A1(n7388), .A2(n7389), .ZN(n7404) );
  INV_X1 U9026 ( .A(n7388), .ZN(n7391) );
  INV_X1 U9027 ( .A(n7389), .ZN(n7390) );
  NAND2_X1 U9028 ( .A1(n7391), .A2(n7390), .ZN(n7392) );
  NAND2_X1 U9029 ( .A1(n7404), .A2(n7392), .ZN(n7398) );
  AOI211_X1 U9030 ( .C1(n7398), .C2(n7397), .A(n7810), .B(n4385), .ZN(n7403)
         );
  AOI22_X1 U9031 ( .A1(n7795), .A2(n8042), .B1(n7794), .B2(n7399), .ZN(n7401)
         );
  AOI22_X1 U9032 ( .A1(n7793), .A2(n8041), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n7400) );
  OAI211_X1 U9033 ( .C1(n10039), .C2(n7414), .A(n7401), .B(n7400), .ZN(n7402)
         );
  OR2_X1 U9034 ( .A1(n7403), .A2(n7402), .ZN(P2_U3219) );
  XNOR2_X1 U9035 ( .A(n8555), .B(n7666), .ZN(n7489) );
  NAND2_X1 U9036 ( .A1(n8041), .A2(n10050), .ZN(n7487) );
  XNOR2_X1 U9037 ( .A(n7489), .B(n7487), .ZN(n7405) );
  NAND2_X1 U9038 ( .A1(n7406), .A2(n7405), .ZN(n7491) );
  OAI211_X1 U9039 ( .C1(n7406), .C2(n7405), .A(n7491), .B(n7789), .ZN(n7413)
         );
  OAI22_X1 U9040 ( .A1(n7409), .A2(n7408), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7407), .ZN(n7410) );
  AOI21_X1 U9041 ( .B1(n7411), .B2(n7794), .A(n7410), .ZN(n7412) );
  OAI211_X1 U9042 ( .C1(n7415), .C2(n7414), .A(n7413), .B(n7412), .ZN(P2_U3238) );
  INV_X1 U9043 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7417) );
  AOI211_X1 U9044 ( .C1(n7418), .C2(n7417), .A(n8091), .B(n9983), .ZN(n7428)
         );
  NOR2_X1 U9045 ( .A1(n7419), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7421) );
  NOR2_X1 U9046 ( .A1(n7421), .A2(n7420), .ZN(n8099) );
  XNOR2_X1 U9047 ( .A(n8099), .B(n8100), .ZN(n7422) );
  NOR2_X1 U9048 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7422), .ZN(n8101) );
  AOI21_X1 U9049 ( .B1(n7422), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8101), .ZN(
        n7426) );
  NOR2_X1 U9050 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5939), .ZN(n7423) );
  AOI21_X1 U9051 ( .B1(n9987), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7423), .ZN(
        n7425) );
  NAND2_X1 U9052 ( .A1(n8150), .A2(n8100), .ZN(n7424) );
  OAI211_X1 U9053 ( .C1(n7426), .C2(n8138), .A(n7425), .B(n7424), .ZN(n7427)
         );
  OR2_X1 U9054 ( .A1(n7428), .A2(n7427), .ZN(P2_U3260) );
  OAI222_X1 U9055 ( .A1(n7689), .A2(n7431), .B1(n9512), .B2(n7430), .C1(n7429), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U9056 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7446) );
  NOR2_X1 U9057 ( .A1(n7433), .A2(n7432), .ZN(n7435) );
  AOI211_X1 U9058 ( .C1(n7436), .C2(n9391), .A(n9044), .B(n9885), .ZN(n7437)
         );
  INV_X1 U9059 ( .A(n7437), .ZN(n7445) );
  NAND2_X1 U9060 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8731) );
  INV_X1 U9061 ( .A(n8731), .ZN(n7442) );
  OAI21_X1 U9062 ( .B1(n7439), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7438), .ZN(
        n9048) );
  XNOR2_X1 U9063 ( .A(n9049), .B(n9048), .ZN(n7440) );
  INV_X1 U9064 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9823) );
  NOR2_X1 U9065 ( .A1(n9823), .A2(n7440), .ZN(n9050) );
  AOI211_X1 U9066 ( .C1(n7440), .C2(n9823), .A(n9050), .B(n9898), .ZN(n7441)
         );
  AOI211_X1 U9067 ( .C1(n9912), .C2(n7443), .A(n7442), .B(n7441), .ZN(n7444)
         );
  OAI211_X1 U9068 ( .C1(n9925), .C2(n7446), .A(n7445), .B(n7444), .ZN(P1_U3256) );
  INV_X1 U9069 ( .A(n7548), .ZN(n9832) );
  INV_X1 U9070 ( .A(n7447), .ZN(n7451) );
  AOI21_X1 U9071 ( .B1(n7502), .B2(n7449), .A(n7448), .ZN(n7450) );
  OAI21_X1 U9072 ( .B1(n7451), .B2(n7450), .A(n8717), .ZN(n7458) );
  INV_X1 U9073 ( .A(n7522), .ZN(n7456) );
  INV_X1 U9074 ( .A(n9016), .ZN(n8771) );
  INV_X1 U9075 ( .A(n7452), .ZN(n7453) );
  AOI21_X1 U9076 ( .B1(n8708), .B2(n9017), .A(n7453), .ZN(n7454) );
  OAI21_X1 U9077 ( .B1(n8771), .B2(n8720), .A(n7454), .ZN(n7455) );
  AOI21_X1 U9078 ( .B1(n7456), .B2(n8723), .A(n7455), .ZN(n7457) );
  OAI211_X1 U9079 ( .C1(n9832), .C2(n8726), .A(n7458), .B(n7457), .ZN(P1_U3222) );
  XNOR2_X1 U9080 ( .A(n7459), .B(n7854), .ZN(n10053) );
  NAND2_X1 U9081 ( .A1(n7460), .A2(n10046), .ZN(n7461) );
  NAND2_X1 U9082 ( .A1(n4598), .A2(n7461), .ZN(n10049) );
  INV_X1 U9083 ( .A(n7493), .ZN(n7462) );
  OAI22_X1 U9084 ( .A1(n8438), .A2(n7463), .B1(n7462), .B2(n8440), .ZN(n7464)
         );
  AOI21_X1 U9085 ( .B1(n8450), .B2(n10046), .A(n7464), .ZN(n7465) );
  OAI21_X1 U9086 ( .B1(n10049), .B2(n8446), .A(n7465), .ZN(n7471) );
  XNOR2_X1 U9087 ( .A(n7466), .B(n7854), .ZN(n7469) );
  OAI22_X1 U9088 ( .A1(n7467), .A2(n6188), .B1(n8414), .B2(n8430), .ZN(n7468)
         );
  AOI21_X1 U9089 ( .B1(n7469), .B2(n8434), .A(n7468), .ZN(n10048) );
  NOR2_X1 U9090 ( .A1(n10048), .A2(n8406), .ZN(n7470) );
  AOI211_X1 U9091 ( .C1(n10053), .C2(n8265), .A(n7471), .B(n7470), .ZN(n7472)
         );
  INV_X1 U9092 ( .A(n7472), .ZN(P2_U3284) );
  NAND2_X1 U9093 ( .A1(n4323), .A2(n7473), .ZN(n7474) );
  XNOR2_X1 U9094 ( .A(n7475), .B(n7474), .ZN(n7482) );
  INV_X1 U9095 ( .A(n7476), .ZN(n7478) );
  NOR2_X1 U9096 ( .A1(n8732), .A2(n9797), .ZN(n7477) );
  AOI211_X1 U9097 ( .C1(n8734), .C2(n9770), .A(n7478), .B(n7477), .ZN(n7479)
         );
  OAI21_X1 U9098 ( .B1(n8736), .B2(n9765), .A(n7479), .ZN(n7480) );
  AOI21_X1 U9099 ( .B1(n8738), .B2(n9779), .A(n7480), .ZN(n7481) );
  OAI21_X1 U9100 ( .B1(n7482), .B2(n8740), .A(n7481), .ZN(P1_U3232) );
  XNOR2_X1 U9101 ( .A(n10046), .B(n7650), .ZN(n7483) );
  NAND2_X1 U9102 ( .A1(n8040), .A2(n10050), .ZN(n7484) );
  NAND2_X1 U9103 ( .A1(n7483), .A2(n7484), .ZN(n7534) );
  INV_X1 U9104 ( .A(n7483), .ZN(n7486) );
  INV_X1 U9105 ( .A(n7484), .ZN(n7485) );
  NAND2_X1 U9106 ( .A1(n7486), .A2(n7485), .ZN(n7536) );
  NAND2_X1 U9107 ( .A1(n7534), .A2(n7536), .ZN(n7492) );
  INV_X1 U9108 ( .A(n7487), .ZN(n7488) );
  NAND2_X1 U9109 ( .A1(n7489), .A2(n7488), .ZN(n7490) );
  XOR2_X1 U9110 ( .A(n7492), .B(n7535), .Z(n7498) );
  AOI22_X1 U9111 ( .A1(n7795), .A2(n8041), .B1(n7794), .B2(n7493), .ZN(n7495)
         );
  OAI211_X1 U9112 ( .C1(n8414), .C2(n7803), .A(n7495), .B(n7494), .ZN(n7496)
         );
  AOI21_X1 U9113 ( .B1(n10046), .B2(n4310), .A(n7496), .ZN(n7497) );
  OAI21_X1 U9114 ( .B1(n7498), .B2(n7810), .A(n7497), .ZN(P2_U3226) );
  AND2_X1 U9115 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9039) );
  AOI21_X1 U9116 ( .B1(n8734), .B2(n9773), .A(n9039), .ZN(n7501) );
  INV_X1 U9117 ( .A(n9790), .ZN(n7499) );
  NAND2_X1 U9118 ( .A1(n8723), .A2(n7499), .ZN(n7500) );
  OAI211_X1 U9119 ( .C1(n9799), .C2(n8732), .A(n7501), .B(n7500), .ZN(n7508)
         );
  INV_X1 U9120 ( .A(n7502), .ZN(n7506) );
  AOI21_X1 U9121 ( .B1(n7369), .B2(n7504), .A(n7503), .ZN(n7505) );
  NOR3_X1 U9122 ( .A1(n7506), .A2(n7505), .A3(n8740), .ZN(n7507) );
  AOI211_X1 U9123 ( .C1(n8738), .C2(n9809), .A(n7508), .B(n7507), .ZN(n7509)
         );
  INV_X1 U9124 ( .A(n7509), .ZN(P1_U3234) );
  INV_X1 U9125 ( .A(n7510), .ZN(n7533) );
  AOI22_X1 U9126 ( .A1(n7511), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n8594), .ZN(n7512) );
  OAI21_X1 U9127 ( .B1(n7533), .B2(n7545), .A(n7512), .ZN(P2_U3332) );
  INV_X1 U9128 ( .A(n9017), .ZN(n8756) );
  NAND2_X1 U9129 ( .A1(n9809), .A2(n8756), .ZN(n8768) );
  OR2_X1 U9130 ( .A1(n9809), .A2(n8756), .ZN(n7552) );
  NAND2_X1 U9131 ( .A1(n7553), .A2(n7552), .ZN(n7514) );
  OR2_X1 U9132 ( .A1(n7548), .A2(n9797), .ZN(n8769) );
  NAND2_X1 U9133 ( .A1(n7548), .A2(n9797), .ZN(n8776) );
  NAND2_X1 U9134 ( .A1(n8769), .A2(n8776), .ZN(n8879) );
  XNOR2_X1 U9135 ( .A(n7514), .B(n8879), .ZN(n7515) );
  NAND2_X1 U9136 ( .A1(n7515), .A2(n9768), .ZN(n7517) );
  AOI22_X1 U9137 ( .A1(n9771), .A2(n9016), .B1(n9017), .B2(n9772), .ZN(n7516)
         );
  NAND2_X1 U9138 ( .A1(n7517), .A2(n7516), .ZN(n9834) );
  INV_X1 U9139 ( .A(n9834), .ZN(n7530) );
  OR2_X1 U9140 ( .A1(n9735), .A2(n9018), .ZN(n7519) );
  NAND2_X1 U9141 ( .A1(n9809), .A2(n9017), .ZN(n7520) );
  XOR2_X1 U9142 ( .A(n8879), .B(n7550), .Z(n9835) );
  NAND2_X1 U9143 ( .A1(n9835), .A2(n7521), .ZN(n7529) );
  OAI22_X1 U9144 ( .A1(n9792), .A2(n7523), .B1(n7522), .B2(n9789), .ZN(n7527)
         );
  INV_X1 U9145 ( .A(n9809), .ZN(n9836) );
  NAND2_X1 U9146 ( .A1(n9783), .A2(n9836), .ZN(n9785) );
  INV_X1 U9147 ( .A(n9785), .ZN(n7524) );
  OR2_X2 U9148 ( .A1(n9785), .A2(n7548), .ZN(n9760) );
  OAI211_X1 U9149 ( .C1(n7524), .C2(n9832), .A(n9816), .B(n9760), .ZN(n9831)
         );
  NOR2_X1 U9150 ( .A1(n9831), .A2(n7525), .ZN(n7526) );
  AOI211_X1 U9151 ( .C1(n9810), .C2(n7548), .A(n7527), .B(n7526), .ZN(n7528)
         );
  OAI211_X1 U9152 ( .C1(n9806), .C2(n7530), .A(n7529), .B(n7528), .ZN(P1_U3279) );
  OAI222_X1 U9153 ( .A1(n9512), .A2(n7533), .B1(P1_U3084), .B2(n7532), .C1(
        n7531), .C2(n7689), .ZN(P1_U3327) );
  NAND2_X1 U9154 ( .A1(n7535), .A2(n7534), .ZN(n7537) );
  NAND2_X1 U9155 ( .A1(n7537), .A2(n7536), .ZN(n7592) );
  XNOR2_X1 U9156 ( .A(n8449), .B(n7666), .ZN(n7595) );
  NAND2_X1 U9157 ( .A1(n8039), .A2(n10050), .ZN(n7593) );
  XNOR2_X1 U9158 ( .A(n7595), .B(n7593), .ZN(n7591) );
  XNOR2_X1 U9159 ( .A(n7592), .B(n7591), .ZN(n7542) );
  AOI22_X1 U9160 ( .A1(n7795), .A2(n8040), .B1(n7794), .B2(n8439), .ZN(n7539)
         );
  OAI211_X1 U9161 ( .C1(n8431), .C2(n7803), .A(n7539), .B(n7538), .ZN(n7540)
         );
  AOI21_X1 U9162 ( .B1(n8449), .B2(n4310), .A(n7540), .ZN(n7541) );
  OAI21_X1 U9163 ( .B1(n7542), .B2(n7810), .A(n7541), .ZN(P2_U3236) );
  INV_X1 U9164 ( .A(n7543), .ZN(n7547) );
  AOI22_X1 U9165 ( .A1(n8025), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n8594), .ZN(n7544) );
  OAI21_X1 U9166 ( .B1(n7547), .B2(n7545), .A(n7544), .ZN(P2_U3331) );
  OAI222_X1 U9167 ( .A1(n9512), .A2(n7547), .B1(n6211), .B2(P1_U3084), .C1(
        n7546), .C2(n7689), .ZN(P1_U3326) );
  AND2_X1 U9168 ( .A1(n7548), .A2(n9773), .ZN(n7549) );
  NOR2_X1 U9169 ( .A1(n9779), .A2(n9016), .ZN(n7551) );
  INV_X1 U9170 ( .A(n9779), .ZN(n9825) );
  INV_X1 U9171 ( .A(n9770), .ZN(n9105) );
  NAND2_X1 U9172 ( .A1(n9486), .A2(n9105), .ZN(n8772) );
  NAND2_X1 U9173 ( .A1(n9133), .A2(n8772), .ZN(n7556) );
  XNOR2_X1 U9174 ( .A(n9103), .B(n7556), .ZN(n9488) );
  AND2_X1 U9175 ( .A1(n8769), .A2(n7552), .ZN(n8778) );
  NAND2_X1 U9176 ( .A1(n7553), .A2(n8778), .ZN(n7554) );
  XNOR2_X1 U9177 ( .A(n9779), .B(n9016), .ZN(n9766) );
  NAND2_X1 U9178 ( .A1(n9767), .A2(n9766), .ZN(n7555) );
  NAND2_X1 U9179 ( .A1(n9779), .A2(n8771), .ZN(n8767) );
  OAI211_X1 U9180 ( .C1(n4868), .C2(n7557), .A(n9134), .B(n9768), .ZN(n7559)
         );
  AOI22_X1 U9181 ( .A1(n9771), .A2(n9107), .B1(n9016), .B2(n9772), .ZN(n7558)
         );
  NAND2_X1 U9182 ( .A1(n7559), .A2(n7558), .ZN(n9484) );
  INV_X1 U9183 ( .A(n9761), .ZN(n7560) );
  AOI211_X1 U9184 ( .C1(n9486), .C2(n7560), .A(n9963), .B(n9388), .ZN(n9485)
         );
  NAND2_X1 U9185 ( .A1(n9485), .A2(n9371), .ZN(n7563) );
  INV_X1 U9186 ( .A(n7576), .ZN(n7561) );
  AOI22_X1 U9187 ( .A1(n9806), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7561), .B2(
        n9316), .ZN(n7562) );
  OAI211_X1 U9188 ( .C1(n9104), .C2(n9404), .A(n7563), .B(n7562), .ZN(n7564)
         );
  AOI21_X1 U9189 ( .B1(n9484), .B2(n9792), .A(n7564), .ZN(n7565) );
  OAI21_X1 U9190 ( .B1(n9488), .B2(n9398), .A(n7565), .ZN(P1_U3277) );
  INV_X1 U9191 ( .A(n8616), .ZN(n7690) );
  NAND2_X1 U9192 ( .A1(n8594), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7566) );
  OAI211_X1 U9193 ( .C1(n7690), .C2(n8597), .A(n7567), .B(n7566), .ZN(P2_U3330) );
  NAND2_X1 U9194 ( .A1(n7568), .A2(n7569), .ZN(n7570) );
  XOR2_X1 U9195 ( .A(n7571), .B(n7570), .Z(n7579) );
  INV_X1 U9196 ( .A(n7572), .ZN(n7574) );
  NOR2_X1 U9197 ( .A1(n8732), .A2(n8771), .ZN(n7573) );
  AOI211_X1 U9198 ( .C1(n8734), .C2(n9107), .A(n7574), .B(n7573), .ZN(n7575)
         );
  OAI21_X1 U9199 ( .B1(n8736), .B2(n7576), .A(n7575), .ZN(n7577) );
  AOI21_X1 U9200 ( .B1(n9486), .B2(n8738), .A(n7577), .ZN(n7578) );
  OAI21_X1 U9201 ( .B1(n7579), .B2(n8740), .A(n7578), .ZN(P1_U3213) );
  INV_X1 U9202 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8827) );
  NAND2_X1 U9203 ( .A1(n7583), .A2(n7582), .ZN(n7581) );
  NAND2_X1 U9204 ( .A1(n7581), .A2(n7580), .ZN(n7585) );
  MUX2_X1 U9205 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7824), .Z(n7821) );
  XNOR2_X1 U9206 ( .A(n7821), .B(SI_30_), .ZN(n7586) );
  INV_X1 U9207 ( .A(n8826), .ZN(n8593) );
  OAI222_X1 U9208 ( .A1(n7689), .A2(n8827), .B1(n9512), .B2(n8593), .C1(
        P1_U3084), .C2(n7587), .ZN(P1_U3323) );
  NOR2_X1 U9209 ( .A1(n8196), .A2(n8539), .ZN(n7588) );
  XNOR2_X1 U9210 ( .A(n7588), .B(n7650), .ZN(n7589) );
  XNOR2_X1 U9211 ( .A(n8459), .B(n7589), .ZN(n7676) );
  INV_X1 U9212 ( .A(n7676), .ZN(n7590) );
  NAND2_X1 U9213 ( .A1(n7590), .A2(n7789), .ZN(n7681) );
  NAND2_X1 U9214 ( .A1(n7592), .A2(n7591), .ZN(n7597) );
  INV_X1 U9215 ( .A(n7593), .ZN(n7594) );
  NAND2_X1 U9216 ( .A1(n7595), .A2(n7594), .ZN(n7596) );
  XNOR2_X1 U9217 ( .A(n8538), .B(n7650), .ZN(n7598) );
  NAND2_X1 U9218 ( .A1(n8038), .A2(n10050), .ZN(n7599) );
  NAND2_X1 U9219 ( .A1(n7598), .A2(n7599), .ZN(n7604) );
  INV_X1 U9220 ( .A(n7598), .ZN(n7601) );
  INV_X1 U9221 ( .A(n7599), .ZN(n7600) );
  NAND2_X1 U9222 ( .A1(n7601), .A2(n7600), .ZN(n7602) );
  NAND2_X1 U9223 ( .A1(n7604), .A2(n7602), .ZN(n7702) );
  NOR2_X1 U9224 ( .A1(n8413), .A2(n8539), .ZN(n7801) );
  XNOR2_X1 U9225 ( .A(n8533), .B(n7666), .ZN(n7744) );
  XNOR2_X1 U9226 ( .A(n8524), .B(n7650), .ZN(n7605) );
  NAND2_X1 U9227 ( .A1(n8036), .A2(n10050), .ZN(n7606) );
  NAND2_X1 U9228 ( .A1(n7605), .A2(n7606), .ZN(n7747) );
  OAI21_X1 U9229 ( .B1(n7801), .B2(n7744), .A(n7747), .ZN(n7611) );
  NAND3_X1 U9230 ( .A1(n7747), .A2(n7801), .A3(n7744), .ZN(n7609) );
  INV_X1 U9231 ( .A(n7605), .ZN(n7608) );
  INV_X1 U9232 ( .A(n7606), .ZN(n7607) );
  NAND2_X1 U9233 ( .A1(n7608), .A2(n7607), .ZN(n7746) );
  AND2_X1 U9234 ( .A1(n7609), .A2(n7746), .ZN(n7610) );
  XNOR2_X1 U9235 ( .A(n8521), .B(n7666), .ZN(n7614) );
  NAND2_X1 U9236 ( .A1(n8342), .A2(n10050), .ZN(n7612) );
  XNOR2_X1 U9237 ( .A(n7614), .B(n7612), .ZN(n7754) );
  NAND2_X1 U9238 ( .A1(n7755), .A2(n7754), .ZN(n7616) );
  INV_X1 U9239 ( .A(n7612), .ZN(n7613) );
  NAND2_X1 U9240 ( .A1(n7614), .A2(n7613), .ZN(n7615) );
  NAND2_X1 U9241 ( .A1(n7616), .A2(n7615), .ZN(n7782) );
  XNOR2_X1 U9242 ( .A(n8514), .B(n7666), .ZN(n7619) );
  NAND2_X1 U9243 ( .A1(n8327), .A2(n10050), .ZN(n7617) );
  XNOR2_X1 U9244 ( .A(n7619), .B(n7617), .ZN(n7783) );
  NAND2_X1 U9245 ( .A1(n7782), .A2(n7783), .ZN(n7621) );
  INV_X1 U9246 ( .A(n7617), .ZN(n7618) );
  NAND2_X1 U9247 ( .A1(n7619), .A2(n7618), .ZN(n7620) );
  XNOR2_X1 U9248 ( .A(n8510), .B(n7650), .ZN(n7622) );
  NAND2_X1 U9249 ( .A1(n8344), .A2(n10050), .ZN(n7623) );
  NAND2_X1 U9250 ( .A1(n7622), .A2(n7623), .ZN(n7628) );
  INV_X1 U9251 ( .A(n7622), .ZN(n7625) );
  INV_X1 U9252 ( .A(n7623), .ZN(n7624) );
  NAND2_X1 U9253 ( .A1(n7625), .A2(n7624), .ZN(n7626) );
  NAND2_X1 U9254 ( .A1(n7628), .A2(n7626), .ZN(n7720) );
  XNOR2_X1 U9255 ( .A(n8504), .B(n7666), .ZN(n7629) );
  NOR2_X1 U9256 ( .A1(n7729), .A2(n8539), .ZN(n7630) );
  XNOR2_X1 U9257 ( .A(n7629), .B(n7630), .ZN(n7767) );
  INV_X1 U9258 ( .A(n7629), .ZN(n7632) );
  INV_X1 U9259 ( .A(n7630), .ZN(n7631) );
  XNOR2_X1 U9260 ( .A(n8499), .B(n7666), .ZN(n7635) );
  NAND2_X1 U9261 ( .A1(n8311), .A2(n10050), .ZN(n7633) );
  XNOR2_X1 U9262 ( .A(n7635), .B(n7633), .ZN(n7727) );
  NAND2_X1 U9263 ( .A1(n7726), .A2(n7727), .ZN(n7637) );
  INV_X1 U9264 ( .A(n7633), .ZN(n7634) );
  NAND2_X1 U9265 ( .A1(n7635), .A2(n7634), .ZN(n7636) );
  NAND2_X1 U9266 ( .A1(n7637), .A2(n7636), .ZN(n7640) );
  XNOR2_X1 U9267 ( .A(n8493), .B(n7650), .ZN(n7638) );
  XNOR2_X1 U9268 ( .A(n7640), .B(n7638), .ZN(n7774) );
  NAND2_X1 U9269 ( .A1(n8297), .A2(n10050), .ZN(n7776) );
  NAND2_X1 U9270 ( .A1(n7774), .A2(n7776), .ZN(n7775) );
  INV_X1 U9271 ( .A(n7638), .ZN(n7639) );
  OR2_X1 U9272 ( .A1(n7640), .A2(n7639), .ZN(n7641) );
  NAND2_X2 U9273 ( .A1(n7775), .A2(n7641), .ZN(n7653) );
  XNOR2_X1 U9274 ( .A(n8484), .B(n7650), .ZN(n7642) );
  NAND2_X1 U9275 ( .A1(n7653), .A2(n7642), .ZN(n7708) );
  NOR2_X1 U9276 ( .A1(n8284), .A2(n8539), .ZN(n7649) );
  NAND2_X1 U9277 ( .A1(n7708), .A2(n7649), .ZN(n7643) );
  OR2_X1 U9278 ( .A1(n7653), .A2(n7642), .ZN(n7709) );
  NAND2_X1 U9279 ( .A1(n7643), .A2(n7709), .ZN(n7645) );
  XNOR2_X1 U9280 ( .A(n8479), .B(n7666), .ZN(n7644) );
  NAND2_X1 U9281 ( .A1(n7645), .A2(n7644), .ZN(n7659) );
  NAND2_X1 U9282 ( .A1(n7649), .A2(n7650), .ZN(n7646) );
  OAI21_X1 U9283 ( .B1(n8484), .B2(n7649), .A(n7646), .ZN(n7647) );
  XNOR2_X1 U9284 ( .A(n7647), .B(n8479), .ZN(n7648) );
  OR2_X2 U9285 ( .A1(n7653), .A2(n7648), .ZN(n7655) );
  INV_X1 U9286 ( .A(n7649), .ZN(n7710) );
  MUX2_X1 U9287 ( .A(n8484), .B(n7650), .S(n7710), .Z(n7651) );
  XNOR2_X1 U9288 ( .A(n7651), .B(n8479), .ZN(n7652) );
  NAND2_X1 U9289 ( .A1(n7653), .A2(n7652), .ZN(n7654) );
  INV_X1 U9290 ( .A(n7762), .ZN(n7657) );
  NAND2_X1 U9291 ( .A1(n8035), .A2(n10050), .ZN(n7761) );
  INV_X1 U9292 ( .A(n7761), .ZN(n7656) );
  NAND2_X1 U9293 ( .A1(n7659), .A2(n7658), .ZN(n7737) );
  XNOR2_X1 U9294 ( .A(n8476), .B(n7666), .ZN(n7735) );
  NAND2_X1 U9295 ( .A1(n8034), .A2(n10050), .ZN(n7734) );
  XNOR2_X1 U9296 ( .A(n8471), .B(n7666), .ZN(n7660) );
  NOR2_X1 U9297 ( .A1(n8226), .A2(n8539), .ZN(n7661) );
  NAND2_X1 U9298 ( .A1(n7660), .A2(n7661), .ZN(n7665) );
  INV_X1 U9299 ( .A(n7660), .ZN(n7663) );
  INV_X1 U9300 ( .A(n7661), .ZN(n7662) );
  NAND2_X1 U9301 ( .A1(n7663), .A2(n7662), .ZN(n7664) );
  AND2_X1 U9302 ( .A1(n7665), .A2(n7664), .ZN(n7791) );
  NAND2_X1 U9303 ( .A1(n7790), .A2(n7665), .ZN(n7692) );
  XNOR2_X1 U9304 ( .A(n8464), .B(n7666), .ZN(n7667) );
  NOR2_X1 U9305 ( .A1(n8210), .A2(n8539), .ZN(n7668) );
  NAND2_X1 U9306 ( .A1(n7667), .A2(n7668), .ZN(n7675) );
  INV_X1 U9307 ( .A(n7667), .ZN(n7670) );
  INV_X1 U9308 ( .A(n7668), .ZN(n7669) );
  NAND2_X1 U9309 ( .A1(n7670), .A2(n7669), .ZN(n7671) );
  NAND4_X1 U9310 ( .A1(n7691), .A2(n7789), .A3(n7675), .A4(n7676), .ZN(n7680)
         );
  INV_X1 U9311 ( .A(n7672), .ZN(n8181) );
  AOI22_X1 U9312 ( .A1(n7793), .A2(n8181), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n7674) );
  NAND2_X1 U9313 ( .A1(n7795), .A2(n8180), .ZN(n7673) );
  OAI211_X1 U9314 ( .C1(n8174), .C2(n7805), .A(n7674), .B(n7673), .ZN(n7678)
         );
  NOR3_X1 U9315 ( .A1(n7676), .A2(n7675), .A3(n7810), .ZN(n7677) );
  AOI211_X1 U9316 ( .C1(n8459), .C2(n4310), .A(n7678), .B(n7677), .ZN(n7679)
         );
  OAI211_X1 U9317 ( .C1(n7681), .C2(n7691), .A(n7680), .B(n7679), .ZN(P2_U3222) );
  AOI22_X1 U9318 ( .A1(n10001), .A2(n4310), .B1(n7682), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n7687) );
  INV_X1 U9319 ( .A(n7868), .ZN(n7683) );
  MUX2_X1 U9320 ( .A(n7683), .B(n10001), .S(n8539), .Z(n7684) );
  OAI21_X1 U9321 ( .B1(n7685), .B2(n7684), .A(n7789), .ZN(n7686) );
  OAI211_X1 U9322 ( .C1(n7803), .C2(n5789), .A(n7687), .B(n7686), .ZN(P2_U3234) );
  INV_X1 U9323 ( .A(n8841), .ZN(n8598) );
  INV_X1 U9324 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8842) );
  OAI222_X1 U9325 ( .A1(n9512), .A2(n8598), .B1(P1_U3084), .B2(n7688), .C1(
        n8842), .C2(n7689), .ZN(P1_U3324) );
  INV_X1 U9326 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8617) );
  OAI222_X1 U9327 ( .A1(n9512), .A2(n7690), .B1(P1_U3084), .B2(n4312), .C1(
        n8617), .C2(n7689), .ZN(P1_U3325) );
  OAI211_X1 U9328 ( .C1(n7693), .C2(n7692), .A(n7691), .B(n7789), .ZN(n7698)
         );
  AOI22_X1 U9329 ( .A1(n8032), .A2(n7793), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        n7694), .ZN(n7697) );
  AOI22_X1 U9330 ( .A1(n7795), .A2(n8033), .B1(n7794), .B2(n8190), .ZN(n7696)
         );
  NAND2_X1 U9331 ( .A1(n8464), .A2(n4310), .ZN(n7695) );
  NAND4_X1 U9332 ( .A1(n7698), .A2(n7697), .A3(n7696), .A4(n7695), .ZN(
        P2_U3216) );
  INV_X1 U9333 ( .A(n7699), .ZN(n7700) );
  AOI21_X1 U9334 ( .B1(n7702), .B2(n7701), .A(n7700), .ZN(n7707) );
  AOI22_X1 U9335 ( .A1(n7795), .A2(n8039), .B1(n7794), .B2(n8405), .ZN(n7704)
         );
  OAI211_X1 U9336 ( .C1(n8413), .C2(n7803), .A(n7704), .B(n7703), .ZN(n7705)
         );
  AOI21_X1 U9337 ( .B1(n8538), .B2(n4310), .A(n7705), .ZN(n7706) );
  OAI21_X1 U9338 ( .B1(n7707), .B2(n7810), .A(n7706), .ZN(P2_U3217) );
  NAND2_X1 U9339 ( .A1(n7709), .A2(n7708), .ZN(n7711) );
  XNOR2_X1 U9340 ( .A(n7711), .B(n7710), .ZN(n7717) );
  OAI22_X1 U9341 ( .A1(n7803), .A2(n8258), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7712), .ZN(n7715) );
  INV_X1 U9342 ( .A(n8267), .ZN(n7713) );
  OAI22_X1 U9343 ( .A1(n7806), .A2(n8257), .B1(n7805), .B2(n7713), .ZN(n7714)
         );
  AOI211_X1 U9344 ( .C1(n8484), .C2(n4310), .A(n7715), .B(n7714), .ZN(n7716)
         );
  OAI21_X1 U9345 ( .B1(n7717), .B2(n7810), .A(n7716), .ZN(P2_U3218) );
  INV_X1 U9346 ( .A(n7718), .ZN(n7719) );
  AOI21_X1 U9347 ( .B1(n7721), .B2(n7720), .A(n7719), .ZN(n7725) );
  AOI22_X1 U9348 ( .A1(n7795), .A2(n8327), .B1(n7794), .B2(n8321), .ZN(n7722)
         );
  NAND2_X1 U9349 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8155) );
  OAI211_X1 U9350 ( .C1(n7729), .C2(n7803), .A(n7722), .B(n8155), .ZN(n7723)
         );
  AOI21_X1 U9351 ( .B1(n8510), .B2(n4310), .A(n7723), .ZN(n7724) );
  OAI21_X1 U9352 ( .B1(n7725), .B2(n7810), .A(n7724), .ZN(P2_U3221) );
  XNOR2_X1 U9353 ( .A(n7726), .B(n7727), .ZN(n7733) );
  OAI22_X1 U9354 ( .A1(n7803), .A2(n8257), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9648), .ZN(n7731) );
  INV_X1 U9355 ( .A(n8293), .ZN(n7728) );
  OAI22_X1 U9356 ( .A1(n7806), .A2(n7729), .B1(n7805), .B2(n7728), .ZN(n7730)
         );
  AOI211_X1 U9357 ( .C1(n8499), .C2(n4310), .A(n7731), .B(n7730), .ZN(n7732)
         );
  OAI21_X1 U9358 ( .B1(n7733), .B2(n7810), .A(n7732), .ZN(P2_U3225) );
  XNOR2_X1 U9359 ( .A(n7735), .B(n7734), .ZN(n7736) );
  XNOR2_X1 U9360 ( .A(n7737), .B(n7736), .ZN(n7742) );
  OAI22_X1 U9361 ( .A1(n7806), .A2(n8258), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7738), .ZN(n7740) );
  OAI22_X1 U9362 ( .A1(n7803), .A2(n8226), .B1(n7805), .B2(n8228), .ZN(n7739)
         );
  AOI211_X1 U9363 ( .C1(n8476), .C2(n4310), .A(n7740), .B(n7739), .ZN(n7741)
         );
  OAI21_X1 U9364 ( .B1(n7742), .B2(n7810), .A(n7741), .ZN(P2_U3227) );
  XNOR2_X1 U9365 ( .A(n7743), .B(n7744), .ZN(n7802) );
  INV_X1 U9366 ( .A(n7743), .ZN(n7745) );
  AOI22_X1 U9367 ( .A1(n7802), .A2(n7801), .B1(n7745), .B2(n7744), .ZN(n7749)
         );
  NAND2_X1 U9368 ( .A1(n7747), .A2(n7746), .ZN(n7748) );
  XNOR2_X1 U9369 ( .A(n7749), .B(n7748), .ZN(n7753) );
  AOI22_X1 U9370 ( .A1(n7795), .A2(n8037), .B1(n7794), .B2(n8374), .ZN(n7750)
         );
  NAND2_X1 U9371 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8096) );
  OAI211_X1 U9372 ( .C1(n8369), .C2(n7803), .A(n7750), .B(n8096), .ZN(n7751)
         );
  AOI21_X1 U9373 ( .B1(n8524), .B2(n4310), .A(n7751), .ZN(n7752) );
  OAI21_X1 U9374 ( .B1(n7753), .B2(n7810), .A(n7752), .ZN(P2_U3228) );
  XNOR2_X1 U9375 ( .A(n7755), .B(n7754), .ZN(n7760) );
  OAI22_X1 U9376 ( .A1(n7803), .A2(n8355), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9661), .ZN(n7758) );
  INV_X1 U9377 ( .A(n8359), .ZN(n7756) );
  OAI22_X1 U9378 ( .A1(n7806), .A2(n8393), .B1(n7805), .B2(n7756), .ZN(n7757)
         );
  AOI211_X1 U9379 ( .C1(n8521), .C2(n4310), .A(n7758), .B(n7757), .ZN(n7759)
         );
  OAI21_X1 U9380 ( .B1(n7760), .B2(n7810), .A(n7759), .ZN(P2_U3230) );
  XNOR2_X1 U9381 ( .A(n7762), .B(n7761), .ZN(n7766) );
  OAI22_X1 U9382 ( .A1(n7803), .A2(n8245), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9673), .ZN(n7764) );
  OAI22_X1 U9383 ( .A1(n7806), .A2(n8284), .B1(n7805), .B2(n8238), .ZN(n7763)
         );
  AOI211_X1 U9384 ( .C1(n8479), .C2(n4310), .A(n7764), .B(n7763), .ZN(n7765)
         );
  OAI21_X1 U9385 ( .B1(n7766), .B2(n7810), .A(n7765), .ZN(P2_U3231) );
  XNOR2_X1 U9386 ( .A(n7768), .B(n7767), .ZN(n7773) );
  OAI22_X1 U9387 ( .A1(n7803), .A2(n8283), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9642), .ZN(n7771) );
  INV_X1 U9388 ( .A(n8307), .ZN(n7769) );
  OAI22_X1 U9389 ( .A1(n7806), .A2(n7785), .B1(n7805), .B2(n7769), .ZN(n7770)
         );
  AOI211_X1 U9390 ( .C1(n8504), .C2(n4310), .A(n7771), .B(n7770), .ZN(n7772)
         );
  OAI21_X1 U9391 ( .B1(n7773), .B2(n7810), .A(n7772), .ZN(P2_U3235) );
  OAI21_X1 U9392 ( .B1(n7774), .B2(n7776), .A(n7775), .ZN(n7777) );
  NAND2_X1 U9393 ( .A1(n7777), .A2(n7789), .ZN(n7781) );
  OAI22_X1 U9394 ( .A1(n7803), .A2(n8284), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9606), .ZN(n7779) );
  OAI22_X1 U9395 ( .A1(n7806), .A2(n8283), .B1(n7805), .B2(n8274), .ZN(n7778)
         );
  AOI211_X1 U9396 ( .C1(n8493), .C2(n4310), .A(n7779), .B(n7778), .ZN(n7780)
         );
  NAND2_X1 U9397 ( .A1(n7781), .A2(n7780), .ZN(P2_U3237) );
  XNOR2_X1 U9398 ( .A(n7782), .B(n7783), .ZN(n7788) );
  AOI22_X1 U9399 ( .A1(n7795), .A2(n8342), .B1(n7794), .B2(n8335), .ZN(n7784)
         );
  NAND2_X1 U9400 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8133) );
  OAI211_X1 U9401 ( .C1(n7785), .C2(n7803), .A(n7784), .B(n8133), .ZN(n7786)
         );
  AOI21_X1 U9402 ( .B1(n8514), .B2(n4310), .A(n7786), .ZN(n7787) );
  OAI21_X1 U9403 ( .B1(n7788), .B2(n7810), .A(n7787), .ZN(P2_U3240) );
  OAI211_X1 U9404 ( .C1(n7792), .C2(n7791), .A(n7790), .B(n7789), .ZN(n7800)
         );
  AOI22_X1 U9405 ( .A1(n7793), .A2(n8180), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n7799) );
  AOI22_X1 U9406 ( .A1(n7795), .A2(n8034), .B1(n7794), .B2(n8214), .ZN(n7798)
         );
  NAND2_X1 U9407 ( .A1(n8471), .A2(n4310), .ZN(n7797) );
  NAND4_X1 U9408 ( .A1(n7800), .A2(n7799), .A3(n7798), .A4(n7797), .ZN(
        P2_U3242) );
  XNOR2_X1 U9409 ( .A(n7802), .B(n7801), .ZN(n7811) );
  OAI22_X1 U9410 ( .A1(n7803), .A2(n8393), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5939), .ZN(n7808) );
  INV_X1 U9411 ( .A(n8387), .ZN(n7804) );
  OAI22_X1 U9412 ( .A1(n7806), .A2(n8431), .B1(n7805), .B2(n7804), .ZN(n7807)
         );
  AOI211_X1 U9413 ( .C1(n8533), .C2(n4310), .A(n7808), .B(n7807), .ZN(n7809)
         );
  OAI21_X1 U9414 ( .B1(n7811), .B2(n7810), .A(n7809), .ZN(P2_U3243) );
  NAND2_X1 U9415 ( .A1(n8826), .A2(n7828), .ZN(n7814) );
  NAND2_X1 U9416 ( .A1(n7812), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7813) );
  NOR2_X1 U9417 ( .A1(n8159), .A2(n7815), .ZN(n7817) );
  INV_X1 U9418 ( .A(n8005), .ZN(n7816) );
  AOI21_X1 U9419 ( .B1(n9754), .B2(n7817), .A(n7816), .ZN(n7819) );
  NOR2_X1 U9420 ( .A1(n9754), .A2(n6187), .ZN(n8007) );
  INV_X1 U9421 ( .A(n7817), .ZN(n7818) );
  AOI22_X1 U9422 ( .A1(n7820), .A2(n7819), .B1(n8007), .B2(n7818), .ZN(n7832)
         );
  INV_X1 U9423 ( .A(n7821), .ZN(n7822) );
  MUX2_X1 U9424 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7824), .Z(n7825) );
  INV_X1 U9425 ( .A(SI_31_), .ZN(n9658) );
  XNOR2_X1 U9426 ( .A(n7825), .B(n9658), .ZN(n7826) );
  NAND2_X1 U9427 ( .A1(n8836), .A2(n7828), .ZN(n7830) );
  NAND2_X1 U9428 ( .A1(n5821), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7829) );
  INV_X1 U9429 ( .A(n8159), .ZN(n7831) );
  OR2_X1 U9430 ( .A1(n9749), .A2(n7831), .ZN(n8013) );
  NAND2_X1 U9431 ( .A1(n9754), .A2(n6187), .ZN(n8006) );
  NAND2_X1 U9432 ( .A1(n8013), .A2(n8006), .ZN(n8011) );
  NAND2_X1 U9433 ( .A1(n9749), .A2(n7831), .ZN(n8014) );
  OAI21_X1 U9434 ( .B1(n7832), .B2(n8011), .A(n8014), .ZN(n7834) );
  XNOR2_X1 U9435 ( .A(n7834), .B(n7833), .ZN(n7835) );
  INV_X1 U9436 ( .A(n8007), .ZN(n7837) );
  NAND2_X1 U9437 ( .A1(n8014), .A2(n7837), .ZN(n8010) );
  INV_X1 U9438 ( .A(n8367), .ZN(n7942) );
  NOR2_X1 U9439 ( .A1(n7839), .A2(n7838), .ZN(n7846) );
  NOR2_X1 U9440 ( .A1(n6160), .A2(n7840), .ZN(n7845) );
  NAND3_X1 U9441 ( .A1(n6158), .A2(n7868), .A3(n7841), .ZN(n7842) );
  NOR2_X1 U9442 ( .A1(n7871), .A2(n7842), .ZN(n7844) );
  NAND4_X1 U9443 ( .A1(n7846), .A2(n7845), .A3(n7844), .A4(n7843), .ZN(n7848)
         );
  NOR3_X1 U9444 ( .A1(n7848), .A2(n5878), .A3(n7847), .ZN(n7852) );
  AND4_X1 U9445 ( .A1(n7852), .A2(n7851), .A3(n7850), .A4(n7849), .ZN(n7853)
         );
  NAND4_X1 U9446 ( .A1(n7932), .A2(n8423), .A3(n7854), .A4(n7853), .ZN(n7855)
         );
  NOR2_X1 U9447 ( .A1(n8391), .A2(n7855), .ZN(n7856) );
  NAND4_X1 U9448 ( .A1(n8339), .A2(n8352), .A3(n7942), .A4(n7856), .ZN(n7857)
         );
  NOR2_X1 U9449 ( .A1(n8317), .A2(n7857), .ZN(n7858) );
  NAND4_X1 U9450 ( .A1(n8279), .A2(n4824), .A3(n4698), .A4(n7858), .ZN(n7859)
         );
  NOR4_X1 U9451 ( .A1(n8224), .A2(n8243), .A3(n7975), .A4(n7859), .ZN(n7860)
         );
  NAND4_X1 U9452 ( .A1(n7861), .A2(n4701), .A3(n7860), .A4(n7987), .ZN(n7862)
         );
  NOR4_X1 U9453 ( .A1(n8011), .A2(n8010), .A3(n7996), .A4(n7862), .ZN(n7863)
         );
  XNOR2_X1 U9454 ( .A(n7863), .B(n8152), .ZN(n8018) );
  NAND2_X1 U9455 ( .A1(n8019), .A2(n8152), .ZN(n7864) );
  INV_X1 U9456 ( .A(n7960), .ZN(n7972) );
  NAND2_X1 U9457 ( .A1(n6158), .A2(n7868), .ZN(n7866) );
  NAND3_X1 U9458 ( .A1(n7872), .A2(n7866), .A3(n7865), .ZN(n7867) );
  NAND2_X1 U9459 ( .A1(n7867), .A2(n7869), .ZN(n7875) );
  AND2_X1 U9460 ( .A1(n7868), .A2(n8019), .ZN(n7870) );
  OAI211_X1 U9461 ( .C1(n7871), .C2(n7870), .A(n7869), .B(n6158), .ZN(n7873)
         );
  NAND2_X1 U9462 ( .A1(n7873), .A2(n7872), .ZN(n7874) );
  MUX2_X1 U9463 ( .A(n7875), .B(n7874), .S(n8012), .Z(n7880) );
  NAND2_X1 U9464 ( .A1(n7889), .A2(n7890), .ZN(n7877) );
  NAND2_X1 U9465 ( .A1(n7883), .A2(n7881), .ZN(n7876) );
  MUX2_X1 U9466 ( .A(n7877), .B(n7876), .S(n8000), .Z(n7892) );
  INV_X1 U9467 ( .A(n7892), .ZN(n7878) );
  NAND3_X1 U9468 ( .A1(n7880), .A2(n7879), .A3(n7878), .ZN(n7887) );
  AND2_X1 U9469 ( .A1(n7882), .A2(n7881), .ZN(n7884) );
  OAI211_X1 U9470 ( .C1(n7892), .C2(n7884), .A(n7883), .B(n7897), .ZN(n7885)
         );
  NAND2_X1 U9471 ( .A1(n7885), .A2(n8012), .ZN(n7886) );
  NAND2_X1 U9472 ( .A1(n7887), .A2(n7886), .ZN(n7895) );
  AND2_X1 U9473 ( .A1(n7889), .A2(n7888), .ZN(n7891) );
  OAI211_X1 U9474 ( .C1(n7892), .C2(n7891), .A(n7890), .B(n7894), .ZN(n7893)
         );
  AOI22_X1 U9475 ( .A1(n7895), .A2(n7894), .B1(n8000), .B2(n7893), .ZN(n7903)
         );
  OAI21_X1 U9476 ( .B1(n7897), .B2(n8012), .A(n7896), .ZN(n7902) );
  MUX2_X1 U9477 ( .A(n7899), .B(n7898), .S(n8012), .Z(n7900) );
  OAI211_X1 U9478 ( .C1(n7903), .C2(n7902), .A(n7901), .B(n7900), .ZN(n7908)
         );
  MUX2_X1 U9479 ( .A(n7905), .B(n7904), .S(n8012), .Z(n7906) );
  NAND3_X1 U9480 ( .A1(n7908), .A2(n7907), .A3(n7906), .ZN(n7913) );
  NAND2_X1 U9481 ( .A1(n7916), .A2(n7915), .ZN(n7910) );
  INV_X1 U9482 ( .A(n7914), .ZN(n7911) );
  NAND2_X1 U9483 ( .A1(n7913), .A2(n7919), .ZN(n7923) );
  AND2_X1 U9484 ( .A1(n7925), .A2(n7914), .ZN(n7921) );
  INV_X1 U9485 ( .A(n7915), .ZN(n7918) );
  NAND2_X1 U9486 ( .A1(n7924), .A2(n7916), .ZN(n7917) );
  AOI21_X1 U9487 ( .B1(n7919), .B2(n7918), .A(n7917), .ZN(n7920) );
  NAND2_X1 U9488 ( .A1(n7923), .A2(n7922), .ZN(n7927) );
  MUX2_X1 U9489 ( .A(n7930), .B(n7929), .S(n8012), .Z(n7931) );
  NAND3_X1 U9490 ( .A1(n7933), .A2(n7932), .A3(n7931), .ZN(n7938) );
  MUX2_X1 U9491 ( .A(n7935), .B(n7934), .S(n8000), .Z(n7936) );
  NAND3_X1 U9492 ( .A1(n7938), .A2(n7937), .A3(n7936), .ZN(n7943) );
  MUX2_X1 U9493 ( .A(n7940), .B(n7939), .S(n8000), .Z(n7941) );
  MUX2_X1 U9494 ( .A(n7945), .B(n7944), .S(n8012), .Z(n7946) );
  INV_X1 U9495 ( .A(n7947), .ZN(n7950) );
  NAND2_X1 U9496 ( .A1(n7955), .A2(n7948), .ZN(n7949) );
  MUX2_X1 U9497 ( .A(n7950), .B(n7949), .S(n8000), .Z(n7952) );
  INV_X1 U9498 ( .A(n7956), .ZN(n7951) );
  NOR2_X1 U9499 ( .A1(n7952), .A2(n7951), .ZN(n7953) );
  NAND2_X1 U9500 ( .A1(n7954), .A2(n7953), .ZN(n7957) );
  INV_X1 U9501 ( .A(n7967), .ZN(n7964) );
  NAND3_X1 U9502 ( .A1(n7960), .A2(n7959), .A3(n8280), .ZN(n7963) );
  INV_X1 U9503 ( .A(n7965), .ZN(n7961) );
  OAI21_X1 U9504 ( .B1(n7968), .B2(n7961), .A(n7960), .ZN(n7962) );
  OAI21_X1 U9505 ( .B1(n7964), .B2(n7963), .A(n7962), .ZN(n7970) );
  NAND2_X1 U9506 ( .A1(n7978), .A2(n7976), .ZN(n7977) );
  NAND2_X1 U9507 ( .A1(n7984), .A2(n7980), .ZN(n7983) );
  NAND2_X1 U9508 ( .A1(n4701), .A2(n7981), .ZN(n7982) );
  MUX2_X1 U9509 ( .A(n7983), .B(n7982), .S(n8012), .Z(n7988) );
  MUX2_X1 U9510 ( .A(n7985), .B(n7984), .S(n8012), .Z(n7986) );
  OAI211_X1 U9511 ( .C1(n7989), .C2(n7988), .A(n7987), .B(n7986), .ZN(n7995)
         );
  INV_X1 U9512 ( .A(n7998), .ZN(n7990) );
  AOI21_X1 U9513 ( .B1(n8210), .B2(n8464), .A(n7990), .ZN(n7991) );
  MUX2_X1 U9514 ( .A(n7992), .B(n7991), .S(n8012), .Z(n7993) );
  NAND3_X1 U9515 ( .A1(n7995), .A2(n7994), .A3(n7993), .ZN(n7999) );
  AOI21_X1 U9516 ( .B1(n7999), .B2(n8196), .A(n7996), .ZN(n8003) );
  INV_X1 U9517 ( .A(n8004), .ZN(n7997) );
  NOR2_X1 U9518 ( .A1(n7997), .A2(n8012), .ZN(n8002) );
  OAI211_X1 U9519 ( .C1(n8000), .C2(n8459), .A(n7999), .B(n7998), .ZN(n8001)
         );
  OAI21_X1 U9520 ( .B1(n8003), .B2(n8002), .A(n8001), .ZN(n8009) );
  MUX2_X1 U9521 ( .A(n8005), .B(n8004), .S(n8012), .Z(n8008) );
  MUX2_X1 U9522 ( .A(n8011), .B(n8010), .S(n8012), .Z(n8016) );
  MUX2_X1 U9523 ( .A(n8014), .B(n8013), .S(n8012), .Z(n8015) );
  INV_X1 U9524 ( .A(n8017), .ZN(n8022) );
  OAI211_X1 U9525 ( .C1(n8022), .C2(n10002), .A(n8021), .B(n8020), .ZN(n8023)
         );
  NAND4_X1 U9526 ( .A1(n9994), .A2(n8025), .A3(n8341), .A4(n8024), .ZN(n8026)
         );
  OAI211_X1 U9527 ( .C1(n8027), .C2(n8029), .A(n8026), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8028) );
  OAI21_X1 U9528 ( .B1(n8030), .B2(n8029), .A(n8028), .ZN(P2_U3244) );
  MUX2_X1 U9529 ( .A(n8031), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8049), .Z(
        P2_U3582) );
  MUX2_X1 U9530 ( .A(n8181), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8049), .Z(
        P2_U3581) );
  MUX2_X1 U9531 ( .A(n8032), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8049), .Z(
        P2_U3580) );
  MUX2_X1 U9532 ( .A(n8180), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8049), .Z(
        P2_U3579) );
  MUX2_X1 U9533 ( .A(n8033), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8049), .Z(
        P2_U3578) );
  MUX2_X1 U9534 ( .A(n8034), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8049), .Z(
        P2_U3577) );
  MUX2_X1 U9535 ( .A(n8035), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8049), .Z(
        P2_U3576) );
  MUX2_X1 U9536 ( .A(n8297), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8049), .Z(
        P2_U3574) );
  MUX2_X1 U9537 ( .A(n8311), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8049), .Z(
        P2_U3573) );
  MUX2_X1 U9538 ( .A(n4560), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8049), .Z(
        P2_U3572) );
  MUX2_X1 U9539 ( .A(n8344), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8049), .Z(
        P2_U3571) );
  MUX2_X1 U9540 ( .A(n8327), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8049), .Z(
        P2_U3570) );
  MUX2_X1 U9541 ( .A(n8342), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8049), .Z(
        P2_U3569) );
  MUX2_X1 U9542 ( .A(n8036), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8049), .Z(
        P2_U3568) );
  MUX2_X1 U9543 ( .A(n8037), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8049), .Z(
        P2_U3567) );
  MUX2_X1 U9544 ( .A(n8038), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8049), .Z(
        P2_U3566) );
  MUX2_X1 U9545 ( .A(n8039), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8049), .Z(
        P2_U3565) );
  MUX2_X1 U9546 ( .A(n8040), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8049), .Z(
        P2_U3564) );
  MUX2_X1 U9547 ( .A(n8041), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8049), .Z(
        P2_U3563) );
  MUX2_X1 U9548 ( .A(n4587), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8049), .Z(
        P2_U3562) );
  MUX2_X1 U9549 ( .A(n8042), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8049), .Z(
        P2_U3561) );
  MUX2_X1 U9550 ( .A(n8043), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8049), .Z(
        P2_U3560) );
  MUX2_X1 U9551 ( .A(n8044), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8049), .Z(
        P2_U3559) );
  MUX2_X1 U9552 ( .A(n8045), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8049), .Z(
        P2_U3558) );
  MUX2_X1 U9553 ( .A(n8046), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8049), .Z(
        P2_U3557) );
  MUX2_X1 U9554 ( .A(n8047), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8049), .Z(
        P2_U3556) );
  MUX2_X1 U9555 ( .A(n6674), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8049), .Z(
        P2_U3555) );
  MUX2_X1 U9556 ( .A(n8048), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8049), .Z(
        P2_U3554) );
  MUX2_X1 U9557 ( .A(n6673), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8049), .Z(
        P2_U3553) );
  OAI211_X1 U9558 ( .C1(n8052), .C2(n8051), .A(n9986), .B(n8050), .ZN(n8062)
         );
  NOR2_X1 U9559 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9659), .ZN(n8053) );
  AOI21_X1 U9560 ( .B1(n9987), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8053), .ZN(
        n8061) );
  NAND2_X1 U9561 ( .A1(n8150), .A2(n8054), .ZN(n8060) );
  AOI21_X1 U9562 ( .B1(n8057), .B2(n8056), .A(n8055), .ZN(n8058) );
  NAND2_X1 U9563 ( .A1(n9981), .A2(n8058), .ZN(n8059) );
  NAND4_X1 U9564 ( .A1(n8062), .A2(n8061), .A3(n8060), .A4(n8059), .ZN(
        P2_U3253) );
  OAI211_X1 U9565 ( .C1(n8065), .C2(n8064), .A(n9986), .B(n8063), .ZN(n8076)
         );
  INV_X1 U9566 ( .A(n8066), .ZN(n8067) );
  AOI21_X1 U9567 ( .B1(n9987), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8067), .ZN(
        n8075) );
  NAND2_X1 U9568 ( .A1(n8150), .A2(n8068), .ZN(n8074) );
  AOI21_X1 U9569 ( .B1(n8071), .B2(n8070), .A(n8069), .ZN(n8072) );
  NAND2_X1 U9570 ( .A1(n9981), .A2(n8072), .ZN(n8073) );
  NAND4_X1 U9571 ( .A1(n8076), .A2(n8075), .A3(n8074), .A4(n8073), .ZN(
        P2_U3254) );
  OAI211_X1 U9572 ( .C1(n8079), .C2(n8078), .A(n9986), .B(n8077), .ZN(n8088)
         );
  NOR2_X1 U9573 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9604), .ZN(n8080) );
  AOI21_X1 U9574 ( .B1(n9987), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n8080), .ZN(
        n8087) );
  NAND2_X1 U9575 ( .A1(n8150), .A2(n8081), .ZN(n8086) );
  AOI21_X1 U9576 ( .B1(n8083), .B2(n4332), .A(n8082), .ZN(n8084) );
  NAND2_X1 U9577 ( .A1(n9981), .A2(n8084), .ZN(n8085) );
  NAND4_X1 U9578 ( .A1(n8088), .A2(n8087), .A3(n8086), .A4(n8085), .ZN(
        P2_U3255) );
  NOR2_X1 U9579 ( .A1(n8090), .A2(n8089), .ZN(n8092) );
  NOR2_X1 U9580 ( .A1(n8092), .A2(n8091), .ZN(n8094) );
  INV_X1 U9581 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8531) );
  XNOR2_X1 U9582 ( .A(n8116), .B(n8531), .ZN(n8093) );
  NAND2_X1 U9583 ( .A1(n8093), .A2(n8094), .ZN(n8115) );
  OAI21_X1 U9584 ( .B1(n8094), .B2(n8093), .A(n8115), .ZN(n8095) );
  NAND2_X1 U9585 ( .A1(n8095), .A2(n9981), .ZN(n8108) );
  INV_X1 U9586 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8097) );
  OAI21_X1 U9587 ( .B1(n8157), .B2(n8097), .A(n8096), .ZN(n8098) );
  AOI21_X1 U9588 ( .B1(n8150), .B2(n8116), .A(n8098), .ZN(n8107) );
  NOR2_X1 U9589 ( .A1(n8100), .A2(n8099), .ZN(n8102) );
  NOR2_X1 U9590 ( .A1(n8102), .A2(n8101), .ZN(n8105) );
  MUX2_X1 U9591 ( .A(n8376), .B(P2_REG2_REG_16__SCAN_IN), .S(n8116), .Z(n8103)
         );
  INV_X1 U9592 ( .A(n8103), .ZN(n8104) );
  NAND2_X1 U9593 ( .A1(n8104), .A2(n8105), .ZN(n8109) );
  OAI211_X1 U9594 ( .C1(n8105), .C2(n8104), .A(n9986), .B(n8109), .ZN(n8106)
         );
  NAND3_X1 U9595 ( .A1(n8108), .A2(n8107), .A3(n8106), .ZN(P2_U3261) );
  NAND2_X1 U9596 ( .A1(n8116), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8110) );
  NAND2_X1 U9597 ( .A1(n8110), .A2(n8109), .ZN(n8113) );
  XNOR2_X1 U9598 ( .A(n8128), .B(n8111), .ZN(n8112) );
  NAND2_X1 U9599 ( .A1(n8112), .A2(n8113), .ZN(n8124) );
  OAI211_X1 U9600 ( .C1(n8113), .C2(n8112), .A(n9986), .B(n8124), .ZN(n8123)
         );
  NOR2_X1 U9601 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9661), .ZN(n8114) );
  AOI21_X1 U9602 ( .B1(n9987), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8114), .ZN(
        n8122) );
  NAND2_X1 U9603 ( .A1(n8150), .A2(n8128), .ZN(n8121) );
  XNOR2_X1 U9604 ( .A(n8128), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8118) );
  OAI21_X1 U9605 ( .B1(n8116), .B2(P2_REG1_REG_16__SCAN_IN), .A(n8115), .ZN(
        n8117) );
  NOR2_X1 U9606 ( .A1(n8118), .A2(n8117), .ZN(n8127) );
  AOI21_X1 U9607 ( .B1(n8118), .B2(n8117), .A(n8127), .ZN(n8119) );
  NAND2_X1 U9608 ( .A1(n9981), .A2(n8119), .ZN(n8120) );
  NAND4_X1 U9609 ( .A1(n8123), .A2(n8122), .A3(n8121), .A4(n8120), .ZN(
        P2_U3262) );
  NAND2_X1 U9610 ( .A1(n8128), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8125) );
  NAND2_X1 U9611 ( .A1(n8125), .A2(n8124), .ZN(n8140) );
  XNOR2_X1 U9612 ( .A(n8145), .B(n8140), .ZN(n8126) );
  NOR2_X1 U9613 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8126), .ZN(n8142) );
  AOI21_X1 U9614 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8126), .A(n8142), .ZN(
        n8139) );
  INV_X1 U9615 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8129) );
  AOI22_X1 U9616 ( .A1(n8145), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n8129), .B2(
        n8134), .ZN(n8130) );
  OAI21_X1 U9617 ( .B1(n8131), .B2(n8130), .A(n8144), .ZN(n8136) );
  NAND2_X1 U9618 ( .A1(n9987), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n8132) );
  OAI211_X1 U9619 ( .C1(n9982), .C2(n8134), .A(n8133), .B(n8132), .ZN(n8135)
         );
  AOI21_X1 U9620 ( .B1(n8136), .B2(n9981), .A(n8135), .ZN(n8137) );
  OAI21_X1 U9621 ( .B1(n8139), .B2(n8138), .A(n8137), .ZN(P2_U3263) );
  INV_X1 U9622 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8158) );
  NOR2_X1 U9623 ( .A1(n8145), .A2(n8140), .ZN(n8141) );
  NOR2_X1 U9624 ( .A1(n8142), .A2(n8141), .ZN(n8143) );
  XOR2_X1 U9625 ( .A(n8143), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8148) );
  AOI22_X1 U9626 ( .A1(n8148), .A2(n9986), .B1(n8146), .B2(n9981), .ZN(n8154)
         );
  INV_X1 U9627 ( .A(n8146), .ZN(n8151) );
  NOR2_X1 U9628 ( .A1(n8148), .A2(n8147), .ZN(n8149) );
  AOI211_X1 U9629 ( .C1(n9981), .C2(n8151), .A(n8150), .B(n8149), .ZN(n8153)
         );
  MUX2_X1 U9630 ( .A(n8154), .B(n8153), .S(n8152), .Z(n8156) );
  OAI211_X1 U9631 ( .C1(n8158), .C2(n8157), .A(n8156), .B(n8155), .ZN(P2_U3264) );
  INV_X1 U9632 ( .A(n9754), .ZN(n8164) );
  AND2_X1 U9633 ( .A1(n8160), .A2(n8159), .ZN(n9753) );
  NAND2_X1 U9634 ( .A1(n8438), .A2(n9753), .ZN(n8166) );
  OAI21_X1 U9635 ( .B1(n8161), .B2(n8438), .A(n8166), .ZN(n8162) );
  AOI21_X1 U9636 ( .B1(n9749), .B2(n8450), .A(n8162), .ZN(n8163) );
  OAI21_X1 U9637 ( .B1(n9747), .B2(n8446), .A(n8163), .ZN(P2_U3265) );
  OAI21_X1 U9638 ( .B1(n8165), .B2(n8164), .A(n4314), .ZN(n9751) );
  INV_X1 U9639 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8167) );
  OAI21_X1 U9640 ( .B1(n8438), .B2(n8167), .A(n8166), .ZN(n8168) );
  AOI21_X1 U9641 ( .B1(n9754), .B2(n8450), .A(n8168), .ZN(n8169) );
  OAI21_X1 U9642 ( .B1(n9751), .B2(n8446), .A(n8169), .ZN(P2_U3266) );
  OAI21_X1 U9643 ( .B1(n8171), .B2(n8178), .A(n8170), .ZN(n8172) );
  INV_X1 U9644 ( .A(n8172), .ZN(n8463) );
  AOI21_X1 U9645 ( .B1(n8459), .B2(n4877), .A(n8173), .ZN(n8460) );
  INV_X1 U9646 ( .A(n8459), .ZN(n8177) );
  INV_X1 U9647 ( .A(n8174), .ZN(n8175) );
  AOI22_X1 U9648 ( .A1(n8175), .A2(n8404), .B1(n8406), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8176) );
  OAI21_X1 U9649 ( .B1(n8177), .B2(n8408), .A(n8176), .ZN(n8184) );
  XNOR2_X1 U9650 ( .A(n8179), .B(n8178), .ZN(n8182) );
  AOI222_X1 U9651 ( .A1(n8434), .A2(n8182), .B1(n8181), .B2(n8343), .C1(n8180), 
        .C2(n8341), .ZN(n8462) );
  NOR2_X1 U9652 ( .A1(n8462), .A2(n8406), .ZN(n8183) );
  AOI211_X1 U9653 ( .C1(n8460), .C2(n8420), .A(n8184), .B(n8183), .ZN(n8185)
         );
  OAI21_X1 U9654 ( .B1(n8463), .B2(n8422), .A(n8185), .ZN(P2_U3268) );
  OAI21_X1 U9655 ( .B1(n8187), .B2(n8194), .A(n8186), .ZN(n8188) );
  INV_X1 U9656 ( .A(n8188), .ZN(n8468) );
  INV_X1 U9657 ( .A(n4877), .ZN(n8189) );
  AOI21_X1 U9658 ( .B1(n8464), .B2(n8211), .A(n8189), .ZN(n8465) );
  AOI22_X1 U9659 ( .A1(n8406), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8190), .B2(
        n8404), .ZN(n8191) );
  OAI21_X1 U9660 ( .B1(n8192), .B2(n8408), .A(n8191), .ZN(n8201) );
  INV_X1 U9661 ( .A(n8193), .ZN(n8195) );
  AOI21_X1 U9662 ( .B1(n8195), .B2(n8194), .A(n8410), .ZN(n8199) );
  OAI22_X1 U9663 ( .A1(n8196), .A2(n8430), .B1(n8226), .B2(n6188), .ZN(n8197)
         );
  AOI21_X1 U9664 ( .B1(n8199), .B2(n8198), .A(n8197), .ZN(n8467) );
  NOR2_X1 U9665 ( .A1(n8467), .A2(n8406), .ZN(n8200) );
  AOI211_X1 U9666 ( .C1(n8420), .C2(n8465), .A(n8201), .B(n8200), .ZN(n8202)
         );
  OAI21_X1 U9667 ( .B1(n8468), .B2(n8422), .A(n8202), .ZN(P2_U3269) );
  OAI21_X1 U9668 ( .B1(n8204), .B2(n8208), .A(n8203), .ZN(n8205) );
  INV_X1 U9669 ( .A(n8205), .ZN(n8473) );
  AOI21_X1 U9670 ( .B1(n8208), .B2(n8207), .A(n8206), .ZN(n8209) );
  OAI222_X1 U9671 ( .A1(n8430), .A2(n8210), .B1(n6188), .B2(n8245), .C1(n8410), 
        .C2(n8209), .ZN(n8469) );
  INV_X1 U9672 ( .A(n8227), .ZN(n8213) );
  INV_X1 U9673 ( .A(n8211), .ZN(n8212) );
  AOI211_X1 U9674 ( .C1(n8471), .C2(n8213), .A(n10050), .B(n8212), .ZN(n8470)
         );
  NAND2_X1 U9675 ( .A1(n8470), .A2(n8358), .ZN(n8216) );
  AOI22_X1 U9676 ( .A1(n8406), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8214), .B2(
        n8404), .ZN(n8215) );
  OAI211_X1 U9677 ( .C1(n8217), .C2(n8408), .A(n8216), .B(n8215), .ZN(n8218)
         );
  AOI21_X1 U9678 ( .B1(n8469), .B2(n8438), .A(n8218), .ZN(n8219) );
  OAI21_X1 U9679 ( .B1(n8473), .B2(n8422), .A(n8219), .ZN(P2_U3270) );
  OAI21_X1 U9680 ( .B1(n8221), .B2(n8224), .A(n8220), .ZN(n8222) );
  INV_X1 U9681 ( .A(n8222), .ZN(n8478) );
  XNOR2_X1 U9682 ( .A(n8223), .B(n8224), .ZN(n8225) );
  OAI222_X1 U9683 ( .A1(n8430), .A2(n8226), .B1(n6188), .B2(n8258), .C1(n8410), 
        .C2(n8225), .ZN(n8474) );
  INV_X1 U9684 ( .A(n8476), .ZN(n8232) );
  AOI211_X1 U9685 ( .C1(n8476), .C2(n8236), .A(n10050), .B(n8227), .ZN(n8475)
         );
  NAND2_X1 U9686 ( .A1(n8475), .A2(n8358), .ZN(n8231) );
  INV_X1 U9687 ( .A(n8228), .ZN(n8229) );
  AOI22_X1 U9688 ( .A1(n8406), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8229), .B2(
        n8404), .ZN(n8230) );
  OAI211_X1 U9689 ( .C1(n8232), .C2(n8408), .A(n8231), .B(n8230), .ZN(n8233)
         );
  AOI21_X1 U9690 ( .B1(n8474), .B2(n8438), .A(n8233), .ZN(n8234) );
  OAI21_X1 U9691 ( .B1(n8478), .B2(n8422), .A(n8234), .ZN(P2_U3271) );
  XNOR2_X1 U9692 ( .A(n8235), .B(n8243), .ZN(n8483) );
  INV_X1 U9693 ( .A(n8236), .ZN(n8237) );
  AOI21_X1 U9694 ( .B1(n8479), .B2(n4324), .A(n8237), .ZN(n8480) );
  INV_X1 U9695 ( .A(n8479), .ZN(n8241) );
  INV_X1 U9696 ( .A(n8238), .ZN(n8239) );
  AOI22_X1 U9697 ( .A1(n8406), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8239), .B2(
        n8404), .ZN(n8240) );
  OAI21_X1 U9698 ( .B1(n8241), .B2(n8408), .A(n8240), .ZN(n8250) );
  NOR2_X1 U9699 ( .A1(n8242), .A2(n8410), .ZN(n8248) );
  OAI21_X1 U9700 ( .B1(n8256), .B2(n8244), .A(n8243), .ZN(n8247) );
  OAI22_X1 U9701 ( .A1(n8245), .A2(n8430), .B1(n8284), .B2(n6188), .ZN(n8246)
         );
  AOI21_X1 U9702 ( .B1(n8248), .B2(n8247), .A(n8246), .ZN(n8482) );
  NOR2_X1 U9703 ( .A1(n8482), .A2(n8406), .ZN(n8249) );
  AOI211_X1 U9704 ( .C1(n8480), .C2(n8420), .A(n8250), .B(n8249), .ZN(n8251)
         );
  OAI21_X1 U9705 ( .B1(n8422), .B2(n8483), .A(n8251), .ZN(P2_U3272) );
  AOI21_X1 U9706 ( .B1(n8253), .B2(n8254), .A(n8261), .ZN(n8255) );
  OR2_X1 U9707 ( .A1(n8256), .A2(n8255), .ZN(n8260) );
  OAI22_X1 U9708 ( .A1(n8258), .A2(n8430), .B1(n8257), .B2(n6188), .ZN(n8259)
         );
  AOI21_X1 U9709 ( .B1(n8260), .B2(n8434), .A(n8259), .ZN(n8487) );
  NAND2_X1 U9710 ( .A1(n8262), .A2(n8261), .ZN(n8263) );
  NAND2_X1 U9711 ( .A1(n8489), .A2(n8265), .ZN(n8272) );
  NAND2_X1 U9712 ( .A1(n8494), .A2(n8484), .ZN(n8266) );
  AND2_X1 U9713 ( .A1(n4324), .A2(n8266), .ZN(n8485) );
  AOI22_X1 U9714 ( .A1(n8406), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8267), .B2(
        n8404), .ZN(n8268) );
  OAI21_X1 U9715 ( .B1(n8269), .B2(n8408), .A(n8268), .ZN(n8270) );
  AOI21_X1 U9716 ( .B1(n8485), .B2(n8420), .A(n8270), .ZN(n8271) );
  OAI211_X1 U9717 ( .C1(n8406), .C2(n8487), .A(n8272), .B(n8271), .ZN(P2_U3273) );
  XNOR2_X1 U9718 ( .A(n8273), .B(n6036), .ZN(n8498) );
  OAI22_X1 U9719 ( .A1(n8438), .A2(n8275), .B1(n8274), .B2(n8440), .ZN(n8278)
         );
  NOR2_X1 U9720 ( .A1(n8291), .A2(n8276), .ZN(n8492) );
  NOR3_X1 U9721 ( .A1(n8492), .A2(n4607), .A3(n8446), .ZN(n8277) );
  AOI211_X1 U9722 ( .C1(n8450), .C2(n8493), .A(n8278), .B(n8277), .ZN(n8288)
         );
  INV_X1 U9723 ( .A(n8253), .ZN(n8282) );
  AOI21_X1 U9724 ( .B1(n8296), .B2(n8280), .A(n8279), .ZN(n8281) );
  NOR3_X1 U9725 ( .A1(n8282), .A2(n8281), .A3(n8410), .ZN(n8286) );
  OAI22_X1 U9726 ( .A1(n8284), .A2(n8430), .B1(n8283), .B2(n6188), .ZN(n8285)
         );
  NOR2_X1 U9727 ( .A1(n8286), .A2(n8285), .ZN(n8497) );
  OR2_X1 U9728 ( .A1(n8497), .A2(n8406), .ZN(n8287) );
  OAI211_X1 U9729 ( .C1(n8498), .C2(n8422), .A(n8288), .B(n8287), .ZN(P2_U3274) );
  XNOR2_X1 U9730 ( .A(n8290), .B(n8289), .ZN(n8503) );
  INV_X1 U9731 ( .A(n8305), .ZN(n8292) );
  AOI21_X1 U9732 ( .B1(n8499), .B2(n8292), .A(n8291), .ZN(n8500) );
  AOI22_X1 U9733 ( .A1(n8406), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8293), .B2(
        n8404), .ZN(n8294) );
  OAI21_X1 U9734 ( .B1(n8295), .B2(n8408), .A(n8294), .ZN(n8300) );
  OAI21_X1 U9735 ( .B1(n4340), .B2(n4698), .A(n8296), .ZN(n8298) );
  AOI222_X1 U9736 ( .A1(n8434), .A2(n8298), .B1(n8297), .B2(n8343), .C1(n4560), 
        .C2(n8341), .ZN(n8502) );
  NOR2_X1 U9737 ( .A1(n8502), .A2(n8406), .ZN(n8299) );
  AOI211_X1 U9738 ( .C1(n8500), .C2(n8420), .A(n8300), .B(n8299), .ZN(n8301)
         );
  OAI21_X1 U9739 ( .B1(n8422), .B2(n8503), .A(n8301), .ZN(P2_U3275) );
  OAI21_X1 U9740 ( .B1(n8304), .B2(n8303), .A(n8302), .ZN(n8508) );
  AOI21_X1 U9741 ( .B1(n8504), .B2(n8306), .A(n8305), .ZN(n8505) );
  AOI22_X1 U9742 ( .A1(n8406), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8307), .B2(
        n8404), .ZN(n8308) );
  OAI21_X1 U9743 ( .B1(n4561), .B2(n8408), .A(n8308), .ZN(n8314) );
  NAND2_X1 U9744 ( .A1(n8324), .A2(n8309), .ZN(n8310) );
  XNOR2_X1 U9745 ( .A(n8310), .B(n4824), .ZN(n8312) );
  AOI222_X1 U9746 ( .A1(n8434), .A2(n8312), .B1(n8344), .B2(n8341), .C1(n8311), 
        .C2(n8343), .ZN(n8507) );
  NOR2_X1 U9747 ( .A1(n8507), .A2(n8406), .ZN(n8313) );
  AOI211_X1 U9748 ( .C1(n8505), .C2(n8420), .A(n8314), .B(n8313), .ZN(n8315)
         );
  OAI21_X1 U9749 ( .B1(n8422), .B2(n8508), .A(n8315), .ZN(P2_U3276) );
  OAI21_X1 U9750 ( .B1(n8318), .B2(n8317), .A(n8316), .ZN(n8513) );
  XNOR2_X1 U9751 ( .A(n8319), .B(n8510), .ZN(n8320) );
  NOR2_X1 U9752 ( .A1(n8320), .A2(n10050), .ZN(n8509) );
  INV_X1 U9753 ( .A(n8510), .ZN(n8323) );
  AOI22_X1 U9754 ( .A1(n8406), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8321), .B2(
        n8404), .ZN(n8322) );
  OAI21_X1 U9755 ( .B1(n8323), .B2(n8408), .A(n8322), .ZN(n8330) );
  OAI21_X1 U9756 ( .B1(n8326), .B2(n8325), .A(n8324), .ZN(n8328) );
  AOI222_X1 U9757 ( .A1(n8434), .A2(n8328), .B1(n4560), .B2(n8343), .C1(n8327), 
        .C2(n8341), .ZN(n8512) );
  NOR2_X1 U9758 ( .A1(n8512), .A2(n8406), .ZN(n8329) );
  AOI211_X1 U9759 ( .C1(n8509), .C2(n8358), .A(n8330), .B(n8329), .ZN(n8331)
         );
  OAI21_X1 U9760 ( .B1(n8422), .B2(n8513), .A(n8331), .ZN(P2_U3277) );
  XNOR2_X1 U9761 ( .A(n8332), .B(n8339), .ZN(n8518) );
  INV_X1 U9762 ( .A(n8356), .ZN(n8334) );
  INV_X1 U9763 ( .A(n8319), .ZN(n8333) );
  AOI21_X1 U9764 ( .B1(n8514), .B2(n8334), .A(n8333), .ZN(n8515) );
  AOI22_X1 U9765 ( .A1(n8406), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8335), .B2(
        n8404), .ZN(n8336) );
  OAI21_X1 U9766 ( .B1(n8337), .B2(n8408), .A(n8336), .ZN(n8347) );
  OAI21_X1 U9767 ( .B1(n8340), .B2(n8339), .A(n8338), .ZN(n8345) );
  AOI222_X1 U9768 ( .A1(n8434), .A2(n8345), .B1(n8344), .B2(n8343), .C1(n8342), 
        .C2(n8341), .ZN(n8517) );
  NOR2_X1 U9769 ( .A1(n8517), .A2(n8406), .ZN(n8346) );
  AOI211_X1 U9770 ( .C1(n8515), .C2(n8420), .A(n8347), .B(n8346), .ZN(n8348)
         );
  OAI21_X1 U9771 ( .B1(n8518), .B2(n8422), .A(n8348), .ZN(P2_U3278) );
  INV_X1 U9772 ( .A(n8349), .ZN(n8350) );
  AOI21_X1 U9773 ( .B1(n8352), .B2(n8351), .A(n8350), .ZN(n8523) );
  XNOR2_X1 U9774 ( .A(n8353), .B(n5978), .ZN(n8354) );
  OAI222_X1 U9775 ( .A1(n6188), .A2(n8393), .B1(n8430), .B2(n8355), .C1(n8354), 
        .C2(n8410), .ZN(n8519) );
  INV_X1 U9776 ( .A(n8377), .ZN(n8357) );
  AOI211_X1 U9777 ( .C1(n8521), .C2(n8357), .A(n10050), .B(n8356), .ZN(n8520)
         );
  NAND2_X1 U9778 ( .A1(n8520), .A2(n8358), .ZN(n8361) );
  AOI22_X1 U9779 ( .A1(n8406), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8359), .B2(
        n8404), .ZN(n8360) );
  OAI211_X1 U9780 ( .C1(n8362), .C2(n8408), .A(n8361), .B(n8360), .ZN(n8363)
         );
  AOI21_X1 U9781 ( .B1(n8519), .B2(n8438), .A(n8363), .ZN(n8364) );
  OAI21_X1 U9782 ( .B1(n8523), .B2(n8422), .A(n8364), .ZN(P2_U3279) );
  OAI21_X1 U9783 ( .B1(n8366), .B2(n8367), .A(n8365), .ZN(n8528) );
  OR2_X1 U9784 ( .A1(n8528), .A2(n8427), .ZN(n8373) );
  XNOR2_X1 U9785 ( .A(n8368), .B(n8367), .ZN(n8371) );
  OAI22_X1 U9786 ( .A1(n8413), .A2(n6188), .B1(n8369), .B2(n8430), .ZN(n8370)
         );
  AOI21_X1 U9787 ( .B1(n8371), .B2(n8434), .A(n8370), .ZN(n8372) );
  NAND2_X1 U9788 ( .A1(n8373), .A2(n8372), .ZN(n8530) );
  NAND2_X1 U9789 ( .A1(n8530), .A2(n8438), .ZN(n8382) );
  INV_X1 U9790 ( .A(n8374), .ZN(n8375) );
  OAI22_X1 U9791 ( .A1(n8438), .A2(n8376), .B1(n8375), .B2(n8440), .ZN(n8380)
         );
  AND2_X1 U9792 ( .A1(n8386), .A2(n8524), .ZN(n8378) );
  OR2_X1 U9793 ( .A1(n8378), .A2(n8377), .ZN(n8525) );
  NOR2_X1 U9794 ( .A1(n8525), .A2(n8446), .ZN(n8379) );
  AOI211_X1 U9795 ( .C1(n8450), .C2(n8524), .A(n8380), .B(n8379), .ZN(n8381)
         );
  OAI211_X1 U9796 ( .C1(n8528), .C2(n8453), .A(n8382), .B(n8381), .ZN(P2_U3280) );
  OAI21_X1 U9797 ( .B1(n8384), .B2(n8391), .A(n8383), .ZN(n8385) );
  INV_X1 U9798 ( .A(n8385), .ZN(n8537) );
  AOI21_X1 U9799 ( .B1(n8533), .B2(n8402), .A(n4604), .ZN(n8534) );
  INV_X1 U9800 ( .A(n8533), .ZN(n8389) );
  AOI22_X1 U9801 ( .A1(n8406), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8387), .B2(
        n8404), .ZN(n8388) );
  OAI21_X1 U9802 ( .B1(n8389), .B2(n8408), .A(n8388), .ZN(n8398) );
  INV_X1 U9803 ( .A(n8390), .ZN(n8392) );
  AOI21_X1 U9804 ( .B1(n8392), .B2(n8391), .A(n8410), .ZN(n8396) );
  OAI22_X1 U9805 ( .A1(n8431), .A2(n6188), .B1(n8393), .B2(n8430), .ZN(n8394)
         );
  AOI21_X1 U9806 ( .B1(n8396), .B2(n8395), .A(n8394), .ZN(n8536) );
  NOR2_X1 U9807 ( .A1(n8536), .A2(n8406), .ZN(n8397) );
  AOI211_X1 U9808 ( .C1(n8534), .C2(n8420), .A(n8398), .B(n8397), .ZN(n8399)
         );
  OAI21_X1 U9809 ( .B1(n8537), .B2(n8422), .A(n8399), .ZN(P2_U3281) );
  NAND2_X1 U9810 ( .A1(n8426), .A2(n8400), .ZN(n8401) );
  XNOR2_X1 U9811 ( .A(n8401), .B(n8411), .ZN(n8543) );
  INV_X1 U9812 ( .A(n8445), .ZN(n8403) );
  AOI21_X1 U9813 ( .B1(n8538), .B2(n8403), .A(n4599), .ZN(n8540) );
  AOI22_X1 U9814 ( .A1(n8406), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8405), .B2(
        n8404), .ZN(n8407) );
  OAI21_X1 U9815 ( .B1(n8409), .B2(n8408), .A(n8407), .ZN(n8419) );
  AOI21_X1 U9816 ( .B1(n8412), .B2(n8411), .A(n8410), .ZN(n8417) );
  OAI22_X1 U9817 ( .A1(n8414), .A2(n6188), .B1(n8413), .B2(n8430), .ZN(n8415)
         );
  AOI21_X1 U9818 ( .B1(n8417), .B2(n8416), .A(n8415), .ZN(n8542) );
  NOR2_X1 U9819 ( .A1(n8542), .A2(n8406), .ZN(n8418) );
  AOI211_X1 U9820 ( .C1(n8540), .C2(n8420), .A(n8419), .B(n8418), .ZN(n8421)
         );
  OAI21_X1 U9821 ( .B1(n8422), .B2(n8543), .A(n8421), .ZN(P2_U3282) );
  NAND2_X1 U9822 ( .A1(n8424), .A2(n8423), .ZN(n8425) );
  NAND2_X1 U9823 ( .A1(n8426), .A2(n8425), .ZN(n8548) );
  OR2_X1 U9824 ( .A1(n8548), .A2(n8427), .ZN(n8437) );
  XNOR2_X1 U9825 ( .A(n8429), .B(n8428), .ZN(n8435) );
  OAI22_X1 U9826 ( .A1(n8432), .A2(n6188), .B1(n8431), .B2(n8430), .ZN(n8433)
         );
  AOI21_X1 U9827 ( .B1(n8435), .B2(n8434), .A(n8433), .ZN(n8436) );
  NAND2_X1 U9828 ( .A1(n8437), .A2(n8436), .ZN(n8550) );
  NAND2_X1 U9829 ( .A1(n8550), .A2(n8438), .ZN(n8452) );
  INV_X1 U9830 ( .A(n8439), .ZN(n8441) );
  OAI22_X1 U9831 ( .A1(n8438), .A2(n8442), .B1(n8441), .B2(n8440), .ZN(n8448)
         );
  NOR2_X1 U9832 ( .A1(n8443), .A2(n8544), .ZN(n8444) );
  OR2_X1 U9833 ( .A1(n8445), .A2(n8444), .ZN(n8545) );
  NOR2_X1 U9834 ( .A1(n8545), .A2(n8446), .ZN(n8447) );
  AOI211_X1 U9835 ( .C1(n8450), .C2(n8449), .A(n8448), .B(n8447), .ZN(n8451)
         );
  OAI211_X1 U9836 ( .C1(n8548), .C2(n8453), .A(n8452), .B(n8451), .ZN(P2_U3283) );
  AOI21_X1 U9837 ( .B1(n10045), .B2(n8455), .A(n8454), .ZN(n8456) );
  MUX2_X1 U9838 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8563), .S(n10069), .Z(
        P2_U3549) );
  AOI22_X1 U9839 ( .A1(n8460), .A2(n8539), .B1(n10045), .B2(n8459), .ZN(n8461)
         );
  OAI211_X1 U9840 ( .C1(n8463), .C2(n10028), .A(n8462), .B(n8461), .ZN(n8564)
         );
  MUX2_X1 U9841 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8564), .S(n10069), .Z(
        P2_U3548) );
  AOI22_X1 U9842 ( .A1(n8465), .A2(n8539), .B1(n10045), .B2(n8464), .ZN(n8466)
         );
  OAI211_X1 U9843 ( .C1(n8468), .C2(n10028), .A(n8467), .B(n8466), .ZN(n8565)
         );
  MUX2_X1 U9844 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8565), .S(n10069), .Z(
        P2_U3547) );
  AOI211_X1 U9845 ( .C1(n10045), .C2(n8471), .A(n8470), .B(n8469), .ZN(n8472)
         );
  OAI21_X1 U9846 ( .B1(n10028), .B2(n8473), .A(n8472), .ZN(n8566) );
  MUX2_X1 U9847 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8566), .S(n10069), .Z(
        P2_U3546) );
  AOI211_X1 U9848 ( .C1(n10045), .C2(n8476), .A(n8475), .B(n8474), .ZN(n8477)
         );
  OAI21_X1 U9849 ( .B1(n10028), .B2(n8478), .A(n8477), .ZN(n8567) );
  MUX2_X1 U9850 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8567), .S(n10069), .Z(
        P2_U3545) );
  AOI22_X1 U9851 ( .A1(n8480), .A2(n8539), .B1(n10045), .B2(n8479), .ZN(n8481)
         );
  OAI211_X1 U9852 ( .C1(n8483), .C2(n10028), .A(n8482), .B(n8481), .ZN(n8568)
         );
  MUX2_X1 U9853 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8568), .S(n10069), .Z(
        P2_U3544) );
  INV_X1 U9854 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8490) );
  AOI22_X1 U9855 ( .A1(n8485), .A2(n8539), .B1(n10045), .B2(n8484), .ZN(n8486)
         );
  NAND2_X1 U9856 ( .A1(n8487), .A2(n8486), .ZN(n8488) );
  AOI21_X1 U9857 ( .B1(n8489), .B2(n10052), .A(n8488), .ZN(n8569) );
  MUX2_X1 U9858 ( .A(n8490), .B(n8569), .S(n10069), .Z(n8491) );
  INV_X1 U9859 ( .A(n8491), .ZN(P2_U3543) );
  NOR2_X1 U9860 ( .A1(n8492), .A2(n10050), .ZN(n8495) );
  AOI22_X1 U9861 ( .A1(n8495), .A2(n8494), .B1(n10045), .B2(n8493), .ZN(n8496)
         );
  OAI211_X1 U9862 ( .C1(n8498), .C2(n10028), .A(n8497), .B(n8496), .ZN(n8572)
         );
  MUX2_X1 U9863 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8572), .S(n10069), .Z(
        P2_U3542) );
  AOI22_X1 U9864 ( .A1(n8500), .A2(n8539), .B1(n10045), .B2(n8499), .ZN(n8501)
         );
  OAI211_X1 U9865 ( .C1(n8503), .C2(n10028), .A(n8502), .B(n8501), .ZN(n8573)
         );
  MUX2_X1 U9866 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8573), .S(n10069), .Z(
        P2_U3541) );
  AOI22_X1 U9867 ( .A1(n8505), .A2(n8539), .B1(n10045), .B2(n8504), .ZN(n8506)
         );
  OAI211_X1 U9868 ( .C1(n8508), .C2(n10028), .A(n8507), .B(n8506), .ZN(n8574)
         );
  MUX2_X1 U9869 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8574), .S(n10069), .Z(
        P2_U3540) );
  AOI21_X1 U9870 ( .B1(n10045), .B2(n8510), .A(n8509), .ZN(n8511) );
  OAI211_X1 U9871 ( .C1(n8513), .C2(n10028), .A(n8512), .B(n8511), .ZN(n8575)
         );
  MUX2_X1 U9872 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8575), .S(n10069), .Z(
        P2_U3539) );
  AOI22_X1 U9873 ( .A1(n8515), .A2(n8539), .B1(n10045), .B2(n8514), .ZN(n8516)
         );
  OAI211_X1 U9874 ( .C1(n8518), .C2(n10028), .A(n8517), .B(n8516), .ZN(n8576)
         );
  MUX2_X1 U9875 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8576), .S(n10069), .Z(
        P2_U3538) );
  AOI211_X1 U9876 ( .C1(n10045), .C2(n8521), .A(n8520), .B(n8519), .ZN(n8522)
         );
  OAI21_X1 U9877 ( .B1(n8523), .B2(n10028), .A(n8522), .ZN(n8577) );
  MUX2_X1 U9878 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8577), .S(n10069), .Z(
        P2_U3537) );
  INV_X1 U9879 ( .A(n10045), .ZN(n10038) );
  OAI22_X1 U9880 ( .A1(n8525), .A2(n10050), .B1(n4603), .B2(n10038), .ZN(n8526) );
  INV_X1 U9881 ( .A(n8526), .ZN(n8527) );
  OAI21_X1 U9882 ( .B1(n8528), .B2(n10031), .A(n8527), .ZN(n8529) );
  NOR2_X1 U9883 ( .A1(n8530), .A2(n8529), .ZN(n8578) );
  MUX2_X1 U9884 ( .A(n8531), .B(n8578), .S(n10069), .Z(n8532) );
  INV_X1 U9885 ( .A(n8532), .ZN(P2_U3536) );
  AOI22_X1 U9886 ( .A1(n8534), .A2(n8539), .B1(n10045), .B2(n8533), .ZN(n8535)
         );
  OAI211_X1 U9887 ( .C1(n8537), .C2(n10028), .A(n8536), .B(n8535), .ZN(n8581)
         );
  MUX2_X1 U9888 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8581), .S(n10069), .Z(
        P2_U3535) );
  AOI22_X1 U9889 ( .A1(n8540), .A2(n8539), .B1(n10045), .B2(n8538), .ZN(n8541)
         );
  OAI211_X1 U9890 ( .C1(n8543), .C2(n10028), .A(n8542), .B(n8541), .ZN(n8582)
         );
  MUX2_X1 U9891 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8582), .S(n10069), .Z(
        P2_U3534) );
  OAI22_X1 U9892 ( .A1(n8545), .A2(n10050), .B1(n8544), .B2(n10038), .ZN(n8546) );
  INV_X1 U9893 ( .A(n8546), .ZN(n8547) );
  OAI21_X1 U9894 ( .B1(n8548), .B2(n10031), .A(n8547), .ZN(n8549) );
  NOR2_X1 U9895 ( .A1(n8550), .A2(n8549), .ZN(n8584) );
  MUX2_X1 U9896 ( .A(n8584), .B(n8551), .S(n10067), .Z(n8552) );
  INV_X1 U9897 ( .A(n8552), .ZN(P2_U3533) );
  AOI211_X1 U9898 ( .C1(n10045), .C2(n8555), .A(n8554), .B(n8553), .ZN(n8556)
         );
  OAI21_X1 U9899 ( .B1(n8557), .B2(n10028), .A(n8556), .ZN(n8586) );
  MUX2_X1 U9900 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n8586), .S(n10069), .Z(
        P2_U3531) );
  AOI21_X1 U9901 ( .B1(n10045), .B2(n8559), .A(n8558), .ZN(n8560) );
  OAI211_X1 U9902 ( .C1(n8562), .C2(n10031), .A(n8561), .B(n8560), .ZN(n8587)
         );
  MUX2_X1 U9903 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n8587), .S(n10069), .Z(
        P2_U3529) );
  MUX2_X1 U9904 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8563), .S(n10055), .Z(
        P2_U3517) );
  MUX2_X1 U9905 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8564), .S(n10055), .Z(
        P2_U3516) );
  MUX2_X1 U9906 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8565), .S(n10055), .Z(
        P2_U3515) );
  MUX2_X1 U9907 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8566), .S(n10055), .Z(
        P2_U3514) );
  MUX2_X1 U9908 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8567), .S(n10055), .Z(
        P2_U3513) );
  MUX2_X1 U9909 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8568), .S(n10055), .Z(
        P2_U3512) );
  INV_X1 U9910 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8570) );
  MUX2_X1 U9911 ( .A(n8570), .B(n8569), .S(n10055), .Z(n8571) );
  INV_X1 U9912 ( .A(n8571), .ZN(P2_U3511) );
  MUX2_X1 U9913 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8572), .S(n10055), .Z(
        P2_U3510) );
  MUX2_X1 U9914 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8573), .S(n10055), .Z(
        P2_U3509) );
  MUX2_X1 U9915 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8574), .S(n10055), .Z(
        P2_U3508) );
  MUX2_X1 U9916 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8575), .S(n10055), .Z(
        P2_U3507) );
  MUX2_X1 U9917 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8576), .S(n10055), .Z(
        P2_U3505) );
  MUX2_X1 U9918 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8577), .S(n10055), .Z(
        P2_U3502) );
  MUX2_X1 U9919 ( .A(n8579), .B(n8578), .S(n10055), .Z(n8580) );
  INV_X1 U9920 ( .A(n8580), .ZN(P2_U3499) );
  MUX2_X1 U9921 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8581), .S(n10055), .Z(
        P2_U3496) );
  MUX2_X1 U9922 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8582), .S(n10055), .Z(
        P2_U3493) );
  MUX2_X1 U9923 ( .A(n8584), .B(n8583), .S(n10054), .Z(n8585) );
  INV_X1 U9924 ( .A(n8585), .ZN(P2_U3490) );
  MUX2_X1 U9925 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n8586), .S(n10055), .Z(
        P2_U3484) );
  MUX2_X1 U9926 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n8587), .S(n10055), .Z(
        P2_U3478) );
  INV_X1 U9927 ( .A(n8836), .ZN(n9513) );
  NOR4_X1 U9928 ( .A1(n4848), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8588), .A4(
        P2_U3152), .ZN(n8589) );
  AOI21_X1 U9929 ( .B1(n8594), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8589), .ZN(
        n8590) );
  OAI21_X1 U9930 ( .B1(n9513), .B2(n8597), .A(n8590), .ZN(P2_U3327) );
  AOI22_X1 U9931 ( .A1(n8591), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8594), .ZN(n8592) );
  OAI21_X1 U9932 ( .B1(n8593), .B2(n8597), .A(n8592), .ZN(P2_U3328) );
  AOI22_X1 U9933 ( .A1(n8595), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8594), .ZN(n8596) );
  OAI21_X1 U9934 ( .B1(n8598), .B2(n8597), .A(n8596), .ZN(P2_U3329) );
  MUX2_X1 U9935 ( .A(n8599), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U9936 ( .A(n8679), .ZN(n8603) );
  AOI21_X1 U9937 ( .B1(n8601), .B2(n8678), .A(n8600), .ZN(n8602) );
  AOI21_X1 U9938 ( .B1(n8603), .B2(n8678), .A(n8602), .ZN(n8608) );
  NAND2_X1 U9939 ( .A1(n9120), .A2(n8734), .ZN(n8605) );
  AOI22_X1 U9940 ( .A1(n9114), .A2(n8708), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8604) );
  OAI211_X1 U9941 ( .C1(n8736), .C2(n9253), .A(n8605), .B(n8604), .ZN(n8606)
         );
  AOI21_X1 U9942 ( .B1(n9444), .B2(n8738), .A(n8606), .ZN(n8607) );
  OAI21_X1 U9943 ( .B1(n8608), .B2(n8740), .A(n8607), .ZN(P1_U3214) );
  OAI21_X1 U9944 ( .B1(n8610), .B2(n4367), .A(n8609), .ZN(n8611) );
  NAND2_X1 U9945 ( .A1(n8611), .A2(n8717), .ZN(n8615) );
  NAND2_X1 U9946 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9091) );
  OAI21_X1 U9947 ( .B1(n8720), .B2(n9284), .A(n9091), .ZN(n8613) );
  NOR2_X1 U9948 ( .A1(n8736), .A2(n9315), .ZN(n8612) );
  AOI211_X1 U9949 ( .C1(n8708), .C2(n9322), .A(n8613), .B(n8612), .ZN(n8614)
         );
  OAI211_X1 U9950 ( .C1(n9319), .C2(n8726), .A(n8615), .B(n8614), .ZN(P1_U3217) );
  NAND2_X1 U9951 ( .A1(n8616), .A2(n8840), .ZN(n8619) );
  OR2_X1 U9952 ( .A1(n5057), .A2(n8617), .ZN(n8618) );
  NAND2_X1 U9953 ( .A1(n9421), .A2(n8620), .ZN(n8622) );
  NAND2_X1 U9954 ( .A1(n9157), .A2(n5215), .ZN(n8621) );
  NAND2_X1 U9955 ( .A1(n8622), .A2(n8621), .ZN(n8623) );
  XNOR2_X1 U9956 ( .A(n8623), .B(n5031), .ZN(n8627) );
  NAND2_X1 U9957 ( .A1(n9421), .A2(n5215), .ZN(n8624) );
  OAI21_X1 U9958 ( .B1(n9192), .B2(n8625), .A(n8624), .ZN(n8626) );
  XNOR2_X1 U9959 ( .A(n8627), .B(n8626), .ZN(n8628) );
  INV_X1 U9960 ( .A(n8628), .ZN(n8639) );
  NAND3_X1 U9961 ( .A1(n8639), .A2(n8717), .A3(n8638), .ZN(n8644) );
  NAND3_X1 U9962 ( .A1(n8645), .A2(n8717), .A3(n8628), .ZN(n8643) );
  INV_X1 U9963 ( .A(n8629), .ZN(n9181) );
  AOI22_X1 U9964 ( .A1(n9181), .A2(n8723), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8637) );
  OR2_X1 U9965 ( .A1(n9162), .A2(n5012), .ZN(n8635) );
  INV_X1 U9966 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8632) );
  NAND2_X1 U9967 ( .A1(n5477), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8631) );
  NAND2_X1 U9968 ( .A1(n8830), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8630) );
  OAI211_X1 U9969 ( .C1(n8632), .C2(n5685), .A(n8631), .B(n8630), .ZN(n8633)
         );
  INV_X1 U9970 ( .A(n8633), .ZN(n8634) );
  NAND2_X1 U9971 ( .A1(n8635), .A2(n8634), .ZN(n9012) );
  NAND2_X1 U9972 ( .A1(n9012), .A2(n8734), .ZN(n8636) );
  OAI211_X1 U9973 ( .C1(n9210), .C2(n8732), .A(n8637), .B(n8636), .ZN(n8641)
         );
  NOR3_X1 U9974 ( .A1(n8639), .A2(n8740), .A3(n8638), .ZN(n8640) );
  AOI211_X1 U9975 ( .C1(n8738), .C2(n9421), .A(n8641), .B(n8640), .ZN(n8642)
         );
  OAI211_X1 U9976 ( .C1(n8645), .C2(n8644), .A(n8643), .B(n8642), .ZN(P1_U3218) );
  XOR2_X1 U9977 ( .A(n8646), .B(n8647), .Z(n8652) );
  AOI22_X1 U9978 ( .A1(n9114), .A2(n8734), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8649) );
  NAND2_X1 U9979 ( .A1(n8723), .A2(n9287), .ZN(n8648) );
  OAI211_X1 U9980 ( .C1(n9284), .C2(n8732), .A(n8649), .B(n8648), .ZN(n8650)
         );
  AOI21_X1 U9981 ( .B1(n9454), .B2(n8738), .A(n8650), .ZN(n8651) );
  OAI21_X1 U9982 ( .B1(n8652), .B2(n8740), .A(n8651), .ZN(P1_U3221) );
  AOI21_X1 U9983 ( .B1(n4343), .B2(n8653), .A(n8715), .ZN(n8658) );
  NAND2_X1 U9984 ( .A1(n9125), .A2(n8734), .ZN(n8655) );
  AOI22_X1 U9985 ( .A1(n9120), .A2(n8708), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8654) );
  OAI211_X1 U9986 ( .C1(n8736), .C2(n9226), .A(n8655), .B(n8654), .ZN(n8656)
         );
  AOI21_X1 U9987 ( .B1(n9434), .B2(n8738), .A(n8656), .ZN(n8657) );
  OAI21_X1 U9988 ( .B1(n8658), .B2(n8740), .A(n8657), .ZN(P1_U3223) );
  OAI21_X1 U9989 ( .B1(n8661), .B2(n8660), .A(n8659), .ZN(n8662) );
  NAND2_X1 U9990 ( .A1(n8662), .A2(n8717), .ZN(n8667) );
  INV_X1 U9991 ( .A(n9367), .ZN(n8665) );
  AOI22_X1 U9992 ( .A1(n8708), .A2(n9107), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n8663) );
  OAI21_X1 U9993 ( .B1(n9376), .B2(n8720), .A(n8663), .ZN(n8664) );
  AOI21_X1 U9994 ( .B1(n8665), .B2(n8723), .A(n8664), .ZN(n8666) );
  OAI211_X1 U9995 ( .C1(n4502), .C2(n8726), .A(n8667), .B(n8666), .ZN(P1_U3224) );
  OAI21_X1 U9996 ( .B1(n8670), .B2(n8669), .A(n8668), .ZN(n8671) );
  NAND2_X1 U9997 ( .A1(n8671), .A2(n8717), .ZN(n8676) );
  OAI22_X1 U9998 ( .A1(n8732), .A2(n9359), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8672), .ZN(n8674) );
  NOR2_X1 U9999 ( .A1(n8736), .A2(n9352), .ZN(n8673) );
  AOI211_X1 U10000 ( .C1(n8734), .C2(n9322), .A(n8674), .B(n8673), .ZN(n8675)
         );
  OAI211_X1 U10001 ( .C1(n9351), .C2(n8726), .A(n8676), .B(n8675), .ZN(
        P1_U3226) );
  AND3_X1 U10002 ( .A1(n8679), .A2(n8678), .A3(n8677), .ZN(n8680) );
  OAI21_X1 U10003 ( .B1(n8681), .B2(n8680), .A(n8717), .ZN(n8685) );
  AOI22_X1 U10004 ( .A1(n9116), .A2(n8708), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8682) );
  OAI21_X1 U10005 ( .B1(n9238), .B2(n8720), .A(n8682), .ZN(n8683) );
  AOI21_X1 U10006 ( .B1(n9240), .B2(n8723), .A(n8683), .ZN(n8684) );
  OAI211_X1 U10007 ( .C1(n9243), .C2(n8726), .A(n8685), .B(n8684), .ZN(
        P1_U3227) );
  NAND2_X1 U10008 ( .A1(n8688), .A2(n8687), .ZN(n8689) );
  XNOR2_X1 U10009 ( .A(n8686), .B(n8689), .ZN(n8695) );
  OAI22_X1 U10010 ( .A1(n9306), .A2(n8720), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8690), .ZN(n8691) );
  AOI21_X1 U10011 ( .B1(n8708), .B2(n9333), .A(n8691), .ZN(n8692) );
  OAI21_X1 U10012 ( .B1(n8736), .B2(n9296), .A(n8692), .ZN(n8693) );
  AOI21_X1 U10013 ( .B1(n9457), .B2(n8738), .A(n8693), .ZN(n8694) );
  OAI21_X1 U10014 ( .B1(n8695), .B2(n8740), .A(n8694), .ZN(P1_U3231) );
  NAND2_X1 U10015 ( .A1(n8696), .A2(n4362), .ZN(n8698) );
  XNOR2_X1 U10016 ( .A(n8698), .B(n8697), .ZN(n8703) );
  AOI22_X1 U10017 ( .A1(n9116), .A2(n8734), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8700) );
  NAND2_X1 U10018 ( .A1(n9015), .A2(n8708), .ZN(n8699) );
  OAI211_X1 U10019 ( .C1(n8736), .C2(n9268), .A(n8700), .B(n8699), .ZN(n8701)
         );
  AOI21_X1 U10020 ( .B1(n9449), .B2(n8738), .A(n8701), .ZN(n8702) );
  OAI21_X1 U10021 ( .B1(n8703), .B2(n8740), .A(n8702), .ZN(P1_U3233) );
  NAND2_X1 U10022 ( .A1(n4316), .A2(n8704), .ZN(n8705) );
  XOR2_X1 U10023 ( .A(n8706), .B(n8705), .Z(n8712) );
  NAND2_X1 U10024 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9909) );
  OAI21_X1 U10025 ( .B1(n8720), .B2(n9305), .A(n9909), .ZN(n8707) );
  AOI21_X1 U10026 ( .B1(n8708), .B2(n9332), .A(n8707), .ZN(n8709) );
  OAI21_X1 U10027 ( .B1(n8736), .B2(n9340), .A(n8709), .ZN(n8710) );
  AOI21_X1 U10028 ( .B1(n9468), .B2(n8738), .A(n8710), .ZN(n8711) );
  OAI21_X1 U10029 ( .B1(n8712), .B2(n8740), .A(n8711), .ZN(P1_U3236) );
  OAI21_X1 U10030 ( .B1(n8715), .B2(n8714), .A(n8713), .ZN(n8716) );
  NAND3_X1 U10031 ( .A1(n8718), .A2(n8717), .A3(n8716), .ZN(n8725) );
  OAI22_X1 U10032 ( .A1(n9238), .A2(n8732), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8719), .ZN(n8722) );
  NOR2_X1 U10033 ( .A1(n9210), .A2(n8720), .ZN(n8721) );
  AOI211_X1 U10034 ( .C1(n9213), .C2(n8723), .A(n8722), .B(n8721), .ZN(n8724)
         );
  OAI211_X1 U10035 ( .C1(n9216), .C2(n8726), .A(n8725), .B(n8724), .ZN(
        P1_U3238) );
  NAND2_X1 U10036 ( .A1(n8728), .A2(n8727), .ZN(n8729) );
  XOR2_X1 U10037 ( .A(n8730), .B(n8729), .Z(n8741) );
  OAI21_X1 U10038 ( .B1(n8732), .B2(n9105), .A(n8731), .ZN(n8733) );
  AOI21_X1 U10039 ( .B1(n8734), .B2(n9385), .A(n8733), .ZN(n8735) );
  OAI21_X1 U10040 ( .B1(n8736), .B2(n9390), .A(n8735), .ZN(n8737) );
  AOI21_X1 U10041 ( .B1(n9393), .B2(n8738), .A(n8737), .ZN(n8739) );
  OAI21_X1 U10042 ( .B1(n8741), .B2(n8740), .A(n8739), .ZN(P1_U3239) );
  OR2_X1 U10043 ( .A1(n9439), .A2(n9250), .ZN(n8863) );
  NAND2_X1 U10044 ( .A1(n8863), .A2(n9145), .ZN(n8987) );
  NAND2_X1 U10045 ( .A1(n9439), .A2(n9250), .ZN(n8862) );
  NAND2_X1 U10046 ( .A1(n8987), .A2(n8862), .ZN(n8742) );
  AND2_X1 U10047 ( .A1(n8946), .A2(n8742), .ZN(n8746) );
  NAND2_X1 U10048 ( .A1(n9434), .A2(n9238), .ZN(n8861) );
  NAND2_X1 U10049 ( .A1(n8861), .A2(n8862), .ZN(n9146) );
  NAND2_X1 U10050 ( .A1(n9444), .A2(n9265), .ZN(n8988) );
  INV_X1 U10051 ( .A(n8988), .ZN(n8743) );
  AND2_X1 U10052 ( .A1(n8863), .A2(n8743), .ZN(n8744) );
  NOR2_X1 U10053 ( .A1(n9146), .A2(n8744), .ZN(n8745) );
  INV_X1 U10054 ( .A(n8850), .ZN(n8800) );
  MUX2_X1 U10055 ( .A(n8746), .B(n8745), .S(n8800), .Z(n8809) );
  NAND2_X1 U10056 ( .A1(n7126), .A2(n8915), .ZN(n8747) );
  AND2_X1 U10057 ( .A1(n8974), .A2(n8967), .ZN(n8908) );
  NAND2_X1 U10058 ( .A1(n8747), .A2(n8908), .ZN(n8748) );
  NAND2_X1 U10059 ( .A1(n8748), .A2(n8918), .ZN(n8751) );
  INV_X1 U10060 ( .A(n8918), .ZN(n8749) );
  OAI21_X1 U10061 ( .B1(n8964), .B2(n8749), .A(n8974), .ZN(n8750) );
  MUX2_X1 U10062 ( .A(n8751), .B(n8750), .S(n8850), .Z(n8761) );
  NAND2_X1 U10063 ( .A1(n8920), .A2(n8919), .ZN(n8752) );
  OAI211_X1 U10064 ( .C1(n8761), .C2(n8752), .A(n8769), .B(n8898), .ZN(n8755)
         );
  NAND2_X1 U10065 ( .A1(n8776), .A2(n8753), .ZN(n8754) );
  MUX2_X1 U10066 ( .A(n8755), .B(n8754), .S(n8850), .Z(n8757) );
  XNOR2_X1 U10067 ( .A(n9809), .B(n8756), .ZN(n9793) );
  NOR2_X1 U10068 ( .A1(n8757), .A2(n9793), .ZN(n8766) );
  INV_X1 U10069 ( .A(n8758), .ZN(n8760) );
  OAI211_X1 U10070 ( .C1(n8761), .C2(n8760), .A(n8759), .B(n8919), .ZN(n8763)
         );
  NAND3_X1 U10071 ( .A1(n8763), .A2(n8897), .A3(n8762), .ZN(n8764) );
  MUX2_X1 U10072 ( .A(n8897), .B(n8764), .S(n8850), .Z(n8765) );
  NAND2_X1 U10073 ( .A1(n8766), .A2(n8765), .ZN(n8779) );
  AND2_X1 U10074 ( .A1(n8772), .A2(n8767), .ZN(n8925) );
  NAND2_X1 U10075 ( .A1(n8776), .A2(n8768), .ZN(n8922) );
  NAND2_X1 U10076 ( .A1(n8922), .A2(n8769), .ZN(n8770) );
  NAND3_X1 U10077 ( .A1(n8779), .A2(n8925), .A3(n8770), .ZN(n8775) );
  OR2_X1 U10078 ( .A1(n9779), .A2(n8771), .ZN(n8899) );
  NAND2_X1 U10079 ( .A1(n9133), .A2(n8899), .ZN(n8773) );
  NAND2_X1 U10080 ( .A1(n8773), .A2(n8772), .ZN(n8774) );
  NAND2_X1 U10081 ( .A1(n8775), .A2(n8774), .ZN(n8782) );
  INV_X1 U10082 ( .A(n8776), .ZN(n8777) );
  OR2_X1 U10083 ( .A1(n8778), .A2(n8777), .ZN(n8900) );
  NAND3_X1 U10084 ( .A1(n8779), .A2(n8900), .A3(n8899), .ZN(n8780) );
  INV_X1 U10085 ( .A(n9133), .ZN(n8902) );
  AOI21_X1 U10086 ( .B1(n8780), .B2(n8925), .A(n8902), .ZN(n8781) );
  MUX2_X1 U10087 ( .A(n8782), .B(n8781), .S(n8850), .Z(n8784) );
  INV_X1 U10088 ( .A(n9107), .ZN(n9375) );
  OR2_X1 U10089 ( .A1(n9393), .A2(n9375), .ZN(n8904) );
  NAND2_X1 U10090 ( .A1(n9393), .A2(n9375), .ZN(n8923) );
  NAND2_X1 U10091 ( .A1(n8904), .A2(n8923), .ZN(n9381) );
  NAND2_X1 U10092 ( .A1(n9481), .A2(n9359), .ZN(n9137) );
  NAND2_X1 U10093 ( .A1(n9136), .A2(n9137), .ZN(n9364) );
  INV_X1 U10094 ( .A(n9364), .ZN(n9372) );
  MUX2_X1 U10095 ( .A(n8904), .B(n8923), .S(n8800), .Z(n8783) );
  OAI211_X1 U10096 ( .C1(n8784), .C2(n9381), .A(n9372), .B(n8783), .ZN(n8786)
         );
  XNOR2_X1 U10097 ( .A(n9351), .B(n9376), .ZN(n9347) );
  MUX2_X1 U10098 ( .A(n9136), .B(n9137), .S(n8850), .Z(n8785) );
  NAND3_X1 U10099 ( .A1(n8786), .A2(n9347), .A3(n8785), .ZN(n8790) );
  NAND2_X1 U10100 ( .A1(n9468), .A2(n9360), .ZN(n9139) );
  AND2_X1 U10101 ( .A1(n9476), .A2(n9376), .ZN(n9138) );
  INV_X1 U10102 ( .A(n9138), .ZN(n8787) );
  AND2_X1 U10103 ( .A1(n9139), .A2(n8787), .ZN(n8896) );
  OR2_X1 U10104 ( .A1(n9468), .A2(n9360), .ZN(n8866) );
  OR2_X1 U10105 ( .A1(n9476), .A2(n9376), .ZN(n9328) );
  NAND2_X1 U10106 ( .A1(n8866), .A2(n9328), .ZN(n9140) );
  INV_X1 U10107 ( .A(n9140), .ZN(n8788) );
  MUX2_X1 U10108 ( .A(n8896), .B(n8788), .S(n8850), .Z(n8789) );
  NAND2_X1 U10109 ( .A1(n8790), .A2(n8789), .ZN(n8794) );
  NAND2_X1 U10110 ( .A1(n9462), .A2(n9305), .ZN(n8933) );
  NAND3_X1 U10111 ( .A1(n8794), .A2(n8933), .A3(n9139), .ZN(n8793) );
  OR2_X1 U10112 ( .A1(n9462), .A2(n9305), .ZN(n8934) );
  NAND4_X1 U10113 ( .A1(n8865), .A2(n9303), .A3(n8934), .A4(n8850), .ZN(n8791)
         );
  NOR2_X1 U10114 ( .A1(n9143), .A2(n8791), .ZN(n8792) );
  NAND2_X1 U10115 ( .A1(n8793), .A2(n8792), .ZN(n8807) );
  NAND3_X1 U10116 ( .A1(n8794), .A2(n8934), .A3(n8866), .ZN(n8796) );
  NAND2_X1 U10117 ( .A1(n9449), .A2(n9285), .ZN(n8864) );
  NAND2_X1 U10118 ( .A1(n9454), .A2(n9306), .ZN(n9261) );
  AND2_X1 U10119 ( .A1(n8864), .A2(n9261), .ZN(n9144) );
  NAND2_X1 U10120 ( .A1(n9457), .A2(n9284), .ZN(n9142) );
  AND4_X1 U10121 ( .A1(n9144), .A2(n8800), .A3(n9142), .A4(n8933), .ZN(n8795)
         );
  NAND2_X1 U10122 ( .A1(n8796), .A2(n8795), .ZN(n8806) );
  INV_X1 U10123 ( .A(n8987), .ZN(n8943) );
  INV_X1 U10124 ( .A(n8862), .ZN(n9220) );
  OR3_X1 U10125 ( .A1(n9143), .A2(n9144), .A3(n8800), .ZN(n8803) );
  INV_X1 U10126 ( .A(n9142), .ZN(n8797) );
  NAND2_X1 U10127 ( .A1(n8865), .A2(n8797), .ZN(n8929) );
  NOR2_X1 U10128 ( .A1(n8929), .A2(n8800), .ZN(n8799) );
  NAND2_X1 U10129 ( .A1(n9143), .A2(n8850), .ZN(n8798) );
  OAI21_X1 U10130 ( .B1(n9143), .B2(n8799), .A(n8798), .ZN(n8802) );
  NAND2_X1 U10131 ( .A1(n8865), .A2(n9303), .ZN(n8937) );
  NAND3_X1 U10132 ( .A1(n9144), .A2(n8800), .A3(n8937), .ZN(n8801) );
  NAND4_X1 U10133 ( .A1(n8803), .A2(n8802), .A3(n8988), .A4(n8801), .ZN(n8804)
         );
  NOR2_X1 U10134 ( .A1(n9220), .A2(n8804), .ZN(n8805) );
  NAND4_X1 U10135 ( .A1(n8807), .A2(n8806), .A3(n8943), .A4(n8805), .ZN(n8808)
         );
  NAND2_X1 U10136 ( .A1(n8809), .A2(n8808), .ZN(n8817) );
  NAND2_X1 U10137 ( .A1(n8817), .A2(n8946), .ZN(n8810) );
  AOI21_X1 U10138 ( .B1(n8810), .B2(n9216), .A(n9125), .ZN(n8813) );
  NAND2_X1 U10139 ( .A1(n8817), .A2(n8861), .ZN(n8811) );
  AOI21_X1 U10140 ( .B1(n8811), .B2(n9224), .A(n9429), .ZN(n8812) );
  MUX2_X1 U10141 ( .A(n8813), .B(n8812), .S(n8850), .Z(n8823) );
  INV_X1 U10142 ( .A(n8946), .ZN(n9206) );
  NAND2_X1 U10143 ( .A1(n9422), .A2(n9210), .ZN(n8949) );
  OAI21_X1 U10144 ( .B1(n9216), .B2(n9206), .A(n8949), .ZN(n8816) );
  NAND2_X1 U10145 ( .A1(n8861), .A2(n9125), .ZN(n8814) );
  NAND2_X1 U10146 ( .A1(n8945), .A2(n8814), .ZN(n8815) );
  MUX2_X1 U10147 ( .A(n8816), .B(n8815), .S(n8850), .Z(n8820) );
  INV_X1 U10148 ( .A(n8817), .ZN(n8818) );
  NAND2_X1 U10149 ( .A1(n8818), .A2(n9128), .ZN(n8819) );
  AND2_X1 U10150 ( .A1(n8820), .A2(n8819), .ZN(n8822) );
  NAND2_X1 U10151 ( .A1(n9421), .A2(n9192), .ZN(n8950) );
  MUX2_X1 U10152 ( .A(n8945), .B(n8949), .S(n8850), .Z(n8821) );
  OAI211_X1 U10153 ( .C1(n8823), .C2(n8822), .A(n9171), .B(n8821), .ZN(n8825)
         );
  MUX2_X1 U10154 ( .A(n8950), .B(n9150), .S(n8850), .Z(n8824) );
  NAND2_X1 U10155 ( .A1(n8825), .A2(n8824), .ZN(n8853) );
  NAND2_X1 U10156 ( .A1(n8826), .A2(n8840), .ZN(n8829) );
  OR2_X1 U10157 ( .A1(n5057), .A2(n8827), .ZN(n8828) );
  INV_X1 U10158 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8833) );
  NAND2_X1 U10159 ( .A1(n8830), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8832) );
  NAND2_X1 U10160 ( .A1(n5477), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8831) );
  OAI211_X1 U10161 ( .C1(n5685), .C2(n8833), .A(n8832), .B(n8831), .ZN(n9155)
         );
  NAND2_X1 U10162 ( .A1(n9096), .A2(n9155), .ZN(n8834) );
  NAND2_X1 U10163 ( .A1(n9099), .A2(n8834), .ZN(n8849) );
  INV_X1 U10164 ( .A(n8849), .ZN(n8955) );
  NOR2_X1 U10165 ( .A1(n8853), .A2(n8955), .ZN(n8839) );
  INV_X1 U10166 ( .A(n9155), .ZN(n8859) );
  NAND2_X1 U10167 ( .A1(n8839), .A2(n8851), .ZN(n8845) );
  INV_X1 U10168 ( .A(n9012), .ZN(n9177) );
  OAI21_X1 U10169 ( .B1(n8845), .B2(n9177), .A(n8851), .ZN(n8847) );
  NAND2_X1 U10170 ( .A1(n8841), .A2(n8840), .ZN(n8844) );
  OR2_X1 U10171 ( .A1(n5057), .A2(n8842), .ZN(n8843) );
  INV_X1 U10172 ( .A(n9412), .ZN(n9166) );
  NOR2_X1 U10173 ( .A1(n9743), .A2(n9096), .ZN(n8998) );
  OAI22_X1 U10174 ( .A1(n8845), .A2(n9166), .B1(n8998), .B2(n8849), .ZN(n8846)
         );
  NOR2_X1 U10175 ( .A1(n9412), .A2(n9012), .ZN(n8854) );
  NAND2_X1 U10176 ( .A1(n9012), .A2(n8850), .ZN(n8848) );
  OAI211_X1 U10177 ( .C1(n9166), .C2(n8850), .A(n8849), .B(n8848), .ZN(n8852)
         );
  AOI211_X1 U10178 ( .C1(n8854), .C2(n8853), .A(n8852), .B(n8959), .ZN(n8855)
         );
  AND2_X1 U10179 ( .A1(n9743), .A2(n9096), .ZN(n8858) );
  INV_X1 U10180 ( .A(n8858), .ZN(n8957) );
  NAND2_X1 U10181 ( .A1(n9099), .A2(n8859), .ZN(n8860) );
  NAND2_X1 U10182 ( .A1(n8957), .A2(n8860), .ZN(n8962) );
  XNOR2_X1 U10183 ( .A(n9216), .B(n9125), .ZN(n9207) );
  NAND2_X1 U10184 ( .A1(n8863), .A2(n8862), .ZN(n9236) );
  NAND2_X1 U10185 ( .A1(n9145), .A2(n8988), .ZN(n9247) );
  INV_X1 U10186 ( .A(n9143), .ZN(n8940) );
  NAND2_X1 U10187 ( .A1(n8940), .A2(n8864), .ZN(n9262) );
  INV_X1 U10188 ( .A(n9335), .ZN(n8883) );
  INV_X1 U10189 ( .A(n9347), .ZN(n9356) );
  INV_X1 U10190 ( .A(n9381), .ZN(n9379) );
  INV_X1 U10191 ( .A(n8867), .ZN(n8869) );
  NAND4_X1 U10192 ( .A1(n8871), .A2(n8870), .A3(n8869), .A4(n8868), .ZN(n8873)
         );
  NOR4_X1 U10193 ( .A1(n8873), .A2(n7105), .A3(n8872), .A4(n6501), .ZN(n8877)
         );
  NAND4_X1 U10194 ( .A1(n8877), .A2(n8876), .A3(n8875), .A4(n8874), .ZN(n8880)
         );
  NOR4_X1 U10195 ( .A1(n8880), .A2(n8879), .A3(n9793), .A4(n8878), .ZN(n8881)
         );
  NAND4_X1 U10196 ( .A1(n9379), .A2(n7557), .A3(n8881), .A4(n9766), .ZN(n8882)
         );
  NOR4_X1 U10197 ( .A1(n8883), .A2(n9356), .A3(n9364), .A4(n8882), .ZN(n8884)
         );
  NAND4_X1 U10198 ( .A1(n9280), .A2(n9300), .A3(n9320), .A4(n8884), .ZN(n8885)
         );
  OR4_X1 U10199 ( .A1(n9236), .A2(n9247), .A3(n9262), .A4(n8885), .ZN(n8886)
         );
  NOR4_X1 U10200 ( .A1(n9191), .A2(n9207), .A3(n9222), .A4(n8886), .ZN(n8887)
         );
  NAND4_X1 U10201 ( .A1(n8993), .A2(n9171), .A3(n8887), .A4(n9152), .ZN(n8888)
         );
  NOR3_X1 U10202 ( .A1(n8998), .A2(n8962), .A3(n8888), .ZN(n8889) );
  NOR2_X1 U10203 ( .A1(n8889), .A2(n5663), .ZN(n8894) );
  NAND3_X1 U10204 ( .A1(n8957), .A2(n5663), .A3(n4515), .ZN(n8891) );
  INV_X1 U10205 ( .A(n8894), .ZN(n8961) );
  OR2_X1 U10206 ( .A1(n9412), .A2(n9177), .ZN(n8895) );
  NAND2_X1 U10207 ( .A1(n8895), .A2(n9150), .ZN(n8992) );
  INV_X1 U10208 ( .A(n8896), .ZN(n8927) );
  AND2_X1 U10209 ( .A1(n8898), .A2(n8897), .ZN(n8901) );
  OAI211_X1 U10210 ( .C1(n8901), .C2(n8922), .A(n8900), .B(n8899), .ZN(n8903)
         );
  AOI21_X1 U10211 ( .B1(n8925), .B2(n8903), .A(n8902), .ZN(n8905) );
  INV_X1 U10212 ( .A(n8923), .ZN(n9135) );
  OAI211_X1 U10213 ( .C1(n8905), .C2(n9135), .A(n9136), .B(n8904), .ZN(n8906)
         );
  NAND2_X1 U10214 ( .A1(n8906), .A2(n9137), .ZN(n8907) );
  NOR2_X1 U10215 ( .A1(n8927), .A2(n8907), .ZN(n8978) );
  INV_X1 U10216 ( .A(n8908), .ZN(n8909) );
  NOR2_X1 U10217 ( .A1(n8978), .A2(n8909), .ZN(n8932) );
  NOR2_X1 U10218 ( .A1(n8911), .A2(n4619), .ZN(n8917) );
  AND2_X1 U10219 ( .A1(n8913), .A2(n8912), .ZN(n8972) );
  INV_X1 U10220 ( .A(n8972), .ZN(n8916) );
  OAI211_X1 U10221 ( .C1(n8917), .C2(n8916), .A(n8915), .B(n8914), .ZN(n8931)
         );
  NAND3_X1 U10222 ( .A1(n8920), .A2(n8919), .A3(n8918), .ZN(n8921) );
  NOR2_X1 U10223 ( .A1(n8922), .A2(n8921), .ZN(n8924) );
  NAND4_X1 U10224 ( .A1(n9137), .A2(n8925), .A3(n8924), .A4(n8923), .ZN(n8926)
         );
  NOR2_X1 U10225 ( .A1(n8927), .A2(n8926), .ZN(n8963) );
  NAND4_X1 U10226 ( .A1(n8932), .A2(n8972), .A3(n8973), .A4(n7043), .ZN(n8928)
         );
  OAI21_X1 U10227 ( .B1(n8978), .B2(n8963), .A(n8928), .ZN(n8930) );
  NAND2_X1 U10228 ( .A1(n9144), .A2(n8929), .ZN(n8939) );
  INV_X1 U10229 ( .A(n8933), .ZN(n9141) );
  OR2_X1 U10230 ( .A1(n8939), .A2(n9141), .ZN(n8985) );
  AOI211_X1 U10231 ( .C1(n8932), .C2(n8931), .A(n8930), .B(n8985), .ZN(n8942)
         );
  NAND3_X1 U10232 ( .A1(n8933), .A2(n9139), .A3(n9140), .ZN(n8935) );
  NAND2_X1 U10233 ( .A1(n8935), .A2(n8934), .ZN(n8936) );
  NOR2_X1 U10234 ( .A1(n8937), .A2(n8936), .ZN(n8938) );
  OR2_X1 U10235 ( .A1(n8939), .A2(n8938), .ZN(n8941) );
  NAND2_X1 U10236 ( .A1(n8941), .A2(n8940), .ZN(n8983) );
  OAI21_X1 U10237 ( .B1(n8942), .B2(n8983), .A(n8988), .ZN(n8944) );
  AOI21_X1 U10238 ( .B1(n8944), .B2(n8943), .A(n9146), .ZN(n8948) );
  INV_X1 U10239 ( .A(n8945), .ZN(n9149) );
  OR2_X1 U10240 ( .A1(n9429), .A2(n9224), .ZN(n8947) );
  NAND2_X1 U10241 ( .A1(n8947), .A2(n8946), .ZN(n9148) );
  NOR4_X1 U10242 ( .A1(n8992), .A2(n8948), .A3(n9149), .A4(n9148), .ZN(n8956)
         );
  NAND2_X1 U10243 ( .A1(n9429), .A2(n9224), .ZN(n9147) );
  OAI211_X1 U10244 ( .C1(n9149), .C2(n9147), .A(n8950), .B(n8949), .ZN(n8951)
         );
  INV_X1 U10245 ( .A(n8951), .ZN(n8952) );
  OR2_X1 U10246 ( .A1(n8992), .A2(n8952), .ZN(n8954) );
  NAND2_X1 U10247 ( .A1(n9412), .A2(n9177), .ZN(n8953) );
  NAND2_X1 U10248 ( .A1(n8954), .A2(n8953), .ZN(n8995) );
  NOR3_X1 U10249 ( .A1(n8956), .A2(n8955), .A3(n8995), .ZN(n8958) );
  OAI211_X1 U10250 ( .C1(n8959), .C2(n8958), .A(n5663), .B(n8957), .ZN(n8960)
         );
  INV_X1 U10251 ( .A(n8962), .ZN(n8997) );
  INV_X1 U10252 ( .A(n8963), .ZN(n8981) );
  INV_X1 U10253 ( .A(n8964), .ZN(n8977) );
  INV_X1 U10254 ( .A(n8965), .ZN(n8968) );
  NAND2_X1 U10255 ( .A1(n9403), .A2(n9026), .ZN(n8966) );
  AND4_X1 U10256 ( .A1(n8968), .A2(n8967), .A3(n5663), .A4(n8966), .ZN(n8971)
         );
  NAND2_X1 U10257 ( .A1(n8969), .A2(n6500), .ZN(n8970) );
  NAND4_X1 U10258 ( .A1(n8973), .A2(n8972), .A3(n8971), .A4(n8970), .ZN(n8976)
         );
  INV_X1 U10259 ( .A(n8974), .ZN(n8975) );
  AOI21_X1 U10260 ( .B1(n8977), .B2(n8976), .A(n8975), .ZN(n8980) );
  INV_X1 U10261 ( .A(n8978), .ZN(n8979) );
  OAI21_X1 U10262 ( .B1(n8981), .B2(n8980), .A(n8979), .ZN(n8982) );
  INV_X1 U10263 ( .A(n8982), .ZN(n8986) );
  INV_X1 U10264 ( .A(n8983), .ZN(n8984) );
  OAI21_X1 U10265 ( .B1(n8986), .B2(n8985), .A(n8984), .ZN(n8989) );
  AOI21_X1 U10266 ( .B1(n8989), .B2(n8988), .A(n8987), .ZN(n8990) );
  OAI211_X1 U10267 ( .C1(n8990), .C2(n9146), .A(n9128), .B(n4626), .ZN(n8991)
         );
  NOR2_X1 U10268 ( .A1(n8992), .A2(n8991), .ZN(n8994) );
  OAI21_X1 U10269 ( .B1(n8995), .B2(n8994), .A(n8993), .ZN(n8996) );
  NAND2_X1 U10270 ( .A1(n8997), .A2(n8996), .ZN(n9000) );
  INV_X1 U10271 ( .A(n8998), .ZN(n8999) );
  NAND2_X1 U10272 ( .A1(n9000), .A2(n8999), .ZN(n9004) );
  NOR3_X1 U10273 ( .A1(n9004), .A2(n9002), .A3(n9001), .ZN(n9003) );
  AOI211_X1 U10274 ( .C1(n9005), .C2(n9004), .A(n9010), .B(n9003), .ZN(n9006)
         );
  NAND3_X1 U10275 ( .A1(n9008), .A2(n9505), .A3(n9007), .ZN(n9009) );
  OAI211_X1 U10276 ( .C1(n5662), .C2(n9010), .A(n9009), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9011) );
  MUX2_X1 U10277 ( .A(n9155), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9027), .Z(
        P1_U3585) );
  MUX2_X1 U10278 ( .A(n9012), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9027), .Z(
        P1_U3584) );
  MUX2_X1 U10279 ( .A(n9157), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9027), .Z(
        P1_U3583) );
  MUX2_X1 U10280 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9013), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10281 ( .A(n9125), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9027), .Z(
        P1_U3581) );
  MUX2_X1 U10282 ( .A(n9014), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9027), .Z(
        P1_U3580) );
  MUX2_X1 U10283 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9120), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10284 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9116), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10285 ( .A(n9114), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9027), .Z(
        P1_U3577) );
  MUX2_X1 U10286 ( .A(n9015), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9027), .Z(
        P1_U3576) );
  MUX2_X1 U10287 ( .A(n9323), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9027), .Z(
        P1_U3575) );
  MUX2_X1 U10288 ( .A(n9333), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9027), .Z(
        P1_U3574) );
  MUX2_X1 U10289 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9322), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10290 ( .A(n9332), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9027), .Z(
        P1_U3572) );
  MUX2_X1 U10291 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9385), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10292 ( .A(n9107), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9027), .Z(
        P1_U3570) );
  MUX2_X1 U10293 ( .A(n9770), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9027), .Z(
        P1_U3569) );
  MUX2_X1 U10294 ( .A(n9016), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9027), .Z(
        P1_U3568) );
  MUX2_X1 U10295 ( .A(n9773), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9027), .Z(
        P1_U3567) );
  MUX2_X1 U10296 ( .A(n9017), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9027), .Z(
        P1_U3566) );
  MUX2_X1 U10297 ( .A(n9018), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9027), .Z(
        P1_U3565) );
  MUX2_X1 U10298 ( .A(n9019), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9027), .Z(
        P1_U3564) );
  MUX2_X1 U10299 ( .A(n9020), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9027), .Z(
        P1_U3563) );
  MUX2_X1 U10300 ( .A(n9021), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9027), .Z(
        P1_U3562) );
  MUX2_X1 U10301 ( .A(n9022), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9027), .Z(
        P1_U3561) );
  MUX2_X1 U10302 ( .A(n9023), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9027), .Z(
        P1_U3560) );
  MUX2_X1 U10303 ( .A(n9024), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9027), .Z(
        P1_U3559) );
  MUX2_X1 U10304 ( .A(n9025), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9027), .Z(
        P1_U3558) );
  MUX2_X1 U10305 ( .A(n9026), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9027), .Z(
        P1_U3557) );
  MUX2_X1 U10306 ( .A(n6500), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9027), .Z(
        P1_U3556) );
  MUX2_X1 U10307 ( .A(n9028), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9027), .Z(
        P1_U3555) );
  OAI21_X1 U10308 ( .B1(n9031), .B2(n9030), .A(n9029), .ZN(n9032) );
  NAND2_X1 U10309 ( .A1(n9032), .A2(n9921), .ZN(n9042) );
  OAI21_X1 U10310 ( .B1(n9035), .B2(n9034), .A(n9033), .ZN(n9036) );
  NAND2_X1 U10311 ( .A1(n9036), .A2(n9920), .ZN(n9041) );
  INV_X1 U10312 ( .A(n9925), .ZN(n9906) );
  NOR2_X1 U10313 ( .A1(n9057), .A2(n9037), .ZN(n9038) );
  AOI211_X1 U10314 ( .C1(n9906), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n9039), .B(
        n9038), .ZN(n9040) );
  NAND3_X1 U10315 ( .A1(n9042), .A2(n9041), .A3(n9040), .ZN(P1_U3252) );
  NOR2_X1 U10316 ( .A1(n9043), .A2(n9049), .ZN(n9045) );
  NAND2_X1 U10317 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9068), .ZN(n9046) );
  OAI21_X1 U10318 ( .B1(n9068), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9046), .ZN(
        n9047) );
  AOI211_X1 U10319 ( .C1(n4375), .C2(n9047), .A(n9067), .B(n9885), .ZN(n9060)
         );
  NOR2_X1 U10320 ( .A1(n9049), .A2(n9048), .ZN(n9051) );
  NOR2_X1 U10321 ( .A1(n9051), .A2(n9050), .ZN(n9053) );
  XNOR2_X1 U10322 ( .A(n9068), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9052) );
  NOR2_X1 U10323 ( .A1(n9053), .A2(n9052), .ZN(n9061) );
  AOI211_X1 U10324 ( .C1(n9053), .C2(n9052), .A(n9061), .B(n9898), .ZN(n9059)
         );
  NAND2_X1 U10325 ( .A1(n9906), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9055) );
  NAND2_X1 U10326 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n9054) );
  OAI211_X1 U10327 ( .C1(n9057), .C2(n9056), .A(n9055), .B(n9054), .ZN(n9058)
         );
  OR3_X1 U10328 ( .A1(n9060), .A2(n9059), .A3(n9058), .ZN(P1_U3257) );
  INV_X1 U10329 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9076) );
  XNOR2_X1 U10330 ( .A(n9083), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9063) );
  AOI21_X1 U10331 ( .B1(n9068), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9061), .ZN(
        n9062) );
  NOR2_X1 U10332 ( .A1(n9062), .A2(n9063), .ZN(n9082) );
  AOI21_X1 U10333 ( .B1(n9063), .B2(n9062), .A(n9082), .ZN(n9064) );
  NAND2_X1 U10334 ( .A1(n9920), .A2(n9064), .ZN(n9066) );
  NAND2_X1 U10335 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n9065) );
  NAND2_X1 U10336 ( .A1(n9066), .A2(n9065), .ZN(n9074) );
  AOI21_X1 U10337 ( .B1(n9068), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9067), .ZN(
        n9072) );
  NOR2_X1 U10338 ( .A1(n9083), .A2(n9069), .ZN(n9070) );
  AOI21_X1 U10339 ( .B1(n9069), .B2(n9083), .A(n9070), .ZN(n9071) );
  NOR2_X1 U10340 ( .A1(n9072), .A2(n9071), .ZN(n9077) );
  AOI211_X1 U10341 ( .C1(n9072), .C2(n9071), .A(n9077), .B(n9885), .ZN(n9073)
         );
  AOI211_X1 U10342 ( .C1(n9912), .C2(n9083), .A(n9074), .B(n9073), .ZN(n9075)
         );
  OAI21_X1 U10343 ( .B1(n9925), .B2(n9076), .A(n9075), .ZN(P1_U3258) );
  INV_X1 U10344 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9092) );
  NAND2_X1 U10345 ( .A1(n9911), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9078) );
  OAI21_X1 U10346 ( .B1(n9911), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9078), .ZN(
        n9914) );
  NOR2_X1 U10347 ( .A1(n9915), .A2(n9914), .ZN(n9913) );
  AOI21_X1 U10348 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9911), .A(n9913), .ZN(
        n9079) );
  XNOR2_X1 U10349 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9079), .ZN(n9088) );
  AOI22_X1 U10350 ( .A1(n9911), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9081), .B2(
        n9080), .ZN(n9918) );
  AOI21_X1 U10351 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9083), .A(n9082), .ZN(
        n9917) );
  NAND2_X1 U10352 ( .A1(n9918), .A2(n9917), .ZN(n9916) );
  OAI21_X1 U10353 ( .B1(n9911), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9916), .ZN(
        n9085) );
  XOR2_X1 U10354 ( .A(n9085), .B(n9084), .Z(n9086) );
  AOI22_X1 U10355 ( .A1(n9088), .A2(n9921), .B1(n9920), .B2(n9086), .ZN(n9090)
         );
  INV_X1 U10356 ( .A(n9086), .ZN(n9089) );
  OR2_X2 U10357 ( .A1(n9365), .A2(n9476), .ZN(n9349) );
  NAND2_X1 U10358 ( .A1(n9338), .A2(n9319), .ZN(n9312) );
  OR2_X2 U10359 ( .A1(n9312), .A2(n9457), .ZN(n9294) );
  NOR2_X2 U10360 ( .A1(n9239), .A2(n9434), .ZN(n9225) );
  AND2_X2 U10361 ( .A1(n9225), .A2(n9216), .ZN(n9211) );
  NAND2_X1 U10362 ( .A1(n9160), .A2(n9814), .ZN(n9093) );
  XNOR2_X1 U10363 ( .A(n9743), .B(n9093), .ZN(n9745) );
  NAND2_X1 U10364 ( .A1(n9745), .A2(n9787), .ZN(n9098) );
  AND2_X1 U10365 ( .A1(n9094), .A2(P1_B_REG_SCAN_IN), .ZN(n9095) );
  NOR2_X1 U10366 ( .A1(n9796), .A2(n9095), .ZN(n9156) );
  NAND2_X1 U10367 ( .A1(n9156), .A2(n9096), .ZN(n9813) );
  NOR2_X1 U10368 ( .A1(n9806), .A2(n9813), .ZN(n9100) );
  AOI21_X1 U10369 ( .B1(n9806), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9100), .ZN(
        n9097) );
  OAI211_X1 U10370 ( .C1(n9404), .C2(n9743), .A(n9098), .B(n9097), .ZN(
        P1_U3261) );
  XNOR2_X1 U10371 ( .A(n9160), .B(n9099), .ZN(n9817) );
  NAND2_X1 U10372 ( .A1(n9817), .A2(n9787), .ZN(n9102) );
  AOI21_X1 U10373 ( .B1(n9806), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9100), .ZN(
        n9101) );
  OAI211_X1 U10374 ( .C1(n9814), .C2(n9404), .A(n9102), .B(n9101), .ZN(
        P1_U3262) );
  NAND2_X1 U10375 ( .A1(n9486), .A2(n9770), .ZN(n9106) );
  NAND2_X1 U10376 ( .A1(n9380), .A2(n9108), .ZN(n9109) );
  NAND2_X1 U10377 ( .A1(n9109), .A2(n4873), .ZN(n9363) );
  NAND2_X1 U10378 ( .A1(n9363), .A2(n9364), .ZN(n9111) );
  NOR2_X1 U10379 ( .A1(n9299), .A2(n9284), .ZN(n9113) );
  INV_X1 U10380 ( .A(n9454), .ZN(n9290) );
  NAND2_X1 U10381 ( .A1(n9257), .A2(n9265), .ZN(n9118) );
  NAND2_X1 U10382 ( .A1(n9233), .A2(n9119), .ZN(n9122) );
  NAND2_X1 U10383 ( .A1(n9243), .A2(n9250), .ZN(n9121) );
  NAND2_X1 U10384 ( .A1(n9122), .A2(n9121), .ZN(n9219) );
  NAND2_X1 U10385 ( .A1(n9216), .A2(n9224), .ZN(n9124) );
  NAND2_X1 U10386 ( .A1(n9205), .A2(n9124), .ZN(n9127) );
  NAND2_X1 U10387 ( .A1(n9429), .A2(n9125), .ZN(n9126) );
  NAND2_X1 U10388 ( .A1(n9201), .A2(n9210), .ZN(n9129) );
  NAND2_X1 U10389 ( .A1(n9130), .A2(n9175), .ZN(n9173) );
  NAND2_X1 U10390 ( .A1(n9421), .A2(n9157), .ZN(n9131) );
  NAND2_X1 U10391 ( .A1(n9173), .A2(n9131), .ZN(n9132) );
  XNOR2_X1 U10392 ( .A(n9132), .B(n9152), .ZN(n9411) );
  INV_X1 U10393 ( .A(n9411), .ZN(n9169) );
  INV_X1 U10394 ( .A(n9171), .ZN(n9175) );
  INV_X1 U10395 ( .A(n9150), .ZN(n9151) );
  NOR2_X1 U10396 ( .A1(n9174), .A2(n9151), .ZN(n9154) );
  XNOR2_X1 U10397 ( .A(n9154), .B(n9153), .ZN(n9159) );
  AOI22_X1 U10398 ( .A1(n9157), .A2(n9772), .B1(n9156), .B2(n9155), .ZN(n9158)
         );
  OAI21_X1 U10399 ( .B1(n9159), .B2(n9802), .A(n9158), .ZN(n9415) );
  NOR2_X1 U10400 ( .A1(n9806), .A2(n9161), .ZN(n9355) );
  NAND2_X1 U10401 ( .A1(n9414), .A2(n9355), .ZN(n9165) );
  INV_X1 U10402 ( .A(n9162), .ZN(n9163) );
  AOI22_X1 U10403 ( .A1(n9163), .A2(n9316), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9806), .ZN(n9164) );
  OAI211_X1 U10404 ( .C1(n9166), .C2(n9404), .A(n9165), .B(n9164), .ZN(n9167)
         );
  AOI21_X1 U10405 ( .B1(n9415), .B2(n9792), .A(n9167), .ZN(n9168) );
  OAI21_X1 U10406 ( .B1(n9169), .B2(n9398), .A(n9168), .ZN(P1_U3355) );
  NAND2_X1 U10407 ( .A1(n9170), .A2(n9171), .ZN(n9172) );
  INV_X1 U10408 ( .A(n9418), .ZN(n9187) );
  OAI22_X1 U10409 ( .A1(n9210), .A2(n9798), .B1(n9177), .B2(n9796), .ZN(n9178)
         );
  INV_X1 U10410 ( .A(n9421), .ZN(n9184) );
  INV_X1 U10411 ( .A(n9179), .ZN(n9180) );
  AOI211_X1 U10412 ( .C1(n9421), .C2(n9195), .A(n9963), .B(n9180), .ZN(n9420)
         );
  NAND2_X1 U10413 ( .A1(n9420), .A2(n9355), .ZN(n9183) );
  AOI22_X1 U10414 ( .A1(n9181), .A2(n9316), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9806), .ZN(n9182) );
  OAI211_X1 U10415 ( .C1(n9184), .C2(n9404), .A(n9183), .B(n9182), .ZN(n9185)
         );
  AOI21_X1 U10416 ( .B1(n9419), .B2(n9792), .A(n9185), .ZN(n9186) );
  OAI21_X1 U10417 ( .B1(n9187), .B2(n9398), .A(n9186), .ZN(P1_U3263) );
  XNOR2_X1 U10418 ( .A(n9188), .B(n9191), .ZN(n9426) );
  AOI211_X1 U10419 ( .C1(n9191), .C2(n9190), .A(n9802), .B(n9189), .ZN(n9194)
         );
  OAI22_X1 U10420 ( .A1(n9192), .A2(n9796), .B1(n9224), .B2(n9798), .ZN(n9193)
         );
  NOR2_X1 U10421 ( .A1(n9194), .A2(n9193), .ZN(n9425) );
  INV_X1 U10422 ( .A(n9425), .ZN(n9203) );
  INV_X1 U10423 ( .A(n9211), .ZN(n9197) );
  INV_X1 U10424 ( .A(n9195), .ZN(n9196) );
  AOI21_X1 U10425 ( .B1(n9422), .B2(n9197), .A(n9196), .ZN(n9423) );
  NAND2_X1 U10426 ( .A1(n9423), .A2(n9787), .ZN(n9200) );
  AOI22_X1 U10427 ( .A1(n9198), .A2(n9316), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9806), .ZN(n9199) );
  OAI211_X1 U10428 ( .C1(n9201), .C2(n9404), .A(n9200), .B(n9199), .ZN(n9202)
         );
  AOI21_X1 U10429 ( .B1(n9203), .B2(n9792), .A(n9202), .ZN(n9204) );
  OAI21_X1 U10430 ( .B1(n9426), .B2(n9398), .A(n9204), .ZN(P1_U3264) );
  XNOR2_X1 U10431 ( .A(n9205), .B(n9207), .ZN(n9431) );
  XNOR2_X1 U10432 ( .A(n9208), .B(n9207), .ZN(n9209) );
  OAI222_X1 U10433 ( .A1(n9796), .A2(n9210), .B1(n9798), .B2(n9238), .C1(n9209), .C2(n9802), .ZN(n9427) );
  INV_X1 U10434 ( .A(n9225), .ZN(n9212) );
  AOI211_X1 U10435 ( .C1(n9429), .C2(n9212), .A(n9963), .B(n9211), .ZN(n9428)
         );
  NAND2_X1 U10436 ( .A1(n9428), .A2(n9355), .ZN(n9215) );
  AOI22_X1 U10437 ( .A1(n9213), .A2(n9316), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9806), .ZN(n9214) );
  OAI211_X1 U10438 ( .C1(n9216), .C2(n9404), .A(n9215), .B(n9214), .ZN(n9217)
         );
  AOI21_X1 U10439 ( .B1(n9427), .B2(n9792), .A(n9217), .ZN(n9218) );
  OAI21_X1 U10440 ( .B1(n9431), .B2(n9398), .A(n9218), .ZN(P1_U3265) );
  XOR2_X1 U10441 ( .A(n9222), .B(n9219), .Z(n9436) );
  NOR2_X1 U10442 ( .A1(n9234), .A2(n9220), .ZN(n9221) );
  XOR2_X1 U10443 ( .A(n9222), .B(n9221), .Z(n9223) );
  OAI222_X1 U10444 ( .A1(n9796), .A2(n9224), .B1(n9798), .B2(n9250), .C1(n9223), .C2(n9802), .ZN(n9432) );
  AOI211_X1 U10445 ( .C1(n9434), .C2(n9239), .A(n9963), .B(n9225), .ZN(n9433)
         );
  NAND2_X1 U10446 ( .A1(n9433), .A2(n9355), .ZN(n9229) );
  INV_X1 U10447 ( .A(n9226), .ZN(n9227) );
  AOI22_X1 U10448 ( .A1(n9227), .A2(n9316), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9806), .ZN(n9228) );
  OAI211_X1 U10449 ( .C1(n9230), .C2(n9404), .A(n9229), .B(n9228), .ZN(n9231)
         );
  AOI21_X1 U10450 ( .B1(n9432), .B2(n9792), .A(n9231), .ZN(n9232) );
  OAI21_X1 U10451 ( .B1(n9436), .B2(n9398), .A(n9232), .ZN(P1_U3266) );
  XOR2_X1 U10452 ( .A(n9233), .B(n9236), .Z(n9441) );
  AOI21_X1 U10453 ( .B1(n9236), .B2(n9235), .A(n9234), .ZN(n9237) );
  OAI222_X1 U10454 ( .A1(n9796), .A2(n9238), .B1(n9798), .B2(n9265), .C1(n9802), .C2(n9237), .ZN(n9437) );
  AOI211_X1 U10455 ( .C1(n9439), .C2(n9251), .A(n9963), .B(n4506), .ZN(n9438)
         );
  NAND2_X1 U10456 ( .A1(n9438), .A2(n9355), .ZN(n9242) );
  AOI22_X1 U10457 ( .A1(n9240), .A2(n9316), .B1(n9806), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n9241) );
  OAI211_X1 U10458 ( .C1(n9243), .C2(n9404), .A(n9242), .B(n9241), .ZN(n9244)
         );
  AOI21_X1 U10459 ( .B1(n9437), .B2(n9792), .A(n9244), .ZN(n9245) );
  OAI21_X1 U10460 ( .B1(n9441), .B2(n9398), .A(n9245), .ZN(P1_U3267) );
  XNOR2_X1 U10461 ( .A(n9246), .B(n9247), .ZN(n9446) );
  XNOR2_X1 U10462 ( .A(n9248), .B(n9247), .ZN(n9249) );
  OAI222_X1 U10463 ( .A1(n9796), .A2(n9250), .B1(n9798), .B2(n9285), .C1(n9802), .C2(n9249), .ZN(n9442) );
  INV_X1 U10464 ( .A(n9266), .ZN(n9252) );
  AOI211_X1 U10465 ( .C1(n9444), .C2(n9252), .A(n9963), .B(n4507), .ZN(n9443)
         );
  NAND2_X1 U10466 ( .A1(n9443), .A2(n9355), .ZN(n9256) );
  INV_X1 U10467 ( .A(n9253), .ZN(n9254) );
  AOI22_X1 U10468 ( .A1(n9806), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9254), .B2(
        n9316), .ZN(n9255) );
  OAI211_X1 U10469 ( .C1(n9257), .C2(n9404), .A(n9256), .B(n9255), .ZN(n9258)
         );
  AOI21_X1 U10470 ( .B1(n9442), .B2(n9792), .A(n9258), .ZN(n9259) );
  OAI21_X1 U10471 ( .B1(n9446), .B2(n9398), .A(n9259), .ZN(P1_U3268) );
  XNOR2_X1 U10472 ( .A(n9260), .B(n9262), .ZN(n9451) );
  NAND2_X1 U10473 ( .A1(n9278), .A2(n9261), .ZN(n9263) );
  XNOR2_X1 U10474 ( .A(n9263), .B(n9262), .ZN(n9264) );
  OAI222_X1 U10475 ( .A1(n9796), .A2(n9265), .B1(n9798), .B2(n9306), .C1(n9264), .C2(n9802), .ZN(n9447) );
  INV_X1 U10476 ( .A(n9286), .ZN(n9267) );
  AOI211_X1 U10477 ( .C1(n9449), .C2(n9267), .A(n9963), .B(n9266), .ZN(n9448)
         );
  NAND2_X1 U10478 ( .A1(n9448), .A2(n9355), .ZN(n9271) );
  INV_X1 U10479 ( .A(n9268), .ZN(n9269) );
  AOI22_X1 U10480 ( .A1(n9806), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9269), .B2(
        n9316), .ZN(n9270) );
  OAI211_X1 U10481 ( .C1(n9272), .C2(n9404), .A(n9271), .B(n9270), .ZN(n9273)
         );
  AOI21_X1 U10482 ( .B1(n9447), .B2(n9792), .A(n9273), .ZN(n9274) );
  OAI21_X1 U10483 ( .B1(n9451), .B2(n9398), .A(n9274), .ZN(P1_U3269) );
  INV_X1 U10484 ( .A(n9275), .ZN(n9277) );
  INV_X1 U10485 ( .A(n9280), .ZN(n9276) );
  OAI21_X1 U10486 ( .B1(n9277), .B2(n9276), .A(n4370), .ZN(n9456) );
  INV_X1 U10487 ( .A(n9278), .ZN(n9282) );
  AOI21_X1 U10488 ( .B1(n9279), .B2(n9303), .A(n9280), .ZN(n9281) );
  NOR2_X1 U10489 ( .A1(n9282), .A2(n9281), .ZN(n9283) );
  OAI222_X1 U10490 ( .A1(n9796), .A2(n9285), .B1(n9798), .B2(n9284), .C1(n9802), .C2(n9283), .ZN(n9452) );
  AOI211_X1 U10491 ( .C1(n9454), .C2(n9294), .A(n9963), .B(n9286), .ZN(n9453)
         );
  NAND2_X1 U10492 ( .A1(n9453), .A2(n9355), .ZN(n9289) );
  AOI22_X1 U10493 ( .A1(n9806), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9287), .B2(
        n9316), .ZN(n9288) );
  OAI211_X1 U10494 ( .C1(n9290), .C2(n9404), .A(n9289), .B(n9288), .ZN(n9291)
         );
  AOI21_X1 U10495 ( .B1(n9452), .B2(n9792), .A(n9291), .ZN(n9292) );
  OAI21_X1 U10496 ( .B1(n9456), .B2(n9398), .A(n9292), .ZN(P1_U3270) );
  XOR2_X1 U10497 ( .A(n9300), .B(n9293), .Z(n9461) );
  INV_X1 U10498 ( .A(n9294), .ZN(n9295) );
  AOI21_X1 U10499 ( .B1(n9457), .B2(n9312), .A(n9295), .ZN(n9458) );
  INV_X1 U10500 ( .A(n9296), .ZN(n9297) );
  AOI22_X1 U10501 ( .A1(n9806), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9297), .B2(
        n9316), .ZN(n9298) );
  OAI21_X1 U10502 ( .B1(n9299), .B2(n9404), .A(n9298), .ZN(n9310) );
  INV_X1 U10503 ( .A(n9279), .ZN(n9304) );
  NOR2_X1 U10504 ( .A1(n9301), .A2(n9300), .ZN(n9302) );
  AOI211_X1 U10505 ( .C1(n9304), .C2(n9303), .A(n9802), .B(n9302), .ZN(n9308)
         );
  OAI22_X1 U10506 ( .A1(n9306), .A2(n9796), .B1(n9305), .B2(n9798), .ZN(n9307)
         );
  NOR2_X1 U10507 ( .A1(n9308), .A2(n9307), .ZN(n9460) );
  NOR2_X1 U10508 ( .A1(n9460), .A2(n9806), .ZN(n9309) );
  AOI211_X1 U10509 ( .C1(n9458), .C2(n9787), .A(n9310), .B(n9309), .ZN(n9311)
         );
  OAI21_X1 U10510 ( .B1(n9461), .B2(n9398), .A(n9311), .ZN(P1_U3271) );
  XNOR2_X1 U10511 ( .A(n4372), .B(n9320), .ZN(n9466) );
  INV_X1 U10512 ( .A(n9338), .ZN(n9314) );
  INV_X1 U10513 ( .A(n9312), .ZN(n9313) );
  AOI21_X1 U10514 ( .B1(n9462), .B2(n9314), .A(n9313), .ZN(n9463) );
  INV_X1 U10515 ( .A(n9315), .ZN(n9317) );
  AOI22_X1 U10516 ( .A1(n9806), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9317), .B2(
        n9316), .ZN(n9318) );
  OAI21_X1 U10517 ( .B1(n9319), .B2(n9404), .A(n9318), .ZN(n9326) );
  XNOR2_X1 U10518 ( .A(n9321), .B(n9320), .ZN(n9324) );
  AOI222_X1 U10519 ( .A1(n9768), .A2(n9324), .B1(n9323), .B2(n9771), .C1(n9322), .C2(n9772), .ZN(n9465) );
  NOR2_X1 U10520 ( .A1(n9465), .A2(n9806), .ZN(n9325) );
  AOI211_X1 U10521 ( .C1(n9463), .C2(n9787), .A(n9326), .B(n9325), .ZN(n9327)
         );
  OAI21_X1 U10522 ( .B1(n9466), .B2(n9398), .A(n9327), .ZN(P1_U3272) );
  INV_X1 U10523 ( .A(n9328), .ZN(n9329) );
  NOR2_X1 U10524 ( .A1(n9330), .A2(n9329), .ZN(n9331) );
  XNOR2_X1 U10525 ( .A(n9331), .B(n9335), .ZN(n9334) );
  AOI222_X1 U10526 ( .A1(n9768), .A2(n9334), .B1(n9333), .B2(n9771), .C1(n9332), .C2(n9772), .ZN(n9471) );
  NAND2_X1 U10527 ( .A1(n9336), .A2(n9335), .ZN(n9467) );
  NAND3_X1 U10528 ( .A1(n4649), .A2(n9337), .A3(n9467), .ZN(n9345) );
  AOI21_X1 U10529 ( .B1(n9468), .B2(n9349), .A(n9338), .ZN(n9469) );
  INV_X1 U10530 ( .A(n9468), .ZN(n9339) );
  NOR2_X1 U10531 ( .A1(n9339), .A2(n9404), .ZN(n9343) );
  OAI22_X1 U10532 ( .A1(n9792), .A2(n9341), .B1(n9340), .B2(n9789), .ZN(n9342)
         );
  AOI211_X1 U10533 ( .C1(n9469), .C2(n9787), .A(n9343), .B(n9342), .ZN(n9344)
         );
  OAI211_X1 U10534 ( .C1(n9806), .C2(n9471), .A(n9345), .B(n9344), .ZN(
        P1_U3273) );
  XNOR2_X1 U10535 ( .A(n9348), .B(n9347), .ZN(n9478) );
  INV_X1 U10536 ( .A(n9349), .ZN(n9350) );
  AOI211_X1 U10537 ( .C1(n9476), .C2(n9365), .A(n9963), .B(n9350), .ZN(n9475)
         );
  NOR2_X1 U10538 ( .A1(n9351), .A2(n9404), .ZN(n9354) );
  OAI22_X1 U10539 ( .A1(n9792), .A2(n9069), .B1(n9352), .B2(n9789), .ZN(n9353)
         );
  AOI211_X1 U10540 ( .C1(n9475), .C2(n9355), .A(n9354), .B(n9353), .ZN(n9362)
         );
  XNOR2_X1 U10541 ( .A(n9357), .B(n9356), .ZN(n9358) );
  OAI222_X1 U10542 ( .A1(n9796), .A2(n9360), .B1(n9798), .B2(n9359), .C1(n9358), .C2(n9802), .ZN(n9474) );
  NAND2_X1 U10543 ( .A1(n9474), .A2(n9792), .ZN(n9361) );
  OAI211_X1 U10544 ( .C1(n9478), .C2(n9398), .A(n9362), .B(n9361), .ZN(
        P1_U3274) );
  XNOR2_X1 U10545 ( .A(n9363), .B(n9364), .ZN(n9483) );
  INV_X1 U10546 ( .A(n9365), .ZN(n9366) );
  AOI211_X1 U10547 ( .C1(n9481), .C2(n4374), .A(n9963), .B(n9366), .ZN(n9480)
         );
  NOR2_X1 U10548 ( .A1(n4502), .A2(n9404), .ZN(n9370) );
  OAI22_X1 U10549 ( .A1(n9792), .A2(n9368), .B1(n9367), .B2(n9789), .ZN(n9369)
         );
  AOI211_X1 U10550 ( .C1(n9480), .C2(n9371), .A(n9370), .B(n9369), .ZN(n9378)
         );
  XNOR2_X1 U10551 ( .A(n9373), .B(n9372), .ZN(n9374) );
  OAI222_X1 U10552 ( .A1(n9796), .A2(n9376), .B1(n9798), .B2(n9375), .C1(n9374), .C2(n9802), .ZN(n9479) );
  NAND2_X1 U10553 ( .A1(n9479), .A2(n9792), .ZN(n9377) );
  OAI211_X1 U10554 ( .C1(n9483), .C2(n9398), .A(n9378), .B(n9377), .ZN(
        P1_U3275) );
  XNOR2_X1 U10555 ( .A(n9380), .B(n9379), .ZN(n9822) );
  INV_X1 U10556 ( .A(n9822), .ZN(n9399) );
  AND2_X1 U10557 ( .A1(n9382), .A2(n9381), .ZN(n9383) );
  OAI21_X1 U10558 ( .B1(n9384), .B2(n9383), .A(n9768), .ZN(n9387) );
  AOI22_X1 U10559 ( .A1(n9385), .A2(n9771), .B1(n9772), .B2(n9770), .ZN(n9386)
         );
  NAND2_X1 U10560 ( .A1(n9387), .A2(n9386), .ZN(n9821) );
  OR2_X1 U10561 ( .A1(n9388), .A2(n9818), .ZN(n9389) );
  NAND2_X1 U10562 ( .A1(n4374), .A2(n9389), .ZN(n9819) );
  OAI22_X1 U10563 ( .A1(n9792), .A2(n9391), .B1(n9390), .B2(n9789), .ZN(n9392)
         );
  AOI21_X1 U10564 ( .B1(n9393), .B2(n9810), .A(n9392), .ZN(n9394) );
  OAI21_X1 U10565 ( .B1(n9819), .B2(n9395), .A(n9394), .ZN(n9396) );
  AOI21_X1 U10566 ( .B1(n9821), .B2(n9792), .A(n9396), .ZN(n9397) );
  OAI21_X1 U10567 ( .B1(n9399), .B2(n9398), .A(n9397), .ZN(P1_U3276) );
  MUX2_X1 U10568 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9400), .S(n9792), .Z(n9401)
         );
  INV_X1 U10569 ( .A(n9401), .ZN(n9410) );
  OAI22_X1 U10570 ( .A1(n9404), .A2(n9403), .B1(n9789), .B2(n9402), .ZN(n9405)
         );
  AOI21_X1 U10571 ( .B1(n9787), .B2(n9406), .A(n9405), .ZN(n9409) );
  NAND2_X1 U10572 ( .A1(n9407), .A2(n9788), .ZN(n9408) );
  NAND3_X1 U10573 ( .A1(n9410), .A2(n9409), .A3(n9408), .ZN(P1_U3289) );
  NAND2_X1 U10574 ( .A1(n9411), .A2(n9967), .ZN(n9417) );
  NAND2_X1 U10575 ( .A1(n9417), .A2(n9416), .ZN(n9489) );
  MUX2_X1 U10576 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9489), .S(n9980), .Z(
        P1_U3552) );
  MUX2_X1 U10577 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9490), .S(n9980), .Z(
        P1_U3551) );
  AOI22_X1 U10578 ( .A1(n9423), .A2(n9816), .B1(n9935), .B2(n9422), .ZN(n9424)
         );
  OAI211_X1 U10579 ( .C1(n9426), .C2(n9932), .A(n9425), .B(n9424), .ZN(n9491)
         );
  MUX2_X1 U10580 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9491), .S(n9980), .Z(
        P1_U3550) );
  OAI21_X1 U10581 ( .B1(n9431), .B2(n9932), .A(n9430), .ZN(n9492) );
  MUX2_X1 U10582 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9492), .S(n9980), .Z(
        P1_U3549) );
  AOI211_X1 U10583 ( .C1(n9935), .C2(n9434), .A(n9433), .B(n9432), .ZN(n9435)
         );
  OAI21_X1 U10584 ( .B1(n9436), .B2(n9932), .A(n9435), .ZN(n9493) );
  MUX2_X1 U10585 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9493), .S(n9980), .Z(
        P1_U3548) );
  AOI211_X1 U10586 ( .C1(n9935), .C2(n9439), .A(n9438), .B(n9437), .ZN(n9440)
         );
  OAI21_X1 U10587 ( .B1(n9441), .B2(n9932), .A(n9440), .ZN(n9494) );
  MUX2_X1 U10588 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9494), .S(n9980), .Z(
        P1_U3547) );
  AOI211_X1 U10589 ( .C1(n9935), .C2(n9444), .A(n9443), .B(n9442), .ZN(n9445)
         );
  OAI21_X1 U10590 ( .B1(n9446), .B2(n9932), .A(n9445), .ZN(n9495) );
  MUX2_X1 U10591 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9495), .S(n9980), .Z(
        P1_U3546) );
  AOI211_X1 U10592 ( .C1(n9935), .C2(n9449), .A(n9448), .B(n9447), .ZN(n9450)
         );
  OAI21_X1 U10593 ( .B1(n9451), .B2(n9932), .A(n9450), .ZN(n9496) );
  MUX2_X1 U10594 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9496), .S(n9980), .Z(
        P1_U3545) );
  AOI211_X1 U10595 ( .C1(n9935), .C2(n9454), .A(n9453), .B(n9452), .ZN(n9455)
         );
  OAI21_X1 U10596 ( .B1(n9456), .B2(n9932), .A(n9455), .ZN(n9497) );
  MUX2_X1 U10597 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9497), .S(n9980), .Z(
        P1_U3544) );
  AOI22_X1 U10598 ( .A1(n9458), .A2(n9816), .B1(n9935), .B2(n9457), .ZN(n9459)
         );
  OAI211_X1 U10599 ( .C1(n9461), .C2(n9932), .A(n9460), .B(n9459), .ZN(n9498)
         );
  MUX2_X1 U10600 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9498), .S(n9980), .Z(
        P1_U3543) );
  AOI22_X1 U10601 ( .A1(n9463), .A2(n9816), .B1(n9935), .B2(n9462), .ZN(n9464)
         );
  OAI211_X1 U10602 ( .C1(n9466), .C2(n9932), .A(n9465), .B(n9464), .ZN(n9499)
         );
  MUX2_X1 U10603 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9499), .S(n9980), .Z(
        P1_U3542) );
  NAND2_X1 U10604 ( .A1(n9467), .A2(n9967), .ZN(n9472) );
  AOI22_X1 U10605 ( .A1(n9469), .A2(n9816), .B1(n9935), .B2(n9468), .ZN(n9470)
         );
  OAI211_X1 U10606 ( .C1(n9473), .C2(n9472), .A(n9471), .B(n9470), .ZN(n9500)
         );
  MUX2_X1 U10607 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9500), .S(n9980), .Z(
        P1_U3541) );
  AOI211_X1 U10608 ( .C1(n9935), .C2(n9476), .A(n9475), .B(n9474), .ZN(n9477)
         );
  OAI21_X1 U10609 ( .B1(n9478), .B2(n9932), .A(n9477), .ZN(n9501) );
  MUX2_X1 U10610 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9501), .S(n9980), .Z(
        P1_U3540) );
  AOI211_X1 U10611 ( .C1(n9935), .C2(n9481), .A(n9480), .B(n9479), .ZN(n9482)
         );
  OAI21_X1 U10612 ( .B1(n9483), .B2(n9932), .A(n9482), .ZN(n9502) );
  MUX2_X1 U10613 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9502), .S(n9980), .Z(
        P1_U3539) );
  AOI211_X1 U10614 ( .C1(n9935), .C2(n9486), .A(n9485), .B(n9484), .ZN(n9487)
         );
  OAI21_X1 U10615 ( .B1(n9488), .B2(n9932), .A(n9487), .ZN(n9503) );
  MUX2_X1 U10616 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9503), .S(n9980), .Z(
        P1_U3537) );
  MUX2_X1 U10617 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9489), .S(n9971), .Z(
        P1_U3520) );
  MUX2_X1 U10618 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9490), .S(n9971), .Z(
        P1_U3519) );
  MUX2_X1 U10619 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9491), .S(n9971), .Z(
        P1_U3518) );
  MUX2_X1 U10620 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9492), .S(n9971), .Z(
        P1_U3517) );
  MUX2_X1 U10621 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9493), .S(n9971), .Z(
        P1_U3516) );
  MUX2_X1 U10622 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9494), .S(n9971), .Z(
        P1_U3515) );
  MUX2_X1 U10623 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9495), .S(n9971), .Z(
        P1_U3514) );
  MUX2_X1 U10624 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9496), .S(n9971), .Z(
        P1_U3513) );
  MUX2_X1 U10625 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9497), .S(n9971), .Z(
        P1_U3512) );
  MUX2_X1 U10626 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9498), .S(n9971), .Z(
        P1_U3511) );
  MUX2_X1 U10627 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9499), .S(n9971), .Z(
        P1_U3510) );
  MUX2_X1 U10628 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9500), .S(n9971), .Z(
        P1_U3508) );
  MUX2_X1 U10629 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9501), .S(n9971), .Z(
        P1_U3505) );
  MUX2_X1 U10630 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9502), .S(n9971), .Z(
        P1_U3502) );
  MUX2_X1 U10631 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9503), .S(n9971), .Z(
        P1_U3496) );
  NAND2_X1 U10632 ( .A1(n9505), .A2(n9504), .ZN(n9926) );
  MUX2_X1 U10633 ( .A(n9506), .B(P1_D_REG_0__SCAN_IN), .S(n9926), .Z(P1_U3440)
         );
  NOR4_X1 U10634 ( .A1(n9508), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9507), .ZN(n9509) );
  AOI21_X1 U10635 ( .B1(n9510), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9509), .ZN(
        n9511) );
  OAI21_X1 U10636 ( .B1(n9513), .B2(n9512), .A(n9511), .ZN(P1_U3322) );
  MUX2_X1 U10637 ( .A(n9514), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10638 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10107) );
  NOR2_X1 U10639 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9515) );
  AOI21_X1 U10640 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9515), .ZN(n10077) );
  NOR2_X1 U10641 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9516) );
  AOI21_X1 U10642 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9516), .ZN(n10080) );
  NOR2_X1 U10643 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9517) );
  AOI21_X1 U10644 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9517), .ZN(n10083) );
  NOR2_X1 U10645 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9518) );
  AOI21_X1 U10646 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9518), .ZN(n10086) );
  NOR2_X1 U10647 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9519) );
  AOI21_X1 U10648 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9519), .ZN(n10089) );
  INV_X1 U10649 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9881) );
  NOR2_X1 U10650 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9526) );
  XOR2_X1 U10651 ( .A(n9866), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10117) );
  NAND2_X1 U10652 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9524) );
  XOR2_X1 U10653 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10115) );
  NAND2_X1 U10654 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9522) );
  XNOR2_X1 U10655 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n9520), .ZN(n10103) );
  AOI21_X1 U10656 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10070) );
  NAND3_X1 U10657 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10072) );
  OAI21_X1 U10658 ( .B1(n10070), .B2(n10074), .A(n10072), .ZN(n10102) );
  NAND2_X1 U10659 ( .A1(n10103), .A2(n10102), .ZN(n9521) );
  NAND2_X1 U10660 ( .A1(n9522), .A2(n9521), .ZN(n10114) );
  NAND2_X1 U10661 ( .A1(n10115), .A2(n10114), .ZN(n9523) );
  NAND2_X1 U10662 ( .A1(n9524), .A2(n9523), .ZN(n10116) );
  NAND2_X1 U10663 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10112), .ZN(n9527) );
  NOR2_X1 U10664 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10112), .ZN(n10111) );
  NAND2_X1 U10665 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n9528), .ZN(n9530) );
  XOR2_X1 U10666 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n9528), .Z(n10110) );
  NAND2_X1 U10667 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10110), .ZN(n9529) );
  NAND2_X1 U10668 ( .A1(n9530), .A2(n9529), .ZN(n9531) );
  NAND2_X1 U10669 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9531), .ZN(n9533) );
  XOR2_X1 U10670 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9531), .Z(n10109) );
  NAND2_X1 U10671 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10109), .ZN(n9532) );
  NAND2_X1 U10672 ( .A1(n9533), .A2(n9532), .ZN(n9534) );
  NAND2_X1 U10673 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9534), .ZN(n9536) );
  XOR2_X1 U10674 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9534), .Z(n10104) );
  NAND2_X1 U10675 ( .A1(n10104), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n9535) );
  NAND2_X1 U10676 ( .A1(n9536), .A2(n9535), .ZN(n9537) );
  AND2_X1 U10677 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9537), .ZN(n9538) );
  XNOR2_X1 U10678 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9537), .ZN(n10101) );
  NAND2_X1 U10679 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9539) );
  OAI21_X1 U10680 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9539), .ZN(n10097) );
  NAND2_X1 U10681 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9540) );
  OAI21_X1 U10682 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9540), .ZN(n10094) );
  NOR2_X1 U10683 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9541) );
  AOI21_X1 U10684 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9541), .ZN(n10091) );
  NAND2_X1 U10685 ( .A1(n10092), .A2(n10091), .ZN(n10090) );
  OAI21_X1 U10686 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10090), .ZN(n10088) );
  NAND2_X1 U10687 ( .A1(n10089), .A2(n10088), .ZN(n10087) );
  OAI21_X1 U10688 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10087), .ZN(n10085) );
  NAND2_X1 U10689 ( .A1(n10086), .A2(n10085), .ZN(n10084) );
  OAI21_X1 U10690 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10084), .ZN(n10082) );
  NAND2_X1 U10691 ( .A1(n10083), .A2(n10082), .ZN(n10081) );
  OAI21_X1 U10692 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10081), .ZN(n10079) );
  NAND2_X1 U10693 ( .A1(n10080), .A2(n10079), .ZN(n10078) );
  OAI21_X1 U10694 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10078), .ZN(n10076) );
  NAND2_X1 U10695 ( .A1(n10077), .A2(n10076), .ZN(n10075) );
  OAI21_X1 U10696 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10075), .ZN(n10106) );
  NOR2_X1 U10697 ( .A1(n10107), .A2(n10106), .ZN(n9542) );
  NAND2_X1 U10698 ( .A1(n10107), .A2(n10106), .ZN(n10105) );
  OAI21_X1 U10699 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n9542), .A(n10105), .ZN(
        n9729) );
  AOI22_X1 U10700 ( .A1(SI_31_), .A2(keyinput_f1), .B1(SI_14_), .B2(
        keyinput_f18), .ZN(n9543) );
  OAI221_X1 U10701 ( .B1(SI_31_), .B2(keyinput_f1), .C1(SI_14_), .C2(
        keyinput_f18), .A(n9543), .ZN(n9550) );
  AOI22_X1 U10702 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(SI_0_), .B2(keyinput_f32), .ZN(n9544) );
  OAI221_X1 U10703 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        SI_0_), .C2(keyinput_f32), .A(n9544), .ZN(n9549) );
  AOI22_X1 U10704 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_f42), .B1(SI_9_), .B2(keyinput_f23), .ZN(n9545) );
  OAI221_X1 U10705 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .C1(
        SI_9_), .C2(keyinput_f23), .A(n9545), .ZN(n9548) );
  AOI22_X1 U10706 ( .A1(SI_12_), .A2(keyinput_f20), .B1(SI_20_), .B2(
        keyinput_f12), .ZN(n9546) );
  OAI221_X1 U10707 ( .B1(SI_12_), .B2(keyinput_f20), .C1(SI_20_), .C2(
        keyinput_f12), .A(n9546), .ZN(n9547) );
  NOR4_X1 U10708 ( .A1(n9550), .A2(n9549), .A3(n9548), .A4(n9547), .ZN(n9578)
         );
  XOR2_X1 U10709 ( .A(n7712), .B(keyinput_f38), .Z(n9557) );
  AOI22_X1 U10710 ( .A1(SI_2_), .A2(keyinput_f30), .B1(n5939), .B2(
        keyinput_f63), .ZN(n9551) );
  OAI221_X1 U10711 ( .B1(SI_2_), .B2(keyinput_f30), .C1(n5939), .C2(
        keyinput_f63), .A(n9551), .ZN(n9556) );
  AOI22_X1 U10712 ( .A1(SI_11_), .A2(keyinput_f21), .B1(SI_16_), .B2(
        keyinput_f16), .ZN(n9552) );
  OAI221_X1 U10713 ( .B1(SI_11_), .B2(keyinput_f21), .C1(SI_16_), .C2(
        keyinput_f16), .A(n9552), .ZN(n9555) );
  AOI22_X1 U10714 ( .A1(SI_7_), .A2(keyinput_f25), .B1(SI_24_), .B2(
        keyinput_f8), .ZN(n9553) );
  OAI221_X1 U10715 ( .B1(SI_7_), .B2(keyinput_f25), .C1(SI_24_), .C2(
        keyinput_f8), .A(n9553), .ZN(n9554) );
  NOR4_X1 U10716 ( .A1(n9557), .A2(n9556), .A3(n9555), .A4(n9554), .ZN(n9577)
         );
  AOI22_X1 U10717 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(n7738), 
        .B2(keyinput_f47), .ZN(n9558) );
  OAI221_X1 U10718 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(n7738), .C2(keyinput_f47), .A(n9558), .ZN(n9566) );
  AOI22_X1 U10719 ( .A1(SI_30_), .A2(keyinput_f2), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(keyinput_f59), .ZN(n9559) );
  OAI221_X1 U10720 ( .B1(SI_30_), .B2(keyinput_f2), .C1(P2_REG3_REG_2__SCAN_IN), .C2(keyinput_f59), .A(n9559), .ZN(n9565) );
  AOI22_X1 U10721 ( .A1(SI_25_), .A2(keyinput_f7), .B1(SI_27_), .B2(
        keyinput_f5), .ZN(n9560) );
  OAI221_X1 U10722 ( .B1(SI_25_), .B2(keyinput_f7), .C1(SI_27_), .C2(
        keyinput_f5), .A(n9560), .ZN(n9564) );
  XNOR2_X1 U10723 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_f62), .ZN(n9562)
         );
  XNOR2_X1 U10724 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_f54), .ZN(n9561)
         );
  NAND2_X1 U10725 ( .A1(n9562), .A2(n9561), .ZN(n9563) );
  NOR4_X1 U10726 ( .A1(n9566), .A2(n9565), .A3(n9564), .A4(n9563), .ZN(n9576)
         );
  AOI22_X1 U10727 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_f52), .B1(SI_6_), 
        .B2(keyinput_f26), .ZN(n9567) );
  OAI221_X1 U10728 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .C1(SI_6_), .C2(keyinput_f26), .A(n9567), .ZN(n9574) );
  AOI22_X1 U10729 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_f60), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .ZN(n9568) );
  OAI221_X1 U10730 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_f34), .A(n9568), .ZN(n9573) );
  AOI22_X1 U10731 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_f53), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput_f37), .ZN(n9569) );
  OAI221_X1 U10732 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_f37), .A(n9569), .ZN(n9572) );
  AOI22_X1 U10733 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_f45), .B1(
        SI_21_), .B2(keyinput_f11), .ZN(n9570) );
  OAI221_X1 U10734 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .C1(
        SI_21_), .C2(keyinput_f11), .A(n9570), .ZN(n9571) );
  NOR4_X1 U10735 ( .A1(n9574), .A2(n9573), .A3(n9572), .A4(n9571), .ZN(n9575)
         );
  NAND4_X1 U10736 ( .A1(n9578), .A2(n9577), .A3(n9576), .A4(n9575), .ZN(n9628)
         );
  AOI22_X1 U10737 ( .A1(n9580), .A2(keyinput_f10), .B1(keyinput_f51), .B2(
        n9673), .ZN(n9579) );
  OAI221_X1 U10738 ( .B1(n9580), .B2(keyinput_f10), .C1(n9673), .C2(
        keyinput_f51), .A(n9579), .ZN(n9589) );
  AOI22_X1 U10739 ( .A1(n9582), .A2(keyinput_f48), .B1(keyinput_f3), .B2(n7582), .ZN(n9581) );
  OAI221_X1 U10740 ( .B1(n9582), .B2(keyinput_f48), .C1(n7582), .C2(
        keyinput_f3), .A(n9581), .ZN(n9588) );
  AOI22_X1 U10741 ( .A1(n9642), .A2(keyinput_f55), .B1(keyinput_f56), .B2(
        n9633), .ZN(n9583) );
  OAI221_X1 U10742 ( .B1(n9642), .B2(keyinput_f55), .C1(n9633), .C2(
        keyinput_f56), .A(n9583), .ZN(n9587) );
  XOR2_X1 U10743 ( .A(n6084), .B(keyinput_f36), .Z(n9585) );
  XNOR2_X1 U10744 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_f44), .ZN(n9584)
         );
  NAND2_X1 U10745 ( .A1(n9585), .A2(n9584), .ZN(n9586) );
  NOR4_X1 U10746 ( .A1(n9589), .A2(n9588), .A3(n9587), .A4(n9586), .ZN(n9626)
         );
  AOI22_X1 U10747 ( .A1(n9591), .A2(keyinput_f9), .B1(keyinput_f35), .B2(n5852), .ZN(n9590) );
  OAI221_X1 U10748 ( .B1(n9591), .B2(keyinput_f9), .C1(n5852), .C2(
        keyinput_f35), .A(n9590), .ZN(n9600) );
  AOI22_X1 U10749 ( .A1(n9593), .A2(keyinput_f6), .B1(keyinput_f41), .B2(n5996), .ZN(n9592) );
  OAI221_X1 U10750 ( .B1(n9593), .B2(keyinput_f6), .C1(n5996), .C2(
        keyinput_f41), .A(n9592), .ZN(n9599) );
  XNOR2_X1 U10751 ( .A(SI_18_), .B(keyinput_f14), .ZN(n9597) );
  XNOR2_X1 U10752 ( .A(SI_3_), .B(keyinput_f29), .ZN(n9596) );
  XNOR2_X1 U10753 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_f33), .ZN(n9595) );
  XNOR2_X1 U10754 ( .A(SI_5_), .B(keyinput_f27), .ZN(n9594) );
  NAND4_X1 U10755 ( .A1(n9597), .A2(n9596), .A3(n9595), .A4(n9594), .ZN(n9598)
         );
  NOR3_X1 U10756 ( .A1(n9600), .A2(n9599), .A3(n9598), .ZN(n9625) );
  INV_X1 U10757 ( .A(SI_13_), .ZN(n9634) );
  INV_X1 U10758 ( .A(SI_15_), .ZN(n9602) );
  AOI22_X1 U10759 ( .A1(n9634), .A2(keyinput_f19), .B1(n9602), .B2(
        keyinput_f17), .ZN(n9601) );
  OAI221_X1 U10760 ( .B1(n9634), .B2(keyinput_f19), .C1(n9602), .C2(
        keyinput_f17), .A(n9601), .ZN(n9612) );
  AOI22_X1 U10761 ( .A1(n6561), .A2(keyinput_f49), .B1(n9604), .B2(
        keyinput_f39), .ZN(n9603) );
  OAI221_X1 U10762 ( .B1(n6561), .B2(keyinput_f49), .C1(n9604), .C2(
        keyinput_f39), .A(n9603), .ZN(n9611) );
  AOI22_X1 U10763 ( .A1(n9606), .A2(keyinput_f57), .B1(keyinput_f50), .B2(
        n9661), .ZN(n9605) );
  OAI221_X1 U10764 ( .B1(n9606), .B2(keyinput_f57), .C1(n9661), .C2(
        keyinput_f50), .A(n9605), .ZN(n9610) );
  XNOR2_X1 U10765 ( .A(SI_1_), .B(keyinput_f31), .ZN(n9608) );
  XNOR2_X1 U10766 ( .A(SI_4_), .B(keyinput_f28), .ZN(n9607) );
  NAND2_X1 U10767 ( .A1(n9608), .A2(n9607), .ZN(n9609) );
  NOR4_X1 U10768 ( .A1(n9612), .A2(n9611), .A3(n9610), .A4(n9609), .ZN(n9624)
         );
  INV_X1 U10769 ( .A(SI_19_), .ZN(n9614) );
  INV_X1 U10770 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9852) );
  AOI22_X1 U10771 ( .A1(n9614), .A2(keyinput_f13), .B1(keyinput_f0), .B2(n9852), .ZN(n9613) );
  OAI221_X1 U10772 ( .B1(n9614), .B2(keyinput_f13), .C1(n9852), .C2(
        keyinput_f0), .A(n9613), .ZN(n9622) );
  AOI22_X1 U10773 ( .A1(n6098), .A2(keyinput_f4), .B1(keyinput_f61), .B2(n9694), .ZN(n9615) );
  OAI221_X1 U10774 ( .B1(n6098), .B2(keyinput_f4), .C1(n9694), .C2(
        keyinput_f61), .A(n9615), .ZN(n9621) );
  AOI22_X1 U10775 ( .A1(n9659), .A2(keyinput_f43), .B1(n9651), .B2(
        keyinput_f22), .ZN(n9616) );
  OAI221_X1 U10776 ( .B1(n9659), .B2(keyinput_f43), .C1(n9651), .C2(
        keyinput_f22), .A(n9616), .ZN(n9620) );
  AOI22_X1 U10777 ( .A1(n7407), .A2(keyinput_f58), .B1(n9618), .B2(
        keyinput_f15), .ZN(n9617) );
  OAI221_X1 U10778 ( .B1(n7407), .B2(keyinput_f58), .C1(n9618), .C2(
        keyinput_f15), .A(n9617), .ZN(n9619) );
  NOR4_X1 U10779 ( .A1(n9622), .A2(n9621), .A3(n9620), .A4(n9619), .ZN(n9623)
         );
  NAND4_X1 U10780 ( .A1(n9626), .A2(n9625), .A3(n9624), .A4(n9623), .ZN(n9627)
         );
  OAI22_X1 U10781 ( .A1(keyinput_f24), .A2(n9727), .B1(n9628), .B2(n9627), 
        .ZN(n9629) );
  AOI21_X1 U10782 ( .B1(keyinput_f24), .B2(n9727), .A(n9629), .ZN(n9726) );
  AOI22_X1 U10783 ( .A1(n7712), .A2(keyinput_g38), .B1(keyinput_g58), .B2(
        n7407), .ZN(n9630) );
  OAI221_X1 U10784 ( .B1(n7712), .B2(keyinput_g38), .C1(n7407), .C2(
        keyinput_g58), .A(n9630), .ZN(n9640) );
  AOI22_X1 U10785 ( .A1(n6098), .A2(keyinput_g4), .B1(keyinput_g49), .B2(n6561), .ZN(n9631) );
  OAI221_X1 U10786 ( .B1(n6098), .B2(keyinput_g4), .C1(n6561), .C2(
        keyinput_g49), .A(n9631), .ZN(n9639) );
  AOI22_X1 U10787 ( .A1(n9634), .A2(keyinput_g19), .B1(keyinput_g56), .B2(
        n9633), .ZN(n9632) );
  OAI221_X1 U10788 ( .B1(n9634), .B2(keyinput_g19), .C1(n9633), .C2(
        keyinput_g56), .A(n9632), .ZN(n9638) );
  XNOR2_X1 U10789 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_g54), .ZN(n9636)
         );
  XNOR2_X1 U10790 ( .A(SI_11_), .B(keyinput_g21), .ZN(n9635) );
  NAND2_X1 U10791 ( .A1(n9636), .A2(n9635), .ZN(n9637) );
  NOR4_X1 U10792 ( .A1(n9640), .A2(n9639), .A3(n9638), .A4(n9637), .ZN(n9685)
         );
  AOI22_X1 U10793 ( .A1(n9643), .A2(keyinput_g12), .B1(keyinput_g55), .B2(
        n9642), .ZN(n9641) );
  OAI221_X1 U10794 ( .B1(n9643), .B2(keyinput_g12), .C1(n9642), .C2(
        keyinput_g55), .A(n9641), .ZN(n9656) );
  AOI22_X1 U10795 ( .A1(n9646), .A2(keyinput_g11), .B1(n9645), .B2(keyinput_g5), .ZN(n9644) );
  OAI221_X1 U10796 ( .B1(n9646), .B2(keyinput_g11), .C1(n9645), .C2(
        keyinput_g5), .A(n9644), .ZN(n9655) );
  AOI22_X1 U10797 ( .A1(n9649), .A2(keyinput_g27), .B1(keyinput_g45), .B2(
        n9648), .ZN(n9647) );
  OAI221_X1 U10798 ( .B1(n9649), .B2(keyinput_g27), .C1(n9648), .C2(
        keyinput_g45), .A(n9647), .ZN(n9654) );
  INV_X1 U10799 ( .A(SI_12_), .ZN(n9652) );
  AOI22_X1 U10800 ( .A1(n9652), .A2(keyinput_g20), .B1(keyinput_g22), .B2(
        n9651), .ZN(n9650) );
  OAI221_X1 U10801 ( .B1(n9652), .B2(keyinput_g20), .C1(n9651), .C2(
        keyinput_g22), .A(n9650), .ZN(n9653) );
  NOR4_X1 U10802 ( .A1(n9656), .A2(n9655), .A3(n9654), .A4(n9653), .ZN(n9684)
         );
  AOI22_X1 U10803 ( .A1(n9659), .A2(keyinput_g43), .B1(keyinput_g1), .B2(n9658), .ZN(n9657) );
  OAI221_X1 U10804 ( .B1(n9659), .B2(keyinput_g43), .C1(n9658), .C2(
        keyinput_g1), .A(n9657), .ZN(n9669) );
  AOI22_X1 U10805 ( .A1(n6752), .A2(keyinput_g40), .B1(n9661), .B2(
        keyinput_g50), .ZN(n9660) );
  OAI221_X1 U10806 ( .B1(n6752), .B2(keyinput_g40), .C1(n9661), .C2(
        keyinput_g50), .A(n9660), .ZN(n9668) );
  AOI22_X1 U10807 ( .A1(P2_U3152), .A2(keyinput_g34), .B1(n9663), .B2(
        keyinput_g7), .ZN(n9662) );
  OAI221_X1 U10808 ( .B1(P2_U3152), .B2(keyinput_g34), .C1(n9663), .C2(
        keyinput_g7), .A(n9662), .ZN(n9667) );
  XNOR2_X1 U10809 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_g57), .ZN(n9665)
         );
  XNOR2_X1 U10810 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_g44), .ZN(n9664)
         );
  NAND2_X1 U10811 ( .A1(n9665), .A2(n9664), .ZN(n9666) );
  NOR4_X1 U10812 ( .A1(n9669), .A2(n9668), .A3(n9667), .A4(n9666), .ZN(n9683)
         );
  AOI22_X1 U10813 ( .A1(n5852), .A2(keyinput_g35), .B1(keyinput_g52), .B2(
        n9671), .ZN(n9670) );
  OAI221_X1 U10814 ( .B1(n5852), .B2(keyinput_g35), .C1(n9671), .C2(
        keyinput_g52), .A(n9670), .ZN(n9681) );
  AOI22_X1 U10815 ( .A1(n9674), .A2(keyinput_g28), .B1(keyinput_g51), .B2(
        n9673), .ZN(n9672) );
  OAI221_X1 U10816 ( .B1(n9674), .B2(keyinput_g28), .C1(n9673), .C2(
        keyinput_g51), .A(n9672), .ZN(n9680) );
  XOR2_X1 U10817 ( .A(n7738), .B(keyinput_g47), .Z(n9678) );
  XNOR2_X1 U10818 ( .A(SI_1_), .B(keyinput_g31), .ZN(n9677) );
  XNOR2_X1 U10819 ( .A(SI_18_), .B(keyinput_g14), .ZN(n9676) );
  XNOR2_X1 U10820 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_g33), .ZN(n9675) );
  NAND4_X1 U10821 ( .A1(n9678), .A2(n9677), .A3(n9676), .A4(n9675), .ZN(n9679)
         );
  NOR3_X1 U10822 ( .A1(n9681), .A2(n9680), .A3(n9679), .ZN(n9682) );
  NAND4_X1 U10823 ( .A1(n9685), .A2(n9684), .A3(n9683), .A4(n9682), .ZN(n9724)
         );
  AOI22_X1 U10824 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_g39), .B1(
        SI_26_), .B2(keyinput_g6), .ZN(n9686) );
  OAI221_X1 U10825 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .C1(
        SI_26_), .C2(keyinput_g6), .A(n9686), .ZN(n9693) );
  AOI22_X1 U10826 ( .A1(SI_6_), .A2(keyinput_g26), .B1(SI_22_), .B2(
        keyinput_g10), .ZN(n9687) );
  OAI221_X1 U10827 ( .B1(SI_6_), .B2(keyinput_g26), .C1(SI_22_), .C2(
        keyinput_g10), .A(n9687), .ZN(n9692) );
  AOI22_X1 U10828 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_g53), .B1(SI_17_), .B2(keyinput_g15), .ZN(n9688) );
  OAI221_X1 U10829 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_g53), .C1(
        SI_17_), .C2(keyinput_g15), .A(n9688), .ZN(n9691) );
  AOI22_X1 U10830 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_g41), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .ZN(n9689) );
  OAI221_X1 U10831 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_g36), .A(n9689), .ZN(n9690) );
  NOR4_X1 U10832 ( .A1(n9693), .A2(n9692), .A3(n9691), .A4(n9690), .ZN(n9722)
         );
  XNOR2_X1 U10833 ( .A(n9694), .B(keyinput_g61), .ZN(n9701) );
  AOI22_X1 U10834 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_g37), .B1(
        SI_23_), .B2(keyinput_g9), .ZN(n9695) );
  OAI221_X1 U10835 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .C1(
        SI_23_), .C2(keyinput_g9), .A(n9695), .ZN(n9700) );
  AOI22_X1 U10836 ( .A1(SI_14_), .A2(keyinput_g18), .B1(SI_24_), .B2(
        keyinput_g8), .ZN(n9696) );
  OAI221_X1 U10837 ( .B1(SI_14_), .B2(keyinput_g18), .C1(SI_24_), .C2(
        keyinput_g8), .A(n9696), .ZN(n9699) );
  AOI22_X1 U10838 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n9697) );
  OAI221_X1 U10839 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n9697), .ZN(n9698) );
  NOR4_X1 U10840 ( .A1(n9701), .A2(n9700), .A3(n9699), .A4(n9698), .ZN(n9721)
         );
  AOI22_X1 U10841 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(SI_15_), 
        .B2(keyinput_g17), .ZN(n9702) );
  OAI221_X1 U10842 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(SI_15_), 
        .C2(keyinput_g17), .A(n9702), .ZN(n9710) );
  AOI22_X1 U10843 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_g42), .B1(
        SI_19_), .B2(keyinput_g13), .ZN(n9703) );
  OAI221_X1 U10844 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .C1(
        SI_19_), .C2(keyinput_g13), .A(n9703), .ZN(n9709) );
  AOI22_X1 U10845 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_g46), .B1(n9705), .B2(keyinput_g23), .ZN(n9704) );
  OAI221_X1 U10846 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .C1(
        n9705), .C2(keyinput_g23), .A(n9704), .ZN(n9708) );
  AOI22_X1 U10847 ( .A1(SI_30_), .A2(keyinput_g2), .B1(SI_0_), .B2(
        keyinput_g32), .ZN(n9706) );
  OAI221_X1 U10848 ( .B1(SI_30_), .B2(keyinput_g2), .C1(SI_0_), .C2(
        keyinput_g32), .A(n9706), .ZN(n9707) );
  NOR4_X1 U10849 ( .A1(n9710), .A2(n9709), .A3(n9708), .A4(n9707), .ZN(n9720)
         );
  AOI22_X1 U10850 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_g62), .B1(SI_3_), .B2(keyinput_g29), .ZN(n9711) );
  OAI221_X1 U10851 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .C1(
        SI_3_), .C2(keyinput_g29), .A(n9711), .ZN(n9718) );
  AOI22_X1 U10852 ( .A1(SI_2_), .A2(keyinput_g30), .B1(SI_16_), .B2(
        keyinput_g16), .ZN(n9712) );
  OAI221_X1 U10853 ( .B1(SI_2_), .B2(keyinput_g30), .C1(SI_16_), .C2(
        keyinput_g16), .A(n9712), .ZN(n9717) );
  AOI22_X1 U10854 ( .A1(SI_29_), .A2(keyinput_g3), .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n9713) );
  OAI221_X1 U10855 ( .B1(SI_29_), .B2(keyinput_g3), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n9713), .ZN(n9716) );
  AOI22_X1 U10856 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_g48), .B1(SI_7_), .B2(keyinput_g25), .ZN(n9714) );
  OAI221_X1 U10857 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .C1(
        SI_7_), .C2(keyinput_g25), .A(n9714), .ZN(n9715) );
  NOR4_X1 U10858 ( .A1(n9718), .A2(n9717), .A3(n9716), .A4(n9715), .ZN(n9719)
         );
  NAND4_X1 U10859 ( .A1(n9722), .A2(n9721), .A3(n9720), .A4(n9719), .ZN(n9723)
         );
  OAI22_X1 U10860 ( .A1(keyinput_g24), .A2(n9727), .B1(n9724), .B2(n9723), 
        .ZN(n9725) );
  AOI211_X1 U10861 ( .C1(keyinput_g24), .C2(n9727), .A(n9726), .B(n9725), .ZN(
        n9728) );
  XNOR2_X1 U10862 ( .A(n9729), .B(n9728), .ZN(n9733) );
  NOR2_X1 U10863 ( .A1(n9731), .A2(n9730), .ZN(n9732) );
  XOR2_X1 U10864 ( .A(n9733), .B(n9732), .Z(ADD_1071_U4) );
  AOI21_X1 U10865 ( .B1(n9935), .B2(n9735), .A(n9734), .ZN(n9736) );
  OAI211_X1 U10866 ( .C1(n9738), .C2(n9824), .A(n9737), .B(n9736), .ZN(n9739)
         );
  AOI21_X1 U10867 ( .B1(n9805), .B2(n9740), .A(n9739), .ZN(n9742) );
  INV_X1 U10868 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9741) );
  AOI22_X1 U10869 ( .A1(n9971), .A2(n9742), .B1(n9741), .B2(n9969), .ZN(
        P1_U3484) );
  AOI22_X1 U10870 ( .A1(n9980), .A2(n9742), .B1(n5188), .B2(n9978), .ZN(
        P1_U3533) );
  OAI21_X1 U10871 ( .B1(n9743), .B2(n9961), .A(n9813), .ZN(n9744) );
  AOI21_X1 U10872 ( .B1(n9745), .B2(n9816), .A(n9744), .ZN(n9746) );
  AOI22_X1 U10873 ( .A1(n9980), .A2(n9746), .B1(n6291), .B2(n9978), .ZN(
        P1_U3554) );
  AOI22_X1 U10874 ( .A1(n9971), .A2(n9746), .B1(n6288), .B2(n9969), .ZN(
        P1_U3522) );
  NOR2_X1 U10875 ( .A1(n9747), .A2(n6936), .ZN(n9748) );
  INV_X1 U10876 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9750) );
  AOI22_X1 U10877 ( .A1(n10069), .A2(n9756), .B1(n9750), .B2(n10067), .ZN(
        P2_U3551) );
  NOR2_X1 U10878 ( .A1(n9751), .A2(n10050), .ZN(n9752) );
  INV_X1 U10879 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9755) );
  AOI22_X1 U10880 ( .A1(n10069), .A2(n9757), .B1(n9755), .B2(n10067), .ZN(
        P2_U3550) );
  AOI22_X1 U10881 ( .A1(n10055), .A2(n9756), .B1(n6301), .B2(n10054), .ZN(
        P2_U3519) );
  AOI22_X1 U10882 ( .A1(n10055), .A2(n9757), .B1(n6185), .B2(n10054), .ZN(
        P2_U3518) );
  INV_X1 U10883 ( .A(n9766), .ZN(n9759) );
  XNOR2_X1 U10884 ( .A(n9758), .B(n9759), .ZN(n9828) );
  AND2_X1 U10885 ( .A1(n9760), .A2(n9779), .ZN(n9762) );
  OR2_X1 U10886 ( .A1(n9762), .A2(n9761), .ZN(n9826) );
  INV_X1 U10887 ( .A(n9826), .ZN(n9763) );
  AOI22_X1 U10888 ( .A1(n9828), .A2(n9788), .B1(n9787), .B2(n9763), .ZN(n9781)
         );
  NAND2_X1 U10889 ( .A1(n9806), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9764) );
  OAI21_X1 U10890 ( .B1(n9789), .B2(n9765), .A(n9764), .ZN(n9778) );
  XNOR2_X1 U10891 ( .A(n9767), .B(n9766), .ZN(n9769) );
  NAND2_X1 U10892 ( .A1(n9769), .A2(n9768), .ZN(n9775) );
  AOI22_X1 U10893 ( .A1(n9773), .A2(n9772), .B1(n9771), .B2(n9770), .ZN(n9774)
         );
  NAND2_X1 U10894 ( .A1(n9775), .A2(n9774), .ZN(n9776) );
  AOI21_X1 U10895 ( .B1(n9828), .B2(n9805), .A(n9776), .ZN(n9830) );
  NOR2_X1 U10896 ( .A1(n9830), .A2(n9806), .ZN(n9777) );
  AOI211_X1 U10897 ( .C1(n9810), .C2(n9779), .A(n9778), .B(n9777), .ZN(n9780)
         );
  NAND2_X1 U10898 ( .A1(n9781), .A2(n9780), .ZN(P1_U3278) );
  XNOR2_X1 U10899 ( .A(n9782), .B(n9793), .ZN(n9839) );
  OR2_X1 U10900 ( .A1(n9783), .A2(n9836), .ZN(n9784) );
  NAND2_X1 U10901 ( .A1(n9785), .A2(n9784), .ZN(n9837) );
  INV_X1 U10902 ( .A(n9837), .ZN(n9786) );
  AOI22_X1 U10903 ( .A1(n9839), .A2(n9788), .B1(n9787), .B2(n9786), .ZN(n9812)
         );
  OAI22_X1 U10904 ( .A1(n9792), .A2(n9791), .B1(n9790), .B2(n9789), .ZN(n9808)
         );
  INV_X1 U10905 ( .A(n9793), .ZN(n9794) );
  XNOR2_X1 U10906 ( .A(n9795), .B(n9794), .ZN(n9803) );
  OAI22_X1 U10907 ( .A1(n9799), .A2(n9798), .B1(n9797), .B2(n9796), .ZN(n9800)
         );
  INV_X1 U10908 ( .A(n9800), .ZN(n9801) );
  OAI21_X1 U10909 ( .B1(n9803), .B2(n9802), .A(n9801), .ZN(n9804) );
  AOI21_X1 U10910 ( .B1(n9839), .B2(n9805), .A(n9804), .ZN(n9841) );
  NOR2_X1 U10911 ( .A1(n9841), .A2(n9806), .ZN(n9807) );
  AOI211_X1 U10912 ( .C1(n9810), .C2(n9809), .A(n9808), .B(n9807), .ZN(n9811)
         );
  NAND2_X1 U10913 ( .A1(n9812), .A2(n9811), .ZN(P1_U3280) );
  OAI21_X1 U10914 ( .B1(n9814), .B2(n9961), .A(n9813), .ZN(n9815) );
  AOI21_X1 U10915 ( .B1(n9817), .B2(n9816), .A(n9815), .ZN(n9843) );
  AOI22_X1 U10916 ( .A1(n9980), .A2(n9843), .B1(n8833), .B2(n9978), .ZN(
        P1_U3553) );
  OAI22_X1 U10917 ( .A1(n9819), .A2(n9963), .B1(n9818), .B2(n9961), .ZN(n9820)
         );
  AOI211_X1 U10918 ( .C1(n9822), .C2(n9967), .A(n9821), .B(n9820), .ZN(n9845)
         );
  AOI22_X1 U10919 ( .A1(n9980), .A2(n9845), .B1(n9823), .B2(n9978), .ZN(
        P1_U3538) );
  INV_X1 U10920 ( .A(n9824), .ZN(n9960) );
  OAI22_X1 U10921 ( .A1(n9826), .A2(n9963), .B1(n9825), .B2(n9961), .ZN(n9827)
         );
  AOI21_X1 U10922 ( .B1(n9828), .B2(n9960), .A(n9827), .ZN(n9829) );
  AOI22_X1 U10923 ( .A1(n9980), .A2(n9847), .B1(n5271), .B2(n9978), .ZN(
        P1_U3536) );
  OAI21_X1 U10924 ( .B1(n9832), .B2(n9961), .A(n9831), .ZN(n9833) );
  AOI211_X1 U10925 ( .C1(n9835), .C2(n9967), .A(n9834), .B(n9833), .ZN(n9849)
         );
  AOI22_X1 U10926 ( .A1(n9980), .A2(n9849), .B1(n6567), .B2(n9978), .ZN(
        P1_U3535) );
  OAI22_X1 U10927 ( .A1(n9837), .A2(n9963), .B1(n9836), .B2(n9961), .ZN(n9838)
         );
  AOI21_X1 U10928 ( .B1(n9839), .B2(n9960), .A(n9838), .ZN(n9840) );
  AOI22_X1 U10929 ( .A1(n9980), .A2(n9851), .B1(n5206), .B2(n9978), .ZN(
        P1_U3534) );
  INV_X1 U10930 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9842) );
  AOI22_X1 U10931 ( .A1(n9971), .A2(n9843), .B1(n9842), .B2(n9969), .ZN(
        P1_U3521) );
  INV_X1 U10932 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9844) );
  AOI22_X1 U10933 ( .A1(n9971), .A2(n9845), .B1(n9844), .B2(n9969), .ZN(
        P1_U3499) );
  INV_X1 U10934 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9846) );
  AOI22_X1 U10935 ( .A1(n9971), .A2(n9847), .B1(n9846), .B2(n9969), .ZN(
        P1_U3493) );
  INV_X1 U10936 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9848) );
  AOI22_X1 U10937 ( .A1(n9971), .A2(n9849), .B1(n9848), .B2(n9969), .ZN(
        P1_U3490) );
  INV_X1 U10938 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9850) );
  AOI22_X1 U10939 ( .A1(n9971), .A2(n9851), .B1(n9850), .B2(n9969), .ZN(
        P1_U3487) );
  XOR2_X1 U10940 ( .A(n9852), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  OAI21_X1 U10941 ( .B1(n9855), .B2(n9854), .A(n9853), .ZN(n9860) );
  OAI21_X1 U10942 ( .B1(n9858), .B2(n9857), .A(n9856), .ZN(n9859) );
  AOI22_X1 U10943 ( .A1(n9921), .A2(n9860), .B1(n9920), .B2(n9859), .ZN(n9865)
         );
  AOI211_X1 U10944 ( .C1(n9912), .C2(n9863), .A(n9862), .B(n9861), .ZN(n9864)
         );
  OAI211_X1 U10945 ( .C1(n9925), .C2(n9866), .A(n9865), .B(n9864), .ZN(
        P1_U3245) );
  NAND2_X1 U10946 ( .A1(n9912), .A2(n9867), .ZN(n9874) );
  AOI21_X1 U10947 ( .B1(n9870), .B2(n9869), .A(n9868), .ZN(n9872) );
  AOI21_X1 U10948 ( .B1(n9920), .B2(n9872), .A(n9871), .ZN(n9873) );
  AND2_X1 U10949 ( .A1(n9874), .A2(n9873), .ZN(n9880) );
  OAI21_X1 U10950 ( .B1(n9877), .B2(n9876), .A(n9875), .ZN(n9878) );
  NAND2_X1 U10951 ( .A1(n9921), .A2(n9878), .ZN(n9879) );
  OAI211_X1 U10952 ( .C1(n9881), .C2(n9925), .A(n9880), .B(n9879), .ZN(
        P1_U3246) );
  OAI21_X1 U10953 ( .B1(n9884), .B2(n9883), .A(n9882), .ZN(n9891) );
  AOI211_X1 U10954 ( .C1(n9888), .C2(n9887), .A(n9886), .B(n9885), .ZN(n9889)
         );
  AOI211_X1 U10955 ( .C1(n9920), .C2(n9891), .A(n9890), .B(n9889), .ZN(n9894)
         );
  AOI22_X1 U10956 ( .A1(n9906), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n9892), .B2(
        n9912), .ZN(n9893) );
  NAND2_X1 U10957 ( .A1(n9894), .A2(n9893), .ZN(P1_U3247) );
  OAI21_X1 U10958 ( .B1(n9897), .B2(n9896), .A(n9895), .ZN(n9904) );
  AOI211_X1 U10959 ( .C1(n9901), .C2(n9900), .A(n9899), .B(n9898), .ZN(n9902)
         );
  AOI211_X1 U10960 ( .C1(n9921), .C2(n9904), .A(n9903), .B(n9902), .ZN(n9908)
         );
  AOI22_X1 U10961 ( .A1(n9906), .A2(P1_ADDR_REG_8__SCAN_IN), .B1(n9905), .B2(
        n9912), .ZN(n9907) );
  NAND2_X1 U10962 ( .A1(n9908), .A2(n9907), .ZN(P1_U3249) );
  INV_X1 U10963 ( .A(n9909), .ZN(n9910) );
  AOI21_X1 U10964 ( .B1(n9912), .B2(n9911), .A(n9910), .ZN(n9924) );
  AOI21_X1 U10965 ( .B1(n9915), .B2(n9914), .A(n9913), .ZN(n9922) );
  OAI21_X1 U10966 ( .B1(n9918), .B2(n9917), .A(n9916), .ZN(n9919) );
  AOI22_X1 U10967 ( .A1(n9922), .A2(n9921), .B1(n9920), .B2(n9919), .ZN(n9923)
         );
  OAI211_X1 U10968 ( .C1(n9925), .C2(n10107), .A(n9924), .B(n9923), .ZN(
        P1_U3259) );
  AND2_X1 U10969 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9926), .ZN(P1_U3292) );
  AND2_X1 U10970 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9926), .ZN(P1_U3293) );
  AND2_X1 U10971 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9926), .ZN(P1_U3294) );
  AND2_X1 U10972 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9926), .ZN(P1_U3295) );
  AND2_X1 U10973 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9926), .ZN(P1_U3296) );
  AND2_X1 U10974 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9926), .ZN(P1_U3297) );
  AND2_X1 U10975 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9926), .ZN(P1_U3298) );
  AND2_X1 U10976 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9926), .ZN(P1_U3299) );
  AND2_X1 U10977 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9926), .ZN(P1_U3300) );
  AND2_X1 U10978 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9926), .ZN(P1_U3301) );
  AND2_X1 U10979 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9926), .ZN(P1_U3302) );
  AND2_X1 U10980 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9926), .ZN(P1_U3303) );
  AND2_X1 U10981 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9926), .ZN(P1_U3304) );
  AND2_X1 U10982 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9926), .ZN(P1_U3305) );
  AND2_X1 U10983 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9926), .ZN(P1_U3306) );
  AND2_X1 U10984 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9926), .ZN(P1_U3307) );
  AND2_X1 U10985 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9926), .ZN(P1_U3308) );
  AND2_X1 U10986 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9926), .ZN(P1_U3309) );
  AND2_X1 U10987 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9926), .ZN(P1_U3310) );
  AND2_X1 U10988 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9926), .ZN(P1_U3311) );
  AND2_X1 U10989 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9926), .ZN(P1_U3312) );
  AND2_X1 U10990 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9926), .ZN(P1_U3313) );
  AND2_X1 U10991 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9926), .ZN(P1_U3314) );
  AND2_X1 U10992 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9926), .ZN(P1_U3315) );
  AND2_X1 U10993 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9926), .ZN(P1_U3316) );
  AND2_X1 U10994 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9926), .ZN(P1_U3317) );
  AND2_X1 U10995 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9926), .ZN(P1_U3318) );
  AND2_X1 U10996 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9926), .ZN(P1_U3319) );
  AND2_X1 U10997 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9926), .ZN(P1_U3320) );
  AND2_X1 U10998 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9926), .ZN(P1_U3321) );
  OAI22_X1 U10999 ( .A1(n9928), .A2(n9963), .B1(n9927), .B2(n9961), .ZN(n9930)
         );
  AOI211_X1 U11000 ( .C1(n9960), .C2(n9931), .A(n9930), .B(n9929), .ZN(n9972)
         );
  AOI22_X1 U11001 ( .A1(n9971), .A2(n9972), .B1(n4989), .B2(n9969), .ZN(
        P1_U3463) );
  OR2_X1 U11002 ( .A1(n9933), .A2(n9932), .ZN(n9940) );
  NAND2_X1 U11003 ( .A1(n9935), .A2(n9934), .ZN(n9936) );
  AND2_X1 U11004 ( .A1(n9937), .A2(n9936), .ZN(n9938) );
  AND3_X1 U11005 ( .A1(n9940), .A2(n9939), .A3(n9938), .ZN(n9973) );
  INV_X1 U11006 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9941) );
  AOI22_X1 U11007 ( .A1(n9971), .A2(n9973), .B1(n9941), .B2(n9969), .ZN(
        P1_U3469) );
  OAI22_X1 U11008 ( .A1(n9943), .A2(n9963), .B1(n9942), .B2(n9961), .ZN(n9945)
         );
  AOI211_X1 U11009 ( .C1(n9960), .C2(n9946), .A(n9945), .B(n9944), .ZN(n9974)
         );
  INV_X1 U11010 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9947) );
  AOI22_X1 U11011 ( .A1(n9971), .A2(n9974), .B1(n9947), .B2(n9969), .ZN(
        P1_U3472) );
  OAI21_X1 U11012 ( .B1(n9949), .B2(n9961), .A(n9948), .ZN(n9951) );
  AOI211_X1 U11013 ( .C1(n9967), .C2(n9952), .A(n9951), .B(n9950), .ZN(n9975)
         );
  INV_X1 U11014 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9953) );
  AOI22_X1 U11015 ( .A1(n9971), .A2(n9975), .B1(n9953), .B2(n9969), .ZN(
        P1_U3475) );
  INV_X1 U11016 ( .A(n9954), .ZN(n9959) );
  OAI22_X1 U11017 ( .A1(n9956), .A2(n9963), .B1(n9955), .B2(n9961), .ZN(n9958)
         );
  AOI211_X1 U11018 ( .C1(n9960), .C2(n9959), .A(n9958), .B(n9957), .ZN(n9977)
         );
  AOI22_X1 U11019 ( .A1(n9971), .A2(n9977), .B1(n5124), .B2(n9969), .ZN(
        P1_U3478) );
  OAI22_X1 U11020 ( .A1(n9964), .A2(n9963), .B1(n9962), .B2(n9961), .ZN(n9966)
         );
  AOI211_X1 U11021 ( .C1(n9968), .C2(n9967), .A(n9966), .B(n9965), .ZN(n9979)
         );
  INV_X1 U11022 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9970) );
  AOI22_X1 U11023 ( .A1(n9971), .A2(n9979), .B1(n9970), .B2(n9969), .ZN(
        P1_U3481) );
  AOI22_X1 U11024 ( .A1(n9980), .A2(n9972), .B1(n4988), .B2(n9978), .ZN(
        P1_U3526) );
  AOI22_X1 U11025 ( .A1(n9980), .A2(n9973), .B1(n5047), .B2(n9978), .ZN(
        P1_U3528) );
  AOI22_X1 U11026 ( .A1(n9980), .A2(n9974), .B1(n5070), .B2(n9978), .ZN(
        P1_U3529) );
  AOI22_X1 U11027 ( .A1(n9980), .A2(n9975), .B1(n5096), .B2(n9978), .ZN(
        P1_U3530) );
  INV_X1 U11028 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9976) );
  AOI22_X1 U11029 ( .A1(n9980), .A2(n9977), .B1(n9976), .B2(n9978), .ZN(
        P1_U3531) );
  AOI22_X1 U11030 ( .A1(n9980), .A2(n9979), .B1(n6217), .B2(n9978), .ZN(
        P1_U3532) );
  AOI22_X1 U11031 ( .A1(n9986), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9981), .ZN(n9991) );
  INV_X1 U11032 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9985) );
  OAI21_X1 U11033 ( .B1(n9983), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9982), .ZN(
        n9984) );
  AOI21_X1 U11034 ( .B1(n9986), .B2(n9985), .A(n9984), .ZN(n9989) );
  AOI22_X1 U11035 ( .A1(n9987), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9988) );
  OAI221_X1 U11036 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9991), .C1(n9990), .C2(
        n9989), .A(n9988), .ZN(P2_U3245) );
  INV_X1 U11037 ( .A(n9992), .ZN(n9993) );
  AND2_X1 U11038 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9997), .ZN(P2_U3297) );
  AND2_X1 U11039 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9997), .ZN(P2_U3298) );
  AND2_X1 U11040 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9997), .ZN(P2_U3299) );
  AND2_X1 U11041 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9997), .ZN(P2_U3300) );
  AND2_X1 U11042 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9997), .ZN(P2_U3301) );
  AND2_X1 U11043 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9997), .ZN(P2_U3302) );
  AND2_X1 U11044 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9997), .ZN(P2_U3303) );
  AND2_X1 U11045 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9997), .ZN(P2_U3304) );
  AND2_X1 U11046 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9997), .ZN(P2_U3305) );
  AND2_X1 U11047 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9997), .ZN(P2_U3306) );
  AND2_X1 U11048 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9997), .ZN(P2_U3307) );
  AND2_X1 U11049 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9997), .ZN(P2_U3308) );
  AND2_X1 U11050 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9997), .ZN(P2_U3309) );
  AND2_X1 U11051 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9997), .ZN(P2_U3310) );
  AND2_X1 U11052 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9997), .ZN(P2_U3311) );
  AND2_X1 U11053 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9997), .ZN(P2_U3312) );
  AND2_X1 U11054 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9997), .ZN(P2_U3313) );
  AND2_X1 U11055 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9997), .ZN(P2_U3314) );
  AND2_X1 U11056 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9997), .ZN(P2_U3315) );
  AND2_X1 U11057 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9997), .ZN(P2_U3316) );
  AND2_X1 U11058 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9997), .ZN(P2_U3317) );
  AND2_X1 U11059 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9997), .ZN(P2_U3318) );
  AND2_X1 U11060 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9997), .ZN(P2_U3319) );
  AND2_X1 U11061 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9997), .ZN(P2_U3320) );
  AND2_X1 U11062 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9997), .ZN(P2_U3321) );
  AND2_X1 U11063 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9997), .ZN(P2_U3322) );
  AND2_X1 U11064 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9997), .ZN(P2_U3323) );
  AND2_X1 U11065 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9997), .ZN(P2_U3324) );
  AND2_X1 U11066 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9997), .ZN(P2_U3325) );
  AND2_X1 U11067 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9997), .ZN(P2_U3326) );
  AOI22_X1 U11068 ( .A1(n10000), .A2(n9996), .B1(n9995), .B2(n9997), .ZN(
        P2_U3437) );
  AOI22_X1 U11069 ( .A1(n10000), .A2(n9999), .B1(n9998), .B2(n9997), .ZN(
        P2_U3438) );
  AOI22_X1 U11070 ( .A1(n10003), .A2(n10052), .B1(n10002), .B2(n10001), .ZN(
        n10004) );
  AND2_X1 U11071 ( .A1(n10005), .A2(n10004), .ZN(n10057) );
  INV_X1 U11072 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10006) );
  AOI22_X1 U11073 ( .A1(n10055), .A2(n10057), .B1(n10006), .B2(n10054), .ZN(
        P2_U3451) );
  OAI211_X1 U11074 ( .C1(n10009), .C2(n10038), .A(n10008), .B(n10007), .ZN(
        n10010) );
  AOI21_X1 U11075 ( .B1(n10052), .B2(n10011), .A(n10010), .ZN(n10058) );
  INV_X1 U11076 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10012) );
  AOI22_X1 U11077 ( .A1(n10055), .A2(n10058), .B1(n10012), .B2(n10054), .ZN(
        P2_U3457) );
  OAI21_X1 U11078 ( .B1(n10014), .B2(n10038), .A(n10013), .ZN(n10016) );
  AOI211_X1 U11079 ( .C1(n10052), .C2(n10017), .A(n10016), .B(n10015), .ZN(
        n10060) );
  AOI22_X1 U11080 ( .A1(n10055), .A2(n10060), .B1(n5816), .B2(n10054), .ZN(
        P2_U3463) );
  OAI21_X1 U11081 ( .B1(n10019), .B2(n10038), .A(n10018), .ZN(n10021) );
  AOI211_X1 U11082 ( .C1(n10052), .C2(n10022), .A(n10021), .B(n10020), .ZN(
        n10062) );
  AOI22_X1 U11083 ( .A1(n10055), .A2(n10062), .B1(n5827), .B2(n10054), .ZN(
        P2_U3466) );
  AOI21_X1 U11084 ( .B1(n10045), .B2(n10024), .A(n10023), .ZN(n10025) );
  OAI211_X1 U11085 ( .C1(n10028), .C2(n10027), .A(n10026), .B(n10025), .ZN(
        n10029) );
  INV_X1 U11086 ( .A(n10029), .ZN(n10064) );
  INV_X1 U11087 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10030) );
  AOI22_X1 U11088 ( .A1(n10055), .A2(n10064), .B1(n10030), .B2(n10054), .ZN(
        P2_U3469) );
  INV_X1 U11089 ( .A(n10031), .ZN(n10044) );
  OAI22_X1 U11090 ( .A1(n10033), .A2(n10050), .B1(n10032), .B2(n10038), .ZN(
        n10035) );
  AOI211_X1 U11091 ( .C1(n10044), .C2(n10036), .A(n10035), .B(n10034), .ZN(
        n10065) );
  AOI22_X1 U11092 ( .A1(n10055), .A2(n10065), .B1(n5869), .B2(n10054), .ZN(
        P2_U3475) );
  INV_X1 U11093 ( .A(n10037), .ZN(n10043) );
  OAI22_X1 U11094 ( .A1(n10040), .A2(n10050), .B1(n10039), .B2(n10038), .ZN(
        n10042) );
  AOI211_X1 U11095 ( .C1(n10044), .C2(n10043), .A(n10042), .B(n10041), .ZN(
        n10066) );
  AOI22_X1 U11096 ( .A1(n10055), .A2(n10066), .B1(n5899), .B2(n10054), .ZN(
        P2_U3481) );
  NAND2_X1 U11097 ( .A1(n10046), .A2(n10045), .ZN(n10047) );
  OAI211_X1 U11098 ( .C1(n10050), .C2(n10049), .A(n10048), .B(n10047), .ZN(
        n10051) );
  AOI21_X1 U11099 ( .B1(n10053), .B2(n10052), .A(n10051), .ZN(n10068) );
  AOI22_X1 U11100 ( .A1(n10055), .A2(n10068), .B1(n5928), .B2(n10054), .ZN(
        P2_U3487) );
  AOI22_X1 U11101 ( .A1(n10069), .A2(n10057), .B1(n10056), .B2(n10067), .ZN(
        P2_U3520) );
  AOI22_X1 U11102 ( .A1(n10069), .A2(n10058), .B1(n6607), .B2(n10067), .ZN(
        P2_U3522) );
  INV_X1 U11103 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10059) );
  AOI22_X1 U11104 ( .A1(n10069), .A2(n10060), .B1(n10059), .B2(n10067), .ZN(
        P2_U3524) );
  INV_X1 U11105 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10061) );
  AOI22_X1 U11106 ( .A1(n10069), .A2(n10062), .B1(n10061), .B2(n10067), .ZN(
        P2_U3525) );
  INV_X1 U11107 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10063) );
  AOI22_X1 U11108 ( .A1(n10069), .A2(n10064), .B1(n10063), .B2(n10067), .ZN(
        P2_U3526) );
  AOI22_X1 U11109 ( .A1(n10069), .A2(n10065), .B1(n6733), .B2(n10067), .ZN(
        P2_U3528) );
  AOI22_X1 U11110 ( .A1(n10069), .A2(n10066), .B1(n6735), .B2(n10067), .ZN(
        P2_U3530) );
  AOI22_X1 U11111 ( .A1(n10069), .A2(n10068), .B1(n6827), .B2(n10067), .ZN(
        P2_U3532) );
  INV_X1 U11112 ( .A(n10070), .ZN(n10071) );
  NAND2_X1 U11113 ( .A1(n10072), .A2(n10071), .ZN(n10073) );
  XOR2_X1 U11114 ( .A(n10074), .B(n10073), .Z(ADD_1071_U5) );
  XOR2_X1 U11115 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11116 ( .B1(n10077), .B2(n10076), .A(n10075), .ZN(ADD_1071_U56) );
  OAI21_X1 U11117 ( .B1(n10080), .B2(n10079), .A(n10078), .ZN(ADD_1071_U57) );
  OAI21_X1 U11118 ( .B1(n10083), .B2(n10082), .A(n10081), .ZN(ADD_1071_U58) );
  OAI21_X1 U11119 ( .B1(n10086), .B2(n10085), .A(n10084), .ZN(ADD_1071_U59) );
  OAI21_X1 U11120 ( .B1(n10089), .B2(n10088), .A(n10087), .ZN(ADD_1071_U60) );
  OAI21_X1 U11121 ( .B1(n10092), .B2(n10091), .A(n10090), .ZN(ADD_1071_U61) );
  AOI21_X1 U11122 ( .B1(n10095), .B2(n10094), .A(n10093), .ZN(ADD_1071_U62) );
  AOI21_X1 U11123 ( .B1(n10098), .B2(n10097), .A(n10096), .ZN(ADD_1071_U63) );
  AOI21_X1 U11124 ( .B1(n10101), .B2(n10100), .A(n10099), .ZN(ADD_1071_U47) );
  XOR2_X1 U11125 ( .A(n10103), .B(n10102), .Z(ADD_1071_U54) );
  XOR2_X1 U11126 ( .A(n10104), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  OAI21_X1 U11127 ( .B1(n10107), .B2(n10106), .A(n10105), .ZN(n10108) );
  XNOR2_X1 U11128 ( .A(n10108), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11129 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10109), .Z(ADD_1071_U49) );
  XOR2_X1 U11130 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10110), .Z(ADD_1071_U50) );
  AOI21_X1 U11131 ( .B1(n10112), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n10111), .ZN(
        n10113) );
  XOR2_X1 U11132 ( .A(n10113), .B(P1_ADDR_REG_5__SCAN_IN), .Z(ADD_1071_U51) );
  XOR2_X1 U11133 ( .A(n10115), .B(n10114), .Z(ADD_1071_U53) );
  XNOR2_X1 U11134 ( .A(n10117), .B(n10116), .ZN(ADD_1071_U52) );
  CLKBUF_X3 U4818 ( .A(n4987), .Z(n8830) );
  CLKBUF_X3 U4852 ( .A(n4949), .Z(n8837) );
  CLKBUF_X1 U4887 ( .A(n5676), .Z(n4312) );
endmodule

