

module b21_C_SARLock_k_128_10 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4451, n4452,
         n4453, n4454, n4455, n4456, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341;

  INV_X2 U4948 ( .A(n9738), .ZN(n10031) );
  OR2_X1 U4949 ( .A1(n9596), .A2(n9584), .ZN(n9580) );
  OAI21_X1 U4950 ( .B1(n7724), .B2(n4634), .A(n4631), .ZN(n6042) );
  INV_X1 U4952 ( .A(n6228), .ZN(n8202) );
  CLKBUF_X2 U4953 ( .A(n5130), .Z(n6888) );
  BUF_X1 U4954 ( .A(n5101), .Z(n7001) );
  INV_X1 U4955 ( .A(n8787), .ZN(n8771) );
  NAND2_X1 U4956 ( .A1(n4709), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4708) );
  INV_X1 U4957 ( .A(n5042), .ZN(n5044) );
  INV_X1 U4958 ( .A(n5844), .ZN(n5802) );
  INV_X1 U4959 ( .A(n5802), .ZN(n6270) );
  OR2_X1 U4960 ( .A1(n10016), .A2(n7699), .ZN(n7790) );
  INV_X1 U4962 ( .A(n5075), .ZN(n6838) );
  AND2_X1 U4963 ( .A1(n4899), .A2(n4490), .ZN(n4905) );
  INV_X1 U4964 ( .A(n5130), .ZN(n8599) );
  AND3_X1 U4966 ( .A1(n5217), .A2(n5216), .A3(n5215), .ZN(n10239) );
  NAND2_X1 U4967 ( .A1(n5073), .A2(n5074), .ZN(n5075) );
  OAI21_X1 U4968 ( .B1(n6365), .B2(n5700), .A(n5699), .ZN(n6360) );
  NAND2_X1 U4969 ( .A1(n5396), .A2(n5395), .ZN(n9350) );
  INV_X1 U4970 ( .A(n9075), .ZN(n9064) );
  NAND2_X1 U4971 ( .A1(n9222), .A2(n9007), .ZN(n9205) );
  INV_X1 U4972 ( .A(n5884), .ZN(n6460) );
  NAND3_X1 U4973 ( .A1(n4466), .A2(n5777), .A3(n5776), .ZN(n5785) );
  NAND2_X1 U4974 ( .A1(n5766), .A2(n5778), .ZN(n8289) );
  NAND2_X1 U4975 ( .A1(n7579), .A2(n5246), .ZN(n7666) );
  INV_X1 U4976 ( .A(n5867), .ZN(n4442) );
  NAND2_X1 U4977 ( .A1(n4546), .A2(n9833), .ZN(n5867) );
  NAND2_X2 U4978 ( .A1(n7272), .A2(n8658), .ZN(n7028) );
  NOR3_X2 U4979 ( .A1(n9719), .A2(n4689), .A3(n9781), .ZN(n4688) );
  NAND2_X2 U4980 ( .A1(n7639), .A2(n8676), .ZN(n7641) );
  NAND2_X2 U4981 ( .A1(n7523), .A2(n4724), .ZN(n7639) );
  AOI21_X2 U4982 ( .B1(n8416), .B2(n8415), .A(n8414), .ZN(n8421) );
  NAND2_X2 U4983 ( .A1(n9082), .A2(n9027), .ZN(n9030) );
  NAND2_X2 U4984 ( .A1(n9026), .A2(n9025), .ZN(n9082) );
  AND4_X2 U4985 ( .A1(n6952), .A2(n6951), .A3(n6950), .A4(n6949), .ZN(n7026)
         );
  OAI21_X2 U4986 ( .B1(n4511), .B2(n4540), .A(n5406), .ZN(n8183) );
  NAND3_X2 U4987 ( .A1(n7641), .A2(n7640), .A3(n7642), .ZN(n7674) );
  XNOR2_X2 U4988 ( .A(n5770), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5775) );
  OR2_X2 U4989 ( .A1(n9825), .A2(n9826), .ZN(n5770) );
  OR2_X2 U4990 ( .A1(n5043), .A2(n5044), .ZN(n5130) );
  XNOR2_X2 U4991 ( .A(n4600), .B(n4599), .ZN(n9833) );
  NAND2_X1 U4992 ( .A1(n7422), .A2(n5079), .ZN(n4443) );
  BUF_X8 U4994 ( .A(n6838), .Z(n4445) );
  OR2_X1 U4995 ( .A1(n8799), .A2(n10218), .ZN(n4446) );
  INV_X2 U4996 ( .A(n8611), .ZN(n6340) );
  CLKBUF_X1 U4997 ( .A(n5130), .Z(n4447) );
  NAND2_X1 U4998 ( .A1(n9162), .A2(n4472), .ZN(n4720) );
  NAND2_X1 U4999 ( .A1(n5530), .A2(n8832), .ZN(n8835) );
  INV_X1 U5000 ( .A(n4563), .ZN(n9223) );
  CLKBUF_X2 U5001 ( .A(n5842), .Z(n6226) );
  NAND2_X2 U5002 ( .A1(n8661), .A2(n8659), .ZN(n8613) );
  INV_X1 U5003 ( .A(n8912), .ZN(n4556) );
  INV_X1 U5004 ( .A(n8827), .ZN(n8911) );
  INV_X1 U5005 ( .A(n8822), .ZN(n7275) );
  OR2_X1 U5006 ( .A1(n5130), .A2(n7625), .ZN(n6949) );
  CLKBUF_X1 U5008 ( .A(n5075), .Z(n8228) );
  NOR2_X1 U5009 ( .A1(n6271), .A2(n6273), .ZN(n6325) );
  NAND2_X1 U5010 ( .A1(n6275), .A2(n6274), .ZN(n9384) );
  OAI21_X1 U5011 ( .B1(n4917), .B2(n4916), .A(n6364), .ZN(n5696) );
  OR2_X1 U5012 ( .A1(n6201), .A2(n6200), .ZN(n5023) );
  AOI21_X1 U5013 ( .B1(n8843), .B2(n5595), .A(n4920), .ZN(n4919) );
  NAND2_X1 U5014 ( .A1(n8835), .A2(n5534), .ZN(n5557) );
  NAND2_X1 U5015 ( .A1(n9014), .A2(n5016), .ZN(n9179) );
  NAND2_X1 U5016 ( .A1(n8770), .A2(n8597), .ZN(n9057) );
  AND2_X1 U5017 ( .A1(n8470), .A2(n8471), .ZN(n9567) );
  AND2_X1 U5018 ( .A1(n9133), .A2(n9132), .ZN(n9135) );
  NAND2_X1 U5019 ( .A1(n9223), .A2(n9226), .ZN(n9222) );
  OAI211_X1 U5020 ( .C1(n4581), .C2(n9730), .A(n4580), .B(n8296), .ZN(n9686)
         );
  INV_X1 U5021 ( .A(n4560), .ZN(n4559) );
  AOI21_X1 U5022 ( .B1(n4560), .B2(n9262), .A(n4783), .ZN(n4558) );
  OAI21_X1 U5023 ( .B1(n5561), .B2(n5560), .A(n5559), .ZN(n5570) );
  OAI21_X1 U5024 ( .B1(n5537), .B2(n5536), .A(n5540), .ZN(n5561) );
  NAND2_X1 U5025 ( .A1(n6131), .A2(n6130), .ZN(n9803) );
  NAND2_X1 U5026 ( .A1(n6111), .A2(n6110), .ZN(n9740) );
  NAND2_X1 U5027 ( .A1(n5438), .A2(n5437), .ZN(n9247) );
  AND2_X1 U5028 ( .A1(n4573), .A2(n4571), .ZN(n7762) );
  NAND2_X1 U5029 ( .A1(n6029), .A2(n6028), .ZN(n7915) );
  NAND2_X1 U5030 ( .A1(n7526), .A2(n8619), .ZN(n7646) );
  AOI21_X1 U5031 ( .B1(n5386), .B2(n4812), .A(n4809), .ZN(n4808) );
  AOI21_X1 U5032 ( .B1(n7563), .B2(n8620), .A(n8670), .ZN(n7526) );
  NAND2_X1 U5033 ( .A1(n6010), .A2(n6009), .ZN(n8028) );
  NAND2_X1 U5034 ( .A1(n5318), .A2(n5317), .ZN(n5337) );
  INV_X2 U5035 ( .A(n10292), .ZN(n4449) );
  OR2_X1 U5036 ( .A1(n5314), .A2(n5313), .ZN(n5318) );
  CLKBUF_X1 U5037 ( .A(n6437), .Z(n10128) );
  AND2_X1 U5038 ( .A1(n6437), .A2(n5784), .ZN(n5842) );
  NAND2_X1 U5040 ( .A1(n4810), .A2(n5432), .ZN(n4809) );
  AND2_X1 U5041 ( .A1(n5797), .A2(n7253), .ZN(n5844) );
  BUF_X2 U5042 ( .A(n5702), .Z(n4462) );
  NAND2_X1 U5043 ( .A1(n4812), .A2(n4814), .ZN(n4810) );
  AND4_X1 U5044 ( .A1(n5841), .A2(n5840), .A3(n5839), .A4(n5838), .ZN(n7387)
         );
  AND3_X2 U5045 ( .A1(n5123), .A2(n5122), .A3(n5121), .ZN(n8826) );
  AND4_X1 U5046 ( .A1(n5134), .A2(n5133), .A3(n5132), .A4(n5131), .ZN(n8827)
         );
  AND2_X2 U5047 ( .A1(n6928), .A2(n6469), .ZN(n10089) );
  NAND2_X1 U5048 ( .A1(n5144), .A2(n5143), .ZN(n5163) );
  INV_X1 U5049 ( .A(n6438), .ZN(n8556) );
  OR2_X1 U5050 ( .A1(n8289), .A2(n6468), .ZN(n5784) );
  INV_X2 U5051 ( .A(n4456), .ZN(n4459) );
  INV_X2 U5052 ( .A(n4456), .ZN(n4458) );
  NAND2_X1 U5053 ( .A1(n5056), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5061) );
  INV_X2 U5054 ( .A(n5110), .ZN(n8233) );
  INV_X2 U5055 ( .A(n6308), .ZN(n5807) );
  NAND2_X1 U5056 ( .A1(n8158), .A2(n5761), .ZN(n5797) );
  NAND2_X1 U5057 ( .A1(n5101), .A2(n8228), .ZN(n5110) );
  INV_X1 U5058 ( .A(n5101), .ZN(n4711) );
  NAND2_X1 U5059 ( .A1(n5054), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5455) );
  OR2_X1 U5060 ( .A1(n9372), .A2(n9374), .ZN(n5036) );
  XNOR2_X1 U5061 ( .A(n4601), .B(n5070), .ZN(n8809) );
  XNOR2_X1 U5062 ( .A(n5063), .B(n4940), .ZN(n8635) );
  OAI21_X1 U5063 ( .B1(n4624), .B2(n5743), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5744) );
  NAND2_X1 U5064 ( .A1(n4602), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4601) );
  INV_X2 U5065 ( .A(n7985), .ZN(n4451) );
  CLKBUF_X1 U5066 ( .A(n5857), .Z(n5892) );
  OR2_X1 U5067 ( .A1(n5034), .A2(n4512), .ZN(n4478) );
  AND2_X1 U5068 ( .A1(n5005), .A2(n6293), .ZN(n4468) );
  OAI21_X2 U5069 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        n5072), .ZN(n5074) );
  AND2_X1 U5070 ( .A1(n4960), .A2(n5025), .ZN(n4898) );
  AND2_X1 U5071 ( .A1(n5739), .A2(n5006), .ZN(n5005) );
  AND4_X1 U5072 ( .A1(n4714), .A2(n4713), .A3(n5273), .A4(n5213), .ZN(n4712)
         );
  OR2_X1 U5073 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(n5033), .ZN(n5034) );
  AND2_X1 U5074 ( .A1(n5735), .A2(n5734), .ZN(n5854) );
  AND2_X1 U5075 ( .A1(n5091), .A2(n4715), .ZN(n5026) );
  NOR3_X1 U5076 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .A3(
        P1_IR_REG_22__SCAN_IN), .ZN(n5739) );
  INV_X1 U5077 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5213) );
  INV_X1 U5078 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5945) );
  NOR2_X1 U5079 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5734) );
  NOR2_X1 U5080 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5735) );
  NOR2_X1 U5081 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5730) );
  INV_X1 U5082 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5035) );
  INV_X1 U5083 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5055) );
  INV_X1 U5084 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5048) );
  INV_X1 U5085 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5391) );
  INV_X1 U5086 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5059) );
  NOR2_X1 U5087 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4714) );
  OR2_X1 U5088 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5033) );
  INV_X1 U5089 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5057) );
  NOR2_X1 U5090 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n4713) );
  INV_X1 U5091 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5273) );
  INV_X1 U5092 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5362) );
  OAI211_X2 U5093 ( .C1(n5110), .C2(n6844), .A(n4708), .B(n4710), .ZN(n7037)
         );
  NAND2_X1 U5094 ( .A1(n5775), .A2(n9833), .ZN(n5872) );
  INV_X1 U5095 ( .A(n8256), .ZN(n10049) );
  NAND3_X1 U5096 ( .A1(n5812), .A2(n5811), .A3(n4497), .ZN(n6375) );
  NAND2_X2 U5097 ( .A1(n7619), .A2(n7025), .ZN(n7272) );
  AOI211_X1 U5098 ( .C1(n7630), .C2(n7629), .A(n8868), .B(n7575), .ZN(n7635)
         );
  OAI21_X2 U5099 ( .B1(n7575), .B2(n5223), .A(n7576), .ZN(n7579) );
  NOR2_X2 U5100 ( .A1(n7630), .A2(n7629), .ZN(n7575) );
  OAI21_X2 U5101 ( .B1(n4780), .B2(n4559), .A(n4558), .ZN(n4563) );
  NAND2_X2 U5102 ( .A1(n4726), .A2(n4489), .ZN(n4780) );
  INV_X1 U5103 ( .A(n5844), .ZN(n6265) );
  INV_X1 U5104 ( .A(n5101), .ZN(n4452) );
  NOR2_X2 U5105 ( .A1(n5661), .A2(n4478), .ZN(n9372) );
  NAND2_X1 U5106 ( .A1(n5045), .A2(n5044), .ZN(n4453) );
  NAND2_X1 U5107 ( .A1(n5045), .A2(n5044), .ZN(n4454) );
  NAND2_X1 U5108 ( .A1(n7026), .A2(n7037), .ZN(n8658) );
  AND2_X1 U5109 ( .A1(n5042), .A2(n5043), .ZN(n5128) );
  CLKBUF_X1 U5110 ( .A(n5479), .Z(n4455) );
  XNOR2_X1 U5111 ( .A(n5061), .B(P2_IR_REG_19__SCAN_IN), .ZN(n5479) );
  INV_X1 U5114 ( .A(n5522), .ZN(n4460) );
  INV_X2 U5115 ( .A(n5522), .ZN(n4461) );
  NAND2_X4 U5116 ( .A1(n8807), .A2(n5044), .ZN(n5522) );
  NOR2_X1 U5117 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5032) );
  OR2_X1 U5118 ( .A1(n9584), .A2(n9589), .ZN(n8470) );
  AOI21_X1 U5119 ( .B1(n5338), .B2(n5339), .A(n4833), .ZN(n4832) );
  NAND2_X1 U5120 ( .A1(n4789), .A2(n4484), .ZN(n5255) );
  OR2_X1 U5121 ( .A1(n9325), .A2(n9175), .ZN(n8745) );
  NAND2_X1 U5122 ( .A1(n9593), .A2(n6408), .ZN(n9568) );
  NAND2_X1 U5123 ( .A1(n6064), .A2(n4445), .ZN(n5834) );
  AOI21_X1 U5124 ( .B1(n8358), .B2(n4545), .A(n6384), .ZN(n4544) );
  NAND2_X1 U5125 ( .A1(n8357), .A2(n8482), .ZN(n4543) );
  MUX2_X1 U5126 ( .A(n8463), .B(n8462), .S(n4545), .Z(n8465) );
  OR2_X1 U5127 ( .A1(n9295), .A2(n9072), .ZN(n8761) );
  NOR2_X1 U5128 ( .A1(n5496), .A2(n4806), .ZN(n4805) );
  INV_X1 U5129 ( .A(n5474), .ZN(n4806) );
  INV_X1 U5130 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5319) );
  AND2_X1 U5131 ( .A1(n8675), .A2(n7645), .ZN(n4961) );
  NOR2_X1 U5132 ( .A1(n9316), .A2(n8900), .ZN(n9020) );
  INV_X1 U5133 ( .A(n9019), .ZN(n4722) );
  INV_X1 U5134 ( .A(n8289), .ZN(n8500) );
  OR2_X1 U5135 ( .A1(n9756), .A2(n9575), .ZN(n8467) );
  NAND2_X1 U5136 ( .A1(n4504), .A2(n4667), .ZN(n4663) );
  OR2_X1 U5137 ( .A1(n8060), .A2(n9427), .ZN(n8411) );
  XNOR2_X1 U5138 ( .A(n6375), .B(n10092), .ZN(n8256) );
  NAND2_X1 U5139 ( .A1(n6337), .A2(n6336), .ZN(n6423) );
  AND2_X1 U5140 ( .A1(n5517), .A2(n5500), .ZN(n5515) );
  NOR2_X1 U5141 ( .A1(n4794), .A2(n4791), .ZN(n4790) );
  INV_X1 U5142 ( .A(n5234), .ZN(n4794) );
  INV_X1 U5143 ( .A(n5209), .ZN(n4791) );
  INV_X1 U5144 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5072) );
  NAND2_X1 U5145 ( .A1(n4919), .A2(n4918), .ZN(n4915) );
  OR2_X1 U5146 ( .A1(n5224), .A2(n8926), .ZN(n5282) );
  NOR2_X1 U5147 ( .A1(n6774), .A2(n4926), .ZN(n4925) );
  INV_X1 U5148 ( .A(n5494), .ZN(n4926) );
  NAND2_X1 U5149 ( .A1(n4912), .A2(n4910), .ZN(n4916) );
  NAND2_X1 U5150 ( .A1(n4908), .A2(n5616), .ZN(n4917) );
  OR2_X1 U5151 ( .A1(n6326), .A2(n4911), .ZN(n4910) );
  NAND2_X1 U5152 ( .A1(n4948), .A2(n4952), .ZN(n4946) );
  AND2_X1 U5153 ( .A1(n4949), .A2(n4950), .ZN(n4948) );
  NOR2_X1 U5154 ( .A1(n9119), .A2(n4782), .ZN(n4781) );
  INV_X1 U5155 ( .A(n9023), .ZN(n4782) );
  NAND2_X1 U5156 ( .A1(n4956), .A2(n4500), .ZN(n9170) );
  INV_X1 U5157 ( .A(n9173), .ZN(n4959) );
  NAND2_X1 U5158 ( .A1(n9179), .A2(n9186), .ZN(n4557) );
  OR2_X1 U5159 ( .A1(n9254), .A2(n9345), .ZN(n9235) );
  NAND2_X1 U5160 ( .A1(n8006), .A2(n4496), .ZN(n8007) );
  INV_X1 U5161 ( .A(n7443), .ZN(n4555) );
  AND4_X2 U5162 ( .A1(n5090), .A2(n5089), .A3(n5088), .A4(n5087), .ZN(n8822)
         );
  OR2_X1 U5163 ( .A1(n4447), .A2(n7429), .ZN(n5087) );
  AND2_X1 U5164 ( .A1(n7022), .A2(n7021), .ZN(n7127) );
  AND2_X1 U5165 ( .A1(n4471), .A2(n4728), .ZN(n4727) );
  NOR2_X1 U5166 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n4728) );
  XNOR2_X1 U5167 ( .A(n5981), .B(n5982), .ZN(n7707) );
  OR2_X1 U5168 ( .A1(n9876), .A2(n8245), .ZN(n8544) );
  CLKBUF_X1 U5169 ( .A(n6308), .Z(n6416) );
  NOR2_X1 U5170 ( .A1(n9545), .A2(n4834), .ZN(n9546) );
  AND2_X1 U5171 ( .A1(n9548), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4834) );
  NAND2_X1 U5172 ( .A1(n9730), .A2(n8419), .ZN(n4767) );
  AOI21_X1 U5173 ( .B1(n4469), .B2(n4885), .A(n4506), .ZN(n4880) );
  INV_X1 U5174 ( .A(n4886), .ZN(n4885) );
  INV_X1 U5175 ( .A(n5878), .ZN(n6144) );
  AOI21_X1 U5176 ( .B1(n7380), .B2(n8361), .A(n6386), .ZN(n7479) );
  NAND2_X1 U5177 ( .A1(n7390), .A2(n8255), .ZN(n4857) );
  AND4_X1 U5178 ( .A1(n5853), .A2(n5852), .A3(n5851), .A4(n5850), .ZN(n7364)
         );
  NAND2_X1 U5179 ( .A1(n6430), .A2(n6429), .ZN(n8483) );
  INV_X1 U5180 ( .A(n4878), .ZN(n4867) );
  OAI22_X1 U5181 ( .A1(n9589), .A2(n6463), .B1(n6465), .B2(n6464), .ZN(n4878)
         );
  NAND2_X1 U5182 ( .A1(n4465), .A2(n10050), .ZN(n4866) );
  NAND2_X1 U5183 ( .A1(n4594), .A2(n4592), .ZN(n4598) );
  NAND2_X1 U5184 ( .A1(n9568), .A2(n4501), .ZN(n4870) );
  NAND2_X1 U5185 ( .A1(n4879), .A2(n4875), .ZN(n4874) );
  NAND2_X1 U5186 ( .A1(n9567), .A2(n4876), .ZN(n4875) );
  AND2_X1 U5187 ( .A1(n6931), .A2(n8546), .ZN(n10149) );
  INV_X1 U5188 ( .A(n4811), .ZN(n5431) );
  AOI21_X1 U5189 ( .B1(n5386), .B2(n4816), .A(n4814), .ZN(n4811) );
  OAI21_X1 U5190 ( .B1(n4902), .B2(n7976), .A(n8141), .ZN(n4540) );
  NAND2_X1 U5191 ( .A1(n4865), .A2(n4877), .ZN(n4871) );
  NOR2_X1 U5192 ( .A1(n4879), .A2(n9567), .ZN(n4877) );
  INV_X1 U5193 ( .A(n9568), .ZN(n4865) );
  AOI21_X1 U5194 ( .B1(n8395), .B2(n8394), .A(n8393), .ZN(n8400) );
  NOR2_X1 U5195 ( .A1(n8787), .A2(n4740), .ZN(n4739) );
  AOI21_X1 U5196 ( .B1(n8697), .B2(n8696), .A(n8695), .ZN(n4743) );
  AND2_X1 U5197 ( .A1(n8702), .A2(n8787), .ZN(n4742) );
  MUX2_X1 U5198 ( .A(n8352), .B(n8351), .S(n8482), .Z(n8454) );
  AOI211_X1 U5199 ( .C1(n8734), .C2(n8745), .A(n8747), .B(n8733), .ZN(n4748)
         );
  OR2_X1 U5200 ( .A1(n8735), .A2(n8771), .ZN(n4745) );
  NAND2_X1 U5201 ( .A1(n8735), .A2(n4747), .ZN(n4746) );
  NOR2_X1 U5202 ( .A1(n8743), .A2(n8787), .ZN(n4747) );
  AND2_X1 U5203 ( .A1(n8458), .A2(n8444), .ZN(n8529) );
  NAND2_X1 U5204 ( .A1(n4863), .A2(n6390), .ZN(n4862) );
  INV_X1 U5205 ( .A(n6389), .ZN(n4863) );
  INV_X1 U5206 ( .A(SI_10_), .ZN(n6668) );
  OR2_X1 U5207 ( .A1(n8483), .A2(n9574), .ZN(n8292) );
  NAND2_X1 U5208 ( .A1(n5340), .A2(n6594), .ZN(n5360) );
  NOR2_X1 U5209 ( .A1(n4820), .A2(n4824), .ZN(n4819) );
  OAI21_X1 U5210 ( .B1(n5021), .B2(n4824), .A(n5020), .ZN(n4823) );
  NAND2_X1 U5211 ( .A1(n5269), .A2(n6668), .ZN(n5294) );
  INV_X1 U5212 ( .A(n5252), .ZN(n4653) );
  NOR2_X1 U5213 ( .A1(n5906), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5943) );
  AND4_X1 U5214 ( .A1(n4518), .A2(n8783), .A3(n4675), .A4(n4486), .ZN(n8633)
         );
  OR2_X1 U5215 ( .A1(n9047), .A2(n8899), .ZN(n8779) );
  NOR2_X1 U5216 ( .A1(n9057), .A2(n4680), .ZN(n4679) );
  AND2_X1 U5217 ( .A1(n9075), .A2(n4681), .ZN(n4680) );
  NAND2_X1 U5218 ( .A1(n4955), .A2(n4951), .ZN(n4950) );
  INV_X1 U5219 ( .A(n9097), .ZN(n4951) );
  OR2_X1 U5220 ( .A1(n9304), .A2(n9136), .ZN(n9024) );
  NOR2_X1 U5221 ( .A1(n9316), .A2(n9311), .ZN(n4608) );
  AND2_X1 U5222 ( .A1(n8698), .A2(n4567), .ZN(n4566) );
  NAND2_X1 U5223 ( .A1(n8700), .A2(n8686), .ZN(n4567) );
  NOR2_X1 U5224 ( .A1(n7919), .A2(n7849), .ZN(n4615) );
  NAND2_X1 U5225 ( .A1(n7646), .A2(n4961), .ZN(n7676) );
  NOR2_X1 U5226 ( .A1(n4607), .A2(n9304), .ZN(n4606) );
  INV_X1 U5227 ( .A(n4608), .ZN(n4607) );
  NAND2_X1 U5228 ( .A1(n7028), .A2(n7027), .ZN(n7270) );
  AOI21_X1 U5229 ( .B1(n10199), .B2(n10214), .A(n10215), .ZN(n7420) );
  INV_X1 U5230 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4960) );
  XNOR2_X1 U5231 ( .A(n5979), .B(n8200), .ZN(n5981) );
  NAND2_X1 U5232 ( .A1(n7699), .A2(n6256), .ZN(n5978) );
  OAI21_X1 U5233 ( .B1(n9443), .B2(n4510), .A(n4476), .ZN(n6201) );
  NOR2_X1 U5234 ( .A1(n6060), .A2(n8134), .ZN(n4981) );
  INV_X1 U5235 ( .A(n7907), .ZN(n4980) );
  INV_X1 U5236 ( .A(n4635), .ZN(n4634) );
  AOI21_X1 U5237 ( .B1(n4633), .B2(n4635), .A(n4632), .ZN(n4631) );
  INV_X1 U5238 ( .A(n4636), .ZN(n4633) );
  INV_X1 U5239 ( .A(n9833), .ZN(n5774) );
  NOR2_X1 U5240 ( .A1(n9761), .A2(n4701), .ZN(n4700) );
  OR2_X1 U5241 ( .A1(n9768), .A2(n9772), .ZN(n4701) );
  INV_X1 U5242 ( .A(n4663), .ZN(n4659) );
  OR2_X1 U5243 ( .A1(n9798), .A2(n9708), .ZN(n8427) );
  NAND2_X1 U5244 ( .A1(n9913), .A2(n4707), .ZN(n4706) );
  AND2_X1 U5245 ( .A1(n4862), .A2(n4864), .ZN(n4859) );
  INV_X1 U5246 ( .A(n6390), .ZN(n4864) );
  NAND2_X1 U5247 ( .A1(n4770), .A2(n8385), .ZN(n7785) );
  NOR2_X1 U5248 ( .A1(n6448), .A2(n8366), .ZN(n4768) );
  OR2_X1 U5249 ( .A1(n7699), .A2(n7787), .ZN(n8385) );
  NOR2_X1 U5250 ( .A1(n8512), .A2(n4759), .ZN(n4758) );
  INV_X1 U5251 ( .A(n8310), .ZN(n4587) );
  NAND2_X1 U5252 ( .A1(n7367), .A2(n9496), .ZN(n8354) );
  INV_X1 U5253 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U5254 ( .A1(n6427), .A2(n6426), .ZN(n8219) );
  NAND2_X1 U5255 ( .A1(n6423), .A2(n6422), .ZN(n6427) );
  NAND2_X1 U5256 ( .A1(n5640), .A2(n5639), .ZN(n6335) );
  NAND2_X1 U5257 ( .A1(n5572), .A2(n5571), .ZN(n5601) );
  NAND2_X1 U5258 ( .A1(n5570), .A2(n5569), .ZN(n5572) );
  AOI21_X1 U5259 ( .B1(n4802), .B2(n4804), .A(n4801), .ZN(n4800) );
  AOI21_X1 U5260 ( .B1(n5470), .B2(n4805), .A(n4803), .ZN(n4802) );
  INV_X1 U5261 ( .A(n5495), .ZN(n4803) );
  INV_X1 U5262 ( .A(n4805), .ZN(n4804) );
  NAND2_X1 U5263 ( .A1(n5321), .A2(n5320), .ZN(n5339) );
  INV_X1 U5264 ( .A(SI_9_), .ZN(n5256) );
  OAI21_X1 U5265 ( .B1(n4445), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n4541), .ZN(
        n5164) );
  NAND2_X1 U5266 ( .A1(n4444), .A2(n6852), .ZN(n4541) );
  AOI21_X1 U5267 ( .B1(n4933), .B2(n4932), .A(n4931), .ZN(n4930) );
  INV_X1 U5268 ( .A(n7747), .ZN(n4931) );
  INV_X1 U5269 ( .A(n4936), .ZN(n4932) );
  OR2_X1 U5270 ( .A1(n5282), .A2(n5281), .ZN(n5302) );
  AND2_X1 U5271 ( .A1(n5447), .A2(n5428), .ZN(n4939) );
  AND2_X1 U5272 ( .A1(n5697), .A2(n5636), .ZN(n6364) );
  INV_X1 U5273 ( .A(n6326), .ZN(n4914) );
  NAND2_X1 U5274 ( .A1(n5376), .A2(n5404), .ZN(n4904) );
  AND3_X1 U5275 ( .A1(n5614), .A2(n5613), .A3(n5612), .ZN(n8851) );
  AOI21_X1 U5276 ( .B1(n9030), .B2(n4553), .A(n4552), .ZN(n4551) );
  OAI21_X1 U5277 ( .B1(n4554), .B2(n9075), .A(n9057), .ZN(n4552) );
  OR2_X1 U5278 ( .A1(n9074), .A2(n4678), .ZN(n4676) );
  INV_X1 U5279 ( .A(n4679), .ZN(n4678) );
  AOI21_X1 U5280 ( .B1(n4679), .B2(n8772), .A(n8773), .ZN(n4677) );
  AND2_X1 U5281 ( .A1(n9045), .A2(n5710), .ZN(n9055) );
  INV_X1 U5282 ( .A(n4619), .ZN(n4617) );
  OR2_X1 U5283 ( .A1(n9301), .A2(n8851), .ZN(n9085) );
  NAND2_X1 U5284 ( .A1(n5575), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5610) );
  AND4_X1 U5285 ( .A1(n5509), .A2(n5508), .A3(n5507), .A4(n5506), .ZN(n9175)
         );
  NAND2_X1 U5286 ( .A1(n8592), .A2(n4957), .ZN(n4956) );
  NOR2_X1 U5287 ( .A1(n9186), .A2(n4958), .ZN(n4957) );
  INV_X1 U5288 ( .A(n8740), .ZN(n4958) );
  OR2_X1 U5289 ( .A1(n9013), .A2(n9012), .ZN(n5016) );
  OR2_X1 U5290 ( .A1(n9332), .A2(n9210), .ZN(n9011) );
  NAND2_X1 U5291 ( .A1(n5482), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5503) );
  INV_X1 U5292 ( .A(n5483), .ZN(n5482) );
  AND2_X1 U5293 ( .A1(n8737), .A2(n8740), .ZN(n9197) );
  NOR2_X1 U5294 ( .A1(n9235), .A2(n4611), .ZN(n9216) );
  INV_X1 U5295 ( .A(n4613), .ZN(n4611) );
  NOR2_X1 U5296 ( .A1(n8718), .A2(n4561), .ZN(n4560) );
  INV_X1 U5297 ( .A(n8168), .ZN(n4561) );
  OR2_X1 U5298 ( .A1(n9350), .A2(n8901), .ZN(n8168) );
  AND2_X1 U5299 ( .A1(n8720), .A2(n9224), .ZN(n8718) );
  NOR2_X1 U5300 ( .A1(n8172), .A2(n8711), .ZN(n9253) );
  NAND2_X1 U5301 ( .A1(n4963), .A2(n4962), .ZN(n8162) );
  AND2_X1 U5302 ( .A1(n8010), .A2(n8009), .ZN(n4962) );
  NAND2_X1 U5303 ( .A1(n7961), .A2(n7960), .ZN(n8006) );
  AND4_X1 U5304 ( .A1(n5308), .A2(n5307), .A3(n5306), .A4(n5305), .ZN(n7927)
         );
  NAND2_X1 U5305 ( .A1(n7674), .A2(n4730), .ZN(n4734) );
  NOR2_X1 U5306 ( .A1(n7852), .A2(n4735), .ZN(n4730) );
  INV_X1 U5307 ( .A(n7673), .ZN(n4735) );
  NAND2_X1 U5308 ( .A1(n4732), .A2(n4734), .ZN(n7921) );
  NOR2_X1 U5309 ( .A1(n7857), .A2(n4733), .ZN(n4732) );
  INV_X1 U5310 ( .A(n8623), .ZN(n4733) );
  NAND2_X1 U5311 ( .A1(n7859), .A2(n8689), .ZN(n7924) );
  AOI21_X1 U5312 ( .B1(n7851), .B2(n4572), .A(n7759), .ZN(n4571) );
  NAND2_X1 U5313 ( .A1(n4725), .A2(n8641), .ZN(n4724) );
  AND2_X1 U5314 ( .A1(n7569), .A2(n7571), .ZN(n7656) );
  XNOR2_X1 U5315 ( .A(n7571), .B(n8641), .ZN(n8620) );
  NAND2_X1 U5316 ( .A1(n8911), .A2(n7600), .ZN(n8639) );
  NAND2_X1 U5317 ( .A1(n8639), .A2(n8637), .ZN(n7455) );
  AND2_X1 U5318 ( .A1(n8809), .A2(n6972), .ZN(n9266) );
  NOR2_X1 U5319 ( .A1(n7469), .A2(n7037), .ZN(n7433) );
  INV_X1 U5320 ( .A(n9228), .ZN(n9269) );
  AND2_X1 U5321 ( .A1(n10231), .A2(n4455), .ZN(n7019) );
  INV_X1 U5322 ( .A(n9266), .ZN(n9231) );
  NOR2_X1 U5323 ( .A1(n4483), .A2(n4718), .ZN(n4717) );
  NAND2_X1 U5324 ( .A1(n9126), .A2(n4719), .ZN(n4718) );
  INV_X1 U5325 ( .A(n9020), .ZN(n4719) );
  NAND2_X1 U5326 ( .A1(n5502), .A2(n5501), .ZN(n9325) );
  NAND2_X1 U5327 ( .A1(n8233), .A2(n4749), .ZN(n5168) );
  INV_X1 U5328 ( .A(n6862), .ZN(n4749) );
  AND2_X1 U5329 ( .A1(n7127), .A2(n7023), .ZN(n7421) );
  NAND2_X1 U5330 ( .A1(n4513), .A2(n4474), .ZN(n4785) );
  INV_X1 U5331 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5070) );
  NAND2_X1 U5332 ( .A1(n4513), .A2(n5065), .ZN(n4788) );
  AND2_X1 U5333 ( .A1(n4471), .A2(n5065), .ZN(n4729) );
  NAND2_X1 U5334 ( .A1(n5689), .A2(n5688), .ZN(n5687) );
  AOI21_X1 U5335 ( .B1(n8197), .B2(n5003), .A(n8198), .ZN(n5002) );
  INV_X1 U5336 ( .A(n6274), .ZN(n5003) );
  INV_X1 U5337 ( .A(n5002), .ZN(n5000) );
  NOR2_X1 U5338 ( .A1(n5911), .A2(n5910), .ZN(n5931) );
  INV_X1 U5339 ( .A(n4977), .ZN(n4974) );
  NAND2_X1 U5340 ( .A1(n7317), .A2(n7318), .ZN(n5924) );
  NOR2_X1 U5341 ( .A1(n4976), .A2(n4973), .ZN(n4972) );
  INV_X1 U5342 ( .A(n5923), .ZN(n4973) );
  NOR2_X1 U5343 ( .A1(n7538), .A2(n5941), .ZN(n4976) );
  NAND2_X1 U5344 ( .A1(n5964), .A2(n5963), .ZN(n7609) );
  NAND2_X1 U5345 ( .A1(n6441), .A2(n5844), .ZN(n5800) );
  NOR2_X1 U5346 ( .A1(n4487), .A2(n9401), .ZN(n4657) );
  INV_X1 U5347 ( .A(n4984), .ZN(n4983) );
  OAI21_X1 U5348 ( .B1(n4987), .B2(n5967), .A(n4515), .ZN(n4984) );
  XNOR2_X1 U5349 ( .A(n4967), .B(n8200), .ZN(n5827) );
  NAND2_X1 U5350 ( .A1(n4970), .A2(n4968), .ZN(n4967) );
  NAND2_X1 U5351 ( .A1(n4969), .A2(n6256), .ZN(n4968) );
  NAND2_X1 U5352 ( .A1(n5785), .A2(n5844), .ZN(n4970) );
  NAND2_X1 U5353 ( .A1(n4516), .A2(n4989), .ZN(n4988) );
  NAND2_X1 U5354 ( .A1(n4994), .A2(n8119), .ZN(n4989) );
  AND3_X1 U5355 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5886) );
  OAI21_X1 U5356 ( .B1(n8493), .B2(n10044), .A(n6468), .ZN(n4826) );
  CLKBUF_X1 U5357 ( .A(n5867), .Z(n5868) );
  OR2_X1 U5358 ( .A1(n6460), .A2(n5909), .ZN(n5915) );
  NAND2_X1 U5359 ( .A1(n4442), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U5360 ( .A1(n4546), .A2(n5774), .ZN(n5871) );
  OR2_X1 U5361 ( .A1(n9516), .A2(n9515), .ZN(n4838) );
  NAND2_X1 U5362 ( .A1(n4838), .A2(n4837), .ZN(n4836) );
  NAND2_X1 U5363 ( .A1(n9537), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4837) );
  AND2_X1 U5364 ( .A1(n4836), .A2(n4835), .ZN(n9545) );
  INV_X1 U5365 ( .A(n9539), .ZN(n4835) );
  AND4_X1 U5366 ( .A1(n6312), .A2(n6311), .A3(n6310), .A4(n6309), .ZN(n9575)
         );
  NOR2_X1 U5367 ( .A1(n9654), .A2(n9772), .ZN(n9643) );
  NOR2_X1 U5368 ( .A1(n6401), .A2(n4893), .ZN(n4892) );
  INV_X1 U5369 ( .A(n6398), .ZN(n4893) );
  OR2_X1 U5370 ( .A1(n9793), .A2(n9484), .ZN(n4667) );
  NOR2_X1 U5371 ( .A1(n6396), .A2(n4665), .ZN(n4664) );
  INV_X1 U5372 ( .A(n6395), .ZN(n4665) );
  AOI21_X1 U5373 ( .B1(n4765), .B2(n4763), .A(n4762), .ZN(n4761) );
  INV_X1 U5374 ( .A(n8419), .ZN(n4763) );
  NOR2_X1 U5375 ( .A1(n9713), .A2(n4766), .ZN(n4765) );
  INV_X1 U5376 ( .A(n6453), .ZN(n4766) );
  NAND2_X1 U5377 ( .A1(n8427), .A2(n8425), .ZN(n9713) );
  NAND2_X1 U5378 ( .A1(n4590), .A2(n4588), .ZN(n6452) );
  AOI21_X1 U5379 ( .B1(n4481), .B2(n8266), .A(n4589), .ZN(n4588) );
  OR2_X1 U5380 ( .A1(n9740), .A2(n9486), .ZN(n4887) );
  NAND2_X1 U5381 ( .A1(n9740), .A2(n9486), .ZN(n4886) );
  NAND2_X1 U5382 ( .A1(n8052), .A2(n6394), .ZN(n9728) );
  NOR2_X1 U5383 ( .A1(n8408), .A2(n4642), .ZN(n4641) );
  INV_X1 U5384 ( .A(n6393), .ZN(n4642) );
  NAND2_X1 U5385 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(n6030), .ZN(n6048) );
  NAND2_X1 U5386 ( .A1(n7805), .A2(n8301), .ZN(n7870) );
  AND2_X1 U5387 ( .A1(n6011), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U5388 ( .A1(n5987), .A2(n5986), .ZN(n7796) );
  AOI21_X1 U5389 ( .B1(n7480), .B2(n4648), .A(n4646), .ZN(n7784) );
  NAND2_X1 U5390 ( .A1(n4647), .A2(n4495), .ZN(n4646) );
  NOR2_X1 U5391 ( .A1(n10025), .A2(n4644), .ZN(n4648) );
  NAND2_X1 U5392 ( .A1(n10021), .A2(n8377), .ZN(n4769) );
  NAND2_X1 U5393 ( .A1(n7304), .A2(n6385), .ZN(n7380) );
  NAND2_X1 U5394 ( .A1(n7386), .A2(n8310), .ZN(n4760) );
  AND2_X1 U5395 ( .A1(n8354), .A2(n8353), .ZN(n7353) );
  NAND2_X1 U5396 ( .A1(n6762), .A2(n4889), .ZN(n4888) );
  INV_X1 U5397 ( .A(n5004), .ZN(n5781) );
  AND2_X1 U5398 ( .A1(n6302), .A2(n8492), .ZN(n10046) );
  NAND2_X1 U5399 ( .A1(n6204), .A2(n6203), .ZN(n9776) );
  INV_X1 U5400 ( .A(n7399), .ZN(n10111) );
  OR2_X1 U5401 ( .A1(n7244), .A2(n6468), .ZN(n10154) );
  OR2_X1 U5402 ( .A1(n5834), .A2(n6844), .ZN(n5813) );
  INV_X1 U5403 ( .A(n10149), .ZN(n10136) );
  AND4_X1 U5404 ( .A1(n6929), .A2(n6928), .A3(n6927), .A4(n6926), .ZN(n7243)
         );
  NAND2_X1 U5405 ( .A1(n5012), .A2(n5769), .ZN(n5011) );
  INV_X1 U5406 ( .A(n5743), .ZN(n5012) );
  INV_X1 U5407 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5755) );
  XNOR2_X1 U5408 ( .A(n5497), .B(n5496), .ZN(n7703) );
  NAND2_X1 U5409 ( .A1(n4807), .A2(n5474), .ZN(n5497) );
  XNOR2_X1 U5410 ( .A(n5293), .B(n5020), .ZN(n6906) );
  INV_X1 U5411 ( .A(n4821), .ZN(n5293) );
  AOI21_X1 U5412 ( .B1(n4789), .B2(n4491), .A(n4651), .ZN(n4821) );
  NAND2_X1 U5413 ( .A1(n4652), .A2(n5268), .ZN(n4651) );
  NAND2_X1 U5414 ( .A1(n4623), .A2(n5187), .ZN(n5189) );
  NAND2_X1 U5415 ( .A1(n5095), .A2(n5094), .ZN(n5098) );
  INV_X1 U5416 ( .A(n5591), .ZN(n5568) );
  NAND2_X1 U5417 ( .A1(n8563), .A2(n5490), .ZN(n8575) );
  INV_X1 U5418 ( .A(n9164), .ZN(n9017) );
  NAND2_X1 U5419 ( .A1(n5417), .A2(n5416), .ZN(n9345) );
  NAND2_X1 U5420 ( .A1(n4923), .A2(n5105), .ZN(n4921) );
  NAND2_X1 U5421 ( .A1(n5336), .A2(n7899), .ZN(n7977) );
  NAND2_X1 U5422 ( .A1(n4924), .A2(n5104), .ZN(n8820) );
  INV_X1 U5423 ( .A(n4923), .ZN(n5104) );
  XNOR2_X1 U5424 ( .A(n8609), .B(n7032), .ZN(n4686) );
  AND2_X1 U5425 ( .A1(n4964), .A2(n4526), .ZN(n8609) );
  NAND2_X1 U5426 ( .A1(n4752), .A2(n4508), .ZN(n4685) );
  OR2_X1 U5427 ( .A1(n8797), .A2(n4753), .ZN(n4752) );
  OR2_X1 U5428 ( .A1(n6970), .A2(n5690), .ZN(n10200) );
  INV_X1 U5429 ( .A(n9264), .ZN(n9233) );
  INV_X1 U5430 ( .A(n8635), .ZN(n8800) );
  INV_X1 U5431 ( .A(n8186), .ZN(n8901) );
  AOI21_X1 U5432 ( .B1(n4577), .B2(n9269), .A(n4574), .ZN(n9287) );
  NAND2_X1 U5433 ( .A1(n4576), .A2(n4575), .ZN(n4574) );
  XNOR2_X1 U5434 ( .A(n4578), .B(n9057), .ZN(n4577) );
  NAND2_X1 U5435 ( .A1(n9058), .A2(n9266), .ZN(n4576) );
  NAND2_X1 U5436 ( .A1(n5624), .A2(n5623), .ZN(n9295) );
  XNOR2_X1 U5437 ( .A(n7271), .B(n4555), .ZN(n7592) );
  AND2_X1 U5438 ( .A1(n9238), .A2(n4539), .ZN(n9246) );
  INV_X1 U5439 ( .A(n9218), .ZN(n9272) );
  INV_X1 U5440 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5068) );
  NAND2_X1 U5441 ( .A1(n5058), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5060) );
  OR2_X1 U5442 ( .A1(n6869), .A2(n5834), .ZN(n5908) );
  NAND2_X1 U5443 ( .A1(n6046), .A2(n6045), .ZN(n9808) );
  AND4_X1 U5444 ( .A1(n5958), .A2(n5957), .A3(n5956), .A4(n5955), .ZN(n7711)
         );
  AND4_X1 U5445 ( .A1(n6137), .A2(n6136), .A3(n6135), .A4(n6134), .ZN(n9717)
         );
  OAI21_X1 U5446 ( .B1(n9554), .B2(n9953), .A(n9553), .ZN(n4850) );
  OAI22_X1 U5447 ( .A1(n9550), .A2(n10003), .B1(n9552), .B2(n9969), .ZN(n4853)
         );
  INV_X1 U5448 ( .A(n9999), .ZN(n10013) );
  NAND2_X1 U5449 ( .A1(n8244), .A2(n8243), .ZN(n9876) );
  INV_X1 U5450 ( .A(n4870), .ZN(n4869) );
  INV_X1 U5451 ( .A(n4776), .ZN(n4775) );
  AOI21_X1 U5452 ( .B1(n8586), .B2(n9720), .A(n8585), .ZN(n4776) );
  INV_X1 U5453 ( .A(n4694), .ZN(n8586) );
  NAND2_X1 U5454 ( .A1(n4866), .A2(n4867), .ZN(n4777) );
  OR2_X1 U5455 ( .A1(n9570), .A2(n9569), .ZN(n9747) );
  NOR2_X1 U5456 ( .A1(n9568), .A2(n9567), .ZN(n9570) );
  NAND2_X1 U5457 ( .A1(n6412), .A2(n6411), .ZN(n9584) );
  NAND2_X1 U5458 ( .A1(n7352), .A2(n6383), .ZN(n7306) );
  OR2_X1 U5459 ( .A1(n6862), .A2(n5834), .ZN(n5880) );
  NAND2_X1 U5460 ( .A1(n4866), .A2(n4475), .ZN(n4629) );
  NAND2_X1 U5461 ( .A1(n8483), .A2(n10149), .ZN(n4693) );
  NAND2_X1 U5462 ( .A1(n4464), .A2(n4871), .ZN(n4627) );
  AOI21_X1 U5463 ( .B1(n8371), .B2(n8365), .A(n8364), .ZN(n8374) );
  NAND2_X1 U5464 ( .A1(n4751), .A2(n4750), .ZN(n8654) );
  NAND2_X1 U5465 ( .A1(n8645), .A2(n8771), .ZN(n4750) );
  OR2_X1 U5466 ( .A1(n8638), .A2(n8771), .ZN(n4751) );
  AND2_X1 U5467 ( .A1(n8407), .A2(n8408), .ZN(n4547) );
  OAI21_X1 U5468 ( .B1(n4743), .B2(n8703), .A(n4742), .ZN(n4741) );
  OAI21_X1 U5469 ( .B1(n4743), .B2(n8699), .A(n4739), .ZN(n4738) );
  NOR2_X1 U5470 ( .A1(n8708), .A2(n8707), .ZN(n4736) );
  OAI21_X1 U5471 ( .B1(n8755), .B2(n4744), .A(n4507), .ZN(n8760) );
  OAI21_X1 U5472 ( .B1(n4748), .B2(n4746), .A(n4745), .ZN(n4744) );
  AND2_X1 U5473 ( .A1(n9345), .A2(n9267), .ZN(n4783) );
  INV_X1 U5474 ( .A(n7908), .ZN(n4632) );
  OR2_X1 U5475 ( .A1(n9594), .A2(n8347), .ZN(n8533) );
  INV_X1 U5476 ( .A(n5515), .ZN(n4801) );
  INV_X1 U5477 ( .A(n4813), .ZN(n4812) );
  OAI21_X1 U5478 ( .B1(n4814), .B2(n4816), .A(n5430), .ZN(n4813) );
  INV_X1 U5479 ( .A(n4479), .ZN(n4833) );
  INV_X1 U5480 ( .A(n4920), .ZN(n4911) );
  INV_X1 U5481 ( .A(n5590), .ZN(n4909) );
  NAND2_X1 U5482 ( .A1(n8843), .A2(n4494), .ZN(n4912) );
  INV_X1 U5483 ( .A(n5595), .ZN(n4913) );
  NOR2_X1 U5484 ( .A1(n9047), .A2(n4619), .ZN(n4618) );
  NAND2_X1 U5485 ( .A1(n9033), .A2(n9071), .ZN(n4619) );
  INV_X1 U5486 ( .A(n8758), .ZN(n4949) );
  NAND2_X1 U5487 ( .A1(n4955), .A2(n4953), .ZN(n4952) );
  INV_X1 U5488 ( .A(n4954), .ZN(n4953) );
  NAND2_X1 U5489 ( .A1(n9119), .A2(n8752), .ZN(n4954) );
  AOI21_X1 U5490 ( .B1(n9170), .B2(n8593), .A(n4579), .ZN(n9133) );
  INV_X1 U5491 ( .A(n8735), .ZN(n4579) );
  NAND2_X1 U5492 ( .A1(n4613), .A2(n9013), .ZN(n4612) );
  AND2_X1 U5493 ( .A1(n5015), .A2(n8725), .ZN(n4668) );
  NOR2_X1 U5494 ( .A1(n9336), .A2(n9247), .ZN(n4613) );
  AND2_X1 U5495 ( .A1(n8162), .A2(n8161), .ZN(n4673) );
  INV_X1 U5496 ( .A(n8678), .ZN(n4572) );
  AND2_X1 U5497 ( .A1(n8643), .A2(n8639), .ZN(n8638) );
  NAND2_X1 U5498 ( .A1(n7520), .A2(n8910), .ZN(n8643) );
  AND2_X1 U5499 ( .A1(n7433), .A2(n7268), .ZN(n7279) );
  NAND2_X1 U5500 ( .A1(n9147), .A2(n4604), .ZN(n9104) );
  NOR2_X1 U5501 ( .A1(n9301), .A2(n4605), .ZN(n4604) );
  INV_X1 U5502 ( .A(n4606), .ZN(n4605) );
  INV_X1 U5503 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5688) );
  INV_X1 U5504 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5025) );
  NAND2_X1 U5505 ( .A1(n4625), .A2(n7707), .ZN(n4987) );
  NAND2_X1 U5506 ( .A1(n7611), .A2(n5967), .ZN(n4625) );
  INV_X1 U5507 ( .A(n4987), .ZN(n4986) );
  INV_X1 U5508 ( .A(n6142), .ZN(n4990) );
  NAND2_X1 U5509 ( .A1(n8291), .A2(n9876), .ZN(n8486) );
  NOR2_X1 U5510 ( .A1(n7740), .A2(n4846), .ZN(n7995) );
  AND2_X1 U5511 ( .A1(n7741), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4846) );
  NOR2_X1 U5512 ( .A1(n9571), .A2(n4774), .ZN(n4773) );
  INV_X1 U5513 ( .A(n8467), .ZN(n4774) );
  NAND2_X1 U5514 ( .A1(n4690), .A2(n6467), .ZN(n4689) );
  INV_X1 U5515 ( .A(n4691), .ZN(n4690) );
  AND2_X1 U5516 ( .A1(P1_REG3_REG_21__SCAN_IN), .A2(n6172), .ZN(n6189) );
  OR2_X1 U5517 ( .A1(n9793), .A2(n9798), .ZN(n4691) );
  NAND2_X1 U5518 ( .A1(n4884), .A2(n4886), .ZN(n4883) );
  INV_X1 U5519 ( .A(n4887), .ZN(n4884) );
  INV_X1 U5520 ( .A(n8409), .ZN(n4589) );
  NOR2_X1 U5521 ( .A1(n8086), .A2(n6093), .ZN(n6112) );
  OR2_X1 U5522 ( .A1(n7870), .A2(n8266), .ZN(n4591) );
  NOR2_X1 U5523 ( .A1(n7790), .A2(n7796), .ZN(n7791) );
  NAND2_X1 U5524 ( .A1(n8261), .A2(n6387), .ZN(n4644) );
  NAND2_X1 U5525 ( .A1(n8261), .A2(n4463), .ZN(n4647) );
  NAND2_X1 U5526 ( .A1(n8492), .A2(n4550), .ZN(n6300) );
  NOR2_X1 U5527 ( .A1(n8347), .A2(n8463), .ZN(n4595) );
  NOR2_X1 U5528 ( .A1(n4771), .A2(n4593), .ZN(n4592) );
  INV_X1 U5529 ( .A(n8293), .ZN(n4593) );
  NAND2_X1 U5530 ( .A1(n8471), .A2(n4772), .ZN(n4771) );
  NAND2_X1 U5531 ( .A1(n4597), .A2(n8471), .ZN(n4596) );
  INV_X1 U5532 ( .A(n4773), .ZN(n4597) );
  AND2_X1 U5533 ( .A1(n9584), .A2(n9482), .ZN(n6421) );
  INV_X1 U5534 ( .A(n6421), .ZN(n4876) );
  NOR3_X1 U5535 ( .A1(n7872), .A2(n9808), .A3(n8046), .ZN(n8056) );
  NOR2_X1 U5536 ( .A1(n7872), .A2(n9808), .ZN(n8042) );
  NOR2_X1 U5537 ( .A1(n7483), .A2(n7535), .ZN(n10017) );
  OAI21_X1 U5538 ( .B1(n8219), .B2(n8218), .A(n8217), .ZN(n8227) );
  INV_X1 U5539 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5742) );
  AND2_X1 U5540 ( .A1(n6336), .A2(n5644), .ZN(n6334) );
  OAI21_X1 U5541 ( .B1(n5619), .B2(n5618), .A(n5617), .ZN(n5638) );
  AND2_X1 U5542 ( .A1(n5639), .A2(n5622), .ZN(n5637) );
  NOR2_X1 U5543 ( .A1(n5408), .A2(n4817), .ZN(n4816) );
  INV_X1 U5544 ( .A(n5384), .ZN(n4817) );
  NAND2_X1 U5545 ( .A1(n4815), .A2(n5407), .ZN(n4814) );
  NAND2_X1 U5546 ( .A1(n4816), .A2(n5385), .ZN(n4815) );
  AND2_X1 U5547 ( .A1(n6026), .A2(n6025), .ZN(n6044) );
  NOR2_X1 U5548 ( .A1(n6007), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n6026) );
  OR2_X1 U5549 ( .A1(n5984), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6007) );
  XNOR2_X1 U5550 ( .A(n5315), .B(SI_11_), .ZN(n5312) );
  INV_X1 U5551 ( .A(n4823), .ZN(n4822) );
  NAND2_X1 U5552 ( .A1(n5021), .A2(n4820), .ZN(n4652) );
  AND2_X1 U5553 ( .A1(n5943), .A2(n5942), .ZN(n5946) );
  AOI21_X1 U5554 ( .B1(n5234), .B2(n4793), .A(n4514), .ZN(n4792) );
  INV_X1 U5555 ( .A(n5212), .ZN(n4793) );
  INV_X1 U5556 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U5557 ( .A1(n4755), .A2(n6850), .ZN(n4569) );
  NAND2_X1 U5558 ( .A1(n4755), .A2(n4757), .ZN(n4754) );
  NAND2_X1 U5559 ( .A1(n5077), .A2(n5795), .ZN(n5096) );
  NAND2_X1 U5560 ( .A1(n4905), .A2(n4906), .ZN(n4902) );
  OR2_X1 U5561 ( .A1(n5503), .A2(n6775), .ZN(n5524) );
  OR3_X1 U5562 ( .A1(n5349), .A2(n5348), .A3(n5347), .ZN(n5369) );
  NAND2_X1 U5563 ( .A1(n5523), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5548) );
  INV_X1 U5564 ( .A(n5524), .ZN(n5523) );
  NAND2_X1 U5565 ( .A1(n5301), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5349) );
  INV_X1 U5566 ( .A(n5302), .ZN(n5301) );
  OAI21_X1 U5567 ( .B1(n7716), .B2(n4935), .A(n5292), .ZN(n4934) );
  NAND2_X1 U5568 ( .A1(n7664), .A2(n7663), .ZN(n4935) );
  NAND2_X1 U5569 ( .A1(n7215), .A2(n4938), .ZN(n8881) );
  AND2_X1 U5570 ( .A1(n5174), .A2(n5152), .ZN(n4938) );
  OR2_X1 U5571 ( .A1(n5397), .A2(n8145), .ZN(n5419) );
  NAND2_X1 U5572 ( .A1(n4674), .A2(n8778), .ZN(n8604) );
  AND2_X1 U5573 ( .A1(n8635), .A2(n8598), .ZN(n8794) );
  AND2_X1 U5574 ( .A1(n8792), .A2(n5014), .ZN(n4753) );
  AND2_X1 U5575 ( .A1(n5655), .A2(n5654), .ZN(n9031) );
  AND4_X1 U5576 ( .A1(n5403), .A2(n5402), .A3(n5401), .A4(n5400), .ZN(n8186)
         );
  NAND2_X1 U5577 ( .A1(n5052), .A2(n5051), .ZN(n5414) );
  NOR2_X1 U5578 ( .A1(n5050), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n5051) );
  INV_X1 U5579 ( .A(n5343), .ZN(n5052) );
  AND2_X1 U5580 ( .A1(n9091), .A2(n4616), .ZN(n9000) );
  AND2_X1 U5581 ( .A1(n9880), .A2(n4618), .ZN(n4616) );
  NAND2_X1 U5582 ( .A1(n4682), .A2(n4681), .ZN(n4578) );
  NAND2_X1 U5583 ( .A1(n9059), .A2(n9264), .ZN(n4575) );
  AND2_X1 U5584 ( .A1(n5632), .A2(n5631), .ZN(n9072) );
  NOR2_X1 U5585 ( .A1(n9104), .A2(n9295), .ZN(n9091) );
  INV_X1 U5586 ( .A(n9027), .ZN(n9087) );
  OR2_X1 U5587 ( .A1(n9301), .A2(n9120), .ZN(n9025) );
  OAI21_X1 U5588 ( .B1(n9135), .B2(n4952), .A(n4950), .ZN(n9103) );
  OR2_X1 U5589 ( .A1(n9135), .A2(n4954), .ZN(n9118) );
  NAND2_X1 U5590 ( .A1(n9147), .A2(n4608), .ZN(n9141) );
  NOR2_X1 U5591 ( .A1(n9180), .A2(n9017), .ZN(n9147) );
  NAND2_X1 U5592 ( .A1(n9147), .A2(n9154), .ZN(n9148) );
  AOI21_X1 U5593 ( .B1(n9205), .B2(n9010), .A(n9009), .ZN(n9192) );
  NAND2_X1 U5594 ( .A1(n4670), .A2(n4669), .ZN(n9208) );
  NAND2_X1 U5595 ( .A1(n4671), .A2(n8725), .ZN(n4669) );
  NAND2_X1 U5596 ( .A1(n4668), .A2(n4673), .ZN(n4670) );
  NAND2_X1 U5597 ( .A1(n4480), .A2(n8591), .ZN(n4671) );
  OR2_X1 U5598 ( .A1(n5459), .A2(n5458), .ZN(n5483) );
  AND2_X1 U5599 ( .A1(n8731), .A2(n8730), .ZN(n9207) );
  AND2_X1 U5600 ( .A1(n4672), .A2(n4480), .ZN(n9225) );
  NAND2_X1 U5601 ( .A1(n4673), .A2(n5015), .ZN(n4672) );
  INV_X1 U5602 ( .A(n4673), .ZN(n9263) );
  NAND2_X1 U5603 ( .A1(n4963), .A2(n8009), .ZN(n8011) );
  NAND2_X1 U5604 ( .A1(n7767), .A2(n4536), .ZN(n8172) );
  AOI21_X1 U5605 ( .B1(n4566), .B2(n4568), .A(n4740), .ZN(n4565) );
  INV_X1 U5606 ( .A(n8700), .ZN(n4568) );
  NAND2_X1 U5607 ( .A1(n7767), .A2(n4470), .ZN(n7970) );
  NAND2_X1 U5608 ( .A1(n7767), .A2(n4615), .ZN(n7928) );
  AND4_X1 U5609 ( .A1(n5287), .A2(n5286), .A3(n5285), .A4(n5284), .ZN(n7861)
         );
  AND2_X1 U5610 ( .A1(n7767), .A2(n10260), .ZN(n7862) );
  AND2_X1 U5611 ( .A1(n8689), .A2(n8688), .ZN(n7761) );
  NOR2_X1 U5612 ( .A1(n7683), .A2(n7688), .ZN(n7767) );
  AND2_X1 U5613 ( .A1(n8683), .A2(n8691), .ZN(n7851) );
  NAND2_X1 U5614 ( .A1(n7674), .A2(n7673), .ZN(n7853) );
  AND4_X1 U5615 ( .A1(n5251), .A2(n5250), .A3(n5249), .A4(n5248), .ZN(n7754)
         );
  NAND2_X1 U5616 ( .A1(n7646), .A2(n7645), .ZN(n7647) );
  NOR2_X1 U5617 ( .A1(n7497), .A2(n10187), .ZN(n7569) );
  AND4_X1 U5618 ( .A1(n5160), .A2(n5159), .A3(n5158), .A4(n5157), .ZN(n7565)
         );
  NAND2_X1 U5619 ( .A1(n7494), .A2(n8614), .ZN(n7522) );
  INV_X1 U5620 ( .A(n8646), .ZN(n7453) );
  NAND2_X1 U5621 ( .A1(n7270), .A2(n7269), .ZN(n4778) );
  NAND2_X1 U5622 ( .A1(n4778), .A2(n8613), .ZN(n7442) );
  NAND2_X1 U5623 ( .A1(n5646), .A2(n5645), .ZN(n9290) );
  NAND2_X1 U5624 ( .A1(n5574), .A2(n5573), .ZN(n9304) );
  NOR3_X1 U5625 ( .A1(n4716), .A2(n4483), .A3(n9020), .ZN(n9127) );
  INV_X1 U5626 ( .A(n4720), .ZN(n4716) );
  OR2_X1 U5627 ( .A1(n6853), .A2(n5110), .ZN(n5146) );
  OR3_X1 U5628 ( .A1(n8789), .A2(n8800), .A3(n7032), .ZN(n10245) );
  INV_X1 U5629 ( .A(n10231), .ZN(n10273) );
  INV_X1 U5630 ( .A(n10272), .ZN(n10230) );
  INV_X1 U5631 ( .A(n8794), .ZN(n10218) );
  INV_X1 U5632 ( .A(n4788), .ZN(n4786) );
  NAND2_X1 U5633 ( .A1(n5031), .A2(n5065), .ZN(n5062) );
  OR2_X1 U5634 ( .A1(n5230), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5232) );
  OR2_X1 U5635 ( .A1(n5232), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5272) );
  NOR2_X1 U5636 ( .A1(n5137), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5190) );
  NOR2_X1 U5637 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4715) );
  INV_X1 U5638 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U5639 ( .A1(n6042), .A2(n7907), .ZN(n4982) );
  NAND2_X1 U5640 ( .A1(n4982), .A2(n6059), .ZN(n8135) );
  INV_X1 U5641 ( .A(n9410), .ZN(n5007) );
  OR2_X1 U5642 ( .A1(n9443), .A2(n6169), .ZN(n5008) );
  INV_X1 U5643 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8086) );
  XNOR2_X1 U5644 ( .A(n5843), .B(n6226), .ZN(n5845) );
  OAI22_X1 U5645 ( .A1(n7263), .A2(n8199), .B1(n7387), .B2(n5802), .ZN(n5843)
         );
  NAND2_X1 U5646 ( .A1(n6922), .A2(n6921), .ZN(n6920) );
  NOR2_X1 U5647 ( .A1(n6024), .A2(n4637), .ZN(n4636) );
  INV_X1 U5648 ( .A(n6006), .ZN(n4637) );
  NAND2_X1 U5649 ( .A1(n4638), .A2(n4498), .ZN(n4635) );
  NAND2_X1 U5650 ( .A1(n4993), .A2(n4485), .ZN(n4992) );
  INV_X1 U5651 ( .A(n9426), .ZN(n4993) );
  AND2_X1 U5652 ( .A1(n6273), .A2(n6272), .ZN(n6274) );
  NAND2_X1 U5653 ( .A1(n6060), .A2(n8134), .ZN(n4978) );
  AND4_X1 U5654 ( .A1(n5936), .A2(n5935), .A3(n5934), .A4(n5933), .ZN(n7612)
         );
  OR2_X1 U5655 ( .A1(n6824), .A2(n6823), .ZN(n4845) );
  NAND2_X1 U5656 ( .A1(n4845), .A2(n4844), .ZN(n9988) );
  NAND2_X1 U5657 ( .A1(n6796), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4844) );
  NOR2_X1 U5658 ( .A1(n6829), .A2(n4531), .ZN(n10006) );
  NOR2_X1 U5659 ( .A1(n10006), .A2(n10005), .ZN(n10004) );
  AND2_X1 U5660 ( .A1(n9507), .A2(n6785), .ZN(n6790) );
  NOR2_X1 U5661 ( .A1(n7164), .A2(n4842), .ZN(n7165) );
  AND2_X1 U5662 ( .A1(n7171), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4842) );
  NAND2_X1 U5663 ( .A1(n7165), .A2(n7166), .ZN(n7334) );
  XNOR2_X1 U5664 ( .A(n7995), .B(n7994), .ZN(n7742) );
  NOR2_X1 U5665 ( .A1(n8483), .A2(n9580), .ZN(n9562) );
  INV_X1 U5666 ( .A(n8282), .ZN(n4879) );
  NAND2_X1 U5667 ( .A1(n9608), .A2(n6405), .ZN(n9595) );
  NAND2_X1 U5668 ( .A1(n9595), .A2(n9594), .ZN(n9593) );
  NAND2_X1 U5669 ( .A1(n4700), .A2(n9598), .ZN(n4699) );
  AND4_X1 U5670 ( .A1(n6420), .A2(n6419), .A3(n6418), .A4(n6417), .ZN(n9589)
         );
  NOR2_X1 U5671 ( .A1(n9654), .A2(n4698), .ZN(n9612) );
  INV_X1 U5672 ( .A(n4700), .ZN(n4698) );
  NOR2_X1 U5673 ( .A1(n9654), .A2(n4701), .ZN(n9622) );
  AND2_X1 U5674 ( .A1(n8458), .A2(n8459), .ZN(n9632) );
  AND2_X1 U5675 ( .A1(n6205), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U5676 ( .A1(n6219), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6241) );
  NOR2_X1 U5677 ( .A1(n9719), .A2(n4689), .ZN(n9689) );
  INV_X1 U5678 ( .A(n4662), .ZN(n4661) );
  OAI21_X1 U5679 ( .B1(n4664), .B2(n4663), .A(n6397), .ZN(n4662) );
  OR2_X1 U5680 ( .A1(n8248), .A2(n8247), .ZN(n9675) );
  NAND2_X1 U5681 ( .A1(n4765), .A2(n8329), .ZN(n4581) );
  OR2_X1 U5682 ( .A1(n4761), .A2(n4582), .ZN(n4580) );
  NOR2_X1 U5683 ( .A1(n9719), .A2(n4691), .ZN(n9697) );
  NOR2_X1 U5684 ( .A1(n9719), .A2(n9798), .ZN(n9718) );
  INV_X1 U5685 ( .A(n6132), .ZN(n6133) );
  NOR2_X1 U5686 ( .A1(n4705), .A2(n4706), .ZN(n4703) );
  OR2_X1 U5687 ( .A1(n8046), .A2(n9740), .ZN(n4705) );
  AOI21_X1 U5688 ( .B1(n4641), .B2(n4467), .A(n4509), .ZN(n4640) );
  NAND2_X1 U5689 ( .A1(n4591), .A2(n4481), .ZN(n8049) );
  AND2_X1 U5690 ( .A1(n4591), .A2(n8403), .ZN(n8035) );
  AND4_X1 U5691 ( .A1(n6097), .A2(n6096), .A3(n6095), .A4(n6094), .ZN(n9427)
         );
  INV_X1 U5692 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6716) );
  OR2_X1 U5693 ( .A1(n7811), .A2(n7915), .ZN(n7872) );
  NAND2_X1 U5694 ( .A1(n7807), .A2(n6451), .ZN(n7805) );
  AOI21_X1 U5695 ( .B1(n8265), .B2(n4859), .A(n4505), .ZN(n4860) );
  AND4_X1 U5696 ( .A1(n6016), .A2(n6015), .A3(n6014), .A4(n6013), .ZN(n7912)
         );
  NAND2_X1 U5697 ( .A1(n10017), .A2(n10030), .ZN(n10016) );
  OR2_X1 U5698 ( .A1(n5952), .A2(n5951), .ZN(n5971) );
  NAND2_X1 U5699 ( .A1(n4758), .A2(n4587), .ZN(n4586) );
  INV_X1 U5700 ( .A(n4758), .ZN(n4583) );
  NAND2_X1 U5701 ( .A1(n4585), .A2(n4584), .ZN(n7372) );
  NAND2_X1 U5702 ( .A1(n10137), .A2(n4687), .ZN(n7483) );
  OR2_X1 U5703 ( .A1(n6865), .A2(n5834), .ZN(n5894) );
  AND2_X1 U5704 ( .A1(n8370), .A2(n8308), .ZN(n8359) );
  NAND2_X1 U5705 ( .A1(n8307), .A2(n8509), .ZN(n7255) );
  OR2_X1 U5706 ( .A1(n9499), .A2(n5816), .ZN(n6377) );
  NAND2_X1 U5707 ( .A1(n8256), .A2(n10038), .ZN(n6376) );
  INV_X1 U5708 ( .A(n9499), .ZN(n7289) );
  OR2_X1 U5709 ( .A1(n4695), .A2(n9562), .ZN(n4694) );
  INV_X1 U5710 ( .A(n4696), .ZN(n4695) );
  AOI21_X1 U5711 ( .B1(n9580), .B2(n8483), .A(n10154), .ZN(n4696) );
  NAND2_X1 U5712 ( .A1(n6407), .A2(n6406), .ZN(n9756) );
  NAND2_X1 U5713 ( .A1(n6217), .A2(n6216), .ZN(n9772) );
  NAND2_X1 U5714 ( .A1(n7480), .A2(n6387), .ZN(n10026) );
  OR2_X1 U5715 ( .A1(n5834), .A2(n6846), .ZN(n5754) );
  XNOR2_X1 U5716 ( .A(n8227), .B(n8226), .ZN(n8588) );
  XNOR2_X1 U5717 ( .A(n8219), .B(n6428), .ZN(n9378) );
  XNOR2_X1 U5718 ( .A(n6335), .B(n6334), .ZN(n8576) );
  XNOR2_X1 U5719 ( .A(n5601), .B(n5596), .ZN(n8020) );
  XNOR2_X1 U5720 ( .A(n5780), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6438) );
  NAND2_X1 U5721 ( .A1(n5778), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U5722 ( .A1(n5762), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U5723 ( .A1(n5765), .A2(n5764), .ZN(n5778) );
  INV_X1 U5724 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5764) );
  INV_X1 U5725 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U5726 ( .A1(n4799), .A2(n4802), .ZN(n5516) );
  OR2_X1 U5727 ( .A1(n5472), .A2(n4804), .ZN(n4799) );
  OAI21_X1 U5728 ( .B1(n5386), .B2(n5385), .A(n5384), .ZN(n5409) );
  XNOR2_X1 U5729 ( .A(n5386), .B(n5381), .ZN(n7194) );
  NAND2_X1 U5730 ( .A1(n4831), .A2(n5339), .ZN(n5359) );
  NAND2_X1 U5731 ( .A1(n5255), .A2(n5254), .ZN(n5267) );
  OR2_X1 U5732 ( .A1(n5892), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5906) );
  XNOR2_X1 U5733 ( .A(n5141), .B(SI_3_), .ZN(n5139) );
  OAI211_X1 U5734 ( .C1(n5074), .C2(n6845), .A(n4895), .B(n4894), .ZN(n5094)
         );
  NAND2_X1 U5735 ( .A1(n4896), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4895) );
  INV_X1 U5736 ( .A(n5073), .ZN(n4896) );
  AND4_X1 U5737 ( .A1(n5229), .A2(n5228), .A3(n5227), .A4(n5226), .ZN(n7677)
         );
  OR2_X1 U5738 ( .A1(n8868), .A2(n6340), .ZN(n8892) );
  OAI21_X1 U5739 ( .B1(n7666), .B2(n7664), .A(n7663), .ZN(n7717) );
  INV_X1 U5740 ( .A(n4915), .ZN(n6327) );
  NAND2_X1 U5741 ( .A1(n7215), .A2(n5152), .ZN(n6814) );
  AND4_X1 U5742 ( .A1(n5424), .A2(n5423), .A3(n5422), .A4(n5421), .ZN(n9232)
         );
  INV_X1 U5743 ( .A(n9247), .ZN(n9006) );
  NAND2_X1 U5744 ( .A1(n5429), .A2(n5428), .ZN(n6766) );
  OR2_X1 U5745 ( .A1(n8570), .A2(n9233), .ZN(n8875) );
  NAND2_X1 U5746 ( .A1(n8575), .A2(n5494), .ZN(n6773) );
  NAND2_X1 U5747 ( .A1(n4929), .A2(n4933), .ZN(n7748) );
  NAND2_X1 U5748 ( .A1(n7666), .A2(n4936), .ZN(n4929) );
  NAND2_X1 U5749 ( .A1(n5103), .A2(n5105), .ZN(n4923) );
  NAND2_X1 U5750 ( .A1(n7976), .A2(n4903), .ZN(n4901) );
  INV_X1 U5751 ( .A(n4904), .ZN(n4903) );
  OAI211_X1 U5752 ( .C1(n6888), .C2(n5580), .A(n5579), .B(n5578), .ZN(n9136)
         );
  INV_X1 U5753 ( .A(n7927), .ZN(n8904) );
  INV_X1 U5754 ( .A(n7677), .ZN(n8907) );
  NAND2_X1 U5755 ( .A1(n8807), .A2(n4473), .ZN(n4941) );
  INV_X2 U5756 ( .A(P2_U3966), .ZN(n8913) );
  NAND2_X1 U5757 ( .A1(n8236), .A2(n8235), .ZN(n9275) );
  XNOR2_X1 U5758 ( .A(n9000), .B(n8237), .ZN(n9277) );
  INV_X1 U5759 ( .A(n9275), .ZN(n8237) );
  NAND2_X1 U5760 ( .A1(n4676), .A2(n4677), .ZN(n9037) );
  INV_X1 U5761 ( .A(n9290), .ZN(n9071) );
  INV_X1 U5762 ( .A(n9304), .ZN(n9117) );
  NAND2_X1 U5763 ( .A1(n9309), .A2(n9023), .ZN(n9113) );
  NAND2_X1 U5764 ( .A1(n5567), .A2(n5566), .ZN(n9311) );
  OAI21_X1 U5765 ( .B1(n4721), .B2(n4723), .A(n9019), .ZN(n9146) );
  INV_X1 U5766 ( .A(n9162), .ZN(n4721) );
  AND2_X1 U5767 ( .A1(n5520), .A2(n5519), .ZN(n9164) );
  NAND2_X1 U5768 ( .A1(n4956), .A2(n8745), .ZN(n9172) );
  NAND2_X1 U5769 ( .A1(n8592), .A2(n8740), .ZN(n9185) );
  NAND2_X1 U5770 ( .A1(n5481), .A2(n5480), .ZN(n9332) );
  NOR2_X1 U5771 ( .A1(n9235), .A2(n9247), .ZN(n9214) );
  NAND2_X1 U5772 ( .A1(n4562), .A2(n8168), .ZN(n8169) );
  AND2_X1 U5773 ( .A1(n4562), .A2(n4560), .ZN(n9005) );
  NAND2_X1 U5774 ( .A1(n4780), .A2(n4779), .ZN(n4562) );
  INV_X1 U5775 ( .A(n4780), .ZN(n9252) );
  INV_X1 U5776 ( .A(n4726), .ZN(n8167) );
  NAND2_X1 U5777 ( .A1(n7924), .A2(n8700), .ZN(n7965) );
  AND2_X1 U5778 ( .A1(n4734), .A2(n4731), .ZN(n7858) );
  INV_X1 U5779 ( .A(n7857), .ZN(n4731) );
  OR2_X1 U5780 ( .A1(n7598), .A2(n10273), .ZN(n9218) );
  AND2_X1 U5781 ( .A1(n5193), .A2(n5192), .ZN(n4683) );
  OR2_X1 U5782 ( .A1(n6865), .A2(n5110), .ZN(n4684) );
  CLKBUF_X1 U5783 ( .A(n7493), .Z(n7448) );
  XNOR2_X1 U5784 ( .A(n7454), .B(n4555), .ZN(n7277) );
  AND2_X1 U5785 ( .A1(n7036), .A2(n4603), .ZN(n7623) );
  INV_X1 U5786 ( .A(n7433), .ZN(n4603) );
  OR2_X1 U5787 ( .A1(n7129), .A2(n7128), .ZN(n10292) );
  AND2_X2 U5788 ( .A1(n7024), .A2(n7421), .ZN(n10281) );
  AND2_X1 U5789 ( .A1(n6895), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10216) );
  NOR2_X1 U5790 ( .A1(n5034), .A2(n4785), .ZN(n4784) );
  NAND2_X1 U5791 ( .A1(n5031), .A2(n4787), .ZN(n4602) );
  NOR2_X1 U5792 ( .A1(n4788), .A2(n5034), .ZN(n4787) );
  NAND2_X1 U5793 ( .A1(n5672), .A2(n5671), .ZN(n8182) );
  INV_X1 U5794 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8023) );
  XNOR2_X1 U5795 ( .A(n5666), .B(n5665), .ZN(n8025) );
  INV_X1 U5796 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7880) );
  INV_X1 U5797 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7802) );
  INV_X1 U5798 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7734) );
  INV_X1 U5799 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7706) );
  INV_X1 U5800 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7359) );
  INV_X1 U5801 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7213) );
  INV_X1 U5802 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7193) );
  INV_X1 U5803 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6916) );
  INV_X1 U5804 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6905) );
  INV_X1 U5805 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6874) );
  INV_X1 U5806 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6870) );
  INV_X1 U5807 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6863) );
  OR2_X1 U5808 ( .A1(n5797), .A2(n6760), .ZN(n6807) );
  AND4_X1 U5809 ( .A1(n5891), .A2(n5890), .A3(n5889), .A4(n5888), .ZN(n7344)
         );
  AND4_X1 U5810 ( .A1(n6264), .A2(n6263), .A3(n6262), .A4(n6261), .ZN(n9634)
         );
  AND2_X1 U5811 ( .A1(n9384), .A2(n8197), .ZN(n9386) );
  OR2_X1 U5812 ( .A1(n4982), .A2(n6059), .ZN(n8137) );
  NAND2_X1 U5813 ( .A1(n7609), .A2(n5967), .ZN(n7708) );
  NOR2_X1 U5814 ( .A1(n9463), .A2(n9468), .ZN(n9403) );
  AND4_X1 U5815 ( .A1(n6436), .A2(n6435), .A3(n6434), .A4(n6433), .ZN(n9574)
         );
  NOR2_X1 U5816 ( .A1(n8205), .A2(n5000), .ZN(n4997) );
  OAI22_X1 U5817 ( .A1(n5000), .A2(n4999), .B1(n8205), .B2(n5002), .ZN(n4998)
         );
  NOR2_X1 U5818 ( .A1(n8197), .A2(n8205), .ZN(n4999) );
  NAND2_X1 U5819 ( .A1(n8197), .A2(n8205), .ZN(n5001) );
  NAND2_X1 U5820 ( .A1(n4974), .A2(n5941), .ZN(n7537) );
  INV_X1 U5821 ( .A(n5008), .ZN(n9411) );
  AND4_X1 U5822 ( .A1(n6035), .A2(n6034), .A3(n6033), .A4(n6032), .ZN(n7887)
         );
  NAND2_X1 U5823 ( .A1(n7725), .A2(n6006), .ZN(n7776) );
  AND4_X1 U5824 ( .A1(n6076), .A2(n6075), .A3(n6074), .A4(n6073), .ZN(n8133)
         );
  NAND2_X1 U5825 ( .A1(n4995), .A2(n8120), .ZN(n9425) );
  AND4_X1 U5826 ( .A1(n6213), .A2(n6212), .A3(n6211), .A4(n6210), .ZN(n9456)
         );
  INV_X1 U5827 ( .A(n7538), .ZN(n4975) );
  AND2_X1 U5828 ( .A1(n4487), .A2(n9401), .ZN(n4656) );
  NAND2_X1 U5829 ( .A1(n4630), .A2(n4635), .ZN(n7910) );
  NAND2_X1 U5830 ( .A1(n7725), .A2(n4636), .ZN(n4630) );
  AND4_X1 U5831 ( .A1(n5976), .A2(n5975), .A3(n5974), .A4(n5973), .ZN(n7787)
         );
  CLKBUF_X1 U5832 ( .A(n7724), .Z(n7725) );
  AND2_X1 U5833 ( .A1(n9430), .A2(n10149), .ZN(n9459) );
  NAND2_X1 U5834 ( .A1(n6317), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9472) );
  NAND2_X1 U5835 ( .A1(n6318), .A2(n6788), .ZN(n9455) );
  INV_X1 U5836 ( .A(n9461), .ZN(n9467) );
  CLKBUF_X1 U5837 ( .A(n6301), .Z(n6302) );
  AOI21_X1 U5838 ( .B1(n4829), .B2(n8494), .A(n4826), .ZN(n4825) );
  AND2_X1 U5839 ( .A1(n8544), .A2(n5019), .ZN(n8494) );
  NAND4_X1 U5840 ( .A1(n5916), .A2(n5915), .A3(n5914), .A4(n5913), .ZN(n9493)
         );
  NAND2_X1 U5841 ( .A1(n5788), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5792) );
  XNOR2_X1 U5842 ( .A(n4848), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9966) );
  NAND2_X1 U5843 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4848) );
  AND2_X1 U5844 ( .A1(n5751), .A2(n5832), .ZN(n9984) );
  INV_X1 U5845 ( .A(n4845), .ZN(n6822) );
  OAI22_X1 U5846 ( .A1(n9988), .A2(n9989), .B1(n4889), .B2(
        P1_REG2_REG_4__SCAN_IN), .ZN(n6831) );
  NOR2_X1 U5847 ( .A1(n10004), .A2(n4839), .ZN(n6877) );
  NOR2_X1 U5848 ( .A1(n4841), .A2(n4840), .ZN(n4839) );
  INV_X1 U5849 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n4840) );
  INV_X1 U5850 ( .A(n10011), .ZN(n4841) );
  NAND2_X1 U5851 ( .A1(n6877), .A2(n6876), .ZN(n6875) );
  AND2_X1 U5852 ( .A1(n6790), .A2(n6789), .ZN(n7070) );
  NOR2_X1 U5853 ( .A1(n7074), .A2(n7073), .ZN(n7164) );
  NOR2_X1 U5854 ( .A1(n4843), .A2(n7070), .ZN(n7074) );
  AND2_X1 U5855 ( .A1(n7071), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4843) );
  NOR2_X1 U5856 ( .A1(n7513), .A2(n7512), .ZN(n7740) );
  NOR2_X1 U5857 ( .A1(n7510), .A2(n4847), .ZN(n7513) );
  AND2_X1 U5858 ( .A1(n7511), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4847) );
  INV_X1 U5859 ( .A(n4838), .ZN(n9536) );
  INV_X1 U5860 ( .A(n4836), .ZN(n9540) );
  INV_X1 U5861 ( .A(n8286), .ZN(n9901) );
  NAND2_X1 U5862 ( .A1(n6455), .A2(n8458), .ZN(n9605) );
  NAND2_X1 U5863 ( .A1(n6399), .A2(n6398), .ZN(n9638) );
  NAND2_X1 U5864 ( .A1(n4660), .A2(n4667), .ZN(n9684) );
  NAND2_X1 U5865 ( .A1(n4666), .A2(n4664), .ZN(n4660) );
  OAI21_X1 U5866 ( .B1(n9730), .B2(n4764), .A(n4761), .ZN(n9705) );
  NAND2_X1 U5867 ( .A1(n4666), .A2(n6395), .ZN(n9696) );
  NAND2_X1 U5868 ( .A1(n4767), .A2(n6453), .ZN(n9712) );
  NAND2_X1 U5869 ( .A1(n9728), .A2(n4887), .ZN(n4882) );
  NAND2_X1 U5870 ( .A1(n6092), .A2(n6091), .ZN(n8060) );
  NAND2_X1 U5871 ( .A1(n4643), .A2(n6393), .ZN(n8039) );
  OR2_X1 U5872 ( .A1(n7869), .A2(n4467), .ZN(n4643) );
  NAND2_X1 U5873 ( .A1(n7784), .A2(n6389), .ZN(n4861) );
  NAND2_X1 U5874 ( .A1(n4769), .A2(n8376), .ZN(n7693) );
  NAND2_X1 U5875 ( .A1(n4620), .A2(n5969), .ZN(n7699) );
  NAND2_X1 U5876 ( .A1(n6906), .A2(n8283), .ZN(n4620) );
  AOI21_X1 U5877 ( .B1(n7480), .B2(n4649), .A(n4463), .ZN(n4645) );
  NOR2_X1 U5878 ( .A1(n10025), .A2(n4650), .ZN(n4649) );
  NAND2_X1 U5879 ( .A1(n4855), .A2(n4854), .ZN(n4856) );
  NAND2_X1 U5880 ( .A1(n8355), .A2(n6382), .ZN(n4854) );
  INV_X1 U5881 ( .A(n9746), .ZN(n9611) );
  NAND2_X1 U5882 ( .A1(n4857), .A2(n6382), .ZN(n7354) );
  NAND2_X1 U5883 ( .A1(n4890), .A2(n4502), .ZN(n7399) );
  NAND2_X1 U5884 ( .A1(n4692), .A2(n8283), .ZN(n4890) );
  INV_X1 U5885 ( .A(n6853), .ZN(n4692) );
  AOI211_X1 U5886 ( .C1(n10149), .C2(n9876), .A(n9903), .B(n9875), .ZN(n9878)
         );
  OR2_X1 U5887 ( .A1(n9747), .A2(n10141), .ZN(n9753) );
  AND2_X2 U5888 ( .A1(n7243), .A2(n6930), .ZN(n10160) );
  AND2_X1 U5889 ( .A1(n5797), .A2(n6295), .ZN(n6928) );
  NAND2_X1 U5890 ( .A1(n5010), .A2(n4599), .ZN(n5009) );
  INV_X1 U5891 ( .A(n5011), .ZN(n5010) );
  CLKBUF_X1 U5892 ( .A(n6461), .Z(n9977) );
  XNOR2_X1 U5893 ( .A(n5757), .B(P1_IR_REG_26__SCAN_IN), .ZN(n8158) );
  INV_X1 U5894 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8021) );
  INV_X1 U5895 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7993) );
  XNOR2_X1 U5896 ( .A(n5570), .B(n5569), .ZN(n7989) );
  INV_X1 U5897 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7878) );
  INV_X1 U5898 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7783) );
  INV_X1 U5899 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7704) );
  INV_X1 U5900 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7467) );
  INV_X1 U5901 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7384) );
  INV_X1 U5902 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7195) );
  INV_X1 U5903 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7204) );
  INV_X1 U5904 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7042) );
  INV_X1 U5905 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6917) );
  INV_X1 U5906 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6900) );
  INV_X1 U5907 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6872) );
  INV_X1 U5908 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6868) );
  NAND2_X1 U5909 ( .A1(n5189), .A2(n5209), .ZN(n4795) );
  INV_X1 U5910 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6861) );
  NAND2_X1 U5911 ( .A1(n4621), .A2(n5166), .ZN(n5184) );
  INV_X1 U5912 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6852) );
  INV_X1 U5913 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6848) );
  NOR2_X1 U5914 ( .A1(n7842), .A2(n10331), .ZN(n10321) );
  AOI21_X1 U5915 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10319), .ZN(n10318) );
  NOR2_X1 U5916 ( .A1(n10318), .A2(n10317), .ZN(n10316) );
  INV_X1 U5917 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8998) );
  OR2_X1 U5918 ( .A1(n6374), .A2(n6373), .ZN(P2_U3242) );
  NAND2_X1 U5919 ( .A1(n9295), .A2(n8890), .ZN(n6372) );
  AOI21_X1 U5920 ( .B1(n4686), .B2(n8798), .A(n4685), .ZN(n8804) );
  NOR2_X1 U5921 ( .A1(n9287), .A2(n10198), .ZN(n9060) );
  NOR2_X1 U5922 ( .A1(n6807), .A2(P1_U3084), .ZN(P1_U4006) );
  AOI21_X1 U5923 ( .B1(n10013), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9555), .ZN(
        n4851) );
  NAND2_X1 U5924 ( .A1(n4853), .A2(n9644), .ZN(n4852) );
  NAND2_X1 U5925 ( .A1(n4850), .A2(n10044), .ZN(n4849) );
  AOI21_X1 U5926 ( .B1(n4777), .B2(n10031), .A(n4775), .ZN(n8587) );
  NOR2_X1 U5927 ( .A1(n4869), .A2(n4872), .ZN(n4868) );
  OAI211_X1 U5928 ( .C1(n4627), .C2(n10171), .A(n6478), .B(n4626), .ZN(n6759)
         );
  NAND2_X1 U5929 ( .A1(n4627), .A2(n4628), .ZN(n9812) );
  INV_X1 U5930 ( .A(n4629), .ZN(n4628) );
  NOR2_X1 U5931 ( .A1(n10150), .A2(n9492), .ZN(n4463) );
  AND3_X1 U5932 ( .A1(n4873), .A2(n4870), .A3(n10156), .ZN(n4464) );
  INV_X2 U5933 ( .A(n5522), .ZN(n5204) );
  XNOR2_X1 U5934 ( .A(n9290), .B(n9031), .ZN(n9075) );
  XNOR2_X1 U5935 ( .A(n6456), .B(n8282), .ZN(n4465) );
  OR2_X1 U5936 ( .A1(n6308), .A2(n7293), .ZN(n4466) );
  AND2_X1 U5937 ( .A1(n9808), .A2(n9488), .ZN(n4467) );
  AND2_X1 U5938 ( .A1(n8249), .A2(n4883), .ZN(n4469) );
  NAND2_X1 U5939 ( .A1(n5380), .A2(n4907), .ZN(n4906) );
  INV_X1 U5940 ( .A(n8361), .ZN(n4584) );
  INV_X1 U5941 ( .A(n6064), .ZN(n6762) );
  AND2_X1 U5942 ( .A1(n4615), .A2(n4614), .ZN(n4470) );
  AND2_X1 U5943 ( .A1(n4513), .A2(n5067), .ZN(n4471) );
  AND2_X1 U5944 ( .A1(n9157), .A2(n9018), .ZN(n4472) );
  AND2_X1 U5945 ( .A1(n5044), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4473) );
  AND2_X1 U5946 ( .A1(n5065), .A2(n5070), .ZN(n4474) );
  NAND2_X1 U5947 ( .A1(n5457), .A2(n5456), .ZN(n9336) );
  AND2_X1 U5948 ( .A1(n4694), .A2(n4503), .ZN(n4475) );
  INV_X1 U5949 ( .A(n8329), .ZN(n4582) );
  XNOR2_X1 U5950 ( .A(n5039), .B(n5038), .ZN(n5042) );
  OR2_X1 U5951 ( .A1(n5007), .A2(n5017), .ZN(n4476) );
  AND2_X1 U5952 ( .A1(n6384), .A2(n6383), .ZN(n4477) );
  INV_X1 U5953 ( .A(n4873), .ZN(n4872) );
  OAI21_X1 U5954 ( .B1(n4879), .B2(n6421), .A(n4874), .ZN(n4873) );
  NAND2_X1 U5955 ( .A1(n7479), .A2(n7478), .ZN(n7480) );
  INV_X1 U5956 ( .A(n10044), .ZN(n9644) );
  INV_X2 U5957 ( .A(n5867), .ZN(n5808) );
  NAND2_X4 U5958 ( .A1(n5045), .A2(n5044), .ZN(n5129) );
  AND2_X1 U5959 ( .A1(n5360), .A2(n5342), .ZN(n4479) );
  OR2_X1 U5960 ( .A1(n8628), .A2(n8716), .ZN(n4480) );
  NAND2_X1 U5961 ( .A1(n6067), .A2(n6066), .ZN(n8046) );
  AND2_X1 U5962 ( .A1(n8408), .A2(n8403), .ZN(n4481) );
  NAND4_X1 U5963 ( .A1(n5109), .A2(n5108), .A3(n5107), .A4(n5106), .ZN(n8912)
         );
  NAND2_X1 U5964 ( .A1(n8575), .A2(n4925), .ZN(n6771) );
  NAND2_X1 U5965 ( .A1(n5026), .A2(n5025), .ZN(n5137) );
  AND2_X1 U5966 ( .A1(n4915), .A2(n4914), .ZN(n4482) );
  AND2_X1 U5967 ( .A1(n9157), .A2(n4722), .ZN(n4483) );
  AND2_X1 U5968 ( .A1(n8377), .A2(n8376), .ZN(n10025) );
  AND2_X1 U5969 ( .A1(n4792), .A2(n4653), .ZN(n4484) );
  NAND2_X1 U5970 ( .A1(n8292), .A2(n8534), .ZN(n8282) );
  NAND2_X1 U5971 ( .A1(n9085), .A2(n8764), .ZN(n9098) );
  INV_X1 U5972 ( .A(n9098), .ZN(n4955) );
  NAND2_X1 U5973 ( .A1(n6445), .A2(n8509), .ZN(n7386) );
  OR2_X1 U5974 ( .A1(n9247), .A2(n8874), .ZN(n8725) );
  NAND2_X1 U5975 ( .A1(n6124), .A2(n6123), .ZN(n4485) );
  INV_X1 U5976 ( .A(n5775), .ZN(n4546) );
  NAND3_X1 U5977 ( .A1(n5046), .A2(n6952), .A3(n6950), .ZN(n7025) );
  NAND2_X1 U5978 ( .A1(n4891), .A2(n6400), .ZN(n9621) );
  NOR4_X1 U5979 ( .A1(n9057), .A2(n8632), .A3(n9075), .A4(n9027), .ZN(n4486)
         );
  NAND3_X1 U5980 ( .A1(n4943), .A2(n5080), .A3(n4941), .ZN(n6954) );
  XNOR2_X1 U5981 ( .A(n8200), .B(n6153), .ZN(n4487) );
  INV_X1 U5982 ( .A(n8641), .ZN(n8909) );
  AND4_X1 U5983 ( .A1(n5182), .A2(n5181), .A3(n5180), .A4(n5179), .ZN(n8641)
         );
  INV_X1 U5984 ( .A(n8701), .ZN(n4740) );
  OR2_X1 U5985 ( .A1(n4975), .A2(n5940), .ZN(n4488) );
  NAND2_X1 U5986 ( .A1(n8467), .A2(n8456), .ZN(n9594) );
  INV_X1 U5987 ( .A(n9594), .ZN(n4772) );
  INV_X1 U5988 ( .A(n6256), .ZN(n8199) );
  NAND2_X1 U5989 ( .A1(n6339), .A2(n6338), .ZN(n8596) );
  INV_X1 U5990 ( .A(n8596), .ZN(n9033) );
  NAND2_X1 U5991 ( .A1(n4871), .A2(n4868), .ZN(n8580) );
  AND2_X1 U5992 ( .A1(n4684), .A2(n4683), .ZN(n7571) );
  INV_X1 U5993 ( .A(n7571), .ZN(n10229) );
  INV_X1 U5994 ( .A(n5404), .ZN(n4907) );
  OR2_X1 U5995 ( .A1(n8711), .A2(n9265), .ZN(n4489) );
  NAND2_X1 U5996 ( .A1(n8779), .A2(n8778), .ZN(n9038) );
  INV_X1 U5997 ( .A(n9038), .ZN(n4675) );
  OR2_X1 U5998 ( .A1(n5380), .A2(n4907), .ZN(n4490) );
  NAND2_X1 U5999 ( .A1(n5238), .A2(n6606), .ZN(n5254) );
  INV_X1 U6000 ( .A(n5254), .ZN(n4820) );
  NAND2_X1 U6001 ( .A1(n5546), .A2(n5545), .ZN(n9316) );
  AND2_X1 U6002 ( .A1(n4484), .A2(n5021), .ZN(n4491) );
  NAND2_X1 U6003 ( .A1(n5004), .A2(n4468), .ZN(n5759) );
  OR2_X1 U6004 ( .A1(n9768), .A2(n9438), .ZN(n8458) );
  AND2_X1 U6005 ( .A1(n5311), .A2(n5310), .ZN(n4492) );
  AND2_X1 U6006 ( .A1(n9591), .A2(n4773), .ZN(n4493) );
  INV_X1 U6007 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9826) );
  INV_X1 U6008 ( .A(n9262), .ZN(n4779) );
  AND2_X1 U6009 ( .A1(n8715), .A2(n8716), .ZN(n9262) );
  NOR2_X1 U6010 ( .A1(n6326), .A2(n4913), .ZN(n4494) );
  NAND2_X1 U6011 ( .A1(n6255), .A2(n6254), .ZN(n9761) );
  NAND2_X1 U6012 ( .A1(n6188), .A2(n6187), .ZN(n9781) );
  OR2_X1 U6013 ( .A1(n7699), .A2(n10023), .ZN(n4495) );
  NAND2_X1 U6014 ( .A1(n5607), .A2(n5606), .ZN(n9301) );
  OR2_X1 U6015 ( .A1(n9891), .A2(n8093), .ZN(n4496) );
  NOR2_X1 U6016 ( .A1(n9654), .A2(n4699), .ZN(n4697) );
  INV_X1 U6017 ( .A(n6387), .ZN(n4650) );
  OR2_X1 U6018 ( .A1(n4448), .A2(n10059), .ZN(n4497) );
  NAND2_X1 U6019 ( .A1(n6171), .A2(n6170), .ZN(n9788) );
  AND2_X1 U6020 ( .A1(n6022), .A2(n7773), .ZN(n4498) );
  INV_X1 U6021 ( .A(n5268), .ZN(n4824) );
  AND2_X1 U6022 ( .A1(n4767), .A2(n4765), .ZN(n4499) );
  AND2_X1 U6023 ( .A1(n4959), .A2(n8745), .ZN(n4500) );
  NAND2_X1 U6024 ( .A1(n9017), .A2(n9187), .ZN(n9018) );
  AND2_X1 U6025 ( .A1(n4879), .A2(n4876), .ZN(n4501) );
  AND2_X1 U6026 ( .A1(n5859), .A2(n4888), .ZN(n4502) );
  INV_X1 U6027 ( .A(n9047), .ZN(n9279) );
  NAND2_X1 U6028 ( .A1(n8213), .A2(n8212), .ZN(n9047) );
  AND2_X1 U6029 ( .A1(n4693), .A2(n4867), .ZN(n4503) );
  OR2_X1 U6030 ( .A1(n9788), .A2(n9678), .ZN(n4504) );
  AND2_X1 U6031 ( .A1(n8028), .A2(n9490), .ZN(n4505) );
  INV_X1 U6032 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5038) );
  INV_X1 U6033 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4599) );
  AND2_X1 U6034 ( .A1(n9803), .A2(n9732), .ZN(n4506) );
  AND2_X1 U6035 ( .A1(n8754), .A2(n9119), .ZN(n4507) );
  INV_X1 U6036 ( .A(n6024), .ZN(n4638) );
  NAND2_X1 U6037 ( .A1(n8797), .A2(n8796), .ZN(n4508) );
  INV_X1 U6038 ( .A(n7611), .ZN(n5963) );
  AND2_X1 U6039 ( .A1(n8046), .A2(n9487), .ZN(n4509) );
  OR2_X1 U6040 ( .A1(n8596), .A2(n8774), .ZN(n8770) );
  INV_X1 U6041 ( .A(n4765), .ZN(n4764) );
  XNOR2_X1 U6042 ( .A(n6423), .B(n6422), .ZN(n6409) );
  OR2_X1 U6043 ( .A1(n5017), .A2(n6169), .ZN(n4510) );
  OR2_X1 U6044 ( .A1(n9316), .A2(n9176), .ZN(n8735) );
  AND2_X1 U6045 ( .A1(n4900), .A2(n7976), .ZN(n4511) );
  INV_X1 U6046 ( .A(n4554), .ZN(n4553) );
  OAI21_X1 U6047 ( .B1(n9064), .B2(n9029), .A(n9032), .ZN(n4554) );
  NAND2_X1 U6048 ( .A1(n5070), .A2(n5038), .ZN(n4512) );
  AND2_X1 U6049 ( .A1(n5032), .A2(n4940), .ZN(n4513) );
  AND2_X1 U6050 ( .A1(n5237), .A2(SI_7_), .ZN(n4514) );
  NAND2_X1 U6051 ( .A1(n5983), .A2(n5982), .ZN(n4515) );
  INV_X1 U6052 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6854) );
  INV_X1 U6053 ( .A(n10137), .ZN(n7379) );
  AND2_X1 U6054 ( .A1(n5908), .A2(n5907), .ZN(n10137) );
  AND2_X1 U6055 ( .A1(n4992), .A2(n4990), .ZN(n4516) );
  AND2_X1 U6056 ( .A1(n8265), .A2(n4862), .ZN(n4517) );
  AND2_X1 U6057 ( .A1(n8788), .A2(n8780), .ZN(n4518) );
  INV_X1 U6058 ( .A(n9880), .ZN(n9001) );
  AOI21_X1 U6059 ( .B1(n8588), .B2(n8233), .A(n8224), .ZN(n9880) );
  NAND2_X1 U6060 ( .A1(n6155), .A2(n6154), .ZN(n9793) );
  AND2_X1 U6061 ( .A1(n4677), .A2(n4675), .ZN(n4519) );
  NAND2_X1 U6062 ( .A1(n6240), .A2(n6239), .ZN(n9768) );
  NAND2_X1 U6063 ( .A1(n4795), .A2(n5212), .ZN(n5235) );
  NOR2_X1 U6064 ( .A1(n4981), .A2(n4980), .ZN(n4520) );
  NOR2_X1 U6065 ( .A1(n6326), .A2(n4909), .ZN(n4521) );
  NOR2_X1 U6066 ( .A1(n9135), .A2(n8594), .ZN(n4522) );
  NAND2_X1 U6067 ( .A1(n8290), .A2(n8289), .ZN(n4523) );
  AND2_X1 U6068 ( .A1(n4659), .A2(n9713), .ZN(n4524) );
  NOR2_X1 U6069 ( .A1(n8618), .A2(n4555), .ZN(n4525) );
  NAND2_X1 U6070 ( .A1(n9275), .A2(n8608), .ZN(n4526) );
  AND2_X1 U6071 ( .A1(n6402), .A2(n6400), .ZN(n4527) );
  AND2_X1 U6072 ( .A1(n8315), .A2(n8322), .ZN(n8408) );
  AND2_X1 U6073 ( .A1(n8678), .A2(n8679), .ZN(n8675) );
  AND2_X1 U6074 ( .A1(n4737), .A2(n4736), .ZN(n4528) );
  AND2_X1 U6075 ( .A1(n10229), .A2(n7521), .ZN(n4529) );
  AND2_X1 U6076 ( .A1(n5008), .A2(n5007), .ZN(n4530) );
  AND2_X1 U6077 ( .A1(n4485), .A2(n8120), .ZN(n4994) );
  INV_X1 U6078 ( .A(n7557), .ZN(n9496) );
  AND4_X1 U6079 ( .A1(n5876), .A2(n5875), .A3(n5874), .A4(n5873), .ZN(n7557)
         );
  NAND2_X1 U6080 ( .A1(n9711), .A2(n9713), .ZN(n4666) );
  INV_X1 U6081 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4940) );
  XNOR2_X1 U6082 ( .A(n5060), .B(n5059), .ZN(n5702) );
  INV_X1 U6083 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4757) );
  AND2_X1 U6084 ( .A1(n6800), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4531) );
  INV_X1 U6085 ( .A(n8425), .ZN(n4762) );
  NAND2_X1 U6086 ( .A1(n6085), .A2(n6084), .ZN(n8118) );
  INV_X1 U6087 ( .A(n6851), .ZN(n4889) );
  NAND2_X1 U6088 ( .A1(n4881), .A2(n4880), .ZN(n9711) );
  NAND2_X1 U6089 ( .A1(n6392), .A2(n6391), .ZN(n7869) );
  NAND2_X1 U6090 ( .A1(n4882), .A2(n4886), .ZN(n8107) );
  OAI211_X1 U6091 ( .C1(n7976), .C2(n4906), .A(n4905), .B(n4901), .ZN(n8142)
         );
  NAND2_X1 U6092 ( .A1(n5345), .A2(n5344), .ZN(n8704) );
  AND2_X1 U6093 ( .A1(n8556), .A2(n10044), .ZN(n8482) );
  INV_X1 U6094 ( .A(n8482), .ZN(n4545) );
  OR3_X1 U6095 ( .A1(n5694), .A2(n9072), .A3(n8892), .ZN(n4532) );
  INV_X1 U6096 ( .A(n9008), .ZN(n9230) );
  INV_X1 U6097 ( .A(n4704), .ZN(n9735) );
  NOR3_X1 U6098 ( .A1(n4706), .A2(n7872), .A3(n8046), .ZN(n4704) );
  NOR3_X1 U6099 ( .A1(n9235), .A2(n9325), .A3(n4612), .ZN(n4609) );
  AND2_X1 U6100 ( .A1(n8135), .A2(n8134), .ZN(n4533) );
  NAND2_X1 U6101 ( .A1(n9147), .A2(n4606), .ZN(n4534) );
  INV_X1 U6102 ( .A(n4610), .ZN(n9195) );
  NOR2_X1 U6103 ( .A1(n9235), .A2(n4612), .ZN(n4610) );
  AND2_X1 U6104 ( .A1(n4643), .A2(n4641), .ZN(n4535) );
  AND2_X1 U6105 ( .A1(n4470), .A2(n9891), .ZN(n4536) );
  NAND2_X1 U6106 ( .A1(n9325), .A2(n9015), .ZN(n4537) );
  OR2_X1 U6107 ( .A1(n5062), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n4538) );
  NAND2_X1 U6108 ( .A1(n5924), .A2(n5923), .ZN(n4977) );
  AND3_X2 U6109 ( .A1(n6477), .A2(n6930), .A3(n6476), .ZN(n10173) );
  NAND2_X1 U6110 ( .A1(n5327), .A2(n5326), .ZN(n7958) );
  INV_X1 U6111 ( .A(n7958), .ZN(n4614) );
  NAND2_X1 U6112 ( .A1(n5031), .A2(n4729), .ZN(n5663) );
  NOR2_X1 U6113 ( .A1(n7348), .A2(n7547), .ZN(n4687) );
  NAND2_X1 U6114 ( .A1(n4857), .A2(n4856), .ZN(n7352) );
  INV_X1 U6115 ( .A(n9808), .ZN(n4707) );
  NAND2_X1 U6116 ( .A1(n7676), .A2(n8678), .ZN(n7760) );
  NAND2_X1 U6117 ( .A1(n4861), .A2(n6390), .ZN(n7881) );
  INV_X1 U6118 ( .A(n4645), .ZN(n7700) );
  INV_X1 U6119 ( .A(n7663), .ZN(n4937) );
  INV_X1 U6120 ( .A(n8511), .ZN(n4759) );
  NAND2_X1 U6121 ( .A1(n7493), .A2(n7492), .ZN(n7494) );
  OAI211_X1 U6122 ( .C1(n7386), .C2(n4583), .A(n8514), .B(n4586), .ZN(n7371)
         );
  INV_X1 U6123 ( .A(n7371), .ZN(n4585) );
  NAND2_X1 U6124 ( .A1(n4971), .A2(n4488), .ZN(n7608) );
  NAND2_X1 U6125 ( .A1(n4977), .A2(n5940), .ZN(n7536) );
  NAND2_X1 U6126 ( .A1(n5031), .A2(n4786), .ZN(n5661) );
  NAND2_X1 U6127 ( .A1(n7641), .A2(n7640), .ZN(n7643) );
  NAND2_X1 U6128 ( .A1(n5004), .A2(n5005), .ZN(n6292) );
  NOR2_X1 U6129 ( .A1(n4462), .A2(n10218), .ZN(n4539) );
  AND2_X1 U6130 ( .A1(n7446), .A2(n7445), .ZN(n7447) );
  INV_X1 U6131 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4797) );
  INV_X1 U6132 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5779) );
  XNOR2_X1 U6133 ( .A(n5767), .B(n5768), .ZN(n8549) );
  INV_X1 U6134 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5006) );
  INV_X1 U6135 ( .A(n8546), .ZN(n4550) );
  INV_X1 U6136 ( .A(n8598), .ZN(n8651) );
  XNOR2_X1 U6137 ( .A(n5066), .B(n5065), .ZN(n8598) );
  NOR2_X1 U6138 ( .A1(n4624), .A2(n5009), .ZN(n9825) );
  AND2_X1 U6139 ( .A1(n8500), .A2(n6438), .ZN(n8492) );
  INV_X1 U6140 ( .A(n8492), .ZN(n6297) );
  INV_X1 U6141 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n4945) );
  NAND2_X2 U6142 ( .A1(n4455), .A2(n8636), .ZN(n8787) );
  OAI211_X1 U6143 ( .C1(n5163), .C2(n4622), .A(n4542), .B(n5183), .ZN(n4623)
         );
  OR2_X1 U6144 ( .A1(n5162), .A2(n4622), .ZN(n4542) );
  AND2_X1 U6145 ( .A1(n4905), .A2(n4904), .ZN(n4900) );
  OR2_X1 U6146 ( .A1(n5376), .A2(n4906), .ZN(n4899) );
  MUX2_X1 U6147 ( .A(n8382), .B(n8381), .S(n4545), .Z(n8384) );
  NAND2_X1 U6148 ( .A1(n4544), .A2(n4543), .ZN(n8371) );
  INV_X1 U6149 ( .A(n7608), .ZN(n5964) );
  INV_X1 U6150 ( .A(n9468), .ZN(n4655) );
  NAND2_X1 U6151 ( .A1(n8391), .A2(n8390), .ZN(n8395) );
  MUX2_X1 U6152 ( .A(n8480), .B(n8479), .S(n4545), .Z(n8491) );
  NAND2_X1 U6153 ( .A1(n8491), .A2(n8490), .ZN(n4829) );
  NAND2_X1 U6154 ( .A1(n4995), .A2(n4994), .ZN(n4991) );
  NAND2_X1 U6155 ( .A1(n4991), .A2(n4992), .ZN(n6143) );
  OAI21_X1 U6156 ( .B1(n8453), .B2(n8454), .A(n8452), .ZN(n4549) );
  NAND2_X1 U6157 ( .A1(n8473), .A2(n8472), .ZN(n8481) );
  OAI21_X1 U6158 ( .B1(n4829), .B2(n6297), .A(n4523), .ZN(n4828) );
  NAND2_X1 U6159 ( .A1(n4442), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5809) );
  NAND2_X1 U6160 ( .A1(n8101), .A2(n5380), .ZN(n5405) );
  AOI21_X1 U6161 ( .B1(n4655), .B2(n4654), .A(n4656), .ZN(n9444) );
  AND3_X4 U6162 ( .A1(n5815), .A2(n5813), .A3(n5814), .ZN(n10092) );
  NAND2_X1 U6163 ( .A1(n4548), .A2(n4547), .ZN(n8416) );
  NAND2_X1 U6164 ( .A1(n8402), .A2(n8401), .ZN(n4548) );
  NAND3_X2 U6165 ( .A1(n5004), .A2(n5740), .A3(n4468), .ZN(n4624) );
  AND2_X2 U6166 ( .A1(n5738), .A2(n5737), .ZN(n5004) );
  NAND2_X4 U6167 ( .A1(n6301), .A2(n6461), .ZN(n6064) );
  NAND2_X1 U6168 ( .A1(n4549), .A2(n8455), .ZN(n8457) );
  NAND2_X1 U6169 ( .A1(n10048), .A2(n10049), .ZN(n10047) );
  NAND2_X1 U6170 ( .A1(n4828), .A2(n10044), .ZN(n4827) );
  NAND2_X1 U6171 ( .A1(n4827), .A2(n4825), .ZN(n8553) );
  OAI21_X1 U6172 ( .B1(n9386), .B2(n9385), .A(n9467), .ZN(n9390) );
  NAND2_X1 U6173 ( .A1(n4985), .A2(n4983), .ZN(n7723) );
  NOR2_X1 U6174 ( .A1(n9444), .A2(n9445), .ZN(n9443) );
  NAND2_X1 U6175 ( .A1(n6201), .A2(n6200), .ZN(n9451) );
  AOI21_X1 U6176 ( .B1(n8118), .B2(n4994), .A(n4988), .ZN(n9465) );
  NAND2_X1 U6177 ( .A1(n6042), .A2(n4520), .ZN(n4979) );
  NAND2_X1 U6178 ( .A1(n4979), .A2(n4978), .ZN(n8063) );
  OAI21_X2 U6179 ( .B1(n5781), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5767) );
  OAI21_X1 U6180 ( .B1(n9030), .B2(n9064), .A(n4553), .ZN(n9053) );
  INV_X1 U6181 ( .A(n4551), .ZN(n9035) );
  NAND2_X1 U6182 ( .A1(n9030), .A2(n9029), .ZN(n9063) );
  INV_X1 U6183 ( .A(n5031), .ZN(n5064) );
  AND2_X4 U6184 ( .A1(n5324), .A2(n5030), .ZN(n5031) );
  AND3_X2 U6185 ( .A1(n4712), .A2(n5026), .A3(n4898), .ZN(n5047) );
  XNOR2_X1 U6186 ( .A(n8826), .B(n4556), .ZN(n7443) );
  NAND2_X2 U6187 ( .A1(n4720), .A2(n4717), .ZN(n9309) );
  AND2_X2 U6188 ( .A1(n4557), .A2(n4537), .ZN(n9162) );
  XNOR2_X2 U6189 ( .A(n5036), .B(n5035), .ZN(n5043) );
  NAND2_X1 U6190 ( .A1(n7859), .A2(n4566), .ZN(n4564) );
  NAND2_X1 U6191 ( .A1(n4564), .A2(n4565), .ZN(n8008) );
  OAI211_X1 U6192 ( .C1(n5073), .C2(P1_DATAO_REG_3__SCAN_IN), .A(n4570), .B(
        n4569), .ZN(n5141) );
  NAND3_X1 U6193 ( .A1(n5074), .A2(n5073), .A3(n6848), .ZN(n4570) );
  NAND3_X1 U6194 ( .A1(n7646), .A2(n4961), .A3(n7851), .ZN(n4573) );
  XNOR2_X1 U6195 ( .A(n5163), .B(n5162), .ZN(n6853) );
  NAND2_X1 U6196 ( .A1(n9686), .A2(n9685), .ZN(n6454) );
  NAND2_X1 U6197 ( .A1(n7870), .A2(n4481), .ZN(n4590) );
  NAND2_X1 U6198 ( .A1(n6455), .A2(n4595), .ZN(n4594) );
  NAND2_X1 U6199 ( .A1(n4594), .A2(n8293), .ZN(n9588) );
  NAND2_X1 U6200 ( .A1(n4598), .A2(n4596), .ZN(n6456) );
  OAI21_X2 U6201 ( .B1(n4624), .B2(n5011), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4600) );
  NAND2_X2 U6202 ( .A1(n6974), .A2(n8809), .ZN(n5101) );
  INV_X1 U6203 ( .A(n4609), .ZN(n9180) );
  AND2_X1 U6204 ( .A1(n9091), .A2(n4617), .ZN(n9054) );
  NAND2_X1 U6205 ( .A1(n9091), .A2(n4618), .ZN(n9043) );
  NAND2_X1 U6206 ( .A1(n9091), .A2(n9071), .ZN(n9065) );
  NAND2_X1 U6207 ( .A1(n5163), .A2(n5162), .ZN(n4621) );
  INV_X1 U6208 ( .A(n5166), .ZN(n4622) );
  NAND2_X2 U6209 ( .A1(n4624), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U6210 ( .A1(n4629), .A2(n10173), .ZN(n4626) );
  NAND2_X1 U6211 ( .A1(n7352), .A2(n4477), .ZN(n7304) );
  NAND2_X1 U6212 ( .A1(n7869), .A2(n4641), .ZN(n4639) );
  NAND2_X1 U6213 ( .A1(n4639), .A2(n4640), .ZN(n8053) );
  NAND2_X1 U6214 ( .A1(n4789), .A2(n4792), .ZN(n5253) );
  NOR2_X1 U6215 ( .A1(n9463), .A2(n4657), .ZN(n4654) );
  NAND2_X1 U6216 ( .A1(n9711), .A2(n4524), .ZN(n4658) );
  NAND2_X1 U6217 ( .A1(n4658), .A2(n4661), .ZN(n9668) );
  NAND2_X1 U6218 ( .A1(n9208), .A2(n9207), .ZN(n9206) );
  OR2_X1 U6219 ( .A1(n9074), .A2(n9075), .ZN(n4682) );
  NAND2_X1 U6220 ( .A1(n4676), .A2(n4519), .ZN(n4674) );
  INV_X1 U6221 ( .A(n4682), .ZN(n9073) );
  INV_X1 U6222 ( .A(n8772), .ZN(n4681) );
  INV_X1 U6223 ( .A(n4688), .ZN(n9669) );
  INV_X2 U6224 ( .A(n5834), .ZN(n8283) );
  INV_X1 U6225 ( .A(n4697), .ZN(n9596) );
  INV_X1 U6226 ( .A(n7872), .ZN(n4702) );
  NAND2_X1 U6227 ( .A1(n4702), .A2(n4703), .ZN(n9736) );
  NAND2_X1 U6228 ( .A1(n7441), .A2(n7442), .ZN(n7446) );
  INV_X2 U6229 ( .A(n5117), .ZN(n4709) );
  INV_X2 U6230 ( .A(n7037), .ZN(n7619) );
  NAND2_X1 U6231 ( .A1(n4452), .A2(n9846), .ZN(n4710) );
  INV_X1 U6232 ( .A(n5026), .ZN(n5135) );
  NOR2_X2 U6233 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5091) );
  INV_X1 U6234 ( .A(n9018), .ZN(n4723) );
  NAND2_X1 U6235 ( .A1(n7522), .A2(n4529), .ZN(n4725) );
  NAND2_X1 U6236 ( .A1(n7522), .A2(n7521), .ZN(n7562) );
  OR2_X2 U6237 ( .A1(n8007), .A2(n8010), .ZN(n4726) );
  AND2_X2 U6238 ( .A1(n5031), .A2(n4727), .ZN(n5670) );
  NAND3_X1 U6239 ( .A1(n4741), .A2(n4738), .A3(n8709), .ZN(n4737) );
  XNOR2_X1 U6240 ( .A(n5184), .B(n5183), .ZN(n6862) );
  INV_X1 U6241 ( .A(n5074), .ZN(n4755) );
  OAI211_X1 U6242 ( .C1(n5073), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n4756), .B(
        n4754), .ZN(n5113) );
  NAND3_X1 U6243 ( .A1(n6842), .A2(n5073), .A3(n5074), .ZN(n4756) );
  NAND2_X1 U6244 ( .A1(n4760), .A2(n8511), .ZN(n8356) );
  NAND2_X1 U6245 ( .A1(n4769), .A2(n4768), .ZN(n4770) );
  OR2_X1 U6246 ( .A1(n9588), .A2(n9594), .ZN(n9591) );
  NAND2_X1 U6247 ( .A1(n9591), .A2(n8467), .ZN(n9572) );
  OAI21_X1 U6248 ( .B1(n8613), .B2(n4778), .A(n7442), .ZN(n10227) );
  NAND2_X1 U6249 ( .A1(n7923), .A2(n7922), .ZN(n7961) );
  AND2_X2 U6250 ( .A1(n7921), .A2(n7920), .ZN(n7923) );
  NAND2_X2 U6251 ( .A1(n5101), .A2(n4445), .ZN(n5117) );
  NAND2_X1 U6252 ( .A1(n9309), .A2(n4781), .ZN(n9111) );
  NAND2_X1 U6253 ( .A1(n5031), .A2(n4784), .ZN(n5037) );
  NAND2_X1 U6254 ( .A1(n7447), .A2(n7455), .ZN(n7493) );
  NAND2_X1 U6255 ( .A1(n9111), .A2(n9024), .ZN(n9096) );
  NAND2_X1 U6256 ( .A1(n5189), .A2(n4790), .ZN(n4789) );
  NAND2_X2 U6257 ( .A1(n4796), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5073) );
  NAND2_X1 U6258 ( .A1(n4797), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4796) );
  NAND2_X1 U6259 ( .A1(n4798), .A2(n4800), .ZN(n5518) );
  NAND2_X1 U6260 ( .A1(n5472), .A2(n4802), .ZN(n4798) );
  NAND2_X1 U6261 ( .A1(n5472), .A2(n5471), .ZN(n4807) );
  INV_X1 U6262 ( .A(n4808), .ZN(n5454) );
  NAND2_X1 U6263 ( .A1(n5255), .A2(n4819), .ZN(n4818) );
  NAND2_X1 U6264 ( .A1(n4818), .A2(n4822), .ZN(n5295) );
  OR2_X1 U6265 ( .A1(n5337), .A2(n5338), .ZN(n4831) );
  NAND2_X1 U6266 ( .A1(n4830), .A2(n4832), .ZN(n5361) );
  NAND2_X1 U6267 ( .A1(n5337), .A2(n5339), .ZN(n4830) );
  NAND3_X1 U6268 ( .A1(n4852), .A2(n4851), .A3(n4849), .ZN(P1_U3260) );
  NAND3_X1 U6269 ( .A1(n9496), .A2(n6382), .A3(n7367), .ZN(n4855) );
  NAND2_X1 U6270 ( .A1(n7784), .A2(n4517), .ZN(n4858) );
  NAND2_X1 U6271 ( .A1(n4858), .A2(n4860), .ZN(n7803) );
  NAND2_X1 U6272 ( .A1(n9728), .A2(n4469), .ZN(n4881) );
  NAND2_X1 U6273 ( .A1(n6399), .A2(n4892), .ZN(n4891) );
  NAND2_X1 U6274 ( .A1(n4891), .A2(n4527), .ZN(n6404) );
  NAND3_X1 U6275 ( .A1(n5074), .A2(n5073), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n4894) );
  NAND3_X1 U6276 ( .A1(n5074), .A2(n5073), .A3(n5076), .ZN(n5795) );
  XNOR2_X1 U6277 ( .A(n5096), .B(n5078), .ZN(n5095) );
  NAND2_X1 U6278 ( .A1(n7157), .A2(n4897), .ZN(n7156) );
  XNOR2_X1 U6279 ( .A(n5083), .B(n5085), .ZN(n4897) );
  OAI21_X1 U6280 ( .B1(n7157), .B2(n4897), .A(n7156), .ZN(n7162) );
  NAND2_X1 U6281 ( .A1(n7976), .A2(n5376), .ZN(n8101) );
  NAND2_X1 U6282 ( .A1(n8811), .A2(n5590), .ZN(n4918) );
  NAND2_X1 U6283 ( .A1(n8811), .A2(n4521), .ZN(n4908) );
  AND2_X1 U6284 ( .A1(n5593), .A2(n5594), .ZN(n4920) );
  INV_X1 U6285 ( .A(n7206), .ZN(n4924) );
  NAND3_X1 U6286 ( .A1(n4922), .A2(n8818), .A3(n4921), .ZN(n7214) );
  NAND2_X1 U6287 ( .A1(n7206), .A2(n5105), .ZN(n4922) );
  NAND2_X1 U6288 ( .A1(n7666), .A2(n4930), .ZN(n4927) );
  NAND2_X1 U6289 ( .A1(n4927), .A2(n4928), .ZN(n7900) );
  AOI21_X1 U6290 ( .B1(n4930), .B2(n4934), .A(n4492), .ZN(n4928) );
  INV_X1 U6291 ( .A(n4934), .ZN(n4933) );
  NOR2_X1 U6292 ( .A1(n7716), .A2(n4937), .ZN(n4936) );
  NAND2_X1 U6293 ( .A1(n8881), .A2(n5195), .ZN(n8880) );
  NAND2_X1 U6294 ( .A1(n5429), .A2(n4939), .ZN(n6763) );
  NAND2_X1 U6295 ( .A1(n6763), .A2(n5448), .ZN(n5469) );
  XNOR2_X2 U6296 ( .A(n5069), .B(n5068), .ZN(n6974) );
  INV_X1 U6297 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n4942) );
  INV_X1 U6298 ( .A(n4944), .ZN(n4943) );
  OAI22_X1 U6299 ( .A1(n5130), .A2(n4945), .B1(n7470), .B2(n4453), .ZN(n4944)
         );
  NAND2_X1 U6300 ( .A1(n4948), .A2(n9135), .ZN(n4947) );
  NAND3_X1 U6301 ( .A1(n4947), .A2(n4946), .A3(n8762), .ZN(n9074) );
  NAND2_X1 U6302 ( .A1(n8008), .A2(n8709), .ZN(n4963) );
  NAND3_X1 U6303 ( .A1(n4966), .A2(n4518), .A3(n4965), .ZN(n4964) );
  NAND2_X1 U6304 ( .A1(n8604), .A2(n8782), .ZN(n4965) );
  OAI21_X1 U6305 ( .B1(n8604), .B2(n9001), .A(n8607), .ZN(n4966) );
  INV_X1 U6306 ( .A(n10098), .ZN(n4969) );
  NAND2_X1 U6307 ( .A1(n5924), .A2(n4972), .ZN(n4971) );
  NAND2_X1 U6308 ( .A1(n5964), .A2(n4986), .ZN(n4985) );
  NAND2_X1 U6309 ( .A1(n6104), .A2(n6103), .ZN(n4995) );
  NAND2_X1 U6310 ( .A1(n6275), .A2(n4997), .ZN(n4996) );
  OAI211_X1 U6311 ( .C1(n6275), .C2(n5001), .A(n4998), .B(n4996), .ZN(n8210)
         );
  INV_X1 U6312 ( .A(n9756), .ZN(n9598) );
  NAND2_X1 U6313 ( .A1(n5695), .A2(n4532), .ZN(n5701) );
  NAND2_X1 U6314 ( .A1(n7444), .A2(n7443), .ZN(n7445) );
  OAI21_X2 U6315 ( .B1(n5454), .B2(n5453), .A(n5452), .ZN(n5472) );
  NAND2_X1 U6316 ( .A1(n7275), .A2(n7268), .ZN(n8661) );
  XNOR2_X1 U6317 ( .A(n9053), .B(n9052), .ZN(n9288) );
  NAND2_X2 U6318 ( .A1(n7977), .A2(n7978), .ZN(n7976) );
  INV_X1 U6319 ( .A(n7010), .ZN(n7013) );
  NAND2_X1 U6320 ( .A1(n6444), .A2(n8503), .ZN(n7254) );
  CLKBUF_X1 U6321 ( .A(n7288), .Z(n8506) );
  INV_X1 U6322 ( .A(n5871), .ZN(n5884) );
  NAND2_X1 U6323 ( .A1(n5037), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5039) );
  NAND2_X2 U6324 ( .A1(n9417), .A2(n9418), .ZN(n6275) );
  CLKBUF_X2 U6325 ( .A(n6375), .Z(n9499) );
  OAI21_X2 U6326 ( .B1(n5601), .B2(n5600), .A(n5599), .ZN(n5619) );
  OR2_X1 U6327 ( .A1(n6321), .A2(n6320), .ZN(n5013) );
  NAND2_X1 U6328 ( .A1(n6440), .A2(n6439), .ZN(n10050) );
  AND2_X1 U6329 ( .A1(n8702), .A2(n8701), .ZN(n8626) );
  AND2_X1 U6330 ( .A1(n6788), .A2(n8492), .ZN(n10045) );
  INV_X1 U6331 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5067) );
  OR2_X1 U6332 ( .A1(n8789), .A2(n8793), .ZN(n5014) );
  NOR2_X1 U6333 ( .A1(n8164), .A2(n8628), .ZN(n5015) );
  AND2_X1 U6334 ( .A1(n6186), .A2(n6185), .ZN(n5017) );
  OR2_X1 U6335 ( .A1(n8211), .A2(n8856), .ZN(n5018) );
  AND2_X1 U6336 ( .A1(n8556), .A2(n8500), .ZN(n5019) );
  AND4_X1 U6337 ( .A1(n5554), .A2(n5553), .A3(n5552), .A4(n5551), .ZN(n9176)
         );
  AND2_X1 U6338 ( .A1(n5294), .A2(n5271), .ZN(n5020) );
  AND2_X1 U6339 ( .A1(n5268), .A2(n5259), .ZN(n5021) );
  AND3_X1 U6340 ( .A1(n5588), .A2(n5587), .A3(n5586), .ZN(n9021) );
  AND2_X1 U6341 ( .A1(n5715), .A2(n5714), .ZN(n8774) );
  AND2_X1 U6342 ( .A1(n8548), .A2(n10044), .ZN(n5022) );
  NAND2_X1 U6343 ( .A1(n8053), .A2(n8271), .ZN(n8052) );
  AND4_X1 U6344 ( .A1(n5529), .A2(n5528), .A3(n5527), .A4(n5526), .ZN(n9016)
         );
  INV_X1 U6345 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5740) );
  OAI21_X1 U6346 ( .B1(n9676), .B2(n8433), .A(n8446), .ZN(n9660) );
  XNOR2_X1 U6347 ( .A(n5827), .B(n5828), .ZN(n7009) );
  AND3_X1 U6348 ( .A1(n6344), .A2(n6345), .A3(n8882), .ZN(n5024) );
  INV_X1 U6349 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5729) );
  AND2_X1 U6350 ( .A1(n4526), .A2(n8782), .ZN(n8783) );
  INV_X1 U6351 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5049) );
  INV_X1 U6352 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5741) );
  OR2_X1 U6353 ( .A1(n5593), .A2(n9136), .ZN(n5589) );
  INV_X1 U6354 ( .A(n7455), .ZN(n7456) );
  AND2_X1 U6355 ( .A1(n5589), .A2(n8810), .ZN(n5590) );
  INV_X1 U6356 ( .A(n5585), .ZN(n5575) );
  OR2_X1 U6357 ( .A1(n5626), .A2(n5625), .ZN(n5649) );
  OR2_X1 U6358 ( .A1(n5583), .A2(n8813), .ZN(n5585) );
  INV_X1 U6359 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5347) );
  INV_X1 U6360 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5053) );
  INV_X1 U6361 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5989) );
  AND2_X1 U6362 ( .A1(n6189), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6205) );
  NOR2_X1 U6363 ( .A1(n6716), .A2(n6048), .ZN(n6068) );
  INV_X1 U6364 ( .A(n8359), .ZN(n6384) );
  INV_X1 U6365 ( .A(n5470), .ZN(n5471) );
  INV_X1 U6366 ( .A(SI_13_), .ZN(n6594) );
  INV_X1 U6367 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5296) );
  INV_X1 U6368 ( .A(SI_8_), .ZN(n6606) );
  INV_X1 U6369 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5348) );
  INV_X1 U6370 ( .A(n5419), .ZN(n5418) );
  OR2_X1 U6371 ( .A1(n5548), .A2(n8862), .ZN(n5583) );
  INV_X1 U6372 ( .A(n6813), .ZN(n5174) );
  OR2_X1 U6373 ( .A1(n5709), .A2(n6348), .ZN(n9045) );
  NAND2_X1 U6374 ( .A1(n5368), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6375 ( .A1(n5204), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5089) );
  AND2_X1 U6376 ( .A1(n7051), .A2(n7050), .ZN(n7053) );
  INV_X1 U6377 ( .A(n9021), .ZN(n9022) );
  INV_X1 U6378 ( .A(n8626), .ZN(n7922) );
  INV_X1 U6379 ( .A(n6059), .ZN(n6060) );
  AND2_X1 U6380 ( .A1(n9382), .A2(n9383), .ZN(n8197) );
  INV_X1 U6381 ( .A(n7722), .ZN(n6000) );
  NOR2_X1 U6382 ( .A1(n5990), .A2(n5989), .ZN(n6011) );
  INV_X1 U6383 ( .A(n6241), .ZN(n6242) );
  NOR2_X1 U6384 ( .A1(n6148), .A2(n9404), .ZN(n6157) );
  NAND2_X1 U6385 ( .A1(n6133), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6148) );
  OR2_X1 U6386 ( .A1(n5971), .A2(n7066), .ZN(n5990) );
  AND2_X1 U6387 ( .A1(n6280), .A2(n6277), .ZN(n5761) );
  OR2_X1 U6388 ( .A1(n6089), .A2(n6088), .ZN(n6109) );
  NAND2_X1 U6389 ( .A1(n5418), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5459) );
  INV_X1 U6390 ( .A(n7436), .ZN(n7268) );
  INV_X1 U6391 ( .A(n5129), .ZN(n6353) );
  OR2_X1 U6392 ( .A1(n4454), .A2(n7618), .ZN(n6950) );
  INV_X1 U6393 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8926) );
  INV_X1 U6394 ( .A(n10200), .ZN(n6894) );
  NOR2_X1 U6395 ( .A1(n9336), .A2(n9008), .ZN(n9009) );
  AND2_X1 U6396 ( .A1(n8800), .A2(n8651), .ZN(n6972) );
  OR2_X1 U6397 ( .A1(n7853), .A2(n7851), .ZN(n7755) );
  INV_X1 U6398 ( .A(n10198), .ZN(n9244) );
  AND2_X1 U6399 ( .A1(n8610), .A2(n8793), .ZN(n9228) );
  INV_X1 U6400 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7066) );
  OR2_X1 U6401 ( .A1(n6308), .A2(n9615), .ZN(n6262) );
  NAND2_X1 U6402 ( .A1(n8285), .A2(n8284), .ZN(n8286) );
  INV_X1 U6403 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U6404 ( .A1(n6377), .A2(n6376), .ZN(n7287) );
  AND2_X1 U6405 ( .A1(n8492), .A2(n8546), .ZN(n6925) );
  AND2_X1 U6406 ( .A1(n8251), .A2(n8250), .ZN(n9729) );
  INV_X1 U6407 ( .A(n10046), .ZN(n9716) );
  AND2_X1 U6408 ( .A1(n5571), .A2(n5565), .ZN(n5569) );
  AND2_X1 U6409 ( .A1(n5432), .A2(n5413), .ZN(n5430) );
  OAI21_X1 U6410 ( .B1(n9071), .B2(n8856), .A(n5721), .ZN(n5722) );
  NAND2_X1 U6411 ( .A1(n6358), .A2(n6357), .ZN(n6359) );
  NAND2_X2 U6412 ( .A1(n6894), .A2(n7019), .ZN(n9241) );
  AND2_X1 U6413 ( .A1(n10272), .A2(n5691), .ZN(n5692) );
  INV_X1 U6414 ( .A(n8868), .ZN(n8882) );
  INV_X1 U6415 ( .A(n8856), .ZN(n8890) );
  INV_X1 U6416 ( .A(n4459), .ZN(n8603) );
  AND4_X1 U6417 ( .A1(n5442), .A2(n5441), .A3(n5440), .A4(n5439), .ZN(n8874)
         );
  AND4_X1 U6418 ( .A1(n5331), .A2(n5330), .A3(n5329), .A4(n5328), .ZN(n7980)
         );
  AND2_X1 U6419 ( .A1(n7003), .A2(n7002), .ZN(n10174) );
  AND2_X1 U6420 ( .A1(n6976), .A2(n8809), .ZN(n9860) );
  AND2_X1 U6421 ( .A1(n5718), .A2(n6972), .ZN(n9264) );
  NAND2_X1 U6422 ( .A1(n7430), .A2(n9241), .ZN(n9238) );
  OR2_X1 U6423 ( .A1(n7420), .A2(n7019), .ZN(n7128) );
  AND2_X1 U6424 ( .A1(n4462), .A2(n8794), .ZN(n10231) );
  NAND2_X1 U6425 ( .A1(n8799), .A2(n8794), .ZN(n10272) );
  INV_X1 U6426 ( .A(n10278), .ZN(n10235) );
  NAND2_X1 U6427 ( .A1(n8170), .A2(n10245), .ZN(n10278) );
  NOR2_X1 U6428 ( .A1(n5673), .A2(n8182), .ZN(n10199) );
  AND2_X1 U6429 ( .A1(n5275), .A2(n5297), .ZN(n6999) );
  XNOR2_X1 U6430 ( .A(n8204), .B(n8203), .ZN(n8205) );
  AND2_X1 U6431 ( .A1(n8551), .A2(n8550), .ZN(n8552) );
  AND4_X1 U6432 ( .A1(n6246), .A2(n6245), .A3(n6244), .A4(n6243), .ZN(n9438)
         );
  AND4_X1 U6433 ( .A1(n6152), .A2(n6151), .A3(n6150), .A4(n6149), .ZN(n9708)
         );
  INV_X1 U6434 ( .A(n10012), .ZN(n9525) );
  INV_X1 U6435 ( .A(n9969), .ZN(n10010) );
  AND2_X1 U6436 ( .A1(n8444), .A2(n9630), .ZN(n9640) );
  INV_X1 U6437 ( .A(n9724), .ZN(n9739) );
  OR2_X1 U6438 ( .A1(n10173), .A2(n6431), .ZN(n6478) );
  OR2_X1 U6439 ( .A1(n10089), .A2(n6473), .ZN(n6477) );
  INV_X1 U6440 ( .A(n10154), .ZN(n10124) );
  AND2_X1 U6441 ( .A1(n10128), .A2(n10106), .ZN(n10141) );
  AND2_X1 U6442 ( .A1(n8482), .A2(n8549), .ZN(n10133) );
  AND2_X1 U6443 ( .A1(n7990), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6295) );
  NOR2_X1 U6444 ( .A1(n5948), .A2(n5947), .ZN(n7071) );
  NOR2_X1 U6445 ( .A1(n10323), .A2(n7831), .ZN(n7832) );
  AND2_X1 U6446 ( .A1(n5686), .A2(n5685), .ZN(n6970) );
  AND2_X1 U6447 ( .A1(n5703), .A2(n9241), .ZN(n8856) );
  NAND2_X1 U6448 ( .A1(n5717), .A2(n5692), .ZN(n8868) );
  NAND2_X1 U6449 ( .A1(n6372), .A2(n6371), .ZN(n6373) );
  INV_X1 U6450 ( .A(n8774), .ZN(n9078) );
  INV_X1 U6451 ( .A(n9016), .ZN(n9187) );
  INV_X1 U6452 ( .A(n9860), .ZN(n10178) );
  INV_X1 U6453 ( .A(n9246), .ZN(n9260) );
  NAND2_X1 U6454 ( .A1(n9238), .A2(n10196), .ZN(n9274) );
  INV_X1 U6455 ( .A(n10281), .ZN(n10279) );
  NOR2_X1 U6456 ( .A1(n10200), .A2(n10199), .ZN(n10210) );
  INV_X1 U6457 ( .A(n10210), .ZN(n10213) );
  INV_X1 U6458 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7987) );
  INV_X1 U6459 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7325) );
  INV_X1 U6460 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6866) );
  INV_X1 U6461 ( .A(n10039), .ZN(n7295) );
  NAND3_X1 U6462 ( .A1(n6297), .A2(n6296), .A3(n10136), .ZN(n9461) );
  NOR2_X1 U6463 ( .A1(n6322), .A2(n5013), .ZN(n6323) );
  INV_X1 U6464 ( .A(n9456), .ZN(n9677) );
  INV_X1 U6465 ( .A(n7612), .ZN(n10022) );
  CLKBUF_X2 U6466 ( .A(P1_U4006), .Z(n9494) );
  OR2_X1 U6467 ( .A1(P1_U3083), .A2(n6808), .ZN(n9999) );
  NAND2_X1 U6468 ( .A1(n10057), .A2(n10042), .ZN(n9724) );
  NAND2_X1 U6469 ( .A1(n10057), .A2(n10027), .ZN(n9746) );
  NAND2_X1 U6470 ( .A1(n7376), .A2(n10036), .ZN(n10057) );
  INV_X1 U6471 ( .A(n10173), .ZN(n10171) );
  INV_X1 U6472 ( .A(n10160), .ZN(n10158) );
  INV_X1 U6473 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8156) );
  INV_X1 U6474 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7732) );
  INV_X1 U6475 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7327) );
  INV_X1 U6476 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6907) );
  NOR2_X1 U6477 ( .A1(n10333), .A2(n10332), .ZN(n10331) );
  NOR2_X1 U6478 ( .A1(n10321), .A2(n10320), .ZN(n10319) );
  AND2_X1 U6479 ( .A1(n6970), .A2(n10216), .ZN(P2_U3966) );
  INV_X2 U6480 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U6481 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5027) );
  NAND4_X1 U6482 ( .A1(n5027), .A2(n5362), .A3(n5048), .A4(n5055), .ZN(n5029)
         );
  NAND4_X1 U6483 ( .A1(n5053), .A2(n5057), .A3(n5391), .A4(n5059), .ZN(n5028)
         );
  NOR2_X1 U6484 ( .A1(n5029), .A2(n5028), .ZN(n5030) );
  INV_X1 U6485 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7625) );
  INV_X1 U6486 ( .A(n6949), .ZN(n5041) );
  NAND2_X1 U6487 ( .A1(n5128), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6951) );
  INV_X1 U6488 ( .A(n6951), .ZN(n5040) );
  NOR2_X1 U6489 ( .A1(n5041), .A2(n5040), .ZN(n5046) );
  BUF_X2 U6490 ( .A(n5043), .Z(n8807) );
  NAND2_X1 U6491 ( .A1(n4460), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6952) );
  INV_X1 U6492 ( .A(n5043), .ZN(n5045) );
  INV_X1 U6493 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7618) );
  BUF_X1 U6494 ( .A(n5047), .Z(n5324) );
  NAND2_X1 U6495 ( .A1(n5047), .A2(n5048), .ZN(n5343) );
  NAND2_X1 U6496 ( .A1(n5391), .A2(n5049), .ZN(n5050) );
  NOR2_X2 U6497 ( .A1(n5414), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U6498 ( .A1(n5434), .A2(n5053), .ZN(n5054) );
  NAND2_X1 U6499 ( .A1(n5455), .A2(n5055), .ZN(n5056) );
  NAND2_X1 U6500 ( .A1(n5061), .A2(n5057), .ZN(n5058) );
  INV_X2 U6501 ( .A(n5479), .ZN(n7032) );
  NAND2_X1 U6502 ( .A1(n5702), .A2(n7032), .ZN(n8799) );
  NAND2_X1 U6503 ( .A1(n5062), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5063) );
  NAND2_X1 U6504 ( .A1(n5064), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5066) );
  INV_X1 U6505 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5065) );
  OR2_X4 U6506 ( .A1(n8799), .A2(n10218), .ZN(n8611) );
  NAND2_X1 U6507 ( .A1(n7025), .A2(n4446), .ZN(n5085) );
  OR2_X2 U6508 ( .A1(n5670), .A2(n9374), .ZN(n5069) );
  NAND2_X1 U6509 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5071) );
  XNOR2_X1 U6510 ( .A(n5071), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9846) );
  INV_X1 U6511 ( .A(n9846), .ZN(n6843) );
  AND2_X1 U6512 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5076) );
  NAND3_X1 U6513 ( .A1(n5075), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n5077) );
  INV_X1 U6514 ( .A(SI_1_), .ZN(n5078) );
  XNOR2_X1 U6515 ( .A(n5094), .B(n5095), .ZN(n6844) );
  INV_X1 U6516 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6845) );
  NAND2_X1 U6517 ( .A1(n4462), .A2(n8651), .ZN(n7422) );
  NAND2_X1 U6518 ( .A1(n5479), .A2(n8800), .ZN(n8793) );
  NAND3_X1 U6519 ( .A1(n8793), .A2(n8598), .A3(n10218), .ZN(n5079) );
  XNOR2_X1 U6520 ( .A(n7037), .B(n4443), .ZN(n5083) );
  INV_X1 U6521 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7470) );
  NAND2_X1 U6522 ( .A1(n5128), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U6523 ( .A1(n8228), .A2(SI_0_), .ZN(n5081) );
  XNOR2_X1 U6524 ( .A(n5081), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9381) );
  MUX2_X1 U6525 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9381), .S(n7001), .Z(n7469) );
  NAND2_X1 U6526 ( .A1(n6954), .A2(n7469), .ZN(n7027) );
  INV_X1 U6527 ( .A(n7027), .ZN(n7030) );
  NAND2_X1 U6528 ( .A1(n7030), .A2(n8611), .ZN(n6955) );
  OR2_X1 U6529 ( .A1(n7469), .A2(n4443), .ZN(n5082) );
  AND2_X1 U6530 ( .A1(n6955), .A2(n5082), .ZN(n7157) );
  INV_X1 U6531 ( .A(n5083), .ZN(n5084) );
  NAND2_X1 U6532 ( .A1(n5085), .A2(n5084), .ZN(n5086) );
  NAND2_X1 U6533 ( .A1(n7156), .A2(n5086), .ZN(n7206) );
  NAND2_X1 U6534 ( .A1(n4459), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5090) );
  INV_X1 U6535 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7434) );
  OR2_X1 U6536 ( .A1(n5129), .A2(n7434), .ZN(n5088) );
  INV_X1 U6537 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7429) );
  NOR2_X1 U6538 ( .A1(n8822), .A2(n6340), .ZN(n5102) );
  INV_X1 U6539 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9374) );
  OR2_X1 U6540 ( .A1(n5091), .A2(n9374), .ZN(n5093) );
  INV_X1 U6541 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5092) );
  NAND2_X1 U6542 ( .A1(n5093), .A2(n5092), .ZN(n5118) );
  OAI21_X1 U6543 ( .B1(n5093), .B2(n5092), .A(n5118), .ZN(n6982) );
  NAND2_X1 U6544 ( .A1(n5096), .A2(SI_1_), .ZN(n5097) );
  NAND2_X1 U6545 ( .A1(n5098), .A2(n5097), .ZN(n5112) );
  INV_X1 U6546 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6842) );
  XNOR2_X1 U6547 ( .A(n5113), .B(SI_2_), .ZN(n5111) );
  XNOR2_X1 U6548 ( .A(n5112), .B(n5111), .ZN(n6846) );
  OR2_X1 U6549 ( .A1(n5110), .A2(n6846), .ZN(n5100) );
  OR2_X1 U6550 ( .A1(n5117), .A2(n4757), .ZN(n5099) );
  OAI211_X1 U6551 ( .C1(n7001), .C2(n6982), .A(n5100), .B(n5099), .ZN(n7436)
         );
  XNOR2_X1 U6552 ( .A(n7436), .B(n4443), .ZN(n8821) );
  OR2_X1 U6553 ( .A1(n5102), .A2(n8821), .ZN(n5103) );
  NAND2_X1 U6554 ( .A1(n5102), .A2(n8821), .ZN(n5105) );
  NAND2_X1 U6555 ( .A1(n4458), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5109) );
  OR2_X1 U6556 ( .A1(n5129), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U6557 ( .A1(n4461), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5107) );
  NAND2_X1 U6558 ( .A1(n8599), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5106) );
  AND2_X1 U6559 ( .A1(n8912), .A2(n8611), .ZN(n5124) );
  NAND2_X1 U6560 ( .A1(n5112), .A2(n5111), .ZN(n5116) );
  INV_X1 U6561 ( .A(n5113), .ZN(n5114) );
  NAND2_X1 U6562 ( .A1(n5114), .A2(SI_2_), .ZN(n5115) );
  NAND2_X1 U6563 ( .A1(n5116), .A2(n5115), .ZN(n5140) );
  INV_X1 U6564 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6850) );
  XNOR2_X1 U6565 ( .A(n5140), .B(n5139), .ZN(n6849) );
  OR2_X1 U6566 ( .A1(n5110), .A2(n6849), .ZN(n5123) );
  OR2_X1 U6567 ( .A1(n5117), .A2(n6850), .ZN(n5122) );
  NAND2_X1 U6568 ( .A1(n5118), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5120) );
  INV_X1 U6569 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5119) );
  XNOR2_X1 U6570 ( .A(n5120), .B(n5119), .ZN(n7118) );
  OR2_X1 U6571 ( .A1(n7001), .A2(n7118), .ZN(n5121) );
  XNOR2_X1 U6573 ( .A(n8826), .B(n5547), .ZN(n7217) );
  NAND2_X1 U6574 ( .A1(n5124), .A2(n7217), .ZN(n5147) );
  INV_X1 U6575 ( .A(n7217), .ZN(n5126) );
  INV_X1 U6576 ( .A(n5124), .ZN(n5125) );
  NAND2_X1 U6577 ( .A1(n5126), .A2(n5125), .ZN(n5127) );
  AND2_X1 U6578 ( .A1(n5147), .A2(n5127), .ZN(n8818) );
  NAND2_X1 U6579 ( .A1(n4458), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5134) );
  INV_X1 U6580 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6984) );
  OR2_X1 U6581 ( .A1(n5522), .A2(n6984), .ZN(n5133) );
  NAND2_X1 U6582 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5155) );
  OAI21_X1 U6583 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n5155), .ZN(n7599) );
  OR2_X1 U6584 ( .A1(n5129), .A2(n7599), .ZN(n5132) );
  INV_X1 U6585 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7596) );
  OR2_X1 U6586 ( .A1(n6888), .A2(n7596), .ZN(n5131) );
  NAND2_X1 U6587 ( .A1(n8911), .A2(n8611), .ZN(n5151) );
  NAND2_X1 U6588 ( .A1(n5135), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5136) );
  MUX2_X1 U6589 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5136), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5138) );
  NAND2_X1 U6590 ( .A1(n5138), .A2(n5137), .ZN(n7103) );
  NAND2_X1 U6591 ( .A1(n5140), .A2(n5139), .ZN(n5144) );
  INV_X1 U6592 ( .A(n5141), .ZN(n5142) );
  NAND2_X1 U6593 ( .A1(n5142), .A2(SI_3_), .ZN(n5143) );
  XNOR2_X1 U6594 ( .A(n5164), .B(SI_4_), .ZN(n5162) );
  OR2_X1 U6595 ( .A1(n5117), .A2(n6854), .ZN(n5145) );
  OAI211_X1 U6596 ( .C1(n7001), .C2(n7103), .A(n5146), .B(n5145), .ZN(n7460)
         );
  XNOR2_X1 U6597 ( .A(n7460), .B(n5169), .ZN(n5149) );
  XNOR2_X1 U6598 ( .A(n5151), .B(n5149), .ZN(n7216) );
  AND2_X1 U6599 ( .A1(n7216), .A2(n5147), .ZN(n5148) );
  NAND2_X1 U6600 ( .A1(n7214), .A2(n5148), .ZN(n7215) );
  INV_X1 U6601 ( .A(n5149), .ZN(n5150) );
  NAND2_X1 U6602 ( .A1(n5151), .A2(n5150), .ZN(n5152) );
  NAND2_X1 U6603 ( .A1(n4459), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5160) );
  INV_X1 U6604 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6988) );
  OR2_X1 U6605 ( .A1(n5522), .A2(n6988), .ZN(n5159) );
  INV_X1 U6606 ( .A(n5155), .ZN(n5153) );
  NAND2_X1 U6607 ( .A1(n5153), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5177) );
  INV_X1 U6608 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U6609 ( .A1(n5155), .A2(n5154), .ZN(n5156) );
  NAND2_X1 U6610 ( .A1(n5177), .A2(n5156), .ZN(n10186) );
  OR2_X1 U6611 ( .A1(n5129), .A2(n10186), .ZN(n5158) );
  INV_X1 U6612 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6959) );
  OR2_X1 U6613 ( .A1(n6888), .A2(n6959), .ZN(n5157) );
  NOR2_X1 U6614 ( .A1(n7565), .A2(n6340), .ZN(n5170) );
  NAND2_X1 U6615 ( .A1(n5137), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5161) );
  XNOR2_X1 U6616 ( .A(n5161), .B(P2_IR_REG_5__SCAN_IN), .ZN(n8918) );
  INV_X1 U6617 ( .A(n8918), .ZN(n6987) );
  INV_X1 U6618 ( .A(n5164), .ZN(n5165) );
  NAND2_X1 U6619 ( .A1(n5165), .A2(SI_4_), .ZN(n5166) );
  MUX2_X1 U6620 ( .A(n6863), .B(n6861), .S(n4444), .Z(n5185) );
  XNOR2_X1 U6621 ( .A(n5185), .B(SI_5_), .ZN(n5183) );
  OR2_X1 U6622 ( .A1(n5117), .A2(n6863), .ZN(n5167) );
  OAI211_X1 U6623 ( .C1(n7001), .C2(n6987), .A(n5168), .B(n5167), .ZN(n10187)
         );
  XNOR2_X1 U6624 ( .A(n10187), .B(n5169), .ZN(n5171) );
  NAND2_X1 U6625 ( .A1(n5170), .A2(n5171), .ZN(n5194) );
  INV_X1 U6626 ( .A(n5170), .ZN(n5172) );
  INV_X1 U6627 ( .A(n5171), .ZN(n8891) );
  NAND2_X1 U6628 ( .A1(n5172), .A2(n8891), .ZN(n5173) );
  NAND2_X1 U6629 ( .A1(n5194), .A2(n5173), .ZN(n6813) );
  NAND2_X1 U6630 ( .A1(n4459), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5182) );
  INV_X1 U6631 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6989) );
  OR2_X1 U6632 ( .A1(n5522), .A2(n6989), .ZN(n5181) );
  INV_X1 U6633 ( .A(n5177), .ZN(n5175) );
  NAND2_X1 U6634 ( .A1(n5175), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5202) );
  INV_X1 U6635 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U6636 ( .A1(n5177), .A2(n5176), .ZN(n5178) );
  NAND2_X1 U6637 ( .A1(n5202), .A2(n5178), .ZN(n8884) );
  OR2_X1 U6638 ( .A1(n5129), .A2(n8884), .ZN(n5180) );
  INV_X1 U6639 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7568) );
  OR2_X1 U6640 ( .A1(n6888), .A2(n7568), .ZN(n5179) );
  NAND2_X1 U6641 ( .A1(n8909), .A2(n8611), .ZN(n5198) );
  INV_X1 U6642 ( .A(n5185), .ZN(n5186) );
  NAND2_X1 U6643 ( .A1(n5186), .A2(SI_5_), .ZN(n5187) );
  INV_X1 U6644 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5188) );
  MUX2_X1 U6645 ( .A(n6866), .B(n5188), .S(n4444), .Z(n5210) );
  XNOR2_X1 U6646 ( .A(n5210), .B(SI_6_), .ZN(n5209) );
  XNOR2_X1 U6647 ( .A(n5189), .B(n5209), .ZN(n6865) );
  OR2_X1 U6648 ( .A1(n8234), .A2(n6866), .ZN(n5193) );
  OR2_X1 U6649 ( .A1(n5190), .A2(n9374), .ZN(n5191) );
  XNOR2_X1 U6650 ( .A(n5191), .B(n5213), .ZN(n7089) );
  OR2_X1 U6651 ( .A1(n7001), .A2(n7089), .ZN(n5192) );
  XNOR2_X1 U6652 ( .A(n7571), .B(n5547), .ZN(n5196) );
  XNOR2_X1 U6653 ( .A(n5198), .B(n5196), .ZN(n8893) );
  AND2_X1 U6654 ( .A1(n8893), .A2(n5194), .ZN(n5195) );
  INV_X1 U6655 ( .A(n5196), .ZN(n5197) );
  NAND2_X1 U6656 ( .A1(n5198), .A2(n5197), .ZN(n5199) );
  NAND2_X1 U6657 ( .A1(n8880), .A2(n5199), .ZN(n7630) );
  INV_X1 U6658 ( .A(n5202), .ZN(n5200) );
  NAND2_X1 U6659 ( .A1(n5200), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5224) );
  INV_X1 U6660 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U6661 ( .A1(n5202), .A2(n5201), .ZN(n5203) );
  NAND2_X1 U6662 ( .A1(n5224), .A2(n5203), .ZN(n7631) );
  OR2_X1 U6663 ( .A1(n5129), .A2(n7631), .ZN(n5208) );
  INV_X1 U6664 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7529) );
  OR2_X1 U6665 ( .A1(n6888), .A2(n7529), .ZN(n5207) );
  NAND2_X1 U6666 ( .A1(n4458), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5206) );
  NAND2_X1 U6667 ( .A1(n5204), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5205) );
  NAND4_X1 U6668 ( .A1(n5208), .A2(n5207), .A3(n5206), .A4(n5205), .ZN(n8908)
         );
  AND2_X1 U6669 ( .A1(n8908), .A2(n8611), .ZN(n5219) );
  INV_X1 U6670 ( .A(n5210), .ZN(n5211) );
  NAND2_X1 U6671 ( .A1(n5211), .A2(SI_6_), .ZN(n5212) );
  MUX2_X1 U6672 ( .A(n6870), .B(n6868), .S(n4445), .Z(n5236) );
  XNOR2_X1 U6673 ( .A(n5236), .B(SI_7_), .ZN(n5234) );
  XNOR2_X1 U6674 ( .A(n5235), .B(n5234), .ZN(n6869) );
  OR2_X1 U6675 ( .A1(n5110), .A2(n6869), .ZN(n5217) );
  OR2_X1 U6676 ( .A1(n8234), .A2(n6870), .ZN(n5216) );
  NAND2_X1 U6677 ( .A1(n5190), .A2(n5213), .ZN(n5230) );
  NAND2_X1 U6678 ( .A1(n5230), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5214) );
  XNOR2_X1 U6679 ( .A(n5214), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6991) );
  INV_X1 U6680 ( .A(n6991), .ZN(n7141) );
  OR2_X1 U6681 ( .A1(n7001), .A2(n7141), .ZN(n5215) );
  XNOR2_X1 U6682 ( .A(n10239), .B(n5547), .ZN(n5218) );
  NAND2_X1 U6683 ( .A1(n5219), .A2(n5218), .ZN(n5222) );
  INV_X1 U6684 ( .A(n5218), .ZN(n7578) );
  INV_X1 U6685 ( .A(n5219), .ZN(n5220) );
  NAND2_X1 U6686 ( .A1(n7578), .A2(n5220), .ZN(n5221) );
  NAND2_X1 U6687 ( .A1(n5222), .A2(n5221), .ZN(n7629) );
  INV_X1 U6688 ( .A(n5222), .ZN(n5223) );
  NAND2_X1 U6689 ( .A1(n4458), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5229) );
  INV_X1 U6690 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6994) );
  OR2_X1 U6691 ( .A1(n5522), .A2(n6994), .ZN(n5228) );
  NAND2_X1 U6692 ( .A1(n5224), .A2(n8926), .ZN(n5225) );
  NAND2_X1 U6693 ( .A1(n5282), .A2(n5225), .ZN(n7654) );
  OR2_X1 U6694 ( .A1(n5129), .A2(n7654), .ZN(n5227) );
  INV_X1 U6695 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7655) );
  OR2_X1 U6696 ( .A1(n6888), .A2(n7655), .ZN(n5226) );
  NAND2_X1 U6697 ( .A1(n8907), .A2(n8611), .ZN(n5243) );
  NAND2_X1 U6698 ( .A1(n5232), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5231) );
  MUX2_X1 U6699 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5231), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5233) );
  NAND2_X1 U6700 ( .A1(n5233), .A2(n5272), .ZN(n8927) );
  INV_X1 U6701 ( .A(n5236), .ZN(n5237) );
  MUX2_X1 U6702 ( .A(n6874), .B(n6872), .S(n4445), .Z(n5238) );
  INV_X1 U6703 ( .A(n5238), .ZN(n5239) );
  NAND2_X1 U6704 ( .A1(n5239), .A2(SI_8_), .ZN(n5240) );
  NAND2_X1 U6705 ( .A1(n5254), .A2(n5240), .ZN(n5252) );
  XNOR2_X1 U6706 ( .A(n5253), .B(n5252), .ZN(n6871) );
  NAND2_X1 U6707 ( .A1(n6871), .A2(n8233), .ZN(n5242) );
  OR2_X1 U6708 ( .A1(n8234), .A2(n6874), .ZN(n5241) );
  OAI211_X1 U6709 ( .C1(n7001), .C2(n8927), .A(n5242), .B(n5241), .ZN(n7672)
         );
  XNOR2_X1 U6710 ( .A(n7672), .B(n5608), .ZN(n5244) );
  XNOR2_X1 U6711 ( .A(n5243), .B(n5244), .ZN(n7576) );
  INV_X1 U6712 ( .A(n5243), .ZN(n5245) );
  NAND2_X1 U6713 ( .A1(n5245), .A2(n5244), .ZN(n5246) );
  NAND2_X1 U6714 ( .A1(n4461), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5251) );
  INV_X1 U6715 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7686) );
  OR2_X1 U6716 ( .A1(n6888), .A2(n7686), .ZN(n5250) );
  INV_X1 U6717 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5280) );
  XNOR2_X1 U6718 ( .A(n5282), .B(n5280), .ZN(n7685) );
  OR2_X1 U6719 ( .A1(n5129), .A2(n7685), .ZN(n5249) );
  INV_X1 U6720 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5247) );
  OR2_X1 U6721 ( .A1(n8603), .A2(n5247), .ZN(n5248) );
  NOR2_X1 U6722 ( .A1(n7754), .A2(n6340), .ZN(n5263) );
  MUX2_X1 U6723 ( .A(n6905), .B(n6900), .S(n4445), .Z(n5257) );
  NAND2_X1 U6724 ( .A1(n5257), .A2(n5256), .ZN(n5268) );
  INV_X1 U6725 ( .A(n5257), .ZN(n5258) );
  NAND2_X1 U6726 ( .A1(n5258), .A2(SI_9_), .ZN(n5259) );
  XNOR2_X1 U6727 ( .A(n5267), .B(n5021), .ZN(n6899) );
  NAND2_X1 U6728 ( .A1(n6899), .A2(n8233), .ZN(n5262) );
  NAND2_X1 U6729 ( .A1(n5272), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5260) );
  XNOR2_X1 U6730 ( .A(n5260), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6996) );
  AOI22_X1 U6731 ( .A1(n4709), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n4711), .B2(
        n6996), .ZN(n5261) );
  NAND2_X1 U6732 ( .A1(n5262), .A2(n5261), .ZN(n7688) );
  XNOR2_X1 U6733 ( .A(n7688), .B(n5608), .ZN(n5264) );
  AND2_X1 U6734 ( .A1(n5263), .A2(n5264), .ZN(n7664) );
  INV_X1 U6735 ( .A(n5263), .ZN(n5266) );
  INV_X1 U6736 ( .A(n5264), .ZN(n5265) );
  NAND2_X1 U6737 ( .A1(n5266), .A2(n5265), .ZN(n7663) );
  MUX2_X1 U6738 ( .A(n6916), .B(n6907), .S(n4445), .Z(n5269) );
  INV_X1 U6739 ( .A(n5269), .ZN(n5270) );
  NAND2_X1 U6740 ( .A1(n5270), .A2(SI_10_), .ZN(n5271) );
  NAND2_X1 U6741 ( .A1(n6906), .A2(n8233), .ZN(n5277) );
  OAI21_X1 U6742 ( .B1(n5272), .B2(P2_IR_REG_9__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5274) );
  OR2_X1 U6743 ( .A1(n5274), .A2(n5273), .ZN(n5275) );
  NAND2_X1 U6744 ( .A1(n5274), .A2(n5273), .ZN(n5297) );
  AOI22_X1 U6745 ( .A1(n4709), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n4711), .B2(
        n6999), .ZN(n5276) );
  NAND2_X1 U6746 ( .A1(n5277), .A2(n5276), .ZN(n7849) );
  XNOR2_X1 U6747 ( .A(n7849), .B(n5547), .ZN(n5288) );
  NAND2_X1 U6748 ( .A1(n5204), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5287) );
  INV_X1 U6749 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5278) );
  OR2_X1 U6750 ( .A1(n8603), .A2(n5278), .ZN(n5286) );
  INV_X1 U6751 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5279) );
  OAI21_X1 U6752 ( .B1(n5282), .B2(n5280), .A(n5279), .ZN(n5283) );
  NAND2_X1 U6753 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5281) );
  NAND2_X1 U6754 ( .A1(n5283), .A2(n5302), .ZN(n7765) );
  OR2_X1 U6755 ( .A1(n5129), .A2(n7765), .ZN(n5285) );
  INV_X1 U6756 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7766) );
  OR2_X1 U6757 ( .A1(n6888), .A2(n7766), .ZN(n5284) );
  INV_X1 U6758 ( .A(n7861), .ZN(n8905) );
  NAND2_X1 U6759 ( .A1(n8905), .A2(n8611), .ZN(n5289) );
  XNOR2_X1 U6760 ( .A(n5288), .B(n5289), .ZN(n7716) );
  INV_X1 U6761 ( .A(n5288), .ZN(n5291) );
  INV_X1 U6762 ( .A(n5289), .ZN(n5290) );
  NAND2_X1 U6763 ( .A1(n5291), .A2(n5290), .ZN(n5292) );
  NAND2_X1 U6764 ( .A1(n5295), .A2(n5294), .ZN(n5314) );
  MUX2_X1 U6765 ( .A(n5296), .B(n6917), .S(n4445), .Z(n5315) );
  XNOR2_X1 U6766 ( .A(n5314), .B(n5312), .ZN(n6908) );
  NAND2_X1 U6767 ( .A1(n6908), .A2(n8233), .ZN(n5300) );
  NAND2_X1 U6768 ( .A1(n5297), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5298) );
  XNOR2_X1 U6769 ( .A(n5298), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7048) );
  AOI22_X1 U6770 ( .A1(n4709), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n4711), .B2(
        n7048), .ZN(n5299) );
  NAND2_X1 U6771 ( .A1(n5300), .A2(n5299), .ZN(n7919) );
  XNOR2_X1 U6772 ( .A(n7919), .B(n5608), .ZN(n5311) );
  NAND2_X1 U6773 ( .A1(n5204), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5308) );
  INV_X1 U6774 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7864) );
  OR2_X1 U6775 ( .A1(n6888), .A2(n7864), .ZN(n5307) );
  INV_X1 U6776 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7749) );
  NAND2_X1 U6777 ( .A1(n5302), .A2(n7749), .ZN(n5303) );
  NAND2_X1 U6778 ( .A1(n5349), .A2(n5303), .ZN(n7863) );
  OR2_X1 U6779 ( .A1(n5129), .A2(n7863), .ZN(n5306) );
  INV_X1 U6780 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5304) );
  OR2_X1 U6781 ( .A1(n8603), .A2(n5304), .ZN(n5305) );
  NAND2_X1 U6782 ( .A1(n8904), .A2(n8611), .ZN(n5309) );
  XNOR2_X1 U6783 ( .A(n5311), .B(n5309), .ZN(n7747) );
  INV_X1 U6784 ( .A(n5309), .ZN(n5310) );
  INV_X1 U6785 ( .A(n5312), .ZN(n5313) );
  INV_X1 U6786 ( .A(n5315), .ZN(n5316) );
  NAND2_X1 U6787 ( .A1(n5316), .A2(SI_11_), .ZN(n5317) );
  MUX2_X1 U6788 ( .A(n5319), .B(n7042), .S(n4445), .Z(n5321) );
  INV_X1 U6789 ( .A(SI_12_), .ZN(n5320) );
  INV_X1 U6790 ( .A(n5321), .ZN(n5322) );
  NAND2_X1 U6791 ( .A1(n5322), .A2(SI_12_), .ZN(n5323) );
  NAND2_X1 U6792 ( .A1(n5339), .A2(n5323), .ZN(n5338) );
  XNOR2_X1 U6793 ( .A(n5337), .B(n5338), .ZN(n6947) );
  NAND2_X1 U6794 ( .A1(n6947), .A2(n8233), .ZN(n5327) );
  OR2_X1 U6795 ( .A1(n5324), .A2(n9374), .ZN(n5325) );
  XNOR2_X1 U6796 ( .A(n5325), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7183) );
  AOI22_X1 U6797 ( .A1(n4709), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n4711), .B2(
        n7183), .ZN(n5326) );
  XNOR2_X1 U6798 ( .A(n7958), .B(n5547), .ZN(n5332) );
  NAND2_X1 U6799 ( .A1(n4458), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5331) );
  INV_X1 U6800 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7045) );
  OR2_X1 U6801 ( .A1(n5522), .A2(n7045), .ZN(n5330) );
  XNOR2_X1 U6802 ( .A(n5349), .B(n5348), .ZN(n7930) );
  OR2_X1 U6803 ( .A1(n5129), .A2(n7930), .ZN(n5329) );
  INV_X1 U6804 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7931) );
  OR2_X1 U6805 ( .A1(n6888), .A2(n7931), .ZN(n5328) );
  INV_X1 U6806 ( .A(n7980), .ZN(n8903) );
  NAND2_X1 U6807 ( .A1(n8903), .A2(n8611), .ZN(n5333) );
  NAND2_X1 U6808 ( .A1(n5332), .A2(n5333), .ZN(n7898) );
  NAND2_X1 U6809 ( .A1(n7900), .A2(n7898), .ZN(n5336) );
  INV_X1 U6810 ( .A(n5332), .ZN(n5335) );
  INV_X1 U6811 ( .A(n5333), .ZN(n5334) );
  NAND2_X1 U6812 ( .A1(n5335), .A2(n5334), .ZN(n7899) );
  MUX2_X1 U6813 ( .A(n7193), .B(n7204), .S(n4445), .Z(n5340) );
  INV_X1 U6814 ( .A(n5340), .ZN(n5341) );
  NAND2_X1 U6815 ( .A1(n5341), .A2(SI_13_), .ZN(n5342) );
  XNOR2_X1 U6816 ( .A(n5359), .B(n4479), .ZN(n7191) );
  NAND2_X1 U6817 ( .A1(n7191), .A2(n8233), .ZN(n5345) );
  NAND2_X1 U6818 ( .A1(n5343), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5363) );
  XNOR2_X1 U6819 ( .A(n5363), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7233) );
  AOI22_X1 U6820 ( .A1(n4709), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n4711), .B2(
        n7233), .ZN(n5344) );
  XNOR2_X1 U6821 ( .A(n8704), .B(n5608), .ZN(n5355) );
  INV_X1 U6822 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5346) );
  OR2_X1 U6823 ( .A1(n5522), .A2(n5346), .ZN(n5354) );
  OAI21_X1 U6824 ( .B1(n5349), .B2(n5348), .A(n5347), .ZN(n5350) );
  NAND2_X1 U6825 ( .A1(n5350), .A2(n5369), .ZN(n7979) );
  OR2_X1 U6826 ( .A1(n5129), .A2(n7979), .ZN(n5353) );
  INV_X1 U6827 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7969) );
  OR2_X1 U6828 ( .A1(n6888), .A2(n7969), .ZN(n5352) );
  NAND2_X1 U6829 ( .A1(n4458), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5351) );
  NAND4_X1 U6830 ( .A1(n5354), .A2(n5353), .A3(n5352), .A4(n5351), .ZN(n8902)
         );
  AND2_X1 U6831 ( .A1(n8902), .A2(n8611), .ZN(n5356) );
  NAND2_X1 U6832 ( .A1(n5355), .A2(n5356), .ZN(n5375) );
  INV_X1 U6833 ( .A(n5355), .ZN(n8094) );
  INV_X1 U6834 ( .A(n5356), .ZN(n5357) );
  NAND2_X1 U6835 ( .A1(n8094), .A2(n5357), .ZN(n5358) );
  AND2_X1 U6836 ( .A1(n5375), .A2(n5358), .ZN(n7978) );
  NAND2_X1 U6837 ( .A1(n5361), .A2(n5360), .ZN(n5386) );
  MUX2_X1 U6838 ( .A(n7213), .B(n7195), .S(n4445), .Z(n5382) );
  XNOR2_X1 U6839 ( .A(n5382), .B(SI_14_), .ZN(n5381) );
  NAND2_X1 U6840 ( .A1(n7194), .A2(n8233), .ZN(n5366) );
  NAND2_X1 U6841 ( .A1(n5363), .A2(n5362), .ZN(n5364) );
  NAND2_X1 U6842 ( .A1(n5364), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5392) );
  XNOR2_X1 U6843 ( .A(n5392), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7412) );
  AOI22_X1 U6844 ( .A1(n4709), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n4711), .B2(
        n7412), .ZN(n5365) );
  NAND2_X2 U6845 ( .A1(n5366), .A2(n5365), .ZN(n8711) );
  XNOR2_X1 U6846 ( .A(n8711), .B(n5608), .ZN(n5377) );
  INV_X1 U6847 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5367) );
  OR2_X1 U6848 ( .A1(n5522), .A2(n5367), .ZN(n5374) );
  INV_X1 U6849 ( .A(n5369), .ZN(n5368) );
  INV_X1 U6850 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U6851 ( .A1(n5369), .A2(n6708), .ZN(n5370) );
  NAND2_X1 U6852 ( .A1(n5397), .A2(n5370), .ZN(n8100) );
  OR2_X1 U6853 ( .A1(n5129), .A2(n8100), .ZN(n5373) );
  INV_X1 U6854 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8015) );
  OR2_X1 U6855 ( .A1(n6888), .A2(n8015), .ZN(n5372) );
  NAND2_X1 U6856 ( .A1(n4459), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5371) );
  NAND4_X1 U6857 ( .A1(n5374), .A2(n5373), .A3(n5372), .A4(n5371), .ZN(n9265)
         );
  NAND2_X1 U6858 ( .A1(n9265), .A2(n8611), .ZN(n5378) );
  XNOR2_X1 U6859 ( .A(n5377), .B(n5378), .ZN(n8105) );
  AND2_X1 U6860 ( .A1(n8105), .A2(n5375), .ZN(n5376) );
  INV_X1 U6861 ( .A(n5377), .ZN(n5379) );
  NAND2_X1 U6862 ( .A1(n5379), .A2(n5378), .ZN(n5380) );
  INV_X1 U6863 ( .A(n5381), .ZN(n5385) );
  INV_X1 U6864 ( .A(n5382), .ZN(n5383) );
  NAND2_X1 U6865 ( .A1(n5383), .A2(SI_14_), .ZN(n5384) );
  MUX2_X1 U6866 ( .A(n7325), .B(n7327), .S(n4445), .Z(n5388) );
  INV_X1 U6867 ( .A(SI_15_), .ZN(n5387) );
  NAND2_X1 U6868 ( .A1(n5388), .A2(n5387), .ZN(n5407) );
  INV_X1 U6869 ( .A(n5388), .ZN(n5389) );
  NAND2_X1 U6870 ( .A1(n5389), .A2(SI_15_), .ZN(n5390) );
  NAND2_X1 U6871 ( .A1(n5407), .A2(n5390), .ZN(n5408) );
  XNOR2_X1 U6872 ( .A(n5409), .B(n5408), .ZN(n7324) );
  NAND2_X1 U6873 ( .A1(n7324), .A2(n8233), .ZN(n5396) );
  NAND2_X1 U6874 ( .A1(n5392), .A2(n5391), .ZN(n5393) );
  NAND2_X1 U6875 ( .A1(n5393), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5394) );
  XNOR2_X1 U6876 ( .A(n5394), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7939) );
  AOI22_X1 U6877 ( .A1(n4709), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n4711), .B2(
        n7939), .ZN(n5395) );
  XNOR2_X1 U6878 ( .A(n9350), .B(n5608), .ZN(n5404) );
  NAND2_X1 U6879 ( .A1(n4458), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5403) );
  INV_X1 U6880 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7414) );
  OR2_X1 U6881 ( .A1(n5522), .A2(n7414), .ZN(n5402) );
  INV_X1 U6882 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8145) );
  NAND2_X1 U6883 ( .A1(n5397), .A2(n8145), .ZN(n5398) );
  NAND2_X1 U6884 ( .A1(n5419), .A2(n5398), .ZN(n9257) );
  OR2_X1 U6885 ( .A1(n5129), .A2(n9257), .ZN(n5401) );
  INV_X1 U6886 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n5399) );
  OR2_X1 U6887 ( .A1(n6888), .A2(n5399), .ZN(n5400) );
  NAND2_X1 U6888 ( .A1(n8901), .A2(n8611), .ZN(n8141) );
  NAND2_X1 U6889 ( .A1(n5405), .A2(n4907), .ZN(n5406) );
  MUX2_X1 U6890 ( .A(n7359), .B(n7384), .S(n4445), .Z(n5411) );
  INV_X1 U6891 ( .A(SI_16_), .ZN(n5410) );
  NAND2_X1 U6892 ( .A1(n5411), .A2(n5410), .ZN(n5432) );
  INV_X1 U6893 ( .A(n5411), .ZN(n5412) );
  NAND2_X1 U6894 ( .A1(n5412), .A2(SI_16_), .ZN(n5413) );
  XNOR2_X1 U6895 ( .A(n5431), .B(n5430), .ZN(n7358) );
  NAND2_X1 U6896 ( .A1(n7358), .A2(n8233), .ZN(n5417) );
  NAND2_X1 U6897 ( .A1(n5414), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5415) );
  XNOR2_X1 U6898 ( .A(n5415), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8961) );
  AOI22_X1 U6899 ( .A1(n4709), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n4711), .B2(
        n8961), .ZN(n5416) );
  XNOR2_X1 U6900 ( .A(n9345), .B(n5608), .ZN(n5425) );
  NAND2_X1 U6901 ( .A1(n4459), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5424) );
  INV_X1 U6902 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n6548) );
  OR2_X1 U6903 ( .A1(n5522), .A2(n6548), .ZN(n5423) );
  INV_X1 U6904 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8955) );
  NAND2_X1 U6905 ( .A1(n5419), .A2(n8955), .ZN(n5420) );
  NAND2_X1 U6906 ( .A1(n5459), .A2(n5420), .ZN(n8185) );
  OR2_X1 U6907 ( .A1(n5129), .A2(n8185), .ZN(n5422) );
  INV_X1 U6908 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8175) );
  OR2_X1 U6909 ( .A1(n6888), .A2(n8175), .ZN(n5421) );
  INV_X1 U6910 ( .A(n9232), .ZN(n9267) );
  NAND2_X1 U6911 ( .A1(n9267), .A2(n8611), .ZN(n5426) );
  XNOR2_X1 U6912 ( .A(n5425), .B(n5426), .ZN(n8184) );
  NAND2_X1 U6913 ( .A1(n8183), .A2(n8184), .ZN(n5429) );
  INV_X1 U6914 ( .A(n5425), .ZN(n5427) );
  NAND2_X1 U6915 ( .A1(n5427), .A2(n5426), .ZN(n5428) );
  INV_X1 U6916 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5433) );
  MUX2_X1 U6917 ( .A(n5433), .B(n7467), .S(n4445), .Z(n5450) );
  XNOR2_X1 U6918 ( .A(n5450), .B(SI_17_), .ZN(n5449) );
  XNOR2_X1 U6919 ( .A(n5454), .B(n5449), .ZN(n7404) );
  NAND2_X1 U6920 ( .A1(n7404), .A2(n8233), .ZN(n5438) );
  INV_X1 U6921 ( .A(n5434), .ZN(n5435) );
  NAND2_X1 U6922 ( .A1(n5435), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5436) );
  XNOR2_X1 U6923 ( .A(n5436), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8971) );
  AOI22_X1 U6924 ( .A1(n4709), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n4711), .B2(
        n8971), .ZN(n5437) );
  XNOR2_X1 U6925 ( .A(n9247), .B(n5608), .ZN(n5443) );
  NAND2_X1 U6926 ( .A1(n4461), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5442) );
  INV_X1 U6927 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n6586) );
  OR2_X1 U6928 ( .A1(n8603), .A2(n6586), .ZN(n5441) );
  INV_X1 U6929 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8969) );
  XNOR2_X1 U6930 ( .A(n5459), .B(n8969), .ZN(n9242) );
  OR2_X1 U6931 ( .A1(n5129), .A2(n9242), .ZN(n5440) );
  INV_X1 U6932 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9243) );
  OR2_X1 U6933 ( .A1(n6888), .A2(n9243), .ZN(n5439) );
  NOR2_X1 U6934 ( .A1(n8874), .A2(n6340), .ZN(n5444) );
  NAND2_X1 U6935 ( .A1(n5443), .A2(n5444), .ZN(n5448) );
  INV_X1 U6936 ( .A(n5443), .ZN(n8870) );
  INV_X1 U6937 ( .A(n5444), .ZN(n5445) );
  NAND2_X1 U6938 ( .A1(n8870), .A2(n5445), .ZN(n5446) );
  NAND2_X1 U6939 ( .A1(n5448), .A2(n5446), .ZN(n6765) );
  INV_X1 U6940 ( .A(n6765), .ZN(n5447) );
  INV_X1 U6941 ( .A(n5449), .ZN(n5453) );
  INV_X1 U6942 ( .A(n5450), .ZN(n5451) );
  NAND2_X1 U6943 ( .A1(n5451), .A2(SI_17_), .ZN(n5452) );
  MUX2_X1 U6944 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4445), .Z(n5473) );
  XNOR2_X1 U6945 ( .A(n5473), .B(SI_18_), .ZN(n5470) );
  XNOR2_X1 U6946 ( .A(n5472), .B(n5470), .ZN(n7606) );
  NAND2_X1 U6947 ( .A1(n7606), .A2(n8233), .ZN(n5457) );
  XNOR2_X1 U6948 ( .A(n5455), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8987) );
  AOI22_X1 U6949 ( .A1(n4709), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n4711), .B2(
        n8987), .ZN(n5456) );
  XNOR2_X1 U6950 ( .A(n9336), .B(n5608), .ZN(n8564) );
  INV_X1 U6951 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7944) );
  OR2_X1 U6952 ( .A1(n5522), .A2(n7944), .ZN(n5464) );
  INV_X1 U6953 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8873) );
  OAI21_X1 U6954 ( .B1(n5459), .B2(n8969), .A(n8873), .ZN(n5460) );
  NAND2_X1 U6955 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_17__SCAN_IN), 
        .ZN(n5458) );
  NAND2_X1 U6956 ( .A1(n5460), .A2(n5483), .ZN(n9212) );
  OR2_X1 U6957 ( .A1(n4454), .A2(n9212), .ZN(n5463) );
  NAND2_X1 U6958 ( .A1(n4459), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U6959 ( .A1(n8599), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5461) );
  NAND4_X1 U6960 ( .A1(n5464), .A2(n5463), .A3(n5462), .A4(n5461), .ZN(n9008)
         );
  AND2_X1 U6961 ( .A1(n9008), .A2(n8611), .ZN(n5465) );
  NAND2_X1 U6962 ( .A1(n8564), .A2(n5465), .ZN(n5489) );
  INV_X1 U6963 ( .A(n8564), .ZN(n5467) );
  INV_X1 U6964 ( .A(n5465), .ZN(n5466) );
  NAND2_X1 U6965 ( .A1(n5467), .A2(n5466), .ZN(n5468) );
  AND2_X1 U6966 ( .A1(n5489), .A2(n5468), .ZN(n8867) );
  NAND2_X1 U6967 ( .A1(n5469), .A2(n8867), .ZN(n8563) );
  NAND2_X1 U6968 ( .A1(n5473), .A2(SI_18_), .ZN(n5474) );
  MUX2_X1 U6969 ( .A(n7706), .B(n7704), .S(n4445), .Z(n5476) );
  INV_X1 U6970 ( .A(SI_19_), .ZN(n5475) );
  NAND2_X1 U6971 ( .A1(n5476), .A2(n5475), .ZN(n5495) );
  INV_X1 U6972 ( .A(n5476), .ZN(n5477) );
  NAND2_X1 U6973 ( .A1(n5477), .A2(SI_19_), .ZN(n5478) );
  NAND2_X1 U6974 ( .A1(n5495), .A2(n5478), .ZN(n5496) );
  NAND2_X1 U6975 ( .A1(n7703), .A2(n8233), .ZN(n5481) );
  AOI22_X1 U6976 ( .A1(n4709), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n4455), .B2(
        n4711), .ZN(n5480) );
  XNOR2_X1 U6977 ( .A(n9332), .B(n5608), .ZN(n5491) );
  NAND2_X1 U6978 ( .A1(n4458), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5488) );
  INV_X1 U6979 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U6980 ( .A1(n5483), .A2(n8569), .ZN(n5484) );
  NAND2_X1 U6981 ( .A1(n5503), .A2(n5484), .ZN(n9193) );
  OR2_X1 U6982 ( .A1(n5129), .A2(n9193), .ZN(n5487) );
  NAND2_X1 U6983 ( .A1(n5204), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U6984 ( .A1(n8599), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5485) );
  NAND4_X1 U6985 ( .A1(n5488), .A2(n5487), .A3(n5486), .A4(n5485), .ZN(n9210)
         );
  NAND2_X1 U6986 ( .A1(n9210), .A2(n4446), .ZN(n5492) );
  XNOR2_X1 U6987 ( .A(n5491), .B(n5492), .ZN(n8566) );
  AND2_X1 U6988 ( .A1(n8566), .A2(n5489), .ZN(n5490) );
  INV_X1 U6989 ( .A(n5491), .ZN(n5493) );
  NAND2_X1 U6990 ( .A1(n5493), .A2(n5492), .ZN(n5494) );
  MUX2_X1 U6991 ( .A(n7734), .B(n7732), .S(n4445), .Z(n5498) );
  INV_X1 U6992 ( .A(SI_20_), .ZN(n6577) );
  NAND2_X1 U6993 ( .A1(n5498), .A2(n6577), .ZN(n5517) );
  INV_X1 U6994 ( .A(n5498), .ZN(n5499) );
  NAND2_X1 U6995 ( .A1(n5499), .A2(SI_20_), .ZN(n5500) );
  XNOR2_X1 U6996 ( .A(n5516), .B(n5515), .ZN(n7731) );
  NAND2_X1 U6997 ( .A1(n7731), .A2(n8233), .ZN(n5502) );
  OR2_X1 U6998 ( .A1(n8234), .A2(n7734), .ZN(n5501) );
  XNOR2_X1 U6999 ( .A(n9325), .B(n5608), .ZN(n5510) );
  NAND2_X1 U7000 ( .A1(n4461), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5509) );
  INV_X1 U7001 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n6556) );
  OR2_X1 U7002 ( .A1(n8603), .A2(n6556), .ZN(n5508) );
  INV_X1 U7003 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6775) );
  NAND2_X1 U7004 ( .A1(n5503), .A2(n6775), .ZN(n5504) );
  NAND2_X1 U7005 ( .A1(n5524), .A2(n5504), .ZN(n9181) );
  OR2_X1 U7006 ( .A1(n4454), .A2(n9181), .ZN(n5507) );
  INV_X1 U7007 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5505) );
  OR2_X1 U7008 ( .A1(n6888), .A2(n5505), .ZN(n5506) );
  NOR2_X1 U7009 ( .A1(n9175), .A2(n6340), .ZN(n5511) );
  NAND2_X1 U7010 ( .A1(n5510), .A2(n5511), .ZN(n5514) );
  INV_X1 U7011 ( .A(n5510), .ZN(n8834) );
  INV_X1 U7012 ( .A(n5511), .ZN(n5512) );
  NAND2_X1 U7013 ( .A1(n8834), .A2(n5512), .ZN(n5513) );
  NAND2_X1 U7014 ( .A1(n5514), .A2(n5513), .ZN(n6774) );
  NAND2_X1 U7015 ( .A1(n6771), .A2(n5514), .ZN(n5530) );
  NAND2_X1 U7016 ( .A1(n5518), .A2(n5517), .ZN(n5537) );
  MUX2_X1 U7017 ( .A(n7802), .B(n7783), .S(n4445), .Z(n5538) );
  XNOR2_X1 U7018 ( .A(n5538), .B(SI_21_), .ZN(n5535) );
  XNOR2_X1 U7019 ( .A(n5537), .B(n5535), .ZN(n7782) );
  NAND2_X1 U7020 ( .A1(n7782), .A2(n8233), .ZN(n5520) );
  OR2_X1 U7021 ( .A1(n8234), .A2(n7802), .ZN(n5519) );
  XNOR2_X1 U7022 ( .A(n9164), .B(n5547), .ZN(n5533) );
  NAND2_X1 U7023 ( .A1(n4458), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5529) );
  INV_X1 U7024 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n5521) );
  OR2_X1 U7025 ( .A1(n5522), .A2(n5521), .ZN(n5528) );
  INV_X1 U7026 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8838) );
  NAND2_X1 U7027 ( .A1(n5524), .A2(n8838), .ZN(n5525) );
  NAND2_X1 U7028 ( .A1(n5548), .A2(n5525), .ZN(n9165) );
  OR2_X1 U7029 ( .A1(n5129), .A2(n9165), .ZN(n5527) );
  INV_X1 U7030 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9166) );
  OR2_X1 U7031 ( .A1(n6888), .A2(n9166), .ZN(n5526) );
  NAND2_X1 U7032 ( .A1(n9187), .A2(n8611), .ZN(n5531) );
  XNOR2_X1 U7033 ( .A(n5533), .B(n5531), .ZN(n8832) );
  INV_X1 U7034 ( .A(n5531), .ZN(n5532) );
  NAND2_X1 U7035 ( .A1(n5533), .A2(n5532), .ZN(n5534) );
  INV_X1 U7036 ( .A(n5535), .ZN(n5536) );
  INV_X1 U7037 ( .A(n5538), .ZN(n5539) );
  NAND2_X1 U7038 ( .A1(n5539), .A2(SI_21_), .ZN(n5540) );
  MUX2_X1 U7039 ( .A(n7880), .B(n7878), .S(n4445), .Z(n5542) );
  INV_X1 U7040 ( .A(SI_22_), .ZN(n5541) );
  NAND2_X1 U7041 ( .A1(n5542), .A2(n5541), .ZN(n5559) );
  INV_X1 U7042 ( .A(n5542), .ZN(n5543) );
  NAND2_X1 U7043 ( .A1(n5543), .A2(SI_22_), .ZN(n5544) );
  NAND2_X1 U7044 ( .A1(n5559), .A2(n5544), .ZN(n5560) );
  XNOR2_X1 U7045 ( .A(n5561), .B(n5560), .ZN(n7877) );
  NAND2_X1 U7046 ( .A1(n7877), .A2(n8233), .ZN(n5546) );
  OR2_X1 U7047 ( .A1(n8234), .A2(n7880), .ZN(n5545) );
  XNOR2_X1 U7048 ( .A(n9316), .B(n5547), .ZN(n5555) );
  XNOR2_X2 U7049 ( .A(n5557), .B(n5555), .ZN(n8859) );
  NAND2_X1 U7050 ( .A1(n4458), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5554) );
  INV_X1 U7051 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6718) );
  OR2_X1 U7052 ( .A1(n5522), .A2(n6718), .ZN(n5553) );
  INV_X1 U7053 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8862) );
  NAND2_X1 U7054 ( .A1(n5548), .A2(n8862), .ZN(n5549) );
  NAND2_X1 U7055 ( .A1(n5583), .A2(n5549), .ZN(n9151) );
  OR2_X1 U7056 ( .A1(n5129), .A2(n9151), .ZN(n5552) );
  INV_X1 U7057 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5550) );
  OR2_X1 U7058 ( .A1(n6888), .A2(n5550), .ZN(n5551) );
  INV_X1 U7059 ( .A(n9176), .ZN(n8900) );
  NAND2_X1 U7060 ( .A1(n8900), .A2(n4446), .ZN(n8858) );
  INV_X1 U7061 ( .A(n5555), .ZN(n5556) );
  NOR2_X1 U7062 ( .A1(n5557), .A2(n5556), .ZN(n5558) );
  AOI21_X2 U7063 ( .B1(n8859), .B2(n8858), .A(n5558), .ZN(n5592) );
  MUX2_X1 U7064 ( .A(n7987), .B(n7993), .S(n4445), .Z(n5563) );
  INV_X1 U7065 ( .A(SI_23_), .ZN(n5562) );
  NAND2_X1 U7066 ( .A1(n5563), .A2(n5562), .ZN(n5571) );
  INV_X1 U7067 ( .A(n5563), .ZN(n5564) );
  NAND2_X1 U7068 ( .A1(n5564), .A2(SI_23_), .ZN(n5565) );
  NAND2_X1 U7069 ( .A1(n7989), .A2(n8233), .ZN(n5567) );
  OR2_X1 U7070 ( .A1(n8234), .A2(n7987), .ZN(n5566) );
  XNOR2_X1 U7071 ( .A(n9311), .B(n5608), .ZN(n5591) );
  XNOR2_X2 U7072 ( .A(n5592), .B(n5568), .ZN(n8811) );
  MUX2_X1 U7073 ( .A(n8023), .B(n8021), .S(n4445), .Z(n5597) );
  XNOR2_X1 U7074 ( .A(n5597), .B(SI_24_), .ZN(n5596) );
  NAND2_X1 U7075 ( .A1(n8020), .A2(n8233), .ZN(n5574) );
  OR2_X1 U7076 ( .A1(n8234), .A2(n8023), .ZN(n5573) );
  XNOR2_X1 U7077 ( .A(n9304), .B(n5608), .ZN(n5593) );
  INV_X1 U7078 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n5580) );
  INV_X1 U7079 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8813) );
  INV_X1 U7080 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7081 ( .A1(n5585), .A2(n5576), .ZN(n5577) );
  NAND2_X1 U7082 ( .A1(n5610), .A2(n5577), .ZN(n9114) );
  OR2_X1 U7083 ( .A1(n9114), .A2(n4454), .ZN(n5579) );
  AOI22_X1 U7084 ( .A1(n4459), .A2(P2_REG0_REG_24__SCAN_IN), .B1(n5204), .B2(
        P2_REG1_REG_24__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7085 ( .A1(n4459), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U7086 ( .A1(n4461), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5581) );
  AND2_X1 U7087 ( .A1(n5582), .A2(n5581), .ZN(n5588) );
  NAND2_X1 U7088 ( .A1(n5583), .A2(n8813), .ZN(n5584) );
  AND2_X1 U7089 ( .A1(n5585), .A2(n5584), .ZN(n8812) );
  NAND2_X1 U7090 ( .A1(n8812), .A2(n6353), .ZN(n5587) );
  NAND2_X1 U7091 ( .A1(n8599), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5586) );
  NOR2_X1 U7092 ( .A1(n9021), .A2(n6340), .ZN(n8810) );
  AND2_X1 U7093 ( .A1(n5592), .A2(n5591), .ZN(n8843) );
  INV_X1 U7094 ( .A(n5593), .ZN(n8845) );
  NAND2_X1 U7095 ( .A1(n9136), .A2(n8611), .ZN(n8849) );
  NAND2_X1 U7096 ( .A1(n8845), .A2(n8849), .ZN(n5595) );
  INV_X1 U7097 ( .A(n8849), .ZN(n5594) );
  INV_X1 U7098 ( .A(n5596), .ZN(n5600) );
  INV_X1 U7099 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U7100 ( .A1(n5598), .A2(SI_24_), .ZN(n5599) );
  INV_X1 U7101 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8151) );
  MUX2_X1 U7102 ( .A(n8151), .B(n8156), .S(n4445), .Z(n5603) );
  INV_X1 U7103 ( .A(SI_25_), .ZN(n5602) );
  NAND2_X1 U7104 ( .A1(n5603), .A2(n5602), .ZN(n5617) );
  INV_X1 U7105 ( .A(n5603), .ZN(n5604) );
  NAND2_X1 U7106 ( .A1(n5604), .A2(SI_25_), .ZN(n5605) );
  NAND2_X1 U7107 ( .A1(n5617), .A2(n5605), .ZN(n5618) );
  XNOR2_X1 U7108 ( .A(n5619), .B(n5618), .ZN(n8150) );
  NAND2_X1 U7109 ( .A1(n8150), .A2(n8233), .ZN(n5607) );
  OR2_X1 U7110 ( .A1(n8234), .A2(n8151), .ZN(n5606) );
  XNOR2_X1 U7111 ( .A(n9301), .B(n5608), .ZN(n6363) );
  INV_X1 U7112 ( .A(n5610), .ZN(n5609) );
  NAND2_X1 U7113 ( .A1(n5609), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5626) );
  INV_X1 U7114 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U7115 ( .A1(n5610), .A2(n6550), .ZN(n5611) );
  NAND2_X1 U7116 ( .A1(n5626), .A2(n5611), .ZN(n9106) );
  OR2_X1 U7117 ( .A1(n9106), .A2(n5129), .ZN(n5614) );
  AOI22_X1 U7118 ( .A1(n4459), .A2(P2_REG0_REG_25__SCAN_IN), .B1(n4461), .B2(
        P2_REG1_REG_25__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7119 ( .A1(n8599), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5612) );
  NOR2_X1 U7120 ( .A1(n8851), .A2(n6340), .ZN(n5615) );
  NAND2_X1 U7121 ( .A1(n6363), .A2(n5615), .ZN(n5616) );
  OAI21_X1 U7122 ( .B1(n6363), .B2(n5615), .A(n5616), .ZN(n6326) );
  INV_X1 U7123 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8180) );
  INV_X1 U7124 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8159) );
  MUX2_X1 U7125 ( .A(n8180), .B(n8159), .S(n4445), .Z(n5620) );
  INV_X1 U7126 ( .A(SI_26_), .ZN(n6653) );
  NAND2_X1 U7127 ( .A1(n5620), .A2(n6653), .ZN(n5639) );
  INV_X1 U7128 ( .A(n5620), .ZN(n5621) );
  NAND2_X1 U7129 ( .A1(n5621), .A2(SI_26_), .ZN(n5622) );
  XNOR2_X1 U7130 ( .A(n5638), .B(n5637), .ZN(n8157) );
  NAND2_X1 U7131 ( .A1(n8157), .A2(n8233), .ZN(n5624) );
  OR2_X1 U7132 ( .A1(n8234), .A2(n8180), .ZN(n5623) );
  XNOR2_X1 U7133 ( .A(n9295), .B(n5608), .ZN(n5633) );
  INV_X1 U7134 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7135 ( .A1(n5626), .A2(n5625), .ZN(n5627) );
  AND2_X1 U7136 ( .A1(n5649), .A2(n5627), .ZN(n6368) );
  NAND2_X1 U7137 ( .A1(n6368), .A2(n6353), .ZN(n5632) );
  INV_X1 U7138 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9083) );
  NAND2_X1 U7139 ( .A1(n4458), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U7140 ( .A1(n5204), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5628) );
  OAI211_X1 U7141 ( .C1(n9083), .C2(n6888), .A(n5629), .B(n5628), .ZN(n5630)
         );
  INV_X1 U7142 ( .A(n5630), .ZN(n5631) );
  NOR2_X1 U7143 ( .A1(n9072), .A2(n6340), .ZN(n5634) );
  NAND2_X1 U7144 ( .A1(n5633), .A2(n5634), .ZN(n5697) );
  INV_X1 U7145 ( .A(n5633), .ZN(n5694) );
  INV_X1 U7146 ( .A(n5634), .ZN(n5635) );
  NAND2_X1 U7147 ( .A1(n5694), .A2(n5635), .ZN(n5636) );
  NAND2_X1 U7148 ( .A1(n5638), .A2(n5637), .ZN(n5640) );
  INV_X1 U7149 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8578) );
  INV_X1 U7150 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8577) );
  MUX2_X1 U7151 ( .A(n8578), .B(n8577), .S(n4445), .Z(n5642) );
  INV_X1 U7152 ( .A(SI_27_), .ZN(n5641) );
  NAND2_X1 U7153 ( .A1(n5642), .A2(n5641), .ZN(n6336) );
  INV_X1 U7154 ( .A(n5642), .ZN(n5643) );
  NAND2_X1 U7155 ( .A1(n5643), .A2(SI_27_), .ZN(n5644) );
  NAND2_X1 U7156 ( .A1(n8576), .A2(n8233), .ZN(n5646) );
  OR2_X1 U7157 ( .A1(n8234), .A2(n8578), .ZN(n5645) );
  XNOR2_X1 U7158 ( .A(n9290), .B(n5608), .ZN(n5656) );
  INV_X1 U7159 ( .A(n5649), .ZN(n5647) );
  NAND2_X1 U7160 ( .A1(n5647), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5709) );
  INV_X1 U7161 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U7162 ( .A1(n5649), .A2(n5648), .ZN(n5650) );
  NAND2_X1 U7163 ( .A1(n5709), .A2(n5650), .ZN(n9068) );
  OR2_X1 U7164 ( .A1(n9068), .A2(n4454), .ZN(n5655) );
  INV_X1 U7165 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6645) );
  NAND2_X1 U7166 ( .A1(n4459), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U7167 ( .A1(n8599), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5651) );
  OAI211_X1 U7168 ( .C1(n5522), .C2(n6645), .A(n5652), .B(n5651), .ZN(n5653)
         );
  INV_X1 U7169 ( .A(n5653), .ZN(n5654) );
  NOR2_X1 U7170 ( .A1(n9031), .A2(n6340), .ZN(n5657) );
  NAND2_X1 U7171 ( .A1(n5656), .A2(n5657), .ZN(n6345) );
  INV_X1 U7172 ( .A(n5656), .ZN(n5659) );
  INV_X1 U7173 ( .A(n5657), .ZN(n5658) );
  NAND2_X1 U7174 ( .A1(n5659), .A2(n5658), .ZN(n5660) );
  NAND2_X1 U7175 ( .A1(n6345), .A2(n5660), .ZN(n5698) );
  NAND2_X1 U7176 ( .A1(n5661), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5662) );
  MUX2_X1 U7177 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5662), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5664) );
  NAND2_X1 U7178 ( .A1(n5664), .A2(n5663), .ZN(n8152) );
  NAND2_X1 U7179 ( .A1(n4538), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U7180 ( .A1(n5687), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5666) );
  INV_X1 U7181 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5665) );
  INV_X1 U7182 ( .A(P2_B_REG_SCAN_IN), .ZN(n5667) );
  XOR2_X1 U7183 ( .A(n8025), .B(n5667), .Z(n5668) );
  AND2_X1 U7184 ( .A1(n8152), .A2(n5668), .ZN(n5673) );
  NAND2_X1 U7185 ( .A1(n5663), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5669) );
  MUX2_X1 U7186 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5669), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5672) );
  INV_X1 U7187 ( .A(n5670), .ZN(n5671) );
  INV_X1 U7188 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10214) );
  AND2_X1 U7189 ( .A1(n8182), .A2(n8152), .ZN(n10215) );
  NOR4_X1 U7190 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n5677) );
  NOR4_X1 U7191 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5676) );
  NOR4_X1 U7192 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5675) );
  NOR4_X1 U7193 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5674) );
  NAND4_X1 U7194 ( .A1(n5677), .A2(n5676), .A3(n5675), .A4(n5674), .ZN(n5683)
         );
  NOR2_X1 U7195 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .ZN(
        n5681) );
  NOR4_X1 U7196 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5680) );
  NOR4_X1 U7197 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n5679) );
  NOR4_X1 U7198 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5678) );
  NAND4_X1 U7199 ( .A1(n5681), .A2(n5680), .A3(n5679), .A4(n5678), .ZN(n5682)
         );
  OAI21_X1 U7200 ( .B1(n5683), .B2(n5682), .A(n10199), .ZN(n7022) );
  INV_X1 U7201 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10211) );
  AND2_X1 U7202 ( .A1(n8182), .A2(n8025), .ZN(n10212) );
  AOI21_X1 U7203 ( .B1(n10199), .B2(n10211), .A(n10212), .ZN(n7126) );
  AND2_X1 U7204 ( .A1(n7022), .A2(n7126), .ZN(n5684) );
  NAND2_X1 U7205 ( .A1(n7420), .A2(n5684), .ZN(n5705) );
  NOR2_X1 U7206 ( .A1(n8182), .A2(n8152), .ZN(n5686) );
  INV_X1 U7207 ( .A(n8025), .ZN(n5685) );
  OAI21_X1 U7208 ( .B1(n5689), .B2(n5688), .A(n5687), .ZN(n6895) );
  INV_X1 U7209 ( .A(n10216), .ZN(n5690) );
  NOR2_X1 U7210 ( .A1(n5705), .A2(n10200), .ZN(n5717) );
  INV_X1 U7211 ( .A(n6972), .ZN(n5691) );
  AOI21_X1 U7212 ( .B1(n5696), .B2(n5698), .A(n8868), .ZN(n5693) );
  INV_X1 U7213 ( .A(n5693), .ZN(n5695) );
  INV_X1 U7214 ( .A(n5696), .ZN(n6365) );
  INV_X1 U7215 ( .A(n5697), .ZN(n5700) );
  INV_X1 U7216 ( .A(n5698), .ZN(n5699) );
  NAND2_X1 U7217 ( .A1(n5701), .A2(n6360), .ZN(n5724) );
  NAND2_X1 U7218 ( .A1(n5717), .A2(n4539), .ZN(n5703) );
  INV_X1 U7219 ( .A(n7019), .ZN(n5704) );
  NAND2_X1 U7220 ( .A1(n5705), .A2(n5704), .ZN(n5708) );
  INV_X1 U7221 ( .A(n6895), .ZN(n5706) );
  AND2_X1 U7222 ( .A1(n8799), .A2(n6972), .ZN(n7020) );
  NOR3_X1 U7223 ( .A1(n6970), .A2(n5706), .A3(n7020), .ZN(n5707) );
  NAND2_X1 U7224 ( .A1(n5708), .A2(n5707), .ZN(n7207) );
  NAND2_X2 U7225 ( .A1(n7207), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8885) );
  NOR2_X1 U7226 ( .A1(n9068), .A2(n8885), .ZN(n5720) );
  INV_X1 U7227 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U7228 ( .A1(n5709), .A2(n6348), .ZN(n5710) );
  NAND2_X1 U7229 ( .A1(n9055), .A2(n6353), .ZN(n5715) );
  INV_X1 U7230 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U7231 ( .A1(n4458), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U7232 ( .A1(n8599), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5711) );
  OAI211_X1 U7233 ( .C1(n5522), .C2(n6666), .A(n5712), .B(n5711), .ZN(n5713)
         );
  INV_X1 U7234 ( .A(n5713), .ZN(n5714) );
  INV_X1 U7235 ( .A(n8799), .ZN(n5716) );
  AND2_X1 U7236 ( .A1(n5717), .A2(n5716), .ZN(n7219) );
  NAND2_X1 U7237 ( .A1(n7219), .A2(n9266), .ZN(n8887) );
  INV_X1 U7238 ( .A(n7219), .ZN(n8570) );
  INV_X1 U7239 ( .A(n8809), .ZN(n5718) );
  OAI22_X1 U7240 ( .A1(n8774), .A2(n8887), .B1(n9072), .B2(n8875), .ZN(n5719)
         );
  AOI211_X1 U7241 ( .C1(P2_REG3_REG_27__SCAN_IN), .C2(P2_U3152), .A(n5720), 
        .B(n5719), .ZN(n5721) );
  INV_X1 U7242 ( .A(n5722), .ZN(n5723) );
  NAND2_X1 U7243 ( .A1(n5724), .A2(n5723), .ZN(P2_U3216) );
  NOR2_X1 U7244 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5728) );
  NOR2_X1 U7245 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5727) );
  NOR2_X1 U7246 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5726) );
  NOR2_X1 U7247 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5725) );
  NAND4_X1 U7248 ( .A1(n5728), .A2(n5727), .A3(n5726), .A4(n5725), .ZN(n5733)
         );
  NOR2_X1 U7249 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5731) );
  NAND4_X1 U7250 ( .A1(n5731), .A2(n5730), .A3(n5945), .A4(n5729), .ZN(n5732)
         );
  NOR2_X1 U7251 ( .A1(n5733), .A2(n5732), .ZN(n5738) );
  NAND2_X1 U7252 ( .A1(n5854), .A2(n5736), .ZN(n5857) );
  INV_X1 U7253 ( .A(n5857), .ZN(n5737) );
  NAND3_X1 U7254 ( .A1(n5742), .A2(n5755), .A3(n5741), .ZN(n5743) );
  XNOR2_X1 U7255 ( .A(n5744), .B(n5769), .ZN(n6301) );
  OAI21_X1 U7256 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5745) );
  NAND2_X1 U7257 ( .A1(n5758), .A2(n5745), .ZN(n5746) );
  XNOR2_X2 U7258 ( .A(n5746), .B(P1_IR_REG_27__SCAN_IN), .ZN(n6461) );
  NAND2_X2 U7259 ( .A1(n6064), .A2(n8228), .ZN(n5878) );
  OR2_X1 U7260 ( .A1(n5878), .A2(n6842), .ZN(n5753) );
  NOR2_X1 U7261 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5749) );
  INV_X1 U7262 ( .A(n5749), .ZN(n5747) );
  NAND2_X1 U7263 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5747), .ZN(n5748) );
  INV_X1 U7264 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5750) );
  MUX2_X1 U7265 ( .A(n5748), .B(P1_IR_REG_31__SCAN_IN), .S(n5750), .Z(n5751)
         );
  NAND2_X1 U7266 ( .A1(n5750), .A2(n5749), .ZN(n5832) );
  INV_X1 U7267 ( .A(n9984), .ZN(n6841) );
  OR2_X1 U7268 ( .A1(n6064), .A2(n6841), .ZN(n5752) );
  AND3_X2 U7269 ( .A1(n5754), .A2(n5753), .A3(n5752), .ZN(n10098) );
  NAND2_X1 U7270 ( .A1(n5758), .A2(n5755), .ZN(n5756) );
  NAND2_X1 U7271 ( .A1(n5756), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5757) );
  XNOR2_X1 U7272 ( .A(n5758), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U7273 ( .A1(n5759), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5760) );
  XNOR2_X1 U7274 ( .A(n5760), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U7275 ( .A1(n5767), .A2(n5768), .ZN(n5762) );
  INV_X1 U7276 ( .A(n5765), .ZN(n5763) );
  NAND2_X1 U7277 ( .A1(n5763), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n5766) );
  INV_X1 U7278 ( .A(n8549), .ZN(n6468) );
  AND2_X4 U7279 ( .A1(n5797), .A2(n5784), .ZN(n6256) );
  INV_X1 U7280 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10163) );
  OR2_X1 U7281 ( .A1(n5871), .A2(n10163), .ZN(n5773) );
  INV_X1 U7282 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5771) );
  OR2_X1 U7283 ( .A1(n5867), .A2(n5771), .ZN(n5772) );
  AND2_X1 U7284 ( .A1(n5773), .A2(n5772), .ZN(n5777) );
  NAND2_X1 U7285 ( .A1(n5788), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5776) );
  NAND2_X2 U7286 ( .A1(n5775), .A2(n5774), .ZN(n6308) );
  INV_X1 U7287 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7293) );
  INV_X1 U7288 ( .A(n5784), .ZN(n7253) );
  NAND2_X1 U7289 ( .A1(n5781), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5782) );
  XNOR2_X2 U7290 ( .A(n5782), .B(P1_IR_REG_19__SCAN_IN), .ZN(n10044) );
  NAND2_X1 U7291 ( .A1(n8549), .A2(n9644), .ZN(n8546) );
  OAI22_X1 U7292 ( .A1(n8556), .A2(n10044), .B1(n8289), .B2(n8546), .ZN(n5783)
         );
  NAND2_X1 U7293 ( .A1(n6300), .A2(n5783), .ZN(n6437) );
  INV_X4 U7294 ( .A(n5842), .ZN(n8200) );
  NAND2_X1 U7295 ( .A1(n8556), .A2(n8289), .ZN(n7244) );
  OR2_X1 U7296 ( .A1(n7244), .A2(n8546), .ZN(n7245) );
  AND2_X4 U7297 ( .A1(n6256), .A2(n7245), .ZN(n6228) );
  NAND2_X1 U7298 ( .A1(n5785), .A2(n6228), .ZN(n5787) );
  OR2_X1 U7299 ( .A1(n10098), .A2(n6265), .ZN(n5786) );
  NAND2_X1 U7300 ( .A1(n5787), .A2(n5786), .ZN(n5828) );
  INV_X1 U7301 ( .A(n7009), .ZN(n5826) );
  INV_X1 U7302 ( .A(n5872), .ZN(n5788) );
  INV_X1 U7303 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9956) );
  OR2_X1 U7304 ( .A1(n5871), .A2(n9956), .ZN(n5791) );
  NAND2_X1 U7305 ( .A1(n5807), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5789) );
  NAND4_X2 U7306 ( .A1(n5792), .A2(n5791), .A3(n5790), .A4(n5789), .ZN(n6441)
         );
  INV_X1 U7307 ( .A(SI_0_), .ZN(n5794) );
  INV_X1 U7308 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5793) );
  OAI21_X1 U7309 ( .B1(n8228), .B2(n5794), .A(n5793), .ZN(n5796) );
  AND2_X1 U7310 ( .A1(n5796), .A2(n5795), .ZN(n9839) );
  MUX2_X1 U7311 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9839), .S(n6064), .Z(n10039)
         );
  NOR2_X1 U7312 ( .A1(n5797), .A2(n9956), .ZN(n5798) );
  AOI21_X1 U7313 ( .B1(n10039), .B2(n6256), .A(n5798), .ZN(n5799) );
  NAND2_X1 U7314 ( .A1(n5800), .A2(n5799), .ZN(n6921) );
  INV_X1 U7315 ( .A(n6921), .ZN(n5801) );
  NAND2_X1 U7316 ( .A1(n5801), .A2(n8200), .ZN(n5806) );
  NAND2_X1 U7317 ( .A1(n6441), .A2(n6228), .ZN(n5805) );
  INV_X1 U7318 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9946) );
  NOR2_X1 U7319 ( .A1(n5797), .A2(n9946), .ZN(n5803) );
  AOI21_X1 U7320 ( .B1(n10039), .B2(n5844), .A(n5803), .ZN(n5804) );
  AND2_X1 U7321 ( .A1(n5805), .A2(n5804), .ZN(n6922) );
  NAND2_X1 U7322 ( .A1(n5806), .A2(n6920), .ZN(n5822) );
  NAND2_X1 U7323 ( .A1(n5807), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5810) );
  AND2_X1 U7324 ( .A1(n5810), .A2(n5809), .ZN(n5812) );
  INV_X1 U7325 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10059) );
  NAND2_X1 U7326 ( .A1(n5884), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U7327 ( .A1(n9499), .A2(n5844), .ZN(n5818) );
  INV_X1 U7328 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6840) );
  OR2_X2 U7329 ( .A1(n5878), .A2(n6840), .ZN(n5815) );
  INV_X1 U7330 ( .A(n9966), .ZN(n6839) );
  OR2_X1 U7331 ( .A1(n6064), .A2(n6839), .ZN(n5814) );
  INV_X1 U7332 ( .A(n10092), .ZN(n5816) );
  NAND2_X1 U7333 ( .A1(n5816), .A2(n6256), .ZN(n5817) );
  NAND2_X1 U7334 ( .A1(n5818), .A2(n5817), .ZN(n5819) );
  XNOR2_X1 U7335 ( .A(n5819), .B(n5842), .ZN(n5823) );
  NAND2_X1 U7336 ( .A1(n5822), .A2(n5823), .ZN(n6941) );
  NAND2_X1 U7337 ( .A1(n9499), .A2(n6228), .ZN(n5821) );
  OR2_X1 U7338 ( .A1(n10092), .A2(n6265), .ZN(n5820) );
  NAND2_X1 U7339 ( .A1(n5821), .A2(n5820), .ZN(n6939) );
  NAND2_X1 U7340 ( .A1(n6941), .A2(n6939), .ZN(n6936) );
  INV_X1 U7341 ( .A(n5822), .ZN(n5825) );
  INV_X1 U7342 ( .A(n5823), .ZN(n5824) );
  NAND2_X1 U7343 ( .A1(n5825), .A2(n5824), .ZN(n6937) );
  AND2_X1 U7344 ( .A1(n6936), .A2(n6937), .ZN(n7010) );
  NAND2_X1 U7345 ( .A1(n5826), .A2(n7010), .ZN(n7011) );
  INV_X1 U7346 ( .A(n5827), .ZN(n5830) );
  INV_X1 U7347 ( .A(n5828), .ZN(n5829) );
  NAND2_X1 U7348 ( .A1(n5830), .A2(n5829), .ZN(n5831) );
  NAND2_X1 U7349 ( .A1(n7011), .A2(n5831), .ZN(n7119) );
  NAND2_X1 U7350 ( .A1(n5832), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5833) );
  XNOR2_X1 U7351 ( .A(n5833), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6796) );
  INV_X1 U7352 ( .A(n6796), .ZN(n6847) );
  OR2_X1 U7353 ( .A1(n5834), .A2(n6849), .ZN(n5836) );
  OR2_X1 U7354 ( .A1(n5878), .A2(n6848), .ZN(n5835) );
  OAI211_X1 U7355 ( .C1(n6064), .C2(n6847), .A(n5836), .B(n5835), .ZN(n10103)
         );
  INV_X1 U7356 ( .A(n10103), .ZN(n7263) );
  NAND2_X1 U7357 ( .A1(n5808), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5841) );
  INV_X1 U7358 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5837) );
  OR2_X1 U7359 ( .A1(n5871), .A2(n5837), .ZN(n5840) );
  INV_X1 U7360 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7262) );
  OR2_X1 U7361 ( .A1(n4448), .A2(n7262), .ZN(n5839) );
  OR2_X1 U7362 ( .A1(n6308), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5838) );
  OAI22_X1 U7363 ( .A1(n7387), .A2(n8202), .B1(n7263), .B2(n5802), .ZN(n5846)
         );
  XNOR2_X1 U7364 ( .A(n5845), .B(n5846), .ZN(n7120) );
  NAND2_X1 U7365 ( .A1(n7119), .A2(n7120), .ZN(n5849) );
  INV_X1 U7366 ( .A(n5845), .ZN(n5847) );
  OR2_X1 U7367 ( .A1(n5847), .A2(n5846), .ZN(n5848) );
  NAND2_X1 U7368 ( .A1(n5849), .A2(n5848), .ZN(n7196) );
  NAND2_X1 U7369 ( .A1(n5808), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5853) );
  INV_X1 U7370 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6797) );
  OR2_X1 U7371 ( .A1(n5871), .A2(n6797), .ZN(n5852) );
  XNOR2_X1 U7372 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7397) );
  OR2_X1 U7373 ( .A1(n6308), .A2(n7397), .ZN(n5851) );
  INV_X1 U7374 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6781) );
  OR2_X1 U7375 ( .A1(n4448), .A2(n6781), .ZN(n5850) );
  NOR2_X1 U7376 ( .A1(n5854), .A2(n9826), .ZN(n5855) );
  MUX2_X1 U7377 ( .A(n9826), .B(n5855), .S(P1_IR_REG_4__SCAN_IN), .Z(n5856) );
  INV_X1 U7378 ( .A(n5856), .ZN(n5858) );
  NAND2_X1 U7379 ( .A1(n5858), .A2(n5892), .ZN(n6851) );
  OR2_X1 U7380 ( .A1(n5878), .A2(n6852), .ZN(n5859) );
  OAI22_X1 U7381 ( .A1(n7364), .A2(n5802), .B1(n10111), .B2(n8199), .ZN(n5860)
         );
  XNOR2_X1 U7382 ( .A(n5860), .B(n6226), .ZN(n5861) );
  OAI22_X1 U7383 ( .A1(n7364), .A2(n8202), .B1(n10111), .B2(n5802), .ZN(n5862)
         );
  XNOR2_X1 U7384 ( .A(n5861), .B(n5862), .ZN(n7197) );
  NAND2_X1 U7385 ( .A1(n7196), .A2(n7197), .ZN(n5865) );
  INV_X1 U7386 ( .A(n5861), .ZN(n5863) );
  OR2_X1 U7387 ( .A1(n5863), .A2(n5862), .ZN(n5864) );
  NAND2_X1 U7388 ( .A1(n5865), .A2(n5864), .ZN(n7360) );
  AOI21_X1 U7389 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5866) );
  NOR2_X1 U7390 ( .A1(n5866), .A2(n5886), .ZN(n7345) );
  NAND2_X1 U7391 ( .A1(n5807), .A2(n7345), .ZN(n5876) );
  INV_X1 U7392 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5869) );
  OR2_X1 U7393 ( .A1(n5868), .A2(n5869), .ZN(n5875) );
  INV_X1 U7394 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5870) );
  OR2_X1 U7395 ( .A1(n5871), .A2(n5870), .ZN(n5874) );
  INV_X1 U7396 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7346) );
  OR2_X1 U7397 ( .A1(n4448), .A2(n7346), .ZN(n5873) );
  OR2_X1 U7398 ( .A1(n7557), .A2(n8202), .ZN(n5882) );
  NAND2_X1 U7399 ( .A1(n5892), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5877) );
  XNOR2_X1 U7400 ( .A(n5877), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6800) );
  INV_X1 U7401 ( .A(n6800), .ZN(n6860) );
  OR2_X1 U7402 ( .A1(n5878), .A2(n6861), .ZN(n5879) );
  OAI211_X1 U7403 ( .C1(n6064), .C2(n6860), .A(n5880), .B(n5879), .ZN(n7351)
         );
  NAND2_X1 U7404 ( .A1(n7351), .A2(n5844), .ZN(n5881) );
  NAND2_X1 U7405 ( .A1(n5882), .A2(n5881), .ZN(n7361) );
  INV_X1 U7406 ( .A(n7351), .ZN(n7367) );
  OAI22_X1 U7407 ( .A1(n7557), .A2(n5802), .B1(n7367), .B2(n8199), .ZN(n5883)
         );
  XNOR2_X1 U7408 ( .A(n5883), .B(n8200), .ZN(n5900) );
  NAND2_X1 U7409 ( .A1(n5788), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5891) );
  INV_X1 U7410 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5885) );
  OR2_X1 U7411 ( .A1(n6460), .A2(n5885), .ZN(n5890) );
  NAND2_X1 U7412 ( .A1(n5886), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5911) );
  OAI21_X1 U7413 ( .B1(n5886), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5911), .ZN(
        n7556) );
  OR2_X1 U7414 ( .A1(n6416), .A2(n7556), .ZN(n5889) );
  INV_X1 U7415 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5887) );
  OR2_X1 U7416 ( .A1(n5868), .A2(n5887), .ZN(n5888) );
  NAND2_X1 U7417 ( .A1(n5906), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5893) );
  XNOR2_X1 U7418 ( .A(n5893), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10011) );
  AOI22_X1 U7419 ( .A1(n6144), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6762), .B2(
        n10011), .ZN(n5895) );
  NAND2_X1 U7420 ( .A1(n5895), .A2(n5894), .ZN(n7547) );
  INV_X1 U7421 ( .A(n7547), .ZN(n7309) );
  OAI22_X1 U7422 ( .A1(n7344), .A2(n5802), .B1(n7309), .B2(n8199), .ZN(n5896)
         );
  XNOR2_X1 U7423 ( .A(n5896), .B(n8200), .ZN(n7551) );
  OR2_X1 U7424 ( .A1(n7344), .A2(n8202), .ZN(n5898) );
  NAND2_X1 U7425 ( .A1(n7547), .A2(n5844), .ZN(n5897) );
  NAND2_X1 U7426 ( .A1(n5898), .A2(n5897), .ZN(n7550) );
  AOI22_X1 U7427 ( .A1(n7361), .A2(n5900), .B1(n7551), .B2(n7550), .ZN(n5899)
         );
  NAND2_X1 U7428 ( .A1(n7360), .A2(n5899), .ZN(n5905) );
  OAI21_X1 U7429 ( .B1(n5900), .B2(n7361), .A(n7550), .ZN(n5903) );
  INV_X1 U7430 ( .A(n7551), .ZN(n5902) );
  INV_X1 U7431 ( .A(n5900), .ZN(n7549) );
  NOR2_X1 U7432 ( .A1(n7361), .A2(n7550), .ZN(n5901) );
  AOI22_X1 U7433 ( .A1(n5903), .A2(n5902), .B1(n7549), .B2(n5901), .ZN(n5904)
         );
  NAND2_X1 U7434 ( .A1(n5905), .A2(n5904), .ZN(n7317) );
  OR2_X1 U7435 ( .A1(n5943), .A2(n9826), .ZN(n5926) );
  XNOR2_X1 U7436 ( .A(n5926), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6867) );
  AOI22_X1 U7437 ( .A1(n6144), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6762), .B2(
        n6867), .ZN(n5907) );
  NAND2_X1 U7438 ( .A1(n5808), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5916) );
  INV_X1 U7439 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5909) );
  AND2_X1 U7440 ( .A1(n5911), .A2(n5910), .ZN(n5912) );
  OR2_X1 U7441 ( .A1(n5912), .A2(n5931), .ZN(n7374) );
  OR2_X1 U7442 ( .A1(n6308), .A2(n7374), .ZN(n5914) );
  INV_X1 U7443 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7375) );
  OR2_X1 U7444 ( .A1(n4448), .A2(n7375), .ZN(n5913) );
  INV_X1 U7445 ( .A(n9493), .ZN(n7543) );
  OAI22_X1 U7446 ( .A1(n10137), .A2(n8199), .B1(n7543), .B2(n5802), .ZN(n5917)
         );
  XNOR2_X1 U7447 ( .A(n5917), .B(n6226), .ZN(n5922) );
  OR2_X1 U7448 ( .A1(n10137), .A2(n5802), .ZN(n5919) );
  NAND2_X1 U7449 ( .A1(n9493), .A2(n6228), .ZN(n5918) );
  NAND2_X1 U7450 ( .A1(n5919), .A2(n5918), .ZN(n5920) );
  XNOR2_X1 U7451 ( .A(n5922), .B(n5920), .ZN(n7318) );
  INV_X1 U7452 ( .A(n5920), .ZN(n5921) );
  NAND2_X1 U7453 ( .A1(n5922), .A2(n5921), .ZN(n5923) );
  NAND2_X1 U7454 ( .A1(n6871), .A2(n8283), .ZN(n5930) );
  INV_X1 U7455 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U7456 ( .A1(n5926), .A2(n5925), .ZN(n5927) );
  NAND2_X1 U7457 ( .A1(n5927), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5928) );
  XNOR2_X1 U7458 ( .A(n5928), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6792) );
  AOI22_X1 U7459 ( .A1(n6144), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6762), .B2(
        n6792), .ZN(n5929) );
  NAND2_X1 U7460 ( .A1(n5930), .A2(n5929), .ZN(n7535) );
  NAND2_X1 U7461 ( .A1(n5808), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5936) );
  INV_X1 U7462 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6803) );
  OR2_X1 U7463 ( .A1(n6460), .A2(n6803), .ZN(n5935) );
  NAND2_X1 U7464 ( .A1(n5931), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5952) );
  OR2_X1 U7465 ( .A1(n5931), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5932) );
  NAND2_X1 U7466 ( .A1(n5952), .A2(n5932), .ZN(n7542) );
  OR2_X1 U7467 ( .A1(n6308), .A2(n7542), .ZN(n5934) );
  INV_X1 U7468 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7482) );
  OR2_X1 U7469 ( .A1(n4448), .A2(n7482), .ZN(n5933) );
  AOI22_X1 U7470 ( .A1(n7535), .A2(n6270), .B1(n10022), .B2(n6228), .ZN(n5940)
         );
  NAND2_X1 U7471 ( .A1(n7535), .A2(n6256), .ZN(n5938) );
  OR2_X1 U7472 ( .A1(n7612), .A2(n5802), .ZN(n5937) );
  NAND2_X1 U7473 ( .A1(n5938), .A2(n5937), .ZN(n5939) );
  XNOR2_X1 U7474 ( .A(n5939), .B(n8200), .ZN(n7538) );
  INV_X1 U7475 ( .A(n5940), .ZN(n5941) );
  NAND2_X1 U7476 ( .A1(n6899), .A2(n8283), .ZN(n5950) );
  NOR2_X1 U7477 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5942) );
  NOR2_X1 U7478 ( .A1(n5946), .A2(n9826), .ZN(n5944) );
  MUX2_X1 U7479 ( .A(n9826), .B(n5944), .S(P1_IR_REG_9__SCAN_IN), .Z(n5948) );
  NAND2_X1 U7480 ( .A1(n5946), .A2(n5945), .ZN(n5984) );
  INV_X1 U7481 ( .A(n5984), .ZN(n5947) );
  AOI22_X1 U7482 ( .A1(n6144), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6762), .B2(
        n7071), .ZN(n5949) );
  NAND2_X1 U7483 ( .A1(n5950), .A2(n5949), .ZN(n10150) );
  NAND2_X1 U7484 ( .A1(n10150), .A2(n6256), .ZN(n5960) );
  NAND2_X1 U7485 ( .A1(n5808), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U7486 ( .A1(n5952), .A2(n5951), .ZN(n5953) );
  NAND2_X1 U7487 ( .A1(n5971), .A2(n5953), .ZN(n10035) );
  OR2_X1 U7488 ( .A1(n6416), .A2(n10035), .ZN(n5957) );
  INV_X1 U7489 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5954) );
  OR2_X1 U7490 ( .A1(n6460), .A2(n5954), .ZN(n5956) );
  INV_X1 U7491 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10018) );
  OR2_X1 U7492 ( .A1(n4448), .A2(n10018), .ZN(n5955) );
  OR2_X1 U7493 ( .A1(n7711), .A2(n5802), .ZN(n5959) );
  NAND2_X1 U7494 ( .A1(n5960), .A2(n5959), .ZN(n5961) );
  XNOR2_X1 U7495 ( .A(n5961), .B(n6226), .ZN(n5966) );
  NOR2_X1 U7496 ( .A1(n7711), .A2(n8202), .ZN(n5962) );
  AOI21_X1 U7497 ( .B1(n10150), .B2(n6270), .A(n5962), .ZN(n5965) );
  XNOR2_X1 U7498 ( .A(n5966), .B(n5965), .ZN(n7611) );
  NAND2_X1 U7499 ( .A1(n5966), .A2(n5965), .ZN(n5967) );
  NAND2_X1 U7500 ( .A1(n5984), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5968) );
  XNOR2_X1 U7501 ( .A(n5968), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7171) );
  AOI22_X1 U7502 ( .A1(n6144), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6762), .B2(
        n7171), .ZN(n5969) );
  NAND2_X1 U7503 ( .A1(n5808), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5976) );
  INV_X1 U7504 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5970) );
  OR2_X1 U7505 ( .A1(n6460), .A2(n5970), .ZN(n5975) );
  INV_X1 U7506 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7695) );
  OR2_X1 U7507 ( .A1(n4448), .A2(n7695), .ZN(n5974) );
  NAND2_X1 U7508 ( .A1(n5971), .A2(n7066), .ZN(n5972) );
  NAND2_X1 U7509 ( .A1(n5990), .A2(n5972), .ZN(n7710) );
  OR2_X1 U7510 ( .A1(n6416), .A2(n7710), .ZN(n5973) );
  OR2_X1 U7511 ( .A1(n7787), .A2(n5802), .ZN(n5977) );
  NAND2_X1 U7512 ( .A1(n5978), .A2(n5977), .ZN(n5979) );
  NOR2_X1 U7513 ( .A1(n7787), .A2(n8202), .ZN(n5980) );
  AOI21_X1 U7514 ( .B1(n7699), .B2(n6270), .A(n5980), .ZN(n5982) );
  INV_X1 U7515 ( .A(n5981), .ZN(n5983) );
  INV_X1 U7516 ( .A(n7723), .ZN(n6001) );
  NAND2_X1 U7517 ( .A1(n6908), .A2(n8283), .ZN(n5987) );
  NAND2_X1 U7518 ( .A1(n6007), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5985) );
  XNOR2_X1 U7519 ( .A(n5985), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7335) );
  AOI22_X1 U7520 ( .A1(n6144), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6762), .B2(
        n7335), .ZN(n5986) );
  NAND2_X1 U7521 ( .A1(n7796), .A2(n6256), .ZN(n5997) );
  NAND2_X1 U7522 ( .A1(n5808), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5995) );
  INV_X1 U7523 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5988) );
  OR2_X1 U7524 ( .A1(n6460), .A2(n5988), .ZN(n5994) );
  AND2_X1 U7525 ( .A1(n5990), .A2(n5989), .ZN(n5991) );
  OR2_X1 U7526 ( .A1(n5991), .A2(n6011), .ZN(n7793) );
  OR2_X1 U7527 ( .A1(n6308), .A2(n7793), .ZN(n5993) );
  INV_X1 U7528 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7794) );
  OR2_X1 U7529 ( .A1(n4448), .A2(n7794), .ZN(n5992) );
  NAND4_X1 U7530 ( .A1(n5995), .A2(n5994), .A3(n5993), .A4(n5992), .ZN(n9491)
         );
  NAND2_X1 U7531 ( .A1(n9491), .A2(n6270), .ZN(n5996) );
  NAND2_X1 U7532 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  XNOR2_X1 U7533 ( .A(n5998), .B(n6226), .ZN(n6002) );
  AND2_X1 U7534 ( .A1(n9491), .A2(n6228), .ZN(n5999) );
  AOI21_X1 U7535 ( .B1(n7796), .B2(n6270), .A(n5999), .ZN(n6003) );
  XNOR2_X1 U7536 ( .A(n6002), .B(n6003), .ZN(n7722) );
  NAND2_X1 U7537 ( .A1(n6001), .A2(n6000), .ZN(n7724) );
  INV_X1 U7538 ( .A(n6002), .ZN(n6005) );
  INV_X1 U7539 ( .A(n6003), .ZN(n6004) );
  NAND2_X1 U7540 ( .A1(n6005), .A2(n6004), .ZN(n6006) );
  NAND2_X1 U7541 ( .A1(n6947), .A2(n8283), .ZN(n6010) );
  OR2_X1 U7542 ( .A1(n6026), .A2(n9826), .ZN(n6008) );
  XNOR2_X1 U7543 ( .A(n6008), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7511) );
  AOI22_X1 U7544 ( .A1(n6144), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6762), .B2(
        n7511), .ZN(n6009) );
  NAND2_X1 U7545 ( .A1(n8028), .A2(n6256), .ZN(n6018) );
  NAND2_X1 U7546 ( .A1(n5808), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6016) );
  INV_X1 U7547 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7329) );
  OR2_X1 U7548 ( .A1(n6460), .A2(n7329), .ZN(n6015) );
  NOR2_X1 U7549 ( .A1(n6011), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6012) );
  OR2_X1 U7550 ( .A1(n6030), .A2(n6012), .ZN(n7891) );
  OR2_X1 U7551 ( .A1(n6308), .A2(n7891), .ZN(n6014) );
  INV_X1 U7552 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7892) );
  OR2_X1 U7553 ( .A1(n4448), .A2(n7892), .ZN(n6013) );
  OR2_X1 U7554 ( .A1(n7912), .A2(n5802), .ZN(n6017) );
  NAND2_X1 U7555 ( .A1(n6018), .A2(n6017), .ZN(n6019) );
  XNOR2_X1 U7556 ( .A(n6019), .B(n8200), .ZN(n7774) );
  INV_X1 U7557 ( .A(n7774), .ZN(n6022) );
  NAND2_X1 U7558 ( .A1(n8028), .A2(n6270), .ZN(n6021) );
  OR2_X1 U7559 ( .A1(n7912), .A2(n8202), .ZN(n6020) );
  NAND2_X1 U7560 ( .A1(n6021), .A2(n6020), .ZN(n6023) );
  INV_X1 U7561 ( .A(n6023), .ZN(n7773) );
  AND2_X1 U7562 ( .A1(n7774), .A2(n6023), .ZN(n6024) );
  NAND2_X1 U7563 ( .A1(n7191), .A2(n8283), .ZN(n6029) );
  INV_X1 U7564 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6025) );
  OR2_X1 U7565 ( .A1(n6044), .A2(n9826), .ZN(n6027) );
  XNOR2_X1 U7566 ( .A(n6027), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7741) );
  AOI22_X1 U7567 ( .A1(n6144), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6762), .B2(
        n7741), .ZN(n6028) );
  NAND2_X1 U7568 ( .A1(n7915), .A2(n6256), .ZN(n6037) );
  NAND2_X1 U7569 ( .A1(n5808), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6035) );
  INV_X1 U7570 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7502) );
  OR2_X1 U7571 ( .A1(n6460), .A2(n7502), .ZN(n6034) );
  OR2_X1 U7572 ( .A1(n6030), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7573 ( .A1(n6031), .A2(n6048), .ZN(n7911) );
  OR2_X1 U7574 ( .A1(n6308), .A2(n7911), .ZN(n6033) );
  INV_X1 U7575 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7812) );
  OR2_X1 U7576 ( .A1(n4448), .A2(n7812), .ZN(n6032) );
  OR2_X1 U7577 ( .A1(n7887), .A2(n5802), .ZN(n6036) );
  NAND2_X1 U7578 ( .A1(n6037), .A2(n6036), .ZN(n6038) );
  XNOR2_X1 U7579 ( .A(n6038), .B(n6226), .ZN(n6041) );
  NOR2_X1 U7580 ( .A1(n7887), .A2(n8202), .ZN(n6039) );
  AOI21_X1 U7581 ( .B1(n7915), .B2(n6270), .A(n6039), .ZN(n6040) );
  OR2_X1 U7582 ( .A1(n6041), .A2(n6040), .ZN(n7908) );
  NAND2_X1 U7583 ( .A1(n6041), .A2(n6040), .ZN(n7907) );
  NAND2_X1 U7584 ( .A1(n7194), .A2(n8283), .ZN(n6046) );
  INV_X1 U7585 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7586 ( .A1(n6044), .A2(n6043), .ZN(n6089) );
  NAND2_X1 U7587 ( .A1(n6089), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6061) );
  XNOR2_X1 U7588 ( .A(n6061), .B(P1_IR_REG_14__SCAN_IN), .ZN(n8000) );
  AOI22_X1 U7589 ( .A1(n8000), .A2(n6762), .B1(n6144), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U7590 ( .A1(n9808), .A2(n6256), .ZN(n6055) );
  NAND2_X1 U7591 ( .A1(n5808), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6053) );
  INV_X1 U7592 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7735) );
  OR2_X1 U7593 ( .A1(n6460), .A2(n7735), .ZN(n6052) );
  INV_X1 U7594 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6047) );
  OR2_X1 U7595 ( .A1(n4448), .A2(n6047), .ZN(n6051) );
  AOI21_X1 U7596 ( .B1(n6716), .B2(n6048), .A(n6068), .ZN(n8129) );
  INV_X1 U7597 ( .A(n8129), .ZN(n6049) );
  OR2_X1 U7598 ( .A1(n6416), .A2(n6049), .ZN(n6050) );
  NAND4_X1 U7599 ( .A1(n6053), .A2(n6052), .A3(n6051), .A4(n6050), .ZN(n9488)
         );
  NAND2_X1 U7600 ( .A1(n9488), .A2(n6270), .ZN(n6054) );
  NAND2_X1 U7601 ( .A1(n6055), .A2(n6054), .ZN(n6056) );
  XNOR2_X1 U7602 ( .A(n6056), .B(n6226), .ZN(n6059) );
  NAND2_X1 U7603 ( .A1(n9808), .A2(n6270), .ZN(n6058) );
  NAND2_X1 U7604 ( .A1(n9488), .A2(n6228), .ZN(n6057) );
  NAND2_X1 U7605 ( .A1(n6058), .A2(n6057), .ZN(n8134) );
  NAND2_X1 U7606 ( .A1(n7324), .A2(n8283), .ZN(n6067) );
  INV_X1 U7607 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7608 ( .A1(n6061), .A2(n6087), .ZN(n6062) );
  NAND2_X1 U7609 ( .A1(n6062), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6063) );
  INV_X1 U7610 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6086) );
  XNOR2_X1 U7611 ( .A(n6063), .B(n6086), .ZN(n8080) );
  OAI22_X1 U7612 ( .A1(n8080), .A2(n6064), .B1(n5878), .B2(n7327), .ZN(n6065)
         );
  INV_X1 U7613 ( .A(n6065), .ZN(n6066) );
  NAND2_X1 U7614 ( .A1(n8046), .A2(n6256), .ZN(n6078) );
  OR2_X1 U7615 ( .A1(n6068), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7616 ( .A1(n6068), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U7617 ( .A1(n6069), .A2(n6093), .ZN(n8069) );
  INV_X1 U7618 ( .A(n8069), .ZN(n6070) );
  NAND2_X1 U7619 ( .A1(n5807), .A2(n6070), .ZN(n6076) );
  INV_X1 U7620 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n6071) );
  OR2_X1 U7621 ( .A1(n5868), .A2(n6071), .ZN(n6075) );
  INV_X1 U7622 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6072) );
  OR2_X1 U7623 ( .A1(n6460), .A2(n6072), .ZN(n6074) );
  INV_X1 U7624 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8040) );
  OR2_X1 U7625 ( .A1(n4448), .A2(n8040), .ZN(n6073) );
  OR2_X1 U7626 ( .A1(n8133), .A2(n6265), .ZN(n6077) );
  NAND2_X1 U7627 ( .A1(n6078), .A2(n6077), .ZN(n6079) );
  XNOR2_X1 U7628 ( .A(n6079), .B(n6226), .ZN(n8065) );
  NOR2_X1 U7629 ( .A1(n8133), .A2(n8202), .ZN(n6080) );
  AOI21_X1 U7630 ( .B1(n8046), .B2(n6270), .A(n6080), .ZN(n8064) );
  NAND2_X1 U7631 ( .A1(n8065), .A2(n8064), .ZN(n6081) );
  NAND2_X1 U7632 ( .A1(n8063), .A2(n6081), .ZN(n6085) );
  INV_X1 U7633 ( .A(n8065), .ZN(n6083) );
  INV_X1 U7634 ( .A(n8064), .ZN(n6082) );
  NAND2_X1 U7635 ( .A1(n6083), .A2(n6082), .ZN(n6084) );
  INV_X1 U7636 ( .A(n8118), .ZN(n6104) );
  NAND2_X1 U7637 ( .A1(n7358), .A2(n8283), .ZN(n6092) );
  NAND2_X1 U7638 ( .A1(n6087), .A2(n6086), .ZN(n6088) );
  NAND2_X1 U7639 ( .A1(n6109), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6090) );
  XNOR2_X1 U7640 ( .A(n6090), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9518) );
  AOI22_X1 U7641 ( .A1(n9518), .A2(n6762), .B1(n6144), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7642 ( .A1(n8060), .A2(n6256), .ZN(n6099) );
  AOI21_X1 U7643 ( .B1(n8086), .B2(n6093), .A(n6112), .ZN(n8055) );
  NAND2_X1 U7644 ( .A1(n8055), .A2(n5807), .ZN(n6097) );
  NAND2_X1 U7645 ( .A1(n5808), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U7646 ( .A1(n5884), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7647 ( .A1(n5788), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6094) );
  OR2_X1 U7648 ( .A1(n9427), .A2(n5802), .ZN(n6098) );
  NAND2_X1 U7649 ( .A1(n6099), .A2(n6098), .ZN(n6100) );
  XNOR2_X1 U7650 ( .A(n6100), .B(n8200), .ZN(n6105) );
  NAND2_X1 U7651 ( .A1(n8060), .A2(n6270), .ZN(n6102) );
  OR2_X1 U7652 ( .A1(n9427), .A2(n8202), .ZN(n6101) );
  NAND2_X1 U7653 ( .A1(n6102), .A2(n6101), .ZN(n6106) );
  AND2_X1 U7654 ( .A1(n6105), .A2(n6106), .ZN(n8119) );
  INV_X1 U7655 ( .A(n8119), .ZN(n6103) );
  INV_X1 U7656 ( .A(n6105), .ZN(n6108) );
  INV_X1 U7657 ( .A(n6106), .ZN(n6107) );
  NAND2_X1 U7658 ( .A1(n6108), .A2(n6107), .ZN(n8120) );
  NAND2_X1 U7659 ( .A1(n7404), .A2(n8283), .ZN(n6111) );
  OAI21_X1 U7660 ( .B1(n6109), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6126) );
  XNOR2_X1 U7661 ( .A(n6126), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9537) );
  AOI22_X1 U7662 ( .A1(n9537), .A2(n6762), .B1(n6144), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U7663 ( .A1(n9740), .A2(n6256), .ZN(n6119) );
  OR2_X1 U7664 ( .A1(n6112), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7665 ( .A1(n6112), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7666 ( .A1(n6113), .A2(n6132), .ZN(n9734) );
  INV_X1 U7667 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9519) );
  NAND2_X1 U7668 ( .A1(n5808), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7669 ( .A1(n5788), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6114) );
  OAI211_X1 U7670 ( .C1(n6460), .C2(n9519), .A(n6115), .B(n6114), .ZN(n6116)
         );
  INV_X1 U7671 ( .A(n6116), .ZN(n6117) );
  OAI21_X1 U7672 ( .B1(n9734), .B2(n6416), .A(n6117), .ZN(n9486) );
  NAND2_X1 U7673 ( .A1(n9486), .A2(n6270), .ZN(n6118) );
  NAND2_X1 U7674 ( .A1(n6119), .A2(n6118), .ZN(n6120) );
  XNOR2_X1 U7675 ( .A(n6120), .B(n8200), .ZN(n6122) );
  AND2_X1 U7676 ( .A1(n9486), .A2(n6228), .ZN(n6121) );
  AOI21_X1 U7677 ( .B1(n9740), .B2(n6270), .A(n6121), .ZN(n6123) );
  XNOR2_X1 U7678 ( .A(n6122), .B(n6123), .ZN(n9426) );
  INV_X1 U7679 ( .A(n6122), .ZN(n6124) );
  NAND2_X1 U7680 ( .A1(n7606), .A2(n8283), .ZN(n6131) );
  INV_X1 U7681 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6125) );
  NAND2_X1 U7682 ( .A1(n6126), .A2(n6125), .ZN(n6127) );
  NAND2_X1 U7683 ( .A1(n6127), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6128) );
  XNOR2_X1 U7684 ( .A(n6128), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9548) );
  INV_X1 U7685 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7638) );
  NOR2_X1 U7686 ( .A1(n5878), .A2(n7638), .ZN(n6129) );
  AOI21_X1 U7687 ( .B1(n9548), .B2(n6762), .A(n6129), .ZN(n6130) );
  NAND2_X1 U7688 ( .A1(n9803), .A2(n6256), .ZN(n6139) );
  NAND2_X1 U7689 ( .A1(n5808), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6137) );
  INV_X1 U7690 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9530) );
  OR2_X1 U7691 ( .A1(n6460), .A2(n9530), .ZN(n6136) );
  OAI21_X1 U7692 ( .B1(P1_REG3_REG_18__SCAN_IN), .B2(n6133), .A(n6148), .ZN(
        n9471) );
  OR2_X1 U7693 ( .A1(n6308), .A2(n9471), .ZN(n6135) );
  INV_X1 U7694 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8109) );
  OR2_X1 U7695 ( .A1(n4448), .A2(n8109), .ZN(n6134) );
  OR2_X1 U7696 ( .A1(n9717), .A2(n5802), .ZN(n6138) );
  NAND2_X1 U7697 ( .A1(n6139), .A2(n6138), .ZN(n6140) );
  XNOR2_X1 U7698 ( .A(n6140), .B(n8200), .ZN(n6142) );
  NOR2_X1 U7699 ( .A1(n9717), .A2(n8202), .ZN(n6141) );
  AOI21_X1 U7700 ( .B1(n9803), .B2(n6270), .A(n6141), .ZN(n9464) );
  NOR2_X1 U7701 ( .A1(n9465), .A2(n9464), .ZN(n9463) );
  AND2_X2 U7702 ( .A1(n6143), .A2(n6142), .ZN(n9468) );
  NAND2_X1 U7703 ( .A1(n7703), .A2(n8283), .ZN(n6146) );
  AOI22_X1 U7704 ( .A1(n6144), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10044), 
        .B2(n6762), .ZN(n6145) );
  NAND2_X2 U7705 ( .A1(n6146), .A2(n6145), .ZN(n9798) );
  NAND2_X1 U7706 ( .A1(n5884), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6152) );
  INV_X1 U7707 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n6147) );
  OR2_X1 U7708 ( .A1(n4448), .A2(n6147), .ZN(n6151) );
  INV_X1 U7709 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n6664) );
  OR2_X1 U7710 ( .A1(n5868), .A2(n6664), .ZN(n6150) );
  INV_X1 U7711 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9404) );
  AOI21_X1 U7712 ( .B1(n6148), .B2(n9404), .A(n6157), .ZN(n9721) );
  INV_X1 U7713 ( .A(n9721), .ZN(n9405) );
  OR2_X1 U7714 ( .A1(n6416), .A2(n9405), .ZN(n6149) );
  INV_X1 U7715 ( .A(n9708), .ZN(n9485) );
  AOI22_X1 U7716 ( .A1(n9798), .A2(n6256), .B1(n6270), .B2(n9485), .ZN(n6153)
         );
  AOI22_X1 U7717 ( .A1(n9798), .A2(n6270), .B1(n6228), .B2(n9485), .ZN(n9401)
         );
  NAND2_X1 U7718 ( .A1(n7731), .A2(n8283), .ZN(n6155) );
  OR2_X1 U7719 ( .A1(n5878), .A2(n7732), .ZN(n6154) );
  NAND2_X1 U7720 ( .A1(n9793), .A2(n6256), .ZN(n6163) );
  NAND2_X1 U7721 ( .A1(n5884), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6161) );
  INV_X1 U7722 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n6156) );
  OR2_X1 U7723 ( .A1(n5868), .A2(n6156), .ZN(n6160) );
  NAND2_X1 U7724 ( .A1(n6157), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6173) );
  OAI21_X1 U7725 ( .B1(P1_REG3_REG_20__SCAN_IN), .B2(n6157), .A(n6173), .ZN(
        n9700) );
  OR2_X1 U7726 ( .A1(n6308), .A2(n9700), .ZN(n6159) );
  INV_X1 U7727 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9701) );
  OR2_X1 U7728 ( .A1(n4448), .A2(n9701), .ZN(n6158) );
  NAND4_X1 U7729 ( .A1(n6161), .A2(n6160), .A3(n6159), .A4(n6158), .ZN(n9484)
         );
  NAND2_X1 U7730 ( .A1(n9484), .A2(n6270), .ZN(n6162) );
  NAND2_X1 U7731 ( .A1(n6163), .A2(n6162), .ZN(n6164) );
  XNOR2_X1 U7732 ( .A(n6164), .B(n6226), .ZN(n6167) );
  AND2_X1 U7733 ( .A1(n9484), .A2(n6228), .ZN(n6165) );
  AOI21_X1 U7734 ( .B1(n9793), .B2(n6270), .A(n6165), .ZN(n6166) );
  NAND2_X1 U7735 ( .A1(n6167), .A2(n6166), .ZN(n6168) );
  OAI21_X1 U7736 ( .B1(n6167), .B2(n6166), .A(n6168), .ZN(n9445) );
  INV_X1 U7737 ( .A(n6168), .ZN(n6169) );
  NAND2_X1 U7738 ( .A1(n7782), .A2(n8283), .ZN(n6171) );
  OR2_X1 U7739 ( .A1(n5878), .A2(n7783), .ZN(n6170) );
  NAND2_X1 U7740 ( .A1(n9788), .A2(n6256), .ZN(n6181) );
  NAND2_X1 U7741 ( .A1(n5808), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6179) );
  INV_X1 U7742 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6728) );
  OR2_X1 U7743 ( .A1(n6460), .A2(n6728), .ZN(n6178) );
  INV_X1 U7744 ( .A(n6173), .ZN(n6172) );
  INV_X1 U7745 ( .A(n6189), .ZN(n6190) );
  INV_X1 U7746 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9412) );
  NAND2_X1 U7747 ( .A1(n9412), .A2(n6173), .ZN(n6174) );
  NAND2_X1 U7748 ( .A1(n6190), .A2(n6174), .ZN(n9691) );
  OR2_X1 U7749 ( .A1(n6416), .A2(n9691), .ZN(n6177) );
  INV_X1 U7750 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n6175) );
  OR2_X1 U7751 ( .A1(n4448), .A2(n6175), .ZN(n6176) );
  NAND4_X1 U7752 ( .A1(n6179), .A2(n6178), .A3(n6177), .A4(n6176), .ZN(n9678)
         );
  NAND2_X1 U7753 ( .A1(n9678), .A2(n6270), .ZN(n6180) );
  NAND2_X1 U7754 ( .A1(n6181), .A2(n6180), .ZN(n6182) );
  XNOR2_X1 U7755 ( .A(n6182), .B(n8200), .ZN(n6183) );
  INV_X1 U7756 ( .A(n9788), .ZN(n6467) );
  INV_X1 U7757 ( .A(n9678), .ZN(n9707) );
  OAI22_X1 U7758 ( .A1(n6467), .A2(n6265), .B1(n9707), .B2(n8202), .ZN(n6184)
         );
  XNOR2_X1 U7759 ( .A(n6183), .B(n6184), .ZN(n9410) );
  INV_X1 U7760 ( .A(n6183), .ZN(n6186) );
  INV_X1 U7761 ( .A(n6184), .ZN(n6185) );
  NAND2_X1 U7762 ( .A1(n7877), .A2(n8283), .ZN(n6188) );
  OR2_X1 U7763 ( .A1(n5878), .A2(n7878), .ZN(n6187) );
  INV_X1 U7764 ( .A(n9781), .ZN(n9674) );
  NAND2_X1 U7765 ( .A1(n5808), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6196) );
  INV_X1 U7766 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6571) );
  OR2_X1 U7767 ( .A1(n6460), .A2(n6571), .ZN(n6195) );
  INV_X1 U7768 ( .A(n6205), .ZN(n6206) );
  INV_X1 U7769 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9454) );
  NAND2_X1 U7770 ( .A1(n6190), .A2(n9454), .ZN(n6191) );
  NAND2_X1 U7771 ( .A1(n6206), .A2(n6191), .ZN(n9671) );
  OR2_X1 U7772 ( .A1(n6308), .A2(n9671), .ZN(n6194) );
  INV_X1 U7773 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n6192) );
  OR2_X1 U7774 ( .A1(n4448), .A2(n6192), .ZN(n6193) );
  NAND4_X1 U7775 ( .A1(n6196), .A2(n6195), .A3(n6194), .A4(n6193), .ZN(n9663)
         );
  INV_X1 U7776 ( .A(n9663), .ZN(n9688) );
  OAI22_X1 U7777 ( .A1(n9674), .A2(n5802), .B1(n9688), .B2(n8202), .ZN(n6200)
         );
  NAND2_X1 U7778 ( .A1(n9781), .A2(n6256), .ZN(n6198) );
  NAND2_X1 U7779 ( .A1(n9663), .A2(n6270), .ZN(n6197) );
  NAND2_X1 U7780 ( .A1(n6198), .A2(n6197), .ZN(n6199) );
  XNOR2_X1 U7781 ( .A(n6199), .B(n6226), .ZN(n9452) );
  NAND2_X1 U7782 ( .A1(n9451), .A2(n9452), .ZN(n6202) );
  NAND2_X1 U7783 ( .A1(n6202), .A2(n5023), .ZN(n6235) );
  NAND2_X1 U7784 ( .A1(n7989), .A2(n8283), .ZN(n6204) );
  OR2_X1 U7785 ( .A1(n5878), .A2(n7993), .ZN(n6203) );
  NAND2_X1 U7786 ( .A1(n5884), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6213) );
  INV_X1 U7787 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n6740) );
  OR2_X1 U7788 ( .A1(n5868), .A2(n6740), .ZN(n6212) );
  INV_X1 U7789 ( .A(n6219), .ZN(n6208) );
  INV_X1 U7790 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9396) );
  NAND2_X1 U7791 ( .A1(n6206), .A2(n9396), .ZN(n6207) );
  NAND2_X1 U7792 ( .A1(n6208), .A2(n6207), .ZN(n9656) );
  OR2_X1 U7793 ( .A1(n6416), .A2(n9656), .ZN(n6211) );
  INV_X1 U7794 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6209) );
  OR2_X1 U7795 ( .A1(n4448), .A2(n6209), .ZN(n6210) );
  AOI22_X1 U7796 ( .A1(n9776), .A2(n6256), .B1(n6270), .B2(n9677), .ZN(n6214)
         );
  XOR2_X1 U7797 ( .A(n8200), .B(n6214), .Z(n6236) );
  INV_X1 U7798 ( .A(n6236), .ZN(n6215) );
  NAND2_X1 U7799 ( .A1(n6235), .A2(n6215), .ZN(n9392) );
  INV_X1 U7800 ( .A(n9776), .ZN(n9659) );
  OAI22_X1 U7801 ( .A1(n9659), .A2(n6265), .B1(n9456), .B2(n8202), .ZN(n9393)
         );
  NAND2_X1 U7802 ( .A1(n9392), .A2(n9393), .ZN(n9435) );
  NAND2_X1 U7803 ( .A1(n8020), .A2(n8283), .ZN(n6217) );
  OR2_X1 U7804 ( .A1(n5878), .A2(n8021), .ZN(n6216) );
  NAND2_X1 U7805 ( .A1(n9772), .A2(n6256), .ZN(n6225) );
  NAND2_X1 U7806 ( .A1(n5808), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6223) );
  INV_X1 U7807 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6218) );
  OR2_X1 U7808 ( .A1(n6460), .A2(n6218), .ZN(n6222) );
  OAI21_X1 U7809 ( .B1(n6219), .B2(P1_REG3_REG_24__SCAN_IN), .A(n6241), .ZN(
        n9646) );
  OR2_X1 U7810 ( .A1(n6308), .A2(n9646), .ZN(n6221) );
  INV_X1 U7811 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9647) );
  OR2_X1 U7812 ( .A1(n4448), .A2(n9647), .ZN(n6220) );
  NAND4_X1 U7813 ( .A1(n6223), .A2(n6222), .A3(n6221), .A4(n6220), .ZN(n9662)
         );
  NAND2_X1 U7814 ( .A1(n9662), .A2(n6270), .ZN(n6224) );
  NAND2_X1 U7815 ( .A1(n6225), .A2(n6224), .ZN(n6227) );
  XNOR2_X1 U7816 ( .A(n6227), .B(n6226), .ZN(n6230) );
  AND2_X1 U7817 ( .A1(n9662), .A2(n6228), .ZN(n6229) );
  AOI21_X1 U7818 ( .B1(n9772), .B2(n6270), .A(n6229), .ZN(n6231) );
  NAND2_X1 U7819 ( .A1(n6230), .A2(n6231), .ZN(n6238) );
  INV_X1 U7820 ( .A(n6230), .ZN(n6233) );
  INV_X1 U7821 ( .A(n6231), .ZN(n6232) );
  NAND2_X1 U7822 ( .A1(n6233), .A2(n6232), .ZN(n6234) );
  AND2_X1 U7823 ( .A1(n6238), .A2(n6234), .ZN(n9434) );
  INV_X1 U7824 ( .A(n6235), .ZN(n6237) );
  NAND2_X1 U7825 ( .A1(n6237), .A2(n6236), .ZN(n9391) );
  NAND3_X1 U7826 ( .A1(n9435), .A2(n9434), .A3(n9391), .ZN(n9433) );
  NAND2_X1 U7827 ( .A1(n9433), .A2(n6238), .ZN(n9417) );
  NAND2_X1 U7828 ( .A1(n8150), .A2(n8283), .ZN(n6240) );
  OR2_X1 U7829 ( .A1(n5878), .A2(n8156), .ZN(n6239) );
  INV_X1 U7830 ( .A(n9768), .ZN(n9624) );
  NAND2_X1 U7831 ( .A1(n5884), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6246) );
  INV_X1 U7832 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n6732) );
  OR2_X1 U7833 ( .A1(n5868), .A2(n6732), .ZN(n6245) );
  NAND2_X1 U7834 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n6242), .ZN(n6259) );
  OAI21_X1 U7835 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n6242), .A(n6259), .ZN(
        n9625) );
  OR2_X1 U7836 ( .A1(n6308), .A2(n9625), .ZN(n6244) );
  INV_X1 U7837 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9626) );
  OR2_X1 U7838 ( .A1(n4448), .A2(n9626), .ZN(n6243) );
  OAI22_X1 U7839 ( .A1(n9624), .A2(n6265), .B1(n9438), .B2(n8202), .ZN(n6251)
         );
  NAND2_X1 U7840 ( .A1(n9768), .A2(n6256), .ZN(n6248) );
  OR2_X1 U7841 ( .A1(n9438), .A2(n6265), .ZN(n6247) );
  NAND2_X1 U7842 ( .A1(n6248), .A2(n6247), .ZN(n6249) );
  XNOR2_X1 U7843 ( .A(n6249), .B(n8200), .ZN(n6250) );
  XOR2_X1 U7844 ( .A(n6251), .B(n6250), .Z(n9418) );
  INV_X1 U7845 ( .A(n6250), .ZN(n6253) );
  INV_X1 U7846 ( .A(n6251), .ZN(n6252) );
  NAND2_X1 U7847 ( .A1(n6253), .A2(n6252), .ZN(n6272) );
  AND2_X1 U7848 ( .A1(n6275), .A2(n6272), .ZN(n6271) );
  NAND2_X1 U7849 ( .A1(n8157), .A2(n8283), .ZN(n6255) );
  OR2_X1 U7850 ( .A1(n5878), .A2(n8159), .ZN(n6254) );
  NAND2_X1 U7851 ( .A1(n9761), .A2(n6256), .ZN(n6267) );
  NAND2_X1 U7852 ( .A1(n5884), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6264) );
  INV_X1 U7853 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n6257) );
  OR2_X1 U7854 ( .A1(n5868), .A2(n6257), .ZN(n6263) );
  INV_X1 U7855 ( .A(n6259), .ZN(n6258) );
  NAND2_X1 U7856 ( .A1(n6258), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6306) );
  INV_X1 U7857 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U7858 ( .A1(n6319), .A2(n6259), .ZN(n6260) );
  NAND2_X1 U7859 ( .A1(n6306), .A2(n6260), .ZN(n9615) );
  INV_X1 U7860 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9616) );
  OR2_X1 U7861 ( .A1(n4448), .A2(n9616), .ZN(n6261) );
  OR2_X1 U7862 ( .A1(n9634), .A2(n6265), .ZN(n6266) );
  NAND2_X1 U7863 ( .A1(n6267), .A2(n6266), .ZN(n6268) );
  XNOR2_X1 U7864 ( .A(n6268), .B(n8200), .ZN(n8194) );
  NOR2_X1 U7865 ( .A1(n9634), .A2(n8202), .ZN(n6269) );
  AOI21_X1 U7866 ( .B1(n9761), .B2(n6270), .A(n6269), .ZN(n8195) );
  XNOR2_X1 U7867 ( .A(n8194), .B(n8195), .ZN(n6273) );
  INV_X1 U7868 ( .A(n6277), .ZN(n8022) );
  INV_X1 U7869 ( .A(n6280), .ZN(n8154) );
  NAND3_X1 U7870 ( .A1(n8154), .A2(P1_B_REG_SCAN_IN), .A3(n8022), .ZN(n6276)
         );
  OAI211_X1 U7871 ( .C1(P1_B_REG_SCAN_IN), .C2(n8022), .A(n8158), .B(n6276), 
        .ZN(n6469) );
  OR2_X1 U7872 ( .A1(n6469), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6279) );
  OR2_X1 U7873 ( .A1(n8158), .A2(n6277), .ZN(n6278) );
  NAND2_X1 U7874 ( .A1(n6279), .A2(n6278), .ZN(n6929) );
  INV_X1 U7875 ( .A(n6929), .ZN(n6857) );
  OR2_X1 U7876 ( .A1(n6469), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6282) );
  OR2_X1 U7877 ( .A1(n8158), .A2(n6280), .ZN(n6281) );
  NAND2_X1 U7878 ( .A1(n6282), .A2(n6281), .ZN(n6475) );
  INV_X1 U7879 ( .A(n6475), .ZN(n7242) );
  NOR4_X1 U7880 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6291) );
  NOR4_X1 U7881 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6290) );
  INV_X1 U7882 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10075) );
  INV_X1 U7883 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10060) );
  INV_X1 U7884 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10076) );
  INV_X1 U7885 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10080) );
  NAND4_X1 U7886 ( .A1(n10075), .A2(n10060), .A3(n10076), .A4(n10080), .ZN(
        n6288) );
  NOR4_X1 U7887 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6286) );
  NOR4_X1 U7888 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6285) );
  NOR4_X1 U7889 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6284) );
  NOR4_X1 U7890 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6283) );
  NAND4_X1 U7891 ( .A1(n6286), .A2(n6285), .A3(n6284), .A4(n6283), .ZN(n6287)
         );
  NOR4_X1 U7892 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6288), .A4(n6287), .ZN(n6289) );
  AND3_X1 U7893 ( .A1(n6291), .A2(n6290), .A3(n6289), .ZN(n6470) );
  OR2_X1 U7894 ( .A1(n6469), .A2(n6470), .ZN(n6926) );
  NAND3_X1 U7895 ( .A1(n6857), .A2(n7242), .A3(n6926), .ZN(n6313) );
  NAND2_X1 U7896 ( .A1(n6292), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6294) );
  INV_X1 U7897 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6293) );
  XNOR2_X1 U7898 ( .A(n6294), .B(n6293), .ZN(n7990) );
  INV_X1 U7899 ( .A(n6928), .ZN(n6472) );
  OR2_X1 U7900 ( .A1(n6313), .A2(n6472), .ZN(n6299) );
  INV_X1 U7901 ( .A(n6299), .ZN(n6296) );
  INV_X1 U7902 ( .A(n7244), .ZN(n6931) );
  NAND2_X1 U7903 ( .A1(n9384), .A2(n9467), .ZN(n6324) );
  INV_X1 U7904 ( .A(n9761), .ZN(n9614) );
  NAND2_X1 U7905 ( .A1(n10133), .A2(n8289), .ZN(n6474) );
  INV_X1 U7906 ( .A(n6474), .ZN(n6298) );
  NAND2_X2 U7907 ( .A1(n6298), .A2(n6928), .ZN(n10036) );
  NAND2_X1 U7908 ( .A1(n6299), .A2(n10036), .ZN(n9430) );
  INV_X1 U7909 ( .A(n9459), .ZN(n9478) );
  NOR2_X1 U7910 ( .A1(n9614), .A2(n9478), .ZN(n6322) );
  INV_X1 U7911 ( .A(n6300), .ZN(n6932) );
  NAND2_X1 U7912 ( .A1(n6928), .A2(n6932), .ZN(n8560) );
  NOR2_X1 U7913 ( .A1(n6313), .A2(n8560), .ZN(n6318) );
  NAND2_X1 U7914 ( .A1(n6318), .A2(n6302), .ZN(n9473) );
  NAND2_X1 U7915 ( .A1(n5808), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6312) );
  INV_X1 U7916 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6303) );
  OR2_X1 U7917 ( .A1(n6460), .A2(n6303), .ZN(n6311) );
  INV_X1 U7918 ( .A(n6306), .ZN(n6304) );
  NAND2_X1 U7919 ( .A1(n6304), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6414) );
  INV_X1 U7920 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U7921 ( .A1(n6306), .A2(n6305), .ZN(n6307) );
  NAND2_X1 U7922 ( .A1(n6414), .A2(n6307), .ZN(n9599) );
  OR2_X1 U7923 ( .A1(n6308), .A2(n9599), .ZN(n6310) );
  INV_X1 U7924 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9600) );
  OR2_X1 U7925 ( .A1(n4448), .A2(n9600), .ZN(n6309) );
  NAND2_X1 U7926 ( .A1(n6313), .A2(n6474), .ZN(n6316) );
  NAND2_X1 U7927 ( .A1(n5797), .A2(n7990), .ZN(n6314) );
  NOR2_X1 U7928 ( .A1(n6314), .A2(n6925), .ZN(n6315) );
  NAND2_X1 U7929 ( .A1(n6316), .A2(n6315), .ZN(n6317) );
  OAI22_X1 U7930 ( .A1(n9473), .A2(n9575), .B1(n9472), .B2(n9615), .ZN(n6321)
         );
  INV_X1 U7931 ( .A(n6302), .ZN(n6788) );
  OAI22_X1 U7932 ( .A1(n9455), .A2(n9438), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6319), .ZN(n6320) );
  OAI21_X1 U7933 ( .B1(n6325), .B2(n6324), .A(n6323), .ZN(P1_U3238) );
  AOI211_X1 U7934 ( .C1(n6327), .C2(n6326), .A(n8868), .B(n4482), .ZN(n6328)
         );
  INV_X1 U7935 ( .A(n6328), .ZN(n6333) );
  INV_X1 U7936 ( .A(n9301), .ZN(n8211) );
  OAI22_X1 U7937 ( .A1(n8885), .A2(n9106), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6550), .ZN(n6329) );
  INV_X1 U7938 ( .A(n6329), .ZN(n6332) );
  INV_X1 U7939 ( .A(n9136), .ZN(n8847) );
  OAI22_X1 U7940 ( .A1(n9072), .A2(n8887), .B1(n8875), .B2(n8847), .ZN(n6330)
         );
  INV_X1 U7941 ( .A(n6330), .ZN(n6331) );
  NAND4_X1 U7942 ( .A1(n6333), .A2(n5018), .A3(n6332), .A4(n6331), .ZN(
        P2_U3227) );
  INV_X1 U7943 ( .A(n6360), .ZN(n6343) );
  NAND2_X1 U7944 ( .A1(n6335), .A2(n6334), .ZN(n6337) );
  MUX2_X1 U7945 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n4445), .Z(n6424) );
  INV_X1 U7946 ( .A(SI_28_), .ZN(n6568) );
  XNOR2_X1 U7947 ( .A(n6424), .B(n6568), .ZN(n6422) );
  NAND2_X1 U7948 ( .A1(n6409), .A2(n8233), .ZN(n6339) );
  INV_X1 U7949 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8808) );
  OR2_X1 U7950 ( .A1(n8234), .A2(n8808), .ZN(n6338) );
  NOR2_X1 U7951 ( .A1(n8774), .A2(n6340), .ZN(n6341) );
  XNOR2_X1 U7952 ( .A(n6341), .B(n5608), .ZN(n6342) );
  XNOR2_X1 U7953 ( .A(n8596), .B(n6342), .ZN(n6346) );
  NAND3_X1 U7954 ( .A1(n6343), .A2(n8882), .A3(n6346), .ZN(n6362) );
  INV_X1 U7955 ( .A(n6346), .ZN(n6344) );
  INV_X1 U7956 ( .A(n6345), .ZN(n6347) );
  NAND3_X1 U7957 ( .A1(n6347), .A2(n8882), .A3(n6346), .ZN(n6358) );
  INV_X1 U7958 ( .A(n9055), .ZN(n6349) );
  OAI22_X1 U7959 ( .A1(n6349), .A2(n8885), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6348), .ZN(n6356) );
  INV_X1 U7960 ( .A(n9045), .ZN(n6354) );
  INV_X1 U7961 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n9044) );
  NAND2_X1 U7962 ( .A1(n4460), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6351) );
  NAND2_X1 U7963 ( .A1(n4459), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6350) );
  OAI211_X1 U7964 ( .C1(n9044), .C2(n4447), .A(n6351), .B(n6350), .ZN(n6352)
         );
  AOI21_X1 U7965 ( .B1(n6354), .B2(n6353), .A(n6352), .ZN(n8899) );
  OAI22_X1 U7966 ( .A1(n8899), .A2(n8887), .B1(n9031), .B2(n8875), .ZN(n6355)
         );
  AOI211_X1 U7967 ( .C1(n8596), .C2(n8890), .A(n6356), .B(n6355), .ZN(n6357)
         );
  AOI21_X1 U7968 ( .B1(n6360), .B2(n5024), .A(n6359), .ZN(n6361) );
  NAND2_X1 U7969 ( .A1(n6362), .A2(n6361), .ZN(P2_U3222) );
  INV_X1 U7970 ( .A(n8892), .ZN(n8857) );
  INV_X1 U7971 ( .A(n8851), .ZN(n9120) );
  NAND3_X1 U7972 ( .A1(n6363), .A2(n8857), .A3(n9120), .ZN(n6367) );
  OAI21_X1 U7973 ( .B1(n4482), .B2(n6364), .A(n8882), .ZN(n6366) );
  AOI21_X1 U7974 ( .B1(n6367), .B2(n6366), .A(n6365), .ZN(n6374) );
  INV_X1 U7975 ( .A(n6368), .ZN(n9084) );
  OAI22_X1 U7976 ( .A1(n9031), .A2(n9231), .B1(n8851), .B2(n9233), .ZN(n9089)
         );
  AOI22_X1 U7977 ( .A1(n9089), .A2(n7219), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n6369) );
  OAI21_X1 U7978 ( .B1(n8885), .B2(n9084), .A(n6369), .ZN(n6370) );
  INV_X1 U7979 ( .A(n6370), .ZN(n6371) );
  NAND2_X1 U7980 ( .A1(n6441), .A2(n10039), .ZN(n10038) );
  XNOR2_X1 U7981 ( .A(n5785), .B(n10098), .ZN(n6443) );
  NAND2_X1 U7982 ( .A1(n7287), .A2(n6443), .ZN(n6379) );
  INV_X1 U7983 ( .A(n5785), .ZN(n8504) );
  NAND2_X1 U7984 ( .A1(n8504), .A2(n10098), .ZN(n6378) );
  NAND2_X1 U7985 ( .A1(n6379), .A2(n6378), .ZN(n7252) );
  INV_X1 U7986 ( .A(n7387), .ZN(n9498) );
  NAND2_X1 U7987 ( .A1(n9498), .A2(n7263), .ZN(n8307) );
  NAND2_X1 U7988 ( .A1(n7387), .A2(n10103), .ZN(n8509) );
  NAND2_X1 U7989 ( .A1(n7252), .A2(n7255), .ZN(n6381) );
  NAND2_X1 U7990 ( .A1(n7387), .A2(n7263), .ZN(n6380) );
  NAND2_X1 U7991 ( .A1(n6381), .A2(n6380), .ZN(n7390) );
  NAND2_X1 U7992 ( .A1(n7364), .A2(n7399), .ZN(n8511) );
  INV_X1 U7993 ( .A(n7364), .ZN(n9497) );
  NAND2_X1 U7994 ( .A1(n9497), .A2(n10111), .ZN(n8310) );
  NAND2_X1 U7995 ( .A1(n8511), .A2(n8310), .ZN(n8255) );
  NAND2_X1 U7996 ( .A1(n7364), .A2(n10111), .ZN(n6382) );
  NAND2_X1 U7997 ( .A1(n7557), .A2(n7351), .ZN(n8353) );
  NAND2_X1 U7998 ( .A1(n9496), .A2(n7351), .ZN(n6383) );
  NAND2_X1 U7999 ( .A1(n7344), .A2(n7547), .ZN(n8370) );
  INV_X1 U8000 ( .A(n7344), .ZN(n9495) );
  NAND2_X1 U8001 ( .A1(n9495), .A2(n7309), .ZN(n8308) );
  NAND2_X1 U8002 ( .A1(n7344), .A2(n7309), .ZN(n6385) );
  NAND2_X1 U8003 ( .A1(n10137), .A2(n9493), .ZN(n8515) );
  NAND2_X1 U8004 ( .A1(n7543), .A2(n7379), .ZN(n8363) );
  NAND2_X1 U8005 ( .A1(n8515), .A2(n8363), .ZN(n8361) );
  NOR2_X1 U8006 ( .A1(n7379), .A2(n9493), .ZN(n6386) );
  OR2_X1 U8007 ( .A1(n7535), .A2(n7612), .ZN(n8372) );
  NAND2_X1 U8008 ( .A1(n7535), .A2(n7612), .ZN(n8375) );
  NAND2_X1 U8009 ( .A1(n8372), .A2(n8375), .ZN(n7478) );
  NAND2_X1 U8010 ( .A1(n7535), .A2(n10022), .ZN(n6387) );
  OR2_X1 U8011 ( .A1(n10150), .A2(n7711), .ZN(n8377) );
  NAND2_X1 U8012 ( .A1(n10150), .A2(n7711), .ZN(n8376) );
  INV_X1 U8013 ( .A(n10025), .ZN(n6388) );
  INV_X1 U8014 ( .A(n7711), .ZN(n9492) );
  NAND2_X1 U8015 ( .A1(n7699), .A2(n7787), .ZN(n8386) );
  NAND2_X1 U8016 ( .A1(n8385), .A2(n8386), .ZN(n8261) );
  INV_X1 U8017 ( .A(n7787), .ZN(n10023) );
  OR2_X1 U8018 ( .A1(n7796), .A2(n9491), .ZN(n6389) );
  NAND2_X1 U8019 ( .A1(n7796), .A2(n9491), .ZN(n6390) );
  OR2_X1 U8020 ( .A1(n8028), .A2(n7912), .ZN(n8392) );
  NAND2_X1 U8021 ( .A1(n8028), .A2(n7912), .ZN(n8389) );
  NAND2_X1 U8022 ( .A1(n8392), .A2(n8389), .ZN(n8265) );
  INV_X1 U8023 ( .A(n7912), .ZN(n9490) );
  OR2_X1 U8024 ( .A1(n7915), .A2(n7887), .ZN(n8316) );
  NAND2_X1 U8025 ( .A1(n7915), .A2(n7887), .ZN(n8301) );
  NAND2_X1 U8026 ( .A1(n8316), .A2(n8301), .ZN(n7804) );
  NAND2_X1 U8027 ( .A1(n7803), .A2(n7804), .ZN(n6392) );
  INV_X1 U8028 ( .A(n7887), .ZN(n9489) );
  NAND2_X1 U8029 ( .A1(n7915), .A2(n9489), .ZN(n6391) );
  OR2_X1 U8030 ( .A1(n9808), .A2(n9488), .ZN(n6393) );
  OR2_X1 U8031 ( .A1(n8046), .A2(n8133), .ZN(n8315) );
  NAND2_X1 U8032 ( .A1(n8046), .A2(n8133), .ZN(n8322) );
  INV_X1 U8033 ( .A(n8133), .ZN(n9487) );
  NAND2_X1 U8034 ( .A1(n8060), .A2(n9427), .ZN(n8412) );
  NAND2_X1 U8035 ( .A1(n8411), .A2(n8412), .ZN(n8271) );
  INV_X1 U8036 ( .A(n9427), .ZN(n9731) );
  NAND2_X1 U8037 ( .A1(n8060), .A2(n9731), .ZN(n6394) );
  OR2_X1 U8038 ( .A1(n9803), .A2(n9717), .ZN(n8424) );
  NAND2_X1 U8039 ( .A1(n9803), .A2(n9717), .ZN(n8331) );
  NAND2_X1 U8040 ( .A1(n8424), .A2(n8331), .ZN(n8249) );
  INV_X1 U8041 ( .A(n9717), .ZN(n9732) );
  NAND2_X1 U8042 ( .A1(n9798), .A2(n9708), .ZN(n8425) );
  NAND2_X1 U8043 ( .A1(n9798), .A2(n9485), .ZN(n6395) );
  AND2_X1 U8044 ( .A1(n9793), .A2(n9484), .ZN(n6396) );
  NAND2_X1 U8045 ( .A1(n9788), .A2(n9678), .ZN(n6397) );
  AND2_X1 U8046 ( .A1(n9781), .A2(n9663), .ZN(n8247) );
  OR2_X1 U8047 ( .A1(n9781), .A2(n9663), .ZN(n8246) );
  OAI21_X1 U8048 ( .B1(n9668), .B2(n8247), .A(n8246), .ZN(n9653) );
  OR2_X1 U8049 ( .A1(n9776), .A2(n9456), .ZN(n8334) );
  NAND2_X1 U8050 ( .A1(n9776), .A2(n9456), .ZN(n8447) );
  NAND2_X1 U8051 ( .A1(n8334), .A2(n8447), .ZN(n9661) );
  NAND2_X1 U8052 ( .A1(n9653), .A2(n9661), .ZN(n6399) );
  OR2_X1 U8053 ( .A1(n9776), .A2(n9677), .ZN(n6398) );
  NOR2_X1 U8054 ( .A1(n9772), .A2(n9662), .ZN(n6401) );
  NAND2_X1 U8055 ( .A1(n9772), .A2(n9662), .ZN(n6400) );
  NAND2_X1 U8056 ( .A1(n9768), .A2(n9438), .ZN(n8459) );
  INV_X1 U8057 ( .A(n9632), .ZN(n6402) );
  INV_X1 U8058 ( .A(n9438), .ZN(n9641) );
  OR2_X1 U8059 ( .A1(n9768), .A2(n9641), .ZN(n6403) );
  NAND2_X1 U8060 ( .A1(n6404), .A2(n6403), .ZN(n9610) );
  OR2_X1 U8061 ( .A1(n9761), .A2(n9634), .ZN(n8460) );
  NAND2_X1 U8062 ( .A1(n9761), .A2(n9634), .ZN(n8293) );
  NAND2_X1 U8063 ( .A1(n8460), .A2(n8293), .ZN(n9609) );
  NAND2_X1 U8064 ( .A1(n9610), .A2(n9609), .ZN(n9608) );
  INV_X1 U8065 ( .A(n9634), .ZN(n9483) );
  OR2_X1 U8066 ( .A1(n9761), .A2(n9483), .ZN(n6405) );
  NAND2_X1 U8067 ( .A1(n8576), .A2(n8283), .ZN(n6407) );
  OR2_X1 U8068 ( .A1(n5878), .A2(n8577), .ZN(n6406) );
  NAND2_X1 U8069 ( .A1(n9756), .A2(n9575), .ZN(n8456) );
  INV_X1 U8070 ( .A(n9575), .ZN(n9606) );
  OR2_X1 U8071 ( .A1(n9756), .A2(n9606), .ZN(n6408) );
  NAND2_X1 U8072 ( .A1(n6409), .A2(n8283), .ZN(n6412) );
  INV_X1 U8073 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n6410) );
  OR2_X1 U8074 ( .A1(n5878), .A2(n6410), .ZN(n6411) );
  NAND2_X1 U8075 ( .A1(n5808), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6420) );
  INV_X1 U8076 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6569) );
  OR2_X1 U8077 ( .A1(n6460), .A2(n6569), .ZN(n6419) );
  INV_X1 U8078 ( .A(n6414), .ZN(n6413) );
  NAND2_X1 U8079 ( .A1(n6413), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8581) );
  INV_X1 U8080 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8206) );
  NAND2_X1 U8081 ( .A1(n6414), .A2(n8206), .ZN(n6415) );
  NAND2_X1 U8082 ( .A1(n8581), .A2(n6415), .ZN(n9581) );
  OR2_X1 U8083 ( .A1(n6416), .A2(n9581), .ZN(n6418) );
  INV_X1 U8084 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9582) );
  OR2_X1 U8085 ( .A1(n4448), .A2(n9582), .ZN(n6417) );
  NAND2_X1 U8086 ( .A1(n9584), .A2(n9589), .ZN(n8471) );
  INV_X1 U8087 ( .A(n9589), .ZN(n9482) );
  INV_X1 U8088 ( .A(n6424), .ZN(n6425) );
  NAND2_X1 U8089 ( .A1(n6425), .A2(n6568), .ZN(n6426) );
  INV_X1 U8090 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9380) );
  INV_X1 U8091 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9832) );
  MUX2_X1 U8092 ( .A(n9380), .B(n9832), .S(n4445), .Z(n8215) );
  XNOR2_X1 U8093 ( .A(n8215), .B(SI_29_), .ZN(n6428) );
  NAND2_X1 U8094 ( .A1(n9378), .A2(n8283), .ZN(n6430) );
  OR2_X1 U8095 ( .A1(n5878), .A2(n9832), .ZN(n6429) );
  NAND2_X1 U8096 ( .A1(n5808), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6436) );
  INV_X1 U8097 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6431) );
  OR2_X1 U8098 ( .A1(n6460), .A2(n6431), .ZN(n6435) );
  OR2_X1 U8099 ( .A1(n6416), .A2(n8581), .ZN(n6434) );
  INV_X1 U8100 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n6432) );
  OR2_X1 U8101 ( .A1(n4448), .A2(n6432), .ZN(n6433) );
  NAND2_X1 U8102 ( .A1(n8483), .A2(n9574), .ZN(n8534) );
  INV_X1 U8103 ( .A(n10133), .ZN(n10106) );
  NAND2_X1 U8104 ( .A1(n6438), .A2(n10044), .ZN(n6440) );
  OR2_X1 U8105 ( .A1(n8289), .A2(n8549), .ZN(n6439) );
  INV_X1 U8106 ( .A(n10050), .ZN(n6466) );
  NOR2_X1 U8107 ( .A1(n6441), .A2(n7295), .ZN(n10048) );
  NAND2_X1 U8108 ( .A1(n7289), .A2(n5816), .ZN(n6442) );
  NAND2_X1 U8109 ( .A1(n10047), .A2(n6442), .ZN(n7288) );
  INV_X1 U8110 ( .A(n6443), .ZN(n8252) );
  NAND2_X1 U8111 ( .A1(n7288), .A2(n8252), .ZN(n6444) );
  NAND2_X1 U8112 ( .A1(n8504), .A2(n4969), .ZN(n8503) );
  INV_X1 U8113 ( .A(n7255), .ZN(n8253) );
  NAND2_X1 U8114 ( .A1(n7254), .A2(n8253), .ZN(n6445) );
  NAND2_X1 U8115 ( .A1(n8370), .A2(n8353), .ZN(n8512) );
  NAND2_X1 U8116 ( .A1(n8308), .A2(n8354), .ZN(n6446) );
  NAND2_X1 U8117 ( .A1(n8370), .A2(n6446), .ZN(n8514) );
  NAND2_X1 U8118 ( .A1(n7372), .A2(n8363), .ZN(n7474) );
  NAND2_X1 U8119 ( .A1(n7474), .A2(n8372), .ZN(n6447) );
  NAND2_X1 U8120 ( .A1(n6447), .A2(n8375), .ZN(n10021) );
  INV_X1 U8121 ( .A(n8386), .ZN(n6448) );
  INV_X1 U8122 ( .A(n9491), .ZN(n7886) );
  NAND2_X1 U8123 ( .A1(n7796), .A2(n7886), .ZN(n6449) );
  AND2_X1 U8124 ( .A1(n8389), .A2(n6449), .ZN(n8394) );
  NAND2_X1 U8125 ( .A1(n7785), .A2(n8394), .ZN(n7807) );
  NOR2_X1 U8126 ( .A1(n7796), .A2(n7886), .ZN(n7882) );
  NAND2_X1 U8127 ( .A1(n8389), .A2(n7882), .ZN(n6450) );
  NAND2_X1 U8128 ( .A1(n6450), .A2(n8392), .ZN(n7806) );
  NOR2_X1 U8129 ( .A1(n7804), .A2(n7806), .ZN(n6451) );
  INV_X1 U8130 ( .A(n9488), .ZN(n8300) );
  XNOR2_X1 U8131 ( .A(n9808), .B(n8300), .ZN(n8266) );
  OR2_X1 U8132 ( .A1(n9808), .A2(n8300), .ZN(n8403) );
  AND2_X1 U8133 ( .A1(n8412), .A2(n8322), .ZN(n8409) );
  NAND2_X1 U8134 ( .A1(n6452), .A2(n8411), .ZN(n9730) );
  INV_X1 U8135 ( .A(n9486), .ZN(n8115) );
  NAND2_X1 U8136 ( .A1(n9740), .A2(n8115), .ZN(n8250) );
  AND2_X1 U8137 ( .A1(n8331), .A2(n8250), .ZN(n8419) );
  OR2_X1 U8138 ( .A1(n9740), .A2(n8115), .ZN(n8251) );
  NAND2_X1 U8139 ( .A1(n8424), .A2(n8251), .ZN(n8417) );
  NAND2_X1 U8140 ( .A1(n8417), .A2(n8331), .ZN(n6453) );
  INV_X1 U8141 ( .A(n9484), .ZN(n9715) );
  OR2_X1 U8142 ( .A1(n9793), .A2(n9715), .ZN(n8329) );
  NAND2_X1 U8143 ( .A1(n9793), .A2(n9715), .ZN(n8296) );
  XNOR2_X1 U8144 ( .A(n9788), .B(n9678), .ZN(n9685) );
  NAND2_X1 U8145 ( .A1(n9788), .A2(n9707), .ZN(n8436) );
  NAND2_X1 U8146 ( .A1(n6454), .A2(n8436), .ZN(n9676) );
  AND2_X1 U8147 ( .A1(n9781), .A2(n9688), .ZN(n8433) );
  OR2_X1 U8148 ( .A1(n9781), .A2(n9688), .ZN(n8446) );
  INV_X1 U8149 ( .A(n9661), .ZN(n9652) );
  INV_X1 U8150 ( .A(n8334), .ZN(n8448) );
  AOI21_X1 U8151 ( .B1(n9660), .B2(n9652), .A(n8448), .ZN(n9639) );
  INV_X1 U8152 ( .A(n9662), .ZN(n9635) );
  OR2_X1 U8153 ( .A1(n9772), .A2(n9635), .ZN(n8444) );
  NAND2_X1 U8154 ( .A1(n9772), .A2(n9635), .ZN(n9630) );
  NAND2_X1 U8155 ( .A1(n9639), .A2(n9640), .ZN(n9629) );
  AND2_X1 U8156 ( .A1(n8459), .A2(n9630), .ZN(n8349) );
  NAND2_X1 U8157 ( .A1(n9629), .A2(n8349), .ZN(n6455) );
  INV_X1 U8158 ( .A(n8460), .ZN(n8347) );
  INV_X1 U8159 ( .A(n9567), .ZN(n9571) );
  INV_X1 U8160 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U8161 ( .A1(n5788), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U8162 ( .A1(n5808), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6457) );
  OAI211_X1 U8163 ( .C1(n6460), .C2(n6459), .A(n6458), .B(n6457), .ZN(n9480)
         );
  INV_X1 U8164 ( .A(n9480), .ZN(n6465) );
  INV_X1 U8165 ( .A(n9977), .ZN(n6804) );
  NAND2_X1 U8166 ( .A1(n6804), .A2(P1_B_REG_SCAN_IN), .ZN(n6462) );
  AND2_X1 U8167 ( .A1(n10046), .A2(n6462), .ZN(n9557) );
  INV_X1 U8168 ( .A(n9557), .ZN(n6464) );
  INV_X1 U8169 ( .A(n10045), .ZN(n6463) );
  INV_X1 U8170 ( .A(n9793), .ZN(n9699) );
  NAND3_X1 U8171 ( .A1(n10092), .A2(n10098), .A3(n7295), .ZN(n7297) );
  OR2_X1 U8172 ( .A1(n7297), .A2(n10103), .ZN(n7394) );
  NOR2_X2 U8173 ( .A1(n7394), .A2(n7399), .ZN(n7395) );
  NAND2_X1 U8174 ( .A1(n7395), .A2(n7367), .ZN(n7348) );
  INV_X1 U8175 ( .A(n10150), .ZN(n10030) );
  INV_X1 U8176 ( .A(n8028), .ZN(n7890) );
  NAND2_X1 U8177 ( .A1(n7791), .A2(n7890), .ZN(n7811) );
  INV_X1 U8178 ( .A(n8046), .ZN(n9918) );
  INV_X1 U8179 ( .A(n8060), .ZN(n9913) );
  OR2_X1 U8180 ( .A1(n9736), .A2(n9803), .ZN(n9719) );
  OR2_X1 U8181 ( .A1(n9776), .A2(n9669), .ZN(n9654) );
  INV_X1 U8182 ( .A(n6470), .ZN(n6471) );
  NOR2_X1 U8183 ( .A1(n6472), .A2(n6471), .ZN(n6473) );
  AND2_X1 U8184 ( .A1(n6475), .A2(n6474), .ZN(n6930) );
  NOR2_X1 U8185 ( .A1(n6929), .A2(n6925), .ZN(n6476) );
  INV_X1 U8186 ( .A(keyinput27), .ZN(n6479) );
  NOR4_X1 U8187 ( .A1(keyinput60), .A2(keyinput77), .A3(keyinput115), .A4(
        n6479), .ZN(n6480) );
  NAND3_X1 U8188 ( .A1(keyinput12), .A2(keyinput33), .A3(n6480), .ZN(n6494) );
  INV_X1 U8189 ( .A(keyinput38), .ZN(n6481) );
  NOR4_X1 U8190 ( .A1(keyinput55), .A2(keyinput111), .A3(keyinput109), .A4(
        n6481), .ZN(n6492) );
  NAND2_X1 U8191 ( .A1(keyinput8), .A2(keyinput34), .ZN(n6482) );
  NOR3_X1 U8192 ( .A1(keyinput70), .A2(keyinput98), .A3(n6482), .ZN(n6491) );
  NOR2_X1 U8193 ( .A1(keyinput74), .A2(keyinput125), .ZN(n6483) );
  NAND3_X1 U8194 ( .A1(keyinput89), .A2(keyinput18), .A3(n6483), .ZN(n6489) );
  NAND4_X1 U8195 ( .A1(keyinput123), .A2(keyinput112), .A3(keyinput124), .A4(
        keyinput107), .ZN(n6488) );
  INV_X1 U8196 ( .A(keyinput41), .ZN(n6484) );
  NAND4_X1 U8197 ( .A1(keyinput0), .A2(keyinput62), .A3(keyinput114), .A4(
        n6484), .ZN(n6487) );
  NOR2_X1 U8198 ( .A1(keyinput73), .A2(keyinput113), .ZN(n6485) );
  NAND3_X1 U8199 ( .A1(keyinput80), .A2(keyinput103), .A3(n6485), .ZN(n6486)
         );
  NOR4_X1 U8200 ( .A1(n6489), .A2(n6488), .A3(n6487), .A4(n6486), .ZN(n6490)
         );
  NAND3_X1 U8201 ( .A1(n6492), .A2(n6491), .A3(n6490), .ZN(n6493) );
  NOR4_X1 U8202 ( .A1(keyinput90), .A2(keyinput42), .A3(n6494), .A4(n6493), 
        .ZN(n6528) );
  NAND2_X1 U8203 ( .A1(keyinput119), .A2(keyinput83), .ZN(n6495) );
  NOR3_X1 U8204 ( .A1(keyinput49), .A2(keyinput106), .A3(n6495), .ZN(n6496) );
  NAND3_X1 U8205 ( .A1(keyinput117), .A2(keyinput56), .A3(n6496), .ZN(n6504)
         );
  NOR4_X1 U8206 ( .A1(keyinput39), .A2(keyinput46), .A3(keyinput121), .A4(
        keyinput16), .ZN(n6502) );
  NAND2_X1 U8207 ( .A1(keyinput19), .A2(keyinput52), .ZN(n6497) );
  NOR3_X1 U8208 ( .A1(keyinput72), .A2(keyinput104), .A3(n6497), .ZN(n6501) );
  NOR4_X1 U8209 ( .A1(keyinput127), .A2(keyinput29), .A3(keyinput82), .A4(
        keyinput21), .ZN(n6500) );
  NAND3_X1 U8210 ( .A1(keyinput37), .A2(keyinput71), .A3(keyinput102), .ZN(
        n6498) );
  NOR2_X1 U8211 ( .A1(keyinput20), .A2(n6498), .ZN(n6499) );
  NAND4_X1 U8212 ( .A1(n6502), .A2(n6501), .A3(n6500), .A4(n6499), .ZN(n6503)
         );
  NOR4_X1 U8213 ( .A1(keyinput40), .A2(keyinput93), .A3(n6504), .A4(n6503), 
        .ZN(n6527) );
  NOR2_X1 U8214 ( .A1(keyinput5), .A2(keyinput13), .ZN(n6505) );
  NAND3_X1 U8215 ( .A1(keyinput101), .A2(keyinput43), .A3(n6505), .ZN(n6512)
         );
  INV_X1 U8216 ( .A(keyinput108), .ZN(n6506) );
  NAND4_X1 U8217 ( .A1(keyinput116), .A2(keyinput24), .A3(keyinput6), .A4(
        n6506), .ZN(n6511) );
  NOR2_X1 U8218 ( .A1(keyinput78), .A2(keyinput17), .ZN(n6507) );
  NAND3_X1 U8219 ( .A1(keyinput86), .A2(keyinput44), .A3(n6507), .ZN(n6510) );
  NOR2_X1 U8220 ( .A1(keyinput97), .A2(keyinput2), .ZN(n6508) );
  NAND3_X1 U8221 ( .A1(keyinput54), .A2(keyinput85), .A3(n6508), .ZN(n6509) );
  NOR4_X1 U8222 ( .A1(n6512), .A2(n6511), .A3(n6510), .A4(n6509), .ZN(n6526)
         );
  INV_X1 U8223 ( .A(keyinput96), .ZN(n6513) );
  NAND4_X1 U8224 ( .A1(keyinput57), .A2(keyinput11), .A3(keyinput66), .A4(
        n6513), .ZN(n6520) );
  NOR2_X1 U8225 ( .A1(keyinput48), .A2(keyinput32), .ZN(n6514) );
  NAND3_X1 U8226 ( .A1(keyinput51), .A2(keyinput36), .A3(n6514), .ZN(n6519) );
  NOR2_X1 U8227 ( .A1(keyinput100), .A2(keyinput28), .ZN(n6515) );
  NAND3_X1 U8228 ( .A1(keyinput35), .A2(keyinput4), .A3(n6515), .ZN(n6518) );
  NOR2_X1 U8229 ( .A1(keyinput79), .A2(keyinput105), .ZN(n6516) );
  NAND3_X1 U8230 ( .A1(keyinput64), .A2(keyinput10), .A3(n6516), .ZN(n6517) );
  NOR4_X1 U8231 ( .A1(n6520), .A2(n6519), .A3(n6518), .A4(n6517), .ZN(n6524)
         );
  INV_X1 U8232 ( .A(keyinput91), .ZN(n6521) );
  NAND4_X1 U8233 ( .A1(keyinput84), .A2(keyinput81), .A3(keyinput110), .A4(
        n6521), .ZN(n6522) );
  NOR3_X1 U8234 ( .A1(keyinput126), .A2(keyinput94), .A3(n6522), .ZN(n6523) );
  AND4_X1 U8235 ( .A1(n6524), .A2(n6523), .A3(keyinput7), .A4(keyinput118), 
        .ZN(n6525) );
  AND4_X1 U8236 ( .A1(n6528), .A2(n6527), .A3(n6526), .A4(n6525), .ZN(n6756)
         );
  NAND2_X1 U8237 ( .A1(keyinput87), .A2(keyinput120), .ZN(n6529) );
  NOR3_X1 U8238 ( .A1(keyinput9), .A2(keyinput31), .A3(n6529), .ZN(n6530) );
  NAND3_X1 U8239 ( .A1(keyinput67), .A2(keyinput30), .A3(n6530), .ZN(n6544) );
  NOR2_X1 U8240 ( .A1(keyinput59), .A2(keyinput45), .ZN(n6531) );
  NAND3_X1 U8241 ( .A1(keyinput58), .A2(keyinput23), .A3(n6531), .ZN(n6532) );
  NOR3_X1 U8242 ( .A1(keyinput68), .A2(keyinput95), .A3(n6532), .ZN(n6542) );
  NOR2_X1 U8243 ( .A1(keyinput65), .A2(keyinput63), .ZN(n6533) );
  NAND3_X1 U8244 ( .A1(keyinput75), .A2(keyinput69), .A3(n6533), .ZN(n6540) );
  NOR3_X1 U8245 ( .A1(keyinput47), .A2(keyinput99), .A3(keyinput88), .ZN(n6534) );
  NAND2_X1 U8246 ( .A1(keyinput15), .A2(n6534), .ZN(n6539) );
  NOR2_X1 U8247 ( .A1(keyinput76), .A2(keyinput22), .ZN(n6535) );
  NAND3_X1 U8248 ( .A1(keyinput25), .A2(keyinput14), .A3(n6535), .ZN(n6538) );
  INV_X1 U8249 ( .A(keyinput122), .ZN(n6536) );
  NAND4_X1 U8250 ( .A1(keyinput92), .A2(keyinput61), .A3(keyinput53), .A4(
        n6536), .ZN(n6537) );
  NOR4_X1 U8251 ( .A1(n6540), .A2(n6539), .A3(n6538), .A4(n6537), .ZN(n6541)
         );
  NAND4_X1 U8252 ( .A1(keyinput50), .A2(keyinput26), .A3(n6542), .A4(n6541), 
        .ZN(n6543) );
  NOR4_X1 U8253 ( .A1(keyinput3), .A2(keyinput1), .A3(n6544), .A4(n6543), .ZN(
        n6755) );
  INV_X1 U8254 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6546) );
  AOI22_X1 U8255 ( .A1(n6546), .A2(keyinput127), .B1(keyinput29), .B2(n6959), 
        .ZN(n6545) );
  OAI221_X1 U8256 ( .B1(n6546), .B2(keyinput127), .C1(n6959), .C2(keyinput29), 
        .A(n6545), .ZN(n6553) );
  AOI22_X1 U8257 ( .A1(n4797), .A2(keyinput51), .B1(keyinput32), .B2(n6548), 
        .ZN(n6547) );
  OAI221_X1 U8258 ( .B1(n4797), .B2(keyinput51), .C1(n6548), .C2(keyinput32), 
        .A(n6547), .ZN(n6552) );
  AOI22_X1 U8259 ( .A1(n5065), .A2(keyinput75), .B1(keyinput65), .B2(n6550), 
        .ZN(n6549) );
  OAI221_X1 U8260 ( .B1(n5065), .B2(keyinput75), .C1(n6550), .C2(keyinput65), 
        .A(n6549), .ZN(n6551) );
  NOR3_X1 U8261 ( .A1(n6553), .A2(n6552), .A3(n6551), .ZN(n6583) );
  AOI22_X1 U8262 ( .A1(n7812), .A2(keyinput35), .B1(keyinput28), .B2(n9956), 
        .ZN(n6554) );
  OAI221_X1 U8263 ( .B1(n7812), .B2(keyinput35), .C1(n9956), .C2(keyinput28), 
        .A(n6554), .ZN(n6558) );
  INV_X1 U8264 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6903) );
  AOI22_X1 U8265 ( .A1(n6903), .A2(keyinput50), .B1(keyinput26), .B2(n6556), 
        .ZN(n6555) );
  OAI221_X1 U8266 ( .B1(n6903), .B2(keyinput50), .C1(n6556), .C2(keyinput26), 
        .A(n6555), .ZN(n6557) );
  NOR2_X1 U8267 ( .A1(n6558), .A2(n6557), .ZN(n6564) );
  INV_X1 U8268 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10208) );
  AOI22_X1 U8269 ( .A1(n10208), .A2(keyinput11), .B1(n7066), .B2(keyinput57), 
        .ZN(n6559) );
  OAI221_X1 U8270 ( .B1(n10208), .B2(keyinput11), .C1(n7066), .C2(keyinput57), 
        .A(n6559), .ZN(n6562) );
  INV_X1 U8271 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9942) );
  AOI22_X1 U8272 ( .A1(n9942), .A2(keyinput47), .B1(n7042), .B2(keyinput15), 
        .ZN(n6560) );
  OAI221_X1 U8273 ( .B1(n9942), .B2(keyinput47), .C1(n7042), .C2(keyinput15), 
        .A(n6560), .ZN(n6561) );
  NOR2_X1 U8274 ( .A1(n6562), .A2(n6561), .ZN(n6563) );
  AND2_X1 U8275 ( .A1(n6564), .A2(n6563), .ZN(n6582) );
  INV_X1 U8276 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n6566) );
  INV_X1 U8277 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U8278 ( .A1(n6566), .A2(keyinput23), .B1(keyinput45), .B2(n10203), 
        .ZN(n6565) );
  OAI221_X1 U8279 ( .B1(n6566), .B2(keyinput23), .C1(n10203), .C2(keyinput45), 
        .A(n6565), .ZN(n6574) );
  AOI22_X1 U8280 ( .A1(n6569), .A2(keyinput100), .B1(n6568), .B2(keyinput4), 
        .ZN(n6567) );
  OAI221_X1 U8281 ( .B1(n6569), .B2(keyinput100), .C1(n6568), .C2(keyinput4), 
        .A(n6567), .ZN(n6573) );
  AOI22_X1 U8282 ( .A1(n10059), .A2(keyinput55), .B1(n6571), .B2(keyinput38), 
        .ZN(n6570) );
  OAI221_X1 U8283 ( .B1(n10059), .B2(keyinput55), .C1(n6571), .C2(keyinput38), 
        .A(n6570), .ZN(n6572) );
  NOR3_X1 U8284 ( .A1(n6574), .A2(n6573), .A3(n6572), .ZN(n6581) );
  AOI22_X1 U8285 ( .A1(n9083), .A2(keyinput25), .B1(keyinput76), .B2(n7429), 
        .ZN(n6575) );
  OAI221_X1 U8286 ( .B1(n9083), .B2(keyinput25), .C1(n7429), .C2(keyinput76), 
        .A(n6575), .ZN(n6579) );
  INV_X1 U8287 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7506) );
  AOI22_X1 U8288 ( .A1(n6577), .A2(keyinput82), .B1(keyinput21), .B2(n7506), 
        .ZN(n6576) );
  OAI221_X1 U8289 ( .B1(n6577), .B2(keyinput82), .C1(n7506), .C2(keyinput21), 
        .A(n6576), .ZN(n6578) );
  NOR2_X1 U8290 ( .A1(n6579), .A2(n6578), .ZN(n6580) );
  NAND4_X1 U8291 ( .A1(n6583), .A2(n6582), .A3(n6581), .A4(n6580), .ZN(n6639)
         );
  AOI22_X1 U8292 ( .A1(n6293), .A2(keyinput70), .B1(keyinput34), .B2(n5925), 
        .ZN(n6584) );
  OAI221_X1 U8293 ( .B1(n6293), .B2(keyinput70), .C1(n5925), .C2(keyinput34), 
        .A(n6584), .ZN(n6591) );
  AOI22_X1 U8294 ( .A1(n6586), .A2(keyinput48), .B1(n7384), .B2(keyinput36), 
        .ZN(n6585) );
  OAI221_X1 U8295 ( .B1(n6586), .B2(keyinput48), .C1(n7384), .C2(keyinput36), 
        .A(n6585), .ZN(n6590) );
  XNOR2_X1 U8296 ( .A(P2_IR_REG_27__SCAN_IN), .B(keyinput92), .ZN(n6588) );
  XNOR2_X1 U8297 ( .A(keyinput109), .B(P2_REG0_REG_10__SCAN_IN), .ZN(n6587) );
  NAND2_X1 U8298 ( .A1(n6588), .A2(n6587), .ZN(n6589) );
  NOR3_X1 U8299 ( .A1(n6591), .A2(n6590), .A3(n6589), .ZN(n6614) );
  INV_X1 U8300 ( .A(keyinput105), .ZN(n6593) );
  AOI22_X1 U8301 ( .A1(n6594), .A2(keyinput64), .B1(SI_29_), .B2(n6593), .ZN(
        n6592) );
  OAI221_X1 U8302 ( .B1(n6594), .B2(keyinput64), .C1(n6593), .C2(SI_29_), .A(
        n6592), .ZN(n6598) );
  INV_X1 U8303 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10201) );
  INV_X1 U8304 ( .A(keyinput14), .ZN(n6596) );
  AOI22_X1 U8305 ( .A1(n10201), .A2(keyinput22), .B1(SI_31_), .B2(n6596), .ZN(
        n6595) );
  OAI221_X1 U8306 ( .B1(n10201), .B2(keyinput22), .C1(n6596), .C2(SI_31_), .A(
        n6595), .ZN(n6597) );
  NOR2_X1 U8307 ( .A1(n6598), .A2(n6597), .ZN(n6613) );
  INV_X1 U8308 ( .A(keyinput68), .ZN(n6600) );
  AOI22_X1 U8309 ( .A1(n6848), .A2(keyinput95), .B1(P1_ADDR_REG_4__SCAN_IN), 
        .B2(n6600), .ZN(n6599) );
  OAI221_X1 U8310 ( .B1(n6848), .B2(keyinput95), .C1(n6600), .C2(
        P1_ADDR_REG_4__SCAN_IN), .A(n6599), .ZN(n6604) );
  INV_X1 U8311 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10072) );
  INV_X1 U8312 ( .A(keyinput99), .ZN(n6602) );
  AOI22_X1 U8313 ( .A1(n10072), .A2(keyinput88), .B1(P1_REG2_REG_31__SCAN_IN), 
        .B2(n6602), .ZN(n6601) );
  OAI221_X1 U8314 ( .B1(n10072), .B2(keyinput88), .C1(n6602), .C2(
        P1_REG2_REG_31__SCAN_IN), .A(n6601), .ZN(n6603) );
  NOR2_X1 U8315 ( .A1(n6604), .A2(n6603), .ZN(n6612) );
  AOI22_X1 U8316 ( .A1(n6606), .A2(keyinput122), .B1(keyinput53), .B2(n9626), 
        .ZN(n6605) );
  OAI221_X1 U8317 ( .B1(n6606), .B2(keyinput122), .C1(n9626), .C2(keyinput53), 
        .A(n6605), .ZN(n6610) );
  INV_X1 U8318 ( .A(keyinput8), .ZN(n6608) );
  AOI22_X1 U8319 ( .A1(n8578), .A2(keyinput98), .B1(P2_ADDR_REG_14__SCAN_IN), 
        .B2(n6608), .ZN(n6607) );
  OAI221_X1 U8320 ( .B1(n8578), .B2(keyinput98), .C1(n6608), .C2(
        P2_ADDR_REG_14__SCAN_IN), .A(n6607), .ZN(n6609) );
  NOR2_X1 U8321 ( .A1(n6610), .A2(n6609), .ZN(n6611) );
  NAND4_X1 U8322 ( .A1(n6614), .A2(n6613), .A3(n6612), .A4(n6611), .ZN(n6638)
         );
  INV_X1 U8323 ( .A(keyinput59), .ZN(n6615) );
  XNOR2_X1 U8324 ( .A(n6615), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(n6620) );
  XNOR2_X1 U8325 ( .A(SI_27_), .B(keyinput71), .ZN(n6618) );
  XNOR2_X1 U8326 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput66), .ZN(n6617) );
  INV_X1 U8327 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10283) );
  XNOR2_X1 U8328 ( .A(keyinput61), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n6616) );
  NAND3_X1 U8329 ( .A1(n6618), .A2(n6617), .A3(n6616), .ZN(n6619) );
  NOR2_X1 U8330 ( .A1(n6620), .A2(n6619), .ZN(n6636) );
  XNOR2_X1 U8331 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput63), .ZN(n6624) );
  XNOR2_X1 U8332 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput58), .ZN(n6623) );
  XNOR2_X1 U8333 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput10), .ZN(n6622) );
  XNOR2_X1 U8334 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(keyinput20), .ZN(n6621) );
  NAND4_X1 U8335 ( .A1(n6624), .A2(n6623), .A3(n6622), .A4(n6621), .ZN(n6630)
         );
  XNOR2_X1 U8336 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput37), .ZN(n6628) );
  XNOR2_X1 U8337 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput111), .ZN(n6627) );
  XNOR2_X1 U8338 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput102), .ZN(n6626) );
  XNOR2_X1 U8339 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput96), .ZN(n6625) );
  NAND4_X1 U8340 ( .A1(n6628), .A2(n6627), .A3(n6626), .A4(n6625), .ZN(n6629)
         );
  NOR2_X1 U8341 ( .A1(n6630), .A2(n6629), .ZN(n6635) );
  INV_X1 U8342 ( .A(keyinput79), .ZN(n6631) );
  XNOR2_X1 U8343 ( .A(n10075), .B(n6631), .ZN(n6634) );
  INV_X1 U8344 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10207) );
  INV_X1 U8345 ( .A(keyinput69), .ZN(n6632) );
  XNOR2_X1 U8346 ( .A(n10207), .B(n6632), .ZN(n6633) );
  NAND4_X1 U8347 ( .A1(n6636), .A2(n6635), .A3(n6634), .A4(n6633), .ZN(n6637)
         );
  NOR3_X1 U8348 ( .A1(n6639), .A2(n6638), .A3(n6637), .ZN(n6676) );
  INV_X1 U8349 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10204) );
  AOI22_X1 U8350 ( .A1(n10204), .A2(keyinput72), .B1(n10060), .B2(keyinput19), 
        .ZN(n6640) );
  OAI221_X1 U8351 ( .B1(n10204), .B2(keyinput72), .C1(n10060), .C2(keyinput19), 
        .A(n6640), .ZN(n6649) );
  INV_X1 U8352 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7090) );
  INV_X1 U8353 ( .A(keyinput52), .ZN(n6642) );
  AOI22_X1 U8354 ( .A1(n7090), .A2(keyinput104), .B1(P1_ADDR_REG_14__SCAN_IN), 
        .B2(n6642), .ZN(n6641) );
  OAI221_X1 U8355 ( .B1(n7090), .B2(keyinput104), .C1(n6642), .C2(
        P1_ADDR_REG_14__SCAN_IN), .A(n6641), .ZN(n6648) );
  AOI22_X1 U8356 ( .A1(n9946), .A2(keyinput121), .B1(keyinput16), .B2(n8838), 
        .ZN(n6643) );
  OAI221_X1 U8357 ( .B1(n9946), .B2(keyinput121), .C1(n8838), .C2(keyinput16), 
        .A(n6643), .ZN(n6647) );
  AOI22_X1 U8358 ( .A1(n5740), .A2(keyinput39), .B1(keyinput46), .B2(n6645), 
        .ZN(n6644) );
  OAI221_X1 U8359 ( .B1(n5740), .B2(keyinput39), .C1(n6645), .C2(keyinput46), 
        .A(n6644), .ZN(n6646) );
  NOR4_X1 U8360 ( .A1(n6649), .A2(n6648), .A3(n6647), .A4(n6646), .ZN(n6675)
         );
  INV_X1 U8361 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10209) );
  INV_X1 U8362 ( .A(keyinput24), .ZN(n6651) );
  AOI22_X1 U8363 ( .A1(n10209), .A2(keyinput6), .B1(P1_ADDR_REG_13__SCAN_IN), 
        .B2(n6651), .ZN(n6650) );
  OAI221_X1 U8364 ( .B1(n10209), .B2(keyinput6), .C1(n6651), .C2(
        P1_ADDR_REG_13__SCAN_IN), .A(n6650), .ZN(n6660) );
  AOI22_X1 U8365 ( .A1(n7568), .A2(keyinput116), .B1(n6653), .B2(keyinput108), 
        .ZN(n6652) );
  OAI221_X1 U8366 ( .B1(n7568), .B2(keyinput116), .C1(n6653), .C2(keyinput108), 
        .A(n6652), .ZN(n6659) );
  INV_X1 U8367 ( .A(keyinput43), .ZN(n6655) );
  AOI22_X1 U8368 ( .A1(n6175), .A2(keyinput13), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n6655), .ZN(n6654) );
  OAI221_X1 U8369 ( .B1(n6175), .B2(keyinput13), .C1(n6655), .C2(
        P1_DATAO_REG_30__SCAN_IN), .A(n6654), .ZN(n6658) );
  AOI22_X1 U8370 ( .A1(n8156), .A2(keyinput5), .B1(keyinput101), .B2(n7359), 
        .ZN(n6656) );
  OAI221_X1 U8371 ( .B1(n8156), .B2(keyinput5), .C1(n7359), .C2(keyinput101), 
        .A(n6656), .ZN(n6657) );
  NOR4_X1 U8372 ( .A1(n6660), .A2(n6659), .A3(n6658), .A4(n6657), .ZN(n6674)
         );
  AOI22_X1 U8373 ( .A1(n5067), .A2(keyinput40), .B1(n10076), .B2(keyinput93), 
        .ZN(n6661) );
  OAI221_X1 U8374 ( .B1(n5067), .B2(keyinput40), .C1(n10076), .C2(keyinput93), 
        .A(n6661), .ZN(n6672) );
  INV_X1 U8375 ( .A(keyinput56), .ZN(n6663) );
  AOI22_X1 U8376 ( .A1(n6664), .A2(keyinput117), .B1(P1_DATAO_REG_29__SCAN_IN), 
        .B2(n6663), .ZN(n6662) );
  OAI221_X1 U8377 ( .B1(n6664), .B2(keyinput117), .C1(n6663), .C2(
        P1_DATAO_REG_29__SCAN_IN), .A(n6662), .ZN(n6671) );
  INV_X1 U8378 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10202) );
  AOI22_X1 U8379 ( .A1(n10202), .A2(keyinput49), .B1(keyinput119), .B2(n6666), 
        .ZN(n6665) );
  OAI221_X1 U8380 ( .B1(n10202), .B2(keyinput49), .C1(n6666), .C2(keyinput119), 
        .A(n6665), .ZN(n6670) );
  INV_X1 U8381 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7284) );
  AOI22_X1 U8382 ( .A1(n7284), .A2(keyinput83), .B1(n6668), .B2(keyinput106), 
        .ZN(n6667) );
  OAI221_X1 U8383 ( .B1(n7284), .B2(keyinput83), .C1(n6668), .C2(keyinput106), 
        .A(n6667), .ZN(n6669) );
  NOR4_X1 U8384 ( .A1(n6672), .A2(n6671), .A3(n6670), .A4(n6669), .ZN(n6673)
         );
  NAND4_X1 U8385 ( .A1(n6676), .A2(n6675), .A3(n6674), .A4(n6673), .ZN(n6753)
         );
  INV_X1 U8386 ( .A(keyinput42), .ZN(n6678) );
  AOI22_X1 U8387 ( .A1(n8569), .A2(keyinput90), .B1(P1_ADDR_REG_3__SCAN_IN), 
        .B2(n6678), .ZN(n6677) );
  OAI221_X1 U8388 ( .B1(n8569), .B2(keyinput90), .C1(n6678), .C2(
        P1_ADDR_REG_3__SCAN_IN), .A(n6677), .ZN(n6687) );
  INV_X1 U8389 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n10206) );
  INV_X1 U8390 ( .A(SI_2_), .ZN(n6680) );
  AOI22_X1 U8391 ( .A1(n10206), .A2(keyinput60), .B1(n6680), .B2(keyinput77), 
        .ZN(n6679) );
  OAI221_X1 U8392 ( .B1(n10206), .B2(keyinput60), .C1(n6680), .C2(keyinput77), 
        .A(n6679), .ZN(n6686) );
  AOI22_X1 U8393 ( .A1(n7204), .A2(keyinput12), .B1(keyinput33), .B2(n6854), 
        .ZN(n6681) );
  OAI221_X1 U8394 ( .B1(n7204), .B2(keyinput12), .C1(n6854), .C2(keyinput33), 
        .A(n6681), .ZN(n6685) );
  INV_X1 U8395 ( .A(keyinput115), .ZN(n6683) );
  AOI22_X1 U8396 ( .A1(n6994), .A2(keyinput27), .B1(P1_ADDR_REG_16__SCAN_IN), 
        .B2(n6683), .ZN(n6682) );
  OAI221_X1 U8397 ( .B1(n6994), .B2(keyinput27), .C1(n6683), .C2(
        P1_ADDR_REG_16__SCAN_IN), .A(n6682), .ZN(n6684) );
  NOR4_X1 U8398 ( .A1(n6687), .A2(n6686), .A3(n6685), .A4(n6684), .ZN(n6726)
         );
  INV_X1 U8399 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6689) );
  AOI22_X1 U8400 ( .A1(n6689), .A2(keyinput73), .B1(n5006), .B2(keyinput80), 
        .ZN(n6688) );
  OAI221_X1 U8401 ( .B1(n6689), .B2(keyinput73), .C1(n5006), .C2(keyinput80), 
        .A(n6688), .ZN(n6699) );
  INV_X1 U8402 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9420) );
  INV_X1 U8403 ( .A(keyinput103), .ZN(n6691) );
  AOI22_X1 U8404 ( .A1(n9420), .A2(keyinput113), .B1(P1_WR_REG_SCAN_IN), .B2(
        n6691), .ZN(n6690) );
  OAI221_X1 U8405 ( .B1(n9420), .B2(keyinput113), .C1(n6691), .C2(
        P1_WR_REG_SCAN_IN), .A(n6690), .ZN(n6698) );
  INV_X1 U8406 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7555) );
  AOI22_X1 U8407 ( .A1(n7325), .A2(keyinput62), .B1(keyinput0), .B2(n7555), 
        .ZN(n6692) );
  OAI221_X1 U8408 ( .B1(n7325), .B2(keyinput62), .C1(n7555), .C2(keyinput0), 
        .A(n6692), .ZN(n6697) );
  INV_X1 U8409 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n6695) );
  INV_X1 U8410 ( .A(keyinput114), .ZN(n6694) );
  AOI22_X1 U8411 ( .A1(n6695), .A2(keyinput41), .B1(P2_REG0_REG_30__SCAN_IN), 
        .B2(n6694), .ZN(n6693) );
  OAI221_X1 U8412 ( .B1(n6695), .B2(keyinput41), .C1(n6694), .C2(
        P2_REG0_REG_30__SCAN_IN), .A(n6693), .ZN(n6696) );
  NOR4_X1 U8413 ( .A1(n6699), .A2(n6698), .A3(n6697), .A4(n6696), .ZN(n6725)
         );
  INV_X1 U8414 ( .A(keyinput120), .ZN(n6701) );
  AOI22_X1 U8415 ( .A1(n6319), .A2(keyinput9), .B1(P2_ADDR_REG_2__SCAN_IN), 
        .B2(n6701), .ZN(n6700) );
  OAI221_X1 U8416 ( .B1(n6319), .B2(keyinput9), .C1(n6701), .C2(
        P2_ADDR_REG_2__SCAN_IN), .A(n6700), .ZN(n6712) );
  INV_X1 U8417 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n6703) );
  AOI22_X1 U8418 ( .A1(n9044), .A2(keyinput87), .B1(n6703), .B2(keyinput31), 
        .ZN(n6702) );
  OAI221_X1 U8419 ( .B1(n9044), .B2(keyinput87), .C1(n6703), .C2(keyinput31), 
        .A(n6702), .ZN(n6711) );
  INV_X1 U8420 ( .A(SI_6_), .ZN(n6706) );
  INV_X1 U8421 ( .A(keyinput30), .ZN(n6705) );
  AOI22_X1 U8422 ( .A1(n6706), .A2(keyinput67), .B1(P2_ADDR_REG_12__SCAN_IN), 
        .B2(n6705), .ZN(n6704) );
  OAI221_X1 U8423 ( .B1(n6706), .B2(keyinput67), .C1(n6705), .C2(
        P2_ADDR_REG_12__SCAN_IN), .A(n6704), .ZN(n6710) );
  AOI22_X1 U8424 ( .A1(n6708), .A2(keyinput3), .B1(n10018), .B2(keyinput1), 
        .ZN(n6707) );
  OAI221_X1 U8425 ( .B1(n6708), .B2(keyinput3), .C1(n10018), .C2(keyinput1), 
        .A(n6707), .ZN(n6709) );
  NOR4_X1 U8426 ( .A1(n6712), .A2(n6711), .A3(n6710), .A4(n6709), .ZN(n6724)
         );
  INV_X1 U8427 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U8428 ( .A1(n10148), .A2(keyinput123), .B1(keyinput112), .B2(n5346), 
        .ZN(n6713) );
  OAI221_X1 U8429 ( .B1(n10148), .B2(keyinput123), .C1(n5346), .C2(keyinput112), .A(n6713), .ZN(n6722) );
  AOI22_X1 U8430 ( .A1(n7195), .A2(keyinput74), .B1(keyinput89), .B2(n8873), 
        .ZN(n6714) );
  OAI221_X1 U8431 ( .B1(n7195), .B2(keyinput74), .C1(n8873), .C2(keyinput89), 
        .A(n6714), .ZN(n6721) );
  AOI22_X1 U8432 ( .A1(n10080), .A2(keyinput125), .B1(keyinput18), .B2(n6716), 
        .ZN(n6715) );
  OAI221_X1 U8433 ( .B1(n10080), .B2(keyinput125), .C1(n6716), .C2(keyinput18), 
        .A(n6715), .ZN(n6720) );
  INV_X1 U8434 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10084) );
  AOI22_X1 U8435 ( .A1(n6718), .A2(keyinput124), .B1(n10084), .B2(keyinput107), 
        .ZN(n6717) );
  OAI221_X1 U8436 ( .B1(n6718), .B2(keyinput124), .C1(n10084), .C2(keyinput107), .A(n6717), .ZN(n6719) );
  NOR4_X1 U8437 ( .A1(n6722), .A2(n6721), .A3(n6720), .A4(n6719), .ZN(n6723)
         );
  NAND4_X1 U8438 ( .A1(n6726), .A2(n6725), .A3(n6724), .A4(n6723), .ZN(n6752)
         );
  INV_X1 U8439 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10244) );
  AOI22_X1 U8440 ( .A1(n10244), .A2(keyinput97), .B1(n6728), .B2(keyinput85), 
        .ZN(n6727) );
  OAI221_X1 U8441 ( .B1(n10244), .B2(keyinput97), .C1(n6728), .C2(keyinput85), 
        .A(n6727), .ZN(n6737) );
  INV_X1 U8442 ( .A(keyinput2), .ZN(n6730) );
  AOI22_X1 U8443 ( .A1(n7638), .A2(keyinput54), .B1(P2_ADDR_REG_1__SCAN_IN), 
        .B2(n6730), .ZN(n6729) );
  OAI221_X1 U8444 ( .B1(n7638), .B2(keyinput54), .C1(n6730), .C2(
        P2_ADDR_REG_1__SCAN_IN), .A(n6729), .ZN(n6736) );
  AOI22_X1 U8445 ( .A1(n6732), .A2(keyinput78), .B1(n6900), .B2(keyinput44), 
        .ZN(n6731) );
  OAI221_X1 U8446 ( .B1(n6732), .B2(keyinput78), .C1(n6900), .C2(keyinput44), 
        .A(n6731), .ZN(n6735) );
  INV_X1 U8447 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n8034) );
  AOI22_X1 U8448 ( .A1(n5779), .A2(keyinput86), .B1(keyinput17), .B2(n8034), 
        .ZN(n6733) );
  OAI221_X1 U8449 ( .B1(n5779), .B2(keyinput86), .C1(n8034), .C2(keyinput17), 
        .A(n6733), .ZN(n6734) );
  NOR4_X1 U8450 ( .A1(n6737), .A2(n6736), .A3(n6735), .A4(n6734), .ZN(n6750)
         );
  INV_X1 U8451 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n10205) );
  AOI22_X1 U8452 ( .A1(n8926), .A2(keyinput81), .B1(n10205), .B2(keyinput84), 
        .ZN(n6738) );
  OAI221_X1 U8453 ( .B1(n8926), .B2(keyinput81), .C1(n10205), .C2(keyinput84), 
        .A(n6738), .ZN(n6748) );
  INV_X1 U8454 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6859) );
  AOI22_X1 U8455 ( .A1(n6740), .A2(keyinput118), .B1(n6859), .B2(keyinput7), 
        .ZN(n6739) );
  OAI221_X1 U8456 ( .B1(n6740), .B2(keyinput118), .C1(n6859), .C2(keyinput7), 
        .A(n6739), .ZN(n6747) );
  INV_X1 U8457 ( .A(SI_14_), .ZN(n6743) );
  INV_X1 U8458 ( .A(keyinput94), .ZN(n6742) );
  AOI22_X1 U8459 ( .A1(n6743), .A2(keyinput126), .B1(P1_REG0_REG_31__SCAN_IN), 
        .B2(n6742), .ZN(n6741) );
  OAI221_X1 U8460 ( .B1(n6743), .B2(keyinput126), .C1(n6742), .C2(
        P1_REG0_REG_31__SCAN_IN), .A(n6741), .ZN(n6746) );
  AOI22_X1 U8461 ( .A1(n6072), .A2(keyinput110), .B1(n8086), .B2(keyinput91), 
        .ZN(n6744) );
  OAI221_X1 U8462 ( .B1(n6072), .B2(keyinput110), .C1(n8086), .C2(keyinput91), 
        .A(n6744), .ZN(n6745) );
  NOR4_X1 U8463 ( .A1(n6748), .A2(n6747), .A3(n6746), .A4(n6745), .ZN(n6749)
         );
  NAND2_X1 U8464 ( .A1(n6750), .A2(n6749), .ZN(n6751) );
  OR3_X1 U8465 ( .A1(n6753), .A2(n6752), .A3(n6751), .ZN(n6754) );
  AOI21_X1 U8466 ( .B1(n6756), .B2(n6755), .A(n6754), .ZN(n6757) );
  INV_X1 U8467 ( .A(n6757), .ZN(n6758) );
  XNOR2_X1 U8468 ( .A(n6759), .B(n6758), .ZN(P1_U3552) );
  INV_X2 U8469 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U8470 ( .A(n7990), .ZN(n6760) );
  NAND2_X1 U8471 ( .A1(n8492), .A2(n7990), .ZN(n6761) );
  NAND2_X1 U8472 ( .A1(n6807), .A2(n6761), .ZN(n6786) );
  OAI21_X1 U8473 ( .B1(n6786), .B2(n6762), .A(P1_STATE_REG_SCAN_IN), .ZN(
        P1_U3083) );
  INV_X1 U8474 ( .A(n6763), .ZN(n6764) );
  AOI211_X1 U8475 ( .C1(n6766), .C2(n6765), .A(n8868), .B(n6764), .ZN(n6770)
         );
  NOR2_X1 U8476 ( .A1(n9006), .A2(n8856), .ZN(n6769) );
  OAI22_X1 U8477 ( .A1(n8885), .A2(n9242), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8969), .ZN(n6768) );
  OAI22_X1 U8478 ( .A1(n9230), .A2(n8887), .B1(n8875), .B2(n9232), .ZN(n6767)
         );
  OR4_X1 U8479 ( .A1(n6770), .A2(n6769), .A3(n6768), .A4(n6767), .ZN(P2_U3230)
         );
  INV_X1 U8480 ( .A(n6771), .ZN(n6772) );
  AOI211_X1 U8481 ( .C1(n6774), .C2(n6773), .A(n8868), .B(n6772), .ZN(n6779)
         );
  INV_X1 U8482 ( .A(n9325), .ZN(n9184) );
  NOR2_X1 U8483 ( .A1(n9184), .A2(n8856), .ZN(n6778) );
  OAI22_X1 U8484 ( .A1(n8885), .A2(n9181), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6775), .ZN(n6777) );
  INV_X1 U8485 ( .A(n9210), .ZN(n9012) );
  OAI22_X1 U8486 ( .A1(n9016), .A2(n8887), .B1(n8875), .B2(n9012), .ZN(n6776)
         );
  OR4_X1 U8487 ( .A1(n6779), .A2(n6778), .A3(n6777), .A4(n6776), .ZN(P2_U3235)
         );
  AND2_X1 U8488 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7614) );
  INV_X1 U8489 ( .A(n6792), .ZN(n9504) );
  AOI22_X1 U8490 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n6792), .B1(n9504), .B2(
        n7482), .ZN(n9509) );
  NOR2_X1 U8491 ( .A1(n6867), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6780) );
  AOI21_X1 U8492 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6867), .A(n6780), .ZN(
        n6876) );
  XNOR2_X1 U8493 ( .A(n6851), .B(n6781), .ZN(n9989) );
  NAND2_X1 U8494 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9979) );
  XNOR2_X1 U8495 ( .A(n9966), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9963) );
  NOR2_X1 U8496 ( .A1(n9979), .A2(n9963), .ZN(n9962) );
  AOI21_X1 U8497 ( .B1(n9966), .B2(P1_REG2_REG_1__SCAN_IN), .A(n9962), .ZN(
        n9976) );
  NAND2_X1 U8498 ( .A1(n9984), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6782) );
  OAI21_X1 U8499 ( .B1(n9984), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6782), .ZN(
        n9975) );
  NOR2_X1 U8500 ( .A1(n9976), .A2(n9975), .ZN(n9974) );
  AOI21_X1 U8501 ( .B1(n9984), .B2(P1_REG2_REG_2__SCAN_IN), .A(n9974), .ZN(
        n6824) );
  NAND2_X1 U8502 ( .A1(n6796), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6783) );
  OAI21_X1 U8503 ( .B1(n6796), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6783), .ZN(
        n6823) );
  NAND2_X1 U8504 ( .A1(n6800), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6784) );
  OAI21_X1 U8505 ( .B1(n6800), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6784), .ZN(
        n6830) );
  NOR2_X1 U8506 ( .A1(n6831), .A2(n6830), .ZN(n6829) );
  XNOR2_X1 U8507 ( .A(n10011), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n10005) );
  OAI21_X1 U8508 ( .B1(n6867), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6875), .ZN(
        n9508) );
  NAND2_X1 U8509 ( .A1(n9509), .A2(n9508), .ZN(n9507) );
  OR2_X1 U8510 ( .A1(n6792), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6785) );
  MUX2_X1 U8511 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10018), .S(n7071), .Z(n6789)
         );
  INV_X1 U8512 ( .A(n6786), .ZN(n9951) );
  NOR2_X1 U8513 ( .A1(n9977), .A2(P1_U3084), .ZN(n6787) );
  AND2_X1 U8514 ( .A1(n9951), .A2(n6787), .ZN(n9551) );
  NAND2_X1 U8515 ( .A1(n9551), .A2(n6788), .ZN(n10003) );
  INV_X1 U8516 ( .A(n10003), .ZN(n9994) );
  OAI21_X1 U8517 ( .B1(n6790), .B2(n6789), .A(n9994), .ZN(n6791) );
  NOR2_X1 U8518 ( .A1(n6791), .A2(n7070), .ZN(n6811) );
  XNOR2_X1 U8519 ( .A(n7071), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n7061) );
  AOI22_X1 U8520 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n6792), .B1(n9504), .B2(
        n6803), .ZN(n9502) );
  NOR2_X1 U8521 ( .A1(n6867), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6793) );
  AOI21_X1 U8522 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n6867), .A(n6793), .ZN(
        n6880) );
  XNOR2_X1 U8523 ( .A(n10011), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n10002) );
  XNOR2_X1 U8524 ( .A(n6851), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9991) );
  NAND2_X1 U8525 ( .A1(n9966), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6794) );
  OAI21_X1 U8526 ( .B1(n9966), .B2(P1_REG1_REG_1__SCAN_IN), .A(n6794), .ZN(
        n9960) );
  NOR3_X1 U8527 ( .A1(n9946), .A2(n9956), .A3(n9960), .ZN(n9959) );
  AOI21_X1 U8528 ( .B1(n9966), .B2(P1_REG1_REG_1__SCAN_IN), .A(n9959), .ZN(
        n9972) );
  XNOR2_X1 U8529 ( .A(n9984), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9971) );
  NOR2_X1 U8530 ( .A1(n9972), .A2(n9971), .ZN(n9970) );
  AOI21_X1 U8531 ( .B1(n9984), .B2(P1_REG1_REG_2__SCAN_IN), .A(n9970), .ZN(
        n6821) );
  NAND2_X1 U8532 ( .A1(n6796), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6795) );
  OAI21_X1 U8533 ( .B1(n6796), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6795), .ZN(
        n6820) );
  NOR2_X1 U8534 ( .A1(n6821), .A2(n6820), .ZN(n6819) );
  AOI21_X1 U8535 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n6796), .A(n6819), .ZN(
        n9990) );
  AOI22_X1 U8536 ( .A1(n9991), .A2(n9990), .B1(n6851), .B2(n6797), .ZN(n6798)
         );
  INV_X1 U8537 ( .A(n6798), .ZN(n6834) );
  NAND2_X1 U8538 ( .A1(n6800), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6799) );
  OAI21_X1 U8539 ( .B1(n6800), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6799), .ZN(
        n6833) );
  NOR2_X1 U8540 ( .A1(n6834), .A2(n6833), .ZN(n6832) );
  AOI21_X1 U8541 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n6800), .A(n6832), .ZN(
        n6801) );
  INV_X1 U8542 ( .A(n6801), .ZN(n10001) );
  OAI22_X1 U8543 ( .A1(n10002), .A2(n10001), .B1(n10011), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n6879) );
  NAND2_X1 U8544 ( .A1(n6880), .A2(n6879), .ZN(n6878) );
  OAI21_X1 U8545 ( .B1(n6867), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6878), .ZN(
        n9501) );
  NAND2_X1 U8546 ( .A1(n9502), .A2(n9501), .ZN(n9500) );
  INV_X1 U8547 ( .A(n9500), .ZN(n6802) );
  AOI21_X1 U8548 ( .B1(n6803), .B2(n9504), .A(n6802), .ZN(n7062) );
  XOR2_X1 U8549 ( .A(n7061), .B(n7062), .Z(n6806) );
  OR2_X1 U8550 ( .A1(n6302), .A2(P1_U3084), .ZN(n9949) );
  NOR2_X1 U8551 ( .A1(n9949), .A2(n6804), .ZN(n6805) );
  NAND2_X1 U8552 ( .A1(n9951), .A2(n6805), .ZN(n9969) );
  NOR2_X1 U8553 ( .A1(n6806), .A2(n9969), .ZN(n6810) );
  AND2_X1 U8554 ( .A1(n9551), .A2(n6302), .ZN(n10012) );
  INV_X1 U8555 ( .A(n7071), .ZN(n6901) );
  INV_X1 U8556 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10333) );
  INV_X1 U8557 ( .A(n6807), .ZN(n6808) );
  OAI22_X1 U8558 ( .A1(n9525), .A2(n6901), .B1(n10333), .B2(n9999), .ZN(n6809)
         );
  OR4_X1 U8559 ( .A1(n7614), .A2(n6811), .A3(n6810), .A4(n6809), .ZN(P1_U3250)
         );
  INV_X1 U8560 ( .A(n8881), .ZN(n6812) );
  AOI211_X1 U8561 ( .C1(n6814), .C2(n6813), .A(n8868), .B(n6812), .ZN(n6818)
         );
  NOR2_X1 U8562 ( .A1(n8875), .A2(n8827), .ZN(n6817) );
  OAI22_X1 U8563 ( .A1(n8887), .A2(n8641), .B1(n8885), .B2(n10186), .ZN(n6816)
         );
  INV_X1 U8564 ( .A(n10187), .ZN(n7520) );
  OAI22_X1 U8565 ( .A1(n8856), .A2(n7520), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5154), .ZN(n6815) );
  OR4_X1 U8566 ( .A1(n6818), .A2(n6817), .A3(n6816), .A4(n6815), .ZN(P2_U3229)
         );
  INV_X1 U8567 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7261) );
  NOR2_X1 U8568 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7261), .ZN(n7122) );
  AOI211_X1 U8569 ( .C1(n6821), .C2(n6820), .A(n6819), .B(n9969), .ZN(n6828)
         );
  AOI211_X1 U8570 ( .C1(n6824), .C2(n6823), .A(n6822), .B(n10003), .ZN(n6827)
         );
  INV_X1 U8571 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6825) );
  OAI22_X1 U8572 ( .A1(n9525), .A2(n6847), .B1(n6825), .B2(n9999), .ZN(n6826)
         );
  OR4_X1 U8573 ( .A1(n7122), .A2(n6828), .A3(n6827), .A4(n6826), .ZN(P1_U3244)
         );
  AND2_X1 U8574 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7366) );
  AOI211_X1 U8575 ( .C1(n6831), .C2(n6830), .A(n6829), .B(n10003), .ZN(n6837)
         );
  AOI211_X1 U8576 ( .C1(n6834), .C2(n6833), .A(n6832), .B(n9969), .ZN(n6836)
         );
  INV_X1 U8577 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10325) );
  OAI22_X1 U8578 ( .A1(n9525), .A2(n6860), .B1(n10325), .B2(n9999), .ZN(n6835)
         );
  OR4_X1 U8579 ( .A1(n7366), .A2(n6837), .A3(n6836), .A4(n6835), .ZN(P1_U3246)
         );
  NAND2_X1 U8580 ( .A1(n8228), .A2(P1_U3084), .ZN(n7992) );
  INV_X1 U8581 ( .A(n7992), .ZN(n9836) );
  INV_X1 U8582 ( .A(n9836), .ZN(n9831) );
  AND2_X1 U8583 ( .A1(n4445), .A2(P1_U3084), .ZN(n7988) );
  OAI222_X1 U8584 ( .A1(n9831), .A2(n6840), .B1(n9835), .B2(n6844), .C1(
        P1_U3084), .C2(n6839), .ZN(P1_U3352) );
  OAI222_X1 U8585 ( .A1(n9831), .A2(n6842), .B1(n9835), .B2(n6846), .C1(
        P1_U3084), .C2(n6841), .ZN(P1_U3351) );
  NOR2_X1 U8586 ( .A1(n8228), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9376) );
  INV_X1 U8587 ( .A(n9376), .ZN(n9379) );
  AND2_X1 U8588 ( .A1(n8228), .A2(P2_U3152), .ZN(n7985) );
  OAI222_X1 U8589 ( .A1(n9379), .A2(n6845), .B1(n4451), .B2(n6844), .C1(
        P2_U3152), .C2(n6843), .ZN(P2_U3357) );
  OAI222_X1 U8590 ( .A1(n9379), .A2(n4757), .B1(n4451), .B2(n6846), .C1(
        P2_U3152), .C2(n6982), .ZN(P2_U3356) );
  OAI222_X1 U8591 ( .A1(n7992), .A2(n6848), .B1(n9835), .B2(n6849), .C1(
        P1_U3084), .C2(n6847), .ZN(P1_U3350) );
  OAI222_X1 U8592 ( .A1(n9379), .A2(n6850), .B1(n4451), .B2(n6849), .C1(
        P2_U3152), .C2(n7118), .ZN(P2_U3355) );
  OAI222_X1 U8593 ( .A1(n9831), .A2(n6852), .B1(n9835), .B2(n6853), .C1(
        P1_U3084), .C2(n6851), .ZN(P1_U3349) );
  OAI222_X1 U8594 ( .A1(n9379), .A2(n6854), .B1(n4451), .B2(n6853), .C1(
        P2_U3152), .C2(n7103), .ZN(P2_U3354) );
  INV_X1 U8595 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6856) );
  NAND2_X1 U8596 ( .A1(n7242), .A2(n6928), .ZN(n6855) );
  OAI21_X1 U8597 ( .B1(n6928), .B2(n6856), .A(n6855), .ZN(P1_U3441) );
  NAND2_X1 U8598 ( .A1(n6857), .A2(n6928), .ZN(n6858) );
  OAI21_X1 U8599 ( .B1(n6928), .B2(n6859), .A(n6858), .ZN(P1_U3440) );
  OAI222_X1 U8600 ( .A1(n9831), .A2(n6861), .B1(n9835), .B2(n6862), .C1(
        P1_U3084), .C2(n6860), .ZN(P1_U3348) );
  OAI222_X1 U8601 ( .A1(n9379), .A2(n6863), .B1(n4451), .B2(n6862), .C1(
        P2_U3152), .C2(n6987), .ZN(P2_U3353) );
  AOI22_X1 U8602 ( .A1(n10011), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9836), .ZN(n6864) );
  OAI21_X1 U8603 ( .B1(n6865), .B2(n9835), .A(n6864), .ZN(P1_U3347) );
  OAI222_X1 U8604 ( .A1(n9379), .A2(n6866), .B1(n4451), .B2(n6865), .C1(
        P2_U3152), .C2(n7089), .ZN(P2_U3352) );
  INV_X1 U8605 ( .A(n6867), .ZN(n6883) );
  OAI222_X1 U8606 ( .A1(n7992), .A2(n6868), .B1(n9835), .B2(n6869), .C1(
        P1_U3084), .C2(n6883), .ZN(P1_U3346) );
  OAI222_X1 U8607 ( .A1(n9379), .A2(n6870), .B1(n4451), .B2(n6869), .C1(
        P2_U3152), .C2(n7141), .ZN(P2_U3351) );
  INV_X1 U8608 ( .A(n6871), .ZN(n6873) );
  OAI222_X1 U8609 ( .A1(n9831), .A2(n6872), .B1(n9835), .B2(n6873), .C1(
        P1_U3084), .C2(n9504), .ZN(P1_U3345) );
  OAI222_X1 U8610 ( .A1(n9379), .A2(n6874), .B1(n4451), .B2(n6873), .C1(
        P2_U3152), .C2(n8927), .ZN(P2_U3350) );
  INV_X1 U8611 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6887) );
  OAI21_X1 U8612 ( .B1(n6877), .B2(n6876), .A(n6875), .ZN(n6885) );
  OAI21_X1 U8613 ( .B1(n6880), .B2(n6879), .A(n6878), .ZN(n6881) );
  AND2_X1 U8614 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7321) );
  AOI21_X1 U8615 ( .B1(n10010), .B2(n6881), .A(n7321), .ZN(n6882) );
  OAI21_X1 U8616 ( .B1(n9525), .B2(n6883), .A(n6882), .ZN(n6884) );
  AOI21_X1 U8617 ( .B1(n9994), .B2(n6885), .A(n6884), .ZN(n6886) );
  OAI21_X1 U8618 ( .B1(n9999), .B2(n6887), .A(n6886), .ZN(P1_U3248) );
  INV_X1 U8619 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6893) );
  INV_X1 U8620 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6891) );
  INV_X1 U8621 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8240) );
  OR2_X1 U8622 ( .A1(n6888), .A2(n8240), .ZN(n6890) );
  NAND2_X1 U8623 ( .A1(n4458), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6889) );
  OAI211_X1 U8624 ( .C1(n5522), .C2(n6891), .A(n6890), .B(n6889), .ZN(n8605)
         );
  NAND2_X1 U8625 ( .A1(n8605), .A2(P2_U3966), .ZN(n6892) );
  OAI21_X1 U8626 ( .B1(n6893), .B2(P2_U3966), .A(n6892), .ZN(P2_U3583) );
  NAND2_X1 U8627 ( .A1(n6894), .A2(n6972), .ZN(n6898) );
  OR2_X1 U8628 ( .A1(n6895), .A2(P2_U3152), .ZN(n8803) );
  NAND2_X1 U8629 ( .A1(n10200), .A2(n8803), .ZN(n6896) );
  NAND2_X1 U8630 ( .A1(n6896), .A2(n4711), .ZN(n6897) );
  AND2_X1 U8631 ( .A1(n6898), .A2(n6897), .ZN(n8999) );
  INV_X1 U8632 ( .A(n8999), .ZN(n10176) );
  NOR2_X1 U8633 ( .A1(n10176), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X2 U8634 ( .A(n7988), .ZN(n9835) );
  INV_X1 U8635 ( .A(n6899), .ZN(n6904) );
  OAI222_X1 U8636 ( .A1(n9835), .A2(n6904), .B1(n6901), .B2(P1_U3084), .C1(
        n6900), .C2(n9831), .ZN(P1_U3344) );
  NAND2_X1 U8637 ( .A1(n6441), .A2(P1_U4006), .ZN(n6902) );
  OAI21_X1 U8638 ( .B1(n9494), .B2(n6903), .A(n6902), .ZN(P1_U3555) );
  INV_X1 U8639 ( .A(n6996), .ZN(n7147) );
  OAI222_X1 U8640 ( .A1(n9379), .A2(n6905), .B1(n4451), .B2(n6904), .C1(n7147), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8641 ( .A(n6906), .ZN(n6915) );
  INV_X1 U8642 ( .A(n7171), .ZN(n7063) );
  OAI222_X1 U8643 ( .A1(n9835), .A2(n6915), .B1(n7063), .B2(P1_U3084), .C1(
        n6907), .C2(n9831), .ZN(P1_U3343) );
  INV_X1 U8644 ( .A(n6908), .ZN(n6918) );
  AOI22_X1 U8645 ( .A1(n7048), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n9376), .ZN(n6909) );
  OAI21_X1 U8646 ( .B1(n6918), .B2(n4451), .A(n6909), .ZN(P2_U3347) );
  INV_X1 U8647 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6914) );
  INV_X1 U8648 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9559) );
  NAND2_X1 U8649 ( .A1(n5884), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6912) );
  INV_X1 U8650 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6910) );
  OR2_X1 U8651 ( .A1(n5868), .A2(n6910), .ZN(n6911) );
  OAI211_X1 U8652 ( .C1(n4448), .C2(n9559), .A(n6912), .B(n6911), .ZN(n9558)
         );
  NAND2_X1 U8653 ( .A1(n9558), .A2(n9494), .ZN(n6913) );
  OAI21_X1 U8654 ( .B1(n9494), .B2(n6914), .A(n6913), .ZN(P1_U3586) );
  INV_X1 U8655 ( .A(n6999), .ZN(n8940) );
  OAI222_X1 U8656 ( .A1(n9379), .A2(n6916), .B1(n4451), .B2(n6915), .C1(n8940), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8657 ( .A(n7335), .ZN(n7169) );
  OAI222_X1 U8658 ( .A1(n9835), .A2(n6918), .B1(n7169), .B2(P1_U3084), .C1(
        n6917), .C2(n9831), .ZN(P1_U3342) );
  INV_X1 U8659 ( .A(n9430), .ZN(n7561) );
  NOR2_X1 U8660 ( .A1(n7561), .A2(n6925), .ZN(n7015) );
  INV_X1 U8661 ( .A(n7015), .ZN(n6919) );
  INV_X1 U8662 ( .A(n9473), .ZN(n8126) );
  AOI22_X1 U8663 ( .A1(n6919), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n8126), .B2(
        n9499), .ZN(n6924) );
  OAI21_X1 U8664 ( .B1(n6922), .B2(n6921), .A(n6920), .ZN(n9978) );
  NAND2_X1 U8665 ( .A1(n9978), .A2(n9467), .ZN(n6923) );
  OAI211_X1 U8666 ( .C1(n9478), .C2(n7295), .A(n6924), .B(n6923), .ZN(P1_U3230) );
  INV_X1 U8667 ( .A(n6925), .ZN(n6927) );
  INV_X1 U8668 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6935) );
  AND2_X1 U8669 ( .A1(n6441), .A2(n7295), .ZN(n8498) );
  NOR2_X1 U8670 ( .A1(n10048), .A2(n8498), .ZN(n8254) );
  NOR3_X1 U8671 ( .A1(n8254), .A2(n6932), .A3(n6931), .ZN(n6933) );
  AOI21_X1 U8672 ( .B1(n10046), .B2(n9499), .A(n6933), .ZN(n7251) );
  OAI21_X1 U8673 ( .B1(n7295), .B2(n7244), .A(n7251), .ZN(n9811) );
  NAND2_X1 U8674 ( .A1(n9811), .A2(n10160), .ZN(n6934) );
  OAI21_X1 U8675 ( .B1(n10160), .B2(n6935), .A(n6934), .ZN(P1_U3454) );
  INV_X1 U8676 ( .A(n6936), .ZN(n6938) );
  NAND2_X1 U8677 ( .A1(n6938), .A2(n6937), .ZN(n6940) );
  AOI22_X1 U8678 ( .A1(n7010), .A2(n6941), .B1(n6940), .B2(n6939), .ZN(n6946)
         );
  INV_X1 U8679 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6943) );
  INV_X1 U8680 ( .A(n9455), .ZN(n9475) );
  AOI22_X1 U8681 ( .A1(n8126), .A2(n5785), .B1(n9475), .B2(n6441), .ZN(n6942)
         );
  OAI21_X1 U8682 ( .B1(n7015), .B2(n6943), .A(n6942), .ZN(n6944) );
  AOI21_X1 U8683 ( .B1(n9459), .B2(n5816), .A(n6944), .ZN(n6945) );
  OAI21_X1 U8684 ( .B1(n6946), .B2(n9461), .A(n6945), .ZN(P1_U3220) );
  INV_X1 U8685 ( .A(n6947), .ZN(n7041) );
  AOI22_X1 U8686 ( .A1(n7183), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n9376), .ZN(n6948) );
  OAI21_X1 U8687 ( .B1(n7041), .B2(n4451), .A(n6948), .ZN(P2_U3346) );
  NOR2_X1 U8688 ( .A1(n7470), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10175) );
  INV_X1 U8689 ( .A(n7469), .ZN(n10217) );
  NOR2_X1 U8690 ( .A1(n8856), .A2(n10217), .ZN(n6953) );
  AOI211_X1 U8691 ( .C1(P2_REG3_REG_0__SCAN_IN), .C2(n7207), .A(n10175), .B(
        n6953), .ZN(n6958) );
  INV_X1 U8692 ( .A(n6954), .ZN(n7159) );
  OAI22_X1 U8693 ( .A1(n8892), .A2(n7159), .B1(n10217), .B2(n8868), .ZN(n6956)
         );
  NAND2_X1 U8694 ( .A1(n6956), .A2(n6955), .ZN(n6957) );
  OAI211_X1 U8695 ( .C1(n7026), .C2(n8887), .A(n6958), .B(n6957), .ZN(P2_U3234) );
  NAND2_X1 U8696 ( .A1(n6996), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6967) );
  NAND2_X1 U8697 ( .A1(n6991), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6964) );
  MUX2_X1 U8698 ( .A(n7529), .B(P2_REG2_REG_7__SCAN_IN), .S(n6991), .Z(n7133)
         );
  INV_X1 U8699 ( .A(n7133), .ZN(n6962) );
  MUX2_X1 U8700 ( .A(n7568), .B(P2_REG2_REG_6__SCAN_IN), .S(n7089), .Z(n7086)
         );
  MUX2_X1 U8701 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n6959), .S(n8918), .Z(n8915)
         );
  NAND2_X1 U8702 ( .A1(n9846), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6961) );
  MUX2_X1 U8703 ( .A(n7625), .B(P2_REG2_REG_1__SCAN_IN), .S(n9846), .Z(n6960)
         );
  INV_X1 U8704 ( .A(n6960), .ZN(n9848) );
  NAND3_X1 U8705 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n9848), .ZN(n9847) );
  NAND2_X1 U8706 ( .A1(n6961), .A2(n9847), .ZN(n9863) );
  MUX2_X1 U8707 ( .A(n7429), .B(P2_REG2_REG_2__SCAN_IN), .S(n6982), .Z(n9862)
         );
  NAND2_X1 U8708 ( .A1(n9863), .A2(n9862), .ZN(n9861) );
  INV_X1 U8709 ( .A(n6982), .ZN(n9859) );
  NAND2_X1 U8710 ( .A1(n9859), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7113) );
  INV_X1 U8711 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7587) );
  MUX2_X1 U8712 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7587), .S(n7118), .Z(n7112)
         );
  AOI21_X1 U8713 ( .B1(n9861), .B2(n7113), .A(n7112), .ZN(n7111) );
  NOR2_X1 U8714 ( .A1(n7118), .A2(n7587), .ZN(n7098) );
  MUX2_X1 U8715 ( .A(n7596), .B(P2_REG2_REG_4__SCAN_IN), .S(n7103), .Z(n7097)
         );
  OAI21_X1 U8716 ( .B1(n7111), .B2(n7098), .A(n7097), .ZN(n7100) );
  OAI21_X1 U8717 ( .B1(n7596), .B2(n7103), .A(n7100), .ZN(n8916) );
  NAND2_X1 U8718 ( .A1(n8915), .A2(n8916), .ZN(n8914) );
  OAI21_X1 U8719 ( .B1(n6987), .B2(n6959), .A(n8914), .ZN(n7085) );
  NAND2_X1 U8720 ( .A1(n7086), .A2(n7085), .ZN(n7084) );
  OAI21_X1 U8721 ( .B1(n7568), .B2(n7089), .A(n7084), .ZN(n7134) );
  NAND2_X1 U8722 ( .A1(n6962), .A2(n7134), .ZN(n6963) );
  NAND2_X1 U8723 ( .A1(n6964), .A2(n6963), .ZN(n8935) );
  MUX2_X1 U8724 ( .A(n7655), .B(P2_REG2_REG_8__SCAN_IN), .S(n8927), .Z(n8934)
         );
  NAND2_X1 U8725 ( .A1(n8935), .A2(n8934), .ZN(n8933) );
  OAI21_X1 U8726 ( .B1(n7655), .B2(n8927), .A(n8933), .ZN(n7145) );
  MUX2_X1 U8727 ( .A(n7686), .B(P2_REG2_REG_9__SCAN_IN), .S(n6996), .Z(n7146)
         );
  INV_X1 U8728 ( .A(n7146), .ZN(n6965) );
  NAND2_X1 U8729 ( .A1(n7145), .A2(n6965), .ZN(n6966) );
  NAND2_X1 U8730 ( .A1(n6967), .A2(n6966), .ZN(n8948) );
  MUX2_X1 U8731 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7766), .S(n6999), .Z(n8947)
         );
  NAND2_X1 U8732 ( .A1(n8948), .A2(n8947), .ZN(n8946) );
  OAI21_X1 U8733 ( .B1(n7766), .B2(n8940), .A(n8946), .ZN(n6969) );
  MUX2_X1 U8734 ( .A(n7864), .B(P2_REG2_REG_11__SCAN_IN), .S(n7048), .Z(n6968)
         );
  NOR2_X1 U8735 ( .A1(n6969), .A2(n6968), .ZN(n7049) );
  AOI21_X1 U8736 ( .B1(n6969), .B2(n6968), .A(n7049), .ZN(n7008) );
  NAND2_X1 U8737 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6970), .ZN(n6971) );
  OAI211_X1 U8738 ( .C1(n10200), .C2(n6972), .A(n6971), .B(n8803), .ZN(n7003)
         );
  NAND2_X1 U8739 ( .A1(n7003), .A2(n7001), .ZN(n6973) );
  NAND2_X1 U8740 ( .A1(n6973), .A2(n8913), .ZN(n6976) );
  NOR2_X1 U8741 ( .A1(n8809), .A2(n6974), .ZN(n6975) );
  NAND2_X1 U8742 ( .A1(n6976), .A2(n6975), .ZN(n8990) );
  INV_X1 U8743 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n6978) );
  OR2_X1 U8744 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7749), .ZN(n6977) );
  OAI21_X1 U8745 ( .B1(n8999), .B2(n6978), .A(n6977), .ZN(n6979) );
  AOI21_X1 U8746 ( .B1(n9860), .B2(n7048), .A(n6979), .ZN(n7007) );
  INV_X1 U8747 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7000) );
  INV_X1 U8748 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6998) );
  INV_X1 U8749 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6993) );
  INV_X1 U8750 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6983) );
  MUX2_X1 U8751 ( .A(n10283), .B(P2_REG1_REG_2__SCAN_IN), .S(n6982), .Z(n9856)
         );
  NAND2_X1 U8752 ( .A1(n9846), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6981) );
  NAND2_X1 U8753 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9844) );
  OAI21_X1 U8754 ( .B1(n9846), .B2(P2_REG1_REG_1__SCAN_IN), .A(n6981), .ZN(
        n9843) );
  NOR2_X1 U8755 ( .A1(n9844), .A2(n9843), .ZN(n9842) );
  INV_X1 U8756 ( .A(n9842), .ZN(n6980) );
  NAND2_X1 U8757 ( .A1(n6981), .A2(n6980), .ZN(n9855) );
  NAND2_X1 U8758 ( .A1(n9856), .A2(n9855), .ZN(n9854) );
  OAI21_X1 U8759 ( .B1(n10283), .B2(n6982), .A(n9854), .ZN(n7106) );
  XNOR2_X1 U8760 ( .A(n7118), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n7107) );
  NAND2_X1 U8761 ( .A1(n7106), .A2(n7107), .ZN(n7105) );
  OAI21_X1 U8762 ( .B1(n6983), .B2(n7118), .A(n7105), .ZN(n7092) );
  XNOR2_X1 U8763 ( .A(n7103), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n7093) );
  NAND2_X1 U8764 ( .A1(n7092), .A2(n7093), .ZN(n7091) );
  OAI21_X1 U8765 ( .B1(n6984), .B2(n7103), .A(n7091), .ZN(n8920) );
  NAND2_X1 U8766 ( .A1(n8918), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6985) );
  OAI21_X1 U8767 ( .B1(n8918), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6985), .ZN(
        n6986) );
  INV_X1 U8768 ( .A(n6986), .ZN(n8921) );
  NAND2_X1 U8769 ( .A1(n8920), .A2(n8921), .ZN(n8919) );
  OAI21_X1 U8770 ( .B1(n6988), .B2(n6987), .A(n8919), .ZN(n7080) );
  XNOR2_X1 U8771 ( .A(n7089), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n7081) );
  NAND2_X1 U8772 ( .A1(n7080), .A2(n7081), .ZN(n7079) );
  OAI21_X1 U8773 ( .B1(n6989), .B2(n7089), .A(n7079), .ZN(n7137) );
  NAND2_X1 U8774 ( .A1(n6991), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6990) );
  OAI21_X1 U8775 ( .B1(n6991), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6990), .ZN(
        n6992) );
  INV_X1 U8776 ( .A(n6992), .ZN(n7138) );
  NAND2_X1 U8777 ( .A1(n7137), .A2(n7138), .ZN(n7136) );
  OAI21_X1 U8778 ( .B1(n6993), .B2(n7141), .A(n7136), .ZN(n8931) );
  MUX2_X1 U8779 ( .A(n6994), .B(P2_REG1_REG_8__SCAN_IN), .S(n8927), .Z(n8932)
         );
  NAND2_X1 U8780 ( .A1(n8931), .A2(n8932), .ZN(n8930) );
  OAI21_X1 U8781 ( .B1(n8927), .B2(n6994), .A(n8930), .ZN(n7151) );
  NAND2_X1 U8782 ( .A1(n6996), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6995) );
  OAI21_X1 U8783 ( .B1(n6996), .B2(P2_REG1_REG_9__SCAN_IN), .A(n6995), .ZN(
        n6997) );
  INV_X1 U8784 ( .A(n6997), .ZN(n7152) );
  NAND2_X1 U8785 ( .A1(n7151), .A2(n7152), .ZN(n7150) );
  OAI21_X1 U8786 ( .B1(n6998), .B2(n7147), .A(n7150), .ZN(n8945) );
  MUX2_X1 U8787 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7000), .S(n6999), .Z(n8944)
         );
  NAND2_X1 U8788 ( .A1(n8945), .A2(n8944), .ZN(n8943) );
  OAI21_X1 U8789 ( .B1(n7000), .B2(n8940), .A(n8943), .ZN(n7005) );
  INV_X1 U8790 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10290) );
  MUX2_X1 U8791 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10290), .S(n7048), .Z(n7004) );
  NAND2_X1 U8792 ( .A1(n7005), .A2(n7004), .ZN(n7043) );
  AND2_X1 U8793 ( .A1(n7001), .A2(n6974), .ZN(n7002) );
  OAI211_X1 U8794 ( .C1(n7005), .C2(n7004), .A(n7043), .B(n10174), .ZN(n7006)
         );
  OAI211_X1 U8795 ( .C1(n7008), .C2(n8990), .A(n7007), .B(n7006), .ZN(P2_U3256) );
  INV_X1 U8796 ( .A(n7011), .ZN(n7012) );
  AOI21_X1 U8797 ( .B1(n7009), .B2(n7013), .A(n7012), .ZN(n7018) );
  AOI22_X1 U8798 ( .A1(n9475), .A2(n9499), .B1(n8126), .B2(n9498), .ZN(n7014)
         );
  OAI21_X1 U8799 ( .B1(n7015), .B2(n7293), .A(n7014), .ZN(n7016) );
  AOI21_X1 U8800 ( .B1(n9459), .B2(n4969), .A(n7016), .ZN(n7017) );
  OAI21_X1 U8801 ( .B1(n7018), .B2(n9461), .A(n7017), .ZN(P1_U3235) );
  INV_X1 U8802 ( .A(n7128), .ZN(n7024) );
  NOR2_X1 U8803 ( .A1(n10200), .A2(n7020), .ZN(n7021) );
  INV_X1 U8804 ( .A(n7126), .ZN(n7023) );
  INV_X1 U8805 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7040) );
  INV_X1 U8806 ( .A(n7028), .ZN(n7031) );
  INV_X1 U8807 ( .A(n7270), .ZN(n7029) );
  AOI21_X1 U8808 ( .B1(n7031), .B2(n7030), .A(n7029), .ZN(n7620) );
  XNOR2_X1 U8809 ( .A(n7422), .B(n8800), .ZN(n9234) );
  NAND2_X1 U8810 ( .A1(n9234), .A2(n7032), .ZN(n8170) );
  INV_X1 U8811 ( .A(n4462), .ZN(n8789) );
  NAND2_X1 U8812 ( .A1(n7159), .A2(n7469), .ZN(n7468) );
  XNOR2_X1 U8813 ( .A(n7028), .B(n7468), .ZN(n7035) );
  NAND2_X1 U8814 ( .A1(n8789), .A2(n8651), .ZN(n8610) );
  NAND2_X1 U8815 ( .A1(n6954), .A2(n9264), .ZN(n7033) );
  OAI21_X1 U8816 ( .B1(n8822), .B2(n9231), .A(n7033), .ZN(n7034) );
  AOI21_X1 U8817 ( .B1(n7035), .B2(n9269), .A(n7034), .ZN(n7624) );
  NAND2_X1 U8818 ( .A1(n7037), .A2(n7469), .ZN(n7036) );
  AOI22_X1 U8819 ( .A1(n7623), .A2(n10231), .B1(n10230), .B2(n7037), .ZN(n7038) );
  OAI211_X1 U8820 ( .C1(n7620), .C2(n10235), .A(n7624), .B(n7038), .ZN(n7130)
         );
  NAND2_X1 U8821 ( .A1(n7130), .A2(n10281), .ZN(n7039) );
  OAI21_X1 U8822 ( .B1(n10281), .B2(n7040), .A(n7039), .ZN(P2_U3454) );
  INV_X1 U8823 ( .A(n7511), .ZN(n7333) );
  OAI222_X1 U8824 ( .A1(n9831), .A2(n7042), .B1(n9835), .B2(n7041), .C1(
        P1_U3084), .C2(n7333), .ZN(P1_U3341) );
  INV_X1 U8825 ( .A(n7043), .ZN(n7044) );
  AOI21_X1 U8826 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7048), .A(n7044), .ZN(
        n7047) );
  MUX2_X1 U8827 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7045), .S(n7183), .Z(n7046)
         );
  NAND2_X1 U8828 ( .A1(n7047), .A2(n7046), .ZN(n7182) );
  OAI21_X1 U8829 ( .B1(n7047), .B2(n7046), .A(n7182), .ZN(n7059) );
  OR2_X1 U8830 ( .A1(n7048), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7051) );
  INV_X1 U8831 ( .A(n7049), .ZN(n7050) );
  MUX2_X1 U8832 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7931), .S(n7183), .Z(n7052)
         );
  NAND2_X1 U8833 ( .A1(n7052), .A2(n7053), .ZN(n7178) );
  OAI21_X1 U8834 ( .B1(n7053), .B2(n7052), .A(n7178), .ZN(n7057) );
  NAND2_X1 U8835 ( .A1(n9860), .A2(n7183), .ZN(n7056) );
  NAND2_X1 U8836 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7902) );
  INV_X1 U8837 ( .A(n7902), .ZN(n7054) );
  AOI21_X1 U8838 ( .B1(n10176), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7054), .ZN(
        n7055) );
  OAI211_X1 U8839 ( .C1(n7057), .C2(n8990), .A(n7056), .B(n7055), .ZN(n7058)
         );
  AOI21_X1 U8840 ( .B1(n7059), .B2(n10174), .A(n7058), .ZN(n7060) );
  INV_X1 U8841 ( .A(n7060), .ZN(P2_U3257) );
  OAI22_X1 U8842 ( .A1(n7062), .A2(n7061), .B1(n7071), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7065) );
  AOI22_X1 U8843 ( .A1(n7171), .A2(P1_REG1_REG_10__SCAN_IN), .B1(n5970), .B2(
        n7063), .ZN(n7064) );
  NAND2_X1 U8844 ( .A1(n7064), .A2(n7065), .ZN(n7170) );
  OAI21_X1 U8845 ( .B1(n7065), .B2(n7064), .A(n7170), .ZN(n7077) );
  INV_X1 U8846 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7069) );
  NAND2_X1 U8847 ( .A1(n10012), .A2(n7171), .ZN(n7068) );
  NOR2_X1 U8848 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7066), .ZN(n7713) );
  INV_X1 U8849 ( .A(n7713), .ZN(n7067) );
  OAI211_X1 U8850 ( .C1(n9999), .C2(n7069), .A(n7068), .B(n7067), .ZN(n7076)
         );
  NAND2_X1 U8851 ( .A1(n7171), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7072) );
  OAI21_X1 U8852 ( .B1(n7171), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7072), .ZN(
        n7073) );
  AOI211_X1 U8853 ( .C1(n7074), .C2(n7073), .A(n10003), .B(n7164), .ZN(n7075)
         );
  AOI211_X1 U8854 ( .C1(n10010), .C2(n7077), .A(n7076), .B(n7075), .ZN(n7078)
         );
  INV_X1 U8855 ( .A(n7078), .ZN(P1_U3251) );
  AND2_X1 U8856 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8889) );
  OAI211_X1 U8857 ( .C1(n7081), .C2(n7080), .A(n10174), .B(n7079), .ZN(n7082)
         );
  INV_X1 U8858 ( .A(n7082), .ZN(n7083) );
  AOI211_X1 U8859 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n10176), .A(n8889), .B(
        n7083), .ZN(n7088) );
  INV_X1 U8860 ( .A(n8990), .ZN(n10177) );
  OAI211_X1 U8861 ( .C1(n7086), .C2(n7085), .A(n10177), .B(n7084), .ZN(n7087)
         );
  OAI211_X1 U8862 ( .C1(n10178), .C2(n7089), .A(n7088), .B(n7087), .ZN(
        P2_U3251) );
  NOR2_X1 U8863 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7090), .ZN(n7096) );
  OAI211_X1 U8864 ( .C1(n7093), .C2(n7092), .A(n10174), .B(n7091), .ZN(n7094)
         );
  INV_X1 U8865 ( .A(n7094), .ZN(n7095) );
  AOI211_X1 U8866 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n10176), .A(n7096), .B(
        n7095), .ZN(n7102) );
  OR3_X1 U8867 ( .A1(n7111), .A2(n7098), .A3(n7097), .ZN(n7099) );
  NAND3_X1 U8868 ( .A1(n10177), .A2(n7100), .A3(n7099), .ZN(n7101) );
  OAI211_X1 U8869 ( .C1(n10178), .C2(n7103), .A(n7102), .B(n7101), .ZN(
        P2_U3249) );
  INV_X1 U8870 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7104) );
  NOR2_X1 U8871 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7104), .ZN(n7110) );
  OAI211_X1 U8872 ( .C1(n7107), .C2(n7106), .A(n10174), .B(n7105), .ZN(n7108)
         );
  INV_X1 U8873 ( .A(n7108), .ZN(n7109) );
  AOI211_X1 U8874 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n10176), .A(n7110), .B(
        n7109), .ZN(n7117) );
  INV_X1 U8875 ( .A(n7111), .ZN(n7115) );
  NAND3_X1 U8876 ( .A1(n9861), .A2(n7113), .A3(n7112), .ZN(n7114) );
  NAND3_X1 U8877 ( .A1(n10177), .A2(n7115), .A3(n7114), .ZN(n7116) );
  OAI211_X1 U8878 ( .C1(n10178), .C2(n7118), .A(n7117), .B(n7116), .ZN(
        P2_U3248) );
  XOR2_X1 U8879 ( .A(n7119), .B(n7120), .Z(n7125) );
  INV_X1 U8880 ( .A(n9472), .ZN(n8130) );
  AOI22_X1 U8881 ( .A1(n9475), .A2(n5785), .B1(n8130), .B2(n7261), .ZN(n7124)
         );
  NOR2_X1 U8882 ( .A1(n9473), .A2(n7364), .ZN(n7121) );
  AOI211_X1 U8883 ( .C1(n9459), .C2(n10103), .A(n7122), .B(n7121), .ZN(n7123)
         );
  OAI211_X1 U8884 ( .C1(n7125), .C2(n9461), .A(n7124), .B(n7123), .ZN(P1_U3216) );
  NAND2_X1 U8885 ( .A1(n7127), .A2(n7126), .ZN(n7129) );
  INV_X1 U8886 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7132) );
  NAND2_X1 U8887 ( .A1(n7130), .A2(n4449), .ZN(n7131) );
  OAI21_X1 U8888 ( .B1(n4449), .B2(n7132), .A(n7131), .ZN(P2_U3521) );
  XNOR2_X1 U8889 ( .A(n7134), .B(n7133), .ZN(n7143) );
  AND2_X1 U8890 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7135) );
  AOI21_X1 U8891 ( .B1(n10176), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7135), .ZN(
        n7140) );
  OAI211_X1 U8892 ( .C1(n7138), .C2(n7137), .A(n10174), .B(n7136), .ZN(n7139)
         );
  OAI211_X1 U8893 ( .C1(n10178), .C2(n7141), .A(n7140), .B(n7139), .ZN(n7142)
         );
  AOI21_X1 U8894 ( .B1(n10177), .B2(n7143), .A(n7142), .ZN(n7144) );
  INV_X1 U8895 ( .A(n7144), .ZN(P2_U3252) );
  XOR2_X1 U8896 ( .A(n7146), .B(n7145), .Z(n7155) );
  NAND2_X1 U8897 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7667) );
  INV_X1 U8898 ( .A(n7667), .ZN(n7149) );
  NOR2_X1 U8899 ( .A1(n10178), .A2(n7147), .ZN(n7148) );
  AOI211_X1 U8900 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n10176), .A(n7149), .B(
        n7148), .ZN(n7154) );
  OAI211_X1 U8901 ( .C1(n7152), .C2(n7151), .A(n10174), .B(n7150), .ZN(n7153)
         );
  OAI211_X1 U8902 ( .C1(n7155), .C2(n8990), .A(n7154), .B(n7153), .ZN(P2_U3254) );
  NAND2_X1 U8903 ( .A1(n7207), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7158) );
  NAND2_X1 U8904 ( .A1(P2_U3152), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9840) );
  OAI211_X1 U8905 ( .C1(n8856), .C2(n7619), .A(n7158), .B(n9840), .ZN(n7161)
         );
  OAI22_X1 U8906 ( .A1(n8822), .A2(n8887), .B1(n8875), .B2(n7159), .ZN(n7160)
         );
  AOI211_X1 U8907 ( .C1(n8882), .C2(n7162), .A(n7161), .B(n7160), .ZN(n7163)
         );
  INV_X1 U8908 ( .A(n7163), .ZN(P2_U3224) );
  AOI22_X1 U8909 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7335), .B1(n7169), .B2(
        n7794), .ZN(n7166) );
  OAI21_X1 U8910 ( .B1(n7166), .B2(n7165), .A(n7334), .ZN(n7167) );
  INV_X1 U8911 ( .A(n7167), .ZN(n7177) );
  AND2_X1 U8912 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3084), .ZN(n7728) );
  NOR2_X1 U8913 ( .A1(n9525), .A2(n7169), .ZN(n7168) );
  AOI211_X1 U8914 ( .C1(P1_ADDR_REG_11__SCAN_IN), .C2(n10013), .A(n7728), .B(
        n7168), .ZN(n7176) );
  AOI22_X1 U8915 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n7335), .B1(n7169), .B2(
        n5988), .ZN(n7173) );
  OAI21_X1 U8916 ( .B1(n7171), .B2(P1_REG1_REG_10__SCAN_IN), .A(n7170), .ZN(
        n7172) );
  NAND2_X1 U8917 ( .A1(n7173), .A2(n7172), .ZN(n7328) );
  OAI21_X1 U8918 ( .B1(n7173), .B2(n7172), .A(n7328), .ZN(n7174) );
  NAND2_X1 U8919 ( .A1(n7174), .A2(n10010), .ZN(n7175) );
  OAI211_X1 U8920 ( .C1(n7177), .C2(n10003), .A(n7176), .B(n7175), .ZN(
        P1_U3252) );
  NAND2_X1 U8921 ( .A1(n7183), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7179) );
  NAND2_X1 U8922 ( .A1(n7179), .A2(n7178), .ZN(n7181) );
  INV_X1 U8923 ( .A(n7233), .ZN(n7192) );
  AOI22_X1 U8924 ( .A1(n7233), .A2(n7969), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7192), .ZN(n7180) );
  NOR2_X1 U8925 ( .A1(n7181), .A2(n7180), .ZN(n7228) );
  AOI21_X1 U8926 ( .B1(n7181), .B2(n7180), .A(n7228), .ZN(n7190) );
  AOI22_X1 U8927 ( .A1(n7233), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n5346), .B2(
        n7192), .ZN(n7185) );
  OAI21_X1 U8928 ( .B1(n7183), .B2(P2_REG1_REG_12__SCAN_IN), .A(n7182), .ZN(
        n7184) );
  NAND2_X1 U8929 ( .A1(n7185), .A2(n7184), .ZN(n7232) );
  OAI21_X1 U8930 ( .B1(n7185), .B2(n7184), .A(n7232), .ZN(n7188) );
  AOI22_X1 U8931 ( .A1(n10176), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3152), .ZN(n7186) );
  OAI21_X1 U8932 ( .B1(n10178), .B2(n7192), .A(n7186), .ZN(n7187) );
  AOI21_X1 U8933 ( .B1(n7188), .B2(n10174), .A(n7187), .ZN(n7189) );
  OAI21_X1 U8934 ( .B1(n7190), .B2(n8990), .A(n7189), .ZN(P2_U3258) );
  INV_X1 U8935 ( .A(n7191), .ZN(n7203) );
  OAI222_X1 U8936 ( .A1(n9379), .A2(n7193), .B1(n4451), .B2(n7203), .C1(n7192), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8937 ( .A(n7194), .ZN(n7212) );
  INV_X1 U8938 ( .A(n8000), .ZN(n7994) );
  OAI222_X1 U8939 ( .A1(n9835), .A2(n7212), .B1(n7994), .B2(P1_U3084), .C1(
        n7195), .C2(n9831), .ZN(P1_U3339) );
  XOR2_X1 U8940 ( .A(n7197), .B(n7196), .Z(n7202) );
  INV_X1 U8941 ( .A(n7397), .ZN(n7198) );
  AOI22_X1 U8942 ( .A1(n9475), .A2(n9498), .B1(n8130), .B2(n7198), .ZN(n7201)
         );
  AND2_X1 U8943 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9996) );
  NOR2_X1 U8944 ( .A1(n9473), .A2(n7557), .ZN(n7199) );
  AOI211_X1 U8945 ( .C1(n9459), .C2(n7399), .A(n9996), .B(n7199), .ZN(n7200)
         );
  OAI211_X1 U8946 ( .C1(n7202), .C2(n9461), .A(n7201), .B(n7200), .ZN(P1_U3228) );
  INV_X1 U8947 ( .A(n7741), .ZN(n7509) );
  OAI222_X1 U8948 ( .A1(n9831), .A2(n7204), .B1(n7509), .B2(P1_U3084), .C1(
        n9835), .C2(n7203), .ZN(P1_U3340) );
  INV_X1 U8949 ( .A(n8820), .ZN(n7205) );
  AOI211_X1 U8950 ( .C1(n7206), .C2(n4923), .A(n8868), .B(n7205), .ZN(n7211)
         );
  INV_X1 U8951 ( .A(n8887), .ZN(n8097) );
  INV_X1 U8952 ( .A(n8875), .ZN(n8894) );
  AOI22_X1 U8953 ( .A1(n8097), .A2(n8912), .B1(n8894), .B2(n7025), .ZN(n7209)
         );
  NOR2_X1 U8954 ( .A1(n7434), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9853) );
  AOI21_X1 U8955 ( .B1(n7207), .B2(P2_REG3_REG_2__SCAN_IN), .A(n9853), .ZN(
        n7208) );
  OAI211_X1 U8956 ( .C1(n7268), .C2(n8856), .A(n7209), .B(n7208), .ZN(n7210)
         );
  OR2_X1 U8957 ( .A1(n7211), .A2(n7210), .ZN(P2_U3239) );
  INV_X1 U8958 ( .A(n7412), .ZN(n7237) );
  OAI222_X1 U8959 ( .A1(n9379), .A2(n7213), .B1(n4451), .B2(n7212), .C1(n7237), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  OAI21_X1 U8960 ( .B1(n7216), .B2(n7214), .A(n7215), .ZN(n7226) );
  INV_X1 U8961 ( .A(n7216), .ZN(n7218) );
  NAND4_X1 U8962 ( .A1(n7218), .A2(n8857), .A3(n7217), .A4(n8912), .ZN(n7224)
         );
  INV_X1 U8963 ( .A(n7565), .ZN(n8910) );
  AOI22_X1 U8964 ( .A1(n8910), .A2(n9266), .B1(n9264), .B2(n8912), .ZN(n7458)
         );
  INV_X1 U8965 ( .A(n7458), .ZN(n7220) );
  AOI22_X1 U8966 ( .A1(n7220), .A2(n7219), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n7223) );
  OR2_X1 U8967 ( .A1(n8885), .A2(n7599), .ZN(n7222) );
  INV_X1 U8968 ( .A(n7460), .ZN(n7600) );
  OR2_X1 U8969 ( .A1(n8856), .A2(n7600), .ZN(n7221) );
  NAND4_X1 U8970 ( .A1(n7224), .A2(n7223), .A3(n7222), .A4(n7221), .ZN(n7225)
         );
  AOI21_X1 U8971 ( .B1(n7226), .B2(n8882), .A(n7225), .ZN(n7227) );
  INV_X1 U8972 ( .A(n7227), .ZN(P2_U3232) );
  NOR2_X1 U8973 ( .A1(n7233), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7229) );
  NOR2_X1 U8974 ( .A1(n7229), .A2(n7228), .ZN(n7231) );
  AOI22_X1 U8975 ( .A1(n7412), .A2(n8015), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7237), .ZN(n7230) );
  NOR2_X1 U8976 ( .A1(n7231), .A2(n7230), .ZN(n7406) );
  AOI21_X1 U8977 ( .B1(n7231), .B2(n7230), .A(n7406), .ZN(n7241) );
  AOI22_X1 U8978 ( .A1(n7412), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n5367), .B2(
        n7237), .ZN(n7235) );
  OAI21_X1 U8979 ( .B1(n7233), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7232), .ZN(
        n7234) );
  NAND2_X1 U8980 ( .A1(n7235), .A2(n7234), .ZN(n7411) );
  OAI21_X1 U8981 ( .B1(n7235), .B2(n7234), .A(n7411), .ZN(n7239) );
  NAND2_X1 U8982 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8098) );
  NAND2_X1 U8983 ( .A1(n10176), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7236) );
  OAI211_X1 U8984 ( .C1(n10178), .C2(n7237), .A(n8098), .B(n7236), .ZN(n7238)
         );
  AOI21_X1 U8985 ( .B1(n7239), .B2(n10174), .A(n7238), .ZN(n7240) );
  OAI21_X1 U8986 ( .B1(n7241), .B2(n8990), .A(n7240), .ZN(P2_U3259) );
  NAND2_X1 U8987 ( .A1(n7243), .A2(n7242), .ZN(n7376) );
  INV_X2 U8988 ( .A(n10057), .ZN(n9738) );
  NOR2_X1 U8989 ( .A1(n7244), .A2(n8549), .ZN(n10042) );
  INV_X1 U8990 ( .A(n7245), .ZN(n7246) );
  NAND2_X1 U8991 ( .A1(n10057), .A2(n7246), .ZN(n10019) );
  AOI21_X1 U8992 ( .B1(n9724), .B2(n10019), .A(n7295), .ZN(n7249) );
  INV_X1 U8993 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9944) );
  INV_X1 U8994 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7247) );
  OAI22_X1 U8995 ( .A1(n10031), .A2(n9944), .B1(n7247), .B2(n10036), .ZN(n7248) );
  NOR2_X1 U8996 ( .A1(n7249), .A2(n7248), .ZN(n7250) );
  OAI21_X1 U8997 ( .B1(n7251), .B2(n9738), .A(n7250), .ZN(P1_U3291) );
  XNOR2_X1 U8998 ( .A(n7252), .B(n7255), .ZN(n7256) );
  INV_X1 U8999 ( .A(n7256), .ZN(n10107) );
  NAND2_X1 U9000 ( .A1(n7253), .A2(n10044), .ZN(n10037) );
  NOR2_X1 U9001 ( .A1(n9738), .A2(n10037), .ZN(n7402) );
  INV_X1 U9002 ( .A(n7402), .ZN(n7303) );
  XNOR2_X1 U9003 ( .A(n7255), .B(n7254), .ZN(n7259) );
  INV_X1 U9004 ( .A(n10128), .ZN(n7391) );
  NAND2_X1 U9005 ( .A1(n7256), .A2(n7391), .ZN(n7258) );
  AOI22_X1 U9006 ( .A1(n9497), .A2(n10046), .B1(n10045), .B2(n5785), .ZN(n7257) );
  OAI211_X1 U9007 ( .C1(n7259), .C2(n6466), .A(n7258), .B(n7257), .ZN(n10109)
         );
  NAND2_X1 U9008 ( .A1(n10109), .A2(n10031), .ZN(n7267) );
  INV_X1 U9009 ( .A(n10019), .ZN(n9682) );
  NAND2_X1 U9010 ( .A1(n7297), .A2(n10103), .ZN(n7260) );
  AND2_X1 U9011 ( .A1(n7394), .A2(n7260), .ZN(n10104) );
  OAI22_X1 U9012 ( .A1(n10057), .A2(n7262), .B1(n10036), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n7265) );
  NOR2_X1 U9013 ( .A1(n9724), .A2(n7263), .ZN(n7264) );
  AOI211_X1 U9014 ( .C1(n9682), .C2(n10104), .A(n7265), .B(n7264), .ZN(n7266)
         );
  OAI211_X1 U9015 ( .C1(n10107), .C2(n7303), .A(n7267), .B(n7266), .ZN(
        P1_U3288) );
  NAND2_X1 U9016 ( .A1(n8822), .A2(n7436), .ZN(n8659) );
  NAND2_X1 U9017 ( .A1(n7026), .A2(n7619), .ZN(n7269) );
  NAND2_X1 U9018 ( .A1(n8822), .A2(n7268), .ZN(n7440) );
  NAND2_X1 U9019 ( .A1(n7442), .A2(n7440), .ZN(n7271) );
  INV_X1 U9020 ( .A(n7592), .ZN(n7282) );
  INV_X1 U9021 ( .A(n8170), .ZN(n7682) );
  NAND2_X1 U9022 ( .A1(n8658), .A2(n7468), .ZN(n8612) );
  NAND2_X1 U9023 ( .A1(n7272), .A2(n8612), .ZN(n7423) );
  INV_X1 U9024 ( .A(n7423), .ZN(n7274) );
  INV_X1 U9025 ( .A(n8613), .ZN(n7273) );
  NAND2_X1 U9026 ( .A1(n7274), .A2(n7273), .ZN(n7425) );
  NAND2_X1 U9027 ( .A1(n7425), .A2(n8659), .ZN(n7454) );
  AOI22_X1 U9028 ( .A1(n9264), .A2(n7275), .B1(n8911), .B2(n9266), .ZN(n7276)
         );
  OAI21_X1 U9029 ( .B1(n7277), .B2(n9228), .A(n7276), .ZN(n7278) );
  AOI21_X1 U9030 ( .B1(n7682), .B2(n7592), .A(n7278), .ZN(n7594) );
  INV_X1 U9031 ( .A(n8826), .ZN(n7452) );
  INV_X1 U9032 ( .A(n7279), .ZN(n7432) );
  NAND2_X1 U9033 ( .A1(n7279), .A2(n8826), .ZN(n7451) );
  INV_X1 U9034 ( .A(n7451), .ZN(n7280) );
  AOI21_X1 U9035 ( .B1(n7452), .B2(n7432), .A(n7280), .ZN(n7589) );
  AOI22_X1 U9036 ( .A1(n7589), .A2(n10231), .B1(n10230), .B2(n7452), .ZN(n7281) );
  OAI211_X1 U9037 ( .C1(n7282), .C2(n10245), .A(n7594), .B(n7281), .ZN(n7285)
         );
  NAND2_X1 U9038 ( .A1(n7285), .A2(n10281), .ZN(n7283) );
  OAI21_X1 U9039 ( .B1(n10281), .B2(n7284), .A(n7283), .ZN(P2_U3460) );
  NAND2_X1 U9040 ( .A1(n7285), .A2(n4449), .ZN(n7286) );
  OAI21_X1 U9041 ( .B1(n4449), .B2(n6983), .A(n7286), .ZN(P2_U3523) );
  XNOR2_X1 U9042 ( .A(n7287), .B(n8252), .ZN(n10097) );
  XNOR2_X1 U9043 ( .A(n8506), .B(n8252), .ZN(n7291) );
  OAI22_X1 U9044 ( .A1(n7289), .A2(n6463), .B1(n7387), .B2(n9716), .ZN(n7290)
         );
  AOI21_X1 U9045 ( .B1(n7291), .B2(n10050), .A(n7290), .ZN(n7292) );
  OAI21_X1 U9046 ( .B1(n10097), .B2(n10128), .A(n7292), .ZN(n10100) );
  NAND2_X1 U9047 ( .A1(n10100), .A2(n10031), .ZN(n7302) );
  INV_X1 U9048 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7294) );
  OAI22_X1 U9049 ( .A1(n10057), .A2(n7294), .B1(n7293), .B2(n10036), .ZN(n7300) );
  NAND2_X1 U9050 ( .A1(n7295), .A2(n10092), .ZN(n7296) );
  NAND2_X1 U9051 ( .A1(n4969), .A2(n7296), .ZN(n7298) );
  NAND2_X1 U9052 ( .A1(n7298), .A2(n7297), .ZN(n10099) );
  NOR2_X1 U9053 ( .A1(n10019), .A2(n10099), .ZN(n7299) );
  AOI211_X1 U9054 ( .C1(n9739), .C2(n4969), .A(n7300), .B(n7299), .ZN(n7301)
         );
  OAI211_X1 U9055 ( .C1(n10097), .C2(n7303), .A(n7302), .B(n7301), .ZN(
        P1_U3289) );
  INV_X1 U9056 ( .A(n7304), .ZN(n7305) );
  AOI21_X1 U9057 ( .B1(n8359), .B2(n7306), .A(n7305), .ZN(n10129) );
  NAND2_X1 U9058 ( .A1(n10128), .A2(n10037), .ZN(n10027) );
  AOI21_X1 U9059 ( .B1(n7547), .B2(n7348), .A(n4687), .ZN(n10125) );
  INV_X1 U9060 ( .A(n7556), .ZN(n7307) );
  INV_X1 U9061 ( .A(n10036), .ZN(n10041) );
  AOI22_X1 U9062 ( .A1(n9738), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7307), .B2(
        n10041), .ZN(n7308) );
  OAI21_X1 U9063 ( .B1(n7309), .B2(n9724), .A(n7308), .ZN(n7310) );
  AOI21_X1 U9064 ( .B1(n10125), .B2(n9682), .A(n7310), .ZN(n7316) );
  NAND2_X1 U9065 ( .A1(n8356), .A2(n8354), .ZN(n7311) );
  NAND2_X1 U9066 ( .A1(n7311), .A2(n8353), .ZN(n8357) );
  XNOR2_X1 U9067 ( .A(n8357), .B(n8359), .ZN(n7312) );
  NAND2_X1 U9068 ( .A1(n7312), .A2(n10050), .ZN(n7314) );
  AOI22_X1 U9069 ( .A1(n9496), .A2(n10045), .B1(n10046), .B2(n9493), .ZN(n7313) );
  NAND2_X1 U9070 ( .A1(n7314), .A2(n7313), .ZN(n10131) );
  NAND2_X1 U9071 ( .A1(n10131), .A2(n10031), .ZN(n7315) );
  OAI211_X1 U9072 ( .C1(n10129), .C2(n9746), .A(n7316), .B(n7315), .ZN(
        P1_U3285) );
  XNOR2_X1 U9073 ( .A(n7317), .B(n7318), .ZN(n7319) );
  NAND2_X1 U9074 ( .A1(n7319), .A2(n9467), .ZN(n7323) );
  OAI22_X1 U9075 ( .A1(n9455), .A2(n7344), .B1(n9472), .B2(n7374), .ZN(n7320)
         );
  AOI211_X1 U9076 ( .C1(n8126), .C2(n10022), .A(n7321), .B(n7320), .ZN(n7322)
         );
  OAI211_X1 U9077 ( .C1(n10137), .C2(n9478), .A(n7323), .B(n7322), .ZN(
        P1_U3211) );
  INV_X1 U9078 ( .A(n7324), .ZN(n7326) );
  INV_X1 U9079 ( .A(n7939), .ZN(n7947) );
  OAI222_X1 U9080 ( .A1(n9379), .A2(n7325), .B1(n4451), .B2(n7326), .C1(
        P2_U3152), .C2(n7947), .ZN(P2_U3343) );
  OAI222_X1 U9081 ( .A1(n9831), .A2(n7327), .B1(n9835), .B2(n7326), .C1(
        P1_U3084), .C2(n8080), .ZN(P1_U3338) );
  OAI21_X1 U9082 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n7335), .A(n7328), .ZN(
        n7331) );
  MUX2_X1 U9083 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7329), .S(n7511), .Z(n7330)
         );
  NAND2_X1 U9084 ( .A1(n7330), .A2(n7331), .ZN(n7503) );
  OAI21_X1 U9085 ( .B1(n7331), .B2(n7330), .A(n7503), .ZN(n7341) );
  NAND2_X1 U9086 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n7777) );
  NAND2_X1 U9087 ( .A1(n10013), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n7332) );
  OAI211_X1 U9088 ( .C1(n9525), .C2(n7333), .A(n7777), .B(n7332), .ZN(n7340)
         );
  OAI21_X1 U9089 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7335), .A(n7334), .ZN(
        n7338) );
  NAND2_X1 U9090 ( .A1(n7511), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7336) );
  OAI21_X1 U9091 ( .B1(n7511), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7336), .ZN(
        n7337) );
  NOR2_X1 U9092 ( .A1(n7337), .A2(n7338), .ZN(n7510) );
  AOI211_X1 U9093 ( .C1(n7338), .C2(n7337), .A(n7510), .B(n10003), .ZN(n7339)
         );
  AOI211_X1 U9094 ( .C1(n10010), .C2(n7341), .A(n7340), .B(n7339), .ZN(n7342)
         );
  INV_X1 U9095 ( .A(n7342), .ZN(P1_U3253) );
  XOR2_X1 U9096 ( .A(n7353), .B(n8356), .Z(n7343) );
  OAI222_X1 U9097 ( .A1(n6463), .A2(n7364), .B1(n9716), .B2(n7344), .C1(n7343), 
        .C2(n6466), .ZN(n10123) );
  INV_X1 U9098 ( .A(n10123), .ZN(n7357) );
  INV_X1 U9099 ( .A(n7345), .ZN(n7363) );
  OAI22_X1 U9100 ( .A1(n10031), .A2(n7346), .B1(n7363), .B2(n10036), .ZN(n7350) );
  OR2_X1 U9101 ( .A1(n7395), .A2(n7367), .ZN(n7347) );
  NAND2_X1 U9102 ( .A1(n7348), .A2(n7347), .ZN(n10119) );
  NOR2_X1 U9103 ( .A1(n10119), .A2(n10019), .ZN(n7349) );
  AOI211_X1 U9104 ( .C1(n9739), .C2(n7351), .A(n7350), .B(n7349), .ZN(n7356)
         );
  NAND2_X1 U9105 ( .A1(n7354), .A2(n7353), .ZN(n10118) );
  NAND3_X1 U9106 ( .A1(n7352), .A2(n10118), .A3(n9611), .ZN(n7355) );
  OAI211_X1 U9107 ( .C1(n7357), .C2(n9738), .A(n7356), .B(n7355), .ZN(P1_U3286) );
  INV_X1 U9108 ( .A(n7358), .ZN(n7383) );
  INV_X1 U9109 ( .A(n8961), .ZN(n7945) );
  OAI222_X1 U9110 ( .A1(n9379), .A2(n7359), .B1(n4451), .B2(n7383), .C1(n7945), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  XNOR2_X1 U9111 ( .A(n7360), .B(n7549), .ZN(n7362) );
  NOR2_X1 U9112 ( .A1(n7362), .A2(n7361), .ZN(n7548) );
  AOI21_X1 U9113 ( .B1(n7362), .B2(n7361), .A(n7548), .ZN(n7370) );
  OAI22_X1 U9114 ( .A1(n9455), .A2(n7364), .B1(n9472), .B2(n7363), .ZN(n7365)
         );
  AOI211_X1 U9115 ( .C1(n8126), .C2(n9495), .A(n7366), .B(n7365), .ZN(n7369)
         );
  NOR2_X1 U9116 ( .A1(n7367), .A2(n10136), .ZN(n10122) );
  NAND2_X1 U9117 ( .A1(n9430), .A2(n10122), .ZN(n7368) );
  OAI211_X1 U9118 ( .C1(n7370), .C2(n9461), .A(n7369), .B(n7368), .ZN(P1_U3225) );
  OAI21_X1 U9119 ( .B1(n4585), .B2(n4584), .A(n7372), .ZN(n7373) );
  AOI222_X1 U9120 ( .A1(n10050), .A2(n7373), .B1(n10022), .B2(n10046), .C1(
        n9495), .C2(n10045), .ZN(n10135) );
  OAI22_X1 U9121 ( .A1(n10031), .A2(n7375), .B1(n7374), .B2(n10036), .ZN(n7378) );
  OAI211_X1 U9122 ( .C1(n4687), .C2(n10137), .A(n10124), .B(n7483), .ZN(n10134) );
  OR2_X1 U9123 ( .A1(n7376), .A2(n10044), .ZN(n8057) );
  NOR2_X1 U9124 ( .A1(n10134), .A2(n8057), .ZN(n7377) );
  AOI211_X1 U9125 ( .C1(n9739), .C2(n7379), .A(n7378), .B(n7377), .ZN(n7382)
         );
  XNOR2_X1 U9126 ( .A(n7380), .B(n8361), .ZN(n10139) );
  NAND2_X1 U9127 ( .A1(n10139), .A2(n9611), .ZN(n7381) );
  OAI211_X1 U9128 ( .C1(n10135), .C2(n9738), .A(n7382), .B(n7381), .ZN(
        P1_U3284) );
  INV_X1 U9129 ( .A(n9518), .ZN(n8089) );
  OAI222_X1 U9130 ( .A1(n9831), .A2(n7384), .B1(n8089), .B2(P1_U3084), .C1(
        n9835), .C2(n7383), .ZN(P1_U3337) );
  INV_X1 U9131 ( .A(n8255), .ZN(n7385) );
  XNOR2_X1 U9132 ( .A(n7386), .B(n7385), .ZN(n7389) );
  OAI22_X1 U9133 ( .A1(n7557), .A2(n9716), .B1(n7387), .B2(n6463), .ZN(n7388)
         );
  AOI21_X1 U9134 ( .B1(n7389), .B2(n10050), .A(n7388), .ZN(n7393) );
  XNOR2_X1 U9135 ( .A(n7390), .B(n8255), .ZN(n10114) );
  NAND2_X1 U9136 ( .A1(n10114), .A2(n7391), .ZN(n7392) );
  AND2_X1 U9137 ( .A1(n7393), .A2(n7392), .ZN(n10116) );
  AND2_X1 U9138 ( .A1(n7394), .A2(n7399), .ZN(n7396) );
  OR2_X1 U9139 ( .A1(n7396), .A2(n7395), .ZN(n10112) );
  OAI22_X1 U9140 ( .A1(n10057), .A2(n6781), .B1(n7397), .B2(n10036), .ZN(n7398) );
  AOI21_X1 U9141 ( .B1(n9739), .B2(n7399), .A(n7398), .ZN(n7400) );
  OAI21_X1 U9142 ( .B1(n10112), .B2(n10019), .A(n7400), .ZN(n7401) );
  AOI21_X1 U9143 ( .B1(n10114), .B2(n7402), .A(n7401), .ZN(n7403) );
  OAI21_X1 U9144 ( .B1(n10116), .B2(n9738), .A(n7403), .ZN(P1_U3287) );
  INV_X1 U9145 ( .A(n7404), .ZN(n7466) );
  AOI22_X1 U9146 ( .A1(n8971), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n9376), .ZN(n7405) );
  OAI21_X1 U9147 ( .B1(n7466), .B2(n4451), .A(n7405), .ZN(P2_U3341) );
  NOR2_X1 U9148 ( .A1(n7412), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7407) );
  NOR2_X1 U9149 ( .A1(n7407), .A2(n7406), .ZN(n7938) );
  XNOR2_X1 U9150 ( .A(n7938), .B(n7939), .ZN(n7408) );
  NOR2_X1 U9151 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7408), .ZN(n7940) );
  AOI21_X1 U9152 ( .B1(n7408), .B2(P2_REG2_REG_15__SCAN_IN), .A(n7940), .ZN(
        n7419) );
  AND2_X1 U9153 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7410) );
  NOR2_X1 U9154 ( .A1(n10178), .A2(n7947), .ZN(n7409) );
  AOI211_X1 U9155 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n10176), .A(n7410), .B(
        n7409), .ZN(n7418) );
  OAI21_X1 U9156 ( .B1(n7412), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7411), .ZN(
        n7946) );
  XNOR2_X1 U9157 ( .A(n7946), .B(n7947), .ZN(n7413) );
  INV_X1 U9158 ( .A(n7413), .ZN(n7416) );
  NOR2_X1 U9159 ( .A1(n7414), .A2(n7413), .ZN(n7948) );
  INV_X1 U9160 ( .A(n7948), .ZN(n7415) );
  OAI211_X1 U9161 ( .C1(n7416), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10174), .B(
        n7415), .ZN(n7417) );
  OAI211_X1 U9162 ( .C1(n7419), .C2(n8990), .A(n7418), .B(n7417), .ZN(P2_U3260) );
  INV_X1 U9163 ( .A(n10227), .ZN(n7439) );
  NAND2_X1 U9164 ( .A1(n7421), .A2(n7420), .ZN(n7430) );
  OR2_X1 U9165 ( .A1(n7422), .A2(n7032), .ZN(n7586) );
  NAND2_X1 U9166 ( .A1(n8170), .A2(n7586), .ZN(n10196) );
  NAND2_X1 U9167 ( .A1(n7423), .A2(n8613), .ZN(n7424) );
  NAND2_X1 U9168 ( .A1(n7425), .A2(n7424), .ZN(n7428) );
  NAND2_X1 U9169 ( .A1(n8912), .A2(n9266), .ZN(n7426) );
  OAI21_X1 U9170 ( .B1(n7026), .B2(n9233), .A(n7426), .ZN(n7427) );
  AOI21_X1 U9171 ( .B1(n7428), .B2(n9269), .A(n7427), .ZN(n10224) );
  MUX2_X1 U9172 ( .A(n7429), .B(n10224), .S(n9244), .Z(n7438) );
  INV_X1 U9173 ( .A(n7430), .ZN(n7431) );
  NAND2_X1 U9174 ( .A1(n7431), .A2(n7032), .ZN(n7598) );
  OAI21_X1 U9175 ( .B1(n7268), .B2(n7433), .A(n7432), .ZN(n10223) );
  OAI22_X1 U9176 ( .A1(n9218), .A2(n10223), .B1(n7434), .B2(n9241), .ZN(n7435)
         );
  AOI21_X1 U9177 ( .B1(n9246), .B2(n7436), .A(n7435), .ZN(n7437) );
  OAI211_X1 U9178 ( .C1(n7439), .C2(n9274), .A(n7438), .B(n7437), .ZN(P2_U3294) );
  INV_X1 U9179 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7463) );
  NAND2_X1 U9180 ( .A1(n4556), .A2(n8826), .ZN(n7444) );
  AND2_X1 U9181 ( .A1(n7440), .A2(n7444), .ZN(n7441) );
  NAND2_X1 U9182 ( .A1(n8827), .A2(n7460), .ZN(n8637) );
  OAI21_X1 U9183 ( .B1(n7447), .B2(n7455), .A(n7448), .ZN(n7449) );
  INV_X1 U9184 ( .A(n7449), .ZN(n7605) );
  OR2_X1 U9185 ( .A1(n7451), .A2(n7460), .ZN(n7497) );
  INV_X1 U9186 ( .A(n7497), .ZN(n7450) );
  AOI211_X1 U9187 ( .C1(n7460), .C2(n7451), .A(n10273), .B(n7450), .ZN(n7602)
         );
  XOR2_X1 U9188 ( .A(n8912), .B(n8826), .Z(n8655) );
  NAND2_X1 U9189 ( .A1(n4556), .A2(n7452), .ZN(n8646) );
  AOI21_X1 U9190 ( .B1(n8655), .B2(n7454), .A(n7453), .ZN(n7457) );
  NAND2_X1 U9191 ( .A1(n7457), .A2(n7456), .ZN(n7524) );
  OAI211_X1 U9192 ( .C1(n7457), .C2(n7456), .A(n7524), .B(n9269), .ZN(n7459)
         );
  NAND2_X1 U9193 ( .A1(n7459), .A2(n7458), .ZN(n7595) );
  AOI211_X1 U9194 ( .C1(n10230), .C2(n7460), .A(n7602), .B(n7595), .ZN(n7461)
         );
  OAI21_X1 U9195 ( .B1(n10235), .B2(n7605), .A(n7461), .ZN(n7464) );
  NAND2_X1 U9196 ( .A1(n7464), .A2(n10281), .ZN(n7462) );
  OAI21_X1 U9197 ( .B1(n10281), .B2(n7463), .A(n7462), .ZN(P2_U3463) );
  NAND2_X1 U9198 ( .A1(n7464), .A2(n4449), .ZN(n7465) );
  OAI21_X1 U9199 ( .B1(n4449), .B2(n6984), .A(n7465), .ZN(P2_U3524) );
  INV_X1 U9200 ( .A(n9537), .ZN(n9524) );
  OAI222_X1 U9201 ( .A1(n9831), .A2(n7467), .B1(n9524), .B2(P1_U3084), .C1(
        n9835), .C2(n7466), .ZN(P1_U3336) );
  NAND2_X1 U9202 ( .A1(n6954), .A2(n10217), .ZN(n8650) );
  AND2_X1 U9203 ( .A1(n7468), .A2(n8650), .ZN(n10219) );
  OAI21_X1 U9204 ( .B1(n9272), .B2(n9246), .A(n7469), .ZN(n7473) );
  OAI22_X1 U9205 ( .A1(n10219), .A2(n9228), .B1(n7026), .B2(n9231), .ZN(n10221) );
  INV_X2 U9206 ( .A(n9238), .ZN(n10198) );
  OAI22_X1 U9207 ( .A1(n9244), .A2(n4945), .B1(n7470), .B2(n9241), .ZN(n7471)
         );
  AOI21_X1 U9208 ( .B1(n10221), .B2(n9238), .A(n7471), .ZN(n7472) );
  OAI211_X1 U9209 ( .C1(n10219), .C2(n9274), .A(n7473), .B(n7472), .ZN(
        P2_U3296) );
  INV_X1 U9210 ( .A(n7478), .ZN(n8258) );
  XNOR2_X1 U9211 ( .A(n7474), .B(n8258), .ZN(n7475) );
  NAND2_X1 U9212 ( .A1(n7475), .A2(n10050), .ZN(n7477) );
  AOI22_X1 U9213 ( .A1(n9492), .A2(n10046), .B1(n10045), .B2(n9493), .ZN(n7476) );
  NAND2_X1 U9214 ( .A1(n7477), .A2(n7476), .ZN(n10146) );
  INV_X1 U9215 ( .A(n10146), .ZN(n7491) );
  NOR2_X1 U9216 ( .A1(n7479), .A2(n7478), .ZN(n10142) );
  INV_X1 U9217 ( .A(n10142), .ZN(n7481) );
  NAND3_X1 U9218 ( .A1(n7481), .A2(n9611), .A3(n7480), .ZN(n7490) );
  OAI22_X1 U9219 ( .A1(n10057), .A2(n7482), .B1(n7542), .B2(n10036), .ZN(n7488) );
  INV_X1 U9220 ( .A(n7535), .ZN(n7486) );
  INV_X1 U9221 ( .A(n7483), .ZN(n7485) );
  INV_X1 U9222 ( .A(n10017), .ZN(n7484) );
  OAI21_X1 U9223 ( .B1(n7486), .B2(n7485), .A(n7484), .ZN(n10144) );
  NOR2_X1 U9224 ( .A1(n10144), .A2(n10019), .ZN(n7487) );
  AOI211_X1 U9225 ( .C1(n9739), .C2(n7535), .A(n7488), .B(n7487), .ZN(n7489)
         );
  OAI211_X1 U9226 ( .C1(n9738), .C2(n7491), .A(n7490), .B(n7489), .ZN(P1_U3283) );
  INV_X1 U9227 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7501) );
  NAND2_X1 U9228 ( .A1(n8827), .A2(n7600), .ZN(n7492) );
  NAND2_X1 U9229 ( .A1(n7565), .A2(n10187), .ZN(n8648) );
  NAND2_X1 U9230 ( .A1(n8648), .A2(n8643), .ZN(n8614) );
  OAI21_X1 U9231 ( .B1(n7494), .B2(n8614), .A(n7522), .ZN(n10195) );
  INV_X1 U9232 ( .A(n10195), .ZN(n7499) );
  NAND2_X1 U9233 ( .A1(n7524), .A2(n8639), .ZN(n7495) );
  XNOR2_X1 U9234 ( .A(n7495), .B(n8614), .ZN(n7496) );
  AOI222_X1 U9235 ( .A1(n9269), .A2(n7496), .B1(n8909), .B2(n9266), .C1(n8911), 
        .C2(n9264), .ZN(n10192) );
  AOI211_X1 U9236 ( .C1(n10187), .C2(n7497), .A(n10273), .B(n7569), .ZN(n10185) );
  AOI21_X1 U9237 ( .B1(n10230), .B2(n10187), .A(n10185), .ZN(n7498) );
  OAI211_X1 U9238 ( .C1(n10235), .C2(n7499), .A(n10192), .B(n7498), .ZN(n7518)
         );
  NAND2_X1 U9239 ( .A1(n7518), .A2(n10281), .ZN(n7500) );
  OAI21_X1 U9240 ( .B1(n10281), .B2(n7501), .A(n7500), .ZN(P2_U3466) );
  MUX2_X1 U9241 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7502), .S(n7741), .Z(n7505)
         );
  OAI21_X1 U9242 ( .B1(n7511), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7503), .ZN(
        n7504) );
  NAND2_X1 U9243 ( .A1(n7505), .A2(n7504), .ZN(n7736) );
  OAI21_X1 U9244 ( .B1(n7505), .B2(n7504), .A(n7736), .ZN(n7516) );
  NOR2_X1 U9245 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7506), .ZN(n7914) );
  INV_X1 U9246 ( .A(n7914), .ZN(n7508) );
  NAND2_X1 U9247 ( .A1(n10013), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n7507) );
  OAI211_X1 U9248 ( .C1(n9525), .C2(n7509), .A(n7508), .B(n7507), .ZN(n7515)
         );
  MUX2_X1 U9249 ( .A(n7812), .B(P1_REG2_REG_13__SCAN_IN), .S(n7741), .Z(n7512)
         );
  AOI211_X1 U9250 ( .C1(n7513), .C2(n7512), .A(n10003), .B(n7740), .ZN(n7514)
         );
  AOI211_X1 U9251 ( .C1(n10010), .C2(n7516), .A(n7515), .B(n7514), .ZN(n7517)
         );
  INV_X1 U9252 ( .A(n7517), .ZN(P1_U3254) );
  NAND2_X1 U9253 ( .A1(n7518), .A2(n4449), .ZN(n7519) );
  OAI21_X1 U9254 ( .B1(n4449), .B2(n6988), .A(n7519), .ZN(P2_U3525) );
  NAND2_X1 U9255 ( .A1(n7565), .A2(n7520), .ZN(n7521) );
  NAND2_X1 U9256 ( .A1(n7562), .A2(n7571), .ZN(n7523) );
  XNOR2_X1 U9257 ( .A(n8908), .B(n10239), .ZN(n8676) );
  XNOR2_X1 U9258 ( .A(n7639), .B(n8676), .ZN(n10243) );
  INV_X1 U9259 ( .A(n10243), .ZN(n7534) );
  NAND2_X1 U9260 ( .A1(n7524), .A2(n8638), .ZN(n7525) );
  NAND2_X1 U9261 ( .A1(n7525), .A2(n8648), .ZN(n7563) );
  NOR2_X1 U9262 ( .A1(n8909), .A2(n7571), .ZN(n8670) );
  INV_X1 U9263 ( .A(n8676), .ZN(n8619) );
  OAI211_X1 U9264 ( .C1(n7526), .C2(n8619), .A(n7646), .B(n9269), .ZN(n7528)
         );
  AOI22_X1 U9265 ( .A1(n9266), .A2(n8907), .B1(n8909), .B2(n9264), .ZN(n7527)
         );
  NAND2_X1 U9266 ( .A1(n7528), .A2(n7527), .ZN(n10241) );
  XNOR2_X1 U9267 ( .A(n7656), .B(n10239), .ZN(n10240) );
  INV_X1 U9268 ( .A(n10239), .ZN(n8671) );
  OAI22_X1 U9269 ( .A1(n9238), .A2(n7529), .B1(n7631), .B2(n9241), .ZN(n7530)
         );
  AOI21_X1 U9270 ( .B1(n9246), .B2(n8671), .A(n7530), .ZN(n7531) );
  OAI21_X1 U9271 ( .B1(n10240), .B2(n9218), .A(n7531), .ZN(n7532) );
  AOI21_X1 U9272 ( .B1(n10241), .B2(n9238), .A(n7532), .ZN(n7533) );
  OAI21_X1 U9273 ( .B1(n7534), .B2(n9274), .A(n7533), .ZN(P2_U3289) );
  NAND2_X1 U9274 ( .A1(n7535), .A2(n10149), .ZN(n10143) );
  NAND2_X1 U9275 ( .A1(n7537), .A2(n7536), .ZN(n7539) );
  XNOR2_X1 U9276 ( .A(n7539), .B(n7538), .ZN(n7540) );
  NAND2_X1 U9277 ( .A1(n7540), .A2(n9467), .ZN(n7546) );
  INV_X1 U9278 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7541) );
  NOR2_X1 U9279 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7541), .ZN(n9506) );
  OAI22_X1 U9280 ( .A1(n9455), .A2(n7543), .B1(n9472), .B2(n7542), .ZN(n7544)
         );
  AOI211_X1 U9281 ( .C1(n8126), .C2(n9492), .A(n9506), .B(n7544), .ZN(n7545)
         );
  OAI211_X1 U9282 ( .C1(n7561), .C2(n10143), .A(n7546), .B(n7545), .ZN(
        P1_U3219) );
  NAND2_X1 U9283 ( .A1(n7547), .A2(n10149), .ZN(n10127) );
  AOI21_X1 U9284 ( .B1(n7549), .B2(n7360), .A(n7548), .ZN(n7553) );
  XNOR2_X1 U9285 ( .A(n7551), .B(n7550), .ZN(n7552) );
  XNOR2_X1 U9286 ( .A(n7553), .B(n7552), .ZN(n7554) );
  NAND2_X1 U9287 ( .A1(n7554), .A2(n9467), .ZN(n7560) );
  NOR2_X1 U9288 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7555), .ZN(n10008) );
  OAI22_X1 U9289 ( .A1(n9455), .A2(n7557), .B1(n9472), .B2(n7556), .ZN(n7558)
         );
  AOI211_X1 U9290 ( .C1(n8126), .C2(n9493), .A(n10008), .B(n7558), .ZN(n7559)
         );
  OAI211_X1 U9291 ( .C1(n7561), .C2(n10127), .A(n7560), .B(n7559), .ZN(
        P1_U3237) );
  XNOR2_X1 U9292 ( .A(n7562), .B(n8620), .ZN(n10236) );
  XNOR2_X1 U9293 ( .A(n7563), .B(n8620), .ZN(n7567) );
  NAND2_X1 U9294 ( .A1(n8908), .A2(n9266), .ZN(n7564) );
  OAI21_X1 U9295 ( .B1(n7565), .B2(n9233), .A(n7564), .ZN(n7566) );
  AOI21_X1 U9296 ( .B1(n7567), .B2(n9269), .A(n7566), .ZN(n10234) );
  MUX2_X1 U9297 ( .A(n10234), .B(n7568), .S(n10198), .Z(n7574) );
  INV_X1 U9298 ( .A(n7569), .ZN(n7570) );
  AOI21_X1 U9299 ( .B1(n10229), .B2(n7570), .A(n7656), .ZN(n10232) );
  OAI22_X1 U9300 ( .A1(n9260), .A2(n7571), .B1(n9241), .B2(n8884), .ZN(n7572)
         );
  AOI21_X1 U9301 ( .B1(n10232), .B2(n9272), .A(n7572), .ZN(n7573) );
  OAI211_X1 U9302 ( .C1(n9274), .C2(n10236), .A(n7574), .B(n7573), .ZN(
        P2_U3290) );
  INV_X1 U9303 ( .A(n7575), .ZN(n7628) );
  INV_X1 U9304 ( .A(n7576), .ZN(n7577) );
  AOI21_X1 U9305 ( .B1(n7628), .B2(n7577), .A(n8868), .ZN(n7581) );
  INV_X1 U9306 ( .A(n8908), .ZN(n8886) );
  NOR3_X1 U9307 ( .A1(n8892), .A2(n7578), .A3(n8886), .ZN(n7580) );
  OAI21_X1 U9308 ( .B1(n7581), .B2(n7580), .A(n7579), .ZN(n7585) );
  OAI22_X1 U9309 ( .A1(n8885), .A2(n7654), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8926), .ZN(n7583) );
  OAI22_X1 U9310 ( .A1(n7754), .A2(n8887), .B1(n8875), .B2(n8886), .ZN(n7582)
         );
  AOI211_X1 U9311 ( .C1(n7672), .C2(n8890), .A(n7583), .B(n7582), .ZN(n7584)
         );
  NAND2_X1 U9312 ( .A1(n7585), .A2(n7584), .ZN(P2_U3223) );
  OR2_X1 U9313 ( .A1(n10198), .A2(n7586), .ZN(n9250) );
  INV_X1 U9314 ( .A(n9250), .ZN(n7691) );
  OAI22_X1 U9315 ( .A1(n9238), .A2(n7587), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9241), .ZN(n7588) );
  AOI21_X1 U9316 ( .B1(n7589), .B2(n9272), .A(n7588), .ZN(n7590) );
  OAI21_X1 U9317 ( .B1(n8826), .B2(n9260), .A(n7590), .ZN(n7591) );
  AOI21_X1 U9318 ( .B1(n7691), .B2(n7592), .A(n7591), .ZN(n7593) );
  OAI21_X1 U9319 ( .B1(n7594), .B2(n10198), .A(n7593), .ZN(P2_U3293) );
  INV_X1 U9320 ( .A(n7595), .ZN(n7597) );
  MUX2_X1 U9321 ( .A(n7597), .B(n7596), .S(n10198), .Z(n7604) );
  INV_X1 U9322 ( .A(n7598), .ZN(n9169) );
  OAI22_X1 U9323 ( .A1(n9260), .A2(n7600), .B1(n9241), .B2(n7599), .ZN(n7601)
         );
  AOI21_X1 U9324 ( .B1(n7602), .B2(n9169), .A(n7601), .ZN(n7603) );
  OAI211_X1 U9325 ( .C1(n7605), .C2(n9274), .A(n7604), .B(n7603), .ZN(P2_U3292) );
  INV_X1 U9326 ( .A(n7606), .ZN(n7637) );
  AOI22_X1 U9327 ( .A1(n8987), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n9376), .ZN(n7607) );
  OAI21_X1 U9328 ( .B1(n7637), .B2(n4451), .A(n7607), .ZN(P2_U3340) );
  INV_X1 U9329 ( .A(n7609), .ZN(n7610) );
  AOI21_X1 U9330 ( .B1(n7611), .B2(n7608), .A(n7610), .ZN(n7617) );
  OAI22_X1 U9331 ( .A1(n9455), .A2(n7612), .B1(n9472), .B2(n10035), .ZN(n7613)
         );
  AOI211_X1 U9332 ( .C1(n8126), .C2(n10023), .A(n7614), .B(n7613), .ZN(n7616)
         );
  NAND2_X1 U9333 ( .A1(n10150), .A2(n9459), .ZN(n7615) );
  OAI211_X1 U9334 ( .C1(n7617), .C2(n9461), .A(n7616), .B(n7615), .ZN(P1_U3229) );
  NOR2_X1 U9335 ( .A1(n9241), .A2(n7618), .ZN(n7622) );
  OAI22_X1 U9336 ( .A1(n7620), .A2(n9274), .B1(n7619), .B2(n9260), .ZN(n7621)
         );
  AOI211_X1 U9337 ( .C1(n9272), .C2(n7623), .A(n7622), .B(n7621), .ZN(n7627)
         );
  MUX2_X1 U9338 ( .A(n7625), .B(n7624), .S(n9244), .Z(n7626) );
  NAND2_X1 U9339 ( .A1(n7627), .A2(n7626), .ZN(P2_U3295) );
  OAI22_X1 U9340 ( .A1(n8887), .A2(n7677), .B1(n7631), .B2(n8885), .ZN(n7634)
         );
  AOI22_X1 U9341 ( .A1(n8890), .A2(n8671), .B1(P2_REG3_REG_7__SCAN_IN), .B2(
        P2_U3152), .ZN(n7632) );
  OAI21_X1 U9342 ( .B1(n8641), .B2(n8875), .A(n7632), .ZN(n7633) );
  OR3_X1 U9343 ( .A1(n7635), .A2(n7634), .A3(n7633), .ZN(P2_U3215) );
  INV_X1 U9344 ( .A(n9548), .ZN(n7636) );
  OAI222_X1 U9345 ( .A1(n9831), .A2(n7638), .B1(n9835), .B2(n7637), .C1(
        P1_U3084), .C2(n7636), .ZN(P1_U3335) );
  NAND2_X1 U9346 ( .A1(n8886), .A2(n10239), .ZN(n7640) );
  NAND2_X1 U9347 ( .A1(n7677), .A2(n7672), .ZN(n8678) );
  INV_X1 U9348 ( .A(n7672), .ZN(n10247) );
  NAND2_X1 U9349 ( .A1(n8907), .A2(n10247), .ZN(n8679) );
  INV_X1 U9350 ( .A(n8675), .ZN(n7642) );
  NAND2_X1 U9351 ( .A1(n7643), .A2(n8675), .ZN(n7644) );
  NAND2_X1 U9352 ( .A1(n7674), .A2(n7644), .ZN(n10246) );
  OR2_X1 U9353 ( .A1(n10246), .A2(n8170), .ZN(n7653) );
  NAND2_X1 U9354 ( .A1(n8908), .A2(n10239), .ZN(n7645) );
  NAND2_X1 U9355 ( .A1(n7647), .A2(n7642), .ZN(n7648) );
  NAND2_X1 U9356 ( .A1(n7676), .A2(n7648), .ZN(n7651) );
  NAND2_X1 U9357 ( .A1(n8908), .A2(n9264), .ZN(n7649) );
  OAI21_X1 U9358 ( .B1(n7754), .B2(n9231), .A(n7649), .ZN(n7650) );
  AOI21_X1 U9359 ( .B1(n7651), .B2(n9269), .A(n7650), .ZN(n7652) );
  NAND2_X1 U9360 ( .A1(n7653), .A2(n7652), .ZN(n10251) );
  NAND2_X1 U9361 ( .A1(n10251), .A2(n9238), .ZN(n7662) );
  OAI22_X1 U9362 ( .A1(n9244), .A2(n7655), .B1(n7654), .B2(n9241), .ZN(n7660)
         );
  NAND2_X1 U9363 ( .A1(n7656), .A2(n10239), .ZN(n7657) );
  OR2_X1 U9364 ( .A1(n7657), .A2(n7672), .ZN(n7683) );
  NAND2_X1 U9365 ( .A1(n7657), .A2(n7672), .ZN(n7658) );
  NAND2_X1 U9366 ( .A1(n7683), .A2(n7658), .ZN(n10248) );
  NOR2_X1 U9367 ( .A1(n10248), .A2(n9218), .ZN(n7659) );
  AOI211_X1 U9368 ( .C1(n9246), .C2(n7672), .A(n7660), .B(n7659), .ZN(n7661)
         );
  OAI211_X1 U9369 ( .C1(n10246), .C2(n9250), .A(n7662), .B(n7661), .ZN(
        P2_U3288) );
  NOR2_X1 U9370 ( .A1(n4937), .A2(n7664), .ZN(n7665) );
  XNOR2_X1 U9371 ( .A(n7666), .B(n7665), .ZN(n7671) );
  AOI22_X1 U9372 ( .A1(n8097), .A2(n8905), .B1(n8894), .B2(n8907), .ZN(n7668)
         );
  OAI211_X1 U9373 ( .C1(n7685), .C2(n8885), .A(n7668), .B(n7667), .ZN(n7669)
         );
  AOI21_X1 U9374 ( .B1(n7688), .B2(n8890), .A(n7669), .ZN(n7670) );
  OAI21_X1 U9375 ( .B1(n7671), .B2(n8868), .A(n7670), .ZN(P2_U3233) );
  NAND2_X1 U9376 ( .A1(n8907), .A2(n7672), .ZN(n7673) );
  NAND2_X1 U9377 ( .A1(n7754), .A2(n7688), .ZN(n8683) );
  INV_X1 U9378 ( .A(n7688), .ZN(n10253) );
  INV_X1 U9379 ( .A(n7754), .ZN(n8906) );
  NAND2_X1 U9380 ( .A1(n10253), .A2(n8906), .ZN(n8691) );
  NAND2_X1 U9381 ( .A1(n7853), .A2(n7851), .ZN(n7675) );
  NAND2_X1 U9382 ( .A1(n7755), .A2(n7675), .ZN(n10256) );
  INV_X1 U9383 ( .A(n7851), .ZN(n8621) );
  XNOR2_X1 U9384 ( .A(n7760), .B(n8621), .ZN(n7680) );
  OAI22_X1 U9385 ( .A1(n7677), .A2(n9233), .B1(n7861), .B2(n9231), .ZN(n7678)
         );
  INV_X1 U9386 ( .A(n7678), .ZN(n7679) );
  OAI21_X1 U9387 ( .B1(n7680), .B2(n9228), .A(n7679), .ZN(n7681) );
  AOI21_X1 U9388 ( .B1(n10256), .B2(n7682), .A(n7681), .ZN(n10258) );
  AND2_X1 U9389 ( .A1(n7683), .A2(n7688), .ZN(n7684) );
  OR2_X1 U9390 ( .A1(n7684), .A2(n7767), .ZN(n10254) );
  OAI22_X1 U9391 ( .A1(n9238), .A2(n7686), .B1(n7685), .B2(n9241), .ZN(n7687)
         );
  AOI21_X1 U9392 ( .B1(n9246), .B2(n7688), .A(n7687), .ZN(n7689) );
  OAI21_X1 U9393 ( .B1(n10254), .B2(n9218), .A(n7689), .ZN(n7690) );
  AOI21_X1 U9394 ( .B1(n10256), .B2(n7691), .A(n7690), .ZN(n7692) );
  OAI21_X1 U9395 ( .B1(n10258), .B2(n10198), .A(n7692), .ZN(P2_U3287) );
  INV_X1 U9396 ( .A(n8261), .ZN(n8383) );
  XNOR2_X1 U9397 ( .A(n7693), .B(n8383), .ZN(n7694) );
  AOI222_X1 U9398 ( .A1(n10050), .A2(n7694), .B1(n9492), .B2(n10045), .C1(
        n9491), .C2(n10046), .ZN(n9868) );
  OAI22_X1 U9399 ( .A1(n10031), .A2(n7695), .B1(n7710), .B2(n10036), .ZN(n7698) );
  INV_X1 U9400 ( .A(n10016), .ZN(n7696) );
  INV_X1 U9401 ( .A(n7699), .ZN(n9869) );
  OAI211_X1 U9402 ( .C1(n7696), .C2(n9869), .A(n10124), .B(n7790), .ZN(n9867)
         );
  NOR2_X1 U9403 ( .A1(n9867), .A2(n8057), .ZN(n7697) );
  AOI211_X1 U9404 ( .C1(n9739), .C2(n7699), .A(n7698), .B(n7697), .ZN(n7702)
         );
  XNOR2_X1 U9405 ( .A(n7700), .B(n8261), .ZN(n9871) );
  NAND2_X1 U9406 ( .A1(n9871), .A2(n9611), .ZN(n7701) );
  OAI211_X1 U9407 ( .C1(n9868), .C2(n9738), .A(n7702), .B(n7701), .ZN(P1_U3281) );
  INV_X1 U9408 ( .A(n7703), .ZN(n7705) );
  OAI222_X1 U9409 ( .A1(n9831), .A2(n7704), .B1(n9835), .B2(n7705), .C1(
        P1_U3084), .C2(n9644), .ZN(P1_U3334) );
  OAI222_X1 U9410 ( .A1(n9379), .A2(n7706), .B1(n4451), .B2(n7705), .C1(
        P2_U3152), .C2(n7032), .ZN(P2_U3339) );
  XNOR2_X1 U9411 ( .A(n7708), .B(n7707), .ZN(n7709) );
  NAND2_X1 U9412 ( .A1(n7709), .A2(n9467), .ZN(n7715) );
  OAI22_X1 U9413 ( .A1(n9455), .A2(n7711), .B1(n9472), .B2(n7710), .ZN(n7712)
         );
  AOI211_X1 U9414 ( .C1(n8126), .C2(n9491), .A(n7713), .B(n7712), .ZN(n7714)
         );
  OAI211_X1 U9415 ( .C1(n9869), .C2(n9478), .A(n7715), .B(n7714), .ZN(P1_U3215) );
  XNOR2_X1 U9416 ( .A(n7717), .B(n7716), .ZN(n7721) );
  AOI22_X1 U9417 ( .A1(n8097), .A2(n8904), .B1(n8894), .B2(n8906), .ZN(n7718)
         );
  NAND2_X1 U9418 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n8939) );
  OAI211_X1 U9419 ( .C1(n7765), .C2(n8885), .A(n7718), .B(n8939), .ZN(n7719)
         );
  AOI21_X1 U9420 ( .B1(n7849), .B2(n8890), .A(n7719), .ZN(n7720) );
  OAI21_X1 U9421 ( .B1(n7721), .B2(n8868), .A(n7720), .ZN(P2_U3219) );
  INV_X1 U9422 ( .A(n7796), .ZN(n9928) );
  AOI21_X1 U9423 ( .B1(n7723), .B2(n7722), .A(n9461), .ZN(n7726) );
  NAND2_X1 U9424 ( .A1(n7726), .A2(n7725), .ZN(n7730) );
  OAI22_X1 U9425 ( .A1(n9455), .A2(n7787), .B1(n9472), .B2(n7793), .ZN(n7727)
         );
  AOI211_X1 U9426 ( .C1(n8126), .C2(n9490), .A(n7728), .B(n7727), .ZN(n7729)
         );
  OAI211_X1 U9427 ( .C1(n9928), .C2(n9478), .A(n7730), .B(n7729), .ZN(P1_U3234) );
  INV_X1 U9428 ( .A(n7731), .ZN(n7733) );
  OAI222_X1 U9429 ( .A1(n9835), .A2(n7733), .B1(n8549), .B2(P1_U3084), .C1(
        n7732), .C2(n9831), .ZN(P1_U3333) );
  OAI222_X1 U9430 ( .A1(n9379), .A2(n7734), .B1(n4451), .B2(n7733), .C1(n4462), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  MUX2_X1 U9431 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7735), .S(n8000), .Z(n7738)
         );
  OAI21_X1 U9432 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n7741), .A(n7736), .ZN(
        n7737) );
  NAND2_X1 U9433 ( .A1(n7737), .A2(n7738), .ZN(n7999) );
  OAI21_X1 U9434 ( .B1(n7738), .B2(n7737), .A(n7999), .ZN(n7745) );
  NAND2_X1 U9435 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n8131) );
  NAND2_X1 U9436 ( .A1(n10013), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n7739) );
  OAI211_X1 U9437 ( .C1(n9525), .C2(n7994), .A(n8131), .B(n7739), .ZN(n7744)
         );
  NOR2_X1 U9438 ( .A1(n6047), .A2(n7742), .ZN(n7996) );
  AOI211_X1 U9439 ( .C1(n7742), .C2(n6047), .A(n7996), .B(n10003), .ZN(n7743)
         );
  AOI211_X1 U9440 ( .C1(n10010), .C2(n7745), .A(n7744), .B(n7743), .ZN(n7746)
         );
  INV_X1 U9441 ( .A(n7746), .ZN(P1_U3255) );
  XNOR2_X1 U9442 ( .A(n7748), .B(n7747), .ZN(n7753) );
  OAI22_X1 U9443 ( .A1(n8885), .A2(n7863), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7749), .ZN(n7751) );
  OAI22_X1 U9444 ( .A1(n7980), .A2(n8887), .B1(n8875), .B2(n7861), .ZN(n7750)
         );
  AOI211_X1 U9445 ( .C1(n7919), .C2(n8890), .A(n7751), .B(n7750), .ZN(n7752)
         );
  OAI21_X1 U9446 ( .B1(n7753), .B2(n8868), .A(n7752), .ZN(P2_U3238) );
  NAND2_X1 U9447 ( .A1(n7754), .A2(n10253), .ZN(n7854) );
  NAND2_X1 U9448 ( .A1(n7755), .A2(n7854), .ZN(n7756) );
  OR2_X1 U9449 ( .A1(n7861), .A2(n7849), .ZN(n8689) );
  NAND2_X1 U9450 ( .A1(n7849), .A2(n7861), .ZN(n8688) );
  OR2_X1 U9451 ( .A1(n7756), .A2(n7761), .ZN(n7758) );
  NAND2_X1 U9452 ( .A1(n7756), .A2(n7761), .ZN(n7757) );
  NAND2_X1 U9453 ( .A1(n7758), .A2(n7757), .ZN(n10259) );
  AOI22_X1 U9454 ( .A1(n9264), .A2(n8906), .B1(n8904), .B2(n9266), .ZN(n7764)
         );
  INV_X1 U9455 ( .A(n8683), .ZN(n7759) );
  INV_X1 U9456 ( .A(n7761), .ZN(n8622) );
  NAND2_X1 U9457 ( .A1(n7762), .A2(n7761), .ZN(n7859) );
  OAI211_X1 U9458 ( .C1(n7762), .C2(n7761), .A(n7859), .B(n9269), .ZN(n7763)
         );
  OAI211_X1 U9459 ( .C1(n10259), .C2(n8170), .A(n7764), .B(n7763), .ZN(n10262)
         );
  NAND2_X1 U9460 ( .A1(n10262), .A2(n9238), .ZN(n7772) );
  OAI22_X1 U9461 ( .A1(n9244), .A2(n7766), .B1(n7765), .B2(n9241), .ZN(n7770)
         );
  INV_X1 U9462 ( .A(n7849), .ZN(n10260) );
  NOR2_X1 U9463 ( .A1(n7767), .A2(n10260), .ZN(n7768) );
  OR2_X1 U9464 ( .A1(n7862), .A2(n7768), .ZN(n10261) );
  NOR2_X1 U9465 ( .A1(n10261), .A2(n9218), .ZN(n7769) );
  AOI211_X1 U9466 ( .C1(n9246), .C2(n7849), .A(n7770), .B(n7769), .ZN(n7771)
         );
  OAI211_X1 U9467 ( .C1(n10259), .C2(n9250), .A(n7772), .B(n7771), .ZN(
        P2_U3286) );
  XNOR2_X1 U9468 ( .A(n7774), .B(n7773), .ZN(n7775) );
  XNOR2_X1 U9469 ( .A(n7776), .B(n7775), .ZN(n7781) );
  OAI21_X1 U9470 ( .B1(n9473), .B2(n7887), .A(n7777), .ZN(n7779) );
  OAI22_X1 U9471 ( .A1(n9455), .A2(n7886), .B1(n9472), .B2(n7891), .ZN(n7778)
         );
  AOI211_X1 U9472 ( .C1(n8028), .C2(n9459), .A(n7779), .B(n7778), .ZN(n7780)
         );
  OAI21_X1 U9473 ( .B1(n7781), .B2(n9461), .A(n7780), .ZN(P1_U3222) );
  INV_X1 U9474 ( .A(n7782), .ZN(n7801) );
  OAI222_X1 U9475 ( .A1(n9835), .A2(n7801), .B1(n8289), .B2(P1_U3084), .C1(
        n7783), .C2(n9831), .ZN(P1_U3332) );
  XNOR2_X1 U9476 ( .A(n7796), .B(n9491), .ZN(n8388) );
  XNOR2_X1 U9477 ( .A(n7784), .B(n8388), .ZN(n9932) );
  INV_X1 U9478 ( .A(n9932), .ZN(n7800) );
  INV_X1 U9479 ( .A(n8388), .ZN(n8264) );
  INV_X1 U9480 ( .A(n7785), .ZN(n7786) );
  NOR2_X1 U9481 ( .A1(n7786), .A2(n8264), .ZN(n7883) );
  AOI211_X1 U9482 ( .C1(n8264), .C2(n7786), .A(n6466), .B(n7883), .ZN(n7789)
         );
  OAI22_X1 U9483 ( .A1(n7912), .A2(n9716), .B1(n7787), .B2(n6463), .ZN(n7788)
         );
  OR2_X1 U9484 ( .A1(n7789), .A2(n7788), .ZN(n9930) );
  INV_X1 U9485 ( .A(n7790), .ZN(n7792) );
  INV_X1 U9486 ( .A(n7791), .ZN(n7889) );
  OAI21_X1 U9487 ( .B1(n9928), .B2(n7792), .A(n7889), .ZN(n9929) );
  OAI22_X1 U9488 ( .A1(n10057), .A2(n7794), .B1(n7793), .B2(n10036), .ZN(n7795) );
  AOI21_X1 U9489 ( .B1(n7796), .B2(n9739), .A(n7795), .ZN(n7797) );
  OAI21_X1 U9490 ( .B1(n9929), .B2(n10019), .A(n7797), .ZN(n7798) );
  AOI21_X1 U9491 ( .B1(n9930), .B2(n10031), .A(n7798), .ZN(n7799) );
  OAI21_X1 U9492 ( .B1(n9746), .B2(n7800), .A(n7799), .ZN(P1_U3280) );
  OAI222_X1 U9493 ( .A1(n9379), .A2(n7802), .B1(n4451), .B2(n7801), .C1(n8598), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  INV_X1 U9494 ( .A(n7804), .ZN(n8269) );
  XNOR2_X1 U9495 ( .A(n7803), .B(n8269), .ZN(n9927) );
  INV_X1 U9496 ( .A(n9927), .ZN(n7817) );
  INV_X1 U9497 ( .A(n7805), .ZN(n7809) );
  INV_X1 U9498 ( .A(n7806), .ZN(n8396) );
  AOI21_X1 U9499 ( .B1(n7807), .B2(n8396), .A(n8269), .ZN(n7808) );
  NOR2_X1 U9500 ( .A1(n7809), .A2(n7808), .ZN(n7810) );
  OAI222_X1 U9501 ( .A1(n9716), .A2(n8300), .B1(n6463), .B2(n7912), .C1(n6466), 
        .C2(n7810), .ZN(n9925) );
  INV_X1 U9502 ( .A(n7811), .ZN(n7888) );
  INV_X1 U9503 ( .A(n7915), .ZN(n9923) );
  OAI21_X1 U9504 ( .B1(n7888), .B2(n9923), .A(n7872), .ZN(n9924) );
  OAI22_X1 U9505 ( .A1(n10057), .A2(n7812), .B1(n7911), .B2(n10036), .ZN(n7813) );
  AOI21_X1 U9506 ( .B1(n7915), .B2(n9739), .A(n7813), .ZN(n7814) );
  OAI21_X1 U9507 ( .B1(n9924), .B2(n10019), .A(n7814), .ZN(n7815) );
  AOI21_X1 U9508 ( .B1(n9925), .B2(n10031), .A(n7815), .ZN(n7816) );
  OAI21_X1 U9509 ( .B1(n7817), .B2(n9746), .A(n7816), .ZN(P1_U3278) );
  INV_X1 U9510 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10329) );
  NOR2_X1 U9511 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7818) );
  AOI21_X1 U9512 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7818), .ZN(n10300) );
  NOR2_X1 U9513 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .ZN(n7819) );
  AOI21_X1 U9514 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n7819), .ZN(n10303) );
  NOR2_X1 U9515 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7820) );
  AOI21_X1 U9516 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7820), .ZN(n10306) );
  NOR2_X1 U9517 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7821) );
  AOI21_X1 U9518 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7821), .ZN(n10309) );
  NOR2_X1 U9519 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .ZN(n7822) );
  AOI21_X1 U9520 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n7822), .ZN(n10312) );
  NOR2_X1 U9521 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7829) );
  XNOR2_X1 U9522 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10341) );
  NAND2_X1 U9523 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7827) );
  XOR2_X1 U9524 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10339) );
  NAND2_X1 U9525 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7825) );
  XOR2_X1 U9526 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10337) );
  AOI21_X1 U9527 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10294) );
  INV_X1 U9528 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7823) );
  NAND3_X1 U9529 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10296) );
  OAI21_X1 U9530 ( .B1(n10294), .B2(n7823), .A(n10296), .ZN(n10336) );
  NAND2_X1 U9531 ( .A1(n10337), .A2(n10336), .ZN(n7824) );
  NAND2_X1 U9532 ( .A1(n7825), .A2(n7824), .ZN(n10338) );
  NAND2_X1 U9533 ( .A1(n10339), .A2(n10338), .ZN(n7826) );
  NAND2_X1 U9534 ( .A1(n7827), .A2(n7826), .ZN(n10340) );
  NOR2_X1 U9535 ( .A1(n10341), .A2(n10340), .ZN(n7828) );
  NOR2_X1 U9536 ( .A1(n7829), .A2(n7828), .ZN(n7830) );
  NOR2_X1 U9537 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7830), .ZN(n10323) );
  AND2_X1 U9538 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7830), .ZN(n10324) );
  NOR2_X1 U9539 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10324), .ZN(n7831) );
  NAND2_X1 U9540 ( .A1(n7832), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7834) );
  XOR2_X1 U9541 ( .A(n7832), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10322) );
  NAND2_X1 U9542 ( .A1(n10322), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7833) );
  NAND2_X1 U9543 ( .A1(n7834), .A2(n7833), .ZN(n7835) );
  NAND2_X1 U9544 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7835), .ZN(n7837) );
  XOR2_X1 U9545 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7835), .Z(n10335) );
  NAND2_X1 U9546 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10335), .ZN(n7836) );
  NAND2_X1 U9547 ( .A1(n7837), .A2(n7836), .ZN(n7838) );
  NAND2_X1 U9548 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7838), .ZN(n7840) );
  XOR2_X1 U9549 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7838), .Z(n10334) );
  NAND2_X1 U9550 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10334), .ZN(n7839) );
  NAND2_X1 U9551 ( .A1(n7840), .A2(n7839), .ZN(n7841) );
  AND2_X1 U9552 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7841), .ZN(n7842) );
  XNOR2_X1 U9553 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7841), .ZN(n10332) );
  NAND2_X1 U9554 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7843) );
  OAI21_X1 U9555 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n7843), .ZN(n10320) );
  NAND2_X1 U9556 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7844) );
  OAI21_X1 U9557 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7844), .ZN(n10317) );
  AOI21_X1 U9558 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10316), .ZN(n10315) );
  NOR2_X1 U9559 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7845) );
  AOI21_X1 U9560 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7845), .ZN(n10314) );
  NAND2_X1 U9561 ( .A1(n10315), .A2(n10314), .ZN(n10313) );
  OAI21_X1 U9562 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10313), .ZN(n10311) );
  NAND2_X1 U9563 ( .A1(n10312), .A2(n10311), .ZN(n10310) );
  OAI21_X1 U9564 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10310), .ZN(n10308) );
  NAND2_X1 U9565 ( .A1(n10309), .A2(n10308), .ZN(n10307) );
  OAI21_X1 U9566 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10307), .ZN(n10305) );
  NAND2_X1 U9567 ( .A1(n10306), .A2(n10305), .ZN(n10304) );
  OAI21_X1 U9568 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10304), .ZN(n10302) );
  NAND2_X1 U9569 ( .A1(n10303), .A2(n10302), .ZN(n10301) );
  OAI21_X1 U9570 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10301), .ZN(n10299) );
  NAND2_X1 U9571 ( .A1(n10300), .A2(n10299), .ZN(n10298) );
  OAI21_X1 U9572 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10298), .ZN(n10328) );
  NOR2_X1 U9573 ( .A1(n10329), .A2(n10328), .ZN(n7846) );
  NAND2_X1 U9574 ( .A1(n10329), .A2(n10328), .ZN(n10327) );
  OAI21_X1 U9575 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7846), .A(n10327), .ZN(
        n7848) );
  XNOR2_X1 U9576 ( .A(n8998), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7847) );
  XNOR2_X1 U9577 ( .A(n7848), .B(n7847), .ZN(ADD_1071_U4) );
  NAND2_X1 U9578 ( .A1(n7849), .A2(n8905), .ZN(n7856) );
  INV_X1 U9579 ( .A(n7856), .ZN(n7850) );
  OR2_X1 U9580 ( .A1(n7851), .A2(n7850), .ZN(n7852) );
  NAND2_X1 U9581 ( .A1(n8622), .A2(n7854), .ZN(n7855) );
  AND2_X1 U9582 ( .A1(n7856), .A2(n7855), .ZN(n7857) );
  OR2_X1 U9583 ( .A1(n7919), .A2(n7927), .ZN(n8690) );
  NAND2_X1 U9584 ( .A1(n7919), .A2(n7927), .ZN(n8700) );
  NAND2_X1 U9585 ( .A1(n8690), .A2(n8700), .ZN(n8623) );
  OAI21_X1 U9586 ( .B1(n7858), .B2(n8623), .A(n7921), .ZN(n10266) );
  XOR2_X1 U9587 ( .A(n7924), .B(n8623), .Z(n7860) );
  OAI222_X1 U9588 ( .A1(n9231), .A2(n7980), .B1(n9233), .B2(n7861), .C1(n9228), 
        .C2(n7860), .ZN(n10269) );
  INV_X1 U9589 ( .A(n7919), .ZN(n10267) );
  OAI21_X1 U9590 ( .B1(n7862), .B2(n10267), .A(n7928), .ZN(n10268) );
  OAI22_X1 U9591 ( .A1(n9244), .A2(n7864), .B1(n7863), .B2(n9241), .ZN(n7865)
         );
  AOI21_X1 U9592 ( .B1(n9246), .B2(n7919), .A(n7865), .ZN(n7866) );
  OAI21_X1 U9593 ( .B1(n10268), .B2(n9218), .A(n7866), .ZN(n7867) );
  AOI21_X1 U9594 ( .B1(n10269), .B2(n9238), .A(n7867), .ZN(n7868) );
  OAI21_X1 U9595 ( .B1(n9274), .B2(n10266), .A(n7868), .ZN(P2_U3285) );
  XNOR2_X1 U9596 ( .A(n7869), .B(n8266), .ZN(n9810) );
  XNOR2_X1 U9597 ( .A(n7870), .B(n8266), .ZN(n7871) );
  OAI222_X1 U9598 ( .A1(n9716), .A2(n8133), .B1(n6463), .B2(n7887), .C1(n6466), 
        .C2(n7871), .ZN(n9806) );
  AOI211_X1 U9599 ( .C1(n9808), .C2(n7872), .A(n10154), .B(n8042), .ZN(n9807)
         );
  INV_X1 U9600 ( .A(n8057), .ZN(n7895) );
  NAND2_X1 U9601 ( .A1(n9807), .A2(n7895), .ZN(n7874) );
  AOI22_X1 U9602 ( .A1(n9738), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8129), .B2(
        n10041), .ZN(n7873) );
  OAI211_X1 U9603 ( .C1(n4707), .C2(n9724), .A(n7874), .B(n7873), .ZN(n7875)
         );
  AOI21_X1 U9604 ( .B1(n9806), .B2(n10031), .A(n7875), .ZN(n7876) );
  OAI21_X1 U9605 ( .B1(n9810), .B2(n9746), .A(n7876), .ZN(P1_U3277) );
  INV_X1 U9606 ( .A(n7877), .ZN(n7879) );
  OAI222_X1 U9607 ( .A1(n9831), .A2(n7878), .B1(n9835), .B2(n7879), .C1(
        P1_U3084), .C2(n8556), .ZN(P1_U3331) );
  OAI222_X1 U9608 ( .A1(n9379), .A2(n7880), .B1(n4451), .B2(n7879), .C1(
        P2_U3152), .C2(n8635), .ZN(P2_U3336) );
  XNOR2_X1 U9609 ( .A(n7881), .B(n8265), .ZN(n8030) );
  NOR2_X1 U9610 ( .A1(n7883), .A2(n7882), .ZN(n7884) );
  XNOR2_X1 U9611 ( .A(n7884), .B(n8265), .ZN(n7885) );
  OAI222_X1 U9612 ( .A1(n9716), .A2(n7887), .B1(n6463), .B2(n7886), .C1(n6466), 
        .C2(n7885), .ZN(n8026) );
  NAND2_X1 U9613 ( .A1(n8026), .A2(n10057), .ZN(n7897) );
  AOI211_X1 U9614 ( .C1(n8028), .C2(n7889), .A(n10154), .B(n7888), .ZN(n8027)
         );
  NOR2_X1 U9615 ( .A1(n7890), .A2(n9724), .ZN(n7894) );
  OAI22_X1 U9616 ( .A1(n10057), .A2(n7892), .B1(n7891), .B2(n10036), .ZN(n7893) );
  AOI211_X1 U9617 ( .C1(n8027), .C2(n7895), .A(n7894), .B(n7893), .ZN(n7896)
         );
  OAI211_X1 U9618 ( .C1(n8030), .C2(n9746), .A(n7897), .B(n7896), .ZN(P1_U3279) );
  NAND2_X1 U9619 ( .A1(n7899), .A2(n7898), .ZN(n7901) );
  XOR2_X1 U9620 ( .A(n7901), .B(n7900), .Z(n7906) );
  AOI22_X1 U9621 ( .A1(n8097), .A2(n8902), .B1(n8894), .B2(n8904), .ZN(n7903)
         );
  OAI211_X1 U9622 ( .C1(n7930), .C2(n8885), .A(n7903), .B(n7902), .ZN(n7904)
         );
  AOI21_X1 U9623 ( .B1(n7958), .B2(n8890), .A(n7904), .ZN(n7905) );
  OAI21_X1 U9624 ( .B1(n7906), .B2(n8868), .A(n7905), .ZN(P2_U3226) );
  NAND2_X1 U9625 ( .A1(n7908), .A2(n7907), .ZN(n7909) );
  XNOR2_X1 U9626 ( .A(n7910), .B(n7909), .ZN(n7918) );
  OAI22_X1 U9627 ( .A1(n9455), .A2(n7912), .B1(n9472), .B2(n7911), .ZN(n7913)
         );
  AOI211_X1 U9628 ( .C1(n8126), .C2(n9488), .A(n7914), .B(n7913), .ZN(n7917)
         );
  NAND2_X1 U9629 ( .A1(n7915), .A2(n9459), .ZN(n7916) );
  OAI211_X1 U9630 ( .C1(n7918), .C2(n9461), .A(n7917), .B(n7916), .ZN(P1_U3232) );
  NAND2_X1 U9631 ( .A1(n7919), .A2(n8904), .ZN(n7920) );
  OR2_X1 U9632 ( .A1(n7958), .A2(n7980), .ZN(n8702) );
  NAND2_X1 U9633 ( .A1(n7958), .A2(n7980), .ZN(n8701) );
  OAI21_X1 U9634 ( .B1(n7923), .B2(n7922), .A(n7961), .ZN(n10277) );
  INV_X1 U9635 ( .A(n10277), .ZN(n7936) );
  INV_X1 U9636 ( .A(n8902), .ZN(n8093) );
  NAND2_X1 U9637 ( .A1(n7965), .A2(n8690), .ZN(n7925) );
  XNOR2_X1 U9638 ( .A(n7925), .B(n8626), .ZN(n7926) );
  OAI222_X1 U9639 ( .A1(n9233), .A2(n7927), .B1(n9231), .B2(n8093), .C1(n9228), 
        .C2(n7926), .ZN(n10275) );
  INV_X1 U9640 ( .A(n7928), .ZN(n7929) );
  OAI21_X1 U9641 ( .B1(n7929), .B2(n4614), .A(n7970), .ZN(n10274) );
  OAI22_X1 U9642 ( .A1(n9244), .A2(n7931), .B1(n7930), .B2(n9241), .ZN(n7932)
         );
  AOI21_X1 U9643 ( .B1(n9246), .B2(n7958), .A(n7932), .ZN(n7933) );
  OAI21_X1 U9644 ( .B1(n10274), .B2(n9218), .A(n7933), .ZN(n7934) );
  AOI21_X1 U9645 ( .B1(n10275), .B2(n9238), .A(n7934), .ZN(n7935) );
  OAI21_X1 U9646 ( .B1(n7936), .B2(n9274), .A(n7935), .ZN(P2_U3284) );
  INV_X1 U9647 ( .A(n8971), .ZN(n7943) );
  XNOR2_X1 U9648 ( .A(n8971), .B(n9243), .ZN(n8967) );
  NAND2_X1 U9649 ( .A1(n8961), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7942) );
  INV_X1 U9650 ( .A(n7942), .ZN(n7937) );
  AOI21_X1 U9651 ( .B1(n8175), .B2(n7945), .A(n7937), .ZN(n8953) );
  NOR2_X1 U9652 ( .A1(n7939), .A2(n7938), .ZN(n7941) );
  NOR2_X1 U9653 ( .A1(n7941), .A2(n7940), .ZN(n8954) );
  NAND2_X1 U9654 ( .A1(n8953), .A2(n8954), .ZN(n8952) );
  NAND2_X1 U9655 ( .A1(n7942), .A2(n8952), .ZN(n8968) );
  NAND2_X1 U9656 ( .A1(n8967), .A2(n8968), .ZN(n8966) );
  OAI21_X1 U9657 ( .B1(n7943), .B2(n9243), .A(n8966), .ZN(n8982) );
  XNOR2_X1 U9658 ( .A(n8982), .B(n8987), .ZN(n8980) );
  XOR2_X1 U9659 ( .A(P2_REG2_REG_18__SCAN_IN), .B(n8980), .Z(n7957) );
  NOR2_X1 U9660 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8873), .ZN(n7954) );
  XNOR2_X1 U9661 ( .A(n8987), .B(n7944), .ZN(n7951) );
  XNOR2_X1 U9662 ( .A(n8971), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8974) );
  XNOR2_X1 U9663 ( .A(n7945), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8958) );
  NOR2_X1 U9664 ( .A1(n7947), .A2(n7946), .ZN(n7949) );
  NOR2_X1 U9665 ( .A1(n7949), .A2(n7948), .ZN(n8959) );
  NAND2_X1 U9666 ( .A1(n8958), .A2(n8959), .ZN(n8957) );
  OAI21_X1 U9667 ( .B1(n8961), .B2(P2_REG1_REG_16__SCAN_IN), .A(n8957), .ZN(
        n8973) );
  NOR2_X1 U9668 ( .A1(n8974), .A2(n8973), .ZN(n8972) );
  AOI21_X1 U9669 ( .B1(n8971), .B2(P2_REG1_REG_17__SCAN_IN), .A(n8972), .ZN(
        n7950) );
  NAND2_X1 U9670 ( .A1(n7951), .A2(n7950), .ZN(n8986) );
  OAI21_X1 U9671 ( .B1(n7951), .B2(n7950), .A(n8986), .ZN(n7952) );
  AND2_X1 U9672 ( .A1(n10174), .A2(n7952), .ZN(n7953) );
  AOI211_X1 U9673 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n10176), .A(n7954), .B(
        n7953), .ZN(n7956) );
  NAND2_X1 U9674 ( .A1(n9860), .A2(n8987), .ZN(n7955) );
  OAI211_X1 U9675 ( .C1(n7957), .C2(n8990), .A(n7956), .B(n7955), .ZN(P2_U3263) );
  OR2_X1 U9676 ( .A1(n7958), .A2(n8903), .ZN(n7962) );
  XNOR2_X1 U9677 ( .A(n8704), .B(n8902), .ZN(n8709) );
  INV_X1 U9678 ( .A(n8709), .ZN(n7959) );
  AND2_X1 U9679 ( .A1(n7962), .A2(n7959), .ZN(n7960) );
  NAND2_X1 U9680 ( .A1(n7961), .A2(n7962), .ZN(n7963) );
  NAND2_X1 U9681 ( .A1(n7963), .A2(n8709), .ZN(n7964) );
  NAND2_X1 U9682 ( .A1(n8006), .A2(n7964), .ZN(n9890) );
  AND2_X1 U9683 ( .A1(n8702), .A2(n8690), .ZN(n8698) );
  XNOR2_X1 U9684 ( .A(n8008), .B(n8709), .ZN(n7967) );
  INV_X1 U9685 ( .A(n9265), .ZN(n8710) );
  OAI22_X1 U9686 ( .A1(n8710), .A2(n9231), .B1(n7980), .B2(n9233), .ZN(n7966)
         );
  AOI21_X1 U9687 ( .B1(n7967), .B2(n9269), .A(n7966), .ZN(n7968) );
  OAI21_X1 U9688 ( .B1(n9890), .B2(n8170), .A(n7968), .ZN(n9893) );
  NAND2_X1 U9689 ( .A1(n9893), .A2(n9238), .ZN(n7975) );
  OAI22_X1 U9690 ( .A1(n9244), .A2(n7969), .B1(n7979), .B2(n9241), .ZN(n7973)
         );
  NAND2_X1 U9691 ( .A1(n7970), .A2(n8704), .ZN(n7971) );
  NAND2_X1 U9692 ( .A1(n8172), .A2(n7971), .ZN(n9892) );
  NOR2_X1 U9693 ( .A1(n9892), .A2(n9218), .ZN(n7972) );
  AOI211_X1 U9694 ( .C1(n9246), .C2(n8704), .A(n7973), .B(n7972), .ZN(n7974)
         );
  OAI211_X1 U9695 ( .C1(n9890), .C2(n9250), .A(n7975), .B(n7974), .ZN(P2_U3283) );
  OAI211_X1 U9696 ( .C1(n7978), .C2(n7977), .A(n7976), .B(n8882), .ZN(n7984)
         );
  OAI22_X1 U9697 ( .A1(n8885), .A2(n7979), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5347), .ZN(n7982) );
  OAI22_X1 U9698 ( .A1(n8710), .A2(n8887), .B1(n8875), .B2(n7980), .ZN(n7981)
         );
  AOI211_X1 U9699 ( .C1(n8704), .C2(n8890), .A(n7982), .B(n7981), .ZN(n7983)
         );
  NAND2_X1 U9700 ( .A1(n7984), .A2(n7983), .ZN(P2_U3236) );
  NAND2_X1 U9701 ( .A1(n7989), .A2(n7985), .ZN(n7986) );
  OAI211_X1 U9702 ( .C1(n7987), .C2(n9379), .A(n7986), .B(n8803), .ZN(P2_U3335) );
  NAND2_X1 U9703 ( .A1(n7989), .A2(n7988), .ZN(n7991) );
  OR2_X1 U9704 ( .A1(n7990), .A2(P1_U3084), .ZN(n8554) );
  OAI211_X1 U9705 ( .C1(n7993), .C2(n7992), .A(n7991), .B(n8554), .ZN(P1_U3330) );
  NOR2_X1 U9706 ( .A1(n7995), .A2(n7994), .ZN(n7997) );
  NOR2_X1 U9707 ( .A1(n7997), .A2(n7996), .ZN(n8074) );
  XNOR2_X1 U9708 ( .A(n8074), .B(n8080), .ZN(n7998) );
  NOR2_X1 U9709 ( .A1(n8040), .A2(n7998), .ZN(n8075) );
  AOI211_X1 U9710 ( .C1(n7998), .C2(n8040), .A(n8075), .B(n10003), .ZN(n8005)
         );
  OAI21_X1 U9711 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n8000), .A(n7999), .ZN(
        n8079) );
  XNOR2_X1 U9712 ( .A(n8080), .B(n8079), .ZN(n8001) );
  NOR2_X1 U9713 ( .A1(n6072), .A2(n8001), .ZN(n8081) );
  AOI211_X1 U9714 ( .C1(n8001), .C2(n6072), .A(n8081), .B(n9969), .ZN(n8004)
         );
  NAND2_X1 U9715 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8068) );
  NAND2_X1 U9716 ( .A1(n10013), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n8002) );
  OAI211_X1 U9717 ( .C1(n9525), .C2(n8080), .A(n8068), .B(n8002), .ZN(n8003)
         );
  OR3_X1 U9718 ( .A1(n8005), .A2(n8004), .A3(n8003), .ZN(P1_U3256) );
  XNOR2_X1 U9719 ( .A(n8711), .B(n9265), .ZN(n8010) );
  INV_X1 U9720 ( .A(n8704), .ZN(n9891) );
  AOI21_X1 U9721 ( .B1(n8010), .B2(n8007), .A(n8167), .ZN(n9884) );
  NAND2_X1 U9722 ( .A1(n8704), .A2(n8093), .ZN(n8009) );
  INV_X1 U9723 ( .A(n8010), .ZN(n8708) );
  NAND2_X1 U9724 ( .A1(n8011), .A2(n8708), .ZN(n8012) );
  NAND3_X1 U9725 ( .A1(n8162), .A2(n9269), .A3(n8012), .ZN(n8014) );
  AOI22_X1 U9726 ( .A1(n8901), .A2(n9266), .B1(n9264), .B2(n8902), .ZN(n8013)
         );
  NAND2_X1 U9727 ( .A1(n8014), .A2(n8013), .ZN(n9888) );
  XNOR2_X1 U9728 ( .A(n8172), .B(n8711), .ZN(n9886) );
  OAI22_X1 U9729 ( .A1(n9244), .A2(n8015), .B1(n8100), .B2(n9241), .ZN(n8016)
         );
  AOI21_X1 U9730 ( .B1(n8711), .B2(n9246), .A(n8016), .ZN(n8017) );
  OAI21_X1 U9731 ( .B1(n9886), .B2(n9218), .A(n8017), .ZN(n8018) );
  AOI21_X1 U9732 ( .B1(n9888), .B2(n9238), .A(n8018), .ZN(n8019) );
  OAI21_X1 U9733 ( .B1(n9884), .B2(n9274), .A(n8019), .ZN(P2_U3282) );
  INV_X1 U9734 ( .A(n8020), .ZN(n8024) );
  OAI222_X1 U9735 ( .A1(n9835), .A2(n8024), .B1(P1_U3084), .B2(n8022), .C1(
        n8021), .C2(n9831), .ZN(P1_U3329) );
  OAI222_X1 U9736 ( .A1(P2_U3152), .A2(n8025), .B1(n4451), .B2(n8024), .C1(
        n8023), .C2(n9379), .ZN(P2_U3334) );
  AOI211_X1 U9737 ( .C1(n10149), .C2(n8028), .A(n8027), .B(n8026), .ZN(n8029)
         );
  OAI21_X1 U9738 ( .B1(n10141), .B2(n8030), .A(n8029), .ZN(n8032) );
  NAND2_X1 U9739 ( .A1(n8032), .A2(n10173), .ZN(n8031) );
  OAI21_X1 U9740 ( .B1(n10173), .B2(n7329), .A(n8031), .ZN(P1_U3535) );
  NAND2_X1 U9741 ( .A1(n8032), .A2(n10160), .ZN(n8033) );
  OAI21_X1 U9742 ( .B1(n10160), .B2(n8034), .A(n8033), .ZN(P1_U3490) );
  OAI21_X1 U9743 ( .B1(n8408), .B2(n8035), .A(n8049), .ZN(n8038) );
  NAND2_X1 U9744 ( .A1(n9488), .A2(n10045), .ZN(n8036) );
  OAI21_X1 U9745 ( .B1(n9427), .B2(n9716), .A(n8036), .ZN(n8037) );
  AOI21_X1 U9746 ( .B1(n8038), .B2(n10050), .A(n8037), .ZN(n9917) );
  AOI21_X1 U9747 ( .B1(n8408), .B2(n8039), .A(n4535), .ZN(n9922) );
  NAND2_X1 U9748 ( .A1(n9922), .A2(n9611), .ZN(n8048) );
  OAI22_X1 U9749 ( .A1(n10057), .A2(n8040), .B1(n8069), .B2(n10036), .ZN(n8045) );
  INV_X1 U9750 ( .A(n8056), .ZN(n8041) );
  OAI211_X1 U9751 ( .C1(n9918), .C2(n8042), .A(n8041), .B(n10124), .ZN(n9916)
         );
  NOR2_X1 U9752 ( .A1(n9738), .A2(n10044), .ZN(n9720) );
  INV_X1 U9753 ( .A(n9720), .ZN(n8043) );
  NOR2_X1 U9754 ( .A1(n9916), .A2(n8043), .ZN(n8044) );
  AOI211_X1 U9755 ( .C1(n9739), .C2(n8046), .A(n8045), .B(n8044), .ZN(n8047)
         );
  OAI211_X1 U9756 ( .C1(n9738), .C2(n9917), .A(n8048), .B(n8047), .ZN(P1_U3276) );
  NAND2_X1 U9757 ( .A1(n8049), .A2(n8322), .ZN(n8050) );
  XOR2_X1 U9758 ( .A(n8271), .B(n8050), .Z(n8051) );
  AOI222_X1 U9759 ( .A1(n10050), .A2(n8051), .B1(n9486), .B2(n10046), .C1(
        n9487), .C2(n10045), .ZN(n9912) );
  OAI21_X1 U9760 ( .B1(n8053), .B2(n8271), .A(n8052), .ZN(n8054) );
  INV_X1 U9761 ( .A(n8054), .ZN(n9915) );
  NAND2_X1 U9762 ( .A1(n9915), .A2(n9611), .ZN(n8062) );
  INV_X1 U9763 ( .A(n8055), .ZN(n8123) );
  OAI22_X1 U9764 ( .A1(n10057), .A2(n6566), .B1(n8123), .B2(n10036), .ZN(n8059) );
  OAI211_X1 U9765 ( .C1(n8056), .C2(n9913), .A(n10124), .B(n9735), .ZN(n9911)
         );
  NOR2_X1 U9766 ( .A1(n9911), .A2(n8057), .ZN(n8058) );
  AOI211_X1 U9767 ( .C1(n9739), .C2(n8060), .A(n8059), .B(n8058), .ZN(n8061)
         );
  OAI211_X1 U9768 ( .C1(n9912), .C2(n9738), .A(n8062), .B(n8061), .ZN(P1_U3275) );
  XNOR2_X1 U9769 ( .A(n8065), .B(n8064), .ZN(n8066) );
  XNOR2_X1 U9770 ( .A(n8063), .B(n8066), .ZN(n8067) );
  NAND2_X1 U9771 ( .A1(n8067), .A2(n9467), .ZN(n8073) );
  INV_X1 U9772 ( .A(n8068), .ZN(n8071) );
  OAI22_X1 U9773 ( .A1(n9455), .A2(n8300), .B1(n9472), .B2(n8069), .ZN(n8070)
         );
  AOI211_X1 U9774 ( .C1(n8126), .C2(n9731), .A(n8071), .B(n8070), .ZN(n8072)
         );
  OAI211_X1 U9775 ( .C1(n9918), .C2(n9478), .A(n8073), .B(n8072), .ZN(P1_U3239) );
  NOR2_X1 U9776 ( .A1(n8074), .A2(n8080), .ZN(n8076) );
  NOR2_X1 U9777 ( .A1(n8076), .A2(n8075), .ZN(n8078) );
  MUX2_X1 U9778 ( .A(n6566), .B(P1_REG2_REG_16__SCAN_IN), .S(n9518), .Z(n8077)
         );
  NOR2_X1 U9779 ( .A1(n8078), .A2(n8077), .ZN(n9514) );
  AOI211_X1 U9780 ( .C1(n8078), .C2(n8077), .A(n10003), .B(n9514), .ZN(n8092)
         );
  NOR2_X1 U9781 ( .A1(n8080), .A2(n8079), .ZN(n8082) );
  NOR2_X1 U9782 ( .A1(n8082), .A2(n8081), .ZN(n8085) );
  INV_X1 U9783 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8083) );
  MUX2_X1 U9784 ( .A(n8083), .B(P1_REG1_REG_16__SCAN_IN), .S(n9518), .Z(n8084)
         );
  NOR2_X1 U9785 ( .A1(n8085), .A2(n8084), .ZN(n9517) );
  AOI211_X1 U9786 ( .C1(n8085), .C2(n8084), .A(n9969), .B(n9517), .ZN(n8091)
         );
  NOR2_X1 U9787 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8086), .ZN(n8125) );
  INV_X1 U9788 ( .A(n8125), .ZN(n8088) );
  NAND2_X1 U9789 ( .A1(n10013), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n8087) );
  OAI211_X1 U9790 ( .C1(n9525), .C2(n8089), .A(n8088), .B(n8087), .ZN(n8090)
         );
  OR3_X1 U9791 ( .A1(n8092), .A2(n8091), .A3(n8090), .ZN(P1_U3257) );
  INV_X1 U9792 ( .A(n7976), .ZN(n8096) );
  NOR3_X1 U9793 ( .A1(n8094), .A2(n8093), .A3(n8892), .ZN(n8095) );
  AOI21_X1 U9794 ( .B1(n8096), .B2(n8882), .A(n8095), .ZN(n8106) );
  AOI22_X1 U9795 ( .A1(n8097), .A2(n8901), .B1(n8894), .B2(n8902), .ZN(n8099)
         );
  OAI211_X1 U9796 ( .C1(n8885), .C2(n8100), .A(n8099), .B(n8098), .ZN(n8103)
         );
  NOR2_X1 U9797 ( .A1(n8101), .A2(n8868), .ZN(n8102) );
  AOI211_X1 U9798 ( .C1(n8711), .C2(n8890), .A(n8103), .B(n8102), .ZN(n8104)
         );
  OAI21_X1 U9799 ( .B1(n8106), .B2(n8105), .A(n8104), .ZN(P2_U3217) );
  XNOR2_X1 U9800 ( .A(n8107), .B(n8249), .ZN(n9805) );
  INV_X1 U9801 ( .A(n9719), .ZN(n8108) );
  AOI211_X1 U9802 ( .C1(n9803), .C2(n9736), .A(n10154), .B(n8108), .ZN(n9802)
         );
  INV_X1 U9803 ( .A(n9803), .ZN(n9479) );
  NOR2_X1 U9804 ( .A1(n9479), .A2(n9724), .ZN(n8111) );
  OAI22_X1 U9805 ( .A1(n10057), .A2(n8109), .B1(n9471), .B2(n10036), .ZN(n8110) );
  AOI211_X1 U9806 ( .C1(n9802), .C2(n9720), .A(n8111), .B(n8110), .ZN(n8117)
         );
  INV_X1 U9807 ( .A(n8251), .ZN(n8112) );
  AOI21_X1 U9808 ( .B1(n9730), .B2(n8250), .A(n8112), .ZN(n8113) );
  XNOR2_X1 U9809 ( .A(n8113), .B(n8249), .ZN(n8114) );
  OAI222_X1 U9810 ( .A1(n6463), .A2(n8115), .B1(n9716), .B2(n9708), .C1(n6466), 
        .C2(n8114), .ZN(n9801) );
  NAND2_X1 U9811 ( .A1(n9801), .A2(n10031), .ZN(n8116) );
  OAI211_X1 U9812 ( .C1(n9805), .C2(n9746), .A(n8117), .B(n8116), .ZN(P1_U3273) );
  NAND2_X1 U9813 ( .A1(n6103), .A2(n8120), .ZN(n8121) );
  XNOR2_X1 U9814 ( .A(n8118), .B(n8121), .ZN(n8122) );
  NAND2_X1 U9815 ( .A1(n8122), .A2(n9467), .ZN(n8128) );
  OAI22_X1 U9816 ( .A1(n9455), .A2(n8133), .B1(n9472), .B2(n8123), .ZN(n8124)
         );
  AOI211_X1 U9817 ( .C1(n8126), .C2(n9486), .A(n8125), .B(n8124), .ZN(n8127)
         );
  OAI211_X1 U9818 ( .C1(n9913), .C2(n9478), .A(n8128), .B(n8127), .ZN(P1_U3224) );
  AOI22_X1 U9819 ( .A1(n9475), .A2(n9489), .B1(n8130), .B2(n8129), .ZN(n8132)
         );
  OAI211_X1 U9820 ( .C1(n8133), .C2(n9473), .A(n8132), .B(n8131), .ZN(n8139)
         );
  AOI21_X1 U9821 ( .B1(n8137), .B2(n8135), .A(n8134), .ZN(n8136) );
  AOI211_X1 U9822 ( .C1(n4533), .C2(n8137), .A(n9461), .B(n8136), .ZN(n8138)
         );
  AOI211_X1 U9823 ( .C1(n9459), .C2(n9808), .A(n8139), .B(n8138), .ZN(n8140)
         );
  INV_X1 U9824 ( .A(n8140), .ZN(P1_U3213) );
  NAND2_X1 U9825 ( .A1(n8857), .A2(n8901), .ZN(n8144) );
  NAND2_X1 U9826 ( .A1(n8882), .A2(n8141), .ZN(n8143) );
  MUX2_X1 U9827 ( .A(n8144), .B(n8143), .S(n8142), .Z(n8149) );
  OAI22_X1 U9828 ( .A1(n8885), .A2(n9257), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8145), .ZN(n8147) );
  OAI22_X1 U9829 ( .A1(n9232), .A2(n8887), .B1(n8875), .B2(n8710), .ZN(n8146)
         );
  AOI211_X1 U9830 ( .C1(n9350), .C2(n8890), .A(n8147), .B(n8146), .ZN(n8148)
         );
  NAND2_X1 U9831 ( .A1(n8149), .A2(n8148), .ZN(P2_U3243) );
  INV_X1 U9832 ( .A(n8150), .ZN(n8155) );
  OAI222_X1 U9833 ( .A1(P2_U3152), .A2(n8152), .B1(n4451), .B2(n8155), .C1(
        n8151), .C2(n9379), .ZN(P2_U3333) );
  OAI222_X1 U9834 ( .A1(n9831), .A2(n8156), .B1(n9835), .B2(n8155), .C1(n8154), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U9835 ( .A(n8157), .ZN(n8181) );
  INV_X1 U9836 ( .A(n8158), .ZN(n8160) );
  OAI222_X1 U9837 ( .A1(n9835), .A2(n8181), .B1(P1_U3084), .B2(n8160), .C1(
        n8159), .C2(n9831), .ZN(P1_U3327) );
  OR2_X1 U9838 ( .A1(n9345), .A2(n9232), .ZN(n8720) );
  NAND2_X1 U9839 ( .A1(n9345), .A2(n9232), .ZN(n9224) );
  OR2_X1 U9840 ( .A1(n8711), .A2(n8710), .ZN(n8161) );
  OR2_X1 U9841 ( .A1(n9350), .A2(n8186), .ZN(n8715) );
  INV_X1 U9842 ( .A(n8715), .ZN(n8164) );
  OR2_X1 U9843 ( .A1(n9263), .A2(n8164), .ZN(n8163) );
  NAND2_X1 U9844 ( .A1(n9350), .A2(n8186), .ZN(n8716) );
  NAND2_X1 U9845 ( .A1(n8163), .A2(n8716), .ZN(n8165) );
  INV_X1 U9846 ( .A(n8718), .ZN(n8628) );
  OAI21_X1 U9847 ( .B1(n8718), .B2(n8165), .A(n9225), .ZN(n8166) );
  INV_X1 U9848 ( .A(n8874), .ZN(n9209) );
  AOI222_X1 U9849 ( .A1(n9269), .A2(n8166), .B1(n9209), .B2(n9266), .C1(n8901), 
        .C2(n9264), .ZN(n9348) );
  INV_X1 U9850 ( .A(n8711), .ZN(n9885) );
  AOI21_X1 U9851 ( .B1(n8718), .B2(n8169), .A(n9005), .ZN(n9344) );
  OAI21_X1 U9852 ( .B1(n10198), .B2(n8170), .A(n9250), .ZN(n8171) );
  NAND2_X1 U9853 ( .A1(n9344), .A2(n8171), .ZN(n8179) );
  INV_X1 U9854 ( .A(n9350), .ZN(n9261) );
  NAND2_X1 U9855 ( .A1(n9253), .A2(n9261), .ZN(n9254) );
  INV_X1 U9856 ( .A(n9235), .ZN(n8173) );
  AOI21_X1 U9857 ( .B1(n9345), .B2(n9254), .A(n8173), .ZN(n9346) );
  INV_X1 U9858 ( .A(n9345), .ZN(n8174) );
  NOR2_X1 U9859 ( .A1(n8174), .A2(n9260), .ZN(n8177) );
  OAI22_X1 U9860 ( .A1(n9244), .A2(n8175), .B1(n8185), .B2(n9241), .ZN(n8176)
         );
  AOI211_X1 U9861 ( .C1(n9346), .C2(n9272), .A(n8177), .B(n8176), .ZN(n8178)
         );
  OAI211_X1 U9862 ( .C1(n10198), .C2(n9348), .A(n8179), .B(n8178), .ZN(
        P2_U3280) );
  OAI222_X1 U9863 ( .A1(n8182), .A2(P2_U3152), .B1(n4451), .B2(n8181), .C1(
        n8180), .C2(n9379), .ZN(P2_U3332) );
  XOR2_X1 U9864 ( .A(n8183), .B(n8184), .Z(n8190) );
  OAI22_X1 U9865 ( .A1(n8885), .A2(n8185), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8955), .ZN(n8188) );
  OAI22_X1 U9866 ( .A1(n8874), .A2(n8887), .B1(n8875), .B2(n8186), .ZN(n8187)
         );
  AOI211_X1 U9867 ( .C1(n9345), .C2(n8890), .A(n8188), .B(n8187), .ZN(n8189)
         );
  OAI21_X1 U9868 ( .B1(n8190), .B2(n8868), .A(n8189), .ZN(P2_U3228) );
  OAI22_X1 U9869 ( .A1(n9598), .A2(n8199), .B1(n9575), .B2(n6265), .ZN(n8191)
         );
  XNOR2_X1 U9870 ( .A(n8191), .B(n8200), .ZN(n8193) );
  OAI22_X1 U9871 ( .A1(n9598), .A2(n6265), .B1(n9575), .B2(n8202), .ZN(n8192)
         );
  NOR2_X1 U9872 ( .A1(n8193), .A2(n8192), .ZN(n8198) );
  AOI21_X1 U9873 ( .B1(n8193), .B2(n8192), .A(n8198), .ZN(n9382) );
  INV_X1 U9874 ( .A(n8194), .ZN(n8196) );
  OR2_X1 U9875 ( .A1(n8196), .A2(n8195), .ZN(n9383) );
  INV_X1 U9876 ( .A(n9584), .ZN(n9748) );
  OAI22_X1 U9877 ( .A1(n9748), .A2(n8199), .B1(n9589), .B2(n6265), .ZN(n8201)
         );
  XNOR2_X1 U9878 ( .A(n8201), .B(n8200), .ZN(n8204) );
  OAI22_X1 U9879 ( .A1(n9748), .A2(n5802), .B1(n9589), .B2(n8202), .ZN(n8203)
         );
  OAI22_X1 U9880 ( .A1(n9455), .A2(n9575), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8206), .ZN(n8208) );
  OAI22_X1 U9881 ( .A1(n9473), .A2(n9574), .B1(n9472), .B2(n9581), .ZN(n8207)
         );
  AOI211_X1 U9882 ( .C1(n9584), .C2(n9459), .A(n8208), .B(n8207), .ZN(n8209)
         );
  OAI21_X1 U9883 ( .B1(n8210), .B2(n9461), .A(n8209), .ZN(P1_U3218) );
  INV_X1 U9884 ( .A(n9336), .ZN(n9213) );
  INV_X1 U9885 ( .A(n9332), .ZN(n9013) );
  INV_X1 U9886 ( .A(n9316), .ZN(n9154) );
  NAND2_X1 U9887 ( .A1(n9378), .A2(n8233), .ZN(n8213) );
  OR2_X1 U9888 ( .A1(n8234), .A2(n9380), .ZN(n8212) );
  INV_X1 U9889 ( .A(SI_29_), .ZN(n8214) );
  AND2_X1 U9890 ( .A1(n8215), .A2(n8214), .ZN(n8218) );
  INV_X1 U9891 ( .A(n8215), .ZN(n8216) );
  NAND2_X1 U9892 ( .A1(n8216), .A2(SI_29_), .ZN(n8217) );
  INV_X1 U9893 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8589) );
  INV_X1 U9894 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8805) );
  MUX2_X1 U9895 ( .A(n8589), .B(n8805), .S(n8228), .Z(n8221) );
  INV_X1 U9896 ( .A(SI_30_), .ZN(n8220) );
  NAND2_X1 U9897 ( .A1(n8221), .A2(n8220), .ZN(n8225) );
  INV_X1 U9898 ( .A(n8221), .ZN(n8222) );
  NAND2_X1 U9899 ( .A1(n8222), .A2(SI_30_), .ZN(n8223) );
  NAND2_X1 U9900 ( .A1(n8225), .A2(n8223), .ZN(n8226) );
  NOR2_X1 U9901 ( .A1(n8234), .A2(n8805), .ZN(n8224) );
  OAI21_X1 U9902 ( .B1(n8227), .B2(n8226), .A(n8225), .ZN(n8232) );
  MUX2_X1 U9903 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8228), .Z(n8230) );
  INV_X1 U9904 ( .A(SI_31_), .ZN(n8229) );
  XNOR2_X1 U9905 ( .A(n8230), .B(n8229), .ZN(n8231) );
  XNOR2_X1 U9906 ( .A(n8232), .B(n8231), .ZN(n9371) );
  NAND2_X1 U9907 ( .A1(n9371), .A2(n8233), .ZN(n8236) );
  OR2_X1 U9908 ( .A1(n8234), .A2(n6914), .ZN(n8235) );
  INV_X1 U9909 ( .A(n6974), .ZN(n8238) );
  NAND2_X1 U9910 ( .A1(n8238), .A2(P2_B_REG_SCAN_IN), .ZN(n8239) );
  AND2_X1 U9911 ( .A1(n9266), .A2(n8239), .ZN(n9040) );
  NAND2_X1 U9912 ( .A1(n8605), .A2(n9040), .ZN(n9879) );
  NOR2_X1 U9913 ( .A1(n10198), .A2(n9879), .ZN(n9002) );
  NOR2_X1 U9914 ( .A1(n9244), .A2(n8240), .ZN(n8241) );
  AOI211_X1 U9915 ( .C1(n9275), .C2(n9246), .A(n9002), .B(n8241), .ZN(n8242)
         );
  OAI21_X1 U9916 ( .B1(n9277), .B2(n9218), .A(n8242), .ZN(P2_U3265) );
  NAND2_X1 U9917 ( .A1(n9371), .A2(n8283), .ZN(n8244) );
  OR2_X1 U9918 ( .A1(n5878), .A2(n6893), .ZN(n8243) );
  INV_X1 U9919 ( .A(n9558), .ZN(n8245) );
  NAND2_X1 U9920 ( .A1(n9876), .A2(n8245), .ZN(n8542) );
  INV_X1 U9921 ( .A(n8246), .ZN(n8248) );
  XNOR2_X1 U9922 ( .A(n9793), .B(n9484), .ZN(n8434) );
  INV_X1 U9923 ( .A(n8434), .ZN(n9704) );
  INV_X1 U9924 ( .A(n9713), .ZN(n8274) );
  INV_X1 U9925 ( .A(n8249), .ZN(n8273) );
  NAND4_X1 U9926 ( .A1(n8254), .A2(n8253), .A3(n8354), .A4(n8252), .ZN(n8257)
         );
  INV_X1 U9927 ( .A(n8308), .ZN(n8360) );
  NOR4_X1 U9928 ( .A1(n8257), .A2(n8256), .A3(n8255), .A4(n8360), .ZN(n8260)
         );
  INV_X1 U9929 ( .A(n8512), .ZN(n8259) );
  NAND4_X1 U9930 ( .A1(n8260), .A2(n8259), .A3(n4584), .A4(n8258), .ZN(n8262)
         );
  OR3_X1 U9931 ( .A1(n8262), .A2(n6388), .A3(n8261), .ZN(n8263) );
  NOR3_X1 U9932 ( .A1(n8265), .A2(n8264), .A3(n8263), .ZN(n8268) );
  INV_X1 U9933 ( .A(n8266), .ZN(n8267) );
  NAND4_X1 U9934 ( .A1(n8408), .A2(n8269), .A3(n8268), .A4(n8267), .ZN(n8270)
         );
  NOR2_X1 U9935 ( .A1(n8271), .A2(n8270), .ZN(n8272) );
  NAND4_X1 U9936 ( .A1(n8274), .A2(n8273), .A3(n9729), .A4(n8272), .ZN(n8275)
         );
  NOR2_X1 U9937 ( .A1(n9704), .A2(n8275), .ZN(n8276) );
  NAND3_X1 U9938 ( .A1(n9675), .A2(n8276), .A3(n9685), .ZN(n8277) );
  NOR2_X1 U9939 ( .A1(n9661), .A2(n8277), .ZN(n8278) );
  NAND3_X1 U9940 ( .A1(n9632), .A2(n9640), .A3(n8278), .ZN(n8279) );
  NOR2_X1 U9941 ( .A1(n9609), .A2(n8279), .ZN(n8280) );
  NAND3_X1 U9942 ( .A1(n9567), .A2(n4772), .A3(n8280), .ZN(n8281) );
  NOR2_X1 U9943 ( .A1(n8282), .A2(n8281), .ZN(n8288) );
  NAND2_X1 U9944 ( .A1(n8588), .A2(n8283), .ZN(n8285) );
  OR2_X1 U9945 ( .A1(n5878), .A2(n8589), .ZN(n8284) );
  OR2_X1 U9946 ( .A1(n8286), .A2(n6465), .ZN(n8538) );
  NAND2_X1 U9947 ( .A1(n8286), .A2(n6465), .ZN(n8539) );
  AND2_X1 U9948 ( .A1(n8538), .A2(n8539), .ZN(n8287) );
  NAND4_X1 U9949 ( .A1(n8544), .A2(n8542), .A3(n8288), .A4(n8287), .ZN(n8290)
         );
  NAND2_X1 U9950 ( .A1(n8538), .A2(n9558), .ZN(n8291) );
  NAND2_X1 U9951 ( .A1(n8292), .A2(n8470), .ZN(n8495) );
  AND2_X1 U9952 ( .A1(n8456), .A2(n8293), .ZN(n8464) );
  INV_X1 U9953 ( .A(n8464), .ZN(n8294) );
  NAND2_X1 U9954 ( .A1(n8294), .A2(n8467), .ZN(n8295) );
  NAND2_X1 U9955 ( .A1(n8471), .A2(n8295), .ZN(n8530) );
  OR2_X1 U9956 ( .A1(n9788), .A2(n9707), .ZN(n8330) );
  INV_X1 U9957 ( .A(n8296), .ZN(n8297) );
  NAND2_X1 U9958 ( .A1(n8330), .A2(n8297), .ZN(n8298) );
  NAND2_X1 U9959 ( .A1(n8298), .A2(n8436), .ZN(n8299) );
  NOR2_X1 U9960 ( .A1(n8433), .A2(n8299), .ZN(n8441) );
  INV_X1 U9961 ( .A(n8441), .ZN(n8336) );
  NOR2_X1 U9962 ( .A1(n8336), .A2(n4762), .ZN(n8496) );
  NAND2_X1 U9963 ( .A1(n9808), .A2(n8300), .ZN(n8317) );
  AND2_X1 U9964 ( .A1(n8317), .A2(n8301), .ZN(n8401) );
  INV_X1 U9965 ( .A(n8401), .ZN(n8404) );
  NAND2_X1 U9966 ( .A1(n8386), .A2(n8376), .ZN(n8302) );
  AND2_X1 U9967 ( .A1(n8302), .A2(n8385), .ZN(n8304) );
  INV_X1 U9968 ( .A(n8394), .ZN(n8303) );
  OR3_X1 U9969 ( .A1(n8404), .A2(n8304), .A3(n8303), .ZN(n8321) );
  NAND2_X1 U9970 ( .A1(n8375), .A2(n8363), .ZN(n8362) );
  NOR2_X1 U9971 ( .A1(n8321), .A2(n8362), .ZN(n8305) );
  AND2_X1 U9972 ( .A1(n8409), .A2(n8305), .ZN(n8306) );
  NAND2_X1 U9973 ( .A1(n8419), .A2(n8306), .ZN(n8497) );
  AND2_X1 U9974 ( .A1(n8310), .A2(n8307), .ZN(n8507) );
  NAND3_X1 U9975 ( .A1(n7254), .A2(n8507), .A3(n8514), .ZN(n8314) );
  NAND2_X1 U9976 ( .A1(n8512), .A2(n8308), .ZN(n8312) );
  NAND2_X1 U9977 ( .A1(n8509), .A2(n8511), .ZN(n8309) );
  NAND4_X1 U9978 ( .A1(n8310), .A2(n8309), .A3(n8308), .A4(n8354), .ZN(n8311)
         );
  AND2_X1 U9979 ( .A1(n8312), .A2(n8311), .ZN(n8313) );
  INV_X1 U9980 ( .A(n8515), .ZN(n8369) );
  AOI21_X1 U9981 ( .B1(n8314), .B2(n8313), .A(n8369), .ZN(n8327) );
  AND2_X1 U9982 ( .A1(n8411), .A2(n8315), .ZN(n8410) );
  AND2_X1 U9983 ( .A1(n8377), .A2(n8372), .ZN(n8367) );
  AND2_X1 U9984 ( .A1(n8385), .A2(n8367), .ZN(n8320) );
  AND2_X1 U9985 ( .A1(n8403), .A2(n8316), .ZN(n8397) );
  INV_X1 U9986 ( .A(n8397), .ZN(n8318) );
  NAND2_X1 U9987 ( .A1(n8318), .A2(n8317), .ZN(n8406) );
  OR2_X1 U9988 ( .A1(n8404), .A2(n8396), .ZN(n8319) );
  OAI211_X1 U9989 ( .C1(n8321), .C2(n8320), .A(n8406), .B(n8319), .ZN(n8323)
         );
  NAND2_X1 U9990 ( .A1(n8323), .A2(n8322), .ZN(n8325) );
  INV_X1 U9991 ( .A(n8412), .ZN(n8324) );
  AOI21_X1 U9992 ( .B1(n8410), .B2(n8325), .A(n8324), .ZN(n8326) );
  NAND2_X1 U9993 ( .A1(n8419), .A2(n8326), .ZN(n8517) );
  OAI21_X1 U9994 ( .B1(n8497), .B2(n8327), .A(n8517), .ZN(n8328) );
  AND2_X1 U9995 ( .A1(n8496), .A2(n8328), .ZN(n8337) );
  NAND2_X1 U9996 ( .A1(n8330), .A2(n8329), .ZN(n8437) );
  NAND2_X1 U9997 ( .A1(n8425), .A2(n8331), .ZN(n8428) );
  INV_X1 U9998 ( .A(n8417), .ZN(n8332) );
  OAI21_X1 U9999 ( .B1(n8428), .B2(n8332), .A(n8427), .ZN(n8333) );
  NOR2_X1 U10000 ( .A1(n8437), .A2(n8333), .ZN(n8335) );
  OAI211_X1 U10001 ( .C1(n8336), .C2(n8335), .A(n8334), .B(n8446), .ZN(n8525)
         );
  OAI21_X1 U10002 ( .B1(n8337), .B2(n8525), .A(n8447), .ZN(n8338) );
  NAND2_X1 U10003 ( .A1(n8338), .A2(n8444), .ZN(n8339) );
  NAND2_X1 U10004 ( .A1(n8339), .A2(n8349), .ZN(n8340) );
  AND4_X1 U10005 ( .A1(n8467), .A2(n8458), .A3(n8460), .A4(n8340), .ZN(n8341)
         );
  NOR2_X1 U10006 ( .A1(n8530), .A2(n8341), .ZN(n8343) );
  NAND2_X1 U10007 ( .A1(n9480), .A2(n9558), .ZN(n8342) );
  NAND2_X1 U10008 ( .A1(n8286), .A2(n8342), .ZN(n8487) );
  OAI211_X1 U10009 ( .C1(n8495), .C2(n8343), .A(n8487), .B(n8534), .ZN(n8344)
         );
  NAND2_X1 U10010 ( .A1(n8486), .A2(n8344), .ZN(n8345) );
  NAND3_X1 U10011 ( .A1(n8345), .A2(n8500), .A3(n8544), .ZN(n8346) );
  NAND2_X1 U10012 ( .A1(n4523), .A2(n8346), .ZN(n8493) );
  NAND2_X1 U10013 ( .A1(n8533), .A2(n4545), .ZN(n8455) );
  NAND2_X1 U10014 ( .A1(n9630), .A2(n8448), .ZN(n8348) );
  NAND2_X1 U10015 ( .A1(n8529), .A2(n8348), .ZN(n8352) );
  INV_X1 U10016 ( .A(n8444), .ZN(n8350) );
  OAI21_X1 U10017 ( .B1(n8350), .B2(n8447), .A(n8349), .ZN(n8351) );
  INV_X1 U10018 ( .A(n8353), .ZN(n8355) );
  OAI21_X1 U10019 ( .B1(n8356), .B2(n8355), .A(n8354), .ZN(n8358) );
  NOR2_X1 U10020 ( .A1(n8361), .A2(n8360), .ZN(n8365) );
  MUX2_X1 U10021 ( .A(n8363), .B(n8362), .S(n8482), .Z(n8364) );
  INV_X1 U10022 ( .A(n8374), .ZN(n8368) );
  INV_X1 U10023 ( .A(n8376), .ZN(n8366) );
  AOI21_X1 U10024 ( .B1(n8368), .B2(n8367), .A(n8366), .ZN(n8382) );
  AOI21_X1 U10025 ( .B1(n8371), .B2(n8370), .A(n8369), .ZN(n8373) );
  OAI21_X1 U10026 ( .B1(n8374), .B2(n8373), .A(n8372), .ZN(n8380) );
  AND2_X1 U10027 ( .A1(n8376), .A2(n8375), .ZN(n8379) );
  INV_X1 U10028 ( .A(n8377), .ZN(n8378) );
  AOI21_X1 U10029 ( .B1(n8380), .B2(n8379), .A(n8378), .ZN(n8381) );
  NAND2_X1 U10030 ( .A1(n8384), .A2(n8383), .ZN(n8391) );
  MUX2_X1 U10031 ( .A(n8386), .B(n8385), .S(n8482), .Z(n8387) );
  AND3_X1 U10032 ( .A1(n8389), .A2(n8388), .A3(n8387), .ZN(n8390) );
  INV_X1 U10033 ( .A(n8392), .ZN(n8393) );
  INV_X1 U10034 ( .A(n8395), .ZN(n8399) );
  NAND3_X1 U10035 ( .A1(n8397), .A2(n8396), .A3(n4545), .ZN(n8398) );
  OAI22_X1 U10036 ( .A1(n8400), .A2(n4545), .B1(n8399), .B2(n8398), .ZN(n8402)
         );
  NAND2_X1 U10037 ( .A1(n8404), .A2(n8403), .ZN(n8405) );
  MUX2_X1 U10038 ( .A(n8406), .B(n8405), .S(n4545), .Z(n8407) );
  MUX2_X1 U10039 ( .A(n8410), .B(n8409), .S(n8482), .Z(n8415) );
  MUX2_X1 U10040 ( .A(n8412), .B(n8411), .S(n8482), .Z(n8413) );
  INV_X1 U10041 ( .A(n8413), .ZN(n8414) );
  INV_X1 U10042 ( .A(n9740), .ZN(n9737) );
  AOI21_X1 U10043 ( .B1(n8421), .B2(n9737), .A(n8417), .ZN(n8418) );
  MUX2_X1 U10044 ( .A(n8419), .B(n8418), .S(n4545), .Z(n8423) );
  MUX2_X1 U10045 ( .A(n8482), .B(n9740), .S(n9486), .Z(n8420) );
  AOI21_X1 U10046 ( .B1(n8421), .B2(n8420), .A(n9713), .ZN(n8422) );
  NAND2_X1 U10047 ( .A1(n8423), .A2(n8422), .ZN(n8432) );
  NAND2_X1 U10048 ( .A1(n8427), .A2(n8424), .ZN(n8426) );
  NAND2_X1 U10049 ( .A1(n8426), .A2(n8425), .ZN(n8430) );
  NAND2_X1 U10050 ( .A1(n8428), .A2(n8427), .ZN(n8429) );
  MUX2_X1 U10051 ( .A(n8430), .B(n8429), .S(n4545), .Z(n8431) );
  NAND2_X1 U10052 ( .A1(n8432), .A2(n8431), .ZN(n8435) );
  INV_X1 U10053 ( .A(n8433), .ZN(n8440) );
  NAND4_X1 U10054 ( .A1(n8435), .A2(n8440), .A3(n9685), .A4(n8434), .ZN(n8445)
         );
  NAND2_X1 U10055 ( .A1(n8437), .A2(n8436), .ZN(n8438) );
  NAND2_X1 U10056 ( .A1(n8446), .A2(n8438), .ZN(n8439) );
  NAND2_X1 U10057 ( .A1(n8440), .A2(n8439), .ZN(n8442) );
  MUX2_X1 U10058 ( .A(n8442), .B(n8441), .S(n4545), .Z(n8443) );
  NAND3_X1 U10059 ( .A1(n8445), .A2(n8444), .A3(n8443), .ZN(n8451) );
  OR2_X1 U10060 ( .A1(n8446), .A2(n8482), .ZN(n8450) );
  NAND2_X1 U10061 ( .A1(n9630), .A2(n8447), .ZN(n8523) );
  OR2_X1 U10062 ( .A1(n8523), .A2(n8448), .ZN(n8449) );
  AOI21_X1 U10063 ( .B1(n8451), .B2(n8450), .A(n8449), .ZN(n8453) );
  INV_X1 U10064 ( .A(n9609), .ZN(n8452) );
  NAND2_X1 U10065 ( .A1(n8457), .A2(n8456), .ZN(n8466) );
  INV_X1 U10066 ( .A(n8458), .ZN(n8463) );
  INV_X1 U10067 ( .A(n8459), .ZN(n8527) );
  NAND2_X1 U10068 ( .A1(n8460), .A2(n8527), .ZN(n8461) );
  NOR2_X1 U10069 ( .A1(n9594), .A2(n8461), .ZN(n8462) );
  OAI22_X1 U10070 ( .A1(n8466), .A2(n8465), .B1(n8464), .B2(n4545), .ZN(n8469)
         );
  OR2_X1 U10071 ( .A1(n8467), .A2(n4545), .ZN(n8468) );
  NAND3_X1 U10072 ( .A1(n8469), .A2(n9567), .A3(n8468), .ZN(n8473) );
  MUX2_X1 U10073 ( .A(n8471), .B(n8470), .S(n4545), .Z(n8472) );
  INV_X1 U10074 ( .A(n8481), .ZN(n8476) );
  INV_X1 U10075 ( .A(n9574), .ZN(n9481) );
  AND2_X1 U10076 ( .A1(n8487), .A2(n9481), .ZN(n8475) );
  INV_X1 U10077 ( .A(n8486), .ZN(n8474) );
  AOI21_X1 U10078 ( .B1(n8476), .B2(n8475), .A(n8474), .ZN(n8480) );
  NAND2_X1 U10079 ( .A1(n8486), .A2(n8483), .ZN(n8477) );
  OAI21_X1 U10080 ( .B1(n8481), .B2(n8477), .A(n8487), .ZN(n8478) );
  NAND2_X1 U10081 ( .A1(n8478), .A2(n8542), .ZN(n8479) );
  INV_X1 U10082 ( .A(n8483), .ZN(n8584) );
  NAND3_X1 U10083 ( .A1(n8481), .A2(n8584), .A3(n9574), .ZN(n8488) );
  MUX2_X1 U10084 ( .A(n9481), .B(n8483), .S(n8482), .Z(n8484) );
  INV_X1 U10085 ( .A(n8484), .ZN(n8485) );
  NAND4_X1 U10086 ( .A1(n8488), .A2(n8487), .A3(n8486), .A4(n8485), .ZN(n8489)
         );
  AND2_X1 U10087 ( .A1(n8489), .A2(n8544), .ZN(n8490) );
  INV_X1 U10088 ( .A(n8495), .ZN(n8537) );
  INV_X1 U10089 ( .A(n8496), .ZN(n8522) );
  INV_X1 U10090 ( .A(n8497), .ZN(n8520) );
  INV_X1 U10091 ( .A(n8498), .ZN(n8501) );
  NAND2_X1 U10092 ( .A1(n9499), .A2(n10092), .ZN(n8499) );
  NAND3_X1 U10093 ( .A1(n8501), .A2(n8500), .A3(n8499), .ZN(n8502) );
  NAND2_X1 U10094 ( .A1(n8503), .A2(n8502), .ZN(n8505) );
  OAI22_X1 U10095 ( .A1(n8506), .A2(n8505), .B1(n8504), .B2(n4969), .ZN(n8510)
         );
  INV_X1 U10096 ( .A(n8507), .ZN(n8508) );
  AOI21_X1 U10097 ( .B1(n8510), .B2(n8509), .A(n8508), .ZN(n8513) );
  OR3_X1 U10098 ( .A1(n8513), .A2(n4759), .A3(n8512), .ZN(n8516) );
  NAND3_X1 U10099 ( .A1(n8516), .A2(n8515), .A3(n8514), .ZN(n8519) );
  INV_X1 U10100 ( .A(n8517), .ZN(n8518) );
  AOI21_X1 U10101 ( .B1(n8520), .B2(n8519), .A(n8518), .ZN(n8521) );
  NOR2_X1 U10102 ( .A1(n8522), .A2(n8521), .ZN(n8526) );
  INV_X1 U10103 ( .A(n8523), .ZN(n8524) );
  OAI21_X1 U10104 ( .B1(n8526), .B2(n8525), .A(n8524), .ZN(n8528) );
  AOI21_X1 U10105 ( .B1(n8529), .B2(n8528), .A(n8527), .ZN(n8532) );
  INV_X1 U10106 ( .A(n8530), .ZN(n8531) );
  OAI21_X1 U10107 ( .B1(n8533), .B2(n8532), .A(n8531), .ZN(n8536) );
  INV_X1 U10108 ( .A(n8534), .ZN(n8535) );
  AOI21_X1 U10109 ( .B1(n8537), .B2(n8536), .A(n8535), .ZN(n8541) );
  INV_X1 U10110 ( .A(n8538), .ZN(n8540) );
  OAI21_X1 U10111 ( .B1(n8541), .B2(n8540), .A(n8539), .ZN(n8543) );
  NAND2_X1 U10112 ( .A1(n8543), .A2(n8542), .ZN(n8545) );
  NAND2_X1 U10113 ( .A1(n8545), .A2(n8544), .ZN(n8548) );
  INV_X1 U10114 ( .A(n8548), .ZN(n8547) );
  AOI21_X1 U10115 ( .B1(n8547), .B2(n4550), .A(n8554), .ZN(n8551) );
  NAND2_X1 U10116 ( .A1(n5022), .A2(n8549), .ZN(n8550) );
  NAND2_X1 U10117 ( .A1(n8553), .A2(n8552), .ZN(n8562) );
  OR2_X1 U10118 ( .A1(n6302), .A2(n9977), .ZN(n8559) );
  INV_X1 U10119 ( .A(n8554), .ZN(n8557) );
  INV_X1 U10120 ( .A(P1_B_REG_SCAN_IN), .ZN(n8555) );
  AOI21_X1 U10121 ( .B1(n8557), .B2(n8556), .A(n8555), .ZN(n8558) );
  OAI21_X1 U10122 ( .B1(n8560), .B2(n8559), .A(n8558), .ZN(n8561) );
  NAND2_X1 U10123 ( .A1(n8562), .A2(n8561), .ZN(P1_U3240) );
  NAND3_X1 U10124 ( .A1(n8564), .A2(n8857), .A3(n9008), .ZN(n8565) );
  OAI21_X1 U10125 ( .B1(n8563), .B2(n8868), .A(n8565), .ZN(n8568) );
  INV_X1 U10126 ( .A(n8566), .ZN(n8567) );
  NAND2_X1 U10127 ( .A1(n8568), .A2(n8567), .ZN(n8574) );
  NOR2_X1 U10128 ( .A1(n8885), .A2(n9193), .ZN(n8572) );
  INV_X1 U10129 ( .A(n9175), .ZN(n9015) );
  AOI22_X1 U10130 ( .A1(n9015), .A2(n9266), .B1(n9264), .B2(n9008), .ZN(n9199)
         );
  OAI22_X1 U10131 ( .A1(n8570), .A2(n9199), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8569), .ZN(n8571) );
  AOI211_X1 U10132 ( .C1(n9332), .C2(n8890), .A(n8572), .B(n8571), .ZN(n8573)
         );
  OAI211_X1 U10133 ( .C1(n8868), .C2(n8575), .A(n8574), .B(n8573), .ZN(
        P2_U3221) );
  INV_X1 U10134 ( .A(n8576), .ZN(n8579) );
  OAI222_X1 U10135 ( .A1(n9835), .A2(n8579), .B1(P1_U3084), .B2(n9977), .C1(
        n8577), .C2(n9831), .ZN(P1_U3326) );
  OAI222_X1 U10136 ( .A1(n6974), .A2(P2_U3152), .B1(n4451), .B2(n8579), .C1(
        n8578), .C2(n9379), .ZN(P2_U3331) );
  INV_X1 U10137 ( .A(n8581), .ZN(n8582) );
  AOI22_X1 U10138 ( .A1(n9738), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8582), .B2(
        n10041), .ZN(n8583) );
  OAI21_X1 U10139 ( .B1(n8584), .B2(n9724), .A(n8583), .ZN(n8585) );
  OAI21_X1 U10140 ( .B1(n8580), .B2(n9746), .A(n8587), .ZN(P1_U3355) );
  INV_X1 U10141 ( .A(n8588), .ZN(n8806) );
  OAI222_X1 U10142 ( .A1(n9831), .A2(n8589), .B1(n9835), .B2(n8806), .C1(
        P1_U3084), .C2(n4546), .ZN(P1_U3323) );
  NAND2_X1 U10143 ( .A1(n9247), .A2(n8874), .ZN(n8724) );
  NAND2_X1 U10144 ( .A1(n8725), .A2(n8724), .ZN(n9226) );
  INV_X1 U10145 ( .A(n9224), .ZN(n8590) );
  NOR2_X1 U10146 ( .A1(n9226), .A2(n8590), .ZN(n8591) );
  OR2_X1 U10147 ( .A1(n9336), .A2(n9230), .ZN(n8731) );
  NAND2_X1 U10148 ( .A1(n9336), .A2(n9230), .ZN(n8730) );
  NAND2_X1 U10149 ( .A1(n9206), .A2(n8730), .ZN(n9198) );
  OR2_X1 U10150 ( .A1(n9332), .A2(n9012), .ZN(n8737) );
  NAND2_X1 U10151 ( .A1(n9332), .A2(n9012), .ZN(n8740) );
  NAND2_X1 U10152 ( .A1(n9198), .A2(n9197), .ZN(n8592) );
  NAND2_X1 U10153 ( .A1(n9325), .A2(n9175), .ZN(n8741) );
  NAND2_X1 U10154 ( .A1(n8745), .A2(n8741), .ZN(n9186) );
  XNOR2_X1 U10155 ( .A(n9017), .B(n9016), .ZN(n9173) );
  NAND2_X1 U10156 ( .A1(n9316), .A2(n9176), .ZN(n8750) );
  NAND2_X1 U10157 ( .A1(n8735), .A2(n8750), .ZN(n9157) );
  AND2_X1 U10158 ( .A1(n9017), .A2(n9016), .ZN(n8747) );
  NOR2_X1 U10159 ( .A1(n9157), .A2(n8747), .ZN(n8593) );
  OR2_X1 U10160 ( .A1(n9311), .A2(n9021), .ZN(n8753) );
  NAND2_X1 U10161 ( .A1(n9311), .A2(n9021), .ZN(n8752) );
  NAND2_X1 U10162 ( .A1(n8753), .A2(n8752), .ZN(n9126) );
  INV_X1 U10163 ( .A(n9126), .ZN(n9132) );
  INV_X1 U10164 ( .A(n8752), .ZN(n8594) );
  NAND2_X1 U10165 ( .A1(n9304), .A2(n9136), .ZN(n8595) );
  NAND2_X1 U10166 ( .A1(n9024), .A2(n8595), .ZN(n9119) );
  NAND2_X1 U10167 ( .A1(n9117), .A2(n9136), .ZN(n9097) );
  NAND2_X1 U10168 ( .A1(n9301), .A2(n8851), .ZN(n8764) );
  NAND2_X1 U10169 ( .A1(n8761), .A2(n9085), .ZN(n8758) );
  NAND2_X1 U10170 ( .A1(n9295), .A2(n9072), .ZN(n8762) );
  NOR2_X1 U10171 ( .A1(n9290), .A2(n9031), .ZN(n8772) );
  NAND2_X1 U10172 ( .A1(n8596), .A2(n8774), .ZN(n8597) );
  NAND2_X1 U10173 ( .A1(n9047), .A2(n8899), .ZN(n8778) );
  NOR2_X1 U10174 ( .A1(n8605), .A2(n8598), .ZN(n8607) );
  INV_X1 U10175 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8602) );
  NAND2_X1 U10176 ( .A1(n5204), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8601) );
  NAND2_X1 U10177 ( .A1(n8599), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8600) );
  OAI211_X1 U10178 ( .C1(n8603), .C2(n8602), .A(n8601), .B(n8600), .ZN(n9039)
         );
  INV_X1 U10179 ( .A(n9039), .ZN(n8606) );
  OR2_X1 U10180 ( .A1(n9001), .A2(n8606), .ZN(n8782) );
  INV_X1 U10181 ( .A(n8605), .ZN(n8608) );
  OR2_X1 U10182 ( .A1(n9275), .A2(n8608), .ZN(n8788) );
  NAND2_X1 U10183 ( .A1(n9001), .A2(n8606), .ZN(n8780) );
  NAND2_X1 U10184 ( .A1(n4446), .A2(n8610), .ZN(n8798) );
  NOR2_X1 U10185 ( .A1(n8612), .A2(n4462), .ZN(n8617) );
  NAND2_X1 U10186 ( .A1(n7272), .A2(n8650), .ZN(n8660) );
  NOR2_X1 U10187 ( .A1(n8613), .A2(n8660), .ZN(n8616) );
  INV_X1 U10188 ( .A(n8614), .ZN(n8615) );
  NAND4_X1 U10189 ( .A1(n8617), .A2(n8616), .A3(n8615), .A4(n7456), .ZN(n8618)
         );
  NAND4_X1 U10190 ( .A1(n4525), .A2(n8675), .A3(n8620), .A4(n8619), .ZN(n8624)
         );
  NOR4_X1 U10191 ( .A1(n8624), .A2(n8623), .A3(n8622), .A4(n8621), .ZN(n8625)
         );
  NAND4_X1 U10192 ( .A1(n9262), .A2(n8626), .A3(n8625), .A4(n8709), .ZN(n8627)
         );
  NOR4_X1 U10193 ( .A1(n9226), .A2(n8628), .A3(n8708), .A4(n8627), .ZN(n8629)
         );
  NAND3_X1 U10194 ( .A1(n9197), .A2(n9207), .A3(n8629), .ZN(n8630) );
  NOR4_X1 U10195 ( .A1(n9157), .A2(n9173), .A3(n9186), .A4(n8630), .ZN(n8631)
         );
  NAND4_X1 U10196 ( .A1(n4955), .A2(n9132), .A3(n8631), .A4(n9119), .ZN(n8632)
         );
  NAND2_X1 U10197 ( .A1(n8761), .A2(n8762), .ZN(n9027) );
  XNOR2_X1 U10198 ( .A(n8633), .B(n7032), .ZN(n8634) );
  NAND2_X1 U10199 ( .A1(n8634), .A2(n8598), .ZN(n8792) );
  AND2_X1 U10200 ( .A1(n8635), .A2(n8651), .ZN(n8636) );
  NAND2_X1 U10201 ( .A1(n8648), .A2(n8637), .ZN(n8645) );
  INV_X1 U10202 ( .A(n8639), .ZN(n8640) );
  AOI21_X1 U10203 ( .B1(n8826), .B2(n8912), .A(n8640), .ZN(n8644) );
  NOR2_X1 U10204 ( .A1(n8641), .A2(n10229), .ZN(n8664) );
  INV_X1 U10205 ( .A(n8664), .ZN(n8642) );
  OAI211_X1 U10206 ( .C1(n8654), .C2(n8644), .A(n8643), .B(n8642), .ZN(n8668)
         );
  INV_X1 U10207 ( .A(n8645), .ZN(n8647) );
  AOI22_X1 U10208 ( .A1(n8654), .A2(n8648), .B1(n8647), .B2(n8646), .ZN(n8649)
         );
  OAI21_X1 U10209 ( .B1(n8649), .B2(n8670), .A(n8787), .ZN(n8666) );
  AOI21_X1 U10210 ( .B1(n8651), .B2(n8650), .A(n8612), .ZN(n8653) );
  NAND2_X1 U10211 ( .A1(n7272), .A2(n8661), .ZN(n8652) );
  OAI211_X1 U10212 ( .C1(n8653), .C2(n8652), .A(n8659), .B(n8787), .ZN(n8657)
         );
  INV_X1 U10213 ( .A(n8654), .ZN(n8656) );
  NAND3_X1 U10214 ( .A1(n8657), .A2(n8656), .A3(n8655), .ZN(n8665) );
  NAND3_X1 U10215 ( .A1(n8660), .A2(n8659), .A3(n8658), .ZN(n8662) );
  AND3_X1 U10216 ( .A1(n8662), .A2(n8771), .A3(n8661), .ZN(n8663) );
  AOI211_X1 U10217 ( .C1(n8666), .C2(n8665), .A(n8664), .B(n8663), .ZN(n8667)
         );
  AOI21_X1 U10218 ( .B1(n8771), .B2(n8668), .A(n8667), .ZN(n8669) );
  AOI21_X1 U10219 ( .B1(n8771), .B2(n8670), .A(n8669), .ZN(n8677) );
  NAND2_X1 U10220 ( .A1(n8671), .A2(n8771), .ZN(n8673) );
  NAND2_X1 U10221 ( .A1(n10239), .A2(n8787), .ZN(n8672) );
  MUX2_X1 U10222 ( .A(n8673), .B(n8672), .S(n8908), .Z(n8674) );
  OAI211_X1 U10223 ( .C1(n8677), .C2(n8676), .A(n8675), .B(n8674), .ZN(n8681)
         );
  MUX2_X1 U10224 ( .A(n8679), .B(n8678), .S(n8787), .Z(n8680) );
  NAND2_X1 U10225 ( .A1(n8681), .A2(n8680), .ZN(n8682) );
  NAND2_X1 U10226 ( .A1(n8682), .A2(n8683), .ZN(n8697) );
  INV_X1 U10227 ( .A(n8691), .ZN(n8685) );
  NAND2_X1 U10228 ( .A1(n8688), .A2(n8683), .ZN(n8684) );
  MUX2_X1 U10229 ( .A(n8685), .B(n8684), .S(n8787), .Z(n8687) );
  INV_X1 U10230 ( .A(n8689), .ZN(n8686) );
  OR2_X1 U10231 ( .A1(n8687), .A2(n8686), .ZN(n8692) );
  INV_X1 U10232 ( .A(n8692), .ZN(n8696) );
  NAND2_X1 U10233 ( .A1(n8700), .A2(n8688), .ZN(n8694) );
  OAI211_X1 U10234 ( .C1(n8692), .C2(n8691), .A(n8690), .B(n8689), .ZN(n8693)
         );
  MUX2_X1 U10235 ( .A(n8694), .B(n8693), .S(n8787), .Z(n8695) );
  INV_X1 U10236 ( .A(n8698), .ZN(n8699) );
  NAND2_X1 U10237 ( .A1(n8701), .A2(n8700), .ZN(n8703) );
  AND2_X1 U10238 ( .A1(n8704), .A2(n8771), .ZN(n8706) );
  NOR2_X1 U10239 ( .A1(n8704), .A2(n8771), .ZN(n8705) );
  MUX2_X1 U10240 ( .A(n8706), .B(n8705), .S(n8902), .Z(n8707) );
  NAND2_X1 U10241 ( .A1(n9265), .A2(n8771), .ZN(n8713) );
  NAND2_X1 U10242 ( .A1(n8710), .A2(n8787), .ZN(n8712) );
  MUX2_X1 U10243 ( .A(n8713), .B(n8712), .S(n8711), .Z(n8714) );
  NAND2_X1 U10244 ( .A1(n9262), .A2(n8714), .ZN(n8719) );
  MUX2_X1 U10245 ( .A(n8716), .B(n8715), .S(n8787), .Z(n8717) );
  OAI211_X1 U10246 ( .C1(n4528), .C2(n8719), .A(n8718), .B(n8717), .ZN(n8723)
         );
  INV_X1 U10247 ( .A(n9226), .ZN(n8722) );
  MUX2_X1 U10248 ( .A(n8720), .B(n9224), .S(n8787), .Z(n8721) );
  AND3_X1 U10249 ( .A1(n8723), .A2(n8722), .A3(n8721), .ZN(n8729) );
  INV_X1 U10250 ( .A(n8724), .ZN(n8727) );
  NAND2_X1 U10251 ( .A1(n8731), .A2(n8725), .ZN(n8726) );
  MUX2_X1 U10252 ( .A(n8727), .B(n8726), .S(n8787), .Z(n8728) );
  OR2_X1 U10253 ( .A1(n8729), .A2(n8728), .ZN(n8736) );
  INV_X1 U10254 ( .A(n8730), .ZN(n8738) );
  OAI211_X1 U10255 ( .C1(n8736), .C2(n8738), .A(n8737), .B(n8731), .ZN(n8732)
         );
  NAND2_X1 U10256 ( .A1(n8732), .A2(n8740), .ZN(n8734) );
  INV_X1 U10257 ( .A(n8741), .ZN(n8733) );
  NOR2_X1 U10258 ( .A1(n9017), .A2(n9016), .ZN(n8743) );
  INV_X1 U10259 ( .A(n8736), .ZN(n8739) );
  OAI21_X1 U10260 ( .B1(n8739), .B2(n8738), .A(n8737), .ZN(n8742) );
  NAND3_X1 U10261 ( .A1(n8742), .A2(n8741), .A3(n8740), .ZN(n8746) );
  INV_X1 U10262 ( .A(n8743), .ZN(n8744) );
  NAND3_X1 U10263 ( .A1(n8746), .A2(n8745), .A3(n8744), .ZN(n8748) );
  INV_X1 U10264 ( .A(n8747), .ZN(n9155) );
  NAND3_X1 U10265 ( .A1(n8748), .A2(n8750), .A3(n9155), .ZN(n8749) );
  MUX2_X1 U10266 ( .A(n8750), .B(n8749), .S(n8787), .Z(n8751) );
  NAND2_X1 U10267 ( .A1(n8751), .A2(n9132), .ZN(n8755) );
  MUX2_X1 U10268 ( .A(n8753), .B(n8752), .S(n8787), .Z(n8754) );
  NOR3_X1 U10269 ( .A1(n9117), .A2(n9136), .A3(n8787), .ZN(n8757) );
  NOR3_X1 U10270 ( .A1(n9304), .A2(n8847), .A3(n8771), .ZN(n8756) );
  NOR3_X1 U10271 ( .A1(n9098), .A2(n8757), .A3(n8756), .ZN(n8759) );
  AOI22_X1 U10272 ( .A1(n8760), .A2(n8759), .B1(n8771), .B2(n8758), .ZN(n8768)
         );
  MUX2_X1 U10273 ( .A(n8762), .B(n8761), .S(n8787), .Z(n8763) );
  NAND2_X1 U10274 ( .A1(n9064), .A2(n8763), .ZN(n8767) );
  AOI21_X1 U10275 ( .B1(n9087), .B2(n8764), .A(n8767), .ZN(n8765) );
  AOI211_X1 U10276 ( .C1(n9031), .C2(n9290), .A(n9057), .B(n8765), .ZN(n8766)
         );
  OAI22_X1 U10277 ( .A1(n8768), .A2(n8767), .B1(n8766), .B2(n8771), .ZN(n8769)
         );
  NAND2_X1 U10278 ( .A1(n8769), .A2(n8770), .ZN(n8777) );
  INV_X1 U10279 ( .A(n8770), .ZN(n8773) );
  OAI21_X1 U10280 ( .B1(n8773), .B2(n8772), .A(n8771), .ZN(n8776) );
  NOR3_X1 U10281 ( .A1(n9033), .A2(n9078), .A3(n8787), .ZN(n8775) );
  AOI211_X1 U10282 ( .C1(n8777), .C2(n8776), .A(n8775), .B(n9038), .ZN(n8786)
         );
  MUX2_X1 U10283 ( .A(n8779), .B(n8778), .S(n8787), .Z(n8781) );
  NAND3_X1 U10284 ( .A1(n8782), .A2(n8781), .A3(n8780), .ZN(n8785) );
  MUX2_X1 U10285 ( .A(n4518), .B(n8783), .S(n8787), .Z(n8784) );
  OAI21_X1 U10286 ( .B1(n8786), .B2(n8785), .A(n8784), .ZN(n8791) );
  MUX2_X1 U10287 ( .A(n4526), .B(n8788), .S(n8787), .Z(n8790) );
  AOI21_X1 U10288 ( .B1(n8791), .B2(n8790), .A(n8789), .ZN(n8797) );
  INV_X1 U10289 ( .A(n8793), .ZN(n8795) );
  NOR2_X1 U10290 ( .A1(n8795), .A2(n8794), .ZN(n8796) );
  NOR4_X1 U10291 ( .A1(n9233), .A2(n10200), .A3(n8799), .A4(n6974), .ZN(n8802)
         );
  OAI21_X1 U10292 ( .B1(n8803), .B2(n8800), .A(P2_B_REG_SCAN_IN), .ZN(n8801)
         );
  OAI22_X1 U10293 ( .A1(n8804), .A2(n8803), .B1(n8802), .B2(n8801), .ZN(
        P2_U3244) );
  OAI222_X1 U10294 ( .A1(P2_U3152), .A2(n8807), .B1(n4451), .B2(n8806), .C1(
        n8805), .C2(n9379), .ZN(P2_U3328) );
  INV_X1 U10295 ( .A(n6409), .ZN(n9838) );
  OAI222_X1 U10296 ( .A1(n8809), .A2(P2_U3152), .B1(n4451), .B2(n9838), .C1(
        n8808), .C2(n9379), .ZN(P2_U3330) );
  AOI22_X1 U10297 ( .A1(n8811), .A2(n8882), .B1(n8857), .B2(n9022), .ZN(n8817)
         );
  AND2_X2 U10298 ( .A1(n8811), .A2(n8810), .ZN(n8844) );
  INV_X1 U10299 ( .A(n8812), .ZN(n9129) );
  OAI22_X1 U10300 ( .A1(n8885), .A2(n9129), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8813), .ZN(n8815) );
  OAI22_X1 U10301 ( .A1(n8847), .A2(n8887), .B1(n8875), .B2(n9176), .ZN(n8814)
         );
  AOI211_X1 U10302 ( .C1(n9311), .C2(n8890), .A(n8815), .B(n8814), .ZN(n8816)
         );
  OAI21_X1 U10303 ( .B1(n8817), .B2(n8844), .A(n8816), .ZN(P2_U3218) );
  INV_X1 U10304 ( .A(n8818), .ZN(n8819) );
  AOI21_X1 U10305 ( .B1(n8820), .B2(n8819), .A(n8868), .ZN(n8825) );
  INV_X1 U10306 ( .A(n8821), .ZN(n8823) );
  NOR3_X1 U10307 ( .A1(n8892), .A2(n8823), .A3(n8822), .ZN(n8824) );
  OAI21_X1 U10308 ( .B1(n8825), .B2(n8824), .A(n7214), .ZN(n8831) );
  OAI22_X1 U10309 ( .A1(n8827), .A2(n8887), .B1(n8856), .B2(n8826), .ZN(n8828)
         );
  AOI21_X1 U10310 ( .B1(n8894), .B2(n7275), .A(n8828), .ZN(n8830) );
  MUX2_X1 U10311 ( .A(n8885), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n8829) );
  NAND3_X1 U10312 ( .A1(n8831), .A2(n8830), .A3(n8829), .ZN(P2_U3220) );
  INV_X1 U10313 ( .A(n8832), .ZN(n8833) );
  AOI21_X1 U10314 ( .B1(n6771), .B2(n8833), .A(n8868), .ZN(n8837) );
  NOR3_X1 U10315 ( .A1(n8834), .A2(n9175), .A3(n8892), .ZN(n8836) );
  OAI21_X1 U10316 ( .B1(n8837), .B2(n8836), .A(n8835), .ZN(n8842) );
  OAI22_X1 U10317 ( .A1(n8885), .A2(n9165), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8838), .ZN(n8840) );
  OAI22_X1 U10318 ( .A1(n9176), .A2(n8887), .B1(n8875), .B2(n9175), .ZN(n8839)
         );
  AOI211_X1 U10319 ( .C1(n9017), .C2(n8890), .A(n8840), .B(n8839), .ZN(n8841)
         );
  NAND2_X1 U10320 ( .A1(n8842), .A2(n8841), .ZN(P2_U3225) );
  NOR2_X1 U10321 ( .A1(n8844), .A2(n8843), .ZN(n8846) );
  XNOR2_X1 U10322 ( .A(n8846), .B(n8845), .ZN(n8850) );
  OAI22_X1 U10323 ( .A1(n8850), .A2(n8868), .B1(n8847), .B2(n8892), .ZN(n8848)
         );
  OAI21_X1 U10324 ( .B1(n8850), .B2(n8849), .A(n8848), .ZN(n8855) );
  NOR2_X1 U10325 ( .A1(n8885), .A2(n9114), .ZN(n8853) );
  OAI22_X1 U10326 ( .A1(n8851), .A2(n8887), .B1(n8875), .B2(n9021), .ZN(n8852)
         );
  AOI211_X1 U10327 ( .C1(P2_REG3_REG_24__SCAN_IN), .C2(P2_U3152), .A(n8853), 
        .B(n8852), .ZN(n8854) );
  OAI211_X1 U10328 ( .C1(n9117), .C2(n8856), .A(n8855), .B(n8854), .ZN(
        P2_U3231) );
  NAND2_X1 U10329 ( .A1(n8857), .A2(n8900), .ZN(n8861) );
  NAND2_X1 U10330 ( .A1(n8858), .A2(n8882), .ZN(n8860) );
  MUX2_X1 U10331 ( .A(n8861), .B(n8860), .S(n8859), .Z(n8866) );
  OAI22_X1 U10332 ( .A1(n8885), .A2(n9151), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8862), .ZN(n8864) );
  OAI22_X1 U10333 ( .A1(n9021), .A2(n8887), .B1(n8875), .B2(n9016), .ZN(n8863)
         );
  AOI211_X1 U10334 ( .C1(n9316), .C2(n8890), .A(n8864), .B(n8863), .ZN(n8865)
         );
  NAND2_X1 U10335 ( .A1(n8866), .A2(n8865), .ZN(P2_U3237) );
  INV_X1 U10336 ( .A(n8867), .ZN(n8869) );
  AOI21_X1 U10337 ( .B1(n6763), .B2(n8869), .A(n8868), .ZN(n8872) );
  NOR3_X1 U10338 ( .A1(n8870), .A2(n8874), .A3(n8892), .ZN(n8871) );
  OAI21_X1 U10339 ( .B1(n8872), .B2(n8871), .A(n8563), .ZN(n8879) );
  OAI22_X1 U10340 ( .A1(n8885), .A2(n9212), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8873), .ZN(n8877) );
  OAI22_X1 U10341 ( .A1(n9012), .A2(n8887), .B1(n8875), .B2(n8874), .ZN(n8876)
         );
  AOI211_X1 U10342 ( .C1(n9336), .C2(n8890), .A(n8877), .B(n8876), .ZN(n8878)
         );
  NAND2_X1 U10343 ( .A1(n8879), .A2(n8878), .ZN(P2_U3240) );
  OAI21_X1 U10344 ( .B1(n8893), .B2(n8881), .A(n8880), .ZN(n8883) );
  NAND2_X1 U10345 ( .A1(n8883), .A2(n8882), .ZN(n8898) );
  OAI22_X1 U10346 ( .A1(n8887), .A2(n8886), .B1(n8885), .B2(n8884), .ZN(n8888)
         );
  AOI211_X1 U10347 ( .C1(n10229), .C2(n8890), .A(n8889), .B(n8888), .ZN(n8897)
         );
  NOR3_X1 U10348 ( .A1(n8893), .A2(n8892), .A3(n8891), .ZN(n8895) );
  OAI21_X1 U10349 ( .B1(n8895), .B2(n8894), .A(n8910), .ZN(n8896) );
  NAND3_X1 U10350 ( .A1(n8898), .A2(n8897), .A3(n8896), .ZN(P2_U3241) );
  MUX2_X1 U10351 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n9039), .S(P2_U3966), .Z(
        P2_U3582) );
  INV_X1 U10352 ( .A(n8899), .ZN(n9058) );
  MUX2_X1 U10353 ( .A(n9058), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8913), .Z(
        P2_U3581) );
  MUX2_X1 U10354 ( .A(n9078), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8913), .Z(
        P2_U3580) );
  INV_X1 U10355 ( .A(n9031), .ZN(n9059) );
  MUX2_X1 U10356 ( .A(n9059), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8913), .Z(
        P2_U3579) );
  INV_X1 U10357 ( .A(n9072), .ZN(n9100) );
  MUX2_X1 U10358 ( .A(n9100), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8913), .Z(
        P2_U3578) );
  MUX2_X1 U10359 ( .A(n9120), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8913), .Z(
        P2_U3577) );
  MUX2_X1 U10360 ( .A(n9136), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8913), .Z(
        P2_U3576) );
  MUX2_X1 U10361 ( .A(n9022), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8913), .Z(
        P2_U3575) );
  MUX2_X1 U10362 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8900), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10363 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9187), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10364 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9015), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10365 ( .A(n9210), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8913), .Z(
        P2_U3571) );
  MUX2_X1 U10366 ( .A(n9008), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8913), .Z(
        P2_U3570) );
  MUX2_X1 U10367 ( .A(n9209), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8913), .Z(
        P2_U3569) );
  MUX2_X1 U10368 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9267), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10369 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8901), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10370 ( .A(n9265), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8913), .Z(
        P2_U3566) );
  MUX2_X1 U10371 ( .A(n8902), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8913), .Z(
        P2_U3565) );
  MUX2_X1 U10372 ( .A(n8903), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8913), .Z(
        P2_U3564) );
  MUX2_X1 U10373 ( .A(n8904), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8913), .Z(
        P2_U3563) );
  MUX2_X1 U10374 ( .A(n8905), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8913), .Z(
        P2_U3562) );
  MUX2_X1 U10375 ( .A(n8906), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8913), .Z(
        P2_U3561) );
  MUX2_X1 U10376 ( .A(n8907), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8913), .Z(
        P2_U3560) );
  MUX2_X1 U10377 ( .A(n8908), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8913), .Z(
        P2_U3559) );
  MUX2_X1 U10378 ( .A(n8909), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8913), .Z(
        P2_U3558) );
  MUX2_X1 U10379 ( .A(n8910), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8913), .Z(
        P2_U3557) );
  MUX2_X1 U10380 ( .A(n8911), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8913), .Z(
        P2_U3556) );
  MUX2_X1 U10381 ( .A(n8912), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8913), .Z(
        P2_U3555) );
  MUX2_X1 U10382 ( .A(n7275), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8913), .Z(
        P2_U3554) );
  MUX2_X1 U10383 ( .A(n7025), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8913), .Z(
        P2_U3553) );
  MUX2_X1 U10384 ( .A(n6954), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8913), .Z(
        P2_U3552) );
  OAI211_X1 U10385 ( .C1(n8916), .C2(n8915), .A(n10177), .B(n8914), .ZN(n8925)
         );
  NOR2_X1 U10386 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5154), .ZN(n8917) );
  AOI21_X1 U10387 ( .B1(n10176), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8917), .ZN(
        n8924) );
  NAND2_X1 U10388 ( .A1(n9860), .A2(n8918), .ZN(n8923) );
  OAI211_X1 U10389 ( .C1(n8921), .C2(n8920), .A(n10174), .B(n8919), .ZN(n8922)
         );
  NAND4_X1 U10390 ( .A1(n8925), .A2(n8924), .A3(n8923), .A4(n8922), .ZN(
        P2_U3250) );
  NOR2_X1 U10391 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8926), .ZN(n8929) );
  NOR2_X1 U10392 ( .A1(n10178), .A2(n8927), .ZN(n8928) );
  AOI211_X1 U10393 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n10176), .A(n8929), .B(
        n8928), .ZN(n8938) );
  OAI211_X1 U10394 ( .C1(n8932), .C2(n8931), .A(n10174), .B(n8930), .ZN(n8937)
         );
  OAI211_X1 U10395 ( .C1(n8935), .C2(n8934), .A(n10177), .B(n8933), .ZN(n8936)
         );
  NAND3_X1 U10396 ( .A1(n8938), .A2(n8937), .A3(n8936), .ZN(P2_U3253) );
  INV_X1 U10397 ( .A(n8939), .ZN(n8942) );
  NOR2_X1 U10398 ( .A1(n10178), .A2(n8940), .ZN(n8941) );
  AOI211_X1 U10399 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n10176), .A(n8942), .B(
        n8941), .ZN(n8951) );
  OAI211_X1 U10400 ( .C1(n8945), .C2(n8944), .A(n8943), .B(n10174), .ZN(n8950)
         );
  OAI211_X1 U10401 ( .C1(n8948), .C2(n8947), .A(n8946), .B(n10177), .ZN(n8949)
         );
  NAND3_X1 U10402 ( .A1(n8951), .A2(n8950), .A3(n8949), .ZN(P2_U3255) );
  OAI211_X1 U10403 ( .C1(n8954), .C2(n8953), .A(n10177), .B(n8952), .ZN(n8965)
         );
  NOR2_X1 U10404 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8955), .ZN(n8956) );
  AOI21_X1 U10405 ( .B1(n10176), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8956), .ZN(
        n8964) );
  OAI21_X1 U10406 ( .B1(n8959), .B2(n8958), .A(n8957), .ZN(n8960) );
  NAND2_X1 U10407 ( .A1(n8960), .A2(n10174), .ZN(n8963) );
  NAND2_X1 U10408 ( .A1(n9860), .A2(n8961), .ZN(n8962) );
  NAND4_X1 U10409 ( .A1(n8965), .A2(n8964), .A3(n8963), .A4(n8962), .ZN(
        P2_U3261) );
  OAI211_X1 U10410 ( .C1(n8968), .C2(n8967), .A(n10177), .B(n8966), .ZN(n8979)
         );
  NOR2_X1 U10411 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8969), .ZN(n8970) );
  AOI21_X1 U10412 ( .B1(n10176), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8970), .ZN(
        n8978) );
  NAND2_X1 U10413 ( .A1(n9860), .A2(n8971), .ZN(n8977) );
  AOI21_X1 U10414 ( .B1(n8974), .B2(n8973), .A(n8972), .ZN(n8975) );
  NAND2_X1 U10415 ( .A1(n10174), .A2(n8975), .ZN(n8976) );
  NAND4_X1 U10416 ( .A1(n8979), .A2(n8978), .A3(n8977), .A4(n8976), .ZN(
        P2_U3262) );
  INV_X1 U10417 ( .A(n8980), .ZN(n8981) );
  NAND2_X1 U10418 ( .A1(n8981), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8984) );
  NAND2_X1 U10419 ( .A1(n8982), .A2(n8987), .ZN(n8983) );
  NAND2_X1 U10420 ( .A1(n8984), .A2(n8983), .ZN(n8985) );
  XOR2_X1 U10421 ( .A(n8985), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8991) );
  OAI21_X1 U10422 ( .B1(n8987), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8986), .ZN(
        n8988) );
  XOR2_X1 U10423 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8988), .Z(n8993) );
  INV_X1 U10424 ( .A(n8993), .ZN(n8989) );
  AOI22_X1 U10425 ( .A1(n8991), .A2(n10177), .B1(n8989), .B2(n10174), .ZN(
        n8995) );
  NOR2_X1 U10426 ( .A1(n8991), .A2(n8990), .ZN(n8992) );
  AOI211_X1 U10427 ( .C1(n10174), .C2(n8993), .A(n9860), .B(n8992), .ZN(n8994)
         );
  MUX2_X1 U10428 ( .A(n8995), .B(n8994), .S(n4455), .Z(n8997) );
  NAND2_X1 U10429 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8996) );
  OAI211_X1 U10430 ( .C1(n8999), .C2(n8998), .A(n8997), .B(n8996), .ZN(
        P2_U3264) );
  AOI21_X1 U10431 ( .B1(n9043), .B2(n9001), .A(n9000), .ZN(n9882) );
  NAND2_X1 U10432 ( .A1(n9882), .A2(n9272), .ZN(n9004) );
  AOI21_X1 U10433 ( .B1(n10198), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9002), .ZN(
        n9003) );
  OAI211_X1 U10434 ( .C1(n9880), .C2(n9260), .A(n9004), .B(n9003), .ZN(
        P2_U3266) );
  NAND2_X1 U10435 ( .A1(n9006), .A2(n8874), .ZN(n9007) );
  NAND2_X1 U10436 ( .A1(n9336), .A2(n9008), .ZN(n9010) );
  NAND2_X1 U10437 ( .A1(n9192), .A2(n9011), .ZN(n9014) );
  NAND2_X1 U10438 ( .A1(n9164), .A2(n9016), .ZN(n9019) );
  NAND2_X1 U10439 ( .A1(n9311), .A2(n9022), .ZN(n9023) );
  NAND2_X1 U10440 ( .A1(n9096), .A2(n9098), .ZN(n9026) );
  INV_X1 U10441 ( .A(n9295), .ZN(n9028) );
  NAND2_X1 U10442 ( .A1(n9028), .A2(n9072), .ZN(n9029) );
  NAND2_X1 U10443 ( .A1(n9071), .A2(n9031), .ZN(n9032) );
  NAND2_X1 U10444 ( .A1(n9033), .A2(n8774), .ZN(n9034) );
  NAND2_X1 U10445 ( .A1(n9035), .A2(n9034), .ZN(n9036) );
  XNOR2_X1 U10446 ( .A(n9036), .B(n9038), .ZN(n9278) );
  INV_X1 U10447 ( .A(n9278), .ZN(n9051) );
  XOR2_X1 U10448 ( .A(n9038), .B(n9037), .Z(n9042) );
  AOI22_X1 U10449 ( .A1(n9078), .A2(n9264), .B1(n9040), .B2(n9039), .ZN(n9041)
         );
  OAI21_X1 U10450 ( .B1(n9042), .B2(n9228), .A(n9041), .ZN(n9282) );
  OAI21_X1 U10451 ( .B1(n9054), .B2(n9279), .A(n9043), .ZN(n9280) );
  OAI22_X1 U10452 ( .A1(n9045), .A2(n9241), .B1(n9044), .B2(n9238), .ZN(n9046)
         );
  AOI21_X1 U10453 ( .B1(n9047), .B2(n9246), .A(n9046), .ZN(n9048) );
  OAI21_X1 U10454 ( .B1(n9280), .B2(n9218), .A(n9048), .ZN(n9049) );
  AOI21_X1 U10455 ( .B1(n9282), .B2(n9238), .A(n9049), .ZN(n9050) );
  OAI21_X1 U10456 ( .B1(n9051), .B2(n9274), .A(n9050), .ZN(P2_U3267) );
  INV_X1 U10457 ( .A(n9057), .ZN(n9052) );
  AOI21_X1 U10458 ( .B1(n8596), .B2(n9065), .A(n9054), .ZN(n9285) );
  INV_X1 U10459 ( .A(n9241), .ZN(n10189) );
  AOI22_X1 U10460 ( .A1(n9055), .A2(n10189), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n10198), .ZN(n9056) );
  OAI21_X1 U10461 ( .B1(n9033), .B2(n9260), .A(n9056), .ZN(n9061) );
  AOI211_X1 U10462 ( .C1(n9272), .C2(n9285), .A(n9061), .B(n9060), .ZN(n9062)
         );
  OAI21_X1 U10463 ( .B1(n9288), .B2(n9274), .A(n9062), .ZN(P2_U3268) );
  XNOR2_X1 U10464 ( .A(n9063), .B(n9064), .ZN(n9293) );
  INV_X1 U10465 ( .A(n9091), .ZN(n9067) );
  INV_X1 U10466 ( .A(n9065), .ZN(n9066) );
  AOI211_X1 U10467 ( .C1(n9290), .C2(n9067), .A(n10273), .B(n9066), .ZN(n9289)
         );
  INV_X1 U10468 ( .A(n9068), .ZN(n9069) );
  AOI22_X1 U10469 ( .A1(n9069), .A2(n10189), .B1(n10198), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n9070) );
  OAI21_X1 U10470 ( .B1(n9071), .B2(n9260), .A(n9070), .ZN(n9080) );
  NOR2_X1 U10471 ( .A1(n9072), .A2(n9233), .ZN(n9077) );
  AOI211_X1 U10472 ( .C1(n9075), .C2(n9074), .A(n9228), .B(n9073), .ZN(n9076)
         );
  AOI211_X1 U10473 ( .C1(n9266), .C2(n9078), .A(n9077), .B(n9076), .ZN(n9292)
         );
  NOR2_X1 U10474 ( .A1(n9292), .A2(n10198), .ZN(n9079) );
  AOI211_X1 U10475 ( .C1(n9169), .C2(n9289), .A(n9080), .B(n9079), .ZN(n9081)
         );
  OAI21_X1 U10476 ( .B1(n9293), .B2(n9274), .A(n9081), .ZN(P2_U3269) );
  XNOR2_X1 U10477 ( .A(n9082), .B(n9087), .ZN(n9298) );
  OAI22_X1 U10478 ( .A1(n9084), .A2(n9241), .B1(n9238), .B2(n9083), .ZN(n9094)
         );
  INV_X1 U10479 ( .A(n9085), .ZN(n9086) );
  NOR2_X1 U10480 ( .A1(n9103), .A2(n9086), .ZN(n9088) );
  XNOR2_X1 U10481 ( .A(n9088), .B(n9087), .ZN(n9090) );
  AOI21_X1 U10482 ( .B1(n9090), .B2(n9269), .A(n9089), .ZN(n9297) );
  AOI211_X1 U10483 ( .C1(n9295), .C2(n9104), .A(n10273), .B(n9091), .ZN(n9294)
         );
  NAND2_X1 U10484 ( .A1(n9294), .A2(n7032), .ZN(n9092) );
  AOI21_X1 U10485 ( .B1(n9297), .B2(n9092), .A(n10198), .ZN(n9093) );
  AOI211_X1 U10486 ( .C1(n9246), .C2(n9295), .A(n9094), .B(n9093), .ZN(n9095)
         );
  OAI21_X1 U10487 ( .B1(n9298), .B2(n9274), .A(n9095), .ZN(P2_U3270) );
  XNOR2_X1 U10488 ( .A(n9096), .B(n4955), .ZN(n9303) );
  AOI22_X1 U10489 ( .A1(n9301), .A2(n9246), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n10198), .ZN(n9110) );
  NAND3_X1 U10490 ( .A1(n9118), .A2(n9098), .A3(n9097), .ZN(n9099) );
  NAND2_X1 U10491 ( .A1(n9099), .A2(n9269), .ZN(n9102) );
  AOI22_X1 U10492 ( .A1(n9100), .A2(n9266), .B1(n9264), .B2(n9136), .ZN(n9101)
         );
  OAI21_X1 U10493 ( .B1(n9103), .B2(n9102), .A(n9101), .ZN(n9299) );
  INV_X1 U10494 ( .A(n9104), .ZN(n9105) );
  AOI211_X1 U10495 ( .C1(n9301), .C2(n4534), .A(n10273), .B(n9105), .ZN(n9300)
         );
  INV_X1 U10496 ( .A(n9300), .ZN(n9107) );
  OAI22_X1 U10497 ( .A1(n9107), .A2(n4455), .B1(n9106), .B2(n9241), .ZN(n9108)
         );
  OAI21_X1 U10498 ( .B1(n9299), .B2(n9108), .A(n9238), .ZN(n9109) );
  OAI211_X1 U10499 ( .C1(n9303), .C2(n9274), .A(n9110), .B(n9109), .ZN(
        P2_U3271) );
  INV_X1 U10500 ( .A(n9111), .ZN(n9112) );
  AOI21_X1 U10501 ( .B1(n9119), .B2(n9113), .A(n9112), .ZN(n9308) );
  XNOR2_X1 U10502 ( .A(n9141), .B(n9117), .ZN(n9305) );
  INV_X1 U10503 ( .A(n9114), .ZN(n9115) );
  AOI22_X1 U10504 ( .A1(n10198), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9115), 
        .B2(n10189), .ZN(n9116) );
  OAI21_X1 U10505 ( .B1(n9117), .B2(n9260), .A(n9116), .ZN(n9124) );
  OAI211_X1 U10506 ( .C1(n4522), .C2(n9119), .A(n9118), .B(n9269), .ZN(n9122)
         );
  AOI22_X1 U10507 ( .A1(n9120), .A2(n9266), .B1(n9264), .B2(n9022), .ZN(n9121)
         );
  AND2_X1 U10508 ( .A1(n9122), .A2(n9121), .ZN(n9307) );
  NOR2_X1 U10509 ( .A1(n9307), .A2(n10198), .ZN(n9123) );
  AOI211_X1 U10510 ( .C1(n9305), .C2(n9272), .A(n9124), .B(n9123), .ZN(n9125)
         );
  OAI21_X1 U10511 ( .B1(n9308), .B2(n9274), .A(n9125), .ZN(P2_U3272) );
  OR2_X1 U10512 ( .A1(n9127), .A2(n9126), .ZN(n9310) );
  INV_X1 U10513 ( .A(n9274), .ZN(n9128) );
  NAND3_X1 U10514 ( .A1(n9310), .A2(n9309), .A3(n9128), .ZN(n9145) );
  INV_X1 U10515 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9130) );
  OAI22_X1 U10516 ( .A1(n9244), .A2(n9130), .B1(n9129), .B2(n9241), .ZN(n9131)
         );
  AOI21_X1 U10517 ( .B1(n9311), .B2(n9246), .A(n9131), .ZN(n9144) );
  NOR2_X1 U10518 ( .A1(n9133), .A2(n9132), .ZN(n9134) );
  OR2_X1 U10519 ( .A1(n9135), .A2(n9134), .ZN(n9139) );
  NAND2_X1 U10520 ( .A1(n9136), .A2(n9266), .ZN(n9137) );
  OAI21_X1 U10521 ( .B1(n9176), .B2(n9233), .A(n9137), .ZN(n9138) );
  AOI21_X1 U10522 ( .B1(n9139), .B2(n9269), .A(n9138), .ZN(n9314) );
  OR2_X1 U10523 ( .A1(n9314), .A2(n10198), .ZN(n9143) );
  NAND2_X1 U10524 ( .A1(n9148), .A2(n9311), .ZN(n9140) );
  AND2_X1 U10525 ( .A1(n9141), .A2(n9140), .ZN(n9312) );
  NAND2_X1 U10526 ( .A1(n9312), .A2(n9272), .ZN(n9142) );
  NAND4_X1 U10527 ( .A1(n9145), .A2(n9144), .A3(n9143), .A4(n9142), .ZN(
        P2_U3273) );
  XOR2_X1 U10528 ( .A(n9146), .B(n9157), .Z(n9320) );
  INV_X1 U10529 ( .A(n9147), .ZN(n9150) );
  INV_X1 U10530 ( .A(n9148), .ZN(n9149) );
  AOI21_X1 U10531 ( .B1(n9316), .B2(n9150), .A(n9149), .ZN(n9317) );
  INV_X1 U10532 ( .A(n9151), .ZN(n9152) );
  AOI22_X1 U10533 ( .A1(n10198), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9152), 
        .B2(n10189), .ZN(n9153) );
  OAI21_X1 U10534 ( .B1(n9154), .B2(n9260), .A(n9153), .ZN(n9160) );
  NAND2_X1 U10535 ( .A1(n9170), .A2(n9155), .ZN(n9156) );
  XOR2_X1 U10536 ( .A(n9157), .B(n9156), .Z(n9158) );
  AOI222_X1 U10537 ( .A1(n9269), .A2(n9158), .B1(n9187), .B2(n9264), .C1(n9022), .C2(n9266), .ZN(n9319) );
  NOR2_X1 U10538 ( .A1(n9319), .A2(n10198), .ZN(n9159) );
  AOI211_X1 U10539 ( .C1(n9317), .C2(n9272), .A(n9160), .B(n9159), .ZN(n9161)
         );
  OAI21_X1 U10540 ( .B1(n9320), .B2(n9274), .A(n9161), .ZN(P2_U3274) );
  XOR2_X1 U10541 ( .A(n9162), .B(n9173), .Z(n9324) );
  XNOR2_X1 U10542 ( .A(n9180), .B(n9017), .ZN(n9163) );
  NOR2_X1 U10543 ( .A1(n9163), .A2(n10273), .ZN(n9322) );
  NOR2_X1 U10544 ( .A1(n9164), .A2(n9260), .ZN(n9168) );
  OAI22_X1 U10545 ( .A1(n9244), .A2(n9166), .B1(n9165), .B2(n9241), .ZN(n9167)
         );
  AOI211_X1 U10546 ( .C1(n9322), .C2(n9169), .A(n9168), .B(n9167), .ZN(n9178)
         );
  INV_X1 U10547 ( .A(n9170), .ZN(n9171) );
  AOI21_X1 U10548 ( .B1(n9173), .B2(n9172), .A(n9171), .ZN(n9174) );
  OAI222_X1 U10549 ( .A1(n9231), .A2(n9176), .B1(n9233), .B2(n9175), .C1(n9228), .C2(n9174), .ZN(n9321) );
  NAND2_X1 U10550 ( .A1(n9321), .A2(n9238), .ZN(n9177) );
  OAI211_X1 U10551 ( .C1(n9324), .C2(n9274), .A(n9178), .B(n9177), .ZN(
        P2_U3275) );
  XNOR2_X1 U10552 ( .A(n9179), .B(n9186), .ZN(n9329) );
  AOI21_X1 U10553 ( .B1(n9325), .B2(n9195), .A(n4609), .ZN(n9326) );
  INV_X1 U10554 ( .A(n9181), .ZN(n9182) );
  AOI22_X1 U10555 ( .A1(n10198), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9182), 
        .B2(n10189), .ZN(n9183) );
  OAI21_X1 U10556 ( .B1(n9184), .B2(n9260), .A(n9183), .ZN(n9190) );
  XOR2_X1 U10557 ( .A(n9186), .B(n9185), .Z(n9188) );
  AOI222_X1 U10558 ( .A1(n9269), .A2(n9188), .B1(n9210), .B2(n9264), .C1(n9187), .C2(n9266), .ZN(n9328) );
  NOR2_X1 U10559 ( .A1(n9328), .A2(n10198), .ZN(n9189) );
  AOI211_X1 U10560 ( .C1(n9326), .C2(n9272), .A(n9190), .B(n9189), .ZN(n9191)
         );
  OAI21_X1 U10561 ( .B1(n9329), .B2(n9274), .A(n9191), .ZN(P2_U3276) );
  XOR2_X1 U10562 ( .A(n9192), .B(n9197), .Z(n9334) );
  INV_X1 U10563 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9194) );
  OAI22_X1 U10564 ( .A1(n9238), .A2(n9194), .B1(n9193), .B2(n9241), .ZN(n9203)
         );
  INV_X1 U10565 ( .A(n9216), .ZN(n9196) );
  AOI211_X1 U10566 ( .C1(n9332), .C2(n9196), .A(n10273), .B(n4610), .ZN(n9331)
         );
  XOR2_X1 U10567 ( .A(n9198), .B(n9197), .Z(n9200) );
  OAI21_X1 U10568 ( .B1(n9200), .B2(n9228), .A(n9199), .ZN(n9330) );
  AOI21_X1 U10569 ( .B1(n9331), .B2(n7032), .A(n9330), .ZN(n9201) );
  NOR2_X1 U10570 ( .A1(n9201), .A2(n10198), .ZN(n9202) );
  AOI211_X1 U10571 ( .C1(n9246), .C2(n9332), .A(n9203), .B(n9202), .ZN(n9204)
         );
  OAI21_X1 U10572 ( .B1(n9334), .B2(n9274), .A(n9204), .ZN(P2_U3277) );
  XNOR2_X1 U10573 ( .A(n9205), .B(n9207), .ZN(n9340) );
  OAI21_X1 U10574 ( .B1(n9208), .B2(n9207), .A(n9206), .ZN(n9211) );
  AOI222_X1 U10575 ( .A1(n9269), .A2(n9211), .B1(n9210), .B2(n9266), .C1(n9209), .C2(n9264), .ZN(n9339) );
  OAI21_X1 U10576 ( .B1(n9212), .B2(n9241), .A(n9339), .ZN(n9220) );
  NOR2_X1 U10577 ( .A1(n9214), .A2(n9213), .ZN(n9215) );
  OR2_X1 U10578 ( .A1(n9216), .A2(n9215), .ZN(n9335) );
  AOI22_X1 U10579 ( .A1(n9336), .A2(n9246), .B1(n10198), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n9217) );
  OAI21_X1 U10580 ( .B1(n9335), .B2(n9218), .A(n9217), .ZN(n9219) );
  AOI21_X1 U10581 ( .B1(n9220), .B2(n9238), .A(n9219), .ZN(n9221) );
  OAI21_X1 U10582 ( .B1(n9340), .B2(n9274), .A(n9221), .ZN(P2_U3278) );
  OAI21_X1 U10583 ( .B1(n9223), .B2(n9226), .A(n9222), .ZN(n9341) );
  INV_X1 U10584 ( .A(n9341), .ZN(n9251) );
  NAND2_X1 U10585 ( .A1(n9225), .A2(n9224), .ZN(n9227) );
  XNOR2_X1 U10586 ( .A(n9227), .B(n9226), .ZN(n9229) );
  OAI222_X1 U10587 ( .A1(n9233), .A2(n9232), .B1(n9231), .B2(n9230), .C1(n9229), .C2(n9228), .ZN(n9240) );
  INV_X1 U10588 ( .A(n9234), .ZN(n9237) );
  XOR2_X1 U10589 ( .A(n9247), .B(n9235), .Z(n9236) );
  AOI21_X1 U10590 ( .B1(n10231), .B2(n9236), .A(n9240), .ZN(n9342) );
  OAI21_X1 U10591 ( .B1(n9251), .B2(n9237), .A(n9342), .ZN(n9239) );
  OAI211_X1 U10592 ( .C1(n7032), .C2(n9240), .A(n9239), .B(n9238), .ZN(n9249)
         );
  OAI22_X1 U10593 ( .A1(n9244), .A2(n9243), .B1(n9242), .B2(n9241), .ZN(n9245)
         );
  AOI21_X1 U10594 ( .B1(n9247), .B2(n9246), .A(n9245), .ZN(n9248) );
  OAI211_X1 U10595 ( .C1(n9251), .C2(n9250), .A(n9249), .B(n9248), .ZN(
        P2_U3279) );
  XOR2_X1 U10596 ( .A(n9262), .B(n9252), .Z(n9354) );
  INV_X1 U10597 ( .A(n9253), .ZN(n9256) );
  INV_X1 U10598 ( .A(n9254), .ZN(n9255) );
  AOI21_X1 U10599 ( .B1(n9350), .B2(n9256), .A(n9255), .ZN(n9351) );
  INV_X1 U10600 ( .A(n9257), .ZN(n9258) );
  AOI22_X1 U10601 ( .A1(n10198), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9258), 
        .B2(n10189), .ZN(n9259) );
  OAI21_X1 U10602 ( .B1(n9261), .B2(n9260), .A(n9259), .ZN(n9271) );
  XOR2_X1 U10603 ( .A(n9263), .B(n9262), .Z(n9268) );
  AOI222_X1 U10604 ( .A1(n9269), .A2(n9268), .B1(n9267), .B2(n9266), .C1(n9265), .C2(n9264), .ZN(n9353) );
  NOR2_X1 U10605 ( .A1(n9353), .A2(n10198), .ZN(n9270) );
  AOI211_X1 U10606 ( .C1(n9351), .C2(n9272), .A(n9271), .B(n9270), .ZN(n9273)
         );
  OAI21_X1 U10607 ( .B1(n9354), .B2(n9274), .A(n9273), .ZN(P2_U3281) );
  NAND2_X1 U10608 ( .A1(n9275), .A2(n10230), .ZN(n9276) );
  OAI211_X1 U10609 ( .C1(n9277), .C2(n10273), .A(n9879), .B(n9276), .ZN(n9355)
         );
  MUX2_X1 U10610 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9355), .S(n4449), .Z(
        P2_U3551) );
  NAND2_X1 U10611 ( .A1(n9278), .A2(n10278), .ZN(n9284) );
  OAI22_X1 U10612 ( .A1(n9280), .A2(n10273), .B1(n9279), .B2(n10272), .ZN(
        n9281) );
  NOR2_X1 U10613 ( .A1(n9282), .A2(n9281), .ZN(n9283) );
  NAND2_X1 U10614 ( .A1(n9284), .A2(n9283), .ZN(n9356) );
  MUX2_X1 U10615 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9356), .S(n4449), .Z(
        P2_U3549) );
  AOI22_X1 U10616 ( .A1(n9285), .A2(n10231), .B1(n10230), .B2(n8596), .ZN(
        n9286) );
  OAI211_X1 U10617 ( .C1(n9288), .C2(n10235), .A(n9287), .B(n9286), .ZN(n9357)
         );
  MUX2_X1 U10618 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9357), .S(n4449), .Z(
        P2_U3548) );
  AOI21_X1 U10619 ( .B1(n10230), .B2(n9290), .A(n9289), .ZN(n9291) );
  OAI211_X1 U10620 ( .C1(n9293), .C2(n10235), .A(n9292), .B(n9291), .ZN(n9358)
         );
  MUX2_X1 U10621 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9358), .S(n4449), .Z(
        P2_U3547) );
  AOI21_X1 U10622 ( .B1(n10230), .B2(n9295), .A(n9294), .ZN(n9296) );
  OAI211_X1 U10623 ( .C1(n9298), .C2(n10235), .A(n9297), .B(n9296), .ZN(n9359)
         );
  MUX2_X1 U10624 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9359), .S(n4449), .Z(
        P2_U3546) );
  AOI211_X1 U10625 ( .C1(n10230), .C2(n9301), .A(n9300), .B(n9299), .ZN(n9302)
         );
  OAI21_X1 U10626 ( .B1(n9303), .B2(n10235), .A(n9302), .ZN(n9360) );
  MUX2_X1 U10627 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9360), .S(n4449), .Z(
        P2_U3545) );
  AOI22_X1 U10628 ( .A1(n9305), .A2(n10231), .B1(n10230), .B2(n9304), .ZN(
        n9306) );
  OAI211_X1 U10629 ( .C1(n9308), .C2(n10235), .A(n9307), .B(n9306), .ZN(n9361)
         );
  MUX2_X1 U10630 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9361), .S(n4449), .Z(
        P2_U3544) );
  NAND3_X1 U10631 ( .A1(n9310), .A2(n9309), .A3(n10278), .ZN(n9315) );
  AOI22_X1 U10632 ( .A1(n9312), .A2(n10231), .B1(n10230), .B2(n9311), .ZN(
        n9313) );
  NAND3_X1 U10633 ( .A1(n9315), .A2(n9314), .A3(n9313), .ZN(n9362) );
  MUX2_X1 U10634 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9362), .S(n4449), .Z(
        P2_U3543) );
  AOI22_X1 U10635 ( .A1(n9317), .A2(n10231), .B1(n10230), .B2(n9316), .ZN(
        n9318) );
  OAI211_X1 U10636 ( .C1(n9320), .C2(n10235), .A(n9319), .B(n9318), .ZN(n9363)
         );
  MUX2_X1 U10637 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9363), .S(n4449), .Z(
        P2_U3542) );
  AOI211_X1 U10638 ( .C1(n10230), .C2(n9017), .A(n9322), .B(n9321), .ZN(n9323)
         );
  OAI21_X1 U10639 ( .B1(n9324), .B2(n10235), .A(n9323), .ZN(n9364) );
  MUX2_X1 U10640 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9364), .S(n4449), .Z(
        P2_U3541) );
  AOI22_X1 U10641 ( .A1(n9326), .A2(n10231), .B1(n10230), .B2(n9325), .ZN(
        n9327) );
  OAI211_X1 U10642 ( .C1(n9329), .C2(n10235), .A(n9328), .B(n9327), .ZN(n9365)
         );
  MUX2_X1 U10643 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9365), .S(n4449), .Z(
        P2_U3540) );
  AOI211_X1 U10644 ( .C1(n10230), .C2(n9332), .A(n9331), .B(n9330), .ZN(n9333)
         );
  OAI21_X1 U10645 ( .B1(n9334), .B2(n10235), .A(n9333), .ZN(n9366) );
  MUX2_X1 U10646 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9366), .S(n4449), .Z(
        P2_U3539) );
  INV_X1 U10647 ( .A(n9335), .ZN(n9337) );
  AOI22_X1 U10648 ( .A1(n9337), .A2(n10231), .B1(n10230), .B2(n9336), .ZN(
        n9338) );
  OAI211_X1 U10649 ( .C1(n9340), .C2(n10235), .A(n9339), .B(n9338), .ZN(n9367)
         );
  MUX2_X1 U10650 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9367), .S(n4449), .Z(
        P2_U3538) );
  NAND2_X1 U10651 ( .A1(n9341), .A2(n10278), .ZN(n9343) );
  OAI211_X1 U10652 ( .C1(n9006), .C2(n10272), .A(n9343), .B(n9342), .ZN(n9368)
         );
  MUX2_X1 U10653 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9368), .S(n4449), .Z(
        P2_U3537) );
  INV_X1 U10654 ( .A(n9344), .ZN(n9349) );
  AOI22_X1 U10655 ( .A1(n9346), .A2(n10231), .B1(n10230), .B2(n9345), .ZN(
        n9347) );
  OAI211_X1 U10656 ( .C1(n9349), .C2(n10235), .A(n9348), .B(n9347), .ZN(n9369)
         );
  MUX2_X1 U10657 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9369), .S(n4449), .Z(
        P2_U3536) );
  AOI22_X1 U10658 ( .A1(n9351), .A2(n10231), .B1(n10230), .B2(n9350), .ZN(
        n9352) );
  OAI211_X1 U10659 ( .C1(n9354), .C2(n10235), .A(n9353), .B(n9352), .ZN(n9370)
         );
  MUX2_X1 U10660 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9370), .S(n4449), .Z(
        P2_U3535) );
  MUX2_X1 U10661 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9355), .S(n10281), .Z(
        P2_U3519) );
  MUX2_X1 U10662 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9356), .S(n10281), .Z(
        P2_U3517) );
  MUX2_X1 U10663 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9357), .S(n10281), .Z(
        P2_U3516) );
  MUX2_X1 U10664 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9358), .S(n10281), .Z(
        P2_U3515) );
  MUX2_X1 U10665 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9359), .S(n10281), .Z(
        P2_U3514) );
  MUX2_X1 U10666 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9360), .S(n10281), .Z(
        P2_U3513) );
  MUX2_X1 U10667 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9361), .S(n10281), .Z(
        P2_U3512) );
  MUX2_X1 U10668 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9362), .S(n10281), .Z(
        P2_U3511) );
  MUX2_X1 U10669 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9363), .S(n10281), .Z(
        P2_U3510) );
  MUX2_X1 U10670 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9364), .S(n10281), .Z(
        P2_U3509) );
  MUX2_X1 U10671 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9365), .S(n10281), .Z(
        P2_U3508) );
  MUX2_X1 U10672 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9366), .S(n10281), .Z(
        P2_U3507) );
  MUX2_X1 U10673 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9367), .S(n10281), .Z(
        P2_U3505) );
  MUX2_X1 U10674 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9368), .S(n10281), .Z(
        P2_U3502) );
  MUX2_X1 U10675 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9369), .S(n10281), .Z(
        P2_U3499) );
  MUX2_X1 U10676 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9370), .S(n10281), .Z(
        P2_U3496) );
  INV_X1 U10677 ( .A(n9371), .ZN(n9830) );
  INV_X1 U10678 ( .A(n9372), .ZN(n9373) );
  NOR4_X1 U10679 ( .A1(n9373), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9374), .A4(
        P2_U3152), .ZN(n9375) );
  AOI21_X1 U10680 ( .B1(n9376), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9375), .ZN(
        n9377) );
  OAI21_X1 U10681 ( .B1(n9830), .B2(n4451), .A(n9377), .ZN(P2_U3327) );
  INV_X1 U10682 ( .A(n9378), .ZN(n9834) );
  OAI222_X1 U10683 ( .A1(n5042), .A2(P2_U3152), .B1(n4451), .B2(n9834), .C1(
        n9380), .C2(n9379), .ZN(P2_U3329) );
  MUX2_X1 U10684 ( .A(n9381), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  AOI21_X1 U10685 ( .B1(n9384), .B2(n9383), .A(n9382), .ZN(n9385) );
  NOR2_X1 U10686 ( .A1(n9455), .A2(n9634), .ZN(n9388) );
  OAI22_X1 U10687 ( .A1(n9473), .A2(n9589), .B1(n9472), .B2(n9599), .ZN(n9387)
         );
  AOI211_X1 U10688 ( .C1(P1_REG3_REG_27__SCAN_IN), .C2(P1_U3084), .A(n9388), 
        .B(n9387), .ZN(n9389) );
  OAI211_X1 U10689 ( .C1(n9598), .C2(n9478), .A(n9390), .B(n9389), .ZN(
        P1_U3212) );
  NAND2_X1 U10690 ( .A1(n9391), .A2(n9392), .ZN(n9394) );
  XNOR2_X1 U10691 ( .A(n9394), .B(n9393), .ZN(n9395) );
  NAND2_X1 U10692 ( .A1(n9395), .A2(n9467), .ZN(n9400) );
  OAI22_X1 U10693 ( .A1(n9455), .A2(n9688), .B1(n9472), .B2(n9656), .ZN(n9398)
         );
  OAI22_X1 U10694 ( .A1(n9473), .A2(n9635), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9396), .ZN(n9397) );
  NOR2_X1 U10695 ( .A1(n9398), .A2(n9397), .ZN(n9399) );
  OAI211_X1 U10696 ( .C1(n9659), .C2(n9478), .A(n9400), .B(n9399), .ZN(
        P1_U3214) );
  XNOR2_X1 U10697 ( .A(n4487), .B(n9401), .ZN(n9402) );
  XNOR2_X1 U10698 ( .A(n9403), .B(n9402), .ZN(n9409) );
  NOR2_X1 U10699 ( .A1(n9404), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9555) );
  OAI22_X1 U10700 ( .A1(n9473), .A2(n9715), .B1(n9472), .B2(n9405), .ZN(n9406)
         );
  AOI211_X1 U10701 ( .C1(n9475), .C2(n9732), .A(n9555), .B(n9406), .ZN(n9408)
         );
  NAND2_X1 U10702 ( .A1(n9798), .A2(n9459), .ZN(n9407) );
  OAI211_X1 U10703 ( .C1(n9409), .C2(n9461), .A(n9408), .B(n9407), .ZN(
        P1_U3217) );
  AOI21_X1 U10704 ( .B1(n9411), .B2(n9410), .A(n4530), .ZN(n9416) );
  OAI22_X1 U10705 ( .A1(n9473), .A2(n9688), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9412), .ZN(n9414) );
  OAI22_X1 U10706 ( .A1(n9455), .A2(n9715), .B1(n9472), .B2(n9691), .ZN(n9413)
         );
  AOI211_X1 U10707 ( .C1(n9788), .C2(n9459), .A(n9414), .B(n9413), .ZN(n9415)
         );
  OAI21_X1 U10708 ( .B1(n9416), .B2(n9461), .A(n9415), .ZN(P1_U3221) );
  OAI21_X1 U10709 ( .B1(n9418), .B2(n9417), .A(n6275), .ZN(n9419) );
  NAND2_X1 U10710 ( .A1(n9419), .A2(n9467), .ZN(n9424) );
  OAI22_X1 U10711 ( .A1(n9473), .A2(n9634), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9420), .ZN(n9422) );
  OAI22_X1 U10712 ( .A1(n9455), .A2(n9635), .B1(n9472), .B2(n9625), .ZN(n9421)
         );
  AOI211_X1 U10713 ( .C1(n9768), .C2(n9459), .A(n9422), .B(n9421), .ZN(n9423)
         );
  NAND2_X1 U10714 ( .A1(n9424), .A2(n9423), .ZN(P1_U3223) );
  XOR2_X1 U10715 ( .A(n9426), .B(n9425), .Z(n9432) );
  NOR2_X1 U10716 ( .A1(n9737), .A2(n10136), .ZN(n9905) );
  NAND2_X1 U10717 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9523) );
  OAI21_X1 U10718 ( .B1(n9473), .B2(n9717), .A(n9523), .ZN(n9429) );
  OAI22_X1 U10719 ( .A1(n9455), .A2(n9427), .B1(n9472), .B2(n9734), .ZN(n9428)
         );
  AOI211_X1 U10720 ( .C1(n9905), .C2(n9430), .A(n9429), .B(n9428), .ZN(n9431)
         );
  OAI21_X1 U10721 ( .B1(n9432), .B2(n9461), .A(n9431), .ZN(P1_U3226) );
  INV_X1 U10722 ( .A(n9772), .ZN(n9648) );
  INV_X1 U10723 ( .A(n9433), .ZN(n9437) );
  AOI21_X1 U10724 ( .B1(n9391), .B2(n9435), .A(n9434), .ZN(n9436) );
  OAI21_X1 U10725 ( .B1(n9437), .B2(n9436), .A(n9467), .ZN(n9442) );
  NOR2_X1 U10726 ( .A1(n9473), .A2(n9438), .ZN(n9440) );
  OAI22_X1 U10727 ( .A1(n9455), .A2(n9456), .B1(n9472), .B2(n9646), .ZN(n9439)
         );
  AOI211_X1 U10728 ( .C1(P1_REG3_REG_24__SCAN_IN), .C2(P1_U3084), .A(n9440), 
        .B(n9439), .ZN(n9441) );
  OAI211_X1 U10729 ( .C1(n9648), .C2(n9478), .A(n9442), .B(n9441), .ZN(
        P1_U3227) );
  AOI21_X1 U10730 ( .B1(n9445), .B2(n9444), .A(n9443), .ZN(n9450) );
  INV_X1 U10731 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9446) );
  OAI22_X1 U10732 ( .A1(n9473), .A2(n9707), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9446), .ZN(n9448) );
  OAI22_X1 U10733 ( .A1(n9455), .A2(n9708), .B1(n9472), .B2(n9700), .ZN(n9447)
         );
  AOI211_X1 U10734 ( .C1(n9793), .C2(n9459), .A(n9448), .B(n9447), .ZN(n9449)
         );
  OAI21_X1 U10735 ( .B1(n9450), .B2(n9461), .A(n9449), .ZN(P1_U3231) );
  NAND2_X1 U10736 ( .A1(n5023), .A2(n9451), .ZN(n9453) );
  XNOR2_X1 U10737 ( .A(n9453), .B(n9452), .ZN(n9462) );
  OAI22_X1 U10738 ( .A1(n9455), .A2(n9707), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9454), .ZN(n9458) );
  OAI22_X1 U10739 ( .A1(n9473), .A2(n9456), .B1(n9472), .B2(n9671), .ZN(n9457)
         );
  AOI211_X1 U10740 ( .C1(n9781), .C2(n9459), .A(n9458), .B(n9457), .ZN(n9460)
         );
  OAI21_X1 U10741 ( .B1(n9462), .B2(n9461), .A(n9460), .ZN(P1_U3233) );
  INV_X1 U10742 ( .A(n9463), .ZN(n9469) );
  OAI21_X1 U10743 ( .B1(n9465), .B2(n9468), .A(n9464), .ZN(n9466) );
  OAI211_X1 U10744 ( .C1(n9469), .C2(n9468), .A(n9467), .B(n9466), .ZN(n9477)
         );
  INV_X1 U10745 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9470) );
  NOR2_X1 U10746 ( .A1(n9470), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9533) );
  OAI22_X1 U10747 ( .A1(n9473), .A2(n9708), .B1(n9472), .B2(n9471), .ZN(n9474)
         );
  AOI211_X1 U10748 ( .C1(n9475), .C2(n9486), .A(n9533), .B(n9474), .ZN(n9476)
         );
  OAI211_X1 U10749 ( .C1(n9479), .C2(n9478), .A(n9477), .B(n9476), .ZN(
        P1_U3236) );
  MUX2_X1 U10750 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9480), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10751 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9481), .S(n9494), .Z(
        P1_U3584) );
  MUX2_X1 U10752 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9482), .S(n9494), .Z(
        P1_U3583) );
  MUX2_X1 U10753 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9606), .S(n9494), .Z(
        P1_U3582) );
  MUX2_X1 U10754 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9483), .S(n9494), .Z(
        P1_U3581) );
  MUX2_X1 U10755 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9641), .S(n9494), .Z(
        P1_U3580) );
  MUX2_X1 U10756 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9662), .S(n9494), .Z(
        P1_U3579) );
  MUX2_X1 U10757 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9677), .S(n9494), .Z(
        P1_U3578) );
  MUX2_X1 U10758 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9663), .S(n9494), .Z(
        P1_U3577) );
  MUX2_X1 U10759 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9678), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10760 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9484), .S(n9494), .Z(
        P1_U3575) );
  MUX2_X1 U10761 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9485), .S(n9494), .Z(
        P1_U3574) );
  MUX2_X1 U10762 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9732), .S(n9494), .Z(
        P1_U3573) );
  MUX2_X1 U10763 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9486), .S(n9494), .Z(
        P1_U3572) );
  MUX2_X1 U10764 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9731), .S(n9494), .Z(
        P1_U3571) );
  MUX2_X1 U10765 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9487), .S(n9494), .Z(
        P1_U3570) );
  MUX2_X1 U10766 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9488), .S(n9494), .Z(
        P1_U3569) );
  MUX2_X1 U10767 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9489), .S(n9494), .Z(
        P1_U3568) );
  MUX2_X1 U10768 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9490), .S(n9494), .Z(
        P1_U3567) );
  MUX2_X1 U10769 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9491), .S(n9494), .Z(
        P1_U3566) );
  MUX2_X1 U10770 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n10023), .S(n9494), .Z(
        P1_U3565) );
  MUX2_X1 U10771 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9492), .S(n9494), .Z(
        P1_U3564) );
  MUX2_X1 U10772 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n10022), .S(n9494), .Z(
        P1_U3563) );
  MUX2_X1 U10773 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9493), .S(n9494), .Z(
        P1_U3562) );
  MUX2_X1 U10774 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9495), .S(n9494), .Z(
        P1_U3561) );
  MUX2_X1 U10775 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9496), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10776 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9497), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10777 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9498), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10778 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n5785), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10779 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9499), .S(P1_U4006), .Z(
        P1_U3556) );
  OAI21_X1 U10780 ( .B1(n9502), .B2(n9501), .A(n9500), .ZN(n9503) );
  NAND2_X1 U10781 ( .A1(n9503), .A2(n10010), .ZN(n9513) );
  NOR2_X1 U10782 ( .A1(n9525), .A2(n9504), .ZN(n9505) );
  AOI211_X1 U10783 ( .C1(n10013), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9506), .B(
        n9505), .ZN(n9512) );
  OAI21_X1 U10784 ( .B1(n9509), .B2(n9508), .A(n9507), .ZN(n9510) );
  NAND2_X1 U10785 ( .A1(n9510), .A2(n9994), .ZN(n9511) );
  NAND3_X1 U10786 ( .A1(n9513), .A2(n9512), .A3(n9511), .ZN(P1_U3249) );
  AOI21_X1 U10787 ( .B1(n9518), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9514), .ZN(
        n9516) );
  MUX2_X1 U10788 ( .A(n6703), .B(P1_REG2_REG_17__SCAN_IN), .S(n9537), .Z(n9515) );
  AOI211_X1 U10789 ( .C1(n9516), .C2(n9515), .A(n10003), .B(n9536), .ZN(n9528)
         );
  AOI21_X1 U10790 ( .B1(n9518), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9517), .ZN(
        n9521) );
  MUX2_X1 U10791 ( .A(n9519), .B(P1_REG1_REG_17__SCAN_IN), .S(n9537), .Z(n9520) );
  NOR2_X1 U10792 ( .A1(n9521), .A2(n9520), .ZN(n9529) );
  AOI211_X1 U10793 ( .C1(n9521), .C2(n9520), .A(n9969), .B(n9529), .ZN(n9527)
         );
  NAND2_X1 U10794 ( .A1(n10013), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9522) );
  OAI211_X1 U10795 ( .C1(n9525), .C2(n9524), .A(n9523), .B(n9522), .ZN(n9526)
         );
  OR3_X1 U10796 ( .A1(n9528), .A2(n9527), .A3(n9526), .ZN(P1_U3258) );
  AOI21_X1 U10797 ( .B1(n9537), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9529), .ZN(
        n9532) );
  XNOR2_X1 U10798 ( .A(n9548), .B(n9530), .ZN(n9531) );
  NAND2_X1 U10799 ( .A1(n9531), .A2(n9532), .ZN(n9547) );
  OAI21_X1 U10800 ( .B1(n9532), .B2(n9531), .A(n9547), .ZN(n9543) );
  INV_X1 U10801 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9535) );
  AOI21_X1 U10802 ( .B1(n10012), .B2(n9548), .A(n9533), .ZN(n9534) );
  OAI21_X1 U10803 ( .B1(n9999), .B2(n9535), .A(n9534), .ZN(n9542) );
  NAND2_X1 U10804 ( .A1(n9548), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9538) );
  OAI21_X1 U10805 ( .B1(n9548), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9538), .ZN(
        n9539) );
  AOI211_X1 U10806 ( .C1(n9540), .C2(n9539), .A(n9545), .B(n10003), .ZN(n9541)
         );
  AOI211_X1 U10807 ( .C1(n10010), .C2(n9543), .A(n9542), .B(n9541), .ZN(n9544)
         );
  INV_X1 U10808 ( .A(n9544), .ZN(P1_U3259) );
  XNOR2_X1 U10809 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9546), .ZN(n9554) );
  INV_X1 U10810 ( .A(n9554), .ZN(n9550) );
  OAI21_X1 U10811 ( .B1(n9548), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9547), .ZN(
        n9549) );
  XOR2_X1 U10812 ( .A(n9549), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9552) );
  INV_X1 U10813 ( .A(n9551), .ZN(n9953) );
  AOI21_X1 U10814 ( .B1(n9552), .B2(n10010), .A(n10012), .ZN(n9553) );
  NAND2_X1 U10815 ( .A1(n9901), .A2(n9562), .ZN(n9556) );
  XNOR2_X1 U10816 ( .A(n9876), .B(n9556), .ZN(n9874) );
  AND2_X1 U10817 ( .A1(n9558), .A2(n9557), .ZN(n9903) );
  NAND2_X1 U10818 ( .A1(n10031), .A2(n9903), .ZN(n9563) );
  OAI21_X1 U10819 ( .B1(n10057), .B2(n9559), .A(n9563), .ZN(n9560) );
  AOI21_X1 U10820 ( .B1(n9876), .B2(n9739), .A(n9560), .ZN(n9561) );
  OAI21_X1 U10821 ( .B1(n9874), .B2(n10019), .A(n9561), .ZN(P1_U3261) );
  XNOR2_X1 U10822 ( .A(n9562), .B(n8286), .ZN(n9904) );
  NAND2_X1 U10823 ( .A1(n9904), .A2(n9682), .ZN(n9566) );
  INV_X1 U10824 ( .A(n9563), .ZN(n9564) );
  AOI21_X1 U10825 ( .B1(n9738), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9564), .ZN(
        n9565) );
  OAI211_X1 U10826 ( .C1(n9901), .C2(n9724), .A(n9566), .B(n9565), .ZN(
        P1_U3262) );
  AND2_X1 U10827 ( .A1(n9568), .A2(n9567), .ZN(n9569) );
  AND2_X1 U10828 ( .A1(n9572), .A2(n9571), .ZN(n9573) );
  OAI21_X1 U10829 ( .B1(n4493), .B2(n9573), .A(n10050), .ZN(n9578) );
  OAI22_X1 U10830 ( .A1(n9575), .A2(n6463), .B1(n9574), .B2(n9716), .ZN(n9576)
         );
  INV_X1 U10831 ( .A(n9576), .ZN(n9577) );
  NAND2_X1 U10832 ( .A1(n9578), .A2(n9577), .ZN(n9751) );
  NAND2_X1 U10833 ( .A1(n9596), .A2(n9584), .ZN(n9579) );
  NAND2_X1 U10834 ( .A1(n9580), .A2(n9579), .ZN(n9749) );
  OAI22_X1 U10835 ( .A1(n10057), .A2(n9582), .B1(n9581), .B2(n10036), .ZN(
        n9583) );
  AOI21_X1 U10836 ( .B1(n9584), .B2(n9739), .A(n9583), .ZN(n9585) );
  OAI21_X1 U10837 ( .B1(n9749), .B2(n10019), .A(n9585), .ZN(n9586) );
  AOI21_X1 U10838 ( .B1(n9751), .B2(n10031), .A(n9586), .ZN(n9587) );
  OAI21_X1 U10839 ( .B1(n9747), .B2(n9746), .A(n9587), .ZN(P1_U3263) );
  AOI21_X1 U10840 ( .B1(n9588), .B2(n9594), .A(n6466), .ZN(n9592) );
  OAI22_X1 U10841 ( .A1(n9589), .A2(n9716), .B1(n9634), .B2(n6463), .ZN(n9590)
         );
  AOI21_X1 U10842 ( .B1(n9592), .B2(n9591), .A(n9590), .ZN(n9758) );
  OAI21_X1 U10843 ( .B1(n9595), .B2(n9594), .A(n9593), .ZN(n9754) );
  NAND2_X1 U10844 ( .A1(n9754), .A2(n9611), .ZN(n9604) );
  INV_X1 U10845 ( .A(n9612), .ZN(n9597) );
  AOI211_X1 U10846 ( .C1(n9756), .C2(n9597), .A(n10154), .B(n4697), .ZN(n9755)
         );
  NOR2_X1 U10847 ( .A1(n9598), .A2(n9724), .ZN(n9602) );
  OAI22_X1 U10848 ( .A1(n10031), .A2(n9600), .B1(n9599), .B2(n10036), .ZN(
        n9601) );
  AOI211_X1 U10849 ( .C1(n9755), .C2(n9720), .A(n9602), .B(n9601), .ZN(n9603)
         );
  OAI211_X1 U10850 ( .C1(n9738), .C2(n9758), .A(n9604), .B(n9603), .ZN(
        P1_U3264) );
  XNOR2_X1 U10851 ( .A(n9605), .B(n9609), .ZN(n9607) );
  AOI222_X1 U10852 ( .A1(n10050), .A2(n9607), .B1(n9641), .B2(n10045), .C1(
        n9606), .C2(n10046), .ZN(n9764) );
  OAI21_X1 U10853 ( .B1(n9610), .B2(n9609), .A(n9608), .ZN(n9760) );
  NAND2_X1 U10854 ( .A1(n9760), .A2(n9611), .ZN(n9620) );
  INV_X1 U10855 ( .A(n9622), .ZN(n9613) );
  AOI21_X1 U10856 ( .B1(n9761), .B2(n9613), .A(n9612), .ZN(n9762) );
  NOR2_X1 U10857 ( .A1(n9614), .A2(n9724), .ZN(n9618) );
  OAI22_X1 U10858 ( .A1(n10031), .A2(n9616), .B1(n9615), .B2(n10036), .ZN(
        n9617) );
  AOI211_X1 U10859 ( .C1(n9762), .C2(n9682), .A(n9618), .B(n9617), .ZN(n9619)
         );
  OAI211_X1 U10860 ( .C1(n9738), .C2(n9764), .A(n9620), .B(n9619), .ZN(
        P1_U3265) );
  XOR2_X1 U10861 ( .A(n9621), .B(n9632), .Z(n9770) );
  INV_X1 U10862 ( .A(n9643), .ZN(n9623) );
  AOI211_X1 U10863 ( .C1(n9768), .C2(n9623), .A(n10154), .B(n9622), .ZN(n9767)
         );
  NOR2_X1 U10864 ( .A1(n9624), .A2(n9724), .ZN(n9628) );
  OAI22_X1 U10865 ( .A1(n10057), .A2(n9626), .B1(n9625), .B2(n10036), .ZN(
        n9627) );
  AOI211_X1 U10866 ( .C1(n9767), .C2(n9720), .A(n9628), .B(n9627), .ZN(n9637)
         );
  NAND2_X1 U10867 ( .A1(n9629), .A2(n9630), .ZN(n9631) );
  XOR2_X1 U10868 ( .A(n9632), .B(n9631), .Z(n9633) );
  OAI222_X1 U10869 ( .A1(n6463), .A2(n9635), .B1(n9716), .B2(n9634), .C1(n9633), .C2(n6466), .ZN(n9766) );
  NAND2_X1 U10870 ( .A1(n9766), .A2(n10031), .ZN(n9636) );
  OAI211_X1 U10871 ( .C1(n9770), .C2(n9746), .A(n9637), .B(n9636), .ZN(
        P1_U3266) );
  XNOR2_X1 U10872 ( .A(n9638), .B(n9640), .ZN(n9775) );
  OAI21_X1 U10873 ( .B1(n9640), .B2(n9639), .A(n9629), .ZN(n9642) );
  AOI222_X1 U10874 ( .A1(n10050), .A2(n9642), .B1(n9641), .B2(n10046), .C1(
        n9677), .C2(n10045), .ZN(n9774) );
  AOI211_X1 U10875 ( .C1(n9772), .C2(n9654), .A(n10154), .B(n9643), .ZN(n9771)
         );
  NAND2_X1 U10876 ( .A1(n9771), .A2(n9644), .ZN(n9645) );
  OAI211_X1 U10877 ( .C1(n10036), .C2(n9646), .A(n9774), .B(n9645), .ZN(n9650)
         );
  OAI22_X1 U10878 ( .A1(n9648), .A2(n9724), .B1(n9647), .B2(n10031), .ZN(n9649) );
  AOI21_X1 U10879 ( .B1(n9650), .B2(n10031), .A(n9649), .ZN(n9651) );
  OAI21_X1 U10880 ( .B1(n9775), .B2(n9746), .A(n9651), .ZN(P1_U3267) );
  XNOR2_X1 U10881 ( .A(n9653), .B(n9652), .ZN(n9780) );
  INV_X1 U10882 ( .A(n9654), .ZN(n9655) );
  AOI21_X1 U10883 ( .B1(n9776), .B2(n9669), .A(n9655), .ZN(n9777) );
  INV_X1 U10884 ( .A(n9656), .ZN(n9657) );
  AOI22_X1 U10885 ( .A1(n9738), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9657), .B2(
        n10041), .ZN(n9658) );
  OAI21_X1 U10886 ( .B1(n9659), .B2(n9724), .A(n9658), .ZN(n9666) );
  XNOR2_X1 U10887 ( .A(n9660), .B(n9661), .ZN(n9664) );
  AOI222_X1 U10888 ( .A1(n10050), .A2(n9664), .B1(n9663), .B2(n10045), .C1(
        n9662), .C2(n10046), .ZN(n9779) );
  NOR2_X1 U10889 ( .A1(n9779), .A2(n9738), .ZN(n9665) );
  AOI211_X1 U10890 ( .C1(n9777), .C2(n9682), .A(n9666), .B(n9665), .ZN(n9667)
         );
  OAI21_X1 U10891 ( .B1(n9780), .B2(n9746), .A(n9667), .ZN(P1_U3268) );
  XOR2_X1 U10892 ( .A(n9668), .B(n9675), .Z(n9785) );
  INV_X1 U10893 ( .A(n9689), .ZN(n9670) );
  AOI21_X1 U10894 ( .B1(n9781), .B2(n9670), .A(n4688), .ZN(n9782) );
  INV_X1 U10895 ( .A(n9671), .ZN(n9672) );
  AOI22_X1 U10896 ( .A1(n9738), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9672), .B2(
        n10041), .ZN(n9673) );
  OAI21_X1 U10897 ( .B1(n9674), .B2(n9724), .A(n9673), .ZN(n9681) );
  XNOR2_X1 U10898 ( .A(n9676), .B(n9675), .ZN(n9679) );
  AOI222_X1 U10899 ( .A1(n10050), .A2(n9679), .B1(n9678), .B2(n10045), .C1(
        n9677), .C2(n10046), .ZN(n9784) );
  NOR2_X1 U10900 ( .A1(n9784), .A2(n9738), .ZN(n9680) );
  AOI211_X1 U10901 ( .C1(n9782), .C2(n9682), .A(n9681), .B(n9680), .ZN(n9683)
         );
  OAI21_X1 U10902 ( .B1(n9785), .B2(n9746), .A(n9683), .ZN(P1_U3269) );
  XNOR2_X1 U10903 ( .A(n9684), .B(n9685), .ZN(n9790) );
  AOI22_X1 U10904 ( .A1(n9788), .A2(n9739), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9738), .ZN(n9695) );
  XOR2_X1 U10905 ( .A(n9686), .B(n9685), .Z(n9687) );
  OAI222_X1 U10906 ( .A1(n9716), .A2(n9688), .B1(n6463), .B2(n9715), .C1(n6466), .C2(n9687), .ZN(n9786) );
  INV_X1 U10907 ( .A(n9697), .ZN(n9690) );
  AOI211_X1 U10908 ( .C1(n9788), .C2(n9690), .A(n10154), .B(n9689), .ZN(n9787)
         );
  INV_X1 U10909 ( .A(n9787), .ZN(n9692) );
  OAI22_X1 U10910 ( .A1(n9692), .A2(n10044), .B1(n10036), .B2(n9691), .ZN(
        n9693) );
  OAI21_X1 U10911 ( .B1(n9786), .B2(n9693), .A(n10031), .ZN(n9694) );
  OAI211_X1 U10912 ( .C1(n9790), .C2(n9746), .A(n9695), .B(n9694), .ZN(
        P1_U3270) );
  XNOR2_X1 U10913 ( .A(n9696), .B(n9704), .ZN(n9795) );
  INV_X1 U10914 ( .A(n9718), .ZN(n9698) );
  AOI211_X1 U10915 ( .C1(n9793), .C2(n9698), .A(n10154), .B(n9697), .ZN(n9792)
         );
  NOR2_X1 U10916 ( .A1(n9699), .A2(n9724), .ZN(n9703) );
  OAI22_X1 U10917 ( .A1(n10057), .A2(n9701), .B1(n9700), .B2(n10036), .ZN(
        n9702) );
  AOI211_X1 U10918 ( .C1(n9792), .C2(n9720), .A(n9703), .B(n9702), .ZN(n9710)
         );
  XNOR2_X1 U10919 ( .A(n9705), .B(n9704), .ZN(n9706) );
  OAI222_X1 U10920 ( .A1(n6463), .A2(n9708), .B1(n9716), .B2(n9707), .C1(n6466), .C2(n9706), .ZN(n9791) );
  NAND2_X1 U10921 ( .A1(n9791), .A2(n10057), .ZN(n9709) );
  OAI211_X1 U10922 ( .C1(n9795), .C2(n9746), .A(n9710), .B(n9709), .ZN(
        P1_U3271) );
  XNOR2_X1 U10923 ( .A(n9711), .B(n9713), .ZN(n9800) );
  AOI21_X1 U10924 ( .B1(n9713), .B2(n9712), .A(n4499), .ZN(n9714) );
  OAI222_X1 U10925 ( .A1(n6463), .A2(n9717), .B1(n9716), .B2(n9715), .C1(n6466), .C2(n9714), .ZN(n9796) );
  INV_X1 U10926 ( .A(n9798), .ZN(n9725) );
  AOI211_X1 U10927 ( .C1(n9798), .C2(n9719), .A(n10154), .B(n9718), .ZN(n9797)
         );
  NAND2_X1 U10928 ( .A1(n9797), .A2(n9720), .ZN(n9723) );
  AOI22_X1 U10929 ( .A1(n9738), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9721), .B2(
        n10041), .ZN(n9722) );
  OAI211_X1 U10930 ( .C1(n9725), .C2(n9724), .A(n9723), .B(n9722), .ZN(n9726)
         );
  AOI21_X1 U10931 ( .B1(n9796), .B2(n10031), .A(n9726), .ZN(n9727) );
  OAI21_X1 U10932 ( .B1(n9800), .B2(n9746), .A(n9727), .ZN(P1_U3272) );
  XNOR2_X1 U10933 ( .A(n9728), .B(n9729), .ZN(n9910) );
  INV_X1 U10934 ( .A(n9910), .ZN(n9745) );
  XOR2_X1 U10935 ( .A(n9730), .B(n9729), .Z(n9733) );
  AOI222_X1 U10936 ( .A1(n10050), .A2(n9733), .B1(n9732), .B2(n10046), .C1(
        n9731), .C2(n10045), .ZN(n9907) );
  OAI21_X1 U10937 ( .B1(n9734), .B2(n10036), .A(n9907), .ZN(n9743) );
  OAI21_X1 U10938 ( .B1(n4704), .B2(n9737), .A(n9736), .ZN(n9908) );
  AOI22_X1 U10939 ( .A1(n9740), .A2(n9739), .B1(P1_REG2_REG_17__SCAN_IN), .B2(
        n9738), .ZN(n9741) );
  OAI21_X1 U10940 ( .B1(n9908), .B2(n10019), .A(n9741), .ZN(n9742) );
  AOI21_X1 U10941 ( .B1(n9743), .B2(n10031), .A(n9742), .ZN(n9744) );
  OAI21_X1 U10942 ( .B1(n9746), .B2(n9745), .A(n9744), .ZN(P1_U3274) );
  OAI22_X1 U10943 ( .A1(n9749), .A2(n10154), .B1(n9748), .B2(n10136), .ZN(
        n9750) );
  NOR2_X1 U10944 ( .A1(n9751), .A2(n9750), .ZN(n9752) );
  NAND2_X1 U10945 ( .A1(n9753), .A2(n9752), .ZN(n9813) );
  MUX2_X1 U10946 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9813), .S(n10173), .Z(
        P1_U3551) );
  INV_X1 U10947 ( .A(n9754), .ZN(n9759) );
  AOI21_X1 U10948 ( .B1(n10149), .B2(n9756), .A(n9755), .ZN(n9757) );
  OAI211_X1 U10949 ( .C1(n9759), .C2(n10141), .A(n9758), .B(n9757), .ZN(n9814)
         );
  MUX2_X1 U10950 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9814), .S(n10173), .Z(
        P1_U3550) );
  INV_X1 U10951 ( .A(n9760), .ZN(n9765) );
  AOI22_X1 U10952 ( .A1(n9762), .A2(n10124), .B1(n10149), .B2(n9761), .ZN(
        n9763) );
  OAI211_X1 U10953 ( .C1(n9765), .C2(n10141), .A(n9764), .B(n9763), .ZN(n9815)
         );
  MUX2_X1 U10954 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9815), .S(n10173), .Z(
        P1_U3549) );
  AOI211_X1 U10955 ( .C1(n10149), .C2(n9768), .A(n9767), .B(n9766), .ZN(n9769)
         );
  OAI21_X1 U10956 ( .B1(n9770), .B2(n10141), .A(n9769), .ZN(n9816) );
  MUX2_X1 U10957 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9816), .S(n10173), .Z(
        P1_U3548) );
  AOI21_X1 U10958 ( .B1(n10149), .B2(n9772), .A(n9771), .ZN(n9773) );
  OAI211_X1 U10959 ( .C1(n9775), .C2(n10141), .A(n9774), .B(n9773), .ZN(n9817)
         );
  MUX2_X1 U10960 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9817), .S(n10173), .Z(
        P1_U3547) );
  AOI22_X1 U10961 ( .A1(n9777), .A2(n10124), .B1(n10149), .B2(n9776), .ZN(
        n9778) );
  OAI211_X1 U10962 ( .C1(n9780), .C2(n10141), .A(n9779), .B(n9778), .ZN(n9818)
         );
  MUX2_X1 U10963 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9818), .S(n10173), .Z(
        P1_U3546) );
  AOI22_X1 U10964 ( .A1(n9782), .A2(n10124), .B1(n10149), .B2(n9781), .ZN(
        n9783) );
  OAI211_X1 U10965 ( .C1(n9785), .C2(n10141), .A(n9784), .B(n9783), .ZN(n9819)
         );
  MUX2_X1 U10966 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9819), .S(n10173), .Z(
        P1_U3545) );
  AOI211_X1 U10967 ( .C1(n10149), .C2(n9788), .A(n9787), .B(n9786), .ZN(n9789)
         );
  OAI21_X1 U10968 ( .B1(n9790), .B2(n10141), .A(n9789), .ZN(n9820) );
  MUX2_X1 U10969 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9820), .S(n10173), .Z(
        P1_U3544) );
  AOI211_X1 U10970 ( .C1(n10149), .C2(n9793), .A(n9792), .B(n9791), .ZN(n9794)
         );
  OAI21_X1 U10971 ( .B1(n9795), .B2(n10141), .A(n9794), .ZN(n9821) );
  MUX2_X1 U10972 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9821), .S(n10173), .Z(
        P1_U3543) );
  AOI211_X1 U10973 ( .C1(n10149), .C2(n9798), .A(n9797), .B(n9796), .ZN(n9799)
         );
  OAI21_X1 U10974 ( .B1(n10141), .B2(n9800), .A(n9799), .ZN(n9822) );
  MUX2_X1 U10975 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9822), .S(n10173), .Z(
        P1_U3542) );
  AOI211_X1 U10976 ( .C1(n10149), .C2(n9803), .A(n9802), .B(n9801), .ZN(n9804)
         );
  OAI21_X1 U10977 ( .B1(n9805), .B2(n10141), .A(n9804), .ZN(n9823) );
  MUX2_X1 U10978 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9823), .S(n10173), .Z(
        P1_U3541) );
  AOI211_X1 U10979 ( .C1(n10149), .C2(n9808), .A(n9807), .B(n9806), .ZN(n9809)
         );
  OAI21_X1 U10980 ( .B1(n10141), .B2(n9810), .A(n9809), .ZN(n9824) );
  MUX2_X1 U10981 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9824), .S(n10173), .Z(
        P1_U3537) );
  MUX2_X1 U10982 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9811), .S(n10173), .Z(
        P1_U3523) );
  MUX2_X1 U10983 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9812), .S(n10160), .Z(
        P1_U3520) );
  MUX2_X1 U10984 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9813), .S(n10160), .Z(
        P1_U3519) );
  MUX2_X1 U10985 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9814), .S(n10160), .Z(
        P1_U3518) );
  MUX2_X1 U10986 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9815), .S(n10160), .Z(
        P1_U3517) );
  MUX2_X1 U10987 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9816), .S(n10160), .Z(
        P1_U3516) );
  MUX2_X1 U10988 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9817), .S(n10160), .Z(
        P1_U3515) );
  MUX2_X1 U10989 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9818), .S(n10160), .Z(
        P1_U3514) );
  MUX2_X1 U10990 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9819), .S(n10160), .Z(
        P1_U3513) );
  MUX2_X1 U10991 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9820), .S(n10160), .Z(
        P1_U3512) );
  MUX2_X1 U10992 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9821), .S(n10160), .Z(
        P1_U3511) );
  MUX2_X1 U10993 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9822), .S(n10160), .Z(
        P1_U3510) );
  MUX2_X1 U10994 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9823), .S(n10160), .Z(
        P1_U3508) );
  MUX2_X1 U10995 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9824), .S(n10160), .Z(
        P1_U3496) );
  INV_X1 U10996 ( .A(n9825), .ZN(n9827) );
  NOR4_X1 U10997 ( .A1(n9827), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9826), .ZN(n9828) );
  AOI21_X1 U10998 ( .B1(n9836), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9828), .ZN(
        n9829) );
  OAI21_X1 U10999 ( .B1(n9830), .B2(n9835), .A(n9829), .ZN(P1_U3322) );
  OAI222_X1 U11000 ( .A1(n9835), .A2(n9834), .B1(n9833), .B2(P1_U3084), .C1(
        n9832), .C2(n9831), .ZN(P1_U3324) );
  NAND2_X1 U11001 ( .A1(n9836), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9837) );
  OAI211_X1 U11002 ( .C1(n9838), .C2(n9835), .A(n9837), .B(n9949), .ZN(
        P1_U3325) );
  MUX2_X1 U11003 ( .A(n9839), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U11004 ( .A(n9840), .ZN(n9841) );
  AOI21_X1 U11005 ( .B1(n10176), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n9841), .ZN(
        n9852) );
  INV_X1 U11006 ( .A(n10174), .ZN(n10180) );
  AOI211_X1 U11007 ( .C1(n9844), .C2(n9843), .A(n9842), .B(n10180), .ZN(n9845)
         );
  AOI21_X1 U11008 ( .B1(n9860), .B2(n9846), .A(n9845), .ZN(n9851) );
  AND2_X1 U11009 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9849) );
  OAI211_X1 U11010 ( .C1(n9849), .C2(n9848), .A(n10177), .B(n9847), .ZN(n9850)
         );
  NAND3_X1 U11011 ( .A1(n9852), .A2(n9851), .A3(n9850), .ZN(P2_U3246) );
  AOI21_X1 U11012 ( .B1(n10176), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n9853), .ZN(
        n9866) );
  OAI21_X1 U11013 ( .B1(n9856), .B2(n9855), .A(n9854), .ZN(n9857) );
  INV_X1 U11014 ( .A(n9857), .ZN(n9858) );
  AOI22_X1 U11015 ( .A1(n9860), .A2(n9859), .B1(n10174), .B2(n9858), .ZN(n9865) );
  OAI211_X1 U11016 ( .C1(n9863), .C2(n9862), .A(n10177), .B(n9861), .ZN(n9864)
         );
  NAND3_X1 U11017 ( .A1(n9866), .A2(n9865), .A3(n9864), .ZN(P2_U3247) );
  INV_X1 U11018 ( .A(n10141), .ZN(n10156) );
  OAI211_X1 U11019 ( .C1(n9869), .C2(n10136), .A(n9868), .B(n9867), .ZN(n9870)
         );
  AOI21_X1 U11020 ( .B1(n10156), .B2(n9871), .A(n9870), .ZN(n9873) );
  INV_X1 U11021 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9872) );
  AOI22_X1 U11022 ( .A1(n10160), .A2(n9873), .B1(n9872), .B2(n10158), .ZN(
        P1_U3484) );
  AOI22_X1 U11023 ( .A1(n10173), .A2(n9873), .B1(n5970), .B2(n10171), .ZN(
        P1_U3533) );
  NOR2_X1 U11024 ( .A1(n9874), .A2(n10154), .ZN(n9875) );
  INV_X1 U11025 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9877) );
  AOI22_X1 U11026 ( .A1(n10173), .A2(n9878), .B1(n9877), .B2(n10171), .ZN(
        P1_U3554) );
  AOI22_X1 U11027 ( .A1(n10160), .A2(n9878), .B1(n6910), .B2(n10158), .ZN(
        P1_U3522) );
  OAI21_X1 U11028 ( .B1(n9880), .B2(n10272), .A(n9879), .ZN(n9881) );
  AOI21_X1 U11029 ( .B1(n9882), .B2(n10231), .A(n9881), .ZN(n9896) );
  INV_X1 U11030 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9883) );
  AOI22_X1 U11031 ( .A1(n4449), .A2(n9896), .B1(n9883), .B2(n10292), .ZN(
        P2_U3550) );
  INV_X1 U11032 ( .A(n9884), .ZN(n9889) );
  OAI22_X1 U11033 ( .A1(n9886), .A2(n10273), .B1(n9885), .B2(n10272), .ZN(
        n9887) );
  AOI211_X1 U11034 ( .C1(n9889), .C2(n10278), .A(n9888), .B(n9887), .ZN(n9898)
         );
  AOI22_X1 U11035 ( .A1(n4449), .A2(n9898), .B1(n5367), .B2(n10292), .ZN(
        P2_U3534) );
  INV_X1 U11036 ( .A(n10245), .ZN(n10265) );
  INV_X1 U11037 ( .A(n9890), .ZN(n9895) );
  OAI22_X1 U11038 ( .A1(n9892), .A2(n10273), .B1(n9891), .B2(n10272), .ZN(
        n9894) );
  AOI211_X1 U11039 ( .C1(n10265), .C2(n9895), .A(n9894), .B(n9893), .ZN(n9900)
         );
  AOI22_X1 U11040 ( .A1(n4449), .A2(n9900), .B1(n5346), .B2(n10292), .ZN(
        P2_U3533) );
  AOI22_X1 U11041 ( .A1(n10281), .A2(n9896), .B1(n8602), .B2(n10279), .ZN(
        P2_U3518) );
  INV_X1 U11042 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9897) );
  AOI22_X1 U11043 ( .A1(n10281), .A2(n9898), .B1(n9897), .B2(n10279), .ZN(
        P2_U3493) );
  INV_X1 U11044 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9899) );
  AOI22_X1 U11045 ( .A1(n10281), .A2(n9900), .B1(n9899), .B2(n10279), .ZN(
        P2_U3490) );
  NOR2_X1 U11046 ( .A1(n9901), .A2(n10136), .ZN(n9902) );
  AOI211_X1 U11047 ( .C1(n10124), .C2(n9904), .A(n9903), .B(n9902), .ZN(n9934)
         );
  AOI22_X1 U11048 ( .A1(n10173), .A2(n9934), .B1(n6459), .B2(n10171), .ZN(
        P1_U3553) );
  INV_X1 U11049 ( .A(n9905), .ZN(n9906) );
  OAI211_X1 U11050 ( .C1(n10154), .C2(n9908), .A(n9907), .B(n9906), .ZN(n9909)
         );
  AOI21_X1 U11051 ( .B1(n9910), .B2(n10156), .A(n9909), .ZN(n9936) );
  AOI22_X1 U11052 ( .A1(n10173), .A2(n9936), .B1(n9519), .B2(n10171), .ZN(
        P1_U3540) );
  OAI211_X1 U11053 ( .C1(n9913), .C2(n10136), .A(n9912), .B(n9911), .ZN(n9914)
         );
  AOI21_X1 U11054 ( .B1(n9915), .B2(n10156), .A(n9914), .ZN(n9938) );
  AOI22_X1 U11055 ( .A1(n10173), .A2(n9938), .B1(n8083), .B2(n10171), .ZN(
        P1_U3539) );
  OAI211_X1 U11056 ( .C1(n9918), .C2(n10136), .A(n9917), .B(n9916), .ZN(n9921)
         );
  INV_X1 U11057 ( .A(n9922), .ZN(n9919) );
  NOR2_X1 U11058 ( .A1(n9919), .A2(n10128), .ZN(n9920) );
  AOI211_X1 U11059 ( .C1(n9922), .C2(n10133), .A(n9921), .B(n9920), .ZN(n9939)
         );
  AOI22_X1 U11060 ( .A1(n10173), .A2(n9939), .B1(n6072), .B2(n10171), .ZN(
        P1_U3538) );
  OAI22_X1 U11061 ( .A1(n9924), .A2(n10154), .B1(n9923), .B2(n10136), .ZN(
        n9926) );
  AOI211_X1 U11062 ( .C1(n9927), .C2(n10156), .A(n9926), .B(n9925), .ZN(n9941)
         );
  AOI22_X1 U11063 ( .A1(n10173), .A2(n9941), .B1(n7502), .B2(n10171), .ZN(
        P1_U3536) );
  OAI22_X1 U11064 ( .A1(n9929), .A2(n10154), .B1(n9928), .B2(n10136), .ZN(
        n9931) );
  AOI211_X1 U11065 ( .C1(n9932), .C2(n10156), .A(n9931), .B(n9930), .ZN(n9943)
         );
  AOI22_X1 U11066 ( .A1(n10173), .A2(n9943), .B1(n5988), .B2(n10171), .ZN(
        P1_U3534) );
  INV_X1 U11067 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9933) );
  AOI22_X1 U11068 ( .A1(n10160), .A2(n9934), .B1(n9933), .B2(n10158), .ZN(
        P1_U3521) );
  INV_X1 U11069 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9935) );
  AOI22_X1 U11070 ( .A1(n10160), .A2(n9936), .B1(n9935), .B2(n10158), .ZN(
        P1_U3505) );
  INV_X1 U11071 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9937) );
  AOI22_X1 U11072 ( .A1(n10160), .A2(n9938), .B1(n9937), .B2(n10158), .ZN(
        P1_U3502) );
  AOI22_X1 U11073 ( .A1(n10160), .A2(n9939), .B1(n6071), .B2(n10158), .ZN(
        P1_U3499) );
  INV_X1 U11074 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9940) );
  AOI22_X1 U11075 ( .A1(n10160), .A2(n9941), .B1(n9940), .B2(n10158), .ZN(
        P1_U3493) );
  AOI22_X1 U11076 ( .A1(n10160), .A2(n9943), .B1(n9942), .B2(n10158), .ZN(
        P1_U3487) );
  XNOR2_X1 U11077 ( .A(P1_WR_REG_SCAN_IN), .B(P2_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11078 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NOR2_X1 U11079 ( .A1(n9977), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9945) );
  OR2_X1 U11080 ( .A1(n9945), .A2(n6302), .ZN(n9947) );
  NAND2_X1 U11081 ( .A1(n9947), .A2(n9946), .ZN(n9980) );
  OAI21_X1 U11082 ( .B1(n9947), .B2(n9946), .A(n9980), .ZN(n9948) );
  INV_X1 U11083 ( .A(n9948), .ZN(n9955) );
  INV_X1 U11084 ( .A(n9949), .ZN(n9950) );
  NAND3_X1 U11085 ( .A1(n9951), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n9950), .ZN(
        n9952) );
  NAND2_X1 U11086 ( .A1(n9953), .A2(n9952), .ZN(n9954) );
  AOI22_X1 U11087 ( .A1(n10013), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(n9955), .B2(
        n9954), .ZN(n9958) );
  NAND3_X1 U11088 ( .A1(n10010), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9956), .ZN(
        n9957) );
  OAI211_X1 U11089 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n7247), .A(n9958), .B(
        n9957), .ZN(P1_U3241) );
  NAND2_X1 U11090 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9961) );
  AOI211_X1 U11091 ( .C1(n9961), .C2(n9960), .A(n9959), .B(n9969), .ZN(n9965)
         );
  AOI211_X1 U11092 ( .C1(n9979), .C2(n9963), .A(n9962), .B(n10003), .ZN(n9964)
         );
  AOI211_X1 U11093 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(P1_U3084), .A(n9965), 
        .B(n9964), .ZN(n9968) );
  AOI22_X1 U11094 ( .A1(n10013), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(n10012), 
        .B2(n9966), .ZN(n9967) );
  NAND2_X1 U11095 ( .A1(n9968), .A2(n9967), .ZN(P1_U3242) );
  INV_X1 U11096 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9987) );
  AOI211_X1 U11097 ( .C1(n9972), .C2(n9971), .A(n9970), .B(n9969), .ZN(n9973)
         );
  AOI21_X1 U11098 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(P1_U3084), .A(n9973), 
        .ZN(n9986) );
  AOI211_X1 U11099 ( .C1(n9976), .C2(n9975), .A(n9974), .B(n10003), .ZN(n9983)
         );
  MUX2_X1 U11100 ( .A(n9979), .B(n9978), .S(n9977), .Z(n9981) );
  OAI211_X1 U11101 ( .C1(n9981), .C2(n6302), .A(P1_U4006), .B(n9980), .ZN(
        n9982) );
  INV_X1 U11102 ( .A(n9982), .ZN(n9995) );
  AOI211_X1 U11103 ( .C1(n10012), .C2(n9984), .A(n9983), .B(n9995), .ZN(n9985)
         );
  OAI211_X1 U11104 ( .C1(n9999), .C2(n9987), .A(n9986), .B(n9985), .ZN(
        P1_U3243) );
  INV_X1 U11105 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10000) );
  XNOR2_X1 U11106 ( .A(n9989), .B(n9988), .ZN(n9993) );
  XNOR2_X1 U11107 ( .A(n9991), .B(n9990), .ZN(n9992) );
  AOI22_X1 U11108 ( .A1(n9994), .A2(n9993), .B1(n10010), .B2(n9992), .ZN(n9998) );
  AOI211_X1 U11109 ( .C1(n10012), .C2(n4889), .A(n9996), .B(n9995), .ZN(n9997)
         );
  OAI211_X1 U11110 ( .C1(n10000), .C2(n9999), .A(n9998), .B(n9997), .ZN(
        P1_U3245) );
  XNOR2_X1 U11111 ( .A(n10002), .B(n10001), .ZN(n10009) );
  AOI211_X1 U11112 ( .C1(n10006), .C2(n10005), .A(n10004), .B(n10003), .ZN(
        n10007) );
  AOI211_X1 U11113 ( .C1(n10010), .C2(n10009), .A(n10008), .B(n10007), .ZN(
        n10015) );
  AOI22_X1 U11114 ( .A1(n10013), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n10012), 
        .B2(n10011), .ZN(n10014) );
  NAND2_X1 U11115 ( .A1(n10015), .A2(n10014), .ZN(P1_U3247) );
  OAI21_X1 U11116 ( .B1(n10017), .B2(n10030), .A(n10016), .ZN(n10153) );
  OAI22_X1 U11117 ( .A1(n10153), .A2(n10019), .B1(n10018), .B2(n10031), .ZN(
        n10020) );
  INV_X1 U11118 ( .A(n10020), .ZN(n10034) );
  INV_X1 U11119 ( .A(n10042), .ZN(n10029) );
  XNOR2_X1 U11120 ( .A(n10021), .B(n10025), .ZN(n10024) );
  AOI222_X1 U11121 ( .A1(n10050), .A2(n10024), .B1(n10023), .B2(n10046), .C1(
        n10022), .C2(n10045), .ZN(n10152) );
  XNOR2_X1 U11122 ( .A(n10026), .B(n10025), .ZN(n10157) );
  NAND2_X1 U11123 ( .A1(n10157), .A2(n10027), .ZN(n10028) );
  OAI211_X1 U11124 ( .C1(n10030), .C2(n10029), .A(n10152), .B(n10028), .ZN(
        n10032) );
  NAND2_X1 U11125 ( .A1(n10032), .A2(n10031), .ZN(n10033) );
  OAI211_X1 U11126 ( .C1(n10036), .C2(n10035), .A(n10034), .B(n10033), .ZN(
        P1_U3282) );
  INV_X1 U11127 ( .A(n10037), .ZN(n10056) );
  XNOR2_X1 U11128 ( .A(n10049), .B(n10038), .ZN(n10054) );
  INV_X1 U11129 ( .A(n10054), .ZN(n10095) );
  XNOR2_X1 U11130 ( .A(n10092), .B(n10039), .ZN(n10040) );
  NAND2_X1 U11131 ( .A1(n10040), .A2(n10124), .ZN(n10091) );
  AOI22_X1 U11132 ( .A1(n5816), .A2(n10042), .B1(n10041), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n10043) );
  OAI21_X1 U11133 ( .B1(n10091), .B2(n10044), .A(n10043), .ZN(n10055) );
  AOI22_X1 U11134 ( .A1(n10046), .A2(n5785), .B1(n6441), .B2(n10045), .ZN(
        n10053) );
  OAI21_X1 U11135 ( .B1(n10049), .B2(n10048), .A(n10047), .ZN(n10051) );
  NAND2_X1 U11136 ( .A1(n10051), .A2(n10050), .ZN(n10052) );
  OAI211_X1 U11137 ( .C1(n10054), .C2(n10128), .A(n10053), .B(n10052), .ZN(
        n10093) );
  AOI211_X1 U11138 ( .C1(n10056), .C2(n10095), .A(n10055), .B(n10093), .ZN(
        n10058) );
  AOI22_X1 U11139 ( .A1(n9738), .A2(n10059), .B1(n10058), .B2(n10057), .ZN(
        P1_U3290) );
  NOR2_X1 U11140 ( .A1(n10089), .A2(n10060), .ZN(P1_U3292) );
  INV_X1 U11141 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10061) );
  NOR2_X1 U11142 ( .A1(n10089), .A2(n10061), .ZN(P1_U3293) );
  INV_X1 U11143 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10062) );
  NOR2_X1 U11144 ( .A1(n10089), .A2(n10062), .ZN(P1_U3294) );
  INV_X1 U11145 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10063) );
  NOR2_X1 U11146 ( .A1(n10089), .A2(n10063), .ZN(P1_U3295) );
  INV_X1 U11147 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10064) );
  NOR2_X1 U11148 ( .A1(n10089), .A2(n10064), .ZN(P1_U3296) );
  INV_X1 U11149 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10065) );
  NOR2_X1 U11150 ( .A1(n10089), .A2(n10065), .ZN(P1_U3297) );
  INV_X1 U11151 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10066) );
  NOR2_X1 U11152 ( .A1(n10089), .A2(n10066), .ZN(P1_U3298) );
  INV_X1 U11153 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10067) );
  NOR2_X1 U11154 ( .A1(n10089), .A2(n10067), .ZN(P1_U3299) );
  INV_X1 U11155 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10068) );
  NOR2_X1 U11156 ( .A1(n10089), .A2(n10068), .ZN(P1_U3300) );
  INV_X1 U11157 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10069) );
  NOR2_X1 U11158 ( .A1(n10089), .A2(n10069), .ZN(P1_U3301) );
  INV_X1 U11159 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10070) );
  NOR2_X1 U11160 ( .A1(n10089), .A2(n10070), .ZN(P1_U3302) );
  INV_X1 U11161 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10071) );
  NOR2_X1 U11162 ( .A1(n10089), .A2(n10071), .ZN(P1_U3303) );
  NOR2_X1 U11163 ( .A1(n10089), .A2(n10072), .ZN(P1_U3304) );
  INV_X1 U11164 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10073) );
  NOR2_X1 U11165 ( .A1(n10089), .A2(n10073), .ZN(P1_U3305) );
  INV_X1 U11166 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10074) );
  NOR2_X1 U11167 ( .A1(n10089), .A2(n10074), .ZN(P1_U3306) );
  NOR2_X1 U11168 ( .A1(n10089), .A2(n10075), .ZN(P1_U3307) );
  NOR2_X1 U11169 ( .A1(n10089), .A2(n10076), .ZN(P1_U3308) );
  INV_X1 U11170 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10077) );
  NOR2_X1 U11171 ( .A1(n10089), .A2(n10077), .ZN(P1_U3309) );
  INV_X1 U11172 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10078) );
  NOR2_X1 U11173 ( .A1(n10089), .A2(n10078), .ZN(P1_U3310) );
  INV_X1 U11174 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10079) );
  NOR2_X1 U11175 ( .A1(n10089), .A2(n10079), .ZN(P1_U3311) );
  NOR2_X1 U11176 ( .A1(n10089), .A2(n10080), .ZN(P1_U3312) );
  INV_X1 U11177 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10081) );
  NOR2_X1 U11178 ( .A1(n10089), .A2(n10081), .ZN(P1_U3313) );
  INV_X1 U11179 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10082) );
  NOR2_X1 U11180 ( .A1(n10089), .A2(n10082), .ZN(P1_U3314) );
  INV_X1 U11181 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10083) );
  NOR2_X1 U11182 ( .A1(n10089), .A2(n10083), .ZN(P1_U3315) );
  NOR2_X1 U11183 ( .A1(n10089), .A2(n10084), .ZN(P1_U3316) );
  INV_X1 U11184 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10085) );
  NOR2_X1 U11185 ( .A1(n10089), .A2(n10085), .ZN(P1_U3317) );
  INV_X1 U11186 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10086) );
  NOR2_X1 U11187 ( .A1(n10089), .A2(n10086), .ZN(P1_U3318) );
  INV_X1 U11188 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10087) );
  NOR2_X1 U11189 ( .A1(n10089), .A2(n10087), .ZN(P1_U3319) );
  INV_X1 U11190 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10088) );
  NOR2_X1 U11191 ( .A1(n10089), .A2(n10088), .ZN(P1_U3320) );
  INV_X1 U11192 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10090) );
  NOR2_X1 U11193 ( .A1(n10089), .A2(n10090), .ZN(P1_U3321) );
  OAI21_X1 U11194 ( .B1(n10092), .B2(n10136), .A(n10091), .ZN(n10094) );
  AOI211_X1 U11195 ( .C1(n10133), .C2(n10095), .A(n10094), .B(n10093), .ZN(
        n10162) );
  INV_X1 U11196 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10096) );
  AOI22_X1 U11197 ( .A1(n10160), .A2(n10162), .B1(n10096), .B2(n10158), .ZN(
        P1_U3457) );
  INV_X1 U11198 ( .A(n10097), .ZN(n10102) );
  OAI22_X1 U11199 ( .A1(n10099), .A2(n10154), .B1(n10098), .B2(n10136), .ZN(
        n10101) );
  AOI211_X1 U11200 ( .C1(n10133), .C2(n10102), .A(n10101), .B(n10100), .ZN(
        n10164) );
  AOI22_X1 U11201 ( .A1(n10160), .A2(n10164), .B1(n5771), .B2(n10158), .ZN(
        P1_U3460) );
  AOI22_X1 U11202 ( .A1(n10104), .A2(n10124), .B1(n10149), .B2(n10103), .ZN(
        n10105) );
  OAI21_X1 U11203 ( .B1(n10107), .B2(n10106), .A(n10105), .ZN(n10108) );
  NOR2_X1 U11204 ( .A1(n10109), .A2(n10108), .ZN(n10165) );
  INV_X1 U11205 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10110) );
  AOI22_X1 U11206 ( .A1(n10160), .A2(n10165), .B1(n10110), .B2(n10158), .ZN(
        P1_U3463) );
  OAI22_X1 U11207 ( .A1(n10112), .A2(n10154), .B1(n10111), .B2(n10136), .ZN(
        n10113) );
  AOI21_X1 U11208 ( .B1(n10114), .B2(n10133), .A(n10113), .ZN(n10115) );
  AND2_X1 U11209 ( .A1(n10116), .A2(n10115), .ZN(n10166) );
  INV_X1 U11210 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10117) );
  AOI22_X1 U11211 ( .A1(n10160), .A2(n10166), .B1(n10117), .B2(n10158), .ZN(
        P1_U3466) );
  AND3_X1 U11212 ( .A1(n7352), .A2(n10156), .A3(n10118), .ZN(n10121) );
  NOR2_X1 U11213 ( .A1(n10119), .A2(n10154), .ZN(n10120) );
  NOR4_X1 U11214 ( .A1(n10123), .A2(n10122), .A3(n10121), .A4(n10120), .ZN(
        n10167) );
  AOI22_X1 U11215 ( .A1(n10160), .A2(n10167), .B1(n5869), .B2(n10158), .ZN(
        P1_U3469) );
  INV_X1 U11216 ( .A(n10129), .ZN(n10132) );
  NAND2_X1 U11217 ( .A1(n10125), .A2(n10124), .ZN(n10126) );
  OAI211_X1 U11218 ( .C1(n10129), .C2(n10128), .A(n10127), .B(n10126), .ZN(
        n10130) );
  AOI211_X1 U11219 ( .C1(n10133), .C2(n10132), .A(n10131), .B(n10130), .ZN(
        n10168) );
  AOI22_X1 U11220 ( .A1(n10160), .A2(n10168), .B1(n5887), .B2(n10158), .ZN(
        P1_U3472) );
  OAI211_X1 U11221 ( .C1(n10137), .C2(n10136), .A(n10135), .B(n10134), .ZN(
        n10138) );
  AOI21_X1 U11222 ( .B1(n10156), .B2(n10139), .A(n10138), .ZN(n10169) );
  INV_X1 U11223 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10140) );
  AOI22_X1 U11224 ( .A1(n10160), .A2(n10169), .B1(n10140), .B2(n10158), .ZN(
        P1_U3475) );
  NOR2_X1 U11225 ( .A1(n10142), .A2(n10141), .ZN(n10147) );
  OAI21_X1 U11226 ( .B1(n10144), .B2(n10154), .A(n10143), .ZN(n10145) );
  AOI211_X1 U11227 ( .C1(n10147), .C2(n7480), .A(n10146), .B(n10145), .ZN(
        n10170) );
  AOI22_X1 U11228 ( .A1(n10160), .A2(n10170), .B1(n10148), .B2(n10158), .ZN(
        P1_U3478) );
  NAND2_X1 U11229 ( .A1(n10150), .A2(n10149), .ZN(n10151) );
  OAI211_X1 U11230 ( .C1(n10154), .C2(n10153), .A(n10152), .B(n10151), .ZN(
        n10155) );
  AOI21_X1 U11231 ( .B1(n10157), .B2(n10156), .A(n10155), .ZN(n10172) );
  INV_X1 U11232 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10159) );
  AOI22_X1 U11233 ( .A1(n10160), .A2(n10172), .B1(n10159), .B2(n10158), .ZN(
        P1_U3481) );
  INV_X1 U11234 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10161) );
  AOI22_X1 U11235 ( .A1(n10173), .A2(n10162), .B1(n10161), .B2(n10171), .ZN(
        P1_U3524) );
  AOI22_X1 U11236 ( .A1(n10173), .A2(n10164), .B1(n10163), .B2(n10171), .ZN(
        P1_U3525) );
  AOI22_X1 U11237 ( .A1(n10173), .A2(n10165), .B1(n5837), .B2(n10171), .ZN(
        P1_U3526) );
  AOI22_X1 U11238 ( .A1(n10173), .A2(n10166), .B1(n6797), .B2(n10171), .ZN(
        P1_U3527) );
  AOI22_X1 U11239 ( .A1(n10173), .A2(n10167), .B1(n5870), .B2(n10171), .ZN(
        P1_U3528) );
  AOI22_X1 U11240 ( .A1(n10173), .A2(n10168), .B1(n5885), .B2(n10171), .ZN(
        P1_U3529) );
  AOI22_X1 U11241 ( .A1(n10173), .A2(n10169), .B1(n5909), .B2(n10171), .ZN(
        P1_U3530) );
  AOI22_X1 U11242 ( .A1(n10173), .A2(n10170), .B1(n6803), .B2(n10171), .ZN(
        P1_U3531) );
  AOI22_X1 U11243 ( .A1(n10173), .A2(n10172), .B1(n5954), .B2(n10171), .ZN(
        P1_U3532) );
  AOI22_X1 U11244 ( .A1(n10177), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10174), .ZN(n10184) );
  AOI21_X1 U11245 ( .B1(n10176), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n10175), .ZN(
        n10183) );
  NAND2_X1 U11246 ( .A1(n10177), .A2(n4945), .ZN(n10179) );
  OAI211_X1 U11247 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n10180), .A(n10179), .B(
        n10178), .ZN(n10181) );
  NAND2_X1 U11248 ( .A1(n10181), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10182) );
  OAI211_X1 U11249 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n10184), .A(n10183), .B(
        n10182), .ZN(P2_U3245) );
  INV_X1 U11250 ( .A(n10185), .ZN(n10191) );
  INV_X1 U11251 ( .A(n10186), .ZN(n10188) );
  AOI22_X1 U11252 ( .A1(n10189), .A2(n10188), .B1(n10187), .B2(n4539), .ZN(
        n10190) );
  OAI21_X1 U11253 ( .B1(n10191), .B2(n4455), .A(n10190), .ZN(n10194) );
  INV_X1 U11254 ( .A(n10192), .ZN(n10193) );
  AOI211_X1 U11255 ( .C1(n10196), .C2(n10195), .A(n10194), .B(n10193), .ZN(
        n10197) );
  AOI22_X1 U11256 ( .A1(n10198), .A2(n6959), .B1(n10197), .B2(n9244), .ZN(
        P2_U3291) );
  AND2_X1 U11257 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10213), .ZN(P2_U3297) );
  AND2_X1 U11258 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10213), .ZN(P2_U3298) );
  AND2_X1 U11259 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10213), .ZN(P2_U3299) );
  AND2_X1 U11260 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10213), .ZN(P2_U3300) );
  NOR2_X1 U11261 ( .A1(n10210), .A2(n10201), .ZN(P2_U3301) );
  NOR2_X1 U11262 ( .A1(n10210), .A2(n10202), .ZN(P2_U3302) );
  NOR2_X1 U11263 ( .A1(n10210), .A2(n10203), .ZN(P2_U3303) );
  NOR2_X1 U11264 ( .A1(n10210), .A2(n10204), .ZN(P2_U3304) );
  AND2_X1 U11265 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10213), .ZN(P2_U3305) );
  AND2_X1 U11266 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10213), .ZN(P2_U3306) );
  AND2_X1 U11267 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10213), .ZN(P2_U3307) );
  AND2_X1 U11268 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10213), .ZN(P2_U3308) );
  NOR2_X1 U11269 ( .A1(n10210), .A2(n10205), .ZN(P2_U3309) );
  AND2_X1 U11270 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10213), .ZN(P2_U3310) );
  AND2_X1 U11271 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10213), .ZN(P2_U3311) );
  NOR2_X1 U11272 ( .A1(n10210), .A2(n10206), .ZN(P2_U3312) );
  NOR2_X1 U11273 ( .A1(n10210), .A2(n10207), .ZN(P2_U3313) );
  AND2_X1 U11274 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10213), .ZN(P2_U3314) );
  NOR2_X1 U11275 ( .A1(n10210), .A2(n10208), .ZN(P2_U3315) );
  AND2_X1 U11276 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10213), .ZN(P2_U3316) );
  NOR2_X1 U11277 ( .A1(n10210), .A2(n10209), .ZN(P2_U3317) );
  AND2_X1 U11278 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10213), .ZN(P2_U3318) );
  AND2_X1 U11279 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10213), .ZN(P2_U3319) );
  AND2_X1 U11280 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10213), .ZN(P2_U3320) );
  AND2_X1 U11281 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10213), .ZN(P2_U3321) );
  AND2_X1 U11282 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10213), .ZN(P2_U3322) );
  AND2_X1 U11283 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10213), .ZN(P2_U3323) );
  AND2_X1 U11284 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10213), .ZN(P2_U3324) );
  AND2_X1 U11285 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10213), .ZN(P2_U3325) );
  AND2_X1 U11286 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10213), .ZN(P2_U3326) );
  AOI22_X1 U11287 ( .A1(n10216), .A2(n10212), .B1(n10211), .B2(n10213), .ZN(
        P2_U3437) );
  AOI22_X1 U11288 ( .A1(n10216), .A2(n10215), .B1(n10214), .B2(n10213), .ZN(
        P2_U3438) );
  OAI22_X1 U11289 ( .A1(n10219), .A2(n10235), .B1(n10218), .B2(n10217), .ZN(
        n10220) );
  NOR2_X1 U11290 ( .A1(n10221), .A2(n10220), .ZN(n10282) );
  INV_X1 U11291 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10222) );
  AOI22_X1 U11292 ( .A1(n10281), .A2(n10282), .B1(n10222), .B2(n10279), .ZN(
        P2_U3451) );
  OAI22_X1 U11293 ( .A1(n10223), .A2(n10273), .B1(n7268), .B2(n10272), .ZN(
        n10226) );
  INV_X1 U11294 ( .A(n10224), .ZN(n10225) );
  AOI211_X1 U11295 ( .C1(n10278), .C2(n10227), .A(n10226), .B(n10225), .ZN(
        n10284) );
  INV_X1 U11296 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10228) );
  AOI22_X1 U11297 ( .A1(n10281), .A2(n10284), .B1(n10228), .B2(n10279), .ZN(
        P2_U3457) );
  AOI22_X1 U11298 ( .A1(n10232), .A2(n10231), .B1(n10230), .B2(n10229), .ZN(
        n10233) );
  OAI211_X1 U11299 ( .C1(n10236), .C2(n10235), .A(n10234), .B(n10233), .ZN(
        n10237) );
  INV_X1 U11300 ( .A(n10237), .ZN(n10285) );
  INV_X1 U11301 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10238) );
  AOI22_X1 U11302 ( .A1(n10281), .A2(n10285), .B1(n10238), .B2(n10279), .ZN(
        P2_U3469) );
  OAI22_X1 U11303 ( .A1(n10240), .A2(n10273), .B1(n10239), .B2(n10272), .ZN(
        n10242) );
  AOI211_X1 U11304 ( .C1(n10243), .C2(n10278), .A(n10242), .B(n10241), .ZN(
        n10286) );
  AOI22_X1 U11305 ( .A1(n10281), .A2(n10286), .B1(n10244), .B2(n10279), .ZN(
        P2_U3472) );
  NOR2_X1 U11306 ( .A1(n10246), .A2(n10245), .ZN(n10250) );
  OAI22_X1 U11307 ( .A1(n10248), .A2(n10273), .B1(n10247), .B2(n10272), .ZN(
        n10249) );
  NOR3_X1 U11308 ( .A1(n10251), .A2(n10250), .A3(n10249), .ZN(n10287) );
  INV_X1 U11309 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10252) );
  AOI22_X1 U11310 ( .A1(n10281), .A2(n10287), .B1(n10252), .B2(n10279), .ZN(
        P2_U3475) );
  OAI22_X1 U11311 ( .A1(n10254), .A2(n10273), .B1(n10253), .B2(n10272), .ZN(
        n10255) );
  AOI21_X1 U11312 ( .B1(n10256), .B2(n10265), .A(n10255), .ZN(n10257) );
  AND2_X1 U11313 ( .A1(n10258), .A2(n10257), .ZN(n10288) );
  AOI22_X1 U11314 ( .A1(n10281), .A2(n10288), .B1(n5247), .B2(n10279), .ZN(
        P2_U3478) );
  INV_X1 U11315 ( .A(n10259), .ZN(n10264) );
  OAI22_X1 U11316 ( .A1(n10261), .A2(n10273), .B1(n10260), .B2(n10272), .ZN(
        n10263) );
  AOI211_X1 U11317 ( .C1(n10265), .C2(n10264), .A(n10263), .B(n10262), .ZN(
        n10289) );
  AOI22_X1 U11318 ( .A1(n10281), .A2(n10289), .B1(n5278), .B2(n10279), .ZN(
        P2_U3481) );
  INV_X1 U11319 ( .A(n10266), .ZN(n10271) );
  OAI22_X1 U11320 ( .A1(n10268), .A2(n10273), .B1(n10267), .B2(n10272), .ZN(
        n10270) );
  AOI211_X1 U11321 ( .C1(n10271), .C2(n10278), .A(n10270), .B(n10269), .ZN(
        n10291) );
  AOI22_X1 U11322 ( .A1(n10281), .A2(n10291), .B1(n5304), .B2(n10279), .ZN(
        P2_U3484) );
  OAI22_X1 U11323 ( .A1(n10274), .A2(n10273), .B1(n4614), .B2(n10272), .ZN(
        n10276) );
  AOI211_X1 U11324 ( .C1(n10278), .C2(n10277), .A(n10276), .B(n10275), .ZN(
        n10293) );
  INV_X1 U11325 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10280) );
  AOI22_X1 U11326 ( .A1(n10281), .A2(n10293), .B1(n10280), .B2(n10279), .ZN(
        P2_U3487) );
  AOI22_X1 U11327 ( .A1(n4449), .A2(n10282), .B1(n4942), .B2(n10292), .ZN(
        P2_U3520) );
  AOI22_X1 U11328 ( .A1(n4449), .A2(n10284), .B1(n10283), .B2(n10292), .ZN(
        P2_U3522) );
  AOI22_X1 U11329 ( .A1(n4449), .A2(n10285), .B1(n6989), .B2(n10292), .ZN(
        P2_U3526) );
  AOI22_X1 U11330 ( .A1(n4449), .A2(n10286), .B1(n6993), .B2(n10292), .ZN(
        P2_U3527) );
  AOI22_X1 U11331 ( .A1(n4449), .A2(n10287), .B1(n6994), .B2(n10292), .ZN(
        P2_U3528) );
  AOI22_X1 U11332 ( .A1(n4449), .A2(n10288), .B1(n6998), .B2(n10292), .ZN(
        P2_U3529) );
  AOI22_X1 U11333 ( .A1(n4449), .A2(n10289), .B1(n7000), .B2(n10292), .ZN(
        P2_U3530) );
  AOI22_X1 U11334 ( .A1(n4449), .A2(n10291), .B1(n10290), .B2(n10292), .ZN(
        P2_U3531) );
  AOI22_X1 U11335 ( .A1(n4449), .A2(n10293), .B1(n7045), .B2(n10292), .ZN(
        P2_U3532) );
  INV_X1 U11336 ( .A(n10294), .ZN(n10295) );
  NAND2_X1 U11337 ( .A1(n10296), .A2(n10295), .ZN(n10297) );
  XNOR2_X1 U11338 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10297), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11339 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11340 ( .B1(n10300), .B2(n10299), .A(n10298), .ZN(ADD_1071_U56) );
  OAI21_X1 U11341 ( .B1(n10303), .B2(n10302), .A(n10301), .ZN(ADD_1071_U57) );
  OAI21_X1 U11342 ( .B1(n10306), .B2(n10305), .A(n10304), .ZN(ADD_1071_U58) );
  OAI21_X1 U11343 ( .B1(n10309), .B2(n10308), .A(n10307), .ZN(ADD_1071_U59) );
  OAI21_X1 U11344 ( .B1(n10312), .B2(n10311), .A(n10310), .ZN(ADD_1071_U60) );
  OAI21_X1 U11345 ( .B1(n10315), .B2(n10314), .A(n10313), .ZN(ADD_1071_U61) );
  AOI21_X1 U11346 ( .B1(n10318), .B2(n10317), .A(n10316), .ZN(ADD_1071_U62) );
  AOI21_X1 U11347 ( .B1(n10321), .B2(n10320), .A(n10319), .ZN(ADD_1071_U63) );
  XOR2_X1 U11348 ( .A(n10322), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11349 ( .A1(n10324), .A2(n10323), .ZN(n10326) );
  XNOR2_X1 U11350 ( .A(n10326), .B(n10325), .ZN(ADD_1071_U51) );
  OAI21_X1 U11351 ( .B1(n10329), .B2(n10328), .A(n10327), .ZN(n10330) );
  XNOR2_X1 U11352 ( .A(n10330), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11353 ( .B1(n10333), .B2(n10332), .A(n10331), .ZN(ADD_1071_U47) );
  XOR2_X1 U11354 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10334), .Z(ADD_1071_U48) );
  XOR2_X1 U11355 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10335), .Z(ADD_1071_U49) );
  XOR2_X1 U11356 ( .A(n10337), .B(n10336), .Z(ADD_1071_U54) );
  XOR2_X1 U11357 ( .A(n10339), .B(n10338), .Z(ADD_1071_U53) );
  XNOR2_X1 U11358 ( .A(n10341), .B(n10340), .ZN(ADD_1071_U52) );
  INV_X1 U6572 ( .A(n5169), .ZN(n5547) );
  NAND2_X2 U4951 ( .A1(n7422), .A2(n5079), .ZN(n5169) );
  CLKBUF_X1 U4961 ( .A(n6838), .Z(n4444) );
  CLKBUF_X2 U4965 ( .A(n5169), .Z(n5608) );
  CLKBUF_X1 U4993 ( .A(n5117), .Z(n8234) );
  BUF_X2 U5007 ( .A(n5872), .Z(n4448) );
  INV_X1 U5039 ( .A(n5128), .ZN(n4456) );
endmodule

