

module b14_C_AntiSAT_k_256_7 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064;

  CLKBUF_X1 U2479 ( .A(n3738), .Z(n2236) );
  NOR2_X1 U2480 ( .A1(n3125), .A2(U3149), .ZN(n3738) );
  CLKBUF_X1 U2481 ( .A(n3757), .Z(n2237) );
  AOI21_X1 U2482 ( .B1(n3023), .B2(n3017), .A(n4557), .ZN(n3757) );
  INV_X1 U2483 ( .A(n2846), .ZN(n2865) );
  NAND2_X1 U2484 ( .A1(n2572), .A2(n2571), .ZN(n2677) );
  NAND2_X1 U2485 ( .A1(n2648), .A2(n2650), .ZN(n2238) );
  AOI22_X1 U2486 ( .A1(n3404), .A2(n2764), .B1(n3457), .B2(n3514), .ZN(n3463)
         );
  NOR2_X2 U2487 ( .A1(n3415), .A2(n3457), .ZN(n3498) );
  OAI22_X2 U2488 ( .A1(n4120), .A2(n2807), .B1(n4128), .B2(n4293), .ZN(n4101)
         );
  AOI21_X2 U2489 ( .B1(n4147), .B2(n3851), .A(n3852), .ZN(n4120) );
  CLKBUF_X2 U2490 ( .A(n2672), .Z(n2240) );
  BUF_X2 U2491 ( .A(n2672), .Z(n2241) );
  BUF_X1 U2492 ( .A(n2672), .Z(n2242) );
  INV_X2 U2493 ( .A(n2238), .ZN(n2239) );
  NOR2_X1 U2494 ( .A1(n2639), .A2(IR_REG_29__SCAN_IN), .ZN(n2641) );
  NAND4_X1 U2495 ( .A1(n2490), .A2(n2548), .A3(n2499), .A4(n2497), .ZN(n2491)
         );
  INV_X1 U2496 ( .A(IR_REG_19__SCAN_IN), .ZN(n5040) );
  OAI21_X1 U2497 ( .B1(n2925), .B2(n4663), .A(n2378), .ZN(n2923) );
  NAND2_X2 U2498 ( .A1(n2933), .A2(n4134), .ZN(n4402) );
  INV_X2 U2499 ( .A(n4418), .ZN(U4043) );
  INV_X2 U2500 ( .A(n3627), .ZN(n3601) );
  NAND4_X1 U2501 ( .A1(n2668), .A2(n2667), .A3(n2666), .A4(n2665), .ZN(n2971)
         );
  INV_X1 U2502 ( .A(n2238), .ZN(n2244) );
  BUF_X4 U2503 ( .A(n2677), .Z(n2835) );
  AND2_X1 U2504 ( .A1(n2579), .A2(n2578), .ZN(n3928) );
  INV_X1 U2505 ( .A(n2650), .ZN(n2956) );
  NAND2_X1 U2506 ( .A1(n2642), .A2(n2960), .ZN(n2650) );
  OR2_X1 U2507 ( .A1(n2641), .A2(n2959), .ZN(n2638) );
  MUX2_X1 U2508 ( .A(IR_REG_31__SCAN_IN), .B(n2640), .S(IR_REG_29__SCAN_IN), 
        .Z(n2642) );
  AND2_X1 U2509 ( .A1(n2333), .A2(n2434), .ZN(n2573) );
  AND2_X1 U2510 ( .A1(n2489), .A2(n2488), .ZN(n2438) );
  NOR2_X2 U2511 ( .A1(n2491), .A2(IR_REG_17__SCAN_IN), .ZN(n2441) );
  INV_X1 U2512 ( .A(n2502), .ZN(n2489) );
  NAND3_X1 U2513 ( .A1(n2509), .A2(n2390), .A3(n2483), .ZN(n2502) );
  AND4_X1 U2514 ( .A1(n2487), .A2(n2486), .A3(n2485), .A4(n2484), .ZN(n2488)
         );
  INV_X1 U2515 ( .A(IR_REG_14__SCAN_IN), .ZN(n2548) );
  INV_X1 U2516 ( .A(IR_REG_4__SCAN_IN), .ZN(n2483) );
  INV_X1 U2517 ( .A(IR_REG_13__SCAN_IN), .ZN(n2497) );
  INV_X1 U2518 ( .A(IR_REG_16__SCAN_IN), .ZN(n2490) );
  NOR2_X1 U2519 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2390)
         );
  NOR2_X1 U2520 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2487)
         );
  INV_X1 U2521 ( .A(IR_REG_15__SCAN_IN), .ZN(n2499) );
  INV_X1 U2522 ( .A(IR_REG_23__SCAN_IN), .ZN(n2566) );
  INV_X1 U2523 ( .A(IR_REG_20__SCAN_IN), .ZN(n2862) );
  NOR2_X2 U2524 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2509)
         );
  NOR2_X1 U2525 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2486)
         );
  NOR2_X1 U2526 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2484)
         );
  NOR2_X1 U2527 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2485)
         );
  AND2_X4 U2528 ( .A1(n2649), .A2(n2650), .ZN(n2671) );
  AND2_X1 U2529 ( .A1(n2649), .A2(n2956), .ZN(n2672) );
  NAND2_X1 U2530 ( .A1(n2779), .A2(n2423), .ZN(n2422) );
  AOI21_X1 U2531 ( .B1(n2360), .B2(n2359), .A(n3832), .ZN(n2358) );
  INV_X1 U2532 ( .A(n2257), .ZN(n2359) );
  INV_X1 U2533 ( .A(n4103), .ZN(n4107) );
  NOR2_X1 U2534 ( .A1(n4412), .A2(n2265), .ZN(n3014) );
  OR2_X1 U2535 ( .A1(n3013), .A2(n3014), .ZN(n2309) );
  NAND2_X1 U2536 ( .A1(n3196), .A2(n2261), .ZN(n3243) );
  AND2_X1 U2537 ( .A1(n2992), .A2(n2991), .ZN(n3023) );
  INV_X1 U2538 ( .A(n2253), .ZN(n3621) );
  OR2_X1 U2539 ( .A1(n4478), .A2(n4479), .ZN(n2386) );
  NAND2_X1 U2540 ( .A1(n4545), .A2(n4546), .ZN(n4544) );
  NAND2_X1 U2541 ( .A1(n2851), .A2(n2398), .ZN(n2397) );
  NAND2_X1 U2542 ( .A1(n4258), .A2(n2850), .ZN(n2851) );
  AND2_X1 U2543 ( .A1(n2431), .A2(n2830), .ZN(n2429) );
  OAI21_X1 U2544 ( .B1(n2430), .B2(n2428), .A(n2283), .ZN(n2427) );
  INV_X1 U2545 ( .A(n2830), .ZN(n2428) );
  NOR2_X1 U2546 ( .A1(n3541), .A2(n4325), .ZN(n2778) );
  AOI21_X1 U2547 ( .B1(n2406), .B2(n2408), .A(n2281), .ZN(n2403) );
  INV_X1 U2548 ( .A(n4213), .ZN(n4189) );
  NAND2_X1 U2549 ( .A1(n2794), .A2(IR_REG_31__SCAN_IN), .ZN(n2795) );
  AND2_X1 U2550 ( .A1(n2377), .A2(n2438), .ZN(n2627) );
  AND2_X1 U2551 ( .A1(n2258), .A2(n2441), .ZN(n2377) );
  AND2_X1 U2552 ( .A1(n2564), .A2(n2565), .ZN(n2437) );
  INV_X1 U2553 ( .A(n3507), .ZN(n2452) );
  NAND2_X1 U2554 ( .A1(n2466), .A2(n2465), .ZN(n2464) );
  INV_X1 U2555 ( .A(n3742), .ZN(n2465) );
  NAND2_X1 U2556 ( .A1(n3743), .A2(n3742), .ZN(n2462) );
  INV_X2 U2557 ( .A(n3166), .ZN(n3624) );
  NAND2_X1 U2558 ( .A1(n4390), .A2(n2520), .ZN(n2521) );
  NAND2_X1 U2559 ( .A1(n4446), .A2(n2480), .ZN(n2525) );
  OAI22_X1 U2560 ( .A1(n4517), .A2(n4515), .B1(REG2_REG_13__SCAN_IN), .B2(
        n4524), .ZN(n2612) );
  NAND2_X1 U2561 ( .A1(n2385), .A2(n2294), .ZN(n2384) );
  NAND2_X1 U2562 ( .A1(n2384), .A2(n4537), .ZN(n2552) );
  NOR2_X1 U2563 ( .A1(n3956), .A2(n2555), .ZN(n2558) );
  INV_X1 U2564 ( .A(n2358), .ZN(n2356) );
  AOI21_X1 U2565 ( .B1(n2422), .B2(n2425), .A(n2787), .ZN(n2420) );
  NAND2_X1 U2566 ( .A1(n3293), .A2(n3814), .ZN(n3344) );
  NAND2_X1 U2567 ( .A1(n2922), .A2(n3920), .ZN(n3002) );
  INV_X1 U2568 ( .A(IR_REG_28__SCAN_IN), .ZN(n2625) );
  OR2_X1 U2569 ( .A1(n2591), .A2(n2568), .ZN(n2570) );
  INV_X1 U2570 ( .A(n3778), .ZN(n2362) );
  INV_X1 U2571 ( .A(IR_REG_27__SCAN_IN), .ZN(n2568) );
  NAND2_X1 U2572 ( .A1(n2573), .A2(n2566), .ZN(n2584) );
  AND2_X1 U2573 ( .A1(n2254), .A2(n2437), .ZN(n2436) );
  CLKBUF_X1 U2574 ( .A(n2438), .Z(n2434) );
  NOR2_X1 U2575 ( .A1(n2273), .A2(n2302), .ZN(n2301) );
  INV_X1 U2576 ( .A(n3423), .ZN(n2302) );
  OAI21_X1 U2577 ( .B1(n2455), .B2(n2273), .A(n3506), .ZN(n2451) );
  NAND2_X1 U2578 ( .A1(n2301), .A2(n2299), .ZN(n2298) );
  INV_X1 U2579 ( .A(n3421), .ZN(n2299) );
  OR2_X1 U2580 ( .A1(n2824), .A2(n3717), .ZN(n2831) );
  NAND2_X1 U2581 ( .A1(n2469), .A2(n2467), .ZN(n3359) );
  NOR2_X1 U2582 ( .A1(n3312), .A2(n2468), .ZN(n2467) );
  INV_X1 U2583 ( .A(n2470), .ZN(n2468) );
  NAND2_X1 U2584 ( .A1(n3524), .A2(n2471), .ZN(n2469) );
  OR2_X1 U2585 ( .A1(n3522), .A2(n3520), .ZN(n2471) );
  NAND2_X1 U2586 ( .A1(n3444), .A2(n3443), .ZN(n2454) );
  OR2_X1 U2587 ( .A1(n3444), .A2(n3443), .ZN(n2455) );
  NAND2_X1 U2588 ( .A1(n3722), .A2(n2307), .ZN(n2306) );
  NOR2_X1 U2589 ( .A1(n3673), .A2(n2308), .ZN(n2307) );
  NAND2_X1 U2590 ( .A1(n2808), .A2(REG3_REG_22__SCAN_IN), .ZN(n2817) );
  NAND2_X1 U2591 ( .A1(n2309), .A2(n2259), .ZN(n3130) );
  NOR2_X1 U2592 ( .A1(n2831), .A2(n4930), .ZN(n2844) );
  NAND2_X1 U2593 ( .A1(n3547), .A2(n3546), .ZN(n3765) );
  NAND2_X1 U2594 ( .A1(n2590), .A2(n2905), .ZN(n2998) );
  NOR2_X1 U2595 ( .A1(n2917), .A2(n2920), .ZN(n2590) );
  NAND2_X1 U2596 ( .A1(n4391), .A2(REG1_REG_3__SCAN_IN), .ZN(n4390) );
  XNOR2_X1 U2597 ( .A(n2521), .B(n4441), .ZN(n4438) );
  NAND2_X1 U2598 ( .A1(n4438), .A2(REG1_REG_4__SCAN_IN), .ZN(n4437) );
  NAND2_X1 U2599 ( .A1(n4392), .A2(n2597), .ZN(n2598) );
  XNOR2_X1 U2600 ( .A(n2525), .B(n2348), .ZN(n4459) );
  NAND2_X1 U2601 ( .A1(n4459), .A2(REG1_REG_6__SCAN_IN), .ZN(n4458) );
  NAND2_X1 U2602 ( .A1(n2386), .A2(n2263), .ZN(n2329) );
  NAND2_X1 U2603 ( .A1(n2329), .A2(n2328), .ZN(n3085) );
  INV_X1 U2604 ( .A(n3087), .ZN(n2328) );
  XNOR2_X1 U2605 ( .A(n2545), .B(n2347), .ZN(n4506) );
  NOR2_X1 U2606 ( .A1(n4495), .A2(n2389), .ZN(n2545) );
  AND2_X1 U2607 ( .A1(n2748), .A2(REG1_REG_11__SCAN_IN), .ZN(n2389) );
  OR2_X1 U2608 ( .A1(n4506), .A2(n4507), .ZN(n2388) );
  NAND2_X1 U2609 ( .A1(n4500), .A2(n2289), .ZN(n2610) );
  NAND2_X1 U2610 ( .A1(n2352), .A2(REG2_REG_14__SCAN_IN), .ZN(n2350) );
  NAND2_X1 U2611 ( .A1(n2612), .A2(n2613), .ZN(n2352) );
  NOR2_X1 U2612 ( .A1(n2612), .A2(n2613), .ZN(n2614) );
  OAI21_X1 U2613 ( .B1(n4534), .B2(n2326), .A(n2325), .ZN(n3956) );
  NAND2_X1 U2614 ( .A1(n2327), .A2(REG1_REG_14__SCAN_IN), .ZN(n2326) );
  NAND2_X1 U2615 ( .A1(n2553), .A2(n2327), .ZN(n2325) );
  INV_X1 U2616 ( .A(n3957), .ZN(n2327) );
  XNOR2_X1 U2617 ( .A(n2558), .B(n4383), .ZN(n3963) );
  NAND2_X1 U2618 ( .A1(n3963), .A2(n4951), .ZN(n3962) );
  OR2_X1 U2619 ( .A1(n2853), .A2(n4973), .ZN(n3984) );
  INV_X1 U2620 ( .A(n2396), .ZN(n2395) );
  OAI21_X1 U2621 ( .B1(n2397), .B2(n3867), .A(n2852), .ZN(n2396) );
  OR2_X1 U2622 ( .A1(n3985), .A2(n2860), .ZN(n3992) );
  INV_X1 U2623 ( .A(n3845), .ZN(n2364) );
  AOI21_X1 U2624 ( .B1(n2367), .B2(n2369), .A(n3901), .ZN(n2366) );
  OR2_X1 U2625 ( .A1(n2432), .A2(n2823), .ZN(n2430) );
  AOI21_X1 U2626 ( .B1(n4107), .B2(n2816), .A(n2274), .ZN(n2432) );
  AND2_X1 U2627 ( .A1(n2433), .A2(n2816), .ZN(n2431) );
  NAND2_X1 U2628 ( .A1(n4129), .A2(n2815), .ZN(n2816) );
  NOR2_X1 U2629 ( .A1(n2331), .A2(n4128), .ZN(n2330) );
  INV_X1 U2630 ( .A(n2332), .ZN(n2331) );
  OR2_X1 U2631 ( .A1(n4101), .A2(n4107), .ZN(n4102) );
  AOI21_X1 U2632 ( .B1(n4161), .B2(n3849), .A(n3848), .ZN(n4147) );
  AOI21_X1 U2633 ( .B1(n4209), .B2(n4194), .A(n4191), .ZN(n4161) );
  INV_X1 U2634 ( .A(n4184), .ZN(n4194) );
  AND2_X1 U2635 ( .A1(n3509), .A2(n3770), .ZN(n2337) );
  OR2_X1 U2636 ( .A1(n2424), .A2(n2422), .ZN(n2421) );
  AND4_X1 U2637 ( .A1(n2659), .A2(n2658), .A3(n2657), .A4(n2656), .ZN(n3710)
         );
  AOI21_X1 U2638 ( .B1(n2412), .B2(n2733), .A(n2266), .ZN(n2409) );
  INV_X1 U2639 ( .A(n3230), .ZN(n2416) );
  NOR2_X1 U2640 ( .A1(n3363), .A2(n3314), .ZN(n2413) );
  OR2_X1 U2641 ( .A1(n3179), .A2(n2878), .ZN(n2879) );
  OAI21_X1 U2642 ( .B1(n3111), .B2(n2875), .A(n3791), .ZN(n3095) );
  AND2_X1 U2643 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2694) );
  INV_X1 U2644 ( .A(n3031), .ZN(n2402) );
  AND2_X1 U2645 ( .A1(n2901), .A2(n2900), .ZN(n4213) );
  NOR2_X1 U2646 ( .A1(n4000), .A2(n4001), .ZN(n4230) );
  OR2_X1 U2647 ( .A1(n4022), .A2(n3994), .ZN(n4000) );
  OR2_X1 U2648 ( .A1(n4284), .A2(n3592), .ZN(n4091) );
  AND2_X1 U2649 ( .A1(n4216), .A2(n4194), .ZN(n4195) );
  NOR2_X1 U2650 ( .A1(n4315), .A2(n4215), .ZN(n4216) );
  INV_X1 U2651 ( .A(n3541), .ZN(n3770) );
  INV_X1 U2652 ( .A(n3447), .ZN(n3457) );
  OR2_X1 U2653 ( .A1(n3336), .A2(n3429), .ZN(n3415) );
  AND2_X1 U2654 ( .A1(n3074), .A2(n2922), .ZN(n4314) );
  NAND2_X1 U2655 ( .A1(n3021), .A2(n2868), .ZN(n4327) );
  XNOR2_X1 U2656 ( .A(n2863), .B(n2862), .ZN(n2922) );
  NAND2_X1 U2657 ( .A1(n2861), .A2(IR_REG_31__SCAN_IN), .ZN(n2863) );
  INV_X1 U2658 ( .A(n3237), .ZN(n3247) );
  AND2_X1 U2659 ( .A1(n3244), .A2(n3241), .ZN(n3242) );
  INV_X1 U2660 ( .A(n3934), .ZN(n3363) );
  INV_X1 U2661 ( .A(n2971), .ZN(n3024) );
  NAND2_X1 U2662 ( .A1(n2303), .A2(n3423), .ZN(n3446) );
  NAND2_X1 U2663 ( .A1(n3422), .A2(n3421), .ZN(n2303) );
  NAND2_X1 U2664 ( .A1(n3715), .A2(n2311), .ZN(n2310) );
  NAND2_X1 U2665 ( .A1(n3655), .A2(n3600), .ZN(n3715) );
  NAND2_X1 U2666 ( .A1(n2312), .A2(n3605), .ZN(n2311) );
  NAND2_X1 U2667 ( .A1(n3655), .A2(n3603), .ZN(n2312) );
  NAND2_X1 U2668 ( .A1(n3023), .A2(n3020), .ZN(n3768) );
  INV_X1 U2669 ( .A(n3710), .ZN(n4211) );
  INV_X1 U2670 ( .A(n3525), .ZN(n3255) );
  NAND2_X1 U2671 ( .A1(n4393), .A2(REG2_REG_3__SCAN_IN), .ZN(n4392) );
  XNOR2_X1 U2672 ( .A(n2598), .B(n4441), .ZN(n4436) );
  NAND2_X1 U2673 ( .A1(n4450), .A2(n4451), .ZN(n4449) );
  NOR2_X1 U2674 ( .A1(n4497), .A2(n4496), .ZN(n4495) );
  XNOR2_X1 U2675 ( .A(n2610), .B(n2347), .ZN(n4512) );
  NAND2_X1 U2676 ( .A1(n4512), .A2(REG2_REG_12__SCAN_IN), .ZN(n4511) );
  NOR2_X1 U2677 ( .A1(n4521), .A2(n4520), .ZN(n4519) );
  NAND2_X1 U2678 ( .A1(n4547), .A2(n2345), .ZN(n2630) );
  AOI21_X1 U2679 ( .B1(n2340), .B2(n2291), .A(n2341), .ZN(n3977) );
  INV_X1 U2680 ( .A(n4528), .ZN(n4551) );
  OR2_X1 U2681 ( .A1(n2786), .A2(REG1_REG_17__SCAN_IN), .ZN(n2316) );
  NAND2_X1 U2682 ( .A1(n4023), .A2(n3994), .ZN(n3995) );
  AND2_X1 U2683 ( .A1(n2869), .A2(n2918), .ZN(n3074) );
  NAND2_X1 U2684 ( .A1(n2381), .A2(n2379), .ZN(n2925) );
  INV_X1 U2685 ( .A(n4015), .ZN(n2381) );
  INV_X1 U2686 ( .A(n2380), .ZN(n2379) );
  OAI21_X1 U2687 ( .B1(n4017), .B2(n4590), .A(n2249), .ZN(n2380) );
  INV_X1 U2688 ( .A(n3537), .ZN(n3533) );
  INV_X1 U2689 ( .A(n2475), .ZN(n2473) );
  NAND2_X1 U2690 ( .A1(n2566), .A2(n2476), .ZN(n2475) );
  INV_X1 U2691 ( .A(IR_REG_24__SCAN_IN), .ZN(n2476) );
  OAI22_X1 U2692 ( .A1(n3024), .A2(n3623), .B1(n3620), .B2(n4585), .ZN(n3001)
         );
  NOR2_X1 U2693 ( .A1(n3668), .A2(n2458), .ZN(n2457) );
  INV_X1 U2694 ( .A(n2464), .ZN(n2458) );
  INV_X1 U2695 ( .A(n3568), .ZN(n2460) );
  AOI21_X1 U2696 ( .B1(n3898), .B2(n2277), .A(n2368), .ZN(n2367) );
  INV_X1 U2697 ( .A(n3903), .ZN(n2368) );
  INV_X1 U2698 ( .A(n3894), .ZN(n2370) );
  INV_X1 U2699 ( .A(n3898), .ZN(n2369) );
  NOR2_X1 U2700 ( .A1(n4206), .A2(n4079), .ZN(n4164) );
  OAI21_X1 U2701 ( .B1(n3344), .B2(n3817), .A(n3821), .ZN(n3491) );
  OAI22_X1 U2702 ( .A1(n3335), .A2(n2756), .B1(n3426), .B2(n3425), .ZN(n3404)
         );
  AOI21_X1 U2703 ( .B1(n2409), .B2(n2410), .A(n2407), .ZN(n2406) );
  INV_X1 U2704 ( .A(n2409), .ZN(n2408) );
  NOR2_X1 U2705 ( .A1(n2734), .A2(n3362), .ZN(n2742) );
  AOI21_X1 U2706 ( .B1(n2374), .B2(n3798), .A(n2373), .ZN(n2372) );
  INV_X1 U2707 ( .A(n3796), .ZN(n2374) );
  INV_X1 U2708 ( .A(n3795), .ZN(n2373) );
  OR2_X1 U2709 ( .A1(n2879), .A2(n2375), .ZN(n2371) );
  INV_X1 U2710 ( .A(n3798), .ZN(n2375) );
  NOR2_X1 U2711 ( .A1(n3562), .A2(n4292), .ZN(n2332) );
  NOR2_X1 U2712 ( .A1(n3107), .A2(n3167), .ZN(n3100) );
  OAI21_X1 U2713 ( .B1(n2872), .B2(n3075), .A(n2873), .ZN(n3036) );
  NOR2_X1 U2714 ( .A1(n2475), .A2(IR_REG_25__SCAN_IN), .ZN(n2474) );
  INV_X1 U2715 ( .A(n2491), .ZN(n2443) );
  OR2_X1 U2716 ( .A1(n2537), .A2(IR_REG_10__SCAN_IN), .ZN(n2506) );
  INV_X1 U2717 ( .A(IR_REG_9__SCAN_IN), .ZN(n4843) );
  AND2_X1 U2718 ( .A1(n3658), .A2(n3657), .ZN(n3595) );
  INV_X1 U2719 ( .A(n3132), .ZN(n3156) );
  NAND2_X1 U2720 ( .A1(n3741), .A2(n2464), .ZN(n2463) );
  AND2_X1 U2721 ( .A1(n3564), .A2(n3563), .ZN(n3565) );
  AND2_X1 U2722 ( .A1(n3003), .A2(n3002), .ZN(n3627) );
  INV_X1 U2723 ( .A(n3018), .ZN(n3003) );
  INV_X1 U2724 ( .A(n3283), .ZN(n3526) );
  AND2_X1 U2725 ( .A1(n2742), .A2(REG3_REG_11__SCAN_IN), .ZN(n2749) );
  NAND2_X1 U2726 ( .A1(n2447), .A2(n3605), .ZN(n2446) );
  INV_X1 U2727 ( .A(n3603), .ZN(n2447) );
  AND2_X1 U2728 ( .A1(n3603), .A2(n3604), .ZN(n3600) );
  OR2_X1 U2729 ( .A1(n2817), .A2(n3659), .ZN(n2824) );
  NAND2_X1 U2730 ( .A1(n3522), .A2(n3520), .ZN(n2470) );
  INV_X1 U2731 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2726) );
  OR2_X1 U2732 ( .A1(n2727), .A2(n2726), .ZN(n2734) );
  NAND2_X1 U2733 ( .A1(n2456), .A2(n2459), .ZN(n3723) );
  AOI21_X1 U2734 ( .B1(n3567), .B2(n2461), .A(n2460), .ZN(n2459) );
  NAND2_X1 U2735 ( .A1(n3741), .A2(n2457), .ZN(n2456) );
  INV_X1 U2736 ( .A(n2462), .ZN(n2461) );
  AND2_X1 U2737 ( .A1(n3454), .A2(n3453), .ZN(n3507) );
  NAND2_X1 U2738 ( .A1(n2749), .A2(REG3_REG_12__SCAN_IN), .ZN(n2757) );
  INV_X1 U2739 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4836) );
  INV_X1 U2740 ( .A(n3264), .ZN(n3206) );
  OR2_X1 U2741 ( .A1(n2757), .A2(n4836), .ZN(n2772) );
  AND2_X1 U2742 ( .A1(n3928), .A2(n3980), .ZN(n3018) );
  NAND2_X1 U2743 ( .A1(n2509), .A2(n2516), .ZN(n2510) );
  INV_X1 U2744 ( .A(IR_REG_3__SCAN_IN), .ZN(n2512) );
  XNOR2_X1 U2745 ( .A(n2519), .B(n2346), .ZN(n4391) );
  NAND2_X1 U2746 ( .A1(n4437), .A2(n2522), .ZN(n4447) );
  NAND2_X1 U2747 ( .A1(n4449), .A2(n2278), .ZN(n2601) );
  NAND2_X1 U2748 ( .A1(n2315), .A2(n2313), .ZN(n2530) );
  NAND2_X1 U2749 ( .A1(n4476), .A2(n2314), .ZN(n2313) );
  NAND2_X1 U2750 ( .A1(n4458), .A2(n2247), .ZN(n2315) );
  AND2_X1 U2751 ( .A1(n3085), .A2(n2536), .ZN(n2539) );
  NAND2_X1 U2752 ( .A1(n2382), .A2(n2552), .ZN(n4534) );
  NAND2_X1 U2753 ( .A1(n2383), .A2(n2613), .ZN(n2382) );
  AND2_X1 U2754 ( .A1(n2349), .A2(n2350), .ZN(n3953) );
  NOR2_X1 U2755 ( .A1(n4534), .A2(n4533), .ZN(n4532) );
  NAND2_X1 U2756 ( .A1(n3962), .A2(n2559), .ZN(n4545) );
  NAND2_X1 U2757 ( .A1(n4382), .A2(REG2_REG_18__SCAN_IN), .ZN(n2344) );
  INV_X1 U2758 ( .A(n2629), .ZN(n2343) );
  INV_X1 U2759 ( .A(n3974), .ZN(n2324) );
  OAI21_X1 U2760 ( .B1(n2251), .B2(n2323), .A(n2322), .ZN(n2321) );
  NOR2_X1 U2761 ( .A1(n2295), .A2(n2324), .ZN(n2323) );
  NAND2_X1 U2762 ( .A1(n2251), .A2(n3974), .ZN(n2322) );
  AND2_X1 U2763 ( .A1(n2394), .A2(n3992), .ZN(n2393) );
  NAND2_X1 U2764 ( .A1(n2395), .A2(n2397), .ZN(n2394) );
  NAND2_X1 U2765 ( .A1(n2354), .A2(n2353), .ZN(n3987) );
  AOI21_X1 U2766 ( .B1(n2355), .B2(n2361), .A(n3909), .ZN(n2353) );
  NOR2_X1 U2767 ( .A1(n4019), .A2(n2356), .ZN(n2355) );
  INV_X1 U2768 ( .A(n4264), .ZN(n4087) );
  OR2_X1 U2769 ( .A1(n2814), .A2(n3901), .ZN(n4103) );
  AND2_X1 U2770 ( .A1(n2801), .A2(n2800), .ZN(n2808) );
  NAND2_X1 U2771 ( .A1(n2419), .A2(n2417), .ZN(n4192) );
  AOI21_X1 U2772 ( .B1(n2420), .B2(n2418), .A(n2284), .ZN(n2417) );
  INV_X1 U2773 ( .A(n2425), .ZN(n2418) );
  NAND2_X1 U2774 ( .A1(n2887), .A2(n3894), .ZN(n4206) );
  AND4_X1 U2775 ( .A1(n2654), .A2(n2653), .A3(n2652), .A4(n2651), .ZN(n4209)
         );
  INV_X1 U2776 ( .A(n4636), .ZN(n3426) );
  INV_X1 U2777 ( .A(n4633), .ZN(n3384) );
  NAND2_X1 U2778 ( .A1(n2881), .A2(n3812), .ZN(n3293) );
  NAND2_X1 U2779 ( .A1(n2371), .A2(n2372), .ZN(n3225) );
  INV_X1 U2780 ( .A(n3249), .ZN(n3313) );
  OAI21_X1 U2781 ( .B1(n3095), .B2(n3093), .A(n3802), .ZN(n3254) );
  OR2_X1 U2782 ( .A1(n3106), .A2(n3140), .ZN(n3107) );
  NAND2_X1 U2783 ( .A1(n2874), .A2(n3787), .ZN(n3111) );
  NAND2_X1 U2784 ( .A1(n2376), .A2(n3782), .ZN(n3064) );
  NAND2_X1 U2785 ( .A1(n3036), .A2(n3035), .ZN(n2376) );
  NAND2_X1 U2786 ( .A1(n4592), .A2(n4585), .ZN(n3044) );
  CLKBUF_X1 U2787 ( .A(n2871), .Z(n2872) );
  NAND2_X1 U2788 ( .A1(n4036), .A2(n2850), .ZN(n4022) );
  NAND2_X1 U2789 ( .A1(n2357), .A2(n2358), .ZN(n4020) );
  OR2_X1 U2790 ( .A1(n2897), .A2(n2361), .ZN(n2357) );
  NOR2_X1 U2791 ( .A1(n4091), .A2(n2338), .ZN(n4036) );
  NAND2_X1 U2792 ( .A1(n2339), .A2(n4072), .ZN(n2338) );
  NOR2_X1 U2793 ( .A1(n4255), .A2(n4263), .ZN(n2339) );
  NOR3_X1 U2794 ( .A1(n4091), .A2(n4272), .A3(n4263), .ZN(n4048) );
  INV_X1 U2795 ( .A(n4052), .ZN(n4263) );
  NAND2_X1 U2796 ( .A1(n4195), .A2(n2332), .ZN(n4148) );
  NAND2_X1 U2797 ( .A1(n4195), .A2(n4176), .ZN(n4175) );
  NAND2_X1 U2798 ( .A1(n3498), .A2(n2337), .ZN(n3483) );
  AND2_X1 U2799 ( .A1(n3498), .A2(n3509), .ZN(n3496) );
  NAND2_X1 U2800 ( .A1(n3295), .A2(n3384), .ZN(n3336) );
  AND4_X1 U2801 ( .A1(n2747), .A2(n2746), .A3(n2745), .A4(n2744), .ZN(n3393)
         );
  INV_X1 U2802 ( .A(n3429), .ZN(n3425) );
  NAND2_X1 U2803 ( .A1(n2336), .A2(n3314), .ZN(n3274) );
  MUX2_X1 U2804 ( .A(n2740), .B(DATAI_10_), .S(n2835), .Z(n3356) );
  NOR2_X1 U2805 ( .A1(n3274), .A2(n3356), .ZN(n3295) );
  NAND2_X1 U2806 ( .A1(n3183), .A2(n3247), .ZN(n3212) );
  AND2_X1 U2807 ( .A1(n4415), .A2(n2868), .ZN(n4635) );
  MUX2_X1 U2808 ( .A(n4457), .B(DATAI_6_), .S(n2835), .Z(n3264) );
  NOR2_X1 U2809 ( .A1(n3044), .A2(n3059), .ZN(n4602) );
  INV_X1 U2810 ( .A(n4635), .ZN(n4594) );
  AND2_X1 U2811 ( .A1(n2931), .A2(n2919), .ZN(n2924) );
  NAND2_X1 U2812 ( .A1(n2584), .A2(IR_REG_31__SCAN_IN), .ZN(n2585) );
  AND2_X1 U2813 ( .A1(n2436), .A2(n2441), .ZN(n2333) );
  INV_X1 U2814 ( .A(n2441), .ZN(n2439) );
  NAND2_X1 U2815 ( .A1(n2434), .A2(n2435), .ZN(n2440) );
  AND2_X1 U2816 ( .A1(n2254), .A2(n2564), .ZN(n2435) );
  NAND2_X1 U2817 ( .A1(n2795), .A2(n5040), .ZN(n2861) );
  NOR2_X1 U2818 ( .A1(n2491), .A2(IR_REG_17__SCAN_IN), .ZN(n2442) );
  INV_X1 U2819 ( .A(IR_REG_7__SCAN_IN), .ZN(n4844) );
  INV_X1 U2820 ( .A(IR_REG_2__SCAN_IN), .ZN(n2516) );
  INV_X1 U2821 ( .A(n2301), .ZN(n2300) );
  AND2_X1 U2822 ( .A1(n2450), .A2(n2298), .ZN(n2297) );
  INV_X1 U2823 ( .A(n2451), .ZN(n2450) );
  NOR2_X1 U2824 ( .A1(n3735), .A2(n2305), .ZN(n2304) );
  INV_X1 U2825 ( .A(n3674), .ZN(n2305) );
  NAND2_X1 U2826 ( .A1(n3359), .A2(n3358), .ZN(n3381) );
  NAND2_X1 U2827 ( .A1(n3130), .A2(n3129), .ZN(n3153) );
  OR2_X1 U2828 ( .A1(n3128), .A2(n3127), .ZN(n3129) );
  AND2_X1 U2829 ( .A1(n3984), .A2(n2854), .ZN(n4009) );
  NAND2_X1 U2830 ( .A1(n3308), .A2(n3307), .ZN(n3524) );
  OAI21_X1 U2831 ( .B1(n2677), .B2(n2945), .A(n2664), .ZN(n3026) );
  NAND2_X1 U2832 ( .A1(n2677), .A2(DATAI_1_), .ZN(n2664) );
  INV_X1 U2833 ( .A(n4132), .ZN(n4128) );
  NAND2_X1 U2834 ( .A1(n2449), .A2(n2444), .ZN(n3688) );
  INV_X1 U2835 ( .A(n2445), .ZN(n2444) );
  NAND2_X1 U2836 ( .A1(n3656), .A2(n2280), .ZN(n2449) );
  OAI21_X1 U2837 ( .B1(n3600), .B2(n2448), .A(n2446), .ZN(n2445) );
  AND4_X1 U2838 ( .A1(n2691), .A2(n2690), .A3(n2689), .A4(n2688), .ZN(n3171)
         );
  NAND2_X1 U2839 ( .A1(n3169), .A2(n3168), .ZN(n3196) );
  OR2_X1 U2840 ( .A1(n3551), .A2(n3550), .ZN(n3552) );
  NAND2_X1 U2841 ( .A1(n2469), .A2(n2470), .ZN(n3311) );
  NAND2_X1 U2842 ( .A1(n3446), .A2(n2455), .ZN(n2453) );
  NAND2_X1 U2843 ( .A1(n2306), .A2(n3674), .ZN(n3734) );
  AND2_X1 U2844 ( .A1(n2309), .A2(n2255), .ZN(n3055) );
  INV_X1 U2845 ( .A(n3775), .ZN(n4667) );
  AND4_X1 U2846 ( .A1(n2714), .A2(n2713), .A3(n2712), .A4(n2711), .ZN(n3525)
         );
  NAND2_X1 U2847 ( .A1(n3023), .A2(n3022), .ZN(n3760) );
  INV_X1 U2848 ( .A(n3760), .ZN(n4669) );
  NAND2_X1 U2849 ( .A1(n2841), .A2(n2840), .ZN(n4251) );
  AND3_X1 U2850 ( .A1(n2839), .A2(n2838), .A3(n2837), .ZN(n2840) );
  INV_X1 U2851 ( .A(n4328), .ZN(n3514) );
  INV_X1 U2852 ( .A(n3393), .ZN(n3428) );
  INV_X1 U2853 ( .A(n3171), .ZN(n3937) );
  OR2_X1 U2854 ( .A1(n2846), .A2(REG3_REG_3__SCAN_IN), .ZN(n2685) );
  NAND4_X2 U2855 ( .A1(n2663), .A2(n2662), .A3(n2661), .A4(n2660), .ZN(n2669)
         );
  XNOR2_X1 U2856 ( .A(n2518), .B(IR_REG_1__SCAN_IN), .ZN(n3945) );
  XNOR2_X1 U2857 ( .A(n2596), .B(n2346), .ZN(n4393) );
  NAND2_X1 U2858 ( .A1(n4435), .A2(n2599), .ZN(n4450) );
  XNOR2_X1 U2859 ( .A(n2601), .B(n2348), .ZN(n4461) );
  NAND2_X1 U2860 ( .A1(n4458), .A2(n2526), .ZN(n4467) );
  XNOR2_X1 U2861 ( .A(n2530), .B(n4580), .ZN(n4478) );
  INV_X1 U2862 ( .A(n2386), .ZN(n4477) );
  INV_X1 U2863 ( .A(n2329), .ZN(n3088) );
  XNOR2_X1 U2864 ( .A(n2539), .B(n4579), .ZN(n4487) );
  INV_X1 U2865 ( .A(n2388), .ZN(n4505) );
  AND2_X1 U2866 ( .A1(n2388), .A2(n2268), .ZN(n4521) );
  NAND2_X1 U2867 ( .A1(n4511), .A2(n2611), .ZN(n4517) );
  OR2_X1 U2868 ( .A1(n2614), .A2(n2351), .ZN(n4530) );
  INV_X1 U2869 ( .A(n2352), .ZN(n2351) );
  NOR2_X1 U2870 ( .A1(n4531), .A2(n2293), .ZN(n2318) );
  NAND2_X1 U2871 ( .A1(n2321), .A2(n2296), .ZN(n2320) );
  NAND2_X1 U2872 ( .A1(n2392), .A2(n2395), .ZN(n3993) );
  NAND2_X1 U2873 ( .A1(n2363), .A2(n3872), .ZN(n4032) );
  NAND2_X1 U2874 ( .A1(n2897), .A2(n2257), .ZN(n2363) );
  NAND2_X1 U2875 ( .A1(n2897), .A2(n3845), .ZN(n4054) );
  NAND2_X1 U2876 ( .A1(n2426), .A2(n2430), .ZN(n4063) );
  NAND2_X1 U2877 ( .A1(n4101), .A2(n2431), .ZN(n2426) );
  NAND2_X1 U2878 ( .A1(n4102), .A2(n2816), .ZN(n4077) );
  NAND2_X1 U2879 ( .A1(n4195), .A2(n2288), .ZN(n4284) );
  AND2_X1 U2880 ( .A1(n2421), .A2(n2425), .ZN(n4205) );
  NAND2_X1 U2881 ( .A1(n3498), .A2(n2290), .ZN(n4315) );
  INV_X1 U2882 ( .A(n2421), .ZN(n3480) );
  INV_X1 U2883 ( .A(n4324), .ZN(n3509) );
  NAND2_X1 U2884 ( .A1(n2405), .A2(n2409), .ZN(n3292) );
  NAND2_X1 U2885 ( .A1(n3230), .A2(n2412), .ZN(n2405) );
  NAND2_X1 U2886 ( .A1(n2414), .A2(n2411), .ZN(n3273) );
  INV_X1 U2887 ( .A(n2413), .ZN(n2411) );
  NAND2_X1 U2888 ( .A1(n2416), .A2(n2415), .ZN(n2414) );
  NAND2_X1 U2889 ( .A1(n2879), .A2(n3796), .ZN(n3219) );
  AND2_X1 U2890 ( .A1(n4402), .A2(n2936), .ZN(n4201) );
  NAND2_X1 U2891 ( .A1(n3030), .A2(n2681), .ZN(n3063) );
  INV_X1 U2892 ( .A(n4134), .ZN(n4557) );
  OR2_X1 U2893 ( .A1(n3016), .A2(n2932), .ZN(n4134) );
  INV_X1 U2894 ( .A(n4560), .ZN(n4220) );
  INV_X1 U2895 ( .A(n3026), .ZN(n4592) );
  MUX2_X1 U2896 ( .A(n2335), .B(n2334), .S(n2677), .Z(n4585) );
  AOI21_X1 U2897 ( .B1(n4234), .B2(n4233), .A(n4232), .ZN(n4403) );
  AOI211_X1 U2898 ( .C1(n4314), .C2(n4244), .A(n4243), .B(n4242), .ZN(n4245)
         );
  AND2_X2 U2899 ( .A1(n2924), .A2(n2929), .ZN(n4649) );
  NAND2_X1 U2900 ( .A1(n2964), .A2(n3009), .ZN(n4570) );
  INV_X1 U2901 ( .A(n4415), .ZN(n3021) );
  XNOR2_X1 U2902 ( .A(n2580), .B(IR_REG_21__SCAN_IN), .ZN(n3920) );
  AND2_X1 U2903 ( .A1(n2556), .A2(n2501), .ZN(n3950) );
  INV_X1 U2904 ( .A(n2699), .ZN(n4583) );
  XNOR2_X1 U2905 ( .A(n2517), .B(n2516), .ZN(n4434) );
  OR2_X1 U2906 ( .A1(n2509), .A2(n2959), .ZN(n2517) );
  XNOR2_X1 U2907 ( .A(n2310), .B(n2448), .ZN(n3721) );
  OAI211_X1 U2908 ( .C1(n2245), .C2(n2295), .A(n3975), .B(n4553), .ZN(n2387)
         );
  NAND2_X1 U2909 ( .A1(n4553), .A2(n2320), .ZN(n2319) );
  NAND2_X1 U2910 ( .A1(n2245), .A2(n2318), .ZN(n2317) );
  NAND2_X1 U2911 ( .A1(n4663), .A2(n4943), .ZN(n2378) );
  AND2_X1 U2912 ( .A1(n2998), .A2(n3002), .ZN(n3131) );
  AND2_X1 U2913 ( .A1(n4544), .A2(n2316), .ZN(n2245) );
  INV_X1 U2914 ( .A(n2361), .ZN(n2360) );
  NAND2_X1 U2915 ( .A1(n3872), .A2(n2362), .ZN(n2361) );
  INV_X1 U2916 ( .A(n2733), .ZN(n2415) );
  AND3_X1 U2917 ( .A1(n2436), .A2(n2270), .A3(n2441), .ZN(n2246) );
  NAND2_X1 U2918 ( .A1(n2463), .A2(n2462), .ZN(n3666) );
  AND2_X1 U2919 ( .A1(n2526), .A2(n2279), .ZN(n2247) );
  AND2_X1 U2920 ( .A1(n4547), .A2(n2291), .ZN(n2248) );
  AND2_X2 U2921 ( .A1(n2998), .A2(n2997), .ZN(n2253) );
  INV_X1 U2922 ( .A(n3227), .ZN(n3314) );
  NAND2_X1 U2923 ( .A1(n2489), .A2(n2488), .ZN(n2496) );
  NOR2_X1 U2924 ( .A1(n2285), .A2(n2903), .ZN(n2249) );
  AND2_X1 U2925 ( .A1(n2372), .A2(n2287), .ZN(n2250) );
  INV_X1 U2926 ( .A(n2291), .ZN(n2342) );
  XOR2_X1 U2927 ( .A(n3980), .B(REG1_REG_19__SCAN_IN), .Z(n2251) );
  NAND2_X1 U2928 ( .A1(n2251), .A2(n2295), .ZN(n2252) );
  AND3_X1 U2929 ( .A1(n5040), .A2(n2562), .A3(n2862), .ZN(n2254) );
  NAND2_X1 U2930 ( .A1(n3053), .A2(n3052), .ZN(n2255) );
  OR2_X1 U2931 ( .A1(n3938), .A2(n3132), .ZN(n2256) );
  NOR2_X1 U2932 ( .A1(n2898), .A2(n2364), .ZN(n2257) );
  XNOR2_X1 U2933 ( .A(n2638), .B(IR_REG_30__SCAN_IN), .ZN(n2648) );
  AOI21_X1 U2934 ( .B1(n3688), .B2(n3684), .A(n3686), .ZN(n3752) );
  AND2_X1 U2935 ( .A1(n2515), .A2(n2514), .ZN(n4389) );
  INV_X1 U2936 ( .A(n4389), .ZN(n2346) );
  AND3_X1 U2937 ( .A1(n2254), .A2(n2473), .A3(n2437), .ZN(n2258) );
  AND2_X1 U2938 ( .A1(n3056), .A2(n2255), .ZN(n2259) );
  NOR2_X1 U2939 ( .A1(n4532), .A2(n2553), .ZN(n2260) );
  AND2_X1 U2940 ( .A1(n3195), .A2(n2292), .ZN(n2261) );
  AND2_X1 U2941 ( .A1(n2648), .A2(n2956), .ZN(n2262) );
  OR2_X1 U2942 ( .A1(n4580), .A2(n2530), .ZN(n2263) );
  NOR2_X1 U2943 ( .A1(n2637), .A2(n2636), .ZN(n2264) );
  INV_X1 U2944 ( .A(IR_REG_26__SCAN_IN), .ZN(n4842) );
  AND2_X1 U2945 ( .A1(n3004), .A2(n3627), .ZN(n2265) );
  AND2_X1 U2946 ( .A1(n3383), .A2(n3364), .ZN(n2266) );
  INV_X1 U2947 ( .A(IR_REG_25__SCAN_IN), .ZN(n2567) );
  OR2_X1 U2948 ( .A1(n2440), .A2(n2439), .ZN(n2267) );
  NAND2_X1 U2949 ( .A1(n2306), .A2(n2304), .ZN(n3656) );
  AND2_X1 U2950 ( .A1(n4258), .A2(n2899), .ZN(n3909) );
  OR2_X1 U2951 ( .A1(n2545), .A2(n2347), .ZN(n2268) );
  AND3_X1 U2952 ( .A1(n2489), .A2(n2488), .A3(n2254), .ZN(n2269) );
  AND2_X1 U2953 ( .A1(n2474), .A2(n4842), .ZN(n2270) );
  NAND2_X1 U2954 ( .A1(n2269), .A2(n2441), .ZN(n2271) );
  INV_X1 U2955 ( .A(IR_REG_31__SCAN_IN), .ZN(n2959) );
  INV_X1 U2956 ( .A(n4457), .ZN(n2348) );
  NAND2_X1 U2957 ( .A1(n4211), .A2(n3482), .ZN(n2425) );
  INV_X1 U2958 ( .A(n3716), .ZN(n2448) );
  NAND2_X1 U2959 ( .A1(n4195), .A2(n2330), .ZN(n2272) );
  NAND2_X1 U2960 ( .A1(n2454), .A2(n2452), .ZN(n2273) );
  OAI21_X1 U2961 ( .B1(n3422), .B2(n2300), .A(n2297), .ZN(n3535) );
  NAND2_X1 U2962 ( .A1(n2453), .A2(n2454), .ZN(n3508) );
  AND2_X1 U2963 ( .A1(n4276), .A2(n4092), .ZN(n2274) );
  AND3_X1 U2964 ( .A1(n2489), .A2(n2488), .A3(n2443), .ZN(n2494) );
  OR2_X1 U2965 ( .A1(n3716), .A2(n3605), .ZN(n2275) );
  OR2_X1 U2966 ( .A1(n4091), .A2(n4272), .ZN(n2276) );
  INV_X1 U2967 ( .A(n3668), .ZN(n3567) );
  OR2_X1 U2968 ( .A1(n3893), .A2(n2370), .ZN(n2277) );
  INV_X1 U2969 ( .A(n3743), .ZN(n2466) );
  OR2_X1 U2970 ( .A1(n4583), .A2(n2600), .ZN(n2278) );
  NAND2_X1 U2971 ( .A1(n4581), .A2(REG1_REG_7__SCAN_IN), .ZN(n2279) );
  AND2_X1 U2972 ( .A1(n2275), .A2(n3595), .ZN(n2280) );
  AND2_X1 U2973 ( .A1(n3393), .A2(n3384), .ZN(n2281) );
  AND2_X1 U2974 ( .A1(n3666), .A2(n3567), .ZN(n2282) );
  NAND2_X1 U2975 ( .A1(n4087), .A2(n4072), .ZN(n2283) );
  NOR2_X1 U2976 ( .A1(n4187), .A2(n4208), .ZN(n2284) );
  AND2_X1 U2977 ( .A1(n4038), .A2(n4637), .ZN(n2285) );
  INV_X1 U2978 ( .A(n3869), .ZN(n2398) );
  NOR2_X1 U2979 ( .A1(n2350), .A2(n2614), .ZN(n2286) );
  INV_X1 U2980 ( .A(n2823), .ZN(n2433) );
  NOR2_X1 U2981 ( .A1(n4276), .A2(n4092), .ZN(n2823) );
  XNOR2_X1 U2982 ( .A(n2589), .B(IR_REG_26__SCAN_IN), .ZN(n2905) );
  INV_X1 U2983 ( .A(n2755), .ZN(n2347) );
  AND2_X1 U2984 ( .A1(n3892), .A2(n3894), .ZN(n3481) );
  INV_X1 U2985 ( .A(n3481), .ZN(n2423) );
  OAI22_X1 U2986 ( .A1(n3099), .A2(n2700), .B1(n3167), .B2(n3936), .ZN(n3253)
         );
  NAND2_X1 U2987 ( .A1(n2404), .A2(n2403), .ZN(n3335) );
  NAND2_X1 U2988 ( .A1(n3934), .A2(n3314), .ZN(n2287) );
  OAI21_X1 U2989 ( .B1(n3253), .B2(n2706), .A(n2705), .ZN(n3177) );
  OAI21_X1 U2990 ( .B1(n3211), .B2(n2725), .A(n2724), .ZN(n3230) );
  MUX2_X1 U2991 ( .A(n3980), .B(n4981), .S(n2835), .Z(n4176) );
  INV_X1 U2992 ( .A(n3855), .ZN(n2407) );
  AND2_X1 U2993 ( .A1(n2330), .A2(n4112), .ZN(n2288) );
  INV_X1 U2994 ( .A(n2336), .ZN(n3231) );
  NOR2_X1 U2995 ( .A1(n3212), .A2(n3283), .ZN(n2336) );
  NAND2_X1 U2996 ( .A1(n3196), .A2(n3195), .ZN(n3202) );
  INV_X1 U2997 ( .A(n2412), .ZN(n2410) );
  NOR2_X1 U2998 ( .A1(n2413), .A2(n2741), .ZN(n2412) );
  OR2_X1 U2999 ( .A1(n4577), .A2(n2609), .ZN(n2289) );
  AND2_X1 U3000 ( .A1(n2337), .A2(n3700), .ZN(n2290) );
  NAND2_X1 U3001 ( .A1(n2402), .A2(n2679), .ZN(n3030) );
  AND2_X2 U3002 ( .A1(n2924), .A2(n2991), .ZN(n4666) );
  INV_X1 U3003 ( .A(n4666), .ZN(n4663) );
  AND2_X1 U3004 ( .A1(n2345), .A2(n2343), .ZN(n2291) );
  INV_X1 U3005 ( .A(n4042), .ZN(n4255) );
  NAND2_X1 U3006 ( .A1(n2472), .A2(IR_REG_31__SCAN_IN), .ZN(n2591) );
  AND2_X1 U3007 ( .A1(n3100), .A2(n3206), .ZN(n3183) );
  AND2_X1 U3008 ( .A1(n2835), .A2(DATAI_27_), .ZN(n2899) );
  OR2_X1 U3009 ( .A1(n3201), .A2(n3200), .ZN(n2292) );
  INV_X1 U3010 ( .A(n2613), .ZN(n4537) );
  AND2_X1 U3011 ( .A1(n2321), .A2(n2252), .ZN(n2293) );
  NAND2_X1 U3012 ( .A1(n4524), .A2(REG1_REG_13__SCAN_IN), .ZN(n2294) );
  OAI21_X1 U3013 ( .B1(n4549), .B2(n2342), .A(n2344), .ZN(n2341) );
  INV_X1 U3014 ( .A(IR_REG_0__SCAN_IN), .ZN(n2335) );
  INV_X1 U3015 ( .A(DATAI_0_), .ZN(n2334) );
  INV_X1 U3016 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2314) );
  AND2_X1 U3017 ( .A1(n3974), .A2(n2561), .ZN(n2295) );
  OR2_X1 U3018 ( .A1(n2251), .A2(n2324), .ZN(n2296) );
  NAND2_X1 U3019 ( .A1(n3535), .A2(n3534), .ZN(n3539) );
  NAND2_X1 U3020 ( .A1(n3722), .A2(n3726), .ZN(n3678) );
  INV_X1 U3021 ( .A(n3726), .ZN(n2308) );
  INV_X1 U3022 ( .A(n2309), .ZN(n3054) );
  INV_X2 U3023 ( .A(n3131), .ZN(n3620) );
  AND2_X2 U3024 ( .A1(n3000), .A2(n3131), .ZN(n3166) );
  OAI211_X1 U3025 ( .C1(n2245), .C2(n2319), .A(n2317), .B(n3983), .ZN(U3259)
         );
  NAND2_X1 U3026 ( .A1(n2245), .A2(n2295), .ZN(n3975) );
  NAND2_X1 U3027 ( .A1(n2434), .A2(n2246), .ZN(n2472) );
  NAND2_X1 U3028 ( .A1(n2573), .A2(n2474), .ZN(n2588) );
  INV_X1 U3029 ( .A(n4585), .ZN(n4670) );
  NAND2_X1 U3030 ( .A1(n4548), .A2(n4549), .ZN(n4547) );
  INV_X1 U3031 ( .A(n4548), .ZN(n2340) );
  OR2_X1 U3032 ( .A1(n2786), .A2(REG2_REG_17__SCAN_IN), .ZN(n2345) );
  INV_X1 U3033 ( .A(n2614), .ZN(n2349) );
  INV_X1 U3034 ( .A(n2384), .ZN(n2383) );
  NOR2_X1 U3035 ( .A1(n4488), .A2(n4487), .ZN(n4486) );
  NOR2_X1 U3036 ( .A1(n3951), .A2(n2616), .ZN(n2618) );
  NOR2_X1 U3037 ( .A1(n3952), .A2(n3953), .ZN(n3951) );
  XNOR2_X1 U3038 ( .A(n2618), .B(n4383), .ZN(n3968) );
  NAND2_X1 U3039 ( .A1(n2264), .A2(n2387), .ZN(U3258) );
  NAND2_X1 U3040 ( .A1(n4447), .A2(n4448), .ZN(n4446) );
  INV_X1 U3041 ( .A(n4519), .ZN(n2385) );
  INV_X2 U3042 ( .A(n2669), .ZN(n3076) );
  NAND2_X1 U3043 ( .A1(n2873), .A2(n3779), .ZN(n2871) );
  NAND2_X1 U3044 ( .A1(n2669), .A2(n4592), .ZN(n3779) );
  NAND2_X1 U3045 ( .A1(n2897), .A2(n2355), .ZN(n2354) );
  NAND2_X1 U3046 ( .A1(n2365), .A2(n2366), .ZN(n2896) );
  NAND2_X1 U3047 ( .A1(n2887), .A2(n2367), .ZN(n2365) );
  NAND2_X1 U3048 ( .A1(n2371), .A2(n2250), .ZN(n2880) );
  NAND4_X1 U3049 ( .A1(n2438), .A2(n2258), .A3(n2626), .A4(n2441), .ZN(n2639)
         );
  NAND2_X1 U3050 ( .A1(n2639), .A2(IR_REG_31__SCAN_IN), .ZN(n2640) );
  OR2_X1 U3051 ( .A1(n4035), .A2(n2397), .ZN(n2392) );
  NAND2_X1 U3052 ( .A1(n2391), .A2(n2393), .ZN(n3996) );
  NAND2_X1 U3053 ( .A1(n4035), .A2(n2395), .ZN(n2391) );
  AOI21_X1 U3054 ( .B1(n4035), .B2(n3867), .A(n3869), .ZN(n4018) );
  NAND2_X1 U3055 ( .A1(n2256), .A2(n2399), .ZN(n2400) );
  AND2_X1 U3056 ( .A1(n3035), .A2(n2681), .ZN(n2399) );
  INV_X1 U3057 ( .A(n3035), .ZN(n2679) );
  NAND3_X1 U3058 ( .A1(n2401), .A2(n2686), .A3(n2400), .ZN(n3110) );
  NAND3_X1 U3059 ( .A1(n3031), .A2(n2256), .A3(n2681), .ZN(n2401) );
  NAND2_X1 U3060 ( .A1(n3230), .A2(n2406), .ZN(n2404) );
  NAND2_X1 U3061 ( .A1(n2780), .A2(n2420), .ZN(n2419) );
  NAND2_X1 U3062 ( .A1(n2780), .A2(n2779), .ZN(n3479) );
  INV_X1 U3063 ( .A(n2780), .ZN(n2424) );
  AOI21_X1 U3064 ( .B1(n4101), .B2(n2429), .A(n2427), .ZN(n4047) );
  NAND3_X1 U3065 ( .A1(n2489), .A2(n2488), .A3(n2442), .ZN(n2563) );
  NAND2_X1 U3066 ( .A1(n3656), .A2(n3595), .ZN(n3655) );
  NAND2_X1 U3067 ( .A1(n2262), .A2(REG3_REG_1__SCAN_IN), .ZN(n2663) );
  XNOR2_X1 U3068 ( .A(n4077), .B(n4086), .ZN(n4281) );
  NAND2_X1 U3069 ( .A1(n3076), .A2(n3026), .ZN(n2873) );
  OR2_X1 U3070 ( .A1(n2998), .A2(n2967), .ZN(n4418) );
  NAND2_X1 U3071 ( .A1(n2570), .A2(n2569), .ZN(n2572) );
  NAND2_X1 U3072 ( .A1(n2591), .A2(n2625), .ZN(n2569) );
  NOR2_X1 U3073 ( .A1(n4413), .A2(n4414), .ZN(n4412) );
  OR2_X1 U3074 ( .A1(n4007), .A2(n4378), .ZN(n2477) );
  OR2_X1 U3075 ( .A1(n4007), .A2(n4333), .ZN(n2478) );
  OR2_X1 U3076 ( .A1(n4410), .A2(n4416), .ZN(n4531) );
  AND2_X1 U3077 ( .A1(n2634), .A2(n3747), .ZN(n2479) );
  AND3_X1 U3078 ( .A1(n2849), .A2(n2848), .A3(n2847), .ZN(n4258) );
  INV_X1 U3079 ( .A(n4258), .ZN(n4038) );
  AND4_X1 U3080 ( .A1(n2822), .A2(n2821), .A3(n2820), .A4(n2819), .ZN(n4276)
         );
  INV_X1 U3081 ( .A(n4129), .ZN(n3660) );
  OR2_X1 U3082 ( .A1(n4583), .A2(n5043), .ZN(n2480) );
  AND2_X1 U3083 ( .A1(n3139), .A2(n3138), .ZN(n2481) );
  AND2_X1 U3084 ( .A1(n2835), .A2(DATAI_23_), .ZN(n3592) );
  AND2_X1 U3085 ( .A1(n3464), .A2(n2777), .ZN(n2482) );
  NAND2_X1 U3086 ( .A1(n3723), .A2(n3724), .ZN(n3722) );
  NAND2_X1 U3087 ( .A1(n2835), .A2(DATAI_22_), .ZN(n4112) );
  INV_X1 U3088 ( .A(IR_REG_18__SCAN_IN), .ZN(n2562) );
  INV_X1 U3089 ( .A(n3536), .ZN(n3532) );
  NAND2_X1 U3090 ( .A1(n3533), .A2(n3532), .ZN(n3534) );
  INV_X1 U3091 ( .A(IR_REG_21__SCAN_IN), .ZN(n2564) );
  INV_X1 U3092 ( .A(n3193), .ZN(n3194) );
  INV_X1 U3093 ( .A(n4112), .ZN(n2815) );
  INV_X1 U3094 ( .A(IR_REG_22__SCAN_IN), .ZN(n2565) );
  AND2_X1 U3095 ( .A1(n3123), .A2(REG1_REG_0__SCAN_IN), .ZN(n2999) );
  INV_X1 U3096 ( .A(n2899), .ZN(n2850) );
  NOR2_X1 U3097 ( .A1(n2482), .A2(n2778), .ZN(n2779) );
  AND2_X1 U3098 ( .A1(n3372), .A2(n3371), .ZN(n3375) );
  INV_X1 U3099 ( .A(n4012), .ZN(n3994) );
  AND2_X1 U3100 ( .A1(n4185), .A2(n3562), .ZN(n3848) );
  INV_X1 U3101 ( .A(n3997), .ZN(n3998) );
  INV_X1 U3102 ( .A(n3059), .ZN(n3050) );
  AND2_X1 U3103 ( .A1(n3512), .A2(n3511), .ZN(n3536) );
  AND2_X1 U3104 ( .A1(n3357), .A2(n3360), .ZN(n3358) );
  NAND2_X1 U3105 ( .A1(n3305), .A2(n3306), .ZN(n3307) );
  INV_X1 U3106 ( .A(n3482), .ZN(n3700) );
  NAND2_X1 U3107 ( .A1(n2766), .A2(REG3_REG_16__SCAN_IN), .ZN(n2781) );
  NOR2_X1 U3108 ( .A1(n2788), .A2(n4915), .ZN(n2801) );
  OR3_X1 U3109 ( .A1(n2781), .A2(n2646), .A3(n2645), .ZN(n2788) );
  NOR2_X1 U3110 ( .A1(n2772), .A2(n2644), .ZN(n2766) );
  OR2_X1 U3111 ( .A1(n3649), .A2(n2846), .ZN(n2849) );
  AND4_X1 U3112 ( .A1(n2762), .A2(n2761), .A3(n2760), .A4(n2759), .ZN(n4328)
         );
  INV_X1 U3113 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3362) );
  OR2_X1 U3114 ( .A1(n4410), .A2(n4417), .ZN(n4528) );
  NAND2_X1 U3115 ( .A1(n4038), .A2(n2899), .ZN(n2852) );
  INV_X1 U3116 ( .A(n4593), .ZN(n4634) );
  INV_X1 U3117 ( .A(n4327), .ZN(n4637) );
  INV_X1 U3118 ( .A(n4072), .ZN(n4272) );
  AND2_X1 U3119 ( .A1(n2835), .A2(DATAI_20_), .ZN(n4292) );
  NOR2_X1 U3120 ( .A1(n2707), .A2(n2643), .ZN(n2717) );
  INV_X1 U3121 ( .A(n3666), .ZN(n3667) );
  NAND2_X1 U3122 ( .A1(n2694), .A2(REG3_REG_5__SCAN_IN), .ZN(n2707) );
  AOI21_X1 U3123 ( .B1(n3153), .B2(n3152), .A(n2481), .ZN(n3145) );
  OR2_X1 U3124 ( .A1(n3621), .A2(n3019), .ZN(n3927) );
  AND3_X1 U3125 ( .A1(n2857), .A2(n2856), .A3(n2855), .ZN(n2858) );
  AND4_X1 U3126 ( .A1(n2793), .A2(n2792), .A3(n2791), .A4(n2790), .ZN(n4296)
         );
  AND4_X1 U3127 ( .A1(n2776), .A2(n2775), .A3(n2774), .A4(n2773), .ZN(n3769)
         );
  INV_X1 U3128 ( .A(n4556), .ZN(n4538) );
  INV_X1 U3129 ( .A(n4531), .ZN(n4553) );
  OR2_X1 U3130 ( .A1(n3909), .A2(n3834), .ZN(n4019) );
  AND2_X1 U3131 ( .A1(n4402), .A2(n2937), .ZN(n4560) );
  NAND2_X1 U3132 ( .A1(n2835), .A2(DATAI_26_), .ZN(n4042) );
  NAND2_X1 U3133 ( .A1(n2835), .A2(DATAI_24_), .ZN(n4072) );
  INV_X1 U3134 ( .A(n4646), .ZN(n4590) );
  AND3_X1 U3135 ( .A1(n2869), .A2(n3109), .A3(n2922), .ZN(n4617) );
  OAI22_X1 U3136 ( .A1(n2964), .A2(D_REG_0__SCAN_IN), .B1(n2905), .B2(n4381), 
        .ZN(n2929) );
  NAND2_X1 U3137 ( .A1(n2906), .A2(n2905), .ZN(n2964) );
  AND2_X1 U3138 ( .A1(n2529), .A2(n2528), .ZN(n4581) );
  AND2_X1 U3139 ( .A1(n2633), .A2(n2632), .ZN(n4543) );
  OR2_X1 U3140 ( .A1(n3012), .A2(n3011), .ZN(n3775) );
  NAND2_X1 U3141 ( .A1(n2859), .A2(n2858), .ZN(n4023) );
  INV_X1 U3142 ( .A(n4209), .ZN(n4172) );
  INV_X1 U3143 ( .A(n3769), .ZN(n3933) );
  OR2_X1 U3144 ( .A1(n4410), .A2(n3021), .ZN(n4556) );
  INV_X1 U3145 ( .A(n4402), .ZN(n4204) );
  INV_X1 U3146 ( .A(n4402), .ZN(n4566) );
  NAND2_X1 U3147 ( .A1(n4666), .A2(n4314), .ZN(n4333) );
  NAND2_X1 U31480 ( .A1(n4649), .A2(n4314), .ZN(n4378) );
  INV_X1 U31490 ( .A(n4649), .ZN(n4647) );
  INV_X1 U3150 ( .A(n4570), .ZN(n4571) );
  AND2_X1 U3151 ( .A1(n3120), .A2(STATE_REG_SCAN_IN), .ZN(n4572) );
  NOR2_X1 U3152 ( .A1(n2534), .A2(n2533), .ZN(n4384) );
  INV_X2 U3153 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NOR2_X1 U3154 ( .A1(n2494), .A2(n2959), .ZN(n2492) );
  MUX2_X1 U3155 ( .A(n2959), .B(n2492), .S(IR_REG_17__SCAN_IN), .Z(n2493) );
  INV_X1 U3156 ( .A(n2493), .ZN(n2495) );
  AND2_X1 U3157 ( .A1(n2495), .A2(n2563), .ZN(n2786) );
  INV_X1 U3158 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4310) );
  INV_X1 U3159 ( .A(n2786), .ZN(n4574) );
  AOI22_X1 U3160 ( .A1(n2786), .A2(REG1_REG_17__SCAN_IN), .B1(n4310), .B2(
        n4574), .ZN(n4546) );
  NAND2_X1 U3161 ( .A1(n2434), .A2(n2497), .ZN(n2547) );
  INV_X1 U3162 ( .A(n2547), .ZN(n2498) );
  NAND2_X1 U3163 ( .A1(n2498), .A2(n2548), .ZN(n2550) );
  NAND2_X1 U3164 ( .A1(n2550), .A2(IR_REG_31__SCAN_IN), .ZN(n2500) );
  NAND2_X1 U3165 ( .A1(n2500), .A2(n2499), .ZN(n2556) );
  OR2_X1 U3166 ( .A1(n2500), .A2(n2499), .ZN(n2501) );
  NAND2_X1 U3167 ( .A1(n3950), .A2(REG1_REG_15__SCAN_IN), .ZN(n2554) );
  OAI21_X1 U3168 ( .B1(n3950), .B2(REG1_REG_15__SCAN_IN), .A(n2554), .ZN(n3957) );
  OR2_X1 U3169 ( .A1(n2502), .A2(IR_REG_5__SCAN_IN), .ZN(n2523) );
  INV_X1 U3170 ( .A(IR_REG_6__SCAN_IN), .ZN(n2504) );
  INV_X1 U3171 ( .A(IR_REG_8__SCAN_IN), .ZN(n2503) );
  NAND3_X1 U3172 ( .A1(n4844), .A2(n2504), .A3(n2503), .ZN(n2505) );
  NOR2_X1 U3173 ( .A1(n2523), .A2(n2505), .ZN(n2531) );
  NAND2_X1 U3174 ( .A1(n2531), .A2(n4843), .ZN(n2537) );
  NAND2_X1 U3175 ( .A1(n2506), .A2(IR_REG_31__SCAN_IN), .ZN(n2542) );
  XNOR2_X1 U3176 ( .A(n2542), .B(IR_REG_11__SCAN_IN), .ZN(n2748) );
  OAI21_X1 U3177 ( .B1(n2523), .B2(IR_REG_6__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2527) );
  NAND2_X1 U3178 ( .A1(n2527), .A2(n4844), .ZN(n2529) );
  NAND2_X1 U3179 ( .A1(n2529), .A2(IR_REG_31__SCAN_IN), .ZN(n2507) );
  XNOR2_X1 U3180 ( .A(n2507), .B(IR_REG_8__SCAN_IN), .ZN(n2723) );
  INV_X1 U3181 ( .A(n2723), .ZN(n4580) );
  NAND2_X1 U3182 ( .A1(n2502), .A2(IR_REG_31__SCAN_IN), .ZN(n2508) );
  XNOR2_X1 U3183 ( .A(n2508), .B(IR_REG_5__SCAN_IN), .ZN(n2699) );
  INV_X1 U3184 ( .A(REG1_REG_5__SCAN_IN), .ZN(n5043) );
  AOI22_X1 U3185 ( .A1(n2699), .A2(REG1_REG_5__SCAN_IN), .B1(n5043), .B2(n4583), .ZN(n4448) );
  NAND2_X1 U3186 ( .A1(n2510), .A2(IR_REG_31__SCAN_IN), .ZN(n2513) );
  NAND2_X1 U3187 ( .A1(n2513), .A2(n2512), .ZN(n2515) );
  NAND2_X1 U3188 ( .A1(n2515), .A2(IR_REG_31__SCAN_IN), .ZN(n2511) );
  XNOR2_X1 U3189 ( .A(n2511), .B(IR_REG_4__SCAN_IN), .ZN(n4386) );
  OR2_X1 U3190 ( .A1(n2513), .A2(n2512), .ZN(n2514) );
  INV_X1 U3191 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4873) );
  MUX2_X1 U3192 ( .A(n4873), .B(REG1_REG_2__SCAN_IN), .S(n4434), .Z(n4425) );
  INV_X1 U3193 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4652) );
  NAND2_X1 U3194 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2518)
         );
  INV_X1 U3195 ( .A(n3945), .ZN(n2945) );
  MUX2_X1 U3196 ( .A(REG1_REG_1__SCAN_IN), .B(n4652), .S(n3945), .Z(n3941) );
  NAND3_X1 U3197 ( .A1(n3941), .A2(REG1_REG_0__SCAN_IN), .A3(IR_REG_0__SCAN_IN), .ZN(n3940) );
  OAI21_X1 U3198 ( .B1(n4652), .B2(n2945), .A(n3940), .ZN(n4426) );
  NAND2_X1 U3199 ( .A1(n4425), .A2(n4426), .ZN(n4424) );
  OAI21_X1 U3200 ( .B1(n4873), .B2(n4434), .A(n4424), .ZN(n2519) );
  NAND2_X1 U3201 ( .A1(n4389), .A2(n2519), .ZN(n2520) );
  NAND2_X1 U3202 ( .A1(n4386), .A2(n2521), .ZN(n2522) );
  INV_X1 U3203 ( .A(n4386), .ZN(n4441) );
  NAND2_X1 U3204 ( .A1(n2523), .A2(IR_REG_31__SCAN_IN), .ZN(n2524) );
  XNOR2_X1 U3205 ( .A(n2524), .B(IR_REG_6__SCAN_IN), .ZN(n4457) );
  NAND2_X1 U3206 ( .A1(n2525), .A2(n4457), .ZN(n2526) );
  OR2_X1 U3207 ( .A1(n2527), .A2(n4844), .ZN(n2528) );
  INV_X1 U3208 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4479) );
  NOR2_X1 U3209 ( .A1(n2531), .A2(n2959), .ZN(n2532) );
  MUX2_X1 U32100 ( .A(n2959), .B(n2532), .S(IR_REG_9__SCAN_IN), .Z(n2534) );
  INV_X1 U32110 ( .A(n2537), .ZN(n2533) );
  NAND2_X1 U32120 ( .A1(n4384), .A2(REG1_REG_9__SCAN_IN), .ZN(n2536) );
  OR2_X1 U32130 ( .A1(n4384), .A2(REG1_REG_9__SCAN_IN), .ZN(n2535) );
  NAND2_X1 U32140 ( .A1(n2536), .A2(n2535), .ZN(n3087) );
  NAND2_X1 U32150 ( .A1(n2537), .A2(IR_REG_31__SCAN_IN), .ZN(n2538) );
  XNOR2_X1 U32160 ( .A(n2538), .B(IR_REG_10__SCAN_IN), .ZN(n2740) );
  INV_X1 U32170 ( .A(n2740), .ZN(n4579) );
  NOR2_X1 U32180 ( .A1(n2539), .A2(n4579), .ZN(n2540) );
  INV_X1 U32190 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4488) );
  NOR2_X1 U32200 ( .A1(n2540), .A2(n4486), .ZN(n4497) );
  INV_X1 U32210 ( .A(n2748), .ZN(n4577) );
  INV_X1 U32220 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4664) );
  AOI22_X1 U32230 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4577), .B1(n2748), .B2(
        n4664), .ZN(n4496) );
  INV_X1 U32240 ( .A(IR_REG_11__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U32250 ( .A1(n2542), .A2(n2541), .ZN(n2543) );
  NAND2_X1 U32260 ( .A1(n2543), .A2(IR_REG_31__SCAN_IN), .ZN(n2544) );
  XNOR2_X1 U32270 ( .A(n2544), .B(IR_REG_12__SCAN_IN), .ZN(n2755) );
  INV_X1 U32280 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4507) );
  NAND2_X1 U32290 ( .A1(n2496), .A2(IR_REG_31__SCAN_IN), .ZN(n2546) );
  XNOR2_X1 U32300 ( .A(n2546), .B(IR_REG_13__SCAN_IN), .ZN(n4524) );
  INV_X1 U32310 ( .A(n4524), .ZN(n4575) );
  INV_X1 U32320 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3437) );
  AOI22_X1 U32330 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4575), .B1(n4524), .B2(
        n3437), .ZN(n4520) );
  NAND2_X1 U32340 ( .A1(n2547), .A2(IR_REG_31__SCAN_IN), .ZN(n2549) );
  MUX2_X1 U32350 ( .A(n2549), .B(IR_REG_31__SCAN_IN), .S(n2548), .Z(n2551) );
  NAND2_X1 U32360 ( .A1(n2551), .A2(n2550), .ZN(n2613) );
  INV_X1 U32370 ( .A(n2552), .ZN(n2553) );
  INV_X1 U32380 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4533) );
  INV_X1 U32390 ( .A(n2554), .ZN(n2555) );
  NAND2_X1 U32400 ( .A1(n2556), .A2(IR_REG_31__SCAN_IN), .ZN(n2557) );
  XNOR2_X1 U32410 ( .A(n2557), .B(IR_REG_16__SCAN_IN), .ZN(n4383) );
  INV_X1 U32420 ( .A(n4383), .ZN(n2617) );
  NAND2_X1 U32430 ( .A1(n2558), .A2(n2617), .ZN(n2559) );
  INV_X1 U32440 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4951) );
  NAND2_X1 U32450 ( .A1(n2563), .A2(IR_REG_31__SCAN_IN), .ZN(n2560) );
  XNOR2_X1 U32460 ( .A(n2560), .B(IR_REG_18__SCAN_IN), .ZN(n4382) );
  NAND2_X1 U32470 ( .A1(n4382), .A2(REG1_REG_18__SCAN_IN), .ZN(n3974) );
  OR2_X1 U32480 ( .A1(n4382), .A2(REG1_REG_18__SCAN_IN), .ZN(n2561) );
  NAND2_X1 U32490 ( .A1(n2625), .A2(IR_REG_27__SCAN_IN), .ZN(n2571) );
  NOR2_X1 U32500 ( .A1(n2573), .A2(n2959), .ZN(n2574) );
  MUX2_X1 U32510 ( .A(n2959), .B(n2574), .S(IR_REG_23__SCAN_IN), .Z(n2575) );
  INV_X1 U32520 ( .A(n2575), .ZN(n2576) );
  NAND2_X1 U32530 ( .A1(n2576), .A2(n2584), .ZN(n3120) );
  NAND2_X1 U32540 ( .A1(n2267), .A2(IR_REG_31__SCAN_IN), .ZN(n2577) );
  MUX2_X1 U32550 ( .A(IR_REG_31__SCAN_IN), .B(n2577), .S(IR_REG_22__SCAN_IN), 
        .Z(n2579) );
  INV_X1 U32560 ( .A(n2573), .ZN(n2578) );
  NAND2_X1 U32570 ( .A1(n2271), .A2(IR_REG_31__SCAN_IN), .ZN(n2580) );
  NAND2_X1 U32580 ( .A1(n3928), .A2(n3920), .ZN(n3008) );
  INV_X1 U32590 ( .A(n3008), .ZN(n2868) );
  NAND2_X1 U32600 ( .A1(n3120), .A2(n2868), .ZN(n2581) );
  AND2_X1 U32610 ( .A1(n2835), .A2(n2581), .ZN(n2631) );
  INV_X1 U32620 ( .A(n2627), .ZN(n2586) );
  NAND2_X1 U32630 ( .A1(n2586), .A2(IR_REG_31__SCAN_IN), .ZN(n2582) );
  MUX2_X1 U32640 ( .A(n2582), .B(IR_REG_31__SCAN_IN), .S(n2567), .Z(n2583) );
  NAND2_X1 U32650 ( .A1(n2583), .A2(n2588), .ZN(n2917) );
  MUX2_X1 U32660 ( .A(IR_REG_31__SCAN_IN), .B(n2585), .S(IR_REG_24__SCAN_IN), 
        .Z(n2587) );
  NAND2_X1 U32670 ( .A1(n2587), .A2(n2586), .ZN(n2920) );
  NAND2_X1 U32680 ( .A1(n2588), .A2(IR_REG_31__SCAN_IN), .ZN(n2589) );
  NAND2_X1 U32690 ( .A1(n2998), .A2(n4572), .ZN(n3016) );
  OR2_X1 U32700 ( .A1(n3120), .A2(U3149), .ZN(n3931) );
  NAND2_X1 U32710 ( .A1(n3016), .A2(n3931), .ZN(n2632) );
  NAND2_X1 U32720 ( .A1(n2631), .A2(n2632), .ZN(n4410) );
  XNOR2_X1 U32730 ( .A(n2591), .B(n2568), .ZN(n4406) );
  INV_X1 U32740 ( .A(n4406), .ZN(n4416) );
  NOR2_X1 U32750 ( .A1(n2786), .A2(REG2_REG_17__SCAN_IN), .ZN(n2592) );
  AOI21_X1 U32760 ( .B1(REG2_REG_17__SCAN_IN), .B2(n2786), .A(n2592), .ZN(
        n4549) );
  NAND2_X1 U32770 ( .A1(n3950), .A2(REG2_REG_15__SCAN_IN), .ZN(n2615) );
  OAI21_X1 U32780 ( .B1(n3950), .B2(REG2_REG_15__SCAN_IN), .A(n2615), .ZN(
        n3952) );
  INV_X1 U32790 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2609) );
  AOI22_X1 U32800 ( .A1(REG2_REG_11__SCAN_IN), .A2(n2748), .B1(n4577), .B2(
        n2609), .ZN(n4502) );
  NAND2_X1 U32810 ( .A1(n4384), .A2(REG2_REG_9__SCAN_IN), .ZN(n2606) );
  INV_X1 U32820 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2593) );
  MUX2_X1 U32830 ( .A(REG2_REG_9__SCAN_IN), .B(n2593), .S(n4384), .Z(n3083) );
  NAND2_X1 U32840 ( .A1(REG2_REG_7__SCAN_IN), .A2(n4581), .ZN(n2603) );
  INV_X1 U32850 ( .A(n4581), .ZN(n4476) );
  INV_X1 U32860 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3186) );
  AOI22_X1 U32870 ( .A1(REG2_REG_7__SCAN_IN), .A2(n4581), .B1(n4476), .B2(
        n3186), .ZN(n4473) );
  INV_X1 U32880 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2600) );
  AOI22_X1 U32890 ( .A1(n2699), .A2(REG2_REG_5__SCAN_IN), .B1(n2600), .B2(
        n4583), .ZN(n4451) );
  INV_X1 U32900 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2595) );
  MUX2_X1 U32910 ( .A(n2595), .B(REG2_REG_2__SCAN_IN), .S(n4434), .Z(n4430) );
  INV_X1 U32920 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2594) );
  MUX2_X1 U32930 ( .A(REG2_REG_1__SCAN_IN), .B(n2594), .S(n3945), .Z(n3944) );
  NAND3_X1 U32940 ( .A1(n3944), .A2(REG2_REG_0__SCAN_IN), .A3(
        IR_REG_0__SCAN_IN), .ZN(n3943) );
  OAI21_X1 U32950 ( .B1(n2594), .B2(n2945), .A(n3943), .ZN(n4431) );
  NAND2_X1 U32960 ( .A1(n4430), .A2(n4431), .ZN(n4429) );
  OAI21_X1 U32970 ( .B1(n2595), .B2(n4434), .A(n4429), .ZN(n2596) );
  NAND2_X1 U32980 ( .A1(n4389), .A2(n2596), .ZN(n2597) );
  NAND2_X1 U32990 ( .A1(n4386), .A2(n2598), .ZN(n2599) );
  NAND2_X1 U33000 ( .A1(REG2_REG_4__SCAN_IN), .A2(n4436), .ZN(n4435) );
  NAND2_X1 U33010 ( .A1(n2601), .A2(n4457), .ZN(n2602) );
  NAND2_X1 U33020 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4461), .ZN(n4460) );
  NAND2_X1 U33030 ( .A1(n2602), .A2(n4460), .ZN(n4472) );
  NAND2_X1 U33040 ( .A1(n4473), .A2(n4472), .ZN(n4471) );
  NAND2_X1 U33050 ( .A1(n2603), .A2(n4471), .ZN(n2604) );
  NAND2_X1 U33060 ( .A1(n2723), .A2(n2604), .ZN(n2605) );
  XNOR2_X1 U33070 ( .A(n2604), .B(n4580), .ZN(n4483) );
  NAND2_X1 U33080 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4483), .ZN(n4482) );
  NAND2_X1 U33090 ( .A1(n2605), .A2(n4482), .ZN(n3084) );
  NAND2_X1 U33100 ( .A1(n3083), .A2(n3084), .ZN(n3082) );
  NAND2_X1 U33110 ( .A1(n2606), .A2(n3082), .ZN(n2607) );
  NAND2_X1 U33120 ( .A1(n2740), .A2(n2607), .ZN(n2608) );
  XNOR2_X1 U33130 ( .A(n2607), .B(n4579), .ZN(n4492) );
  NAND2_X1 U33140 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4492), .ZN(n4491) );
  NAND2_X1 U33150 ( .A1(n2608), .A2(n4491), .ZN(n4501) );
  NAND2_X1 U33160 ( .A1(n4502), .A2(n4501), .ZN(n4500) );
  NAND2_X1 U33170 ( .A1(n2755), .A2(n2610), .ZN(n2611) );
  INV_X1 U33180 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4978) );
  NOR2_X1 U33190 ( .A1(n4978), .A2(n4575), .ZN(n4515) );
  INV_X1 U33200 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4529) );
  INV_X1 U33210 ( .A(n2615), .ZN(n2616) );
  NAND2_X1 U33220 ( .A1(n2618), .A2(n2617), .ZN(n2619) );
  INV_X1 U33230 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3967) );
  NAND2_X1 U33240 ( .A1(n3968), .A2(n3967), .ZN(n3966) );
  NAND2_X1 U33250 ( .A1(n2619), .A2(n3966), .ZN(n4548) );
  XNOR2_X1 U33260 ( .A(n4382), .B(REG2_REG_18__SCAN_IN), .ZN(n2629) );
  NAND2_X1 U33270 ( .A1(n2568), .A2(n4842), .ZN(n2620) );
  NOR2_X1 U33280 ( .A1(IR_REG_25__SCAN_IN), .A2(n2620), .ZN(n2624) );
  AND2_X1 U33290 ( .A1(n2627), .A2(n2624), .ZN(n2621) );
  NOR2_X1 U33300 ( .A1(n2621), .A2(n2959), .ZN(n2622) );
  MUX2_X1 U33310 ( .A(n2959), .B(n2622), .S(IR_REG_28__SCAN_IN), .Z(n2623) );
  INV_X1 U33320 ( .A(n2623), .ZN(n2628) );
  AND2_X1 U33330 ( .A1(n2625), .A2(n2624), .ZN(n2626) );
  NAND2_X1 U33340 ( .A1(n2628), .A2(n2639), .ZN(n4415) );
  NAND2_X1 U33350 ( .A1(n3021), .A2(n4416), .ZN(n4417) );
  AOI211_X1 U33360 ( .C1(n2630), .C2(n2629), .A(n4528), .B(n2248), .ZN(n2637)
         );
  NAND2_X1 U33370 ( .A1(n4538), .A2(n4382), .ZN(n2635) );
  INV_X1 U33380 ( .A(n2631), .ZN(n2633) );
  INV_X1 U33390 ( .A(n4543), .ZN(n4527) );
  INV_X1 U33400 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n4898) );
  OR2_X1 U33410 ( .A1(n4527), .A2(n4898), .ZN(n2634) );
  NAND2_X1 U33420 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n3747) );
  NAND2_X1 U33430 ( .A1(n2635), .A2(n2479), .ZN(n2636) );
  INV_X1 U33440 ( .A(n2641), .ZN(n2960) );
  INV_X1 U33450 ( .A(n2262), .ZN(n2846) );
  NAND2_X1 U33460 ( .A1(REG3_REG_7__SCAN_IN), .A2(REG3_REG_6__SCAN_IN), .ZN(
        n2643) );
  NAND2_X1 U33470 ( .A1(n2717), .A2(REG3_REG_8__SCAN_IN), .ZN(n2727) );
  NAND2_X1 U33480 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n2644) );
  INV_X1 U33490 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2646) );
  INV_X1 U33500 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2645) );
  OAI21_X1 U33510 ( .B1(n2781), .B2(n2646), .A(n2645), .ZN(n2647) );
  AND2_X1 U33520 ( .A1(n2647), .A2(n2788), .ZN(n4197) );
  NAND2_X1 U3353 ( .A1(n2865), .A2(n4197), .ZN(n2654) );
  INV_X1 U33540 ( .A(n2648), .ZN(n2649) );
  NAND2_X1 U3355 ( .A1(n2671), .A2(REG0_REG_18__SCAN_IN), .ZN(n2653) );
  NAND2_X1 U3356 ( .A1(n2240), .A2(REG1_REG_18__SCAN_IN), .ZN(n2652) );
  NAND2_X1 U3357 ( .A1(n2239), .A2(REG2_REG_18__SCAN_IN), .ZN(n2651) );
  MUX2_X1 U3358 ( .A(n4382), .B(DATAI_18_), .S(n2835), .Z(n4184) );
  MUX2_X1 U3359 ( .A(n4383), .B(DATAI_16_), .S(n2835), .Z(n3482) );
  OR2_X1 U3360 ( .A1(n2766), .A2(REG3_REG_16__SCAN_IN), .ZN(n2655) );
  AND2_X1 U3361 ( .A1(n2781), .A2(n2655), .ZN(n3702) );
  NAND2_X1 U3362 ( .A1(n2865), .A2(n3702), .ZN(n2659) );
  NAND2_X1 U3363 ( .A1(n2244), .A2(REG2_REG_16__SCAN_IN), .ZN(n2658) );
  NAND2_X1 U3364 ( .A1(n2671), .A2(REG0_REG_16__SCAN_IN), .ZN(n2657) );
  NAND2_X1 U3365 ( .A1(n2240), .A2(REG1_REG_16__SCAN_IN), .ZN(n2656) );
  NAND2_X1 U3366 ( .A1(n2239), .A2(REG2_REG_1__SCAN_IN), .ZN(n2662) );
  NAND2_X1 U3367 ( .A1(n2671), .A2(REG0_REG_1__SCAN_IN), .ZN(n2661) );
  NAND2_X1 U3368 ( .A1(n2240), .A2(REG1_REG_1__SCAN_IN), .ZN(n2660) );
  NAND2_X1 U3369 ( .A1(n2262), .A2(REG3_REG_0__SCAN_IN), .ZN(n2668) );
  NAND2_X1 U3370 ( .A1(n2242), .A2(REG1_REG_0__SCAN_IN), .ZN(n2667) );
  NAND2_X1 U3371 ( .A1(n2671), .A2(REG0_REG_0__SCAN_IN), .ZN(n2666) );
  NAND2_X1 U3372 ( .A1(n2244), .A2(REG2_REG_0__SCAN_IN), .ZN(n2665) );
  AND2_X1 U3373 ( .A1(n2971), .A2(n4670), .ZN(n2935) );
  NAND2_X1 U3374 ( .A1(n2871), .A2(n2935), .ZN(n2934) );
  NAND2_X1 U3375 ( .A1(n2669), .A2(n3026), .ZN(n2670) );
  NAND2_X1 U3376 ( .A1(n2934), .A2(n2670), .ZN(n3031) );
  NAND2_X1 U3377 ( .A1(n2262), .A2(REG3_REG_2__SCAN_IN), .ZN(n2676) );
  NAND2_X1 U3378 ( .A1(n2671), .A2(REG0_REG_2__SCAN_IN), .ZN(n2675) );
  NAND2_X1 U3379 ( .A1(n2241), .A2(REG1_REG_2__SCAN_IN), .ZN(n2674) );
  NAND2_X1 U3380 ( .A1(n2239), .A2(REG2_REG_2__SCAN_IN), .ZN(n2673) );
  AND4_X2 U3381 ( .A1(n2676), .A2(n2675), .A3(n2674), .A4(n2673), .ZN(n2680)
         );
  INV_X1 U3382 ( .A(n2680), .ZN(n3939) );
  INV_X1 U3383 ( .A(n4434), .ZN(n2678) );
  MUX2_X1 U3384 ( .A(n2678), .B(DATAI_2_), .S(n2677), .Z(n3059) );
  NAND2_X1 U3385 ( .A1(n3939), .A2(n3050), .ZN(n3785) );
  NAND2_X1 U3386 ( .A1(n2680), .A2(n3059), .ZN(n3782) );
  AND2_X2 U3387 ( .A1(n3785), .A2(n3782), .ZN(n3035) );
  NAND2_X1 U3388 ( .A1(n2680), .A2(n3050), .ZN(n2681) );
  NAND2_X1 U3389 ( .A1(n2240), .A2(REG1_REG_3__SCAN_IN), .ZN(n2684) );
  NAND2_X1 U3390 ( .A1(n2239), .A2(REG2_REG_3__SCAN_IN), .ZN(n2683) );
  NAND2_X1 U3391 ( .A1(n2671), .A2(REG0_REG_3__SCAN_IN), .ZN(n2682) );
  NAND4_X1 U3392 ( .A1(n2685), .A2(n2684), .A3(n2683), .A4(n2682), .ZN(n3938)
         );
  MUX2_X1 U3393 ( .A(n4389), .B(DATAI_3_), .S(n2835), .Z(n3132) );
  NAND2_X1 U3394 ( .A1(n3938), .A2(n3132), .ZN(n2686) );
  NOR2_X1 U3395 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2687) );
  NOR2_X1 U3396 ( .A1(n2694), .A2(n2687), .ZN(n3126) );
  NAND2_X1 U3397 ( .A1(n2262), .A2(n3126), .ZN(n2691) );
  NAND2_X1 U3398 ( .A1(n2671), .A2(REG0_REG_4__SCAN_IN), .ZN(n2690) );
  NAND2_X1 U3399 ( .A1(n2241), .A2(REG1_REG_4__SCAN_IN), .ZN(n2689) );
  NAND2_X1 U3400 ( .A1(n2244), .A2(REG2_REG_4__SCAN_IN), .ZN(n2688) );
  MUX2_X1 U3401 ( .A(n4386), .B(DATAI_4_), .S(n2835), .Z(n3140) );
  NAND2_X1 U3402 ( .A1(n3171), .A2(n3140), .ZN(n3788) );
  INV_X1 U3403 ( .A(n3140), .ZN(n3147) );
  NAND2_X1 U3404 ( .A1(n3937), .A2(n3147), .ZN(n3791) );
  NAND2_X1 U3405 ( .A1(n3788), .A2(n3791), .ZN(n3874) );
  NAND2_X1 U3406 ( .A1(n3110), .A2(n3874), .ZN(n2693) );
  NAND2_X1 U3407 ( .A1(n3937), .A2(n3140), .ZN(n2692) );
  NAND2_X1 U3408 ( .A1(n2693), .A2(n2692), .ZN(n3099) );
  OAI21_X1 U3409 ( .B1(n2694), .B2(REG3_REG_5__SCAN_IN), .A(n2707), .ZN(n3176)
         );
  INV_X1 U3410 ( .A(n3176), .ZN(n3102) );
  NAND2_X1 U3411 ( .A1(n2262), .A2(n3102), .ZN(n2698) );
  NAND2_X1 U3412 ( .A1(n2239), .A2(REG2_REG_5__SCAN_IN), .ZN(n2697) );
  NAND2_X1 U3413 ( .A1(n2671), .A2(REG0_REG_5__SCAN_IN), .ZN(n2696) );
  NAND2_X1 U3414 ( .A1(n2242), .A2(REG1_REG_5__SCAN_IN), .ZN(n2695) );
  NAND4_X1 U3415 ( .A1(n2698), .A2(n2697), .A3(n2696), .A4(n2695), .ZN(n3936)
         );
  MUX2_X1 U3416 ( .A(n2699), .B(DATAI_5_), .S(n2835), .Z(n3167) );
  AND2_X1 U3417 ( .A1(n3936), .A2(n3167), .ZN(n2700) );
  INV_X1 U3418 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3205) );
  XOR2_X1 U3419 ( .A(n2707), .B(n3205), .Z(n4558) );
  NAND2_X1 U3420 ( .A1(n2865), .A2(n4558), .ZN(n2704) );
  NAND2_X1 U3421 ( .A1(n2240), .A2(REG1_REG_6__SCAN_IN), .ZN(n2703) );
  NAND2_X1 U3422 ( .A1(n2244), .A2(REG2_REG_6__SCAN_IN), .ZN(n2702) );
  NAND2_X1 U3423 ( .A1(n2671), .A2(REG0_REG_6__SCAN_IN), .ZN(n2701) );
  NAND4_X1 U3424 ( .A1(n2704), .A2(n2703), .A3(n2702), .A4(n2701), .ZN(n3935)
         );
  NOR2_X1 U3425 ( .A1(n3935), .A2(n3264), .ZN(n2706) );
  NAND2_X1 U3426 ( .A1(n3935), .A2(n3264), .ZN(n2705) );
  INV_X1 U3427 ( .A(n2707), .ZN(n2708) );
  AOI21_X1 U3428 ( .B1(n2708), .B2(REG3_REG_6__SCAN_IN), .A(
        REG3_REG_7__SCAN_IN), .ZN(n2709) );
  OR2_X1 U3429 ( .A1(n2709), .A2(n2717), .ZN(n3252) );
  INV_X1 U3430 ( .A(n3252), .ZN(n2710) );
  NAND2_X1 U3431 ( .A1(n2262), .A2(n2710), .ZN(n2714) );
  NAND2_X1 U3432 ( .A1(n2671), .A2(REG0_REG_7__SCAN_IN), .ZN(n2713) );
  NAND2_X1 U3433 ( .A1(n2241), .A2(REG1_REG_7__SCAN_IN), .ZN(n2712) );
  NAND2_X1 U3434 ( .A1(n2244), .A2(REG2_REG_7__SCAN_IN), .ZN(n2711) );
  MUX2_X1 U3435 ( .A(n4581), .B(DATAI_7_), .S(n2835), .Z(n3237) );
  NAND2_X1 U3436 ( .A1(n3525), .A2(n3237), .ZN(n2877) );
  NAND2_X1 U3437 ( .A1(n3255), .A2(n3247), .ZN(n3796) );
  NAND2_X1 U3438 ( .A1(n2877), .A2(n3796), .ZN(n3178) );
  NAND2_X1 U3439 ( .A1(n3177), .A2(n3178), .ZN(n2716) );
  NAND2_X1 U3440 ( .A1(n3255), .A2(n3237), .ZN(n2715) );
  NAND2_X1 U3441 ( .A1(n2716), .A2(n2715), .ZN(n3211) );
  OR2_X1 U3442 ( .A1(n2717), .A2(REG3_REG_8__SCAN_IN), .ZN(n2718) );
  AND2_X1 U3443 ( .A1(n2727), .A2(n2718), .ZN(n3528) );
  NAND2_X1 U3444 ( .A1(n2865), .A2(n3528), .ZN(n2722) );
  NAND2_X1 U3445 ( .A1(n2244), .A2(REG2_REG_8__SCAN_IN), .ZN(n2721) );
  NAND2_X1 U3446 ( .A1(n2671), .A2(REG0_REG_8__SCAN_IN), .ZN(n2720) );
  NAND2_X1 U3447 ( .A1(n2242), .A2(REG1_REG_8__SCAN_IN), .ZN(n2719) );
  NAND4_X1 U3448 ( .A1(n2722), .A2(n2721), .A3(n2720), .A4(n2719), .ZN(n3249)
         );
  MUX2_X1 U3449 ( .A(n2723), .B(DATAI_8_), .S(n2835), .Z(n3283) );
  AND2_X1 U3450 ( .A1(n3249), .A2(n3283), .ZN(n2725) );
  NAND2_X1 U3451 ( .A1(n3313), .A2(n3526), .ZN(n2724) );
  NAND2_X1 U3452 ( .A1(n2727), .A2(n2726), .ZN(n2728) );
  AND2_X1 U3453 ( .A1(n2734), .A2(n2728), .ZN(n3317) );
  NAND2_X1 U3454 ( .A1(n2865), .A2(n3317), .ZN(n2732) );
  NAND2_X1 U3455 ( .A1(n2671), .A2(REG0_REG_9__SCAN_IN), .ZN(n2731) );
  NAND2_X1 U3456 ( .A1(n2240), .A2(REG1_REG_9__SCAN_IN), .ZN(n2730) );
  NAND2_X1 U3457 ( .A1(n2244), .A2(REG2_REG_9__SCAN_IN), .ZN(n2729) );
  NAND4_X1 U34580 ( .A1(n2732), .A2(n2731), .A3(n2730), .A4(n2729), .ZN(n3934)
         );
  MUX2_X1 U34590 ( .A(n4384), .B(DATAI_9_), .S(n2835), .Z(n3227) );
  NOR2_X1 U3460 ( .A1(n3934), .A2(n3227), .ZN(n2733) );
  AND2_X1 U3461 ( .A1(n2734), .A2(n3362), .ZN(n2735) );
  NOR2_X1 U3462 ( .A1(n2742), .A2(n2735), .ZN(n3275) );
  NAND2_X1 U3463 ( .A1(n2865), .A2(n3275), .ZN(n2739) );
  NAND2_X1 U3464 ( .A1(n2239), .A2(REG2_REG_10__SCAN_IN), .ZN(n2738) );
  NAND2_X1 U3465 ( .A1(n2671), .A2(REG0_REG_10__SCAN_IN), .ZN(n2737) );
  NAND2_X1 U3466 ( .A1(n2242), .A2(REG1_REG_10__SCAN_IN), .ZN(n2736) );
  NAND4_X1 U34670 ( .A1(n2739), .A2(n2738), .A3(n2737), .A4(n2736), .ZN(n4638)
         );
  AND2_X1 U3468 ( .A1(n4638), .A2(n3356), .ZN(n2741) );
  INV_X1 U34690 ( .A(n4638), .ZN(n3383) );
  INV_X1 U3470 ( .A(n3356), .ZN(n3364) );
  NOR2_X1 U34710 ( .A1(n2742), .A2(REG3_REG_11__SCAN_IN), .ZN(n2743) );
  OR2_X1 U3472 ( .A1(n2749), .A2(n2743), .ZN(n3297) );
  INV_X1 U34730 ( .A(n3297), .ZN(n3386) );
  NAND2_X1 U3474 ( .A1(n2865), .A2(n3386), .ZN(n2747) );
  NAND2_X1 U34750 ( .A1(n2239), .A2(REG2_REG_11__SCAN_IN), .ZN(n2746) );
  NAND2_X1 U3476 ( .A1(n2671), .A2(REG0_REG_11__SCAN_IN), .ZN(n2745) );
  NAND2_X1 U34770 ( .A1(n2241), .A2(REG1_REG_11__SCAN_IN), .ZN(n2744) );
  MUX2_X1 U3478 ( .A(n2748), .B(DATAI_11_), .S(n2835), .Z(n4633) );
  NAND2_X1 U34790 ( .A1(n3393), .A2(n4633), .ZN(n3343) );
  NAND2_X1 U3480 ( .A1(n3428), .A2(n3384), .ZN(n3814) );
  NAND2_X1 U34810 ( .A1(n3343), .A2(n3814), .ZN(n3855) );
  OR2_X1 U3482 ( .A1(n2749), .A2(REG3_REG_12__SCAN_IN), .ZN(n2750) );
  AND2_X1 U34830 ( .A1(n2757), .A2(n2750), .ZN(n3432) );
  NAND2_X1 U3484 ( .A1(n2865), .A2(n3432), .ZN(n2754) );
  NAND2_X1 U34850 ( .A1(n2671), .A2(REG0_REG_12__SCAN_IN), .ZN(n2753) );
  NAND2_X1 U3486 ( .A1(n2242), .A2(REG1_REG_12__SCAN_IN), .ZN(n2752) );
  NAND2_X1 U34870 ( .A1(n2244), .A2(REG2_REG_12__SCAN_IN), .ZN(n2751) );
  NAND4_X1 U3488 ( .A1(n2754), .A2(n2753), .A3(n2752), .A4(n2751), .ZN(n4636)
         );
  MUX2_X1 U34890 ( .A(n2755), .B(DATAI_12_), .S(n2835), .Z(n3429) );
  NOR2_X1 U3490 ( .A1(n4636), .A2(n3429), .ZN(n2756) );
  NAND2_X1 U34910 ( .A1(n2757), .A2(n4836), .ZN(n2758) );
  AND2_X1 U3492 ( .A1(n2772), .A2(n2758), .ZN(n3460) );
  NAND2_X1 U34930 ( .A1(n2865), .A2(n3460), .ZN(n2762) );
  NAND2_X1 U3494 ( .A1(n2244), .A2(REG2_REG_13__SCAN_IN), .ZN(n2761) );
  NAND2_X1 U34950 ( .A1(n2671), .A2(REG0_REG_13__SCAN_IN), .ZN(n2760) );
  NAND2_X1 U3496 ( .A1(n2241), .A2(REG1_REG_13__SCAN_IN), .ZN(n2759) );
  INV_X1 U34970 ( .A(DATAI_13_), .ZN(n2763) );
  MUX2_X1 U3498 ( .A(n4575), .B(n2763), .S(n2835), .Z(n3447) );
  NAND2_X1 U34990 ( .A1(n4328), .A2(n3447), .ZN(n2764) );
  INV_X1 U3500 ( .A(n2772), .ZN(n2765) );
  AOI21_X1 U35010 ( .B1(n2765), .B2(REG3_REG_14__SCAN_IN), .A(
        REG3_REG_15__SCAN_IN), .ZN(n2767) );
  NOR2_X1 U3502 ( .A1(n2767), .A2(n2766), .ZN(n3772) );
  NAND2_X1 U35030 ( .A1(n2865), .A2(n3772), .ZN(n2771) );
  NAND2_X1 U3504 ( .A1(n2239), .A2(REG2_REG_15__SCAN_IN), .ZN(n2770) );
  NAND2_X1 U35050 ( .A1(n2671), .A2(REG0_REG_15__SCAN_IN), .ZN(n2769) );
  NAND2_X1 U35060 ( .A1(n2240), .A2(REG1_REG_15__SCAN_IN), .ZN(n2768) );
  NAND4_X1 U35070 ( .A1(n2771), .A2(n2770), .A3(n2769), .A4(n2768), .ZN(n4325)
         );
  MUX2_X1 U35080 ( .A(n3950), .B(DATAI_15_), .S(n2835), .Z(n3541) );
  NAND2_X1 U35090 ( .A1(n4325), .A2(n3541), .ZN(n2777) );
  XNOR2_X1 U35100 ( .A(n2772), .B(REG3_REG_14__SCAN_IN), .ZN(n3517) );
  NAND2_X1 U35110 ( .A1(n2865), .A2(n3517), .ZN(n2776) );
  NAND2_X1 U35120 ( .A1(n2671), .A2(REG0_REG_14__SCAN_IN), .ZN(n2775) );
  NAND2_X1 U35130 ( .A1(n2241), .A2(REG1_REG_14__SCAN_IN), .ZN(n2774) );
  NAND2_X1 U35140 ( .A1(n2239), .A2(REG2_REG_14__SCAN_IN), .ZN(n2773) );
  MUX2_X1 U35150 ( .A(n4537), .B(DATAI_14_), .S(n2835), .Z(n4324) );
  NAND2_X1 U35160 ( .A1(n3769), .A2(n4324), .ZN(n3820) );
  NAND2_X1 U35170 ( .A1(n3933), .A2(n3509), .ZN(n3800) );
  NAND2_X1 U35180 ( .A1(n3820), .A2(n3800), .ZN(n3878) );
  NAND3_X1 U35190 ( .A1(n3463), .A2(n2777), .A3(n3878), .ZN(n2780) );
  NOR2_X1 U35200 ( .A1(n3933), .A2(n4324), .ZN(n3464) );
  NAND2_X1 U35210 ( .A1(n3710), .A2(n3482), .ZN(n3892) );
  NAND2_X1 U35220 ( .A1(n4211), .A2(n3700), .ZN(n3894) );
  XNOR2_X1 U35230 ( .A(n2781), .B(REG3_REG_17__SCAN_IN), .ZN(n4218) );
  NAND2_X1 U35240 ( .A1(n2865), .A2(n4218), .ZN(n2785) );
  NAND2_X1 U35250 ( .A1(n2671), .A2(REG0_REG_17__SCAN_IN), .ZN(n2784) );
  NAND2_X1 U35260 ( .A1(n2242), .A2(REG1_REG_17__SCAN_IN), .ZN(n2783) );
  NAND2_X1 U35270 ( .A1(n2244), .A2(REG2_REG_17__SCAN_IN), .ZN(n2782) );
  NAND4_X1 U35280 ( .A1(n2785), .A2(n2784), .A3(n2783), .A4(n2782), .ZN(n3745)
         );
  MUX2_X1 U35290 ( .A(n2786), .B(DATAI_17_), .S(n2835), .Z(n4215) );
  NOR2_X1 U35300 ( .A1(n3745), .A2(n4215), .ZN(n2787) );
  INV_X1 U35310 ( .A(n3745), .ZN(n4187) );
  INV_X1 U35320 ( .A(n4215), .ZN(n4208) );
  NAND2_X1 U35330 ( .A1(n4209), .A2(n4184), .ZN(n4167) );
  NAND2_X1 U35340 ( .A1(n4172), .A2(n4194), .ZN(n4165) );
  NAND2_X1 U35350 ( .A1(n4167), .A2(n4165), .ZN(n4182) );
  INV_X1 U35360 ( .A(n4182), .ZN(n4193) );
  NOR2_X1 U35370 ( .A1(n4192), .A2(n4193), .ZN(n4191) );
  INV_X1 U35380 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4915) );
  AND2_X1 U35390 ( .A1(n2788), .A2(n4915), .ZN(n2789) );
  NOR2_X1 U35400 ( .A1(n2801), .A2(n2789), .ZN(n4177) );
  NAND2_X1 U35410 ( .A1(n2865), .A2(n4177), .ZN(n2793) );
  NAND2_X1 U35420 ( .A1(n2671), .A2(REG0_REG_19__SCAN_IN), .ZN(n2792) );
  NAND2_X1 U35430 ( .A1(n2241), .A2(REG1_REG_19__SCAN_IN), .ZN(n2791) );
  NAND2_X1 U35440 ( .A1(n2244), .A2(REG2_REG_19__SCAN_IN), .ZN(n2790) );
  OR2_X1 U35450 ( .A1(n2563), .A2(IR_REG_18__SCAN_IN), .ZN(n2794) );
  OAI21_X2 U35460 ( .B1(n2795), .B2(n5040), .A(n2861), .ZN(n3980) );
  INV_X1 U35470 ( .A(DATAI_19_), .ZN(n4981) );
  NAND2_X1 U35480 ( .A1(n4296), .A2(n4176), .ZN(n3849) );
  INV_X1 U35490 ( .A(n4296), .ZN(n4185) );
  INV_X1 U35500 ( .A(n4176), .ZN(n3562) );
  INV_X1 U35510 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3728) );
  XNOR2_X1 U35520 ( .A(n2801), .B(n3728), .ZN(n4153) );
  NAND2_X1 U35530 ( .A1(n2865), .A2(n4153), .ZN(n2799) );
  NAND2_X1 U35540 ( .A1(n2244), .A2(REG2_REG_20__SCAN_IN), .ZN(n2798) );
  NAND2_X1 U35550 ( .A1(n2671), .A2(REG0_REG_20__SCAN_IN), .ZN(n2797) );
  NAND2_X1 U35560 ( .A1(n2240), .A2(REG1_REG_20__SCAN_IN), .ZN(n2796) );
  NAND4_X1 U35570 ( .A1(n2799), .A2(n2798), .A3(n2797), .A4(n2796), .ZN(n4121)
         );
  NAND2_X1 U35580 ( .A1(n4121), .A2(n4292), .ZN(n3851) );
  NOR2_X1 U35590 ( .A1(n4121), .A2(n4292), .ZN(n3852) );
  AND2_X1 U35600 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2800) );
  AOI21_X1 U35610 ( .B1(n2801), .B2(REG3_REG_20__SCAN_IN), .A(
        REG3_REG_21__SCAN_IN), .ZN(n2802) );
  OR2_X1 U35620 ( .A1(n2808), .A2(n2802), .ZN(n4135) );
  INV_X1 U35630 ( .A(n4135), .ZN(n3679) );
  NAND2_X1 U35640 ( .A1(n2865), .A2(n3679), .ZN(n2806) );
  NAND2_X1 U35650 ( .A1(n2671), .A2(REG0_REG_21__SCAN_IN), .ZN(n2805) );
  NAND2_X1 U35660 ( .A1(n2241), .A2(REG1_REG_21__SCAN_IN), .ZN(n2804) );
  NAND2_X1 U35670 ( .A1(n2244), .A2(REG2_REG_21__SCAN_IN), .ZN(n2803) );
  NAND4_X1 U35680 ( .A1(n2806), .A2(n2805), .A3(n2804), .A4(n2803), .ZN(n4293)
         );
  INV_X1 U35690 ( .A(n4293), .ZN(n4108) );
  NAND2_X1 U35700 ( .A1(n2835), .A2(DATAI_21_), .ZN(n4132) );
  NOR2_X1 U35710 ( .A1(n4108), .A2(n4132), .ZN(n2807) );
  OR2_X1 U35720 ( .A1(n2808), .A2(REG3_REG_22__SCAN_IN), .ZN(n2809) );
  AND2_X1 U35730 ( .A1(n2817), .A2(n2809), .ZN(n4113) );
  NAND2_X1 U35740 ( .A1(n2865), .A2(n4113), .ZN(n2813) );
  NAND2_X1 U35750 ( .A1(n2671), .A2(REG0_REG_22__SCAN_IN), .ZN(n2812) );
  NAND2_X1 U35760 ( .A1(n2242), .A2(REG1_REG_22__SCAN_IN), .ZN(n2811) );
  NAND2_X1 U35770 ( .A1(n2239), .A2(REG2_REG_22__SCAN_IN), .ZN(n2810) );
  NAND4_X1 U35780 ( .A1(n2813), .A2(n2812), .A3(n2811), .A4(n2810), .ZN(n4129)
         );
  NAND2_X1 U35790 ( .A1(n4129), .A2(n4112), .ZN(n2895) );
  INV_X1 U35800 ( .A(n2895), .ZN(n2814) );
  NOR2_X1 U35810 ( .A1(n4129), .A2(n4112), .ZN(n3901) );
  INV_X1 U3582 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3659) );
  NAND2_X1 U3583 ( .A1(n2817), .A2(n3659), .ZN(n2818) );
  AND2_X1 U3584 ( .A1(n2824), .A2(n2818), .ZN(n4094) );
  NAND2_X1 U3585 ( .A1(n2865), .A2(n4094), .ZN(n2822) );
  NAND2_X1 U3586 ( .A1(n2671), .A2(REG0_REG_23__SCAN_IN), .ZN(n2821) );
  NAND2_X1 U3587 ( .A1(n2240), .A2(REG1_REG_23__SCAN_IN), .ZN(n2820) );
  NAND2_X1 U3588 ( .A1(n2239), .A2(REG2_REG_23__SCAN_IN), .ZN(n2819) );
  INV_X1 U3589 ( .A(n3592), .ZN(n4092) );
  INV_X1 U3590 ( .A(n4276), .ZN(n4067) );
  INV_X1 U3591 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3717) );
  NAND2_X1 U3592 ( .A1(n2824), .A2(n3717), .ZN(n2825) );
  AND2_X1 U3593 ( .A1(n2831), .A2(n2825), .ZN(n4068) );
  NAND2_X1 U3594 ( .A1(n4068), .A2(n2865), .ZN(n2829) );
  NAND2_X1 U3595 ( .A1(n2239), .A2(REG2_REG_24__SCAN_IN), .ZN(n2828) );
  NAND2_X1 U3596 ( .A1(n2671), .A2(REG0_REG_24__SCAN_IN), .ZN(n2827) );
  NAND2_X1 U3597 ( .A1(n2240), .A2(REG1_REG_24__SCAN_IN), .ZN(n2826) );
  NAND4_X1 U3598 ( .A1(n2829), .A2(n2828), .A3(n2827), .A4(n2826), .ZN(n4264)
         );
  NAND2_X1 U3599 ( .A1(n4264), .A2(n4272), .ZN(n2830) );
  INV_X1 U3600 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4930) );
  AND2_X1 U3601 ( .A1(n2831), .A2(n4930), .ZN(n2832) );
  OR2_X1 U3602 ( .A1(n2832), .A2(n2844), .ZN(n3689) );
  AOI22_X1 U3603 ( .A1(n2242), .A2(REG1_REG_25__SCAN_IN), .B1(n2671), .B2(
        REG0_REG_25__SCAN_IN), .ZN(n2834) );
  NAND2_X1 U3604 ( .A1(n2244), .A2(REG2_REG_25__SCAN_IN), .ZN(n2833) );
  OAI211_X1 U3605 ( .C1(n3689), .C2(n2846), .A(n2834), .B(n2833), .ZN(n4273)
         );
  INV_X1 U3606 ( .A(n4273), .ZN(n3758) );
  NAND2_X1 U3607 ( .A1(n2835), .A2(DATAI_25_), .ZN(n4052) );
  NAND2_X1 U3608 ( .A1(n3758), .A2(n4052), .ZN(n2836) );
  AOI22_X2 U3609 ( .A1(n4047), .A2(n2836), .B1(n4263), .B2(n4273), .ZN(n4035)
         );
  INV_X1 U3610 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3759) );
  XNOR2_X1 U3611 ( .A(n2844), .B(n3759), .ZN(n4039) );
  NAND2_X1 U3612 ( .A1(n4039), .A2(n2865), .ZN(n2841) );
  NAND2_X1 U3613 ( .A1(n2241), .A2(REG1_REG_26__SCAN_IN), .ZN(n2839) );
  NAND2_X1 U3614 ( .A1(n2239), .A2(REG2_REG_26__SCAN_IN), .ZN(n2838) );
  NAND2_X1 U3615 ( .A1(n2671), .A2(REG0_REG_26__SCAN_IN), .ZN(n2837) );
  NAND2_X1 U3616 ( .A1(n4251), .A2(n4255), .ZN(n3867) );
  NOR2_X1 U3617 ( .A1(n4251), .A2(n4255), .ZN(n3869) );
  NAND2_X1 U3618 ( .A1(n2844), .A2(REG3_REG_26__SCAN_IN), .ZN(n2842) );
  INV_X1 U3619 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3650) );
  NAND2_X1 U3620 ( .A1(n2842), .A2(n3650), .ZN(n2845) );
  AND2_X1 U3621 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2843) );
  NAND2_X1 U3622 ( .A1(n2844), .A2(n2843), .ZN(n2853) );
  NAND2_X1 U3623 ( .A1(n2845), .A2(n2853), .ZN(n3649) );
  AOI22_X1 U3624 ( .A1(n2242), .A2(REG1_REG_27__SCAN_IN), .B1(n2671), .B2(
        REG0_REG_27__SCAN_IN), .ZN(n2848) );
  NAND2_X1 U3625 ( .A1(n2244), .A2(REG2_REG_27__SCAN_IN), .ZN(n2847) );
  INV_X1 U3626 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4973) );
  NAND2_X1 U3627 ( .A1(n2853), .A2(n4973), .ZN(n2854) );
  NAND2_X1 U3628 ( .A1(n4009), .A2(n2865), .ZN(n2859) );
  NAND2_X1 U3629 ( .A1(n2241), .A2(REG1_REG_28__SCAN_IN), .ZN(n2857) );
  NAND2_X1 U3630 ( .A1(n2239), .A2(REG2_REG_28__SCAN_IN), .ZN(n2856) );
  NAND2_X1 U3631 ( .A1(n2671), .A2(REG0_REG_28__SCAN_IN), .ZN(n2855) );
  NAND2_X1 U3632 ( .A1(n2835), .A2(DATAI_28_), .ZN(n4012) );
  NOR2_X1 U3633 ( .A1(n4023), .A2(n4012), .ZN(n3985) );
  NAND2_X1 U3634 ( .A1(n4023), .A2(n4012), .ZN(n3986) );
  INV_X1 U3635 ( .A(n3986), .ZN(n2860) );
  XNOR2_X1 U3636 ( .A(n3993), .B(n3992), .ZN(n4017) );
  XNOR2_X1 U3637 ( .A(n3002), .B(n3928), .ZN(n2864) );
  NAND2_X1 U3638 ( .A1(n2864), .A2(n3980), .ZN(n3495) );
  INV_X1 U3639 ( .A(n3928), .ZN(n2869) );
  INV_X1 U3640 ( .A(n3980), .ZN(n3109) );
  INV_X1 U3641 ( .A(n4617), .ZN(n4609) );
  NAND2_X1 U3642 ( .A1(n3495), .A2(n4609), .ZN(n4646) );
  AOI22_X1 U3643 ( .A1(n2244), .A2(REG2_REG_29__SCAN_IN), .B1(n2671), .B2(
        REG0_REG_29__SCAN_IN), .ZN(n2867) );
  NAND2_X1 U3644 ( .A1(n2240), .A2(REG1_REG_29__SCAN_IN), .ZN(n2866) );
  OAI211_X1 U3645 ( .C1(n3984), .C2(n2846), .A(n2867), .B(n2866), .ZN(n4008)
         );
  INV_X1 U3646 ( .A(n4008), .ZN(n2870) );
  INV_X1 U3647 ( .A(n3920), .ZN(n2918) );
  INV_X1 U3648 ( .A(n2922), .ZN(n3923) );
  NAND2_X1 U3649 ( .A1(n3074), .A2(n3923), .ZN(n4593) );
  OAI22_X1 U3650 ( .A1(n2870), .A2(n4594), .B1(n4593), .B2(n4012), .ZN(n2903)
         );
  NAND2_X1 U3651 ( .A1(n3024), .A2(n4670), .ZN(n3075) );
  INV_X1 U3652 ( .A(n3938), .ZN(n3146) );
  NAND2_X1 U3653 ( .A1(n3146), .A2(n3132), .ZN(n3787) );
  NAND2_X1 U3654 ( .A1(n3938), .A2(n3156), .ZN(n3784) );
  AND2_X1 U3655 ( .A1(n3787), .A2(n3784), .ZN(n3873) );
  NAND2_X1 U3656 ( .A1(n3064), .A2(n3873), .ZN(n2874) );
  INV_X1 U3657 ( .A(n3788), .ZN(n2875) );
  INV_X1 U3658 ( .A(n3167), .ZN(n3172) );
  AND2_X1 U3659 ( .A1(n3936), .A2(n3172), .ZN(n3093) );
  INV_X1 U3660 ( .A(n3936), .ZN(n3257) );
  NAND2_X1 U3661 ( .A1(n3257), .A2(n3167), .ZN(n3802) );
  NAND2_X1 U3662 ( .A1(n3935), .A2(n3206), .ZN(n3804) );
  NAND2_X1 U3663 ( .A1(n3254), .A2(n3804), .ZN(n2876) );
  INV_X1 U3664 ( .A(n3935), .ZN(n3246) );
  NAND2_X1 U3665 ( .A1(n3246), .A2(n3264), .ZN(n3793) );
  NAND2_X1 U3666 ( .A1(n2876), .A2(n3793), .ZN(n3179) );
  INV_X1 U3667 ( .A(n2877), .ZN(n2878) );
  NAND2_X1 U3668 ( .A1(n3313), .A2(n3283), .ZN(n3798) );
  NAND2_X1 U3669 ( .A1(n3249), .A2(n3526), .ZN(n3795) );
  NAND2_X1 U3670 ( .A1(n3363), .A2(n3227), .ZN(n3797) );
  NAND2_X1 U3671 ( .A1(n2880), .A2(n3797), .ZN(n3270) );
  NAND2_X1 U3672 ( .A1(n4638), .A2(n3364), .ZN(n3813) );
  NAND2_X1 U3673 ( .A1(n3270), .A2(n3813), .ZN(n2881) );
  NAND2_X1 U3674 ( .A1(n3383), .A2(n3356), .ZN(n3812) );
  NAND2_X1 U3675 ( .A1(n4636), .A2(n3425), .ZN(n3406) );
  NAND2_X1 U3676 ( .A1(n3514), .A2(n3447), .ZN(n3401) );
  NAND2_X1 U3677 ( .A1(n3406), .A2(n3401), .ZN(n3817) );
  NAND2_X1 U3678 ( .A1(n3426), .A2(n3429), .ZN(n3405) );
  NAND2_X1 U3679 ( .A1(n3343), .A2(n3405), .ZN(n2883) );
  INV_X1 U3680 ( .A(n3817), .ZN(n2882) );
  NOR2_X1 U3681 ( .A1(n3514), .A2(n3447), .ZN(n3402) );
  AOI21_X1 U3682 ( .B1(n2883), .B2(n2882), .A(n3402), .ZN(n3821) );
  INV_X1 U3683 ( .A(n3878), .ZN(n3490) );
  NAND2_X1 U3684 ( .A1(n3491), .A2(n3490), .ZN(n3492) );
  INV_X1 U3685 ( .A(n4325), .ZN(n3699) );
  NAND2_X1 U3686 ( .A1(n3699), .A2(n3541), .ZN(n3819) );
  NAND2_X1 U3687 ( .A1(n4325), .A2(n3770), .ZN(n3801) );
  NAND2_X1 U3688 ( .A1(n3819), .A2(n3801), .ZN(n3881) );
  INV_X1 U3689 ( .A(n3820), .ZN(n2884) );
  NOR2_X1 U3690 ( .A1(n3881), .A2(n2884), .ZN(n2885) );
  NAND2_X1 U3691 ( .A1(n3492), .A2(n2885), .ZN(n2886) );
  NAND2_X1 U3692 ( .A1(n2886), .A2(n3801), .ZN(n3475) );
  NAND2_X1 U3693 ( .A1(n3475), .A2(n3481), .ZN(n2887) );
  NAND2_X1 U3694 ( .A1(n4185), .A2(n4176), .ZN(n2888) );
  AND2_X1 U3695 ( .A1(n4165), .A2(n2888), .ZN(n4080) );
  INV_X1 U3696 ( .A(n4292), .ZN(n4149) );
  NAND2_X1 U3697 ( .A1(n4121), .A2(n4149), .ZN(n4081) );
  NAND2_X1 U3698 ( .A1(n3745), .A2(n4208), .ZN(n4078) );
  AND2_X1 U3699 ( .A1(n4081), .A2(n4078), .ZN(n2889) );
  NAND2_X1 U3700 ( .A1(n4080), .A2(n2889), .ZN(n3893) );
  NAND2_X1 U3701 ( .A1(n4187), .A2(n4215), .ZN(n4162) );
  NAND2_X1 U3702 ( .A1(n4167), .A2(n4162), .ZN(n2890) );
  NAND2_X1 U3703 ( .A1(n2890), .A2(n4080), .ZN(n2892) );
  NAND2_X1 U3704 ( .A1(n4296), .A2(n3562), .ZN(n2891) );
  NAND2_X1 U3705 ( .A1(n2892), .A2(n2891), .ZN(n4140) );
  NOR2_X1 U3706 ( .A1(n4121), .A2(n4149), .ZN(n2893) );
  OR2_X1 U3707 ( .A1(n4140), .A2(n2893), .ZN(n2894) );
  NAND2_X1 U3708 ( .A1(n2894), .A2(n4081), .ZN(n3825) );
  NAND2_X1 U3709 ( .A1(n4108), .A2(n4128), .ZN(n4083) );
  AND2_X1 U3710 ( .A1(n3825), .A2(n4083), .ZN(n3898) );
  NAND2_X1 U3711 ( .A1(n4293), .A2(n4132), .ZN(n3903) );
  INV_X1 U3712 ( .A(n3901), .ZN(n4084) );
  OR2_X1 U3713 ( .A1(n4276), .A2(n3592), .ZN(n3847) );
  AND2_X1 U3714 ( .A1(n3847), .A2(n2895), .ZN(n3829) );
  NAND2_X1 U3715 ( .A1(n2896), .A2(n3829), .ZN(n4060) );
  NAND2_X1 U3716 ( .A1(n4087), .A2(n4272), .ZN(n3846) );
  NAND2_X1 U3717 ( .A1(n4276), .A2(n3592), .ZN(n4059) );
  NAND2_X1 U3718 ( .A1(n3846), .A2(n4059), .ZN(n3900) );
  INV_X1 U3719 ( .A(n3900), .ZN(n3827) );
  NAND2_X1 U3720 ( .A1(n4060), .A2(n3827), .ZN(n2897) );
  NAND2_X1 U3721 ( .A1(n4264), .A2(n4072), .ZN(n3845) );
  NAND2_X1 U3722 ( .A1(n4273), .A2(n4052), .ZN(n3871) );
  INV_X1 U3723 ( .A(n3871), .ZN(n2898) );
  OR2_X1 U3724 ( .A1(n4273), .A2(n4052), .ZN(n3872) );
  NOR2_X1 U3725 ( .A1(n4251), .A2(n4042), .ZN(n3778) );
  AND2_X1 U3726 ( .A1(n4251), .A2(n4042), .ZN(n3832) );
  NOR2_X1 U3727 ( .A1(n4258), .A2(n2899), .ZN(n3834) );
  XNOR2_X1 U3728 ( .A(n3987), .B(n3992), .ZN(n2902) );
  NAND2_X1 U3729 ( .A1(n3928), .A2(n3109), .ZN(n2901) );
  NAND2_X1 U3730 ( .A1(n3923), .A2(n3920), .ZN(n2900) );
  NOR2_X1 U3731 ( .A1(n2902), .A2(n4213), .ZN(n4015) );
  NAND2_X1 U3732 ( .A1(n2917), .A2(n2920), .ZN(n2904) );
  MUX2_X1 U3733 ( .A(n2920), .B(n2904), .S(B_REG_SCAN_IN), .Z(n2906) );
  NOR4_X1 U3734 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n2915) );
  NOR4_X1 U3735 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2914) );
  INV_X1 U3736 ( .A(D_REG_17__SCAN_IN), .ZN(n4567) );
  INV_X1 U3737 ( .A(D_REG_14__SCAN_IN), .ZN(n4569) );
  INV_X1 U3738 ( .A(D_REG_19__SCAN_IN), .ZN(n4856) );
  INV_X1 U3739 ( .A(D_REG_15__SCAN_IN), .ZN(n4568) );
  NAND4_X1 U3740 ( .A1(n4567), .A2(n4569), .A3(n4856), .A4(n4568), .ZN(n2912)
         );
  NOR4_X1 U3741 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2910) );
  NOR4_X1 U3742 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2909) );
  NOR4_X1 U3743 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2908) );
  NOR4_X1 U3744 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_22__SCAN_IN), .ZN(n2907) );
  NAND4_X1 U3745 ( .A1(n2910), .A2(n2909), .A3(n2908), .A4(n2907), .ZN(n2911)
         );
  NOR4_X1 U3746 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(n2912), 
        .A4(n2911), .ZN(n2913) );
  AND3_X1 U3747 ( .A1(n2915), .A2(n2914), .A3(n2913), .ZN(n2916) );
  NOR2_X1 U3748 ( .A1(n2964), .A2(n2916), .ZN(n2989) );
  AND2_X1 U3749 ( .A1(n2922), .A2(n3980), .ZN(n3010) );
  NOR2_X1 U3750 ( .A1(n3008), .A2(n3010), .ZN(n3121) );
  OR2_X1 U3751 ( .A1(n3016), .A2(n3121), .ZN(n2994) );
  NOR2_X1 U3752 ( .A1(n2989), .A2(n2994), .ZN(n2931) );
  INV_X1 U3753 ( .A(n2917), .ZN(n4380) );
  OAI22_X1 U3754 ( .A1(n2964), .A2(D_REG_1__SCAN_IN), .B1(n2905), .B2(n4380), 
        .ZN(n2990) );
  NAND2_X1 U3755 ( .A1(n4617), .A2(n2918), .ZN(n2932) );
  AND2_X1 U3756 ( .A1(n2990), .A2(n2932), .ZN(n2919) );
  INV_X1 U3757 ( .A(n2920), .ZN(n4381) );
  INV_X1 U3758 ( .A(n2929), .ZN(n2991) );
  NAND2_X1 U3759 ( .A1(n4602), .A2(n3156), .ZN(n3106) );
  NAND2_X1 U3760 ( .A1(n4022), .A2(n3994), .ZN(n2921) );
  NAND2_X1 U3761 ( .A1(n4000), .A2(n2921), .ZN(n4007) );
  NAND2_X1 U3762 ( .A1(n2923), .A2(n2478), .ZN(U3546) );
  MUX2_X1 U3763 ( .A(REG0_REG_28__SCAN_IN), .B(n2925), .S(n4649), .Z(n2926) );
  INV_X1 U3764 ( .A(n2926), .ZN(n2927) );
  NAND2_X1 U3765 ( .A1(n2927), .A2(n2477), .ZN(U3514) );
  INV_X1 U3766 ( .A(n4572), .ZN(n2967) );
  INV_X1 U3767 ( .A(n3075), .ZN(n3781) );
  XNOR2_X1 U3768 ( .A(n2872), .B(n3781), .ZN(n2928) );
  NOR2_X1 U3769 ( .A1(n2928), .A2(n4213), .ZN(n4600) );
  INV_X1 U3770 ( .A(n2990), .ZN(n2930) );
  NAND3_X1 U3771 ( .A1(n2931), .A2(n2930), .A3(n2929), .ZN(n2933) );
  MUX2_X1 U3772 ( .A(REG2_REG_1__SCAN_IN), .B(n4600), .S(n4402), .Z(n2943) );
  OAI21_X1 U3773 ( .B1(n2872), .B2(n2935), .A(n2934), .ZN(n4591) );
  OR2_X1 U3774 ( .A1(n3002), .A2(n3980), .ZN(n3033) );
  NAND2_X1 U3775 ( .A1(n3495), .A2(n3033), .ZN(n2936) );
  INV_X1 U3776 ( .A(n4201), .ZN(n4223) );
  AND2_X1 U3777 ( .A1(n4402), .A2(n4637), .ZN(n4066) );
  INV_X1 U3778 ( .A(n4066), .ZN(n4156) );
  OAI22_X1 U3779 ( .A1(n4591), .A2(n4223), .B1(n3024), .B2(n4156), .ZN(n2942)
         );
  NAND2_X1 U3780 ( .A1(n4314), .A2(n3980), .ZN(n3000) );
  INV_X1 U3781 ( .A(n3000), .ZN(n2937) );
  NAND2_X1 U3782 ( .A1(n3026), .A2(n4670), .ZN(n2938) );
  NAND2_X1 U3783 ( .A1(n3044), .A2(n2938), .ZN(n4596) );
  INV_X1 U3784 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3029) );
  OAI22_X1 U3785 ( .A1(n4220), .A2(n4596), .B1(n3029), .B2(n4134), .ZN(n2941)
         );
  AND2_X1 U3786 ( .A1(n4402), .A2(n4635), .ZN(n4151) );
  INV_X1 U3787 ( .A(n4151), .ZN(n2939) );
  NAND2_X1 U3788 ( .A1(n4402), .A2(n4634), .ZN(n4071) );
  OAI22_X1 U3789 ( .A1(n2939), .A2(n2680), .B1(n4071), .B2(n4592), .ZN(n2940)
         );
  OR4_X1 U3790 ( .A1(n2943), .A2(n2942), .A3(n2941), .A4(n2940), .ZN(U3289) );
  INV_X1 U3791 ( .A(DATAI_1_), .ZN(n2944) );
  MUX2_X1 U3792 ( .A(n2945), .B(n2944), .S(U3149), .Z(n2946) );
  INV_X1 U3793 ( .A(n2946), .ZN(U3351) );
  INV_X1 U3794 ( .A(DATAI_14_), .ZN(n2948) );
  NAND2_X1 U3795 ( .A1(n4537), .A2(STATE_REG_SCAN_IN), .ZN(n2947) );
  OAI21_X1 U3796 ( .B1(STATE_REG_SCAN_IN), .B2(n2948), .A(n2947), .ZN(U3338)
         );
  INV_X1 U3797 ( .A(DATAI_15_), .ZN(n4957) );
  NAND2_X1 U3798 ( .A1(n3950), .A2(STATE_REG_SCAN_IN), .ZN(n2949) );
  OAI21_X1 U3799 ( .B1(STATE_REG_SCAN_IN), .B2(n4957), .A(n2949), .ZN(U3337)
         );
  INV_X1 U3800 ( .A(DATAI_21_), .ZN(n2951) );
  NAND2_X1 U3801 ( .A1(n3920), .A2(STATE_REG_SCAN_IN), .ZN(n2950) );
  OAI21_X1 U3802 ( .B1(STATE_REG_SCAN_IN), .B2(n2951), .A(n2950), .ZN(U3331)
         );
  MUX2_X1 U3803 ( .A(n3980), .B(n4981), .S(U3149), .Z(n2952) );
  INV_X1 U3804 ( .A(n2952), .ZN(U3333) );
  INV_X1 U3805 ( .A(DATAI_22_), .ZN(n4935) );
  NAND2_X1 U3806 ( .A1(n3928), .A2(STATE_REG_SCAN_IN), .ZN(n2953) );
  OAI21_X1 U3807 ( .B1(STATE_REG_SCAN_IN), .B2(n4935), .A(n2953), .ZN(U3330)
         );
  INV_X1 U3808 ( .A(DATAI_20_), .ZN(n2955) );
  NAND2_X1 U3809 ( .A1(n3923), .A2(STATE_REG_SCAN_IN), .ZN(n2954) );
  OAI21_X1 U3810 ( .B1(STATE_REG_SCAN_IN), .B2(n2955), .A(n2954), .ZN(U3332)
         );
  INV_X1 U3811 ( .A(DATAI_29_), .ZN(n2958) );
  NAND2_X1 U3812 ( .A1(n2956), .A2(STATE_REG_SCAN_IN), .ZN(n2957) );
  OAI21_X1 U3813 ( .B1(STATE_REG_SCAN_IN), .B2(n2958), .A(n2957), .ZN(U3323)
         );
  INV_X1 U3814 ( .A(DATAI_31_), .ZN(n4822) );
  OR4_X1 U3815 ( .A1(n2960), .A2(IR_REG_30__SCAN_IN), .A3(n2959), .A4(U3149), 
        .ZN(n2961) );
  OAI21_X1 U3816 ( .B1(STATE_REG_SCAN_IN), .B2(n4822), .A(n2961), .ZN(U3321)
         );
  INV_X1 U3817 ( .A(DATAI_28_), .ZN(n4821) );
  NAND2_X1 U3818 ( .A1(n3021), .A2(STATE_REG_SCAN_IN), .ZN(n2962) );
  OAI21_X1 U3819 ( .B1(STATE_REG_SCAN_IN), .B2(n4821), .A(n2962), .ZN(U3324)
         );
  INV_X1 U3820 ( .A(DATAI_27_), .ZN(n4982) );
  NAND2_X1 U3821 ( .A1(n4416), .A2(STATE_REG_SCAN_IN), .ZN(n2963) );
  OAI21_X1 U3822 ( .B1(STATE_REG_SCAN_IN), .B2(n4982), .A(n2963), .ZN(U3325)
         );
  INV_X1 U3823 ( .A(n3016), .ZN(n3009) );
  INV_X1 U3824 ( .A(D_REG_1__SCAN_IN), .ZN(n2966) );
  NOR3_X1 U3825 ( .A1(n2967), .A2(n2905), .A3(n4380), .ZN(n2965) );
  AOI21_X1 U3826 ( .B1(n4570), .B2(n2966), .A(n2965), .ZN(U3459) );
  INV_X1 U3827 ( .A(D_REG_0__SCAN_IN), .ZN(n2969) );
  NOR3_X1 U3828 ( .A1(n2967), .A2(n2905), .A3(n4381), .ZN(n2968) );
  AOI21_X1 U3829 ( .B1(n4570), .B2(n2969), .A(n2968), .ZN(U3458) );
  NOR2_X1 U3830 ( .A1(n4543), .A2(U4043), .ZN(U3148) );
  INV_X1 U3831 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n4995) );
  NAND2_X1 U3832 ( .A1(n3428), .A2(U4043), .ZN(n2970) );
  OAI21_X1 U3833 ( .B1(U4043), .B2(n4995), .A(n2970), .ZN(U3561) );
  INV_X1 U3834 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n5024) );
  NAND2_X1 U3835 ( .A1(n2971), .A2(U4043), .ZN(n2972) );
  OAI21_X1 U3836 ( .B1(U4043), .B2(n5024), .A(n2972), .ZN(U3550) );
  INV_X1 U3837 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n4904) );
  NAND2_X1 U3838 ( .A1(n4264), .A2(U4043), .ZN(n2973) );
  OAI21_X1 U3839 ( .B1(U4043), .B2(n4904), .A(n2973), .ZN(U3574) );
  INV_X1 U3840 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n4902) );
  NAND2_X1 U3841 ( .A1(n3249), .A2(U4043), .ZN(n2974) );
  OAI21_X1 U3842 ( .B1(U4043), .B2(n4902), .A(n2974), .ZN(U3558) );
  INV_X1 U3843 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4910) );
  NAND2_X1 U3844 ( .A1(n2241), .A2(REG1_REG_30__SCAN_IN), .ZN(n2977) );
  NAND2_X1 U3845 ( .A1(n2239), .A2(REG2_REG_30__SCAN_IN), .ZN(n2976) );
  NAND2_X1 U3846 ( .A1(n2671), .A2(REG0_REG_30__SCAN_IN), .ZN(n2975) );
  AND3_X1 U3847 ( .A1(n2977), .A2(n2976), .A3(n2975), .ZN(n3989) );
  INV_X1 U3848 ( .A(n3989), .ZN(n2978) );
  NAND2_X1 U3849 ( .A1(n2978), .A2(U4043), .ZN(n2979) );
  OAI21_X1 U3850 ( .B1(U4043), .B2(n4910), .A(n2979), .ZN(U3580) );
  INV_X1 U3851 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n5048) );
  NAND2_X1 U3852 ( .A1(n4067), .A2(U4043), .ZN(n2980) );
  OAI21_X1 U3853 ( .B1(U4043), .B2(n5048), .A(n2980), .ZN(U3573) );
  INV_X1 U3854 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4932) );
  NAND2_X1 U3855 ( .A1(n2239), .A2(REG2_REG_31__SCAN_IN), .ZN(n2983) );
  NAND2_X1 U3856 ( .A1(n2242), .A2(REG1_REG_31__SCAN_IN), .ZN(n2982) );
  NAND2_X1 U3857 ( .A1(n2671), .A2(REG0_REG_31__SCAN_IN), .ZN(n2981) );
  NAND3_X1 U3858 ( .A1(n2983), .A2(n2982), .A3(n2981), .ZN(n3914) );
  NAND2_X1 U3859 ( .A1(n3914), .A2(U4043), .ZN(n2984) );
  OAI21_X1 U3860 ( .B1(U4043), .B2(n4932), .A(n2984), .ZN(U3581) );
  INV_X1 U3861 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n5012) );
  NAND2_X1 U3862 ( .A1(n3514), .A2(U4043), .ZN(n2985) );
  OAI21_X1 U3863 ( .B1(U4043), .B2(n5012), .A(n2985), .ZN(U3563) );
  INV_X1 U3864 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n4998) );
  NAND2_X1 U3865 ( .A1(n3255), .A2(U4043), .ZN(n2986) );
  OAI21_X1 U3866 ( .B1(U4043), .B2(n4998), .A(n2986), .ZN(U3557) );
  INV_X1 U3867 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4996) );
  NAND2_X1 U3868 ( .A1(n4251), .A2(U4043), .ZN(n2987) );
  OAI21_X1 U3869 ( .B1(U4043), .B2(n4996), .A(n2987), .ZN(U3576) );
  INV_X1 U3870 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4929) );
  NAND2_X1 U3871 ( .A1(n3745), .A2(U4043), .ZN(n2988) );
  OAI21_X1 U3872 ( .B1(U4043), .B2(n4929), .A(n2988), .ZN(U3567) );
  INV_X1 U3873 ( .A(n3074), .ZN(n4584) );
  NOR2_X1 U3874 ( .A1(n4584), .A2(n3980), .ZN(n2993) );
  NOR2_X1 U3875 ( .A1(n2990), .A2(n2989), .ZN(n2992) );
  AOI21_X1 U3876 ( .B1(n4593), .B2(n2993), .A(n3023), .ZN(n3124) );
  INV_X1 U3877 ( .A(n3124), .ZN(n2996) );
  INV_X1 U3878 ( .A(n2994), .ZN(n2995) );
  AND2_X1 U3879 ( .A1(n2996), .A2(n2995), .ZN(n4675) );
  INV_X1 U3880 ( .A(n3002), .ZN(n2997) );
  INV_X2 U3881 ( .A(n2253), .ZN(n3623) );
  INV_X1 U3882 ( .A(n2998), .ZN(n3123) );
  NOR2_X1 U3883 ( .A1(n3001), .A2(n2999), .ZN(n4413) );
  AOI222_X1 U3884 ( .A1(n2971), .A2(n3166), .B1(n2253), .B2(n4670), .C1(n3123), 
        .C2(IR_REG_0__SCAN_IN), .ZN(n4414) );
  INV_X1 U3885 ( .A(n3001), .ZN(n3004) );
  OR2_X1 U3886 ( .A1(n3076), .A2(n3624), .ZN(n3006) );
  NAND2_X1 U3887 ( .A1(n3026), .A2(n2253), .ZN(n3005) );
  NAND2_X1 U3888 ( .A1(n3006), .A2(n3005), .ZN(n3052) );
  OAI22_X1 U3889 ( .A1(n3076), .A2(n3623), .B1(n3620), .B2(n4592), .ZN(n3007)
         );
  XNOR2_X1 U3890 ( .A(n3007), .B(n3601), .ZN(n3053) );
  XNOR2_X1 U3891 ( .A(n3052), .B(n3053), .ZN(n3013) );
  INV_X1 U3892 ( .A(n3023), .ZN(n3012) );
  OAI211_X1 U3893 ( .C1(n3010), .C2(n4584), .A(n3009), .B(n3008), .ZN(n3011)
         );
  AOI211_X1 U3894 ( .C1(n3014), .C2(n3013), .A(n3775), .B(n3054), .ZN(n3015)
         );
  INV_X1 U3895 ( .A(n3015), .ZN(n3028) );
  NOR2_X1 U3896 ( .A1(n3016), .A2(n4593), .ZN(n3017) );
  INV_X1 U3897 ( .A(n2237), .ZN(n4671) );
  NAND2_X1 U3898 ( .A1(n4572), .A2(n3018), .ZN(n3019) );
  NOR2_X1 U3899 ( .A1(n3927), .A2(n4415), .ZN(n3020) );
  NOR2_X1 U3900 ( .A1(n3021), .A2(n3927), .ZN(n3022) );
  OAI22_X1 U3901 ( .A1(n3024), .A2(n3768), .B1(n2680), .B2(n3760), .ZN(n3025)
         );
  AOI21_X1 U3902 ( .B1(n3026), .B2(n4671), .A(n3025), .ZN(n3027) );
  OAI211_X1 U3903 ( .C1(n4675), .C2(n3029), .A(n3028), .B(n3027), .ZN(U3219)
         );
  NAND2_X1 U3904 ( .A1(n3031), .A2(n3035), .ZN(n3032) );
  NAND2_X1 U3905 ( .A1(n3030), .A2(n3032), .ZN(n4606) );
  INV_X1 U3906 ( .A(n4606), .ZN(n3049) );
  INV_X1 U3907 ( .A(n3033), .ZN(n3034) );
  NAND2_X1 U3908 ( .A1(n4402), .A2(n3034), .ZN(n3505) );
  XNOR2_X1 U3909 ( .A(n3036), .B(n2679), .ZN(n3042) );
  INV_X1 U3910 ( .A(n3495), .ZN(n3037) );
  NAND2_X1 U3911 ( .A1(n4606), .A2(n3037), .ZN(n3041) );
  AOI22_X1 U3912 ( .A1(n3938), .A2(n4635), .B1(n3059), .B2(n4634), .ZN(n3038)
         );
  OAI21_X1 U3913 ( .B1(n3076), .B2(n4327), .A(n3038), .ZN(n3039) );
  INV_X1 U3914 ( .A(n3039), .ZN(n3040) );
  OAI211_X1 U3915 ( .C1(n3042), .C2(n4213), .A(n3041), .B(n3040), .ZN(n4604)
         );
  MUX2_X1 U3916 ( .A(n4604), .B(REG2_REG_2__SCAN_IN), .S(n4566), .Z(n3043) );
  INV_X1 U3917 ( .A(n3043), .ZN(n3048) );
  INV_X1 U3918 ( .A(n3044), .ZN(n3045) );
  NOR2_X1 U3919 ( .A1(n3045), .A2(n3050), .ZN(n4603) );
  NOR3_X1 U3920 ( .A1(n4220), .A2(n4603), .A3(n4602), .ZN(n3046) );
  AOI21_X1 U3921 ( .B1(n4557), .B2(REG3_REG_2__SCAN_IN), .A(n3046), .ZN(n3047)
         );
  OAI211_X1 U3922 ( .C1(n3049), .C2(n3505), .A(n3048), .B(n3047), .ZN(U3288)
         );
  INV_X1 U3923 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3062) );
  OAI22_X1 U3924 ( .A1(n2680), .A2(n3624), .B1(n3621), .B2(n3050), .ZN(n3127)
         );
  OAI22_X1 U3925 ( .A1(n2680), .A2(n3623), .B1(n3620), .B2(n3050), .ZN(n3051)
         );
  XNOR2_X1 U3926 ( .A(n3051), .B(n3601), .ZN(n3128) );
  XOR2_X1 U3927 ( .A(n3127), .B(n3128), .Z(n3056) );
  OAI21_X1 U3928 ( .B1(n3056), .B2(n3055), .A(n3130), .ZN(n3057) );
  NAND2_X1 U3929 ( .A1(n3057), .A2(n4667), .ZN(n3061) );
  OAI22_X1 U3930 ( .A1(n3146), .A2(n3760), .B1(n3076), .B2(n3768), .ZN(n3058)
         );
  AOI21_X1 U3931 ( .B1(n3059), .B2(n4671), .A(n3058), .ZN(n3060) );
  OAI211_X1 U3932 ( .C1(n4675), .C2(n3062), .A(n3061), .B(n3060), .ZN(U3234)
         );
  XNOR2_X1 U3933 ( .A(n3063), .B(n3873), .ZN(n4610) );
  XNOR2_X1 U3934 ( .A(n3064), .B(n3873), .ZN(n3067) );
  AOI22_X1 U3935 ( .A1(n3937), .A2(n4635), .B1(n4634), .B2(n3132), .ZN(n3065)
         );
  OAI21_X1 U3936 ( .B1(n2680), .B2(n4327), .A(n3065), .ZN(n3066) );
  AOI21_X1 U3937 ( .B1(n3067), .B2(n4189), .A(n3066), .ZN(n3068) );
  OAI21_X1 U3938 ( .B1(n4610), .B2(n3495), .A(n3068), .ZN(n4612) );
  INV_X1 U3939 ( .A(n4612), .ZN(n3073) );
  INV_X1 U3940 ( .A(n4610), .ZN(n3071) );
  INV_X1 U3941 ( .A(n3505), .ZN(n4561) );
  OAI21_X1 U3942 ( .B1(n4602), .B2(n3156), .A(n3106), .ZN(n4608) );
  INV_X1 U3943 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3155) );
  AOI22_X1 U3944 ( .A1(n4566), .A2(REG2_REG_3__SCAN_IN), .B1(n4557), .B2(n3155), .ZN(n3069) );
  OAI21_X1 U3945 ( .B1(n4608), .B2(n4220), .A(n3069), .ZN(n3070) );
  AOI21_X1 U3946 ( .B1(n3071), .B2(n4561), .A(n3070), .ZN(n3072) );
  OAI21_X1 U3947 ( .B1(n3073), .B2(n4204), .A(n3072), .ZN(U3287) );
  NAND2_X1 U3948 ( .A1(n4402), .A2(n3980), .ZN(n4199) );
  INV_X1 U3949 ( .A(n4199), .ZN(n3188) );
  INV_X1 U3950 ( .A(n4071), .ZN(n4152) );
  AOI21_X1 U3951 ( .B1(n3074), .B2(n3188), .A(n4152), .ZN(n3081) );
  NAND2_X1 U3952 ( .A1(n2971), .A2(n4585), .ZN(n3780) );
  NAND2_X1 U3953 ( .A1(n3075), .A2(n3780), .ZN(n4588) );
  INV_X1 U3954 ( .A(n4588), .ZN(n3078) );
  OAI22_X1 U3955 ( .A1(n3078), .A2(n4213), .B1(n3076), .B2(n4594), .ZN(n4586)
         );
  AOI22_X1 U3956 ( .A1(n4566), .A2(REG2_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(n4557), .ZN(n3077) );
  OAI21_X1 U3957 ( .B1(n3078), .B2(n4223), .A(n3077), .ZN(n3079) );
  AOI21_X1 U3958 ( .B1(n4586), .B2(n4402), .A(n3079), .ZN(n3080) );
  OAI21_X1 U3959 ( .B1(n3081), .B2(n4585), .A(n3080), .ZN(U3290) );
  INV_X1 U3960 ( .A(n4384), .ZN(n3092) );
  OAI211_X1 U3961 ( .C1(n3084), .C2(n3083), .A(n4551), .B(n3082), .ZN(n3091)
         );
  AND2_X1 U3962 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3316) );
  INV_X1 U3963 ( .A(n3085), .ZN(n3086) );
  AOI211_X1 U3964 ( .C1(n3088), .C2(n3087), .A(n3086), .B(n4531), .ZN(n3089)
         );
  AOI211_X1 U3965 ( .C1(n4543), .C2(ADDR_REG_9__SCAN_IN), .A(n3316), .B(n3089), 
        .ZN(n3090) );
  OAI211_X1 U3966 ( .C1(n4556), .C2(n3092), .A(n3091), .B(n3090), .ZN(U3249)
         );
  INV_X1 U3967 ( .A(n3093), .ZN(n3790) );
  AND2_X1 U3968 ( .A1(n3790), .A2(n3802), .ZN(n3857) );
  INV_X1 U3969 ( .A(n3857), .ZN(n3094) );
  XNOR2_X1 U3970 ( .A(n3095), .B(n3094), .ZN(n3098) );
  AOI22_X1 U3971 ( .A1(n3935), .A2(n4635), .B1(n4634), .B2(n3167), .ZN(n3096)
         );
  OAI21_X1 U3972 ( .B1(n3171), .B2(n4327), .A(n3096), .ZN(n3097) );
  AOI21_X1 U3973 ( .B1(n3098), .B2(n4189), .A(n3097), .ZN(n4620) );
  XNOR2_X1 U3974 ( .A(n3099), .B(n3857), .ZN(n4623) );
  INV_X1 U3975 ( .A(n3107), .ZN(n3101) );
  INV_X1 U3976 ( .A(n3100), .ZN(n3263) );
  OAI21_X1 U3977 ( .B1(n3101), .B2(n3172), .A(n3263), .ZN(n4621) );
  AOI22_X1 U3978 ( .A1(n4566), .A2(REG2_REG_5__SCAN_IN), .B1(n3102), .B2(n4557), .ZN(n3103) );
  OAI21_X1 U3979 ( .B1(n4621), .B2(n4220), .A(n3103), .ZN(n3104) );
  AOI21_X1 U3980 ( .B1(n4623), .B2(n4201), .A(n3104), .ZN(n3105) );
  OAI21_X1 U3981 ( .B1(n4620), .B2(n4566), .A(n3105), .ZN(U3285) );
  INV_X1 U3982 ( .A(n3106), .ZN(n3108) );
  OAI211_X1 U3983 ( .C1(n3108), .C2(n3147), .A(n4314), .B(n3107), .ZN(n4614)
         );
  NOR2_X1 U3984 ( .A1(n4614), .A2(n3109), .ZN(n3116) );
  XNOR2_X1 U3985 ( .A(n3110), .B(n3874), .ZN(n3117) );
  XOR2_X1 U3986 ( .A(n3874), .B(n3111), .Z(n3114) );
  AOI22_X1 U3987 ( .A1(n3936), .A2(n4635), .B1(n3140), .B2(n4634), .ZN(n3112)
         );
  OAI21_X1 U3988 ( .B1(n3146), .B2(n4327), .A(n3112), .ZN(n3113) );
  AOI21_X1 U3989 ( .B1(n3114), .B2(n4189), .A(n3113), .ZN(n3115) );
  OAI21_X1 U3990 ( .B1(n3495), .B2(n3117), .A(n3115), .ZN(n4615) );
  AOI211_X1 U3991 ( .C1(n4557), .C2(n3126), .A(n3116), .B(n4615), .ZN(n3119)
         );
  INV_X1 U3992 ( .A(n3117), .ZN(n4618) );
  AOI22_X1 U3993 ( .A1(n4618), .A2(n4561), .B1(REG2_REG_4__SCAN_IN), .B2(n4566), .ZN(n3118) );
  OAI21_X1 U3994 ( .B1(n3119), .B2(n4566), .A(n3118), .ZN(U3286) );
  INV_X1 U3995 ( .A(n3120), .ZN(n3122) );
  NOR4_X1 U3996 ( .A1(n3124), .A2(n3123), .A3(n3122), .A4(n3121), .ZN(n3125)
         );
  INV_X1 U3997 ( .A(n2236), .ZN(n3369) );
  INV_X1 U3998 ( .A(n3126), .ZN(n3151) );
  OAI22_X1 U3999 ( .A1(n3146), .A2(n3624), .B1(n3621), .B2(n3156), .ZN(n3137)
         );
  NAND2_X1 U4000 ( .A1(n3938), .A2(n2253), .ZN(n3134) );
  NAND2_X1 U4001 ( .A1(n3132), .A2(n3131), .ZN(n3133) );
  NAND2_X1 U4002 ( .A1(n3134), .A2(n3133), .ZN(n3135) );
  XNOR2_X1 U4003 ( .A(n3135), .B(n3601), .ZN(n3136) );
  XOR2_X1 U4004 ( .A(n3137), .B(n3136), .Z(n3152) );
  INV_X1 U4005 ( .A(n3136), .ZN(n3139) );
  INV_X1 U4006 ( .A(n3137), .ZN(n3138) );
  OR2_X1 U4007 ( .A1(n3171), .A2(n3624), .ZN(n3142) );
  NAND2_X1 U4008 ( .A1(n3140), .A2(n2253), .ZN(n3141) );
  NAND2_X1 U4009 ( .A1(n3142), .A2(n3141), .ZN(n3160) );
  OAI22_X1 U4010 ( .A1(n3171), .A2(n3623), .B1(n3620), .B2(n3147), .ZN(n3143)
         );
  XNOR2_X1 U4011 ( .A(n3143), .B(n3601), .ZN(n3161) );
  XOR2_X1 U4012 ( .A(n3160), .B(n3161), .Z(n3144) );
  NAND2_X1 U4013 ( .A1(n3145), .A2(n3144), .ZN(n3162) );
  OAI211_X1 U4014 ( .C1(n3145), .C2(n3144), .A(n3162), .B(n4667), .ZN(n3150)
         );
  AND2_X1 U4015 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4443) );
  OAI22_X1 U4016 ( .A1(n2237), .A2(n3147), .B1(n3146), .B2(n3768), .ZN(n3148)
         );
  AOI211_X1 U4017 ( .C1(n4669), .C2(n3936), .A(n4443), .B(n3148), .ZN(n3149)
         );
  OAI211_X1 U4018 ( .C1(n3369), .C2(n3151), .A(n3150), .B(n3149), .ZN(U3227)
         );
  XNOR2_X1 U4019 ( .A(n3153), .B(n3152), .ZN(n3154) );
  NAND2_X1 U4020 ( .A1(n3154), .A2(n4667), .ZN(n3159) );
  NOR2_X1 U4021 ( .A1(STATE_REG_SCAN_IN), .A2(n3155), .ZN(n4388) );
  OAI22_X1 U4022 ( .A1(n2237), .A2(n3156), .B1(n2680), .B2(n3768), .ZN(n3157)
         );
  AOI211_X1 U4023 ( .C1(n4669), .C2(n3937), .A(n4388), .B(n3157), .ZN(n3158)
         );
  OAI211_X1 U4024 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3369), .A(n3159), .B(n3158), 
        .ZN(U3215) );
  INV_X1 U4025 ( .A(n3160), .ZN(n3164) );
  INV_X1 U4026 ( .A(n3161), .ZN(n3163) );
  OAI21_X1 U4027 ( .B1(n3164), .B2(n3163), .A(n3162), .ZN(n3169) );
  OAI22_X1 U4028 ( .A1(n3257), .A2(n3623), .B1(n3620), .B2(n3172), .ZN(n3165)
         );
  XNOR2_X1 U4029 ( .A(n3165), .B(n3601), .ZN(n3192) );
  AOI22_X1 U4030 ( .A1(n3936), .A2(n3166), .B1(n2253), .B2(n3167), .ZN(n3193)
         );
  XNOR2_X1 U4031 ( .A(n3192), .B(n3193), .ZN(n3168) );
  OAI211_X1 U4032 ( .C1(n3169), .C2(n3168), .A(n3196), .B(n4667), .ZN(n3175)
         );
  INV_X1 U4033 ( .A(REG3_REG_5__SCAN_IN), .ZN(n3170) );
  NOR2_X1 U4034 ( .A1(STATE_REG_SCAN_IN), .A2(n3170), .ZN(n4455) );
  OAI22_X1 U4035 ( .A1(n2237), .A2(n3172), .B1(n3171), .B2(n3768), .ZN(n3173)
         );
  AOI211_X1 U4036 ( .C1(n4669), .C2(n3935), .A(n4455), .B(n3173), .ZN(n3174)
         );
  OAI211_X1 U4037 ( .C1(n3369), .C2(n3176), .A(n3175), .B(n3174), .ZN(U3224)
         );
  INV_X1 U4038 ( .A(n3178), .ZN(n3856) );
  XNOR2_X1 U4039 ( .A(n3177), .B(n3856), .ZN(n4627) );
  INV_X1 U4040 ( .A(n4627), .ZN(n3191) );
  XNOR2_X1 U4041 ( .A(n3179), .B(n3178), .ZN(n3182) );
  OAI22_X1 U4042 ( .A1(n3313), .A2(n4594), .B1(n4593), .B2(n3247), .ZN(n3180)
         );
  AOI21_X1 U40430 ( .B1(n4637), .B2(n3935), .A(n3180), .ZN(n3181) );
  OAI21_X1 U4044 ( .B1(n3182), .B2(n4213), .A(n3181), .ZN(n4625) );
  NAND2_X1 U4045 ( .A1(n4625), .A2(n4402), .ZN(n3190) );
  INV_X1 U4046 ( .A(n3183), .ZN(n3185) );
  INV_X1 U4047 ( .A(n4314), .ZN(n4641) );
  INV_X1 U4048 ( .A(n3212), .ZN(n3184) );
  AOI211_X1 U4049 ( .C1(n3237), .C2(n3185), .A(n4641), .B(n3184), .ZN(n4626)
         );
  OAI22_X1 U4050 ( .A1(n4402), .A2(n3186), .B1(n3252), .B2(n4134), .ZN(n3187)
         );
  AOI21_X1 U4051 ( .B1(n4626), .B2(n3188), .A(n3187), .ZN(n3189) );
  OAI211_X1 U4052 ( .C1(n3191), .C2(n4223), .A(n3190), .B(n3189), .ZN(U3283)
         );
  NAND2_X1 U4053 ( .A1(n3192), .A2(n3194), .ZN(n3195) );
  NAND2_X1 U4054 ( .A1(n3935), .A2(n2253), .ZN(n3198) );
  NAND2_X1 U4055 ( .A1(n3264), .A2(n3131), .ZN(n3197) );
  NAND2_X1 U4056 ( .A1(n3198), .A2(n3197), .ZN(n3199) );
  XNOR2_X1 U4057 ( .A(n3199), .B(n3627), .ZN(n3201) );
  AOI22_X1 U4058 ( .A1(n3935), .A2(n3166), .B1(n2253), .B2(n3264), .ZN(n3200)
         );
  INV_X1 U4059 ( .A(n3243), .ZN(n3204) );
  NAND2_X1 U4060 ( .A1(n3201), .A2(n3200), .ZN(n3241) );
  NAND2_X1 U4061 ( .A1(n2292), .A2(n3241), .ZN(n3203) );
  AOI22_X1 U4062 ( .A1(n3204), .A2(n3241), .B1(n3202), .B2(n3203), .ZN(n3210)
         );
  OAI22_X1 U4063 ( .A1(n3525), .A2(n3760), .B1(STATE_REG_SCAN_IN), .B2(n3205), 
        .ZN(n3208) );
  OAI22_X1 U4064 ( .A1(n2237), .A2(n3206), .B1(n3257), .B2(n3768), .ZN(n3207)
         );
  AOI211_X1 U4065 ( .C1(n2236), .C2(n4558), .A(n3208), .B(n3207), .ZN(n3209)
         );
  OAI21_X1 U4066 ( .B1(n3210), .B2(n3775), .A(n3209), .ZN(U3236) );
  AND2_X1 U4067 ( .A1(n3798), .A2(n3795), .ZN(n3861) );
  XNOR2_X1 U4068 ( .A(n3211), .B(n3861), .ZN(n3287) );
  NAND2_X1 U4069 ( .A1(n3212), .A2(n3283), .ZN(n3213) );
  NAND2_X1 U4070 ( .A1(n3231), .A2(n3213), .ZN(n3291) );
  INV_X1 U4071 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3215) );
  INV_X1 U4072 ( .A(n3528), .ZN(n3214) );
  OAI22_X1 U4073 ( .A1(n4402), .A2(n3215), .B1(n3214), .B2(n4134), .ZN(n3216)
         );
  AOI21_X1 U4074 ( .B1(n3283), .B2(n4152), .A(n3216), .ZN(n3218) );
  AOI22_X1 U4075 ( .A1(n3255), .A2(n4066), .B1(n4151), .B2(n3934), .ZN(n3217)
         );
  OAI211_X1 U4076 ( .C1(n3291), .C2(n4220), .A(n3218), .B(n3217), .ZN(n3222)
         );
  XOR2_X1 U4077 ( .A(n3861), .B(n3219), .Z(n3220) );
  NAND2_X1 U4078 ( .A1(n3220), .A2(n4189), .ZN(n3285) );
  NOR2_X1 U4079 ( .A1(n3285), .A2(n4566), .ZN(n3221) );
  AOI211_X1 U4080 ( .C1(n3287), .C2(n4201), .A(n3222), .B(n3221), .ZN(n3223)
         );
  INV_X1 U4081 ( .A(n3223), .ZN(U3282) );
  AND2_X1 U4082 ( .A1(n2287), .A2(n3797), .ZN(n3858) );
  INV_X1 U4083 ( .A(n3858), .ZN(n3224) );
  XNOR2_X1 U4084 ( .A(n3225), .B(n3224), .ZN(n3226) );
  NAND2_X1 U4085 ( .A1(n3226), .A2(n4189), .ZN(n3229) );
  AOI22_X1 U4086 ( .A1(n4638), .A2(n4635), .B1(n4634), .B2(n3227), .ZN(n3228)
         );
  OAI211_X1 U4087 ( .C1(n3313), .C2(n4327), .A(n3229), .B(n3228), .ZN(n4630)
         );
  INV_X1 U4088 ( .A(n4630), .ZN(n3236) );
  XOR2_X1 U4089 ( .A(n3230), .B(n3858), .Z(n4632) );
  OAI21_X1 U4090 ( .B1(n2336), .B2(n3314), .A(n3274), .ZN(n4629) );
  NOR2_X1 U4091 ( .A1(n4629), .A2(n4220), .ZN(n3234) );
  INV_X1 U4092 ( .A(n3317), .ZN(n3232) );
  OAI22_X1 U4093 ( .A1(n4402), .A2(n2593), .B1(n3232), .B2(n4134), .ZN(n3233)
         );
  AOI211_X1 U4094 ( .C1(n4632), .C2(n4201), .A(n3234), .B(n3233), .ZN(n3235)
         );
  OAI21_X1 U4095 ( .B1(n4204), .B2(n3236), .A(n3235), .ZN(U3281) );
  AND2_X1 U4096 ( .A1(n3243), .A2(n3241), .ZN(n3245) );
  OR2_X1 U4097 ( .A1(n3525), .A2(n3624), .ZN(n3239) );
  NAND2_X1 U4098 ( .A1(n3237), .A2(n2253), .ZN(n3238) );
  NAND2_X1 U4099 ( .A1(n3239), .A2(n3238), .ZN(n3306) );
  OAI22_X1 U4100 ( .A1(n3525), .A2(n3623), .B1(n3620), .B2(n3247), .ZN(n3240)
         );
  XNOR2_X1 U4101 ( .A(n3240), .B(n3601), .ZN(n3305) );
  XOR2_X1 U4102 ( .A(n3306), .B(n3305), .Z(n3244) );
  NAND2_X1 U4103 ( .A1(n3243), .A2(n3242), .ZN(n3308) );
  OAI211_X1 U4104 ( .C1(n3245), .C2(n3244), .A(n3308), .B(n4667), .ZN(n3251)
         );
  INV_X1 U4105 ( .A(REG3_REG_7__SCAN_IN), .ZN(n5031) );
  NOR2_X1 U4106 ( .A1(STATE_REG_SCAN_IN), .A2(n5031), .ZN(n4469) );
  OAI22_X1 U4107 ( .A1(n2237), .A2(n3247), .B1(n3246), .B2(n3768), .ZN(n3248)
         );
  AOI211_X1 U4108 ( .C1(n4669), .C2(n3249), .A(n4469), .B(n3248), .ZN(n3250)
         );
  OAI211_X1 U4109 ( .C1(n3369), .C2(n3252), .A(n3251), .B(n3250), .ZN(U3210)
         );
  NAND2_X1 U4110 ( .A1(n3793), .A2(n3804), .ZN(n3876) );
  XOR2_X1 U4111 ( .A(n3876), .B(n3253), .Z(n3258) );
  INV_X1 U4112 ( .A(n3258), .ZN(n4562) );
  XOR2_X1 U4113 ( .A(n3876), .B(n3254), .Z(n3261) );
  AOI22_X1 U4114 ( .A1(n3255), .A2(n4635), .B1(n4634), .B2(n3264), .ZN(n3256)
         );
  OAI21_X1 U4115 ( .B1(n3257), .B2(n4327), .A(n3256), .ZN(n3260) );
  NOR2_X1 U4116 ( .A1(n3258), .A2(n3495), .ZN(n3259) );
  AOI211_X1 U4117 ( .C1(n3261), .C2(n4189), .A(n3260), .B(n3259), .ZN(n4565)
         );
  INV_X1 U4118 ( .A(n4565), .ZN(n3262) );
  AOI21_X1 U4119 ( .B1(n4617), .B2(n4562), .A(n3262), .ZN(n3269) );
  AOI21_X1 U4120 ( .B1(n3264), .B2(n3263), .A(n3183), .ZN(n4559) );
  INV_X1 U4121 ( .A(n4378), .ZN(n4336) );
  INV_X1 U4122 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3265) );
  NOR2_X1 U4123 ( .A1(n4649), .A2(n3265), .ZN(n3266) );
  AOI21_X1 U4124 ( .B1(n4559), .B2(n4336), .A(n3266), .ZN(n3267) );
  OAI21_X1 U4125 ( .B1(n3269), .B2(n4647), .A(n3267), .ZN(U3479) );
  INV_X1 U4126 ( .A(n4333), .ZN(n4235) );
  AOI22_X1 U4127 ( .A1(n4559), .A2(n4235), .B1(n4663), .B2(REG1_REG_6__SCAN_IN), .ZN(n3268) );
  OAI21_X1 U4128 ( .B1(n3269), .B2(n4663), .A(n3268), .ZN(U3524) );
  NAND2_X1 U4129 ( .A1(n3812), .A2(n3813), .ZN(n3877) );
  INV_X1 U4130 ( .A(n3877), .ZN(n3272) );
  XNOR2_X1 U4131 ( .A(n3270), .B(n3272), .ZN(n3271) );
  NAND2_X1 U4132 ( .A1(n3271), .A2(n4189), .ZN(n3326) );
  XNOR2_X1 U4133 ( .A(n3273), .B(n3272), .ZN(n3321) );
  NAND2_X1 U4134 ( .A1(n3321), .A2(n4201), .ZN(n3282) );
  AOI21_X1 U4135 ( .B1(n3356), .B2(n3274), .A(n3295), .ZN(n3333) );
  AOI22_X1 U4136 ( .A1(n3428), .A2(n4151), .B1(n4066), .B2(n3934), .ZN(n3279)
         );
  INV_X1 U4137 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3276) );
  INV_X1 U4138 ( .A(n3275), .ZN(n3368) );
  OAI22_X1 U4139 ( .A1(n4402), .A2(n3276), .B1(n3368), .B2(n4134), .ZN(n3277)
         );
  AOI21_X1 U4140 ( .B1(n3356), .B2(n4152), .A(n3277), .ZN(n3278) );
  NAND2_X1 U4141 ( .A1(n3279), .A2(n3278), .ZN(n3280) );
  AOI21_X1 U4142 ( .B1(n3333), .B2(n4560), .A(n3280), .ZN(n3281) );
  OAI211_X1 U4143 ( .C1(n4566), .C2(n3326), .A(n3282), .B(n3281), .ZN(U3280)
         );
  INV_X1 U4144 ( .A(REG0_REG_8__SCAN_IN), .ZN(n5009) );
  AOI22_X1 U4145 ( .A1(n3934), .A2(n4635), .B1(n4634), .B2(n3283), .ZN(n3284)
         );
  OAI211_X1 U4146 ( .C1(n3525), .C2(n4327), .A(n3285), .B(n3284), .ZN(n3286)
         );
  AOI21_X1 U4147 ( .B1(n3287), .B2(n4646), .A(n3286), .ZN(n3289) );
  MUX2_X1 U4148 ( .A(n5009), .B(n3289), .S(n4649), .Z(n3288) );
  OAI21_X1 U4149 ( .B1(n3291), .B2(n4378), .A(n3288), .ZN(U3483) );
  MUX2_X1 U4150 ( .A(n4479), .B(n3289), .S(n4666), .Z(n3290) );
  OAI21_X1 U4151 ( .B1(n3291), .B2(n4333), .A(n3290), .ZN(U3526) );
  XNOR2_X1 U4152 ( .A(n3292), .B(n3855), .ZN(n4645) );
  INV_X1 U4153 ( .A(n4645), .ZN(n3303) );
  XNOR2_X1 U4154 ( .A(n3293), .B(n3855), .ZN(n3294) );
  NOR2_X1 U4155 ( .A1(n3294), .A2(n4213), .ZN(n4643) );
  OR2_X1 U4156 ( .A1(n3295), .A2(n3384), .ZN(n3296) );
  NAND2_X1 U4157 ( .A1(n3336), .A2(n3296), .ZN(n4642) );
  OAI22_X1 U4158 ( .A1(n4402), .A2(n2609), .B1(n3297), .B2(n4134), .ZN(n3298)
         );
  AOI21_X1 U4159 ( .B1(n4633), .B2(n4152), .A(n3298), .ZN(n3300) );
  AOI22_X1 U4160 ( .A1(n4066), .A2(n4638), .B1(n4151), .B2(n4636), .ZN(n3299)
         );
  OAI211_X1 U4161 ( .C1(n4642), .C2(n4220), .A(n3300), .B(n3299), .ZN(n3301)
         );
  AOI21_X1 U4162 ( .B1(n4643), .B2(n4402), .A(n3301), .ZN(n3302) );
  OAI21_X1 U4163 ( .B1(n3303), .B2(n4223), .A(n3302), .ZN(U3279) );
  OAI22_X1 U4164 ( .A1(n3363), .A2(n3623), .B1(n3620), .B2(n3314), .ZN(n3304)
         );
  XNOR2_X1 U4165 ( .A(n3304), .B(n3601), .ZN(n3349) );
  OAI22_X1 U4166 ( .A1(n3363), .A2(n3624), .B1(n3623), .B2(n3314), .ZN(n3350)
         );
  XNOR2_X1 U4167 ( .A(n3349), .B(n3350), .ZN(n3312) );
  OAI22_X1 U4168 ( .A1(n3313), .A2(n3624), .B1(n3623), .B2(n3526), .ZN(n3520)
         );
  OAI22_X1 U4169 ( .A1(n3313), .A2(n3623), .B1(n3620), .B2(n3526), .ZN(n3309)
         );
  XNOR2_X1 U4170 ( .A(n3309), .B(n3601), .ZN(n3522) );
  INV_X1 U4171 ( .A(n3359), .ZN(n3310) );
  AOI21_X1 U4172 ( .B1(n3312), .B2(n3311), .A(n3310), .ZN(n3320) );
  OAI22_X1 U4173 ( .A1(n2237), .A2(n3314), .B1(n3313), .B2(n3768), .ZN(n3315)
         );
  AOI211_X1 U4174 ( .C1(n4669), .C2(n4638), .A(n3316), .B(n3315), .ZN(n3319)
         );
  NAND2_X1 U4175 ( .A1(n2236), .A2(n3317), .ZN(n3318) );
  OAI211_X1 U4176 ( .C1(n3320), .C2(n3775), .A(n3319), .B(n3318), .ZN(U3228)
         );
  NAND2_X1 U4177 ( .A1(n3321), .A2(n4646), .ZN(n3328) );
  NAND2_X1 U4178 ( .A1(n3356), .A2(n4634), .ZN(n3323) );
  NAND2_X1 U4179 ( .A1(n3934), .A2(n4637), .ZN(n3322) );
  OAI211_X1 U4180 ( .C1(n3393), .C2(n4594), .A(n3323), .B(n3322), .ZN(n3324)
         );
  INV_X1 U4181 ( .A(n3324), .ZN(n3325) );
  AND2_X1 U4182 ( .A1(n3326), .A2(n3325), .ZN(n3327) );
  NAND2_X1 U4183 ( .A1(n3328), .A2(n3327), .ZN(n3331) );
  MUX2_X1 U4184 ( .A(REG0_REG_10__SCAN_IN), .B(n3331), .S(n4649), .Z(n3329) );
  AOI21_X1 U4185 ( .B1(n3333), .B2(n4336), .A(n3329), .ZN(n3330) );
  INV_X1 U4186 ( .A(n3330), .ZN(U3487) );
  MUX2_X1 U4187 ( .A(REG1_REG_10__SCAN_IN), .B(n3331), .S(n4666), .Z(n3332) );
  AOI21_X1 U4188 ( .B1(n3333), .B2(n4235), .A(n3332), .ZN(n3334) );
  INV_X1 U4189 ( .A(n3334), .ZN(U3528) );
  AND2_X1 U4190 ( .A1(n3405), .A2(n3406), .ZN(n3862) );
  XOR2_X1 U4191 ( .A(n3862), .B(n3335), .Z(n3395) );
  NAND2_X1 U4192 ( .A1(n3336), .A2(n3429), .ZN(n3337) );
  NAND2_X1 U4193 ( .A1(n3415), .A2(n3337), .ZN(n3400) );
  INV_X1 U4194 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3339) );
  INV_X1 U4195 ( .A(n3432), .ZN(n3338) );
  OAI22_X1 U4196 ( .A1(n4402), .A2(n3339), .B1(n3338), .B2(n4134), .ZN(n3340)
         );
  AOI21_X1 U4197 ( .B1(n3429), .B2(n4152), .A(n3340), .ZN(n3342) );
  AOI22_X1 U4198 ( .A1(n4066), .A2(n3428), .B1(n3514), .B2(n4151), .ZN(n3341)
         );
  OAI211_X1 U4199 ( .C1(n3400), .C2(n4220), .A(n3342), .B(n3341), .ZN(n3347)
         );
  NAND2_X1 U4200 ( .A1(n3344), .A2(n3343), .ZN(n3408) );
  XNOR2_X1 U4201 ( .A(n3408), .B(n3862), .ZN(n3345) );
  NAND2_X1 U4202 ( .A1(n3345), .A2(n4189), .ZN(n3392) );
  NOR2_X1 U4203 ( .A1(n3392), .A2(n4566), .ZN(n3346) );
  AOI211_X1 U4204 ( .C1(n4201), .C2(n3395), .A(n3347), .B(n3346), .ZN(n3348)
         );
  INV_X1 U4205 ( .A(n3348), .ZN(U3278) );
  INV_X1 U4206 ( .A(n3349), .ZN(n3352) );
  INV_X1 U4207 ( .A(n3350), .ZN(n3351) );
  NAND2_X1 U4208 ( .A1(n3352), .A2(n3351), .ZN(n3357) );
  AND2_X1 U4209 ( .A1(n3359), .A2(n3357), .ZN(n3361) );
  NAND2_X1 U4210 ( .A1(n4638), .A2(n2253), .ZN(n3354) );
  NAND2_X1 U4211 ( .A1(n3356), .A2(n3131), .ZN(n3353) );
  NAND2_X1 U4212 ( .A1(n3354), .A2(n3353), .ZN(n3355) );
  XNOR2_X1 U4213 ( .A(n3355), .B(n3601), .ZN(n3377) );
  AOI22_X1 U4214 ( .A1(n4638), .A2(n3166), .B1(n2253), .B2(n3356), .ZN(n3378)
         );
  XNOR2_X1 U4215 ( .A(n3377), .B(n3378), .ZN(n3360) );
  OAI211_X1 U4216 ( .C1(n3361), .C2(n3360), .A(n4667), .B(n3381), .ZN(n3367)
         );
  NOR2_X1 U4217 ( .A1(STATE_REG_SCAN_IN), .A2(n3362), .ZN(n4489) );
  OAI22_X1 U4218 ( .A1(n2237), .A2(n3364), .B1(n3363), .B2(n3768), .ZN(n3365)
         );
  AOI211_X1 U4219 ( .C1(n4669), .C2(n3428), .A(n4489), .B(n3365), .ZN(n3366)
         );
  OAI211_X1 U4220 ( .C1(n3369), .C2(n3368), .A(n3367), .B(n3366), .ZN(U3214)
         );
  OAI22_X1 U4221 ( .A1(n3393), .A2(n3623), .B1(n3620), .B2(n3384), .ZN(n3370)
         );
  XNOR2_X1 U4222 ( .A(n3370), .B(n3627), .ZN(n3376) );
  INV_X1 U4223 ( .A(n3376), .ZN(n3374) );
  OR2_X1 U4224 ( .A1(n3393), .A2(n3624), .ZN(n3372) );
  NAND2_X1 U4225 ( .A1(n4633), .A2(n2253), .ZN(n3371) );
  INV_X1 U4226 ( .A(n3375), .ZN(n3373) );
  NAND2_X1 U4227 ( .A1(n3374), .A2(n3373), .ZN(n3423) );
  NAND2_X1 U4228 ( .A1(n3376), .A2(n3375), .ZN(n3421) );
  NAND2_X1 U4229 ( .A1(n3423), .A2(n3421), .ZN(n3382) );
  INV_X1 U4230 ( .A(n3377), .ZN(n3379) );
  OR2_X1 U4231 ( .A1(n3379), .A2(n3378), .ZN(n3380) );
  NAND2_X1 U4232 ( .A1(n3381), .A2(n3380), .ZN(n3422) );
  XOR2_X1 U4233 ( .A(n3382), .B(n3422), .Z(n3389) );
  INV_X1 U4234 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4934) );
  NOR2_X1 U4235 ( .A1(STATE_REG_SCAN_IN), .A2(n4934), .ZN(n4498) );
  OAI22_X1 U4236 ( .A1(n2237), .A2(n3384), .B1(n3383), .B2(n3768), .ZN(n3385)
         );
  AOI211_X1 U4237 ( .C1(n4669), .C2(n4636), .A(n4498), .B(n3385), .ZN(n3388)
         );
  NAND2_X1 U4238 ( .A1(n2236), .A2(n3386), .ZN(n3387) );
  OAI211_X1 U4239 ( .C1(n3389), .C2(n3775), .A(n3388), .B(n3387), .ZN(U3233)
         );
  INV_X1 U4240 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3396) );
  OAI22_X1 U4241 ( .A1(n4328), .A2(n4594), .B1(n4593), .B2(n3425), .ZN(n3390)
         );
  INV_X1 U4242 ( .A(n3390), .ZN(n3391) );
  OAI211_X1 U4243 ( .C1(n3393), .C2(n4327), .A(n3392), .B(n3391), .ZN(n3394)
         );
  AOI21_X1 U4244 ( .B1(n3395), .B2(n4646), .A(n3394), .ZN(n3398) );
  MUX2_X1 U4245 ( .A(n3396), .B(n3398), .S(n4649), .Z(n3397) );
  OAI21_X1 U4246 ( .B1(n3400), .B2(n4378), .A(n3397), .ZN(U3491) );
  MUX2_X1 U4247 ( .A(n4507), .B(n3398), .S(n4666), .Z(n3399) );
  OAI21_X1 U4248 ( .B1(n3400), .B2(n4333), .A(n3399), .ZN(U3530) );
  INV_X1 U4249 ( .A(n3401), .ZN(n3403) );
  OR2_X1 U4250 ( .A1(n3403), .A2(n3402), .ZN(n3859) );
  XNOR2_X1 U4251 ( .A(n3404), .B(n3859), .ZN(n3414) );
  INV_X1 U4252 ( .A(n3405), .ZN(n3407) );
  OAI21_X1 U4253 ( .B1(n3408), .B2(n3407), .A(n3406), .ZN(n3409) );
  XNOR2_X1 U4254 ( .A(n3409), .B(n3859), .ZN(n3412) );
  AOI22_X1 U4255 ( .A1(n3933), .A2(n4635), .B1(n3457), .B2(n4634), .ZN(n3410)
         );
  OAI21_X1 U4256 ( .B1(n3426), .B2(n4327), .A(n3410), .ZN(n3411) );
  AOI21_X1 U4257 ( .B1(n3412), .B2(n4189), .A(n3411), .ZN(n3413) );
  OAI21_X1 U4258 ( .B1(n3414), .B2(n3495), .A(n3413), .ZN(n3435) );
  INV_X1 U4259 ( .A(n3435), .ZN(n3420) );
  INV_X1 U4260 ( .A(n3414), .ZN(n3436) );
  AND2_X1 U4261 ( .A1(n3415), .A2(n3457), .ZN(n3416) );
  OR2_X1 U4262 ( .A1(n3416), .A2(n3498), .ZN(n3442) );
  AOI22_X1 U4263 ( .A1(n4566), .A2(REG2_REG_13__SCAN_IN), .B1(n3460), .B2(
        n4557), .ZN(n3417) );
  OAI21_X1 U4264 ( .B1(n3442), .B2(n4220), .A(n3417), .ZN(n3418) );
  AOI21_X1 U4265 ( .B1(n3436), .B2(n4561), .A(n3418), .ZN(n3419) );
  OAI21_X1 U4266 ( .B1(n3420), .B2(n4566), .A(n3419), .ZN(U3277) );
  OAI22_X1 U4267 ( .A1(n3426), .A2(n3621), .B1(n3620), .B2(n3425), .ZN(n3424)
         );
  XNOR2_X1 U4268 ( .A(n3424), .B(n3601), .ZN(n3444) );
  INV_X1 U4269 ( .A(n3444), .ZN(n3445) );
  OAI22_X1 U4270 ( .A1(n3426), .A2(n3624), .B1(n3623), .B2(n3425), .ZN(n3443)
         );
  XNOR2_X1 U4271 ( .A(n3445), .B(n3443), .ZN(n3427) );
  XNOR2_X1 U4272 ( .A(n3446), .B(n3427), .ZN(n3434) );
  INV_X1 U4273 ( .A(n3768), .ZN(n3746) );
  AOI22_X1 U4274 ( .A1(n4671), .A2(n3429), .B1(n3428), .B2(n3746), .ZN(n3430)
         );
  NAND2_X1 U4275 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4508) );
  OAI211_X1 U4276 ( .C1(n4328), .C2(n3760), .A(n3430), .B(n4508), .ZN(n3431)
         );
  AOI21_X1 U4277 ( .B1(n2236), .B2(n3432), .A(n3431), .ZN(n3433) );
  OAI21_X1 U4278 ( .B1(n3434), .B2(n3775), .A(n3433), .ZN(U3221) );
  AOI21_X1 U4279 ( .B1(n4617), .B2(n3436), .A(n3435), .ZN(n3439) );
  MUX2_X1 U4280 ( .A(n3437), .B(n3439), .S(n4666), .Z(n3438) );
  OAI21_X1 U4281 ( .B1(n4333), .B2(n3442), .A(n3438), .ZN(U3531) );
  INV_X1 U4282 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3440) );
  MUX2_X1 U4283 ( .A(n3440), .B(n3439), .S(n4649), .Z(n3441) );
  OAI21_X1 U4284 ( .B1(n3442), .B2(n4378), .A(n3441), .ZN(U3493) );
  OAI22_X1 U4285 ( .A1(n4328), .A2(n3621), .B1(n3620), .B2(n3447), .ZN(n3448)
         );
  XNOR2_X1 U4286 ( .A(n3448), .B(n3601), .ZN(n3454) );
  INV_X1 U4287 ( .A(n3454), .ZN(n3452) );
  OR2_X1 U4288 ( .A1(n4328), .A2(n3624), .ZN(n3450) );
  NAND2_X1 U4289 ( .A1(n3457), .A2(n2253), .ZN(n3449) );
  NAND2_X1 U4290 ( .A1(n3450), .A2(n3449), .ZN(n3453) );
  INV_X1 U4291 ( .A(n3453), .ZN(n3451) );
  NAND2_X1 U4292 ( .A1(n3452), .A2(n3451), .ZN(n3506) );
  INV_X1 U4293 ( .A(n3506), .ZN(n3455) );
  NOR2_X1 U4294 ( .A1(n3455), .A2(n3507), .ZN(n3456) );
  XNOR2_X1 U4295 ( .A(n3508), .B(n3456), .ZN(n3462) );
  AOI22_X1 U4296 ( .A1(n4671), .A2(n3457), .B1(n3746), .B2(n4636), .ZN(n3458)
         );
  NAND2_X1 U4297 ( .A1(REG3_REG_13__SCAN_IN), .A2(U3149), .ZN(n4525) );
  OAI211_X1 U4298 ( .C1(n3769), .C2(n3760), .A(n3458), .B(n4525), .ZN(n3459)
         );
  AOI21_X1 U4299 ( .B1(n2236), .B2(n3460), .A(n3459), .ZN(n3461) );
  OAI21_X1 U4300 ( .B1(n3462), .B2(n3775), .A(n3461), .ZN(U3231) );
  INV_X1 U4301 ( .A(n3463), .ZN(n3489) );
  NOR2_X1 U4302 ( .A1(n3489), .A2(n3490), .ZN(n3488) );
  NOR2_X1 U4303 ( .A1(n3488), .A2(n3464), .ZN(n3465) );
  XOR2_X1 U4304 ( .A(n3881), .B(n3465), .Z(n4320) );
  INV_X1 U4305 ( .A(n4320), .ZN(n3474) );
  NAND2_X1 U4306 ( .A1(n3492), .A2(n3820), .ZN(n3466) );
  XNOR2_X1 U4307 ( .A(n3466), .B(n3881), .ZN(n3469) );
  OAI22_X1 U4308 ( .A1(n3710), .A2(n4594), .B1(n3770), .B2(n4593), .ZN(n3467)
         );
  AOI21_X1 U4309 ( .B1(n4637), .B2(n3933), .A(n3467), .ZN(n3468) );
  OAI21_X1 U4310 ( .B1(n3469), .B2(n4213), .A(n3468), .ZN(n4319) );
  OR2_X1 U4311 ( .A1(n3496), .A2(n3770), .ZN(n3470) );
  NAND2_X1 U4312 ( .A1(n3483), .A2(n3470), .ZN(n4375) );
  AOI22_X1 U4313 ( .A1(n4566), .A2(REG2_REG_15__SCAN_IN), .B1(n3772), .B2(
        n4557), .ZN(n3471) );
  OAI21_X1 U4314 ( .B1(n4375), .B2(n4220), .A(n3471), .ZN(n3472) );
  AOI21_X1 U4315 ( .B1(n4319), .B2(n4402), .A(n3472), .ZN(n3473) );
  OAI21_X1 U4316 ( .B1(n3474), .B2(n4223), .A(n3473), .ZN(U3275) );
  XNOR2_X1 U4317 ( .A(n3475), .B(n2423), .ZN(n3478) );
  AOI22_X1 U4318 ( .A1(n3745), .A2(n4635), .B1(n4634), .B2(n3482), .ZN(n3476)
         );
  OAI21_X1 U4319 ( .B1(n3699), .B2(n4327), .A(n3476), .ZN(n3477) );
  AOI21_X1 U4320 ( .B1(n3478), .B2(n4189), .A(n3477), .ZN(n4317) );
  AOI21_X1 U4321 ( .B1(n3481), .B2(n3479), .A(n3480), .ZN(n4312) );
  NAND2_X1 U4322 ( .A1(n3483), .A2(n3482), .ZN(n4313) );
  AND3_X1 U4323 ( .A1(n4315), .A2(n4560), .A3(n4313), .ZN(n3486) );
  INV_X1 U4324 ( .A(n3702), .ZN(n3484) );
  OAI22_X1 U4325 ( .A1(n4402), .A2(n3967), .B1(n3484), .B2(n4134), .ZN(n3485)
         );
  AOI211_X1 U4326 ( .C1(n4312), .C2(n4201), .A(n3486), .B(n3485), .ZN(n3487)
         );
  OAI21_X1 U4327 ( .B1(n4204), .B2(n4317), .A(n3487), .ZN(U3274) );
  AOI21_X1 U4328 ( .B1(n3490), .B2(n3489), .A(n3488), .ZN(n4323) );
  INV_X1 U4329 ( .A(n3491), .ZN(n3891) );
  INV_X1 U4330 ( .A(n3492), .ZN(n3493) );
  AOI21_X1 U4331 ( .B1(n3891), .B2(n3878), .A(n3493), .ZN(n3494) );
  OAI22_X1 U4332 ( .A1(n4323), .A2(n3495), .B1(n4213), .B2(n3494), .ZN(n4329)
         );
  NAND2_X1 U4333 ( .A1(n4329), .A2(n4402), .ZN(n3504) );
  INV_X1 U4334 ( .A(n3496), .ZN(n3497) );
  OAI21_X1 U4335 ( .B1(n3498), .B2(n3509), .A(n3497), .ZN(n4379) );
  INV_X1 U4336 ( .A(n4379), .ZN(n3502) );
  AOI22_X1 U4337 ( .A1(n3514), .A2(n4066), .B1(n4151), .B2(n4325), .ZN(n3500)
         );
  AOI22_X1 U4338 ( .A1(n4566), .A2(REG2_REG_14__SCAN_IN), .B1(n3517), .B2(
        n4557), .ZN(n3499) );
  OAI211_X1 U4339 ( .C1(n3509), .C2(n4071), .A(n3500), .B(n3499), .ZN(n3501)
         );
  AOI21_X1 U4340 ( .B1(n3502), .B2(n4560), .A(n3501), .ZN(n3503) );
  OAI211_X1 U4341 ( .C1(n4323), .C2(n3505), .A(n3504), .B(n3503), .ZN(U3276)
         );
  OAI22_X1 U4342 ( .A1(n3769), .A2(n3623), .B1(n3620), .B2(n3509), .ZN(n3510)
         );
  XNOR2_X1 U4343 ( .A(n3510), .B(n3627), .ZN(n3537) );
  OR2_X1 U4344 ( .A1(n3769), .A2(n3624), .ZN(n3512) );
  NAND2_X1 U4345 ( .A1(n4324), .A2(n2253), .ZN(n3511) );
  XNOR2_X1 U4346 ( .A(n3537), .B(n3536), .ZN(n3513) );
  XNOR2_X1 U4347 ( .A(n3535), .B(n3513), .ZN(n3519) );
  AOI22_X1 U4348 ( .A1(n4671), .A2(n4324), .B1(n3514), .B2(n3746), .ZN(n3515)
         );
  NAND2_X1 U4349 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4539) );
  OAI211_X1 U4350 ( .C1(n3699), .C2(n3760), .A(n3515), .B(n4539), .ZN(n3516)
         );
  AOI21_X1 U4351 ( .B1(n2236), .B2(n3517), .A(n3516), .ZN(n3518) );
  OAI21_X1 U4352 ( .B1(n3519), .B2(n3775), .A(n3518), .ZN(U3212) );
  INV_X1 U4353 ( .A(n3520), .ZN(n3521) );
  XNOR2_X1 U4354 ( .A(n3522), .B(n3521), .ZN(n3523) );
  XNOR2_X1 U4355 ( .A(n3524), .B(n3523), .ZN(n3531) );
  INV_X1 U4356 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4837) );
  NOR2_X1 U4357 ( .A1(STATE_REG_SCAN_IN), .A2(n4837), .ZN(n4481) );
  OAI22_X1 U4358 ( .A1(n2237), .A2(n3526), .B1(n3525), .B2(n3768), .ZN(n3527)
         );
  AOI211_X1 U4359 ( .C1(n4669), .C2(n3934), .A(n4481), .B(n3527), .ZN(n3530)
         );
  NAND2_X1 U4360 ( .A1(n2236), .A2(n3528), .ZN(n3529) );
  OAI211_X1 U4361 ( .C1(n3531), .C2(n3775), .A(n3530), .B(n3529), .ZN(U3218)
         );
  NAND2_X1 U4362 ( .A1(n3537), .A2(n3536), .ZN(n3538) );
  NAND2_X1 U4363 ( .A1(n3539), .A2(n3538), .ZN(n3544) );
  OAI22_X1 U4364 ( .A1(n3699), .A2(n3621), .B1(n3620), .B2(n3770), .ZN(n3540)
         );
  XOR2_X1 U4365 ( .A(n3601), .B(n3540), .Z(n3545) );
  NAND2_X1 U4366 ( .A1(n3544), .A2(n3545), .ZN(n3694) );
  NAND2_X1 U4367 ( .A1(n4325), .A2(n3166), .ZN(n3543) );
  NAND2_X1 U4368 ( .A1(n3541), .A2(n2253), .ZN(n3542) );
  NAND2_X1 U4369 ( .A1(n3543), .A2(n3542), .ZN(n3767) );
  NAND2_X1 U4370 ( .A1(n3694), .A2(n3767), .ZN(n3549) );
  INV_X1 U4371 ( .A(n3544), .ZN(n3547) );
  INV_X1 U4372 ( .A(n3545), .ZN(n3546) );
  OAI22_X1 U4373 ( .A1(n3710), .A2(n3624), .B1(n3621), .B2(n3700), .ZN(n3550)
         );
  OAI22_X1 U4374 ( .A1(n3710), .A2(n3623), .B1(n3620), .B2(n3700), .ZN(n3548)
         );
  XNOR2_X1 U4375 ( .A(n3548), .B(n3601), .ZN(n3551) );
  XOR2_X1 U4376 ( .A(n3550), .B(n3551), .Z(n3697) );
  NAND3_X1 U4377 ( .A1(n3549), .A2(n3765), .A3(n3697), .ZN(n3553) );
  NAND2_X1 U4378 ( .A1(n3553), .A2(n3552), .ZN(n3706) );
  NAND2_X1 U4379 ( .A1(n3745), .A2(n2253), .ZN(n3555) );
  NAND2_X1 U4380 ( .A1(n4215), .A2(n3131), .ZN(n3554) );
  NAND2_X1 U4381 ( .A1(n3555), .A2(n3554), .ZN(n3556) );
  XNOR2_X1 U4382 ( .A(n3556), .B(n3627), .ZN(n3558) );
  AOI22_X1 U4383 ( .A1(n3745), .A2(n3166), .B1(n2253), .B2(n4215), .ZN(n3557)
         );
  OR2_X1 U4384 ( .A1(n3558), .A2(n3557), .ZN(n3708) );
  NAND2_X1 U4385 ( .A1(n3706), .A2(n3708), .ZN(n3559) );
  NAND2_X1 U4386 ( .A1(n3558), .A2(n3557), .ZN(n3707) );
  NAND2_X1 U4387 ( .A1(n3559), .A2(n3707), .ZN(n3741) );
  AOI22_X1 U4388 ( .A1(n4172), .A2(n3166), .B1(n2253), .B2(n4184), .ZN(n3742)
         );
  OAI22_X1 U4389 ( .A1(n4209), .A2(n3621), .B1(n3620), .B2(n4194), .ZN(n3560)
         );
  XOR2_X1 U4390 ( .A(n3601), .B(n3560), .Z(n3743) );
  OAI22_X1 U4391 ( .A1(n4296), .A2(n3621), .B1(n3620), .B2(n4176), .ZN(n3561)
         );
  XNOR2_X1 U4392 ( .A(n3561), .B(n3627), .ZN(n3566) );
  OR2_X1 U4393 ( .A1(n4296), .A2(n3624), .ZN(n3564) );
  NAND2_X1 U4394 ( .A1(n3562), .A2(n2253), .ZN(n3563) );
  NAND2_X1 U4395 ( .A1(n3566), .A2(n3565), .ZN(n3568) );
  OAI21_X1 U4396 ( .B1(n3566), .B2(n3565), .A(n3568), .ZN(n3668) );
  NAND2_X1 U4397 ( .A1(n4121), .A2(n2253), .ZN(n3570) );
  NAND2_X1 U4398 ( .A1(n4292), .A2(n3131), .ZN(n3569) );
  NAND2_X1 U4399 ( .A1(n3570), .A2(n3569), .ZN(n3571) );
  XNOR2_X1 U4400 ( .A(n3571), .B(n3601), .ZN(n3574) );
  NAND2_X1 U4401 ( .A1(n4121), .A2(n3166), .ZN(n3573) );
  NAND2_X1 U4402 ( .A1(n4292), .A2(n2253), .ZN(n3572) );
  NAND2_X1 U4403 ( .A1(n3573), .A2(n3572), .ZN(n3575) );
  NAND2_X1 U4404 ( .A1(n3574), .A2(n3575), .ZN(n3724) );
  INV_X1 U4405 ( .A(n3574), .ZN(n3577) );
  INV_X1 U4406 ( .A(n3575), .ZN(n3576) );
  NAND2_X1 U4407 ( .A1(n3577), .A2(n3576), .ZN(n3726) );
  NAND2_X1 U4408 ( .A1(n4293), .A2(n2253), .ZN(n3579) );
  NAND2_X1 U4409 ( .A1(n4128), .A2(n3131), .ZN(n3578) );
  NAND2_X1 U4410 ( .A1(n3579), .A2(n3578), .ZN(n3580) );
  XNOR2_X1 U4411 ( .A(n3580), .B(n3627), .ZN(n3582) );
  NOR2_X1 U4412 ( .A1(n4132), .A2(n3623), .ZN(n3581) );
  AOI21_X1 U4413 ( .B1(n4293), .B2(n3166), .A(n3581), .ZN(n3583) );
  AND2_X1 U4414 ( .A1(n3582), .A2(n3583), .ZN(n3673) );
  INV_X1 U4415 ( .A(n3582), .ZN(n3585) );
  INV_X1 U4416 ( .A(n3583), .ZN(n3584) );
  NAND2_X1 U4417 ( .A1(n3585), .A2(n3584), .ZN(n3674) );
  OAI22_X1 U4418 ( .A1(n3660), .A2(n3621), .B1(n3620), .B2(n4112), .ZN(n3586)
         );
  XNOR2_X1 U4419 ( .A(n3586), .B(n3601), .ZN(n3587) );
  OAI22_X1 U4420 ( .A1(n3660), .A2(n3624), .B1(n3621), .B2(n4112), .ZN(n3588)
         );
  XNOR2_X1 U4421 ( .A(n3587), .B(n3588), .ZN(n3735) );
  INV_X1 U4422 ( .A(n3587), .ZN(n3590) );
  INV_X1 U4423 ( .A(n3588), .ZN(n3589) );
  NAND2_X1 U4424 ( .A1(n3590), .A2(n3589), .ZN(n3658) );
  OAI22_X1 U4425 ( .A1(n4276), .A2(n3621), .B1(n3620), .B2(n4092), .ZN(n3591)
         );
  XNOR2_X1 U4426 ( .A(n3591), .B(n3627), .ZN(n3596) );
  OR2_X1 U4427 ( .A1(n4276), .A2(n3624), .ZN(n3594) );
  NAND2_X1 U4428 ( .A1(n3592), .A2(n2253), .ZN(n3593) );
  NAND2_X1 U4429 ( .A1(n3594), .A2(n3593), .ZN(n3597) );
  XNOR2_X1 U4430 ( .A(n3596), .B(n3597), .ZN(n3657) );
  INV_X1 U4431 ( .A(n3596), .ZN(n3598) );
  NAND2_X1 U4432 ( .A1(n3598), .A2(n3597), .ZN(n3603) );
  NOR2_X1 U4433 ( .A1(n4072), .A2(n3623), .ZN(n3599) );
  AOI21_X1 U4434 ( .B1(n4264), .B2(n3166), .A(n3599), .ZN(n3604) );
  OAI22_X1 U4435 ( .A1(n4087), .A2(n3621), .B1(n3620), .B2(n4072), .ZN(n3602)
         );
  XNOR2_X1 U4436 ( .A(n3602), .B(n3601), .ZN(n3716) );
  INV_X1 U4437 ( .A(n3604), .ZN(n3605) );
  NAND2_X1 U4438 ( .A1(n4273), .A2(n2253), .ZN(n3607) );
  NAND2_X1 U4439 ( .A1(n4263), .A2(n3131), .ZN(n3606) );
  NAND2_X1 U4440 ( .A1(n3607), .A2(n3606), .ZN(n3608) );
  XNOR2_X1 U4441 ( .A(n3608), .B(n3627), .ZN(n3611) );
  NOR2_X1 U4442 ( .A1(n4052), .A2(n3623), .ZN(n3609) );
  AOI21_X1 U4443 ( .B1(n4273), .B2(n3166), .A(n3609), .ZN(n3610) );
  NAND2_X1 U4444 ( .A1(n3611), .A2(n3610), .ZN(n3684) );
  NOR2_X1 U4445 ( .A1(n3611), .A2(n3610), .ZN(n3686) );
  NAND2_X1 U4446 ( .A1(n4251), .A2(n2253), .ZN(n3613) );
  NAND2_X1 U4447 ( .A1(n4255), .A2(n3131), .ZN(n3612) );
  NAND2_X1 U4448 ( .A1(n3613), .A2(n3612), .ZN(n3614) );
  XNOR2_X1 U4449 ( .A(n3614), .B(n3627), .ZN(n3619) );
  INV_X1 U4450 ( .A(n3619), .ZN(n3617) );
  NOR2_X1 U4451 ( .A1(n4042), .A2(n3623), .ZN(n3615) );
  AOI21_X1 U4452 ( .B1(n4251), .B2(n3166), .A(n3615), .ZN(n3618) );
  INV_X1 U4453 ( .A(n3618), .ZN(n3616) );
  NAND2_X1 U4454 ( .A1(n3617), .A2(n3616), .ZN(n3754) );
  AND2_X1 U4455 ( .A1(n3619), .A2(n3618), .ZN(n3753) );
  AOI21_X1 U4456 ( .B1(n3752), .B2(n3754), .A(n3753), .ZN(n3648) );
  OAI22_X1 U4457 ( .A1(n4258), .A2(n3621), .B1(n3620), .B2(n2850), .ZN(n3622)
         );
  XNOR2_X1 U4458 ( .A(n3622), .B(n3627), .ZN(n3633) );
  OAI22_X1 U4459 ( .A1(n4258), .A2(n3624), .B1(n3623), .B2(n2850), .ZN(n3631)
         );
  XNOR2_X1 U4460 ( .A(n3633), .B(n3631), .ZN(n3647) );
  NAND2_X1 U4461 ( .A1(n3648), .A2(n3647), .ZN(n3646) );
  NAND2_X1 U4462 ( .A1(n4023), .A2(n2253), .ZN(n3626) );
  NAND2_X1 U4463 ( .A1(n3994), .A2(n3131), .ZN(n3625) );
  NAND2_X1 U4464 ( .A1(n3626), .A2(n3625), .ZN(n3628) );
  XNOR2_X1 U4465 ( .A(n3628), .B(n3627), .ZN(n3630) );
  AOI22_X1 U4466 ( .A1(n4023), .A2(n3166), .B1(n2253), .B2(n3994), .ZN(n3629)
         );
  XNOR2_X1 U4467 ( .A(n3630), .B(n3629), .ZN(n3638) );
  NAND2_X1 U4468 ( .A1(n3638), .A2(n4667), .ZN(n3645) );
  INV_X1 U4469 ( .A(n3631), .ZN(n3632) );
  NOR2_X1 U4470 ( .A1(n3633), .A2(n3632), .ZN(n3637) );
  NOR3_X1 U4471 ( .A1(n3637), .A2(n3638), .A3(n3775), .ZN(n3634) );
  NAND2_X1 U4472 ( .A1(n3646), .A2(n3634), .ZN(n3644) );
  AOI22_X1 U4473 ( .A1(n4008), .A2(n4669), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3636) );
  NAND2_X1 U4474 ( .A1(n4671), .A2(n3994), .ZN(n3635) );
  OAI211_X1 U4475 ( .C1(n4258), .C2(n3768), .A(n3636), .B(n3635), .ZN(n3642)
         );
  INV_X1 U4476 ( .A(n3637), .ZN(n3640) );
  INV_X1 U4477 ( .A(n3638), .ZN(n3639) );
  NOR3_X1 U4478 ( .A1(n3640), .A2(n3639), .A3(n3775), .ZN(n3641) );
  AOI211_X1 U4479 ( .C1(n4009), .C2(n2236), .A(n3642), .B(n3641), .ZN(n3643)
         );
  OAI211_X1 U4480 ( .C1(n3646), .C2(n3645), .A(n3644), .B(n3643), .ZN(U3217)
         );
  XNOR2_X1 U4481 ( .A(n3648), .B(n3647), .ZN(n3654) );
  INV_X1 U4482 ( .A(n3649), .ZN(n4024) );
  INV_X1 U4483 ( .A(n4251), .ZN(n4266) );
  OAI22_X1 U4484 ( .A1(n4266), .A2(n3768), .B1(n2237), .B2(n2850), .ZN(n3652)
         );
  INV_X1 U4485 ( .A(n4023), .ZN(n4247) );
  OAI22_X1 U4486 ( .A1(n4247), .A2(n3760), .B1(STATE_REG_SCAN_IN), .B2(n3650), 
        .ZN(n3651) );
  AOI211_X1 U4487 ( .C1(n4024), .C2(n2236), .A(n3652), .B(n3651), .ZN(n3653)
         );
  OAI21_X1 U4488 ( .B1(n3654), .B2(n3775), .A(n3653), .ZN(U3211) );
  NAND2_X1 U4489 ( .A1(n3655), .A2(n4667), .ZN(n3665) );
  AOI21_X1 U4490 ( .B1(n3656), .B2(n3658), .A(n3657), .ZN(n3664) );
  OAI22_X1 U4491 ( .A1(n4087), .A2(n3760), .B1(STATE_REG_SCAN_IN), .B2(n3659), 
        .ZN(n3662) );
  OAI22_X1 U4492 ( .A1(n2237), .A2(n4092), .B1(n3660), .B2(n3768), .ZN(n3661)
         );
  AOI211_X1 U4493 ( .C1(n2236), .C2(n4094), .A(n3662), .B(n3661), .ZN(n3663)
         );
  OAI21_X1 U4494 ( .B1(n3665), .B2(n3664), .A(n3663), .ZN(U3213) );
  AOI21_X1 U4495 ( .B1(n3668), .B2(n3667), .A(n2282), .ZN(n3672) );
  NOR2_X1 U4496 ( .A1(n4915), .A2(STATE_REG_SCAN_IN), .ZN(n3978) );
  OAI22_X1 U4497 ( .A1(n2237), .A2(n4176), .B1(n4209), .B2(n3768), .ZN(n3669)
         );
  AOI211_X1 U4498 ( .C1(n4669), .C2(n4121), .A(n3978), .B(n3669), .ZN(n3671)
         );
  NAND2_X1 U4499 ( .A1(n2236), .A2(n4177), .ZN(n3670) );
  OAI211_X1 U4500 ( .C1(n3672), .C2(n3775), .A(n3671), .B(n3670), .ZN(U3216)
         );
  INV_X1 U4501 ( .A(n3673), .ZN(n3675) );
  NAND2_X1 U4502 ( .A1(n3675), .A2(n3674), .ZN(n3677) );
  OAI211_X1 U4503 ( .C1(n3723), .C2(n2308), .A(n3724), .B(n3677), .ZN(n3676)
         );
  OAI211_X1 U4504 ( .C1(n3678), .C2(n3677), .A(n4667), .B(n3676), .ZN(n3683)
         );
  AOI22_X1 U4505 ( .A1(n4669), .A2(n4129), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3682) );
  AOI22_X1 U4506 ( .A1(n4671), .A2(n4128), .B1(n3746), .B2(n4121), .ZN(n3681)
         );
  NAND2_X1 U4507 ( .A1(n2236), .A2(n3679), .ZN(n3680) );
  NAND4_X1 U4508 ( .A1(n3683), .A2(n3682), .A3(n3681), .A4(n3680), .ZN(U3220)
         );
  INV_X1 U4509 ( .A(n3684), .ZN(n3685) );
  NOR2_X1 U4510 ( .A1(n3686), .A2(n3685), .ZN(n3687) );
  XNOR2_X1 U4511 ( .A(n3688), .B(n3687), .ZN(n3693) );
  INV_X1 U4512 ( .A(n3689), .ZN(n4049) );
  OAI22_X1 U4513 ( .A1(n4266), .A2(n3760), .B1(STATE_REG_SCAN_IN), .B2(n4930), 
        .ZN(n3691) );
  OAI22_X1 U4514 ( .A1(n2237), .A2(n4052), .B1(n4087), .B2(n3768), .ZN(n3690)
         );
  AOI211_X1 U4515 ( .C1(n2236), .C2(n4049), .A(n3691), .B(n3690), .ZN(n3692)
         );
  OAI21_X1 U4516 ( .B1(n3693), .B2(n3775), .A(n3692), .ZN(U3222) );
  INV_X1 U4517 ( .A(n3765), .ZN(n3695) );
  OAI21_X1 U4518 ( .B1(n3695), .B2(n3767), .A(n3694), .ZN(n3696) );
  XOR2_X1 U4519 ( .A(n3697), .B(n3696), .Z(n3705) );
  INV_X1 U4520 ( .A(REG3_REG_16__SCAN_IN), .ZN(n3698) );
  NOR2_X1 U4521 ( .A1(STATE_REG_SCAN_IN), .A2(n3698), .ZN(n3965) );
  OAI22_X1 U4522 ( .A1(n2237), .A2(n3700), .B1(n3699), .B2(n3768), .ZN(n3701)
         );
  AOI211_X1 U4523 ( .C1(n4669), .C2(n3745), .A(n3965), .B(n3701), .ZN(n3704)
         );
  NAND2_X1 U4524 ( .A1(n2236), .A2(n3702), .ZN(n3703) );
  OAI211_X1 U4525 ( .C1(n3705), .C2(n3775), .A(n3704), .B(n3703), .ZN(U3223)
         );
  NAND2_X1 U4526 ( .A1(n3708), .A2(n3707), .ZN(n3709) );
  XNOR2_X1 U4527 ( .A(n3706), .B(n3709), .ZN(n3714) );
  AND2_X1 U4528 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4542) );
  OAI22_X1 U4529 ( .A1(n2237), .A2(n4208), .B1(n3710), .B2(n3768), .ZN(n3711)
         );
  AOI211_X1 U4530 ( .C1(n4669), .C2(n4172), .A(n4542), .B(n3711), .ZN(n3713)
         );
  NAND2_X1 U4531 ( .A1(n2236), .A2(n4218), .ZN(n3712) );
  OAI211_X1 U4532 ( .C1(n3714), .C2(n3775), .A(n3713), .B(n3712), .ZN(U3225)
         );
  OAI22_X1 U4533 ( .A1(n3758), .A2(n3760), .B1(STATE_REG_SCAN_IN), .B2(n3717), 
        .ZN(n3719) );
  OAI22_X1 U4534 ( .A1(n2237), .A2(n4072), .B1(n4276), .B2(n3768), .ZN(n3718)
         );
  AOI211_X1 U4535 ( .C1(n2236), .C2(n4068), .A(n3719), .B(n3718), .ZN(n3720)
         );
  OAI21_X1 U4536 ( .B1(n3721), .B2(n3775), .A(n3720), .ZN(U3226) );
  INV_X1 U4537 ( .A(n3722), .ZN(n3727) );
  AOI21_X1 U4538 ( .B1(n3724), .B2(n3726), .A(n3723), .ZN(n3725) );
  AOI21_X1 U4539 ( .B1(n3727), .B2(n3726), .A(n3725), .ZN(n3732) );
  OAI22_X1 U4540 ( .A1(n4108), .A2(n3760), .B1(STATE_REG_SCAN_IN), .B2(n3728), 
        .ZN(n3730) );
  OAI22_X1 U4541 ( .A1(n2237), .A2(n4149), .B1(n4296), .B2(n3768), .ZN(n3729)
         );
  AOI211_X1 U4542 ( .C1(n2236), .C2(n4153), .A(n3730), .B(n3729), .ZN(n3731)
         );
  OAI21_X1 U4543 ( .B1(n3732), .B2(n3775), .A(n3731), .ZN(U3230) );
  INV_X1 U4544 ( .A(n3656), .ZN(n3733) );
  AOI21_X1 U4545 ( .B1(n3735), .B2(n3734), .A(n3733), .ZN(n3740) );
  INV_X1 U4546 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4975) );
  OAI22_X1 U4547 ( .A1(n4276), .A2(n3760), .B1(STATE_REG_SCAN_IN), .B2(n4975), 
        .ZN(n3737) );
  OAI22_X1 U4548 ( .A1(n2237), .A2(n4112), .B1(n4108), .B2(n3768), .ZN(n3736)
         );
  AOI211_X1 U4549 ( .C1(n2236), .C2(n4113), .A(n3737), .B(n3736), .ZN(n3739)
         );
  OAI21_X1 U4550 ( .B1(n3740), .B2(n3775), .A(n3739), .ZN(U3232) );
  XNOR2_X1 U4551 ( .A(n3743), .B(n3742), .ZN(n3744) );
  XNOR2_X1 U4552 ( .A(n3741), .B(n3744), .ZN(n3751) );
  AOI22_X1 U4553 ( .A1(n4671), .A2(n4184), .B1(n3746), .B2(n3745), .ZN(n3748)
         );
  OAI211_X1 U4554 ( .C1(n4296), .C2(n3760), .A(n3748), .B(n3747), .ZN(n3749)
         );
  AOI21_X1 U4555 ( .B1(n2236), .B2(n4197), .A(n3749), .ZN(n3750) );
  OAI21_X1 U4556 ( .B1(n3751), .B2(n3775), .A(n3750), .ZN(U3235) );
  INV_X1 U4557 ( .A(n3753), .ZN(n3755) );
  NAND2_X1 U4558 ( .A1(n3755), .A2(n3754), .ZN(n3756) );
  XNOR2_X1 U4559 ( .A(n3752), .B(n3756), .ZN(n3764) );
  OAI22_X1 U4560 ( .A1(n3758), .A2(n3768), .B1(n2237), .B2(n4042), .ZN(n3762)
         );
  OAI22_X1 U4561 ( .A1(n4258), .A2(n3760), .B1(STATE_REG_SCAN_IN), .B2(n3759), 
        .ZN(n3761) );
  AOI211_X1 U4562 ( .C1(n2236), .C2(n4039), .A(n3762), .B(n3761), .ZN(n3763)
         );
  OAI21_X1 U4563 ( .B1(n3764), .B2(n3775), .A(n3763), .ZN(U3237) );
  NAND2_X1 U4564 ( .A1(n3765), .A2(n3694), .ZN(n3766) );
  XOR2_X1 U4565 ( .A(n3767), .B(n3766), .Z(n3776) );
  AND2_X1 U4566 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n3955) );
  OAI22_X1 U4567 ( .A1(n2237), .A2(n3770), .B1(n3769), .B2(n3768), .ZN(n3771)
         );
  AOI211_X1 U4568 ( .C1(n4669), .C2(n4211), .A(n3955), .B(n3771), .ZN(n3774)
         );
  NAND2_X1 U4569 ( .A1(n2236), .A2(n3772), .ZN(n3773) );
  OAI211_X1 U4570 ( .C1(n3776), .C2(n3775), .A(n3774), .B(n3773), .ZN(U3238)
         );
  INV_X1 U4571 ( .A(n3872), .ZN(n3777) );
  NOR2_X1 U4572 ( .A1(n3778), .A2(n3777), .ZN(n3905) );
  OAI211_X1 U4573 ( .C1(n3781), .C2(n3920), .A(n3780), .B(n3779), .ZN(n3783)
         );
  NAND3_X1 U4574 ( .A1(n3783), .A2(n3782), .A3(n2873), .ZN(n3786) );
  NAND3_X1 U4575 ( .A1(n3786), .A2(n3785), .A3(n3784), .ZN(n3789) );
  NAND3_X1 U4576 ( .A1(n3789), .A2(n3788), .A3(n3787), .ZN(n3792) );
  NAND4_X1 U4577 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3804), .ZN(n3794)
         );
  AND3_X1 U4578 ( .A1(n3794), .A2(n3856), .A3(n3793), .ZN(n3799) );
  NAND2_X1 U4579 ( .A1(n3796), .A2(n3795), .ZN(n3803) );
  OAI211_X1 U4580 ( .C1(n3799), .C2(n3803), .A(n3798), .B(n3797), .ZN(n3811)
         );
  NAND2_X1 U4581 ( .A1(n3801), .A2(n3800), .ZN(n3807) );
  INV_X1 U4582 ( .A(n3807), .ZN(n3810) );
  INV_X1 U4583 ( .A(n3802), .ZN(n3806) );
  INV_X1 U4584 ( .A(n3803), .ZN(n3805) );
  NAND3_X1 U4585 ( .A1(n3806), .A2(n3805), .A3(n3804), .ZN(n3808) );
  AND2_X1 U4586 ( .A1(n3807), .A2(n3819), .ZN(n3889) );
  AOI21_X1 U4587 ( .B1(n3812), .B2(n3808), .A(n3889), .ZN(n3809) );
  AOI21_X1 U4588 ( .B1(n3811), .B2(n3810), .A(n3809), .ZN(n3818) );
  INV_X1 U4589 ( .A(n3812), .ZN(n3815) );
  OAI211_X1 U4590 ( .C1(n3815), .C2(n2287), .A(n3814), .B(n3813), .ZN(n3816)
         );
  NOR3_X1 U4591 ( .A1(n3818), .A2(n3817), .A3(n3816), .ZN(n3823) );
  AND2_X1 U4592 ( .A1(n3820), .A2(n3819), .ZN(n3890) );
  AOI21_X1 U4593 ( .B1(n3821), .B2(n3890), .A(n3889), .ZN(n3822) );
  OAI21_X1 U4594 ( .B1(n3823), .B2(n3822), .A(n3894), .ZN(n3824) );
  AOI21_X1 U4595 ( .B1(n3824), .B2(n3892), .A(n3893), .ZN(n3826) );
  INV_X1 U4596 ( .A(n3825), .ZN(n4124) );
  OAI21_X1 U4597 ( .B1(n3826), .B2(n4124), .A(n3903), .ZN(n3828) );
  NAND3_X1 U4598 ( .A1(n3828), .A2(n3827), .A3(n4083), .ZN(n3831) );
  OAI211_X1 U4599 ( .C1(n3829), .C2(n3900), .A(n3871), .B(n3845), .ZN(n3906)
         );
  INV_X1 U4600 ( .A(n3906), .ZN(n3830) );
  OAI21_X1 U4601 ( .B1(n3901), .B2(n3831), .A(n3830), .ZN(n3835) );
  NAND2_X1 U4602 ( .A1(n2835), .A2(DATAI_29_), .ZN(n4241) );
  NAND2_X1 U4603 ( .A1(n4008), .A2(n4241), .ZN(n3879) );
  NAND2_X1 U4604 ( .A1(n3879), .A2(n3986), .ZN(n3837) );
  NOR2_X1 U4605 ( .A1(n3832), .A2(n3837), .ZN(n3912) );
  INV_X1 U4606 ( .A(n3912), .ZN(n3833) );
  AOI211_X1 U4607 ( .C1(n3905), .C2(n3835), .A(n3834), .B(n3833), .ZN(n3839)
         );
  NOR2_X1 U4608 ( .A1(n3985), .A2(n3909), .ZN(n3838) );
  AND2_X1 U4609 ( .A1(n2835), .A2(DATAI_30_), .ZN(n4234) );
  NAND2_X1 U4610 ( .A1(n3989), .A2(n4234), .ZN(n3836) );
  NAND2_X1 U4611 ( .A1(n2835), .A2(DATAI_31_), .ZN(n4227) );
  NAND2_X1 U4612 ( .A1(n3914), .A2(n4227), .ZN(n3842) );
  AND2_X1 U4613 ( .A1(n3836), .A2(n3842), .ZN(n3880) );
  OR2_X1 U4614 ( .A1(n4008), .A2(n4241), .ZN(n3904) );
  OAI211_X1 U4615 ( .C1(n3838), .C2(n3837), .A(n3880), .B(n3904), .ZN(n3911)
         );
  OR2_X1 U4616 ( .A1(n3839), .A2(n3911), .ZN(n3844) );
  OR2_X1 U4617 ( .A1(n3989), .A2(n4234), .ZN(n3915) );
  INV_X1 U4618 ( .A(n3914), .ZN(n4226) );
  INV_X1 U4619 ( .A(n4227), .ZN(n3840) );
  NAND2_X1 U4620 ( .A1(n4226), .A2(n3840), .ZN(n3841) );
  NAND2_X1 U4621 ( .A1(n3915), .A2(n3841), .ZN(n3860) );
  NAND2_X1 U4622 ( .A1(n3860), .A2(n3842), .ZN(n3843) );
  NAND2_X1 U4623 ( .A1(n3844), .A2(n3843), .ZN(n3925) );
  AND2_X1 U4624 ( .A1(n3846), .A2(n3845), .ZN(n4064) );
  AND2_X1 U4625 ( .A1(n3847), .A2(n4059), .ZN(n4086) );
  INV_X1 U4626 ( .A(n3848), .ZN(n3850) );
  AND2_X1 U4627 ( .A1(n3850), .A2(n3849), .ZN(n4168) );
  INV_X1 U4628 ( .A(n3851), .ZN(n3853) );
  OR2_X1 U4629 ( .A1(n3853), .A2(n3852), .ZN(n4143) );
  INV_X1 U4630 ( .A(n4143), .ZN(n4146) );
  NAND2_X1 U4631 ( .A1(n4162), .A2(n4078), .ZN(n4207) );
  NOR4_X1 U4632 ( .A1(n4168), .A2(n4146), .A3(n4182), .A4(n4207), .ZN(n3854)
         );
  NAND3_X1 U4633 ( .A1(n4064), .A2(n4086), .A3(n3854), .ZN(n3888) );
  INV_X1 U4634 ( .A(n4019), .ZN(n3913) );
  AND2_X1 U4635 ( .A1(n4083), .A2(n3903), .ZN(n4123) );
  NAND4_X1 U4636 ( .A1(n2407), .A2(n3858), .A3(n3857), .A4(n3856), .ZN(n3866)
         );
  INV_X1 U4637 ( .A(n3859), .ZN(n3864) );
  INV_X1 U4638 ( .A(n3860), .ZN(n3863) );
  NAND4_X1 U4639 ( .A1(n3864), .A2(n3863), .A3(n3862), .A4(n3861), .ZN(n3865)
         );
  NOR2_X1 U4640 ( .A1(n3866), .A2(n3865), .ZN(n3870) );
  INV_X1 U4641 ( .A(n3867), .ZN(n3868) );
  NOR2_X1 U4642 ( .A1(n3869), .A2(n3868), .ZN(n4034) );
  INV_X1 U4643 ( .A(n4034), .ZN(n4031) );
  NAND4_X1 U4644 ( .A1(n3913), .A2(n4123), .A3(n3870), .A4(n4031), .ZN(n3887)
         );
  NAND2_X1 U4645 ( .A1(n3872), .A2(n3871), .ZN(n4053) );
  NOR3_X1 U4646 ( .A1(n3992), .A2(n4103), .A3(n4053), .ZN(n3885) );
  INV_X1 U4647 ( .A(n3873), .ZN(n3875) );
  NOR4_X1 U4648 ( .A1(n2679), .A2(n3875), .A3(n2872), .A4(n3874), .ZN(n3884)
         );
  NOR4_X1 U4649 ( .A1(n2423), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3883)
         );
  NAND2_X1 U4650 ( .A1(n3904), .A2(n3879), .ZN(n3997) );
  INV_X1 U4651 ( .A(n3880), .ZN(n3908) );
  NOR4_X1 U4652 ( .A1(n3997), .A2(n3908), .A3(n3881), .A4(n4588), .ZN(n3882)
         );
  NAND4_X1 U4653 ( .A1(n3885), .A2(n3884), .A3(n3883), .A4(n3882), .ZN(n3886)
         );
  OR3_X1 U4654 ( .A1(n3888), .A2(n3887), .A3(n3886), .ZN(n3922) );
  AOI21_X1 U4655 ( .B1(n3891), .B2(n3890), .A(n3889), .ZN(n3897) );
  INV_X1 U4656 ( .A(n3892), .ZN(n3896) );
  INV_X1 U4657 ( .A(n3893), .ZN(n3895) );
  OAI211_X1 U4658 ( .C1(n3897), .C2(n3896), .A(n3895), .B(n3894), .ZN(n3899)
         );
  NAND2_X1 U4659 ( .A1(n3899), .A2(n3898), .ZN(n3902) );
  AOI211_X1 U4660 ( .C1(n3903), .C2(n3902), .A(n3901), .B(n3900), .ZN(n3907)
         );
  OAI211_X1 U4661 ( .C1(n3907), .C2(n3906), .A(n3905), .B(n3904), .ZN(n3910)
         );
  NOR4_X1 U4662 ( .A1(n3910), .A2(n3985), .A3(n3909), .A4(n3908), .ZN(n3918)
         );
  AOI21_X1 U4663 ( .B1(n3913), .B2(n3912), .A(n3911), .ZN(n3917) );
  AOI21_X1 U4664 ( .B1(n3915), .B2(n3914), .A(n4227), .ZN(n3916) );
  NOR3_X1 U4665 ( .A1(n3918), .A2(n3917), .A3(n3916), .ZN(n3919) );
  AOI21_X1 U4666 ( .B1(n4234), .B2(n4227), .A(n3919), .ZN(n3921) );
  MUX2_X1 U4667 ( .A(n3922), .B(n3921), .S(n3920), .Z(n3924) );
  MUX2_X1 U4668 ( .A(n3925), .B(n3924), .S(n3923), .Z(n3926) );
  XNOR2_X1 U4669 ( .A(n3926), .B(n3980), .ZN(n3932) );
  NOR2_X1 U4670 ( .A1(n4417), .A2(n3927), .ZN(n3930) );
  OAI21_X1 U4671 ( .B1(n3931), .B2(n3928), .A(B_REG_SCAN_IN), .ZN(n3929) );
  OAI22_X1 U4672 ( .A1(n3932), .A2(n3931), .B1(n3930), .B2(n3929), .ZN(U3239)
         );
  MUX2_X1 U4673 ( .A(n4008), .B(DATAO_REG_29__SCAN_IN), .S(n4418), .Z(U3579)
         );
  MUX2_X1 U4674 ( .A(n4023), .B(DATAO_REG_28__SCAN_IN), .S(n4418), .Z(U3578)
         );
  MUX2_X1 U4675 ( .A(DATAO_REG_27__SCAN_IN), .B(n4038), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4676 ( .A(n4273), .B(DATAO_REG_25__SCAN_IN), .S(n4418), .Z(U3575)
         );
  MUX2_X1 U4677 ( .A(n4129), .B(DATAO_REG_22__SCAN_IN), .S(n4418), .Z(U3572)
         );
  MUX2_X1 U4678 ( .A(n4293), .B(DATAO_REG_21__SCAN_IN), .S(n4418), .Z(U3571)
         );
  MUX2_X1 U4679 ( .A(n4121), .B(DATAO_REG_20__SCAN_IN), .S(n4418), .Z(U3570)
         );
  MUX2_X1 U4680 ( .A(DATAO_REG_19__SCAN_IN), .B(n4185), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4681 ( .A(DATAO_REG_18__SCAN_IN), .B(n4172), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4682 ( .A(DATAO_REG_16__SCAN_IN), .B(n4211), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4683 ( .A(n4325), .B(DATAO_REG_15__SCAN_IN), .S(n4418), .Z(U3565)
         );
  MUX2_X1 U4684 ( .A(DATAO_REG_14__SCAN_IN), .B(n3933), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4685 ( .A(n4636), .B(DATAO_REG_12__SCAN_IN), .S(n4418), .Z(U3562)
         );
  MUX2_X1 U4686 ( .A(n4638), .B(DATAO_REG_10__SCAN_IN), .S(n4418), .Z(U3560)
         );
  MUX2_X1 U4687 ( .A(n3934), .B(DATAO_REG_9__SCAN_IN), .S(n4418), .Z(U3559) );
  MUX2_X1 U4688 ( .A(n3935), .B(DATAO_REG_6__SCAN_IN), .S(n4418), .Z(U3556) );
  MUX2_X1 U4689 ( .A(n3936), .B(DATAO_REG_5__SCAN_IN), .S(n4418), .Z(U3555) );
  MUX2_X1 U4690 ( .A(DATAO_REG_4__SCAN_IN), .B(n3937), .S(U4043), .Z(U3554) );
  MUX2_X1 U4691 ( .A(n3938), .B(DATAO_REG_3__SCAN_IN), .S(n4418), .Z(U3553) );
  MUX2_X1 U4692 ( .A(DATAO_REG_2__SCAN_IN), .B(n3939), .S(U4043), .Z(U3552) );
  MUX2_X1 U4693 ( .A(DATAO_REG_1__SCAN_IN), .B(n2669), .S(U4043), .Z(U3551) );
  INV_X1 U4694 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4650) );
  NOR2_X1 U4695 ( .A1(n2335), .A2(n4650), .ZN(n3942) );
  OAI211_X1 U4696 ( .C1(n3942), .C2(n3941), .A(n4553), .B(n3940), .ZN(n3949)
         );
  INV_X1 U4697 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4405) );
  NOR2_X1 U4698 ( .A1(n2335), .A2(n4405), .ZN(n4419) );
  OAI211_X1 U4699 ( .C1(n4419), .C2(n3944), .A(n4551), .B(n3943), .ZN(n3948)
         );
  AOI22_X1 U4700 ( .A1(n4543), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3947) );
  NAND2_X1 U4701 ( .A1(n4538), .A2(n3945), .ZN(n3946) );
  NAND4_X1 U4702 ( .A1(n3949), .A2(n3948), .A3(n3947), .A4(n3946), .ZN(U3241)
         );
  INV_X1 U4703 ( .A(n3950), .ZN(n3961) );
  AOI211_X1 U4704 ( .C1(n3953), .C2(n3952), .A(n3951), .B(n4528), .ZN(n3954)
         );
  AOI211_X1 U4705 ( .C1(n4543), .C2(ADDR_REG_15__SCAN_IN), .A(n3955), .B(n3954), .ZN(n3960) );
  AOI21_X1 U4706 ( .B1(n3957), .B2(n2260), .A(n3956), .ZN(n3958) );
  NAND2_X1 U4707 ( .A1(n4553), .A2(n3958), .ZN(n3959) );
  OAI211_X1 U4708 ( .C1(n4556), .C2(n3961), .A(n3960), .B(n3959), .ZN(U3255)
         );
  OAI21_X1 U4709 ( .B1(n3963), .B2(n4951), .A(n3962), .ZN(n3964) );
  NAND2_X1 U4710 ( .A1(n3964), .A2(n4553), .ZN(n3973) );
  AOI21_X1 U4711 ( .B1(n4543), .B2(ADDR_REG_16__SCAN_IN), .A(n3965), .ZN(n3972) );
  OAI21_X1 U4712 ( .B1(n3968), .B2(n3967), .A(n3966), .ZN(n3969) );
  NAND2_X1 U4713 ( .A1(n3969), .A2(n4551), .ZN(n3971) );
  NAND2_X1 U4714 ( .A1(n4538), .A2(n4383), .ZN(n3970) );
  NAND4_X1 U4715 ( .A1(n3973), .A2(n3972), .A3(n3971), .A4(n3970), .ZN(U3256)
         );
  INV_X1 U4716 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4976) );
  MUX2_X1 U4717 ( .A(n4976), .B(REG2_REG_19__SCAN_IN), .S(n3980), .Z(n3976) );
  XNOR2_X1 U4718 ( .A(n3977), .B(n3976), .ZN(n3982) );
  AOI21_X1 U4719 ( .B1(n4543), .B2(ADDR_REG_19__SCAN_IN), .A(n3978), .ZN(n3979) );
  OAI21_X1 U4720 ( .B1(n3980), .B2(n4556), .A(n3979), .ZN(n3981) );
  AOI21_X1 U4721 ( .B1(n3982), .B2(n4551), .A(n3981), .ZN(n3983) );
  INV_X1 U4722 ( .A(n3984), .ZN(n3991) );
  AOI21_X1 U4723 ( .B1(n3987), .B2(n3986), .A(n3985), .ZN(n3988) );
  XOR2_X1 U4724 ( .A(n3997), .B(n3988), .Z(n3990) );
  INV_X1 U4725 ( .A(B_REG_SCAN_IN), .ZN(n4912) );
  OAI21_X1 U4726 ( .B1(n4912), .B2(n4406), .A(n4635), .ZN(n4225) );
  OAI22_X1 U4727 ( .A1(n3990), .A2(n4213), .B1(n3989), .B2(n4225), .ZN(n4242)
         );
  AOI21_X1 U4728 ( .B1(n3991), .B2(n4557), .A(n4242), .ZN(n4006) );
  NAND2_X1 U4729 ( .A1(n3996), .A2(n3995), .ZN(n3999) );
  XNOR2_X1 U4730 ( .A(n3999), .B(n3998), .ZN(n4240) );
  NAND2_X1 U4731 ( .A1(n4240), .A2(n4201), .ZN(n4005) );
  INV_X1 U4732 ( .A(n4241), .ZN(n4001) );
  AOI21_X1 U4733 ( .B1(n4001), .B2(n4000), .A(n4230), .ZN(n4244) );
  AOI22_X1 U4734 ( .A1(n4023), .A2(n4066), .B1(n4204), .B2(
        REG2_REG_29__SCAN_IN), .ZN(n4002) );
  OAI21_X1 U4735 ( .B1(n4241), .B2(n4071), .A(n4002), .ZN(n4003) );
  AOI21_X1 U4736 ( .B1(n4244), .B2(n4560), .A(n4003), .ZN(n4004) );
  OAI211_X1 U4737 ( .C1(n4566), .C2(n4006), .A(n4005), .B(n4004), .ZN(U3354)
         );
  NOR2_X1 U4738 ( .A1(n4007), .A2(n4220), .ZN(n4014) );
  AOI22_X1 U4739 ( .A1(n4038), .A2(n4066), .B1(n4151), .B2(n4008), .ZN(n4011)
         );
  AOI22_X1 U4740 ( .A1(n4009), .A2(n4557), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4204), .ZN(n4010) );
  OAI211_X1 U4741 ( .C1(n4012), .C2(n4071), .A(n4011), .B(n4010), .ZN(n4013)
         );
  AOI211_X1 U4742 ( .C1(n4015), .C2(n4402), .A(n4014), .B(n4013), .ZN(n4016)
         );
  OAI21_X1 U4743 ( .B1(n4017), .B2(n4223), .A(n4016), .ZN(U3262) );
  XNOR2_X1 U4744 ( .A(n4018), .B(n4019), .ZN(n4254) );
  XNOR2_X1 U4745 ( .A(n4020), .B(n4019), .ZN(n4021) );
  NAND2_X1 U4746 ( .A1(n4021), .A2(n4189), .ZN(n4252) );
  INV_X1 U4747 ( .A(n4252), .ZN(n4029) );
  OAI21_X1 U4748 ( .B1(n4036), .B2(n2850), .A(n4022), .ZN(n4248) );
  NOR2_X1 U4749 ( .A1(n4248), .A2(n4220), .ZN(n4028) );
  AOI22_X1 U4750 ( .A1(n4023), .A2(n4151), .B1(n4066), .B2(n4251), .ZN(n4026)
         );
  AOI22_X1 U4751 ( .A1(n4024), .A2(n4557), .B1(n4204), .B2(
        REG2_REG_27__SCAN_IN), .ZN(n4025) );
  OAI211_X1 U4752 ( .C1(n2850), .C2(n4071), .A(n4026), .B(n4025), .ZN(n4027)
         );
  AOI211_X1 U4753 ( .C1(n4029), .C2(n4402), .A(n4028), .B(n4027), .ZN(n4030)
         );
  OAI21_X1 U4754 ( .B1(n4254), .B2(n4223), .A(n4030), .ZN(U3263) );
  XNOR2_X1 U4755 ( .A(n4032), .B(n4031), .ZN(n4033) );
  NAND2_X1 U4756 ( .A1(n4033), .A2(n4189), .ZN(n4257) );
  XNOR2_X1 U4757 ( .A(n4035), .B(n4034), .ZN(n4260) );
  NAND2_X1 U4758 ( .A1(n4260), .A2(n4201), .ZN(n4046) );
  INV_X1 U4759 ( .A(n4036), .ZN(n4037) );
  OAI21_X1 U4760 ( .B1(n4048), .B2(n4042), .A(n4037), .ZN(n4343) );
  INV_X1 U4761 ( .A(n4343), .ZN(n4044) );
  AOI22_X1 U4762 ( .A1(n4038), .A2(n4151), .B1(n4066), .B2(n4273), .ZN(n4041)
         );
  AOI22_X1 U4763 ( .A1(n4039), .A2(n4557), .B1(n4204), .B2(
        REG2_REG_26__SCAN_IN), .ZN(n4040) );
  OAI211_X1 U4764 ( .C1(n4042), .C2(n4071), .A(n4041), .B(n4040), .ZN(n4043)
         );
  AOI21_X1 U4765 ( .B1(n4044), .B2(n4560), .A(n4043), .ZN(n4045) );
  OAI211_X1 U4766 ( .C1(n4566), .C2(n4257), .A(n4046), .B(n4045), .ZN(U3264)
         );
  XNOR2_X1 U4767 ( .A(n4047), .B(n4053), .ZN(n4271) );
  AOI21_X1 U4768 ( .B1(n4263), .B2(n2276), .A(n4048), .ZN(n4268) );
  AOI22_X1 U4769 ( .A1(n4251), .A2(n4151), .B1(n4066), .B2(n4264), .ZN(n4051)
         );
  AOI22_X1 U4770 ( .A1(n4204), .A2(REG2_REG_25__SCAN_IN), .B1(n4049), .B2(
        n4557), .ZN(n4050) );
  OAI211_X1 U4771 ( .C1(n4052), .C2(n4071), .A(n4051), .B(n4050), .ZN(n4057)
         );
  XNOR2_X1 U4772 ( .A(n4054), .B(n4053), .ZN(n4055) );
  NAND2_X1 U4773 ( .A1(n4055), .A2(n4189), .ZN(n4269) );
  NOR2_X1 U4774 ( .A1(n4269), .A2(n4566), .ZN(n4056) );
  AOI211_X1 U4775 ( .C1(n4268), .C2(n4560), .A(n4057), .B(n4056), .ZN(n4058)
         );
  OAI21_X1 U4776 ( .B1(n4271), .B2(n4223), .A(n4058), .ZN(U3265) );
  NAND2_X1 U4777 ( .A1(n4060), .A2(n4059), .ZN(n4061) );
  XNOR2_X1 U4778 ( .A(n4061), .B(n4064), .ZN(n4062) );
  NAND2_X1 U4779 ( .A1(n4062), .A2(n4189), .ZN(n4275) );
  XOR2_X1 U4780 ( .A(n4064), .B(n4063), .Z(n4278) );
  NAND2_X1 U4781 ( .A1(n4278), .A2(n4201), .ZN(n4076) );
  INV_X1 U4782 ( .A(n4091), .ZN(n4065) );
  OAI21_X1 U4783 ( .B1(n4065), .B2(n4072), .A(n2276), .ZN(n4348) );
  INV_X1 U4784 ( .A(n4348), .ZN(n4074) );
  AOI22_X1 U4785 ( .A1(n4273), .A2(n4151), .B1(n4067), .B2(n4066), .ZN(n4070)
         );
  AOI22_X1 U4786 ( .A1(n4204), .A2(REG2_REG_24__SCAN_IN), .B1(n4068), .B2(
        n4557), .ZN(n4069) );
  OAI211_X1 U4787 ( .C1(n4072), .C2(n4071), .A(n4070), .B(n4069), .ZN(n4073)
         );
  AOI21_X1 U4788 ( .B1(n4074), .B2(n4560), .A(n4073), .ZN(n4075) );
  OAI211_X1 U4789 ( .C1(n4566), .C2(n4275), .A(n4076), .B(n4075), .ZN(U3266)
         );
  INV_X1 U4790 ( .A(n4281), .ZN(n4100) );
  INV_X1 U4791 ( .A(n4078), .ZN(n4079) );
  NAND2_X1 U4792 ( .A1(n4164), .A2(n4080), .ZN(n4142) );
  INV_X1 U4793 ( .A(n4081), .ZN(n4082) );
  NOR2_X1 U4794 ( .A1(n4142), .A2(n4082), .ZN(n4125) );
  OAI21_X1 U4795 ( .B1(n4125), .B2(n4124), .A(n4123), .ZN(n4122) );
  NAND2_X1 U4796 ( .A1(n4122), .A2(n4083), .ZN(n4106) );
  NAND2_X1 U4797 ( .A1(n4106), .A2(n4107), .ZN(n4105) );
  NAND2_X1 U4798 ( .A1(n4105), .A2(n4084), .ZN(n4085) );
  XOR2_X1 U4799 ( .A(n4086), .B(n4085), .Z(n4090) );
  OAI22_X1 U4800 ( .A1(n4087), .A2(n4594), .B1(n4092), .B2(n4593), .ZN(n4088)
         );
  AOI21_X1 U4801 ( .B1(n4637), .B2(n4129), .A(n4088), .ZN(n4089) );
  OAI21_X1 U4802 ( .B1(n4090), .B2(n4213), .A(n4089), .ZN(n4280) );
  INV_X1 U4803 ( .A(n4284), .ZN(n4093) );
  OAI21_X1 U4804 ( .B1(n4093), .B2(n4092), .A(n4091), .ZN(n4352) );
  NOR2_X1 U4805 ( .A1(n4352), .A2(n4220), .ZN(n4098) );
  INV_X1 U4806 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4096) );
  INV_X1 U4807 ( .A(n4094), .ZN(n4095) );
  OAI22_X1 U4808 ( .A1(n4402), .A2(n4096), .B1(n4095), .B2(n4134), .ZN(n4097)
         );
  AOI211_X1 U4809 ( .C1(n4280), .C2(n4402), .A(n4098), .B(n4097), .ZN(n4099)
         );
  OAI21_X1 U4810 ( .B1(n4100), .B2(n4223), .A(n4099), .ZN(U3267) );
  INV_X1 U4811 ( .A(n4101), .ZN(n4104) );
  OAI21_X1 U4812 ( .B1(n4104), .B2(n4103), .A(n4102), .ZN(n4288) );
  OAI21_X1 U4813 ( .B1(n4107), .B2(n4106), .A(n4105), .ZN(n4111) );
  NOR2_X1 U4814 ( .A1(n4108), .A2(n4327), .ZN(n4110) );
  OAI22_X1 U4815 ( .A1(n4276), .A2(n4594), .B1(n4112), .B2(n4593), .ZN(n4109)
         );
  AOI211_X1 U4816 ( .C1(n4111), .C2(n4189), .A(n4110), .B(n4109), .ZN(n4287)
         );
  INV_X1 U4817 ( .A(n4287), .ZN(n4118) );
  NAND2_X1 U4818 ( .A1(n2272), .A2(n2815), .ZN(n4285) );
  AND3_X1 U4819 ( .A1(n4285), .A2(n4560), .A3(n4284), .ZN(n4117) );
  INV_X1 U4820 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4115) );
  INV_X1 U4821 ( .A(n4113), .ZN(n4114) );
  OAI22_X1 U4822 ( .A1(n4402), .A2(n4115), .B1(n4114), .B2(n4134), .ZN(n4116)
         );
  AOI211_X1 U4823 ( .C1(n4118), .C2(n4402), .A(n4117), .B(n4116), .ZN(n4119)
         );
  OAI21_X1 U4824 ( .B1(n4288), .B2(n4223), .A(n4119), .ZN(U3268) );
  XNOR2_X1 U4825 ( .A(n4120), .B(n4123), .ZN(n4290) );
  INV_X1 U4826 ( .A(n4290), .ZN(n4139) );
  INV_X1 U4827 ( .A(n4121), .ZN(n4170) );
  INV_X1 U4828 ( .A(n4122), .ZN(n4127) );
  NOR3_X1 U4829 ( .A1(n4125), .A2(n4124), .A3(n4123), .ZN(n4126) );
  OAI21_X1 U4830 ( .B1(n4127), .B2(n4126), .A(n4189), .ZN(n4131) );
  AOI22_X1 U4831 ( .A1(n4129), .A2(n4635), .B1(n4634), .B2(n4128), .ZN(n4130)
         );
  OAI211_X1 U4832 ( .C1(n4170), .C2(n4327), .A(n4131), .B(n4130), .ZN(n4289)
         );
  INV_X1 U4833 ( .A(n4148), .ZN(n4133) );
  OAI21_X1 U4834 ( .B1(n4133), .B2(n4132), .A(n2272), .ZN(n4357) );
  NOR2_X1 U4835 ( .A1(n4357), .A2(n4220), .ZN(n4137) );
  INV_X1 U4836 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4962) );
  OAI22_X1 U4837 ( .A1(n4402), .A2(n4962), .B1(n4135), .B2(n4134), .ZN(n4136)
         );
  AOI211_X1 U4838 ( .C1(n4289), .C2(n4402), .A(n4137), .B(n4136), .ZN(n4138)
         );
  OAI21_X1 U4839 ( .B1(n4139), .B2(n4223), .A(n4138), .ZN(U3269) );
  INV_X1 U4840 ( .A(n4140), .ZN(n4141) );
  NAND2_X1 U4841 ( .A1(n4142), .A2(n4141), .ZN(n4144) );
  XNOR2_X1 U4842 ( .A(n4144), .B(n4143), .ZN(n4145) );
  NAND2_X1 U4843 ( .A1(n4145), .A2(n4189), .ZN(n4295) );
  XNOR2_X1 U4844 ( .A(n4147), .B(n4146), .ZN(n4298) );
  NAND2_X1 U4845 ( .A1(n4298), .A2(n4201), .ZN(n4160) );
  INV_X1 U4846 ( .A(n4175), .ZN(n4150) );
  OAI21_X1 U4847 ( .B1(n4150), .B2(n4149), .A(n4148), .ZN(n4361) );
  INV_X1 U4848 ( .A(n4361), .ZN(n4158) );
  AOI22_X1 U4849 ( .A1(n4152), .A2(n4292), .B1(n4151), .B2(n4293), .ZN(n4155)
         );
  AOI22_X1 U4850 ( .A1(n4566), .A2(REG2_REG_20__SCAN_IN), .B1(n4153), .B2(
        n4557), .ZN(n4154) );
  OAI211_X1 U4851 ( .C1(n4296), .C2(n4156), .A(n4155), .B(n4154), .ZN(n4157)
         );
  AOI21_X1 U4852 ( .B1(n4158), .B2(n4560), .A(n4157), .ZN(n4159) );
  OAI211_X1 U4853 ( .C1(n4204), .C2(n4295), .A(n4160), .B(n4159), .ZN(U3270)
         );
  XOR2_X1 U4854 ( .A(n4168), .B(n4161), .Z(n4302) );
  INV_X1 U4855 ( .A(n4302), .ZN(n4181) );
  INV_X1 U4856 ( .A(n4162), .ZN(n4163) );
  NOR2_X1 U4857 ( .A1(n4164), .A2(n4163), .ZN(n4183) );
  INV_X1 U4858 ( .A(n4165), .ZN(n4166) );
  AOI21_X1 U4859 ( .B1(n4183), .B2(n4167), .A(n4166), .ZN(n4169) );
  XNOR2_X1 U4860 ( .A(n4169), .B(n4168), .ZN(n4174) );
  OAI22_X1 U4861 ( .A1(n4170), .A2(n4594), .B1(n4593), .B2(n4176), .ZN(n4171)
         );
  AOI21_X1 U4862 ( .B1(n4637), .B2(n4172), .A(n4171), .ZN(n4173) );
  OAI21_X1 U4863 ( .B1(n4174), .B2(n4213), .A(n4173), .ZN(n4301) );
  OAI21_X1 U4864 ( .B1(n4195), .B2(n4176), .A(n4175), .ZN(n4365) );
  AOI22_X1 U4865 ( .A1(n4566), .A2(REG2_REG_19__SCAN_IN), .B1(n4177), .B2(
        n4557), .ZN(n4178) );
  OAI21_X1 U4866 ( .B1(n4365), .B2(n4220), .A(n4178), .ZN(n4179) );
  AOI21_X1 U4867 ( .B1(n4301), .B2(n4402), .A(n4179), .ZN(n4180) );
  OAI21_X1 U4868 ( .B1(n4181), .B2(n4223), .A(n4180), .ZN(U3271) );
  XNOR2_X1 U4869 ( .A(n4183), .B(n4182), .ZN(n4190) );
  AOI22_X1 U4870 ( .A1(n4185), .A2(n4635), .B1(n4634), .B2(n4184), .ZN(n4186)
         );
  OAI21_X1 U4871 ( .B1(n4187), .B2(n4327), .A(n4186), .ZN(n4188) );
  AOI21_X1 U4872 ( .B1(n4190), .B2(n4189), .A(n4188), .ZN(n4306) );
  AOI21_X1 U4873 ( .B1(n4193), .B2(n4192), .A(n4191), .ZN(n4307) );
  INV_X1 U4874 ( .A(n4307), .ZN(n4202) );
  OAI21_X1 U4875 ( .B1(n4216), .B2(n4194), .A(n4314), .ZN(n4196) );
  OR2_X1 U4876 ( .A1(n4196), .A2(n4195), .ZN(n4305) );
  AOI22_X1 U4877 ( .A1(n4566), .A2(REG2_REG_18__SCAN_IN), .B1(n4197), .B2(
        n4557), .ZN(n4198) );
  OAI21_X1 U4878 ( .B1(n4305), .B2(n4199), .A(n4198), .ZN(n4200) );
  AOI21_X1 U4879 ( .B1(n4202), .B2(n4201), .A(n4200), .ZN(n4203) );
  OAI21_X1 U4880 ( .B1(n4204), .B2(n4306), .A(n4203), .ZN(U3272) );
  XNOR2_X1 U4881 ( .A(n4205), .B(n4207), .ZN(n4309) );
  INV_X1 U4882 ( .A(n4309), .ZN(n4224) );
  XOR2_X1 U4883 ( .A(n4207), .B(n4206), .Z(n4214) );
  OAI22_X1 U4884 ( .A1(n4209), .A2(n4594), .B1(n4208), .B2(n4593), .ZN(n4210)
         );
  AOI21_X1 U4885 ( .B1(n4637), .B2(n4211), .A(n4210), .ZN(n4212) );
  OAI21_X1 U4886 ( .B1(n4214), .B2(n4213), .A(n4212), .ZN(n4308) );
  AND2_X1 U4887 ( .A1(n4315), .A2(n4215), .ZN(n4217) );
  OR2_X1 U4888 ( .A1(n4217), .A2(n4216), .ZN(n4370) );
  AOI22_X1 U4889 ( .A1(n4566), .A2(REG2_REG_17__SCAN_IN), .B1(n4218), .B2(
        n4557), .ZN(n4219) );
  OAI21_X1 U4890 ( .B1(n4370), .B2(n4220), .A(n4219), .ZN(n4221) );
  AOI21_X1 U4891 ( .B1(n4308), .B2(n4402), .A(n4221), .ZN(n4222) );
  OAI21_X1 U4892 ( .B1(n4224), .B2(n4223), .A(n4222), .ZN(U3273) );
  INV_X1 U4893 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4950) );
  INV_X1 U4894 ( .A(n4234), .ZN(n4237) );
  NAND2_X1 U4895 ( .A1(n4230), .A2(n4237), .ZN(n4231) );
  XNOR2_X1 U4896 ( .A(n4231), .B(n4227), .ZN(n4399) );
  NAND2_X1 U4897 ( .A1(n4399), .A2(n4235), .ZN(n4229) );
  OR2_X1 U4898 ( .A1(n4226), .A2(n4225), .ZN(n4236) );
  OAI21_X1 U4899 ( .B1(n4227), .B2(n4593), .A(n4236), .ZN(n4398) );
  NAND2_X1 U4900 ( .A1(n4398), .A2(n4666), .ZN(n4228) );
  OAI211_X1 U4901 ( .C1(n4666), .C2(n4950), .A(n4229), .B(n4228), .ZN(U3549)
         );
  INV_X1 U4902 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4886) );
  INV_X1 U4903 ( .A(n4230), .ZN(n4233) );
  INV_X1 U4904 ( .A(n4231), .ZN(n4232) );
  NAND2_X1 U4905 ( .A1(n4403), .A2(n4235), .ZN(n4239) );
  OAI21_X1 U4906 ( .B1(n4237), .B2(n4593), .A(n4236), .ZN(n4401) );
  NAND2_X1 U4907 ( .A1(n4401), .A2(n4666), .ZN(n4238) );
  OAI211_X1 U4908 ( .C1(n4666), .C2(n4886), .A(n4239), .B(n4238), .ZN(U3548)
         );
  NAND2_X1 U4909 ( .A1(n4240), .A2(n4646), .ZN(n4246) );
  OAI22_X1 U4910 ( .A1(n4247), .A2(n4327), .B1(n4593), .B2(n4241), .ZN(n4243)
         );
  NAND2_X1 U4911 ( .A1(n4246), .A2(n4245), .ZN(n4339) );
  MUX2_X1 U4912 ( .A(REG1_REG_29__SCAN_IN), .B(n4339), .S(n4666), .Z(U3547) );
  OAI22_X1 U4913 ( .A1(n4247), .A2(n4594), .B1(n2850), .B2(n4593), .ZN(n4250)
         );
  NOR2_X1 U4914 ( .A1(n4248), .A2(n4641), .ZN(n4249) );
  AOI211_X1 U4915 ( .C1(n4637), .C2(n4251), .A(n4250), .B(n4249), .ZN(n4253)
         );
  OAI211_X1 U4916 ( .C1(n4254), .C2(n4590), .A(n4253), .B(n4252), .ZN(n4340)
         );
  MUX2_X1 U4917 ( .A(REG1_REG_27__SCAN_IN), .B(n4340), .S(n4666), .Z(U3545) );
  INV_X1 U4918 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4261) );
  AOI22_X1 U4919 ( .A1(n4273), .A2(n4637), .B1(n4255), .B2(n4634), .ZN(n4256)
         );
  OAI211_X1 U4920 ( .C1(n4258), .C2(n4594), .A(n4257), .B(n4256), .ZN(n4259)
         );
  AOI21_X1 U4921 ( .B1(n4260), .B2(n4646), .A(n4259), .ZN(n4341) );
  MUX2_X1 U4922 ( .A(n4261), .B(n4341), .S(n4666), .Z(n4262) );
  OAI21_X1 U4923 ( .B1(n4333), .B2(n4343), .A(n4262), .ZN(U3544) );
  AOI22_X1 U4924 ( .A1(n4264), .A2(n4637), .B1(n4263), .B2(n4634), .ZN(n4265)
         );
  OAI21_X1 U4925 ( .B1(n4266), .B2(n4594), .A(n4265), .ZN(n4267) );
  AOI21_X1 U4926 ( .B1(n4268), .B2(n4314), .A(n4267), .ZN(n4270) );
  OAI211_X1 U4927 ( .C1(n4271), .C2(n4590), .A(n4270), .B(n4269), .ZN(n4344)
         );
  MUX2_X1 U4928 ( .A(REG1_REG_25__SCAN_IN), .B(n4344), .S(n4666), .Z(U3543) );
  INV_X1 U4929 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4993) );
  AOI22_X1 U4930 ( .A1(n4273), .A2(n4635), .B1(n4634), .B2(n4272), .ZN(n4274)
         );
  OAI211_X1 U4931 ( .C1(n4276), .C2(n4327), .A(n4275), .B(n4274), .ZN(n4277)
         );
  AOI21_X1 U4932 ( .B1(n4278), .B2(n4646), .A(n4277), .ZN(n4345) );
  MUX2_X1 U4933 ( .A(n4993), .B(n4345), .S(n4666), .Z(n4279) );
  OAI21_X1 U4934 ( .B1(n4333), .B2(n4348), .A(n4279), .ZN(U3542) );
  INV_X1 U4935 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4282) );
  AOI21_X1 U4936 ( .B1(n4281), .B2(n4646), .A(n4280), .ZN(n4349) );
  MUX2_X1 U4937 ( .A(n4282), .B(n4349), .S(n4666), .Z(n4283) );
  OAI21_X1 U4938 ( .B1(n4333), .B2(n4352), .A(n4283), .ZN(U3541) );
  NAND3_X1 U4939 ( .A1(n4285), .A2(n4314), .A3(n4284), .ZN(n4286) );
  OAI211_X1 U4940 ( .C1(n4288), .C2(n4590), .A(n4287), .B(n4286), .ZN(n4353)
         );
  MUX2_X1 U4941 ( .A(REG1_REG_22__SCAN_IN), .B(n4353), .S(n4666), .Z(U3540) );
  INV_X1 U4942 ( .A(REG1_REG_21__SCAN_IN), .ZN(n5042) );
  AOI21_X1 U4943 ( .B1(n4290), .B2(n4646), .A(n4289), .ZN(n4354) );
  MUX2_X1 U4944 ( .A(n5042), .B(n4354), .S(n4666), .Z(n4291) );
  OAI21_X1 U4945 ( .B1(n4333), .B2(n4357), .A(n4291), .ZN(U3539) );
  INV_X1 U4946 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4299) );
  AOI22_X1 U4947 ( .A1(n4293), .A2(n4635), .B1(n4634), .B2(n4292), .ZN(n4294)
         );
  OAI211_X1 U4948 ( .C1(n4296), .C2(n4327), .A(n4295), .B(n4294), .ZN(n4297)
         );
  AOI21_X1 U4949 ( .B1(n4298), .B2(n4646), .A(n4297), .ZN(n4358) );
  MUX2_X1 U4950 ( .A(n4299), .B(n4358), .S(n4666), .Z(n4300) );
  OAI21_X1 U4951 ( .B1(n4333), .B2(n4361), .A(n4300), .ZN(U3538) );
  INV_X1 U4952 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4303) );
  AOI21_X1 U4953 ( .B1(n4302), .B2(n4646), .A(n4301), .ZN(n4362) );
  MUX2_X1 U4954 ( .A(n4303), .B(n4362), .S(n4666), .Z(n4304) );
  OAI21_X1 U4955 ( .B1(n4333), .B2(n4365), .A(n4304), .ZN(U3537) );
  OAI211_X1 U4956 ( .C1(n4307), .C2(n4590), .A(n4306), .B(n4305), .ZN(n4366)
         );
  MUX2_X1 U4957 ( .A(REG1_REG_18__SCAN_IN), .B(n4366), .S(n4666), .Z(U3536) );
  AOI21_X1 U4958 ( .B1(n4309), .B2(n4646), .A(n4308), .ZN(n4367) );
  MUX2_X1 U4959 ( .A(n4310), .B(n4367), .S(n4666), .Z(n4311) );
  OAI21_X1 U4960 ( .B1(n4333), .B2(n4370), .A(n4311), .ZN(U3535) );
  INV_X1 U4961 ( .A(n4312), .ZN(n4318) );
  NAND3_X1 U4962 ( .A1(n4315), .A2(n4314), .A3(n4313), .ZN(n4316) );
  OAI211_X1 U4963 ( .C1(n4318), .C2(n4590), .A(n4317), .B(n4316), .ZN(n4371)
         );
  MUX2_X1 U4964 ( .A(REG1_REG_16__SCAN_IN), .B(n4371), .S(n4666), .Z(U3534) );
  INV_X1 U4965 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4321) );
  AOI21_X1 U4966 ( .B1(n4320), .B2(n4646), .A(n4319), .ZN(n4372) );
  MUX2_X1 U4967 ( .A(n4321), .B(n4372), .S(n4666), .Z(n4322) );
  OAI21_X1 U4968 ( .B1(n4333), .B2(n4375), .A(n4322), .ZN(U3533) );
  INV_X1 U4969 ( .A(n4323), .ZN(n4331) );
  AOI22_X1 U4970 ( .A1(n4325), .A2(n4635), .B1(n4634), .B2(n4324), .ZN(n4326)
         );
  OAI21_X1 U4971 ( .B1(n4328), .B2(n4327), .A(n4326), .ZN(n4330) );
  AOI211_X1 U4972 ( .C1(n4617), .C2(n4331), .A(n4330), .B(n4329), .ZN(n4376)
         );
  MUX2_X1 U4973 ( .A(n4533), .B(n4376), .S(n4666), .Z(n4332) );
  OAI21_X1 U4974 ( .B1(n4333), .B2(n4379), .A(n4332), .ZN(U3532) );
  INV_X1 U4975 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4992) );
  NAND2_X1 U4976 ( .A1(n4399), .A2(n4336), .ZN(n4335) );
  NAND2_X1 U4977 ( .A1(n4398), .A2(n4649), .ZN(n4334) );
  OAI211_X1 U4978 ( .C1(n4649), .C2(n4992), .A(n4335), .B(n4334), .ZN(U3517)
         );
  INV_X1 U4979 ( .A(REG0_REG_30__SCAN_IN), .ZN(n5011) );
  NAND2_X1 U4980 ( .A1(n4403), .A2(n4336), .ZN(n4338) );
  NAND2_X1 U4981 ( .A1(n4401), .A2(n4649), .ZN(n4337) );
  OAI211_X1 U4982 ( .C1(n4649), .C2(n5011), .A(n4338), .B(n4337), .ZN(U3516)
         );
  MUX2_X1 U4983 ( .A(REG0_REG_29__SCAN_IN), .B(n4339), .S(n4649), .Z(U3515) );
  MUX2_X1 U4984 ( .A(REG0_REG_27__SCAN_IN), .B(n4340), .S(n4649), .Z(U3513) );
  INV_X1 U4985 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4862) );
  MUX2_X1 U4986 ( .A(n4862), .B(n4341), .S(n4649), .Z(n4342) );
  OAI21_X1 U4987 ( .B1(n4343), .B2(n4378), .A(n4342), .ZN(U3512) );
  MUX2_X1 U4988 ( .A(REG0_REG_25__SCAN_IN), .B(n4344), .S(n4649), .Z(U3511) );
  INV_X1 U4989 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4346) );
  MUX2_X1 U4990 ( .A(n4346), .B(n4345), .S(n4649), .Z(n4347) );
  OAI21_X1 U4991 ( .B1(n4348), .B2(n4378), .A(n4347), .ZN(U3510) );
  INV_X1 U4992 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4350) );
  MUX2_X1 U4993 ( .A(n4350), .B(n4349), .S(n4649), .Z(n4351) );
  OAI21_X1 U4994 ( .B1(n4352), .B2(n4378), .A(n4351), .ZN(U3509) );
  MUX2_X1 U4995 ( .A(REG0_REG_22__SCAN_IN), .B(n4353), .S(n4649), .Z(U3508) );
  INV_X1 U4996 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4355) );
  MUX2_X1 U4997 ( .A(n4355), .B(n4354), .S(n4649), .Z(n4356) );
  OAI21_X1 U4998 ( .B1(n4357), .B2(n4378), .A(n4356), .ZN(U3507) );
  INV_X1 U4999 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4359) );
  MUX2_X1 U5000 ( .A(n4359), .B(n4358), .S(n4649), .Z(n4360) );
  OAI21_X1 U5001 ( .B1(n4361), .B2(n4378), .A(n4360), .ZN(U3506) );
  INV_X1 U5002 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4363) );
  MUX2_X1 U5003 ( .A(n4363), .B(n4362), .S(n4649), .Z(n4364) );
  OAI21_X1 U5004 ( .B1(n4365), .B2(n4378), .A(n4364), .ZN(U3505) );
  MUX2_X1 U5005 ( .A(REG0_REG_18__SCAN_IN), .B(n4366), .S(n4649), .Z(U3503) );
  INV_X1 U5006 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4368) );
  MUX2_X1 U5007 ( .A(n4368), .B(n4367), .S(n4649), .Z(n4369) );
  OAI21_X1 U5008 ( .B1(n4370), .B2(n4378), .A(n4369), .ZN(U3501) );
  MUX2_X1 U5009 ( .A(REG0_REG_16__SCAN_IN), .B(n4371), .S(n4649), .Z(U3499) );
  INV_X1 U5010 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4373) );
  MUX2_X1 U5011 ( .A(n4373), .B(n4372), .S(n4649), .Z(n4374) );
  OAI21_X1 U5012 ( .B1(n4375), .B2(n4378), .A(n4374), .ZN(U3497) );
  INV_X1 U5013 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4863) );
  MUX2_X1 U5014 ( .A(n4863), .B(n4376), .S(n4649), .Z(n4377) );
  OAI21_X1 U5015 ( .B1(n4379), .B2(n4378), .A(n4377), .ZN(U3495) );
  MUX2_X1 U5016 ( .A(n2648), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U5017 ( .A(n2905), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5018 ( .A(n4380), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U5019 ( .A(n4381), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5020 ( .A(DATAI_18_), .B(n4382), .S(STATE_REG_SCAN_IN), .Z(U3334)
         );
  MUX2_X1 U5021 ( .A(DATAI_16_), .B(n4383), .S(STATE_REG_SCAN_IN), .Z(U3336)
         );
  MUX2_X1 U5022 ( .A(DATAI_9_), .B(n4384), .S(STATE_REG_SCAN_IN), .Z(U3343) );
  MUX2_X1 U5023 ( .A(n4457), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  INV_X1 U5024 ( .A(DATAI_2_), .ZN(n4385) );
  AOI22_X1 U5025 ( .A1(STATE_REG_SCAN_IN), .A2(n4434), .B1(n4385), .B2(U3149), 
        .ZN(U3350) );
  INV_X1 U5026 ( .A(DATAI_3_), .ZN(n4833) );
  AOI22_X1 U5027 ( .A1(STATE_REG_SCAN_IN), .A2(n2346), .B1(n4833), .B2(U3149), 
        .ZN(U3349) );
  OAI22_X1 U5028 ( .A1(U3149), .A2(n4386), .B1(DATAI_4_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4387) );
  INV_X1 U5029 ( .A(n4387), .ZN(U3348) );
  AOI21_X1 U5030 ( .B1(n4543), .B2(ADDR_REG_3__SCAN_IN), .A(n4388), .ZN(n4397)
         );
  NAND2_X1 U5031 ( .A1(n4389), .A2(n4538), .ZN(n4396) );
  OAI211_X1 U5032 ( .C1(REG1_REG_3__SCAN_IN), .C2(n4391), .A(n4553), .B(n4390), 
        .ZN(n4395) );
  OAI211_X1 U5033 ( .C1(REG2_REG_3__SCAN_IN), .C2(n4393), .A(n4551), .B(n4392), 
        .ZN(n4394) );
  NAND4_X1 U5034 ( .A1(n4397), .A2(n4396), .A3(n4395), .A4(n4394), .ZN(U3243)
         );
  INV_X1 U5035 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4892) );
  AOI22_X1 U5036 ( .A1(n4399), .A2(n4560), .B1(n4402), .B2(n4398), .ZN(n4400)
         );
  OAI21_X1 U5037 ( .B1(n4402), .B2(n4892), .A(n4400), .ZN(U3260) );
  INV_X1 U5038 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4891) );
  AOI22_X1 U5039 ( .A1(n4403), .A2(n4560), .B1(n4402), .B2(n4401), .ZN(n4404)
         );
  OAI21_X1 U5040 ( .B1(n4891), .B2(n4402), .A(n4404), .ZN(U3261) );
  NOR2_X1 U5041 ( .A1(n4406), .A2(REG2_REG_0__SCAN_IN), .ZN(n4407) );
  NOR2_X1 U5042 ( .A1(n4415), .A2(n4407), .ZN(n4423) );
  OAI21_X1 U5043 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4416), .A(n4423), .ZN(n4408)
         );
  XNOR2_X1 U5044 ( .A(n4408), .B(n2335), .ZN(n4411) );
  AOI22_X1 U5045 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4543), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4409) );
  OAI21_X1 U5046 ( .B1(n4411), .B2(n4410), .A(n4409), .ZN(U3240) );
  AOI22_X1 U5047 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4543), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4428) );
  AOI21_X1 U5048 ( .B1(n4414), .B2(n4413), .A(n4412), .ZN(n4668) );
  OR3_X1 U5049 ( .A1(n4668), .A2(n4416), .A3(n4415), .ZN(n4422) );
  INV_X1 U5050 ( .A(n4417), .ZN(n4420) );
  AOI21_X1 U5051 ( .B1(n4420), .B2(n4419), .A(n4418), .ZN(n4421) );
  OAI211_X1 U5052 ( .C1(IR_REG_0__SCAN_IN), .C2(n4423), .A(n4422), .B(n4421), 
        .ZN(n4444) );
  OAI211_X1 U5053 ( .C1(n4426), .C2(n4425), .A(n4553), .B(n4424), .ZN(n4427)
         );
  AND3_X1 U5054 ( .A1(n4428), .A2(n4444), .A3(n4427), .ZN(n4433) );
  OAI211_X1 U5055 ( .C1(n4431), .C2(n4430), .A(n4551), .B(n4429), .ZN(n4432)
         );
  OAI211_X1 U5056 ( .C1(n4556), .C2(n4434), .A(n4433), .B(n4432), .ZN(U3242)
         );
  OAI211_X1 U5057 ( .C1(REG2_REG_4__SCAN_IN), .C2(n4436), .A(n4551), .B(n4435), 
        .ZN(n4440) );
  OAI211_X1 U5058 ( .C1(REG1_REG_4__SCAN_IN), .C2(n4438), .A(n4553), .B(n4437), 
        .ZN(n4439) );
  OAI211_X1 U5059 ( .C1(n4556), .C2(n4441), .A(n4440), .B(n4439), .ZN(n4442)
         );
  AOI211_X1 U5060 ( .C1(n4543), .C2(ADDR_REG_4__SCAN_IN), .A(n4443), .B(n4442), 
        .ZN(n4445) );
  NAND2_X1 U5061 ( .A1(n4445), .A2(n4444), .ZN(U3244) );
  OAI211_X1 U5062 ( .C1(n4448), .C2(n4447), .A(n4553), .B(n4446), .ZN(n4453)
         );
  OAI211_X1 U5063 ( .C1(n4451), .C2(n4450), .A(n4551), .B(n4449), .ZN(n4452)
         );
  OAI211_X1 U5064 ( .C1(n4556), .C2(n4583), .A(n4453), .B(n4452), .ZN(n4454)
         );
  AOI211_X1 U5065 ( .C1(n4543), .C2(ADDR_REG_5__SCAN_IN), .A(n4455), .B(n4454), 
        .ZN(n4456) );
  INV_X1 U5066 ( .A(n4456), .ZN(U3245) );
  AOI22_X1 U5067 ( .A1(ADDR_REG_6__SCAN_IN), .A2(n4543), .B1(
        REG3_REG_6__SCAN_IN), .B2(U3149), .ZN(n4465) );
  NAND2_X1 U5068 ( .A1(n4538), .A2(n4457), .ZN(n4464) );
  OAI211_X1 U5069 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4459), .A(n4553), .B(n4458), 
        .ZN(n4463) );
  OAI211_X1 U5070 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4461), .A(n4551), .B(n4460), 
        .ZN(n4462) );
  NAND4_X1 U5071 ( .A1(n4465), .A2(n4464), .A3(n4463), .A4(n4462), .ZN(U3246)
         );
  AOI22_X1 U5072 ( .A1(REG1_REG_7__SCAN_IN), .A2(n4581), .B1(n4476), .B2(n2314), .ZN(n4468) );
  OAI21_X1 U5073 ( .B1(n4468), .B2(n4467), .A(n4553), .ZN(n4466) );
  AOI21_X1 U5074 ( .B1(n4468), .B2(n4467), .A(n4466), .ZN(n4470) );
  AOI211_X1 U5075 ( .C1(n4543), .C2(ADDR_REG_7__SCAN_IN), .A(n4470), .B(n4469), 
        .ZN(n4475) );
  OAI211_X1 U5076 ( .C1(n4473), .C2(n4472), .A(n4551), .B(n4471), .ZN(n4474)
         );
  OAI211_X1 U5077 ( .C1(n4556), .C2(n4476), .A(n4475), .B(n4474), .ZN(U3247)
         );
  AOI211_X1 U5078 ( .C1(n4479), .C2(n4478), .A(n4477), .B(n4531), .ZN(n4480)
         );
  AOI211_X1 U5079 ( .C1(n4543), .C2(ADDR_REG_8__SCAN_IN), .A(n4481), .B(n4480), 
        .ZN(n4485) );
  OAI211_X1 U5080 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4483), .A(n4551), .B(n4482), 
        .ZN(n4484) );
  OAI211_X1 U5081 ( .C1(n4556), .C2(n4580), .A(n4485), .B(n4484), .ZN(U3248)
         );
  AOI211_X1 U5082 ( .C1(n4488), .C2(n4487), .A(n4486), .B(n4531), .ZN(n4490)
         );
  AOI211_X1 U5083 ( .C1(n4543), .C2(ADDR_REG_10__SCAN_IN), .A(n4490), .B(n4489), .ZN(n4494) );
  OAI211_X1 U5084 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4492), .A(n4551), .B(n4491), .ZN(n4493) );
  OAI211_X1 U5085 ( .C1(n4556), .C2(n4579), .A(n4494), .B(n4493), .ZN(U3250)
         );
  AOI211_X1 U5086 ( .C1(n4497), .C2(n4496), .A(n4495), .B(n4531), .ZN(n4499)
         );
  AOI211_X1 U5087 ( .C1(n4543), .C2(ADDR_REG_11__SCAN_IN), .A(n4499), .B(n4498), .ZN(n4504) );
  OAI211_X1 U5088 ( .C1(n4502), .C2(n4501), .A(n4551), .B(n4500), .ZN(n4503)
         );
  OAI211_X1 U5089 ( .C1(n4556), .C2(n4577), .A(n4504), .B(n4503), .ZN(U3251)
         );
  AOI211_X1 U5090 ( .C1(n4507), .C2(n4506), .A(n4505), .B(n4531), .ZN(n4510)
         );
  INV_X1 U5091 ( .A(n4508), .ZN(n4509) );
  AOI211_X1 U5092 ( .C1(n4543), .C2(ADDR_REG_12__SCAN_IN), .A(n4510), .B(n4509), .ZN(n4514) );
  OAI211_X1 U5093 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4512), .A(n4551), .B(n4511), .ZN(n4513) );
  OAI211_X1 U5094 ( .C1(n4556), .C2(n2347), .A(n4514), .B(n4513), .ZN(U3252)
         );
  INV_X1 U5095 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n5008) );
  AOI21_X1 U5096 ( .B1(n4978), .B2(n4575), .A(n4515), .ZN(n4518) );
  OAI21_X1 U5097 ( .B1(n4518), .B2(n4517), .A(n4551), .ZN(n4516) );
  AOI21_X1 U5098 ( .B1(n4518), .B2(n4517), .A(n4516), .ZN(n4523) );
  AOI211_X1 U5099 ( .C1(n4521), .C2(n4520), .A(n4519), .B(n4531), .ZN(n4522)
         );
  AOI211_X1 U5100 ( .C1(n4538), .C2(n4524), .A(n4523), .B(n4522), .ZN(n4526)
         );
  OAI211_X1 U5101 ( .C1(n4527), .C2(n5008), .A(n4526), .B(n4525), .ZN(U3253)
         );
  NAND2_X1 U5102 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4543), .ZN(n4541) );
  AOI211_X1 U5103 ( .C1(n4530), .C2(n4529), .A(n2286), .B(n4528), .ZN(n4536)
         );
  AOI211_X1 U5104 ( .C1(n4534), .C2(n4533), .A(n4532), .B(n4531), .ZN(n4535)
         );
  AOI211_X1 U5105 ( .C1(n4538), .C2(n4537), .A(n4536), .B(n4535), .ZN(n4540)
         );
  NAND3_X1 U5106 ( .A1(n4541), .A2(n4540), .A3(n4539), .ZN(U3254) );
  AOI21_X1 U5107 ( .B1(n4543), .B2(ADDR_REG_17__SCAN_IN), .A(n4542), .ZN(n4555) );
  OAI21_X1 U5108 ( .B1(n4546), .B2(n4545), .A(n4544), .ZN(n4552) );
  OAI21_X1 U5109 ( .B1(n4549), .B2(n4548), .A(n4547), .ZN(n4550) );
  AOI22_X1 U5110 ( .A1(n4553), .A2(n4552), .B1(n4551), .B2(n4550), .ZN(n4554)
         );
  OAI211_X1 U5111 ( .C1(n4574), .C2(n4556), .A(n4555), .B(n4554), .ZN(U3257)
         );
  AOI22_X1 U5112 ( .A1(n4558), .A2(n4557), .B1(REG2_REG_6__SCAN_IN), .B2(n4566), .ZN(n4564) );
  AOI22_X1 U5113 ( .A1(n4562), .A2(n4561), .B1(n4560), .B2(n4559), .ZN(n4563)
         );
  OAI211_X1 U5114 ( .C1(n4566), .C2(n4565), .A(n4564), .B(n4563), .ZN(U3284)
         );
  INV_X1 U5115 ( .A(D_REG_31__SCAN_IN), .ZN(n4965) );
  NOR2_X1 U5116 ( .A1(n4571), .A2(n4965), .ZN(U3291) );
  AND2_X1 U5117 ( .A1(D_REG_30__SCAN_IN), .A2(n4570), .ZN(U3292) );
  AND2_X1 U5118 ( .A1(D_REG_29__SCAN_IN), .A2(n4570), .ZN(U3293) );
  AND2_X1 U5119 ( .A1(D_REG_28__SCAN_IN), .A2(n4570), .ZN(U3294) );
  AND2_X1 U5120 ( .A1(D_REG_27__SCAN_IN), .A2(n4570), .ZN(U3295) );
  AND2_X1 U5121 ( .A1(n4570), .A2(D_REG_26__SCAN_IN), .ZN(U3296) );
  AND2_X1 U5122 ( .A1(D_REG_25__SCAN_IN), .A2(n4570), .ZN(U3297) );
  AND2_X1 U5123 ( .A1(D_REG_24__SCAN_IN), .A2(n4570), .ZN(U3298) );
  INV_X1 U5124 ( .A(D_REG_23__SCAN_IN), .ZN(n5028) );
  NOR2_X1 U5125 ( .A1(n4571), .A2(n5028), .ZN(U3299) );
  AND2_X1 U5126 ( .A1(D_REG_22__SCAN_IN), .A2(n4570), .ZN(U3300) );
  AND2_X1 U5127 ( .A1(D_REG_21__SCAN_IN), .A2(n4570), .ZN(U3301) );
  AND2_X1 U5128 ( .A1(D_REG_20__SCAN_IN), .A2(n4570), .ZN(U3302) );
  NOR2_X1 U5129 ( .A1(n4571), .A2(n4856), .ZN(U3303) );
  INV_X1 U5130 ( .A(D_REG_18__SCAN_IN), .ZN(n4857) );
  NOR2_X1 U5131 ( .A1(n4571), .A2(n4857), .ZN(U3304) );
  NOR2_X1 U5132 ( .A1(n4571), .A2(n4567), .ZN(U3305) );
  AND2_X1 U5133 ( .A1(D_REG_16__SCAN_IN), .A2(n4570), .ZN(U3306) );
  NOR2_X1 U5134 ( .A1(n4571), .A2(n4568), .ZN(U3307) );
  NOR2_X1 U5135 ( .A1(n4571), .A2(n4569), .ZN(U3308) );
  AND2_X1 U5136 ( .A1(D_REG_13__SCAN_IN), .A2(n4570), .ZN(U3309) );
  AND2_X1 U5137 ( .A1(D_REG_12__SCAN_IN), .A2(n4570), .ZN(U3310) );
  AND2_X1 U5138 ( .A1(n4570), .A2(D_REG_11__SCAN_IN), .ZN(U3311) );
  INV_X1 U5139 ( .A(D_REG_10__SCAN_IN), .ZN(n5018) );
  NOR2_X1 U5140 ( .A1(n4571), .A2(n5018), .ZN(U3312) );
  INV_X1 U5141 ( .A(D_REG_9__SCAN_IN), .ZN(n4972) );
  NOR2_X1 U5142 ( .A1(n4571), .A2(n4972), .ZN(U3313) );
  INV_X1 U5143 ( .A(D_REG_8__SCAN_IN), .ZN(n5030) );
  NOR2_X1 U5144 ( .A1(n4571), .A2(n5030), .ZN(U3314) );
  AND2_X1 U5145 ( .A1(D_REG_7__SCAN_IN), .A2(n4570), .ZN(U3315) );
  AND2_X1 U5146 ( .A1(D_REG_6__SCAN_IN), .A2(n4570), .ZN(U3316) );
  AND2_X1 U5147 ( .A1(n4570), .A2(D_REG_5__SCAN_IN), .ZN(U3317) );
  AND2_X1 U5148 ( .A1(D_REG_4__SCAN_IN), .A2(n4570), .ZN(U3318) );
  INV_X1 U5149 ( .A(D_REG_3__SCAN_IN), .ZN(n5027) );
  NOR2_X1 U5150 ( .A1(n4571), .A2(n5027), .ZN(U3319) );
  INV_X1 U5151 ( .A(D_REG_2__SCAN_IN), .ZN(n5015) );
  NOR2_X1 U5152 ( .A1(n4571), .A2(n5015), .ZN(U3320) );
  INV_X1 U5153 ( .A(DATAI_23_), .ZN(n4573) );
  AOI21_X1 U5154 ( .B1(U3149), .B2(n4573), .A(n4572), .ZN(U3329) );
  INV_X1 U5155 ( .A(DATAI_17_), .ZN(n4999) );
  AOI22_X1 U5156 ( .A1(STATE_REG_SCAN_IN), .A2(n4574), .B1(n4999), .B2(U3149), 
        .ZN(U3335) );
  AOI22_X1 U5157 ( .A1(STATE_REG_SCAN_IN), .A2(n4575), .B1(n2763), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5158 ( .A(DATAI_12_), .ZN(n4946) );
  AOI22_X1 U5159 ( .A1(STATE_REG_SCAN_IN), .A2(n2347), .B1(n4946), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5160 ( .A(DATAI_11_), .ZN(n4576) );
  AOI22_X1 U5161 ( .A1(STATE_REG_SCAN_IN), .A2(n4577), .B1(n4576), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5162 ( .A(DATAI_10_), .ZN(n4578) );
  AOI22_X1 U5163 ( .A1(STATE_REG_SCAN_IN), .A2(n4579), .B1(n4578), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5164 ( .A(DATAI_8_), .ZN(n4826) );
  AOI22_X1 U5165 ( .A1(STATE_REG_SCAN_IN), .A2(n4580), .B1(n4826), .B2(U3149), 
        .ZN(U3344) );
  OAI22_X1 U5166 ( .A1(U3149), .A2(n4581), .B1(DATAI_7_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4582) );
  INV_X1 U5167 ( .A(n4582), .ZN(U3345) );
  INV_X1 U5168 ( .A(DATAI_5_), .ZN(n5014) );
  AOI22_X1 U5169 ( .A1(STATE_REG_SCAN_IN), .A2(n4583), .B1(n5014), .B2(U3149), 
        .ZN(U3347) );
  AOI22_X1 U5170 ( .A1(STATE_REG_SCAN_IN), .A2(n2335), .B1(n2334), .B2(U3149), 
        .ZN(U3352) );
  NOR2_X1 U5171 ( .A1(n4585), .A2(n4584), .ZN(n4587) );
  AOI211_X1 U5172 ( .C1(n4646), .C2(n4588), .A(n4587), .B(n4586), .ZN(n4651)
         );
  INV_X1 U5173 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4589) );
  AOI22_X1 U5174 ( .A1(n4649), .A2(n4651), .B1(n4589), .B2(n4647), .ZN(U3467)
         );
  NOR2_X1 U5175 ( .A1(n4591), .A2(n4590), .ZN(n4599) );
  OAI22_X1 U5176 ( .A1(n2680), .A2(n4594), .B1(n4593), .B2(n4592), .ZN(n4598)
         );
  NAND2_X1 U5177 ( .A1(n2971), .A2(n4637), .ZN(n4595) );
  OAI21_X1 U5178 ( .B1(n4596), .B2(n4641), .A(n4595), .ZN(n4597) );
  NOR4_X1 U5179 ( .A1(n4600), .A2(n4599), .A3(n4598), .A4(n4597), .ZN(n4653)
         );
  INV_X1 U5180 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4601) );
  AOI22_X1 U5181 ( .A1(n4649), .A2(n4653), .B1(n4601), .B2(n4647), .ZN(U3469)
         );
  NOR3_X1 U5182 ( .A1(n4603), .A2(n4602), .A3(n4641), .ZN(n4605) );
  AOI211_X1 U5183 ( .C1(n4617), .C2(n4606), .A(n4605), .B(n4604), .ZN(n4654)
         );
  INV_X1 U5184 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4607) );
  AOI22_X1 U5185 ( .A1(n4649), .A2(n4654), .B1(n4607), .B2(n4647), .ZN(U3471)
         );
  OAI22_X1 U5186 ( .A1(n4610), .A2(n4609), .B1(n4641), .B2(n4608), .ZN(n4611)
         );
  NOR2_X1 U5187 ( .A1(n4612), .A2(n4611), .ZN(n4656) );
  INV_X1 U5188 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4613) );
  AOI22_X1 U5189 ( .A1(n4649), .A2(n4656), .B1(n4613), .B2(n4647), .ZN(U3473)
         );
  INV_X1 U5190 ( .A(n4614), .ZN(n4616) );
  AOI211_X1 U5191 ( .C1(n4618), .C2(n4617), .A(n4616), .B(n4615), .ZN(n4658)
         );
  INV_X1 U5192 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4619) );
  AOI22_X1 U5193 ( .A1(n4649), .A2(n4658), .B1(n4619), .B2(n4647), .ZN(U3475)
         );
  OAI21_X1 U5194 ( .B1(n4641), .B2(n4621), .A(n4620), .ZN(n4622) );
  AOI21_X1 U5195 ( .B1(n4623), .B2(n4646), .A(n4622), .ZN(n4659) );
  INV_X1 U5196 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4624) );
  AOI22_X1 U5197 ( .A1(n4649), .A2(n4659), .B1(n4624), .B2(n4647), .ZN(U3477)
         );
  AOI211_X1 U5198 ( .C1(n4627), .C2(n4646), .A(n4626), .B(n4625), .ZN(n4660)
         );
  INV_X1 U5199 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4628) );
  AOI22_X1 U5200 ( .A1(n4649), .A2(n4660), .B1(n4628), .B2(n4647), .ZN(U3481)
         );
  NOR2_X1 U5201 ( .A1(n4629), .A2(n4641), .ZN(n4631) );
  AOI211_X1 U5202 ( .C1(n4646), .C2(n4632), .A(n4631), .B(n4630), .ZN(n4662)
         );
  INV_X1 U5203 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4860) );
  AOI22_X1 U5204 ( .A1(n4649), .A2(n4662), .B1(n4860), .B2(n4647), .ZN(U3485)
         );
  AOI22_X1 U5205 ( .A1(n4636), .A2(n4635), .B1(n4634), .B2(n4633), .ZN(n4640)
         );
  NAND2_X1 U5206 ( .A1(n4638), .A2(n4637), .ZN(n4639) );
  OAI211_X1 U5207 ( .C1(n4642), .C2(n4641), .A(n4640), .B(n4639), .ZN(n4644)
         );
  AOI211_X1 U5208 ( .C1(n4646), .C2(n4645), .A(n4644), .B(n4643), .ZN(n4665)
         );
  INV_X1 U5209 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4648) );
  AOI22_X1 U5210 ( .A1(n4649), .A2(n4665), .B1(n4648), .B2(n4647), .ZN(U3489)
         );
  AOI22_X1 U5211 ( .A1(n4666), .A2(n4651), .B1(n4650), .B2(n4663), .ZN(U3518)
         );
  AOI22_X1 U5212 ( .A1(n4666), .A2(n4653), .B1(n4652), .B2(n4663), .ZN(U3519)
         );
  AOI22_X1 U5213 ( .A1(n4666), .A2(n4654), .B1(n4873), .B2(n4663), .ZN(U3520)
         );
  INV_X1 U5214 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4655) );
  AOI22_X1 U5215 ( .A1(n4666), .A2(n4656), .B1(n4655), .B2(n4663), .ZN(U3521)
         );
  INV_X1 U5216 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4657) );
  AOI22_X1 U5217 ( .A1(n4666), .A2(n4658), .B1(n4657), .B2(n4663), .ZN(U3522)
         );
  AOI22_X1 U5218 ( .A1(n4666), .A2(n4659), .B1(n5043), .B2(n4663), .ZN(U3523)
         );
  AOI22_X1 U5219 ( .A1(n4666), .A2(n4660), .B1(n2314), .B2(n4663), .ZN(U3525)
         );
  INV_X1 U5220 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4661) );
  AOI22_X1 U5221 ( .A1(n4666), .A2(n4662), .B1(n4661), .B2(n4663), .ZN(U3527)
         );
  AOI22_X1 U5222 ( .A1(n4666), .A2(n4665), .B1(n4664), .B2(n4663), .ZN(U3529)
         );
  INV_X1 U5223 ( .A(REG3_REG_0__SCAN_IN), .ZN(n4674) );
  NAND2_X1 U5224 ( .A1(n4668), .A2(n4667), .ZN(n4673) );
  AOI22_X1 U5225 ( .A1(n4671), .A2(n4670), .B1(n2669), .B2(n4669), .ZN(n4672)
         );
  OAI211_X1 U5226 ( .C1(n4675), .C2(n4674), .A(n4673), .B(n4672), .ZN(n5064)
         );
  OAI22_X1 U5227 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput93), .B1(keyinput73), 
        .B2(DATAO_REG_5__SCAN_IN), .ZN(n4676) );
  AOI221_X1 U5228 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput93), .C1(
        DATAO_REG_5__SCAN_IN), .C2(keyinput73), .A(n4676), .ZN(n4683) );
  OAI22_X1 U5229 ( .A1(IR_REG_21__SCAN_IN), .A2(keyinput37), .B1(keyinput25), 
        .B2(REG1_REG_30__SCAN_IN), .ZN(n4677) );
  AOI221_X1 U5230 ( .B1(IR_REG_21__SCAN_IN), .B2(keyinput37), .C1(
        REG1_REG_30__SCAN_IN), .C2(keyinput25), .A(n4677), .ZN(n4682) );
  OAI22_X1 U5231 ( .A1(D_REG_15__SCAN_IN), .A2(keyinput101), .B1(
        D_REG_11__SCAN_IN), .B2(keyinput4), .ZN(n4678) );
  AOI221_X1 U5232 ( .B1(D_REG_15__SCAN_IN), .B2(keyinput101), .C1(keyinput4), 
        .C2(D_REG_11__SCAN_IN), .A(n4678), .ZN(n4681) );
  OAI22_X1 U5233 ( .A1(IR_REG_27__SCAN_IN), .A2(keyinput81), .B1(keyinput12), 
        .B2(REG2_REG_31__SCAN_IN), .ZN(n4679) );
  AOI221_X1 U5234 ( .B1(IR_REG_27__SCAN_IN), .B2(keyinput81), .C1(
        REG2_REG_31__SCAN_IN), .C2(keyinput12), .A(n4679), .ZN(n4680) );
  NAND4_X1 U5235 ( .A1(n4683), .A2(n4682), .A3(n4681), .A4(n4680), .ZN(n4711)
         );
  OAI22_X1 U5236 ( .A1(REG2_REG_5__SCAN_IN), .A2(keyinput61), .B1(keyinput9), 
        .B2(REG1_REG_18__SCAN_IN), .ZN(n4684) );
  AOI221_X1 U5237 ( .B1(REG2_REG_5__SCAN_IN), .B2(keyinput61), .C1(
        REG1_REG_18__SCAN_IN), .C2(keyinput9), .A(n4684), .ZN(n4691) );
  OAI22_X1 U5238 ( .A1(REG0_REG_9__SCAN_IN), .A2(keyinput119), .B1(
        ADDR_REG_18__SCAN_IN), .B2(keyinput88), .ZN(n4685) );
  AOI221_X1 U5239 ( .B1(REG0_REG_9__SCAN_IN), .B2(keyinput119), .C1(keyinput88), .C2(ADDR_REG_18__SCAN_IN), .A(n4685), .ZN(n4690) );
  OAI22_X1 U5240 ( .A1(REG0_REG_14__SCAN_IN), .A2(keyinput33), .B1(
        DATAO_REG_20__SCAN_IN), .B2(keyinput1), .ZN(n4686) );
  AOI221_X1 U5241 ( .B1(REG0_REG_14__SCAN_IN), .B2(keyinput33), .C1(keyinput1), 
        .C2(DATAO_REG_20__SCAN_IN), .A(n4686), .ZN(n4689) );
  OAI22_X1 U5242 ( .A1(IR_REG_15__SCAN_IN), .A2(keyinput17), .B1(keyinput57), 
        .B2(REG1_REG_2__SCAN_IN), .ZN(n4687) );
  AOI221_X1 U5243 ( .B1(IR_REG_15__SCAN_IN), .B2(keyinput17), .C1(
        REG1_REG_2__SCAN_IN), .C2(keyinput57), .A(n4687), .ZN(n4688) );
  NAND4_X1 U5244 ( .A1(n4691), .A2(n4690), .A3(n4689), .A4(n4688), .ZN(n4710)
         );
  OAI22_X1 U5245 ( .A1(IR_REG_11__SCAN_IN), .A2(keyinput122), .B1(keyinput102), 
        .B2(REG2_REG_4__SCAN_IN), .ZN(n4692) );
  AOI221_X1 U5246 ( .B1(IR_REG_11__SCAN_IN), .B2(keyinput122), .C1(
        REG2_REG_4__SCAN_IN), .C2(keyinput102), .A(n4692), .ZN(n4699) );
  OAI22_X1 U5247 ( .A1(IR_REG_4__SCAN_IN), .A2(keyinput98), .B1(keyinput106), 
        .B2(DATAI_7_), .ZN(n4693) );
  AOI221_X1 U5248 ( .B1(IR_REG_4__SCAN_IN), .B2(keyinput98), .C1(DATAI_7_), 
        .C2(keyinput106), .A(n4693), .ZN(n4698) );
  OAI22_X1 U5249 ( .A1(D_REG_26__SCAN_IN), .A2(keyinput22), .B1(keyinput6), 
        .B2(REG3_REG_18__SCAN_IN), .ZN(n4694) );
  AOI221_X1 U5250 ( .B1(D_REG_26__SCAN_IN), .B2(keyinput22), .C1(
        REG3_REG_18__SCAN_IN), .C2(keyinput6), .A(n4694), .ZN(n4697) );
  OAI22_X1 U5251 ( .A1(IR_REG_25__SCAN_IN), .A2(keyinput2), .B1(keyinput18), 
        .B2(REG1_REG_13__SCAN_IN), .ZN(n4695) );
  AOI221_X1 U5252 ( .B1(IR_REG_25__SCAN_IN), .B2(keyinput2), .C1(
        REG1_REG_13__SCAN_IN), .C2(keyinput18), .A(n4695), .ZN(n4696) );
  NAND4_X1 U5253 ( .A1(n4699), .A2(n4698), .A3(n4697), .A4(n4696), .ZN(n4709)
         );
  OAI22_X1 U5254 ( .A1(IR_REG_9__SCAN_IN), .A2(keyinput58), .B1(
        REG3_REG_8__SCAN_IN), .B2(keyinput50), .ZN(n4700) );
  AOI221_X1 U5255 ( .B1(IR_REG_9__SCAN_IN), .B2(keyinput58), .C1(keyinput50), 
        .C2(REG3_REG_8__SCAN_IN), .A(n4700), .ZN(n4707) );
  OAI22_X1 U5256 ( .A1(D_REG_5__SCAN_IN), .A2(keyinput77), .B1(
        REG0_REG_26__SCAN_IN), .B2(keyinput69), .ZN(n4701) );
  AOI221_X1 U5257 ( .B1(D_REG_5__SCAN_IN), .B2(keyinput77), .C1(keyinput69), 
        .C2(REG0_REG_26__SCAN_IN), .A(n4701), .ZN(n4706) );
  OAI22_X1 U5258 ( .A1(D_REG_18__SCAN_IN), .A2(keyinput78), .B1(keyinput82), 
        .B2(DATAI_8_), .ZN(n4702) );
  AOI221_X1 U5259 ( .B1(D_REG_18__SCAN_IN), .B2(keyinput78), .C1(DATAI_8_), 
        .C2(keyinput82), .A(n4702), .ZN(n4705) );
  OAI22_X1 U5260 ( .A1(DATAI_3_), .A2(keyinput86), .B1(keyinput66), .B2(
        REG2_REG_30__SCAN_IN), .ZN(n4703) );
  AOI221_X1 U5261 ( .B1(DATAI_3_), .B2(keyinput86), .C1(REG2_REG_30__SCAN_IN), 
        .C2(keyinput66), .A(n4703), .ZN(n4704) );
  NAND4_X1 U5262 ( .A1(n4707), .A2(n4706), .A3(n4705), .A4(n4704), .ZN(n4708)
         );
  NOR4_X1 U5263 ( .A1(n4711), .A2(n4710), .A3(n4709), .A4(n4708), .ZN(n5062)
         );
  OAI22_X1 U5264 ( .A1(B_REG_SCAN_IN), .A2(keyinput43), .B1(keyinput63), .B2(
        REG3_REG_13__SCAN_IN), .ZN(n4712) );
  AOI221_X1 U5265 ( .B1(B_REG_SCAN_IN), .B2(keyinput43), .C1(
        REG3_REG_13__SCAN_IN), .C2(keyinput63), .A(n4712), .ZN(n4719) );
  OAI22_X1 U5266 ( .A1(REG1_REG_6__SCAN_IN), .A2(keyinput67), .B1(DATAI_13_), 
        .B2(keyinput71), .ZN(n4713) );
  AOI221_X1 U5267 ( .B1(REG1_REG_6__SCAN_IN), .B2(keyinput67), .C1(keyinput71), 
        .C2(DATAI_13_), .A(n4713), .ZN(n4718) );
  OAI22_X1 U5268 ( .A1(D_REG_14__SCAN_IN), .A2(keyinput27), .B1(keyinput23), 
        .B2(REG2_REG_15__SCAN_IN), .ZN(n4714) );
  AOI221_X1 U5269 ( .B1(D_REG_14__SCAN_IN), .B2(keyinput27), .C1(
        REG2_REG_15__SCAN_IN), .C2(keyinput23), .A(n4714), .ZN(n4717) );
  OAI22_X1 U5270 ( .A1(REG3_REG_6__SCAN_IN), .A2(keyinput31), .B1(keyinput39), 
        .B2(REG0_REG_16__SCAN_IN), .ZN(n4715) );
  AOI221_X1 U5271 ( .B1(REG3_REG_6__SCAN_IN), .B2(keyinput31), .C1(
        REG0_REG_16__SCAN_IN), .C2(keyinput39), .A(n4715), .ZN(n4716) );
  NAND4_X1 U5272 ( .A1(n4719), .A2(n4718), .A3(n4717), .A4(n4716), .ZN(n4747)
         );
  OAI22_X1 U5273 ( .A1(D_REG_17__SCAN_IN), .A2(keyinput115), .B1(keyinput111), 
        .B2(REG2_REG_27__SCAN_IN), .ZN(n4720) );
  AOI221_X1 U5274 ( .B1(D_REG_17__SCAN_IN), .B2(keyinput115), .C1(
        REG2_REG_27__SCAN_IN), .C2(keyinput111), .A(n4720), .ZN(n4727) );
  OAI22_X1 U5275 ( .A1(REG2_REG_23__SCAN_IN), .A2(keyinput95), .B1(
        DATAO_REG_30__SCAN_IN), .B2(keyinput91), .ZN(n4721) );
  AOI221_X1 U5276 ( .B1(REG2_REG_23__SCAN_IN), .B2(keyinput95), .C1(keyinput91), .C2(DATAO_REG_30__SCAN_IN), .A(n4721), .ZN(n4726) );
  OAI22_X1 U5277 ( .A1(REG1_REG_7__SCAN_IN), .A2(keyinput79), .B1(keyinput75), 
        .B2(ADDR_REG_8__SCAN_IN), .ZN(n4722) );
  AOI221_X1 U5278 ( .B1(REG1_REG_7__SCAN_IN), .B2(keyinput79), .C1(
        ADDR_REG_8__SCAN_IN), .C2(keyinput75), .A(n4722), .ZN(n4725) );
  OAI22_X1 U5279 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput83), .B1(keyinput87), 
        .B2(DATAI_23_), .ZN(n4723) );
  AOI221_X1 U5280 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput83), .C1(DATAI_23_), 
        .C2(keyinput87), .A(n4723), .ZN(n4724) );
  NAND4_X1 U5281 ( .A1(n4727), .A2(n4726), .A3(n4725), .A4(n4724), .ZN(n4746)
         );
  OAI22_X1 U5282 ( .A1(DATAO_REG_2__SCAN_IN), .A2(keyinput96), .B1(keyinput123), .B2(DATAO_REG_6__SCAN_IN), .ZN(n4728) );
  AOI221_X1 U5283 ( .B1(DATAO_REG_2__SCAN_IN), .B2(keyinput96), .C1(
        DATAO_REG_6__SCAN_IN), .C2(keyinput123), .A(n4728), .ZN(n4735) );
  OAI22_X1 U5284 ( .A1(D_REG_19__SCAN_IN), .A2(keyinput56), .B1(
        DATAO_REG_8__SCAN_IN), .B2(keyinput28), .ZN(n4729) );
  AOI221_X1 U5285 ( .B1(D_REG_19__SCAN_IN), .B2(keyinput56), .C1(keyinput28), 
        .C2(DATAO_REG_8__SCAN_IN), .A(n4729), .ZN(n4734) );
  OAI22_X1 U5286 ( .A1(D_REG_0__SCAN_IN), .A2(keyinput100), .B1(keyinput112), 
        .B2(ADDR_REG_16__SCAN_IN), .ZN(n4730) );
  AOI221_X1 U5287 ( .B1(D_REG_0__SCAN_IN), .B2(keyinput100), .C1(
        ADDR_REG_16__SCAN_IN), .C2(keyinput112), .A(n4730), .ZN(n4733) );
  OAI22_X1 U5288 ( .A1(DATAI_28_), .A2(keyinput116), .B1(keyinput108), .B2(
        REG2_REG_26__SCAN_IN), .ZN(n4731) );
  AOI221_X1 U5289 ( .B1(DATAI_28_), .B2(keyinput116), .C1(REG2_REG_26__SCAN_IN), .C2(keyinput108), .A(n4731), .ZN(n4732) );
  NAND4_X1 U5290 ( .A1(n4735), .A2(n4734), .A3(n4733), .A4(n4732), .ZN(n4745)
         );
  OAI22_X1 U5291 ( .A1(STATE_REG_SCAN_IN), .A2(keyinput20), .B1(DATAI_31_), 
        .B2(keyinput76), .ZN(n4736) );
  AOI221_X1 U5292 ( .B1(STATE_REG_SCAN_IN), .B2(keyinput20), .C1(keyinput76), 
        .C2(DATAI_31_), .A(n4736), .ZN(n4743) );
  OAI22_X1 U5293 ( .A1(IR_REG_26__SCAN_IN), .A2(keyinput3), .B1(keyinput19), 
        .B2(REG2_REG_6__SCAN_IN), .ZN(n4737) );
  AOI221_X1 U5294 ( .B1(IR_REG_26__SCAN_IN), .B2(keyinput3), .C1(
        REG2_REG_6__SCAN_IN), .C2(keyinput19), .A(n4737), .ZN(n4742) );
  OAI22_X1 U5295 ( .A1(IR_REG_7__SCAN_IN), .A2(keyinput92), .B1(
        DATAO_REG_24__SCAN_IN), .B2(keyinput48), .ZN(n4738) );
  AOI221_X1 U5296 ( .B1(IR_REG_7__SCAN_IN), .B2(keyinput92), .C1(keyinput48), 
        .C2(DATAO_REG_24__SCAN_IN), .A(n4738), .ZN(n4741) );
  OAI22_X1 U5297 ( .A1(REG3_REG_15__SCAN_IN), .A2(keyinput84), .B1(
        REG2_REG_1__SCAN_IN), .B2(keyinput8), .ZN(n4739) );
  AOI221_X1 U5298 ( .B1(REG3_REG_15__SCAN_IN), .B2(keyinput84), .C1(keyinput8), 
        .C2(REG2_REG_1__SCAN_IN), .A(n4739), .ZN(n4740) );
  NAND4_X1 U5299 ( .A1(n4743), .A2(n4742), .A3(n4741), .A4(n4740), .ZN(n4744)
         );
  NOR4_X1 U5300 ( .A1(n4747), .A2(n4746), .A3(n4745), .A4(n4744), .ZN(n5061)
         );
  AOI22_X1 U5301 ( .A1(DATAI_30_), .A2(keyinput222), .B1(DATAI_23_), .B2(
        keyinput215), .ZN(n4748) );
  OAI221_X1 U5302 ( .B1(DATAI_30_), .B2(keyinput222), .C1(DATAI_23_), .C2(
        keyinput215), .A(n4748), .ZN(n4755) );
  AOI22_X1 U5303 ( .A1(DATAI_19_), .A2(keyinput182), .B1(DATAI_22_), .B2(
        keyinput181), .ZN(n4749) );
  OAI221_X1 U5304 ( .B1(DATAI_19_), .B2(keyinput182), .C1(DATAI_22_), .C2(
        keyinput181), .A(n4749), .ZN(n4754) );
  AOI22_X1 U5305 ( .A1(DATAI_15_), .A2(keyinput180), .B1(DATAI_7_), .B2(
        keyinput234), .ZN(n4750) );
  OAI221_X1 U5306 ( .B1(DATAI_15_), .B2(keyinput180), .C1(DATAI_7_), .C2(
        keyinput234), .A(n4750), .ZN(n4753) );
  AOI22_X1 U5307 ( .A1(REG3_REG_21__SCAN_IN), .A2(keyinput237), .B1(
        REG3_REG_28__SCAN_IN), .B2(keyinput245), .ZN(n4751) );
  OAI221_X1 U5308 ( .B1(REG3_REG_21__SCAN_IN), .B2(keyinput237), .C1(
        REG3_REG_28__SCAN_IN), .C2(keyinput245), .A(n4751), .ZN(n4752) );
  NOR4_X1 U5309 ( .A1(n4755), .A2(n4754), .A3(n4753), .A4(n4752), .ZN(n4783)
         );
  AOI22_X1 U5310 ( .A1(IR_REG_0__SCAN_IN), .A2(keyinput225), .B1(
        IR_REG_4__SCAN_IN), .B2(keyinput226), .ZN(n4756) );
  OAI221_X1 U5311 ( .B1(IR_REG_0__SCAN_IN), .B2(keyinput225), .C1(
        IR_REG_4__SCAN_IN), .C2(keyinput226), .A(n4756), .ZN(n4763) );
  AOI22_X1 U5312 ( .A1(IR_REG_6__SCAN_IN), .A2(keyinput162), .B1(
        IR_REG_11__SCAN_IN), .B2(keyinput250), .ZN(n4757) );
  OAI221_X1 U5313 ( .B1(IR_REG_6__SCAN_IN), .B2(keyinput162), .C1(
        IR_REG_11__SCAN_IN), .C2(keyinput250), .A(n4757), .ZN(n4762) );
  AOI22_X1 U5314 ( .A1(IR_REG_19__SCAN_IN), .A2(keyinput170), .B1(
        IR_REG_16__SCAN_IN), .B2(keyinput169), .ZN(n4758) );
  OAI221_X1 U5315 ( .B1(IR_REG_19__SCAN_IN), .B2(keyinput170), .C1(
        IR_REG_16__SCAN_IN), .C2(keyinput169), .A(n4758), .ZN(n4761) );
  AOI22_X1 U5316 ( .A1(IR_REG_21__SCAN_IN), .A2(keyinput165), .B1(
        IR_REG_22__SCAN_IN), .B2(keyinput139), .ZN(n4759) );
  OAI221_X1 U5317 ( .B1(IR_REG_21__SCAN_IN), .B2(keyinput165), .C1(
        IR_REG_22__SCAN_IN), .C2(keyinput139), .A(n4759), .ZN(n4760) );
  NOR4_X1 U5318 ( .A1(n4763), .A2(n4762), .A3(n4761), .A4(n4760), .ZN(n4782)
         );
  AOI22_X1 U5319 ( .A1(IR_REG_27__SCAN_IN), .A2(keyinput209), .B1(
        IR_REG_25__SCAN_IN), .B2(keyinput130), .ZN(n4764) );
  OAI221_X1 U5320 ( .B1(IR_REG_27__SCAN_IN), .B2(keyinput209), .C1(
        IR_REG_25__SCAN_IN), .C2(keyinput130), .A(n4764), .ZN(n4771) );
  AOI22_X1 U5321 ( .A1(D_REG_5__SCAN_IN), .A2(keyinput205), .B1(
        D_REG_0__SCAN_IN), .B2(keyinput228), .ZN(n4765) );
  OAI221_X1 U5322 ( .B1(D_REG_5__SCAN_IN), .B2(keyinput205), .C1(
        D_REG_0__SCAN_IN), .C2(keyinput228), .A(n4765), .ZN(n4770) );
  AOI22_X1 U5323 ( .A1(D_REG_11__SCAN_IN), .A2(keyinput132), .B1(
        D_REG_14__SCAN_IN), .B2(keyinput155), .ZN(n4766) );
  OAI221_X1 U5324 ( .B1(D_REG_11__SCAN_IN), .B2(keyinput132), .C1(
        D_REG_14__SCAN_IN), .C2(keyinput155), .A(n4766), .ZN(n4769) );
  AOI22_X1 U5325 ( .A1(D_REG_15__SCAN_IN), .A2(keyinput229), .B1(
        D_REG_17__SCAN_IN), .B2(keyinput243), .ZN(n4767) );
  OAI221_X1 U5326 ( .B1(D_REG_15__SCAN_IN), .B2(keyinput229), .C1(
        D_REG_17__SCAN_IN), .C2(keyinput243), .A(n4767), .ZN(n4768) );
  NOR4_X1 U5327 ( .A1(n4771), .A2(n4770), .A3(n4769), .A4(n4768), .ZN(n4781)
         );
  AOI22_X1 U5328 ( .A1(D_REG_31__SCAN_IN), .A2(keyinput253), .B1(
        D_REG_26__SCAN_IN), .B2(keyinput150), .ZN(n4772) );
  OAI221_X1 U5329 ( .B1(D_REG_31__SCAN_IN), .B2(keyinput253), .C1(
        D_REG_26__SCAN_IN), .C2(keyinput150), .A(n4772), .ZN(n4779) );
  AOI22_X1 U5330 ( .A1(REG0_REG_16__SCAN_IN), .A2(keyinput167), .B1(
        REG0_REG_25__SCAN_IN), .B2(keyinput246), .ZN(n4773) );
  OAI221_X1 U5331 ( .B1(REG0_REG_16__SCAN_IN), .B2(keyinput167), .C1(
        REG0_REG_25__SCAN_IN), .C2(keyinput246), .A(n4773), .ZN(n4778) );
  AOI22_X1 U5332 ( .A1(REG0_REG_31__SCAN_IN), .A2(keyinput183), .B1(
        REG0_REG_30__SCAN_IN), .B2(keyinput227), .ZN(n4774) );
  OAI221_X1 U5333 ( .B1(REG0_REG_31__SCAN_IN), .B2(keyinput183), .C1(
        REG0_REG_30__SCAN_IN), .C2(keyinput227), .A(n4774), .ZN(n4777) );
  AOI22_X1 U5334 ( .A1(REG1_REG_13__SCAN_IN), .A2(keyinput146), .B1(
        REG1_REG_5__SCAN_IN), .B2(keyinput163), .ZN(n4775) );
  OAI221_X1 U5335 ( .B1(REG1_REG_13__SCAN_IN), .B2(keyinput146), .C1(
        REG1_REG_5__SCAN_IN), .C2(keyinput163), .A(n4775), .ZN(n4776) );
  NOR4_X1 U5336 ( .A1(n4779), .A2(n4778), .A3(n4777), .A4(n4776), .ZN(n4780)
         );
  NAND4_X1 U5337 ( .A1(n4783), .A2(n4782), .A3(n4781), .A4(n4780), .ZN(n4927)
         );
  AOI22_X1 U5338 ( .A1(REG1_REG_24__SCAN_IN), .A2(keyinput187), .B1(
        REG1_REG_21__SCAN_IN), .B2(keyinput158), .ZN(n4784) );
  OAI221_X1 U5339 ( .B1(REG1_REG_24__SCAN_IN), .B2(keyinput187), .C1(
        REG1_REG_21__SCAN_IN), .C2(keyinput158), .A(n4784), .ZN(n4791) );
  AOI22_X1 U5340 ( .A1(REG2_REG_1__SCAN_IN), .A2(keyinput136), .B1(
        REG1_REG_25__SCAN_IN), .B2(keyinput142), .ZN(n4785) );
  OAI221_X1 U5341 ( .B1(REG2_REG_1__SCAN_IN), .B2(keyinput136), .C1(
        REG1_REG_25__SCAN_IN), .C2(keyinput142), .A(n4785), .ZN(n4790) );
  AOI22_X1 U5342 ( .A1(REG1_REG_31__SCAN_IN), .A2(keyinput160), .B1(
        REG2_REG_5__SCAN_IN), .B2(keyinput189), .ZN(n4786) );
  OAI221_X1 U5343 ( .B1(REG1_REG_31__SCAN_IN), .B2(keyinput160), .C1(
        REG2_REG_5__SCAN_IN), .C2(keyinput189), .A(n4786), .ZN(n4789) );
  AOI22_X1 U5344 ( .A1(REG2_REG_6__SCAN_IN), .A2(keyinput147), .B1(
        REG2_REG_8__SCAN_IN), .B2(keyinput232), .ZN(n4787) );
  OAI221_X1 U5345 ( .B1(REG2_REG_6__SCAN_IN), .B2(keyinput147), .C1(
        REG2_REG_8__SCAN_IN), .C2(keyinput232), .A(n4787), .ZN(n4788) );
  NOR4_X1 U5346 ( .A1(n4791), .A2(n4790), .A3(n4789), .A4(n4788), .ZN(n4819)
         );
  AOI22_X1 U5347 ( .A1(REG2_REG_15__SCAN_IN), .A2(keyinput151), .B1(
        REG2_REG_13__SCAN_IN), .B2(keyinput152), .ZN(n4792) );
  OAI221_X1 U5348 ( .B1(REG2_REG_15__SCAN_IN), .B2(keyinput151), .C1(
        REG2_REG_13__SCAN_IN), .C2(keyinput152), .A(n4792), .ZN(n4799) );
  AOI22_X1 U5349 ( .A1(REG2_REG_21__SCAN_IN), .A2(keyinput196), .B1(
        REG2_REG_22__SCAN_IN), .B2(keyinput233), .ZN(n4793) );
  OAI221_X1 U5350 ( .B1(REG2_REG_21__SCAN_IN), .B2(keyinput196), .C1(
        REG2_REG_22__SCAN_IN), .C2(keyinput233), .A(n4793), .ZN(n4798) );
  AOI22_X1 U5351 ( .A1(REG2_REG_24__SCAN_IN), .A2(keyinput168), .B1(
        REG2_REG_23__SCAN_IN), .B2(keyinput223), .ZN(n4794) );
  OAI221_X1 U5352 ( .B1(REG2_REG_24__SCAN_IN), .B2(keyinput168), .C1(
        REG2_REG_23__SCAN_IN), .C2(keyinput223), .A(n4794), .ZN(n4797) );
  AOI22_X1 U5353 ( .A1(ADDR_REG_9__SCAN_IN), .A2(keyinput249), .B1(
        ADDR_REG_16__SCAN_IN), .B2(keyinput240), .ZN(n4795) );
  OAI221_X1 U5354 ( .B1(ADDR_REG_9__SCAN_IN), .B2(keyinput249), .C1(
        ADDR_REG_16__SCAN_IN), .C2(keyinput240), .A(n4795), .ZN(n4796) );
  NOR4_X1 U5355 ( .A1(n4799), .A2(n4798), .A3(n4797), .A4(n4796), .ZN(n4818)
         );
  AOI22_X1 U5356 ( .A1(ADDR_REG_1__SCAN_IN), .A2(keyinput213), .B1(
        ADDR_REG_4__SCAN_IN), .B2(keyinput248), .ZN(n4800) );
  OAI221_X1 U5357 ( .B1(ADDR_REG_1__SCAN_IN), .B2(keyinput213), .C1(
        ADDR_REG_4__SCAN_IN), .C2(keyinput248), .A(n4800), .ZN(n4807) );
  AOI22_X1 U5358 ( .A1(DATAO_REG_5__SCAN_IN), .A2(keyinput201), .B1(
        DATAO_REG_0__SCAN_IN), .B2(keyinput135), .ZN(n4801) );
  OAI221_X1 U5359 ( .B1(DATAO_REG_5__SCAN_IN), .B2(keyinput201), .C1(
        DATAO_REG_0__SCAN_IN), .C2(keyinput135), .A(n4801), .ZN(n4806) );
  AOI22_X1 U5360 ( .A1(DATAO_REG_6__SCAN_IN), .A2(keyinput251), .B1(
        DATAO_REG_2__SCAN_IN), .B2(keyinput224), .ZN(n4802) );
  OAI221_X1 U5361 ( .B1(DATAO_REG_6__SCAN_IN), .B2(keyinput251), .C1(
        DATAO_REG_2__SCAN_IN), .C2(keyinput224), .A(n4802), .ZN(n4805) );
  AOI22_X1 U5362 ( .A1(DATAO_REG_20__SCAN_IN), .A2(keyinput129), .B1(
        DATAO_REG_13__SCAN_IN), .B2(keyinput242), .ZN(n4803) );
  OAI221_X1 U5363 ( .B1(DATAO_REG_20__SCAN_IN), .B2(keyinput129), .C1(
        DATAO_REG_13__SCAN_IN), .C2(keyinput242), .A(n4803), .ZN(n4804) );
  NOR4_X1 U5364 ( .A1(n4807), .A2(n4806), .A3(n4805), .A4(n4804), .ZN(n4817)
         );
  AOI22_X1 U5365 ( .A1(DATAO_REG_31__SCAN_IN), .A2(keyinput133), .B1(
        DATAO_REG_23__SCAN_IN), .B2(keyinput175), .ZN(n4808) );
  OAI221_X1 U5366 ( .B1(DATAO_REG_31__SCAN_IN), .B2(keyinput133), .C1(
        DATAO_REG_23__SCAN_IN), .C2(keyinput175), .A(n4808), .ZN(n4815) );
  AOI22_X1 U5367 ( .A1(REG3_REG_6__SCAN_IN), .A2(keyinput159), .B1(
        REG3_REG_15__SCAN_IN), .B2(keyinput212), .ZN(n4809) );
  OAI221_X1 U5368 ( .B1(REG3_REG_6__SCAN_IN), .B2(keyinput159), .C1(
        REG3_REG_15__SCAN_IN), .C2(keyinput212), .A(n4809), .ZN(n4814) );
  AOI22_X1 U5369 ( .A1(REG2_REG_26__SCAN_IN), .A2(keyinput236), .B1(
        REG3_REG_22__SCAN_IN), .B2(keyinput164), .ZN(n4810) );
  OAI221_X1 U5370 ( .B1(REG2_REG_26__SCAN_IN), .B2(keyinput236), .C1(
        REG3_REG_22__SCAN_IN), .C2(keyinput164), .A(n4810), .ZN(n4813) );
  AOI22_X1 U5371 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput221), .B1(
        D_REG_8__SCAN_IN), .B2(keyinput143), .ZN(n4811) );
  OAI221_X1 U5372 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput221), .C1(
        D_REG_8__SCAN_IN), .C2(keyinput143), .A(n4811), .ZN(n4812) );
  NOR4_X1 U5373 ( .A1(n4815), .A2(n4814), .A3(n4813), .A4(n4812), .ZN(n4816)
         );
  NAND4_X1 U5374 ( .A1(n4819), .A2(n4818), .A3(n4817), .A4(n4816), .ZN(n4926)
         );
  AOI22_X1 U5375 ( .A1(n4822), .A2(keyinput204), .B1(n4821), .B2(keyinput244), 
        .ZN(n4820) );
  OAI221_X1 U5376 ( .B1(n4822), .B2(keyinput204), .C1(n4821), .C2(keyinput244), 
        .A(n4820), .ZN(n4830) );
  INV_X1 U5377 ( .A(DATAI_24_), .ZN(n4979) );
  AOI22_X1 U5378 ( .A1(n4982), .A2(keyinput190), .B1(keyinput144), .B2(n4979), 
        .ZN(n4823) );
  OAI221_X1 U5379 ( .B1(n4982), .B2(keyinput190), .C1(n4979), .C2(keyinput144), 
        .A(n4823), .ZN(n4829) );
  INV_X1 U5380 ( .A(DATAI_16_), .ZN(n5002) );
  AOI22_X1 U5381 ( .A1(n4999), .A2(keyinput218), .B1(keyinput198), .B2(n5002), 
        .ZN(n4824) );
  OAI221_X1 U5382 ( .B1(n4999), .B2(keyinput218), .C1(n5002), .C2(keyinput198), 
        .A(n4824), .ZN(n4828) );
  AOI22_X1 U5383 ( .A1(n2763), .A2(keyinput199), .B1(n4826), .B2(keyinput210), 
        .ZN(n4825) );
  OAI221_X1 U5384 ( .B1(n2763), .B2(keyinput199), .C1(n4826), .C2(keyinput210), 
        .A(n4825), .ZN(n4827) );
  NOR4_X1 U5385 ( .A1(n4830), .A2(n4829), .A3(n4828), .A4(n4827), .ZN(n4871)
         );
  AOI22_X1 U5386 ( .A1(n4946), .A2(keyinput217), .B1(keyinput128), .B2(n5014), 
        .ZN(n4831) );
  OAI221_X1 U5387 ( .B1(n4946), .B2(keyinput217), .C1(n5014), .C2(keyinput128), 
        .A(n4831), .ZN(n4841) );
  AOI22_X1 U5388 ( .A1(n4833), .A2(keyinput214), .B1(keyinput141), .B2(n2334), 
        .ZN(n4832) );
  OAI221_X1 U5389 ( .B1(n4833), .B2(keyinput214), .C1(n2334), .C2(keyinput141), 
        .A(n4832), .ZN(n4840) );
  AOI22_X1 U5390 ( .A1(U3149), .A2(keyinput148), .B1(keyinput138), .B2(n5031), 
        .ZN(n4834) );
  OAI221_X1 U5391 ( .B1(U3149), .B2(keyinput148), .C1(n5031), .C2(keyinput138), 
        .A(n4834), .ZN(n4839) );
  AOI22_X1 U5392 ( .A1(n4837), .A2(keyinput178), .B1(n4836), .B2(keyinput191), 
        .ZN(n4835) );
  OAI221_X1 U5393 ( .B1(n4837), .B2(keyinput178), .C1(n4836), .C2(keyinput191), 
        .A(n4835), .ZN(n4838) );
  NOR4_X1 U5394 ( .A1(n4841), .A2(n4840), .A3(n4839), .A4(n4838), .ZN(n4870)
         );
  XNOR2_X1 U5395 ( .A(n4842), .B(keyinput131), .ZN(n4847) );
  XNOR2_X1 U5396 ( .A(n4843), .B(keyinput186), .ZN(n4846) );
  XNOR2_X1 U5397 ( .A(n4844), .B(keyinput220), .ZN(n4845) );
  NOR3_X1 U5398 ( .A1(n4847), .A2(n4846), .A3(n4845), .ZN(n4850) );
  XNOR2_X1 U5399 ( .A(IR_REG_15__SCAN_IN), .B(keyinput145), .ZN(n4849) );
  XNOR2_X1 U5400 ( .A(IR_REG_14__SCAN_IN), .B(keyinput252), .ZN(n4848) );
  NAND3_X1 U5401 ( .A1(n4850), .A2(n4849), .A3(n4848), .ZN(n4854) );
  AOI22_X1 U5402 ( .A1(n5027), .A2(keyinput255), .B1(n5018), .B2(keyinput192), 
        .ZN(n4851) );
  OAI221_X1 U5403 ( .B1(n5027), .B2(keyinput255), .C1(n5018), .C2(keyinput192), 
        .A(n4851), .ZN(n4853) );
  XNOR2_X1 U5404 ( .A(n5015), .B(keyinput231), .ZN(n4852) );
  NOR3_X1 U5405 ( .A1(n4854), .A2(n4853), .A3(n4852), .ZN(n4869) );
  AOI22_X1 U5406 ( .A1(n4857), .A2(keyinput206), .B1(n4856), .B2(keyinput184), 
        .ZN(n4855) );
  OAI221_X1 U5407 ( .B1(n4857), .B2(keyinput206), .C1(n4856), .C2(keyinput184), 
        .A(n4855), .ZN(n4867) );
  AOI22_X1 U5408 ( .A1(n5028), .A2(keyinput254), .B1(keyinput235), .B2(n5009), 
        .ZN(n4858) );
  OAI221_X1 U5409 ( .B1(n5028), .B2(keyinput254), .C1(n5009), .C2(keyinput235), 
        .A(n4858), .ZN(n4866) );
  INV_X1 U5410 ( .A(REG0_REG_10__SCAN_IN), .ZN(n5039) );
  AOI22_X1 U5411 ( .A1(n5039), .A2(keyinput154), .B1(keyinput247), .B2(n4860), 
        .ZN(n4859) );
  OAI221_X1 U5412 ( .B1(n5039), .B2(keyinput154), .C1(n4860), .C2(keyinput247), 
        .A(n4859), .ZN(n4865) );
  AOI22_X1 U5413 ( .A1(n4863), .A2(keyinput161), .B1(n4862), .B2(keyinput197), 
        .ZN(n4861) );
  OAI221_X1 U5414 ( .B1(n4863), .B2(keyinput161), .C1(n4862), .C2(keyinput197), 
        .A(n4861), .ZN(n4864) );
  NOR4_X1 U5415 ( .A1(n4867), .A2(n4866), .A3(n4865), .A4(n4864), .ZN(n4868)
         );
  NAND4_X1 U5416 ( .A1(n4871), .A2(n4870), .A3(n4869), .A4(n4868), .ZN(n4925)
         );
  INV_X1 U5417 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4960) );
  AOI22_X1 U5418 ( .A1(n4960), .A2(keyinput208), .B1(keyinput185), .B2(n4873), 
        .ZN(n4872) );
  OAI221_X1 U5419 ( .B1(n4960), .B2(keyinput208), .C1(n4873), .C2(keyinput185), 
        .A(n4872), .ZN(n4883) );
  INV_X1 U5420 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4875) );
  AOI22_X1 U5421 ( .A1(n4875), .A2(keyinput195), .B1(n2314), .B2(keyinput207), 
        .ZN(n4874) );
  OAI221_X1 U5422 ( .B1(n4875), .B2(keyinput195), .C1(n2314), .C2(keyinput207), 
        .A(n4874), .ZN(n4882) );
  INV_X1 U5423 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4877) );
  AOI22_X1 U5424 ( .A1(n4877), .A2(keyinput137), .B1(n4951), .B2(keyinput188), 
        .ZN(n4876) );
  OAI221_X1 U5425 ( .B1(n4877), .B2(keyinput137), .C1(n4951), .C2(keyinput188), 
        .A(n4876), .ZN(n4881) );
  INV_X1 U5426 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4943) );
  INV_X1 U5427 ( .A(REG1_REG_29__SCAN_IN), .ZN(n4879) );
  AOI22_X1 U5428 ( .A1(n4943), .A2(keyinput193), .B1(n4879), .B2(keyinput173), 
        .ZN(n4878) );
  OAI221_X1 U5429 ( .B1(n4943), .B2(keyinput193), .C1(n4879), .C2(keyinput173), 
        .A(n4878), .ZN(n4880) );
  NOR4_X1 U5430 ( .A1(n4883), .A2(n4882), .A3(n4881), .A4(n4880), .ZN(n4923)
         );
  INV_X1 U5431 ( .A(REG2_REG_4__SCAN_IN), .ZN(n4885) );
  AOI22_X1 U5432 ( .A1(n4886), .A2(keyinput153), .B1(n4885), .B2(keyinput230), 
        .ZN(n4884) );
  OAI221_X1 U5433 ( .B1(n4886), .B2(keyinput153), .C1(n4885), .C2(keyinput230), 
        .A(n4884), .ZN(n4896) );
  INV_X1 U5434 ( .A(REG2_REG_20__SCAN_IN), .ZN(n5044) );
  AOI22_X1 U5435 ( .A1(n4976), .A2(keyinput172), .B1(n5044), .B2(keyinput166), 
        .ZN(n4887) );
  OAI221_X1 U5436 ( .B1(n4976), .B2(keyinput172), .C1(n5044), .C2(keyinput166), 
        .A(n4887), .ZN(n4895) );
  INV_X1 U5437 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4963) );
  INV_X1 U5438 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4889) );
  AOI22_X1 U5439 ( .A1(n4963), .A2(keyinput200), .B1(n4889), .B2(keyinput239), 
        .ZN(n4888) );
  OAI221_X1 U5440 ( .B1(n4963), .B2(keyinput200), .C1(n4889), .C2(keyinput239), 
        .A(n4888), .ZN(n4894) );
  AOI22_X1 U5441 ( .A1(n4892), .A2(keyinput140), .B1(n4891), .B2(keyinput194), 
        .ZN(n4890) );
  OAI221_X1 U5442 ( .B1(n4892), .B2(keyinput140), .C1(n4891), .C2(keyinput194), 
        .A(n4890), .ZN(n4893) );
  NOR4_X1 U5443 ( .A1(n4896), .A2(n4895), .A3(n4894), .A4(n4893), .ZN(n4922)
         );
  AOI22_X1 U5444 ( .A1(n4898), .A2(keyinput216), .B1(keyinput238), .B2(n5008), 
        .ZN(n4897) );
  OAI221_X1 U5445 ( .B1(n4898), .B2(keyinput216), .C1(n5008), .C2(keyinput238), 
        .A(n4897), .ZN(n4908) );
  INV_X1 U5446 ( .A(ADDR_REG_8__SCAN_IN), .ZN(n4900) );
  AOI22_X1 U5447 ( .A1(n4900), .A2(keyinput203), .B1(keyinput202), .B2(n4998), 
        .ZN(n4899) );
  OAI221_X1 U5448 ( .B1(n4900), .B2(keyinput203), .C1(n4998), .C2(keyinput202), 
        .A(n4899), .ZN(n4907) );
  AOI22_X1 U5449 ( .A1(n4902), .A2(keyinput156), .B1(keyinput174), .B2(n4995), 
        .ZN(n4901) );
  OAI221_X1 U5450 ( .B1(n4902), .B2(keyinput156), .C1(n4995), .C2(keyinput174), 
        .A(n4901), .ZN(n4906) );
  AOI22_X1 U5451 ( .A1(n4929), .A2(keyinput149), .B1(keyinput176), .B2(n4904), 
        .ZN(n4903) );
  OAI221_X1 U5452 ( .B1(n4929), .B2(keyinput149), .C1(n4904), .C2(keyinput176), 
        .A(n4903), .ZN(n4905) );
  NOR4_X1 U5453 ( .A1(n4908), .A2(n4907), .A3(n4906), .A4(n4905), .ZN(n4921)
         );
  AOI22_X1 U5454 ( .A1(n4996), .A2(keyinput179), .B1(keyinput219), .B2(n4910), 
        .ZN(n4909) );
  OAI221_X1 U5455 ( .B1(n4996), .B2(keyinput179), .C1(n4910), .C2(keyinput219), 
        .A(n4909), .ZN(n4919) );
  AOI22_X1 U5456 ( .A1(n4912), .A2(keyinput171), .B1(keyinput134), .B2(n2645), 
        .ZN(n4911) );
  OAI221_X1 U5457 ( .B1(n4912), .B2(keyinput171), .C1(n2645), .C2(keyinput134), 
        .A(n4911), .ZN(n4918) );
  AOI22_X1 U5458 ( .A1(n4934), .A2(keyinput177), .B1(n4930), .B2(keyinput157), 
        .ZN(n4913) );
  OAI221_X1 U5459 ( .B1(n4934), .B2(keyinput177), .C1(n4930), .C2(keyinput157), 
        .A(n4913), .ZN(n4917) );
  AOI22_X1 U5460 ( .A1(n4915), .A2(keyinput211), .B1(n4972), .B2(keyinput241), 
        .ZN(n4914) );
  OAI221_X1 U5461 ( .B1(n4915), .B2(keyinput211), .C1(n4972), .C2(keyinput241), 
        .A(n4914), .ZN(n4916) );
  NOR4_X1 U5462 ( .A1(n4919), .A2(n4918), .A3(n4917), .A4(n4916), .ZN(n4920)
         );
  NAND4_X1 U5463 ( .A1(n4923), .A2(n4922), .A3(n4921), .A4(n4920), .ZN(n4924)
         );
  NOR4_X1 U5464 ( .A1(n4927), .A2(n4926), .A3(n4925), .A4(n4924), .ZN(n5059)
         );
  AOI22_X1 U5465 ( .A1(n4930), .A2(keyinput29), .B1(keyinput21), .B2(n4929), 
        .ZN(n4928) );
  OAI221_X1 U5466 ( .B1(n4930), .B2(keyinput29), .C1(n4929), .C2(keyinput21), 
        .A(n4928), .ZN(n4941) );
  AOI22_X1 U5467 ( .A1(n4932), .A2(keyinput5), .B1(n2334), .B2(keyinput13), 
        .ZN(n4931) );
  OAI221_X1 U5468 ( .B1(n4932), .B2(keyinput5), .C1(n2334), .C2(keyinput13), 
        .A(n4931), .ZN(n4940) );
  AOI22_X1 U5469 ( .A1(n4935), .A2(keyinput53), .B1(n4934), .B2(keyinput49), 
        .ZN(n4933) );
  OAI221_X1 U5470 ( .B1(n4935), .B2(keyinput53), .C1(n4934), .C2(keyinput49), 
        .A(n4933), .ZN(n4939) );
  XNOR2_X1 U5471 ( .A(REG1_REG_29__SCAN_IN), .B(keyinput45), .ZN(n4937) );
  XNOR2_X1 U5472 ( .A(IR_REG_16__SCAN_IN), .B(keyinput41), .ZN(n4936) );
  NAND2_X1 U5473 ( .A1(n4937), .A2(n4936), .ZN(n4938) );
  NOR4_X1 U5474 ( .A1(n4941), .A2(n4940), .A3(n4939), .A4(n4938), .ZN(n4990)
         );
  INV_X1 U5475 ( .A(ADDR_REG_1__SCAN_IN), .ZN(n4944) );
  AOI22_X1 U5476 ( .A1(n4944), .A2(keyinput85), .B1(n4943), .B2(keyinput65), 
        .ZN(n4942) );
  OAI221_X1 U5477 ( .B1(n4944), .B2(keyinput85), .C1(n4943), .C2(keyinput65), 
        .A(n4942), .ZN(n4955) );
  AOI22_X1 U5478 ( .A1(n2335), .A2(keyinput97), .B1(keyinput89), .B2(n4946), 
        .ZN(n4945) );
  OAI221_X1 U5479 ( .B1(n2335), .B2(keyinput97), .C1(n4946), .C2(keyinput89), 
        .A(n4945), .ZN(n4954) );
  INV_X1 U5480 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4948) );
  AOI22_X1 U5481 ( .A1(n4948), .A2(keyinput109), .B1(keyinput105), .B2(n4115), 
        .ZN(n4947) );
  OAI221_X1 U5482 ( .B1(n4948), .B2(keyinput109), .C1(n4115), .C2(keyinput105), 
        .A(n4947), .ZN(n4953) );
  AOI22_X1 U5483 ( .A1(n4951), .A2(keyinput60), .B1(keyinput32), .B2(n4950), 
        .ZN(n4949) );
  OAI221_X1 U5484 ( .B1(n4951), .B2(keyinput60), .C1(n4950), .C2(keyinput32), 
        .A(n4949), .ZN(n4952) );
  NOR4_X1 U5485 ( .A1(n4955), .A2(n4954), .A3(n4953), .A4(n4952), .ZN(n4989)
         );
  INV_X1 U5486 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4958) );
  AOI22_X1 U5487 ( .A1(n4958), .A2(keyinput40), .B1(n4957), .B2(keyinput52), 
        .ZN(n4956) );
  OAI221_X1 U5488 ( .B1(n4958), .B2(keyinput40), .C1(n4957), .C2(keyinput52), 
        .A(n4956), .ZN(n4970) );
  AOI22_X1 U5489 ( .A1(n3215), .A2(keyinput104), .B1(n4960), .B2(keyinput80), 
        .ZN(n4959) );
  OAI221_X1 U5490 ( .B1(n3215), .B2(keyinput104), .C1(n4960), .C2(keyinput80), 
        .A(n4959), .ZN(n4969) );
  AOI22_X1 U5491 ( .A1(n4963), .A2(keyinput72), .B1(keyinput68), .B2(n4962), 
        .ZN(n4961) );
  OAI221_X1 U5492 ( .B1(n4963), .B2(keyinput72), .C1(n4962), .C2(keyinput68), 
        .A(n4961), .ZN(n4968) );
  INV_X1 U5493 ( .A(ADDR_REG_9__SCAN_IN), .ZN(n4966) );
  AOI22_X1 U5494 ( .A1(n4966), .A2(keyinput121), .B1(n4965), .B2(keyinput125), 
        .ZN(n4964) );
  OAI221_X1 U5495 ( .B1(n4966), .B2(keyinput121), .C1(n4965), .C2(keyinput125), 
        .A(n4964), .ZN(n4967) );
  NOR4_X1 U5496 ( .A1(n4970), .A2(n4969), .A3(n4968), .A4(n4967), .ZN(n4988)
         );
  AOI22_X1 U5497 ( .A1(n4973), .A2(keyinput117), .B1(n4972), .B2(keyinput113), 
        .ZN(n4971) );
  OAI221_X1 U5498 ( .B1(n4973), .B2(keyinput117), .C1(n4972), .C2(keyinput113), 
        .A(n4971), .ZN(n4986) );
  AOI22_X1 U5499 ( .A1(n4976), .A2(keyinput44), .B1(n4975), .B2(keyinput36), 
        .ZN(n4974) );
  OAI221_X1 U5500 ( .B1(n4976), .B2(keyinput44), .C1(n4975), .C2(keyinput36), 
        .A(n4974), .ZN(n4985) );
  AOI22_X1 U5501 ( .A1(n4979), .A2(keyinput16), .B1(n4978), .B2(keyinput24), 
        .ZN(n4977) );
  OAI221_X1 U5502 ( .B1(n4979), .B2(keyinput16), .C1(n4978), .C2(keyinput24), 
        .A(n4977), .ZN(n4984) );
  AOI22_X1 U5503 ( .A1(n4982), .A2(keyinput62), .B1(keyinput54), .B2(n4981), 
        .ZN(n4980) );
  OAI221_X1 U5504 ( .B1(n4982), .B2(keyinput62), .C1(n4981), .C2(keyinput54), 
        .A(n4980), .ZN(n4983) );
  NOR4_X1 U5505 ( .A1(n4986), .A2(n4985), .A3(n4984), .A4(n4983), .ZN(n4987)
         );
  NAND4_X1 U5506 ( .A1(n4990), .A2(n4989), .A3(n4988), .A4(n4987), .ZN(n5058)
         );
  AOI22_X1 U5507 ( .A1(n4993), .A2(keyinput59), .B1(keyinput55), .B2(n4992), 
        .ZN(n4991) );
  OAI221_X1 U5508 ( .B1(n4993), .B2(keyinput59), .C1(n4992), .C2(keyinput55), 
        .A(n4991), .ZN(n5006) );
  AOI22_X1 U5509 ( .A1(n4996), .A2(keyinput51), .B1(n4995), .B2(keyinput46), 
        .ZN(n4994) );
  OAI221_X1 U5510 ( .B1(n4996), .B2(keyinput51), .C1(n4995), .C2(keyinput46), 
        .A(n4994), .ZN(n5005) );
  AOI22_X1 U5511 ( .A1(n4999), .A2(keyinput90), .B1(keyinput74), .B2(n4998), 
        .ZN(n4997) );
  OAI221_X1 U5512 ( .B1(n4999), .B2(keyinput90), .C1(n4998), .C2(keyinput74), 
        .A(n4997), .ZN(n5004) );
  INV_X1 U5513 ( .A(DATAI_30_), .ZN(n5001) );
  AOI22_X1 U5514 ( .A1(n5002), .A2(keyinput70), .B1(keyinput94), .B2(n5001), 
        .ZN(n5000) );
  OAI221_X1 U5515 ( .B1(n5002), .B2(keyinput70), .C1(n5001), .C2(keyinput94), 
        .A(n5000), .ZN(n5003) );
  NOR4_X1 U5516 ( .A1(n5006), .A2(n5005), .A3(n5004), .A4(n5003), .ZN(n5056)
         );
  AOI22_X1 U5517 ( .A1(n5009), .A2(keyinput107), .B1(keyinput110), .B2(n5008), 
        .ZN(n5007) );
  OAI221_X1 U5518 ( .B1(n5009), .B2(keyinput107), .C1(n5008), .C2(keyinput110), 
        .A(n5007), .ZN(n5022) );
  AOI22_X1 U5519 ( .A1(n5012), .A2(keyinput114), .B1(n5011), .B2(keyinput99), 
        .ZN(n5010) );
  OAI221_X1 U5520 ( .B1(n5012), .B2(keyinput114), .C1(n5011), .C2(keyinput99), 
        .A(n5010), .ZN(n5021) );
  AOI22_X1 U5521 ( .A1(n5015), .A2(keyinput103), .B1(keyinput0), .B2(n5014), 
        .ZN(n5013) );
  OAI221_X1 U5522 ( .B1(n5015), .B2(keyinput103), .C1(n5014), .C2(keyinput0), 
        .A(n5013), .ZN(n5020) );
  INV_X1 U5523 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n5017) );
  AOI22_X1 U5524 ( .A1(n5018), .A2(keyinput64), .B1(keyinput120), .B2(n5017), 
        .ZN(n5016) );
  OAI221_X1 U5525 ( .B1(n5018), .B2(keyinput64), .C1(n5017), .C2(keyinput120), 
        .A(n5016), .ZN(n5019) );
  NOR4_X1 U5526 ( .A1(n5022), .A2(n5021), .A3(n5020), .A4(n5019), .ZN(n5055)
         );
  INV_X1 U5527 ( .A(REG1_REG_25__SCAN_IN), .ZN(n5025) );
  AOI22_X1 U5528 ( .A1(n5025), .A2(keyinput14), .B1(keyinput7), .B2(n5024), 
        .ZN(n5023) );
  OAI221_X1 U5529 ( .B1(n5025), .B2(keyinput14), .C1(n5024), .C2(keyinput7), 
        .A(n5023), .ZN(n5037) );
  AOI22_X1 U5530 ( .A1(n5028), .A2(keyinput126), .B1(keyinput127), .B2(n5027), 
        .ZN(n5026) );
  OAI221_X1 U5531 ( .B1(n5028), .B2(keyinput126), .C1(n5027), .C2(keyinput127), 
        .A(n5026), .ZN(n5036) );
  AOI22_X1 U5532 ( .A1(n5031), .A2(keyinput10), .B1(n5030), .B2(keyinput15), 
        .ZN(n5029) );
  OAI221_X1 U5533 ( .B1(n5031), .B2(keyinput10), .C1(n5030), .C2(keyinput15), 
        .A(n5029), .ZN(n5035) );
  XNOR2_X1 U5534 ( .A(REG0_REG_25__SCAN_IN), .B(keyinput118), .ZN(n5033) );
  XNOR2_X1 U5535 ( .A(IR_REG_14__SCAN_IN), .B(keyinput124), .ZN(n5032) );
  NAND2_X1 U5536 ( .A1(n5033), .A2(n5032), .ZN(n5034) );
  NOR4_X1 U5537 ( .A1(n5037), .A2(n5036), .A3(n5035), .A4(n5034), .ZN(n5054)
         );
  AOI22_X1 U5538 ( .A1(n5040), .A2(keyinput42), .B1(keyinput26), .B2(n5039), 
        .ZN(n5038) );
  OAI221_X1 U5539 ( .B1(n5040), .B2(keyinput42), .C1(n5039), .C2(keyinput26), 
        .A(n5038), .ZN(n5052) );
  AOI22_X1 U5540 ( .A1(n5043), .A2(keyinput35), .B1(n5042), .B2(keyinput30), 
        .ZN(n5041) );
  OAI221_X1 U5541 ( .B1(n5043), .B2(keyinput35), .C1(n5042), .C2(keyinput30), 
        .A(n5041), .ZN(n5051) );
  XOR2_X1 U5542 ( .A(n5044), .B(keyinput38), .Z(n5047) );
  XNOR2_X1 U5543 ( .A(IR_REG_22__SCAN_IN), .B(keyinput11), .ZN(n5046) );
  XNOR2_X1 U5544 ( .A(IR_REG_6__SCAN_IN), .B(keyinput34), .ZN(n5045) );
  NAND3_X1 U5545 ( .A1(n5047), .A2(n5046), .A3(n5045), .ZN(n5050) );
  XNOR2_X1 U5546 ( .A(n5048), .B(keyinput47), .ZN(n5049) );
  NOR4_X1 U5547 ( .A1(n5052), .A2(n5051), .A3(n5050), .A4(n5049), .ZN(n5053)
         );
  NAND4_X1 U5548 ( .A1(n5056), .A2(n5055), .A3(n5054), .A4(n5053), .ZN(n5057)
         );
  NOR3_X1 U5549 ( .A1(n5059), .A2(n5058), .A3(n5057), .ZN(n5060) );
  NAND3_X1 U5550 ( .A1(n5062), .A2(n5061), .A3(n5060), .ZN(n5063) );
  XNOR2_X1 U5551 ( .A(n5064), .B(n5063), .ZN(U3229) );
endmodule

