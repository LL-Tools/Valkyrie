

module b22_C_SARLock_k_64_6 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6435, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208;

  AOI211_X1 U7184 ( .C1(n12532), .C2(n12531), .A(n14939), .B(n12530), .ZN(
        n12534) );
  NAND2_X1 U7185 ( .A1(n12811), .A2(n9704), .ZN(n12864) );
  AND2_X1 U7186 ( .A1(n13820), .A2(n11864), .ZN(n13800) );
  OAI21_X1 U7187 ( .B1(n10442), .B2(n10375), .A(n10374), .ZN(n10373) );
  INV_X2 U7188 ( .A(n12273), .ZN(n12277) );
  INV_X2 U7189 ( .A(n9155), .ZN(n9007) );
  CLKBUF_X2 U7190 ( .A(n8806), .Z(n6460) );
  CLKBUF_X1 U7191 ( .A(n8172), .Z(n8591) );
  XNOR2_X1 U7192 ( .A(n8774), .B(n8773), .ZN(n11907) );
  NAND2_X1 U7193 ( .A1(n8771), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8764) );
  BUF_X1 U7194 ( .A(n8119), .Z(n8577) );
  AND4_X1 U7195 ( .A1(n8063), .A2(n8062), .A3(n8061), .A4(n8060), .ZN(n14516)
         );
  INV_X1 U7196 ( .A(n8119), .ZN(n8590) );
  BUF_X2 U7197 ( .A(n7684), .Z(n6440) );
  OR2_X2 U7198 ( .A1(n8058), .A2(n8056), .ZN(n8462) );
  CLKBUF_X3 U7199 ( .A(n9465), .Z(n6439) );
  INV_X1 U7200 ( .A(n8252), .ZN(n8167) );
  AOI21_X1 U7201 ( .B1(n12370), .B2(n12383), .A(n12369), .ZN(n14923) );
  AND2_X1 U7202 ( .A1(n10147), .A2(n10146), .ZN(n11931) );
  NOR2_X1 U7203 ( .A1(n14271), .A2(n14272), .ZN(n14270) );
  NAND2_X1 U7204 ( .A1(n7226), .A2(n7227), .ZN(n12605) );
  NAND2_X1 U7206 ( .A1(n7597), .A2(n7596), .ZN(n11227) );
  CLKBUF_X2 U7207 ( .A(n8142), .Z(n8392) );
  NAND2_X2 U7208 ( .A1(n9190), .A2(n9191), .ZN(n8829) );
  CLKBUF_X3 U7209 ( .A(n8795), .Z(n6444) );
  NAND2_X1 U7211 ( .A1(n12843), .A2(n9686), .ZN(n9689) );
  INV_X2 U7212 ( .A(n9461), .ZN(n7737) );
  NOR3_X2 U7213 ( .A1(n13172), .A2(n13236), .A3(n6827), .ZN(n13098) );
  NAND2_X1 U7214 ( .A1(n13171), .A2(n13179), .ZN(n13172) );
  CLKBUF_X2 U7215 ( .A(n7009), .Z(n9469) );
  INV_X1 U7216 ( .A(n10598), .ZN(n13360) );
  INV_X1 U7217 ( .A(n8462), .ZN(n8493) );
  AND4_X1 U7218 ( .A1(n8837), .A2(n8836), .A3(n8835), .A4(n8834), .ZN(n10499)
         );
  NAND2_X1 U7219 ( .A1(n12753), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8774) );
  NAND2_X1 U7220 ( .A1(n7629), .A2(n7628), .ZN(n13273) );
  CLKBUF_X3 U7221 ( .A(n9616), .Z(n13190) );
  NAND2_X1 U7222 ( .A1(n7225), .A2(n7224), .ZN(n13835) );
  AND2_X1 U7223 ( .A1(n14089), .A2(n9834), .ZN(n13863) );
  INV_X1 U7224 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8303) );
  AND2_X1 U7225 ( .A1(n8100), .A2(n14556), .ZN(n6435) );
  OR2_X2 U7226 ( .A1(n12398), .A2(n12399), .ZN(n7124) );
  XNOR2_X2 U7227 ( .A(n6688), .B(n9653), .ZN(n11663) );
  NAND2_X2 U7228 ( .A1(n12509), .A2(n7388), .ZN(n12496) );
  NAND2_X2 U7229 ( .A1(n13852), .A2(n11859), .ZN(n13836) );
  INV_X1 U7230 ( .A(n8100), .ZN(n10398) );
  NAND2_X2 U7231 ( .A1(n11871), .A2(n11870), .ZN(n13944) );
  NAND3_X2 U7232 ( .A1(n8805), .A2(n7369), .A3(n8804), .ZN(n14954) );
  OR2_X1 U7233 ( .A1(n9155), .A2(n9758), .ZN(n8804) );
  OAI222_X1 U7234 ( .A1(P3_U3151), .A2(n9190), .B1(n14215), .B2(n12765), .C1(
        n12764), .C2(n14213), .ZN(P3_U3267) );
  NAND2_X2 U7235 ( .A1(n11906), .A2(n9651), .ZN(n6688) );
  AOI21_X2 U7236 ( .B1(n10445), .B2(n10444), .A(n10443), .ZN(n10442) );
  NAND2_X2 U7237 ( .A1(n6462), .A2(n6459), .ZN(n8142) );
  AOI22_X2 U7238 ( .A1(n6752), .A2(n6749), .B1(n6751), .B2(n6496), .ZN(n7580)
         );
  AND4_X2 U7239 ( .A1(n8113), .A2(n8112), .A3(n8111), .A4(n8110), .ZN(n14529)
         );
  INV_X1 U7240 ( .A(n9191), .ZN(n10118) );
  INV_X2 U7241 ( .A(n10396), .ZN(n14535) );
  NOR2_X2 U7242 ( .A1(n11277), .A2(n14793), .ZN(n11276) );
  NAND2_X2 U7243 ( .A1(n8718), .A2(n8717), .ZN(n8885) );
  NAND2_X2 U7244 ( .A1(n7490), .A2(n7489), .ZN(n7697) );
  OAI22_X2 U7245 ( .A1(n14179), .A2(n14178), .B1(P3_ADDR_REG_16__SCAN_IN), 
        .B2(n14464), .ZN(n14180) );
  CLKBUF_X1 U7246 ( .A(n6444), .Z(n6437) );
  NOR2_X2 U7247 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7540) );
  AOI21_X2 U7248 ( .B1(P3_REG1_REG_16__SCAN_IN), .B2(n14288), .A(n14289), .ZN(
        n12421) );
  BUF_X1 U7249 ( .A(n14248), .Z(n6438) );
  NAND2_X2 U7250 ( .A1(n8816), .A2(n14954), .ZN(n9240) );
  NAND2_X1 U7251 ( .A1(n7538), .A2(n7433), .ZN(n7684) );
  XNOR2_X2 U7252 ( .A(n8071), .B(n8067), .ZN(n10867) );
  BUF_X1 U7253 ( .A(n9461), .Z(n6441) );
  NAND2_X2 U7254 ( .A1(n8005), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7399) );
  NAND2_X2 U7255 ( .A1(n6507), .A2(n9302), .ZN(n9588) );
  OAI21_X2 U7256 ( .B1(n12605), .B2(n9044), .A(n9043), .ZN(n12592) );
  XNOR2_X1 U7257 ( .A(n11227), .B(n12891), .ZN(n11223) );
  AOI21_X2 U7258 ( .B1(n12603), .B2(n12606), .A(n12224), .ZN(n12590) );
  OAI21_X2 U7259 ( .B1(n9085), .B2(n7044), .A(n7043), .ZN(n9113) );
  CLKBUF_X1 U7260 ( .A(n8795), .Z(n6442) );
  CLKBUF_X3 U7261 ( .A(n8795), .Z(n6443) );
  AND2_X1 U7262 ( .A1(n11907), .A2(n8778), .ZN(n8795) );
  BUF_X2 U7263 ( .A(n7754), .Z(n6445) );
  BUF_X4 U7264 ( .A(n7754), .Z(n6446) );
  XNOR2_X2 U7265 ( .A(n10630), .B(n10645), .ZN(n10512) );
  NAND4_X4 U7267 ( .A1(n7728), .A2(n7727), .A3(n7726), .A4(n7725), .ZN(n12898)
         );
  NAND4_X4 U7268 ( .A1(n8077), .A2(n8076), .A3(n8075), .A4(n8074), .ZN(n8100)
         );
  NAND2_X2 U7269 ( .A1(n8172), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8075) );
  NAND2_X2 U7270 ( .A1(n9240), .A2(n12145), .ZN(n10236) );
  OR2_X2 U7271 ( .A1(n8053), .A2(n8325), .ZN(n8050) );
  XNOR2_X2 U7272 ( .A(n8105), .B(P1_IR_REG_2__SCAN_IN), .ZN(n13619) );
  XNOR2_X2 U7273 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8801) );
  XNOR2_X2 U7274 ( .A(n8764), .B(n8763), .ZN(n9190) );
  NOR2_X2 U7275 ( .A1(n10962), .A2(n10961), .ZN(n12350) );
  NOR2_X2 U7276 ( .A1(n10959), .A2(n10958), .ZN(n10962) );
  AND2_X2 U7277 ( .A1(n9576), .A2(n10947), .ZN(n14772) );
  AND2_X2 U7278 ( .A1(n9576), .A2(n12997), .ZN(n9303) );
  BUF_X2 U7280 ( .A(n10279), .Z(n6448) );
  XNOR2_X1 U7281 ( .A(n8824), .B(n15098), .ZN(n10279) );
  XNOR2_X2 U7282 ( .A(n8766), .B(n8765), .ZN(n9191) );
  XNOR2_X1 U7283 ( .A(n12330), .B(n12156), .ZN(n12115) );
  XNOR2_X2 U7284 ( .A(n8050), .B(P1_IR_REG_30__SCAN_IN), .ZN(n8058) );
  NAND2_X2 U7285 ( .A1(n8054), .A2(n14079), .ZN(n8056) );
  MUX2_X1 U7286 ( .A(n12475), .B(n12474), .S(n14963), .Z(n12479) );
  OAI21_X1 U7287 ( .B1(n13782), .B2(n13781), .A(n13780), .ZN(n13983) );
  NAND2_X1 U7288 ( .A1(n6900), .A2(n6535), .ZN(n13780) );
  AND2_X1 U7289 ( .A1(n7387), .A2(n7236), .ZN(n7235) );
  NOR2_X2 U7290 ( .A1(n13808), .A2(n13988), .ZN(n13794) );
  OAI21_X1 U7291 ( .B1(n13085), .B2(n13066), .A(n13082), .ZN(n13061) );
  NAND2_X1 U7292 ( .A1(n11664), .A2(n6687), .ZN(n11833) );
  AND2_X1 U7293 ( .A1(n9655), .A2(n7173), .ZN(n6687) );
  NAND2_X1 U7294 ( .A1(n11663), .A2(n9652), .ZN(n11664) );
  OR2_X1 U7295 ( .A1(n6688), .A2(n9654), .ZN(n9655) );
  NAND2_X1 U7296 ( .A1(n11189), .A2(n11188), .ZN(n11352) );
  NAND2_X1 U7297 ( .A1(n10685), .A2(n9610), .ZN(n10678) );
  AND2_X1 U7298 ( .A1(n10801), .A2(n8860), .ZN(n10790) );
  CLKBUF_X2 U7299 ( .A(P2_U3947), .Z(n6451) );
  CLKBUF_X2 U7300 ( .A(n9578), .Z(n13136) );
  NAND2_X1 U7301 ( .A1(n12146), .A2(n12153), .ZN(n7278) );
  INV_X1 U7302 ( .A(n12897), .ZN(n10424) );
  CLKBUF_X2 U7303 ( .A(n8492), .Z(n8589) );
  CLKBUF_X3 U7304 ( .A(n8833), .Z(n12089) );
  INV_X4 U7305 ( .A(n6486), .ZN(n6449) );
  NAND2_X2 U7306 ( .A1(n10407), .A2(n10867), .ZN(n10209) );
  NOR2_X1 U7307 ( .A1(n11907), .A2(n8778), .ZN(n8806) );
  INV_X1 U7309 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10204) );
  INV_X2 U7310 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  OAI21_X1 U7311 ( .B1(n14050), .B2(n14595), .A(n6604), .ZN(n13986) );
  OAI21_X1 U7312 ( .B1(n14050), .B2(n6712), .A(n6605), .ZN(n14051) );
  AND2_X1 U7313 ( .A1(n6506), .A2(n7372), .ZN(n9300) );
  OR2_X1 U7314 ( .A1(n6710), .A2(n11889), .ZN(n14050) );
  NAND2_X1 U7315 ( .A1(n12864), .A2(n6693), .ZN(n12769) );
  AOI21_X1 U7316 ( .B1(n7015), .B2(n14858), .A(n6596), .ZN(n7014) );
  NAND2_X1 U7317 ( .A1(n13787), .A2(n6706), .ZN(n13786) );
  NAND2_X1 U7318 ( .A1(n7020), .A2(n7019), .ZN(n12987) );
  OR2_X1 U7319 ( .A1(n7959), .A2(n9543), .ZN(n7020) );
  AOI21_X1 U7320 ( .B1(n12532), .B2(n7259), .A(n7257), .ZN(n7256) );
  OR2_X1 U7321 ( .A1(n9526), .A2(n9474), .ZN(n9484) );
  NAND2_X1 U7322 ( .A1(n13032), .A2(n7949), .ZN(n13014) );
  NAND2_X1 U7323 ( .A1(n13835), .A2(n6896), .ZN(n13816) );
  AOI21_X1 U7324 ( .B1(n13078), .B2(n7912), .A(n6730), .ZN(n13063) );
  NAND2_X1 U7325 ( .A1(n13862), .A2(n13861), .ZN(n7225) );
  NAND2_X1 U7326 ( .A1(n13905), .A2(n7360), .ZN(n13869) );
  AOI21_X1 U7327 ( .B1(n13013), .B2(n13012), .A(n7999), .ZN(n12960) );
  OAI21_X1 U7328 ( .B1(n7148), .B2(n7146), .A(n7145), .ZN(n7144) );
  NAND2_X1 U7329 ( .A1(n9170), .A2(n9169), .ZN(n9270) );
  NAND2_X1 U7330 ( .A1(n6643), .A2(n6640), .ZN(n13862) );
  NAND2_X1 U7331 ( .A1(n6998), .A2(n6997), .ZN(n13078) );
  AND2_X1 U7332 ( .A1(n9143), .A2(n9142), .ZN(n12680) );
  OR2_X1 U7333 ( .A1(n9168), .A2(n9167), .ZN(n9170) );
  NAND2_X1 U7334 ( .A1(n8617), .A2(n8573), .ZN(n13303) );
  NAND2_X1 U7335 ( .A1(n6715), .A2(n7880), .ZN(n13128) );
  NAND2_X1 U7336 ( .A1(n9153), .A2(n9152), .ZN(n9168) );
  NAND2_X1 U7337 ( .A1(n7152), .A2(n6511), .ZN(n13549) );
  AND2_X1 U7338 ( .A1(n9472), .A2(n9471), .ZN(n13196) );
  NAND2_X1 U7339 ( .A1(n8562), .A2(n8561), .ZN(n13980) );
  NAND2_X1 U7340 ( .A1(n13146), .A2(n7879), .ZN(n6715) );
  NAND2_X1 U7341 ( .A1(n13794), .A2(n14052), .ZN(n13774) );
  NAND2_X1 U7342 ( .A1(n9120), .A2(n9119), .ZN(n12691) );
  OR2_X1 U7343 ( .A1(n9151), .A2(n7378), .ZN(n9153) );
  OR2_X1 U7344 ( .A1(n8572), .A2(n8571), .ZN(n8617) );
  NAND2_X1 U7345 ( .A1(n6716), .A2(n7871), .ZN(n13146) );
  NAND2_X1 U7346 ( .A1(n13571), .A2(n13341), .ZN(n13505) );
  OAI22_X1 U7347 ( .A1(n9377), .A2(n6967), .B1(n9378), .B2(n6966), .ZN(n9382)
         );
  XNOR2_X1 U7348 ( .A(n8565), .B(n8564), .ZN(n13307) );
  NAND2_X1 U7349 ( .A1(n8519), .A2(n8518), .ZN(n13988) );
  NAND2_X1 U7350 ( .A1(n13167), .A2(n7870), .ZN(n6716) );
  OR2_X1 U7351 ( .A1(n14242), .A2(n6634), .ZN(n6635) );
  XNOR2_X1 U7352 ( .A(n7715), .B(n7714), .ZN(n11626) );
  OR2_X1 U7353 ( .A1(n8555), .A2(n11596), .ZN(n8556) );
  NAND2_X1 U7354 ( .A1(n6853), .A2(n6852), .ZN(n12561) );
  INV_X1 U7355 ( .A(n13074), .ZN(n13226) );
  AND2_X1 U7356 ( .A1(n7712), .A2(n7711), .ZN(n13038) );
  AND2_X1 U7357 ( .A1(n7704), .A2(n7703), .ZN(n13074) );
  NAND2_X1 U7358 ( .A1(n9116), .A2(n9115), .ZN(n9117) );
  NAND2_X1 U7359 ( .A1(n8467), .A2(n8466), .ZN(n14001) );
  AND2_X1 U7360 ( .A1(n13085), .A2(n13098), .ZN(n13087) );
  NAND2_X1 U7361 ( .A1(n7498), .A2(n7497), .ZN(n7710) );
  AND2_X1 U7362 ( .A1(n7525), .A2(n7524), .ZN(n13085) );
  OAI21_X1 U7363 ( .B1(n14261), .B2(n7299), .A(n7298), .ZN(n12426) );
  XNOR2_X1 U7364 ( .A(n7702), .B(n7701), .ZN(n11343) );
  NAND2_X1 U7365 ( .A1(n7699), .A2(n7698), .ZN(n7702) );
  NAND2_X1 U7366 ( .A1(n7300), .A2(n7301), .ZN(n7299) );
  INV_X1 U7367 ( .A(n13870), .ZN(n6450) );
  NAND2_X1 U7368 ( .A1(n11740), .A2(n7991), .ZN(n13181) );
  NOR2_X1 U7369 ( .A1(n14262), .A2(n14263), .ZN(n14261) );
  OR2_X1 U7370 ( .A1(n11738), .A2(n11741), .ZN(n11740) );
  AOI22_X1 U7371 ( .A1(n11923), .A2(n11922), .B1(n11921), .B2(n12318), .ZN(
        n12019) );
  NAND2_X1 U7372 ( .A1(n11442), .A2(n7199), .ZN(n11895) );
  NAND2_X1 U7373 ( .A1(n8384), .A2(n8383), .ZN(n13917) );
  OAI21_X1 U7374 ( .B1(n9060), .B2(n7025), .A(n7023), .ZN(n8753) );
  NAND2_X1 U7375 ( .A1(n10982), .A2(n6739), .ZN(n11152) );
  NAND2_X1 U7376 ( .A1(n7687), .A2(n7686), .ZN(n13246) );
  NAND2_X1 U7377 ( .A1(n11537), .A2(n11536), .ZN(n14494) );
  NAND2_X1 U7378 ( .A1(n7693), .A2(n7487), .ZN(n7490) );
  NOR2_X2 U7379 ( .A1(n11751), .A2(n13262), .ZN(n13171) );
  OAI21_X1 U7380 ( .B1(n11703), .B2(n7989), .A(n7988), .ZN(n11716) );
  NAND2_X1 U7381 ( .A1(n10983), .A2(n7072), .ZN(n10982) );
  NAND2_X1 U7382 ( .A1(n11352), .A2(n7356), .ZN(n11537) );
  NAND2_X1 U7383 ( .A1(n7673), .A2(n7672), .ZN(n13253) );
  NAND2_X1 U7384 ( .A1(n7486), .A2(n7485), .ZN(n7693) );
  OAI21_X1 U7385 ( .B1(n11551), .B2(n7080), .A(n7078), .ZN(n11703) );
  OR2_X1 U7386 ( .A1(n7484), .A2(n10535), .ZN(n7485) );
  XNOR2_X1 U7387 ( .A(n12364), .B(n12387), .ZN(n14914) );
  AND3_X1 U7388 ( .A1(n7110), .A2(n7112), .A3(P3_REG1_REG_11__SCAN_IN), .ZN(
        n14900) );
  NAND2_X1 U7389 ( .A1(n7785), .A2(n7018), .ZN(n11220) );
  NAND2_X1 U7390 ( .A1(n8330), .A2(n8329), .ZN(n14362) );
  NOR2_X1 U7391 ( .A1(n12363), .A2(n6817), .ZN(n12364) );
  NAND2_X1 U7392 ( .A1(n7652), .A2(n7651), .ZN(n13269) );
  OR2_X1 U7393 ( .A1(n12350), .A2(n7111), .ZN(n7110) );
  NAND2_X1 U7394 ( .A1(n7637), .A2(n7636), .ZN(n9640) );
  NAND2_X1 U7395 ( .A1(n7475), .A2(n7474), .ZN(n7676) );
  NAND2_X1 U7396 ( .A1(n8308), .A2(n8307), .ZN(n14241) );
  NAND2_X1 U7397 ( .A1(n7661), .A2(n7660), .ZN(n7475) );
  NAND2_X1 U7398 ( .A1(n8317), .A2(n8316), .ZN(n14336) );
  NAND2_X1 U7399 ( .A1(n7530), .A2(n7529), .ZN(n11730) );
  NAND2_X1 U7400 ( .A1(n7612), .A2(n7611), .ZN(n14842) );
  NAND2_X1 U7401 ( .A1(n8273), .A2(n8272), .ZN(n14373) );
  NAND2_X1 U7402 ( .A1(n6713), .A2(n8251), .ZN(n14502) );
  OAI22_X1 U7403 ( .A1(n10760), .A2(n6816), .B1(n6493), .B2(n10953), .ZN(
        n12335) );
  OAI21_X1 U7404 ( .B1(n9318), .B2(n6957), .A(n6956), .ZN(n9323) );
  OR2_X1 U7405 ( .A1(n7613), .A2(n7614), .ZN(n6778) );
  AND2_X1 U7406 ( .A1(n8236), .A2(n8235), .ZN(n11535) );
  AOI21_X1 U7407 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n15155), .A(n14108), .ZN(
        n14127) );
  NAND2_X1 U7408 ( .A1(n7214), .A2(n7216), .ZN(n7613) );
  NAND2_X1 U7409 ( .A1(n6702), .A2(n7439), .ZN(n7598) );
  INV_X1 U7410 ( .A(n9716), .ZN(n9709) );
  NAND2_X1 U7411 ( .A1(n6703), .A2(n7436), .ZN(n7590) );
  NAND2_X1 U7412 ( .A1(n8845), .A2(n8844), .ZN(n12146) );
  AND2_X1 U7413 ( .A1(n8149), .A2(n8148), .ZN(n14569) );
  NAND2_X2 U7414 ( .A1(n13767), .A2(n13952), .ZN(n14543) );
  AND2_X1 U7415 ( .A1(n8116), .A2(n10405), .ZN(n11330) );
  INV_X2 U7416 ( .A(n11931), .ZN(n11980) );
  AND4_X1 U7417 ( .A1(n8867), .A2(n8866), .A3(n8865), .A4(n8864), .ZN(n10902)
         );
  AND4_X1 U7418 ( .A1(n8881), .A2(n8880), .A3(n8879), .A4(n8878), .ZN(n10933)
         );
  NAND2_X1 U7419 ( .A1(n6487), .A2(n7061), .ZN(n12896) );
  NAND4_X1 U7420 ( .A1(n7742), .A2(n6488), .A3(n7741), .A4(n7740), .ZN(n12897)
         );
  NAND4_X1 U7421 ( .A1(n7733), .A2(n7732), .A3(n7731), .A4(n7730), .ZN(n12899)
         );
  NAND4_X1 U7422 ( .A1(n8823), .A2(n8822), .A3(n8821), .A4(n8820), .ZN(n12331)
         );
  INV_X1 U7423 ( .A(n14785), .ZN(n10825) );
  NAND2_X1 U7424 ( .A1(n8005), .A2(n7405), .ZN(n10947) );
  OR2_X1 U7425 ( .A1(n10385), .A2(n10295), .ZN(n10296) );
  NAND3_X1 U7426 ( .A1(n8107), .A2(n6895), .A3(n8106), .ZN(n11339) );
  INV_X1 U7427 ( .A(n8172), .ZN(n8157) );
  INV_X2 U7428 ( .A(n6486), .ZN(n13462) );
  AND3_X1 U7429 ( .A1(n8843), .A2(n8842), .A3(n8841), .ZN(n14976) );
  INV_X2 U7430 ( .A(n13463), .ZN(n13404) );
  NAND2_X1 U7431 ( .A1(n8058), .A2(n8056), .ZN(n8119) );
  NAND2_X2 U7432 ( .A1(n10210), .A2(n10209), .ZN(n13463) );
  NAND2_X4 U7433 ( .A1(n8584), .A2(n8099), .ZN(n8252) );
  NAND2_X1 U7434 ( .A1(n13302), .A2(n7723), .ZN(n9465) );
  NAND2_X1 U7435 ( .A1(n7723), .A2(n7724), .ZN(n9461) );
  AND2_X1 U7436 ( .A1(n6738), .A2(n6735), .ZN(n7723) );
  INV_X1 U7437 ( .A(n7724), .ZN(n13302) );
  XNOR2_X1 U7438 ( .A(n7407), .B(P2_IR_REG_20__SCAN_IN), .ZN(n9723) );
  INV_X1 U7439 ( .A(n10945), .ZN(n10407) );
  XNOR2_X1 U7440 ( .A(n8776), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8778) );
  MUX2_X1 U7441 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8052), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n8054) );
  NAND2_X1 U7442 ( .A1(n8070), .A2(n8669), .ZN(n10945) );
  NAND2_X1 U7443 ( .A1(n7517), .A2(n7720), .ZN(n7971) );
  XNOR2_X1 U7444 ( .A(n8096), .B(P1_IR_REG_19__SCAN_IN), .ZN(n13747) );
  MUX2_X1 U7445 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8068), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n8070) );
  NAND2_X1 U7446 ( .A1(n6872), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8766) );
  MUX2_X1 U7447 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7515), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n7517) );
  INV_X1 U7448 ( .A(n7663), .ZN(n7198) );
  NAND2_X1 U7449 ( .A1(n6498), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8071) );
  NAND2_X1 U7450 ( .A1(n7520), .A2(n7519), .ZN(n13311) );
  INV_X2 U7451 ( .A(n13306), .ZN(n6452) );
  OAI21_X1 U7452 ( .B1(n8013), .B2(n6697), .A(n6558), .ZN(n7520) );
  NAND4_X1 U7453 ( .A1(n7512), .A2(n6747), .A3(n6985), .A4(n6467), .ZN(n7720)
         );
  NOR2_X1 U7454 ( .A1(n7100), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n7099) );
  NOR2_X1 U7455 ( .A1(n7366), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n7365) );
  NAND2_X1 U7456 ( .A1(n6887), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7411) );
  OAI211_X1 U7457 ( .C1(n8802), .C2(n7293), .A(n8803), .B(n7292), .ZN(n10143)
         );
  NAND2_X1 U7458 ( .A1(n6888), .A2(n7410), .ZN(n7412) );
  AND2_X1 U7459 ( .A1(n10274), .A2(n8696), .ZN(n8851) );
  AND4_X1 U7460 ( .A1(n7389), .A2(n6990), .A3(n7390), .A4(n7568), .ZN(n6467)
         );
  AND2_X1 U7461 ( .A1(n6686), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14134) );
  AND2_X1 U7462 ( .A1(n8697), .A2(n7272), .ZN(n7269) );
  AND4_X1 U7463 ( .A1(n8692), .A2(n8691), .A3(n8690), .A4(n8689), .ZN(n7377)
         );
  AND4_X1 U7464 ( .A1(n8694), .A2(n8854), .A3(n8693), .A4(n8926), .ZN(n8695)
         );
  INV_X1 U7465 ( .A(P2_RD_REG_SCAN_IN), .ZN(n6699) );
  INV_X1 U7466 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n6700) );
  INV_X1 U7467 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8697) );
  INV_X1 U7468 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6889) );
  NOR2_X2 U7469 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n10274) );
  INV_X1 U7470 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8854) );
  INV_X1 U7471 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8144) );
  NOR2_X1 U7472 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n8696) );
  INV_X1 U7473 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8048) );
  INV_X1 U7474 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8183) );
  INV_X4 U7475 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7476 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8269) );
  NOR2_X1 U7477 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8692) );
  NOR2_X1 U7478 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n8691) );
  NOR2_X1 U7479 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n8690) );
  NOR2_X1 U7480 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8689) );
  INV_X1 U7481 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n12948) );
  INV_X1 U7482 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8926) );
  NOR2_X1 U7483 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7389) );
  NOR2_X1 U7484 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7390) );
  NOR2_X1 U7485 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n6990) );
  NOR2_X1 U7486 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7621) );
  NOR2_X1 U7487 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7505) );
  INV_X1 U7488 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8028) );
  INV_X1 U7489 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7509) );
  INV_X4 U7490 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  XNOR2_X1 U7491 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n14133) );
  INV_X1 U7492 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7568) );
  AND3_X4 U7493 ( .A1(n8087), .A2(n8086), .A3(n8085), .ZN(n14556) );
  NAND2_X4 U7494 ( .A1(n8079), .A2(n6629), .ZN(n8685) );
  NAND2_X2 U7495 ( .A1(n13860), .A2(n13845), .ZN(n13842) );
  NAND2_X1 U7496 ( .A1(n13905), .A2(n6455), .ZN(n6453) );
  AND2_X2 U7497 ( .A1(n6453), .A2(n6454), .ZN(n13873) );
  OR2_X1 U7498 ( .A1(n6450), .A2(n13871), .ZN(n6454) );
  AND2_X1 U7499 ( .A1(n7360), .A2(n13870), .ZN(n6455) );
  CLKBUF_X1 U7500 ( .A(n6704), .Z(n6456) );
  INV_X1 U7501 ( .A(n6435), .ZN(n6457) );
  BUF_X1 U7502 ( .A(n8051), .Z(n8079) );
  NOR2_X2 U7503 ( .A1(n12592), .A2(n12591), .ZN(n12595) );
  NAND2_X1 U7504 ( .A1(n10398), .A2(n13479), .ZN(n10403) );
  NOR2_X2 U7505 ( .A1(n10947), .A2(n9723), .ZN(n6953) );
  AND2_X1 U7506 ( .A1(n11907), .A2(n12760), .ZN(n8833) );
  OAI222_X1 U7507 ( .A1(P3_U3151), .A2(n11907), .B1(n14215), .B2(n11914), .C1(
        n12085), .C2(n14213), .ZN(P3_U3265) );
  MUX2_X2 U7508 ( .A(n13977), .B(n14046), .S(n14597), .Z(n13978) );
  MUX2_X2 U7509 ( .A(n14047), .B(n14046), .S(n14589), .Z(n14048) );
  INV_X1 U7510 ( .A(n7433), .ZN(n6458) );
  INV_X2 U7511 ( .A(n7433), .ZN(n6459) );
  AND2_X4 U7512 ( .A1(n7412), .A2(n7411), .ZN(n7433) );
  AOI21_X4 U7513 ( .B1(n12708), .B2(n12047), .A(n12549), .ZN(n12541) );
  OR2_X4 U7514 ( .A1(n10209), .A2(n10042), .ZN(n6486) );
  OR2_X1 U7515 ( .A1(n8058), .A2(n8056), .ZN(n6461) );
  NAND2_X1 U7516 ( .A1(n8685), .A2(n8684), .ZN(n6462) );
  NAND2_X1 U7517 ( .A1(n8685), .A2(n8684), .ZN(n6463) );
  INV_X1 U7518 ( .A(n8172), .ZN(n6464) );
  NOR2_X2 U7519 ( .A1(n13934), .A2(n13917), .ZN(n13916) );
  AOI21_X2 U7520 ( .B1(n13803), .B2(n14519), .A(n13802), .ZN(n13992) );
  NAND2_X1 U7521 ( .A1(n7359), .A2(n8058), .ZN(n8492) );
  NAND2_X2 U7522 ( .A1(n6946), .A2(n6945), .ZN(n13808) );
  NOR2_X4 U7523 ( .A1(n13842), .A2(n13827), .ZN(n6946) );
  NOR2_X2 U7524 ( .A1(n13956), .A2(n14034), .ZN(n6944) );
  NAND2_X1 U7525 ( .A1(n7471), .A2(n10031), .ZN(n7474) );
  NOR2_X1 U7526 ( .A1(n12680), .A2(n12309), .ZN(n12267) );
  NAND2_X1 U7527 ( .A1(n6831), .A2(n12179), .ZN(n11375) );
  NAND2_X1 U7528 ( .A1(n13014), .A2(n7950), .ZN(n7959) );
  OR2_X1 U7529 ( .A1(n13209), .A2(n12814), .ZN(n7950) );
  INV_X1 U7530 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6986) );
  NOR2_X1 U7531 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n6987) );
  NOR2_X1 U7532 ( .A1(n11642), .A2(n6901), .ZN(n6637) );
  NAND2_X1 U7533 ( .A1(n6796), .A2(n6801), .ZN(n8555) );
  NAND2_X1 U7534 ( .A1(n6800), .A2(n6797), .ZN(n6796) );
  AND2_X1 U7535 ( .A1(n6806), .A2(n6798), .ZN(n6797) );
  INV_X1 U7536 ( .A(n6803), .ZN(n6798) );
  NOR2_X1 U7537 ( .A1(n9484), .A2(n9477), .ZN(n9478) );
  NAND2_X1 U7538 ( .A1(n13311), .A2(n7971), .ZN(n7538) );
  NOR2_X1 U7539 ( .A1(n13749), .A2(n6899), .ZN(n6898) );
  INV_X1 U7540 ( .A(n11881), .ZN(n6899) );
  NAND2_X1 U7541 ( .A1(n13816), .A2(n7221), .ZN(n13806) );
  NOR2_X1 U7542 ( .A1(n7223), .A2(n7222), .ZN(n7221) );
  INV_X1 U7543 ( .A(n11879), .ZN(n7222) );
  INV_X1 U7544 ( .A(n8574), .ZN(n8147) );
  NAND2_X1 U7545 ( .A1(n9317), .A2(n9320), .ZN(n6956) );
  NOR2_X1 U7546 ( .A1(n9320), .A2(n9317), .ZN(n6957) );
  INV_X1 U7547 ( .A(n7318), .ZN(n7317) );
  NAND2_X1 U7548 ( .A1(n9419), .A2(n6965), .ZN(n6964) );
  AOI21_X1 U7549 ( .B1(n6779), .B2(n6776), .A(n6775), .ZN(n6774) );
  INV_X1 U7550 ( .A(n7448), .ZN(n6776) );
  INV_X1 U7551 ( .A(n7206), .ZN(n6775) );
  AOI21_X1 U7552 ( .B1(n7209), .B2(n7211), .A(n7207), .ZN(n7206) );
  INV_X1 U7553 ( .A(n6779), .ZN(n6777) );
  NAND2_X1 U7554 ( .A1(n6771), .A2(n6774), .ZN(n7640) );
  OR2_X1 U7555 ( .A1(n7613), .A2(n6777), .ZN(n6771) );
  NAND2_X1 U7556 ( .A1(n7556), .A2(n7425), .ZN(n6752) );
  INV_X1 U7557 ( .A(n7557), .ZN(n7425) );
  AOI21_X1 U7558 ( .B1(n12027), .B2(n11944), .A(n6907), .ZN(n6906) );
  INV_X1 U7559 ( .A(n11998), .ZN(n6907) );
  AND2_X1 U7560 ( .A1(n12348), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n12349) );
  NOR2_X1 U7561 ( .A1(n12394), .A2(n12395), .ZN(n12396) );
  NAND2_X1 U7562 ( .A1(n7239), .A2(n7237), .ZN(n7236) );
  INV_X1 U7563 ( .A(n9150), .ZN(n7237) );
  NAND2_X1 U7564 ( .A1(n7265), .A2(n12528), .ZN(n7264) );
  NAND2_X1 U7565 ( .A1(n7265), .A2(n9111), .ZN(n7263) );
  OR2_X1 U7566 ( .A1(n12557), .A2(n12047), .ZN(n12247) );
  NAND2_X1 U7567 ( .A1(n9206), .A2(n7274), .ZN(n6872) );
  NAND2_X1 U7568 ( .A1(n9113), .A2(n9112), .ZN(n9116) );
  INV_X1 U7569 ( .A(n7024), .ZN(n7023) );
  OAI21_X1 U7570 ( .B1(n9059), .B2(n7025), .A(P1_DATAO_REG_20__SCAN_IN), .ZN(
        n7024) );
  INV_X1 U7571 ( .A(n8752), .ZN(n7025) );
  NAND2_X1 U7572 ( .A1(n7058), .A2(n7056), .ZN(n8734) );
  AOI21_X1 U7573 ( .B1(n6586), .B2(n8730), .A(n7057), .ZN(n7056) );
  INV_X1 U7574 ( .A(n8733), .ZN(n7057) );
  XNOR2_X1 U7575 ( .A(n12772), .B(n12958), .ZN(n9543) );
  NAND2_X1 U7576 ( .A1(n13118), .A2(n12797), .ZN(n7007) );
  INV_X1 U7577 ( .A(n13150), .ZN(n7085) );
  OR2_X1 U7578 ( .A1(n11223), .A2(n7076), .ZN(n7075) );
  INV_X1 U7579 ( .A(n7983), .ZN(n7076) );
  NAND2_X1 U7580 ( .A1(n11239), .A2(n7783), .ZN(n7785) );
  OR3_X1 U7581 ( .A1(n9718), .A2(n8032), .A3(n14764), .ZN(n10809) );
  INV_X1 U7582 ( .A(n13297), .ZN(n6737) );
  INV_X1 U7583 ( .A(n7142), .ZN(n7141) );
  OAI21_X1 U7584 ( .B1(n7144), .B2(n7147), .A(n13401), .ZN(n7142) );
  AOI21_X1 U7585 ( .B1(n7150), .B2(n13539), .A(n7149), .ZN(n7148) );
  INV_X1 U7586 ( .A(n13432), .ZN(n7149) );
  NAND2_X1 U7587 ( .A1(n10231), .A2(n13446), .ZN(n10706) );
  AND2_X1 U7588 ( .A1(n6770), .A2(n8597), .ZN(n6766) );
  NAND3_X1 U7589 ( .A1(n6784), .A2(n6782), .A3(n6781), .ZN(n7498) );
  NOR2_X1 U7590 ( .A1(n6786), .A2(n6783), .ZN(n6782) );
  NAND2_X1 U7591 ( .A1(n7470), .A2(n7469), .ZN(n7661) );
  AND2_X1 U7592 ( .A1(n7474), .A2(n7473), .ZN(n7660) );
  NAND2_X1 U7593 ( .A1(n6778), .A2(n7448), .ZN(n7620) );
  NAND2_X1 U7594 ( .A1(n6752), .A2(n7427), .ZN(n7564) );
  NAND2_X1 U7595 ( .A1(n8089), .A2(n7532), .ZN(n7535) );
  NAND2_X1 U7596 ( .A1(n10896), .A2(n10895), .ZN(n12007) );
  NAND2_X1 U7597 ( .A1(n12285), .A2(n7049), .ZN(n7048) );
  NOR2_X1 U7598 ( .A1(n12129), .A2(n12130), .ZN(n7049) );
  AND4_X1 U7599 ( .A1(n9138), .A2(n9137), .A3(n9136), .A4(n9135), .ZN(n12032)
         );
  AND3_X1 U7600 ( .A1(n9071), .A2(n9070), .A3(n9069), .ZN(n12058) );
  AND4_X1 U7601 ( .A1(n8904), .A2(n8903), .A3(n8902), .A4(n8901), .ZN(n10935)
         );
  XNOR2_X1 U7602 ( .A(n6624), .B(n6623), .ZN(n10516) );
  INV_X1 U7603 ( .A(n10955), .ZN(n10956) );
  NOR2_X1 U7604 ( .A1(n12335), .A2(n7282), .ZN(n12336) );
  AND2_X1 U7605 ( .A1(n12348), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7282) );
  XNOR2_X1 U7606 ( .A(n12396), .B(n12412), .ZN(n14268) );
  XNOR2_X1 U7607 ( .A(n12426), .B(n12425), .ZN(n12404) );
  NOR2_X1 U7608 ( .A1(n12403), .A2(n12404), .ZN(n12429) );
  NAND2_X1 U7609 ( .A1(n7240), .A2(n7239), .ZN(n12480) );
  AOI21_X1 U7610 ( .B1(n7245), .B2(n7243), .A(n6563), .ZN(n7242) );
  AOI21_X1 U7611 ( .B1(n7229), .B2(n7232), .A(n6539), .ZN(n7227) );
  INV_X1 U7612 ( .A(n9017), .ZN(n7232) );
  INV_X1 U7613 ( .A(n8968), .ZN(n12083) );
  INV_X1 U7614 ( .A(n8829), .ZN(n9193) );
  AND2_X1 U7615 ( .A1(n6938), .A2(n9217), .ZN(n9802) );
  INV_X1 U7616 ( .A(n12895), .ZN(n10690) );
  NAND2_X1 U7617 ( .A1(n11258), .A2(n9635), .ZN(n11442) );
  NOR2_X1 U7618 ( .A1(n9727), .A2(n14764), .ZN(n9734) );
  NAND2_X1 U7619 ( .A1(n6445), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7740) );
  NAND2_X1 U7620 ( .A1(n12969), .A2(n9528), .ZN(n12984) );
  AND2_X1 U7621 ( .A1(n13209), .A2(n13035), .ZN(n7999) );
  AND2_X1 U7622 ( .A1(n7947), .A2(n7946), .ZN(n12814) );
  AOI21_X1 U7623 ( .B1(n7000), .B2(n7002), .A(n6554), .ZN(n6997) );
  NAND2_X1 U7624 ( .A1(n7994), .A2(n6494), .ZN(n13147) );
  NOR2_X1 U7625 ( .A1(n11718), .A2(n7013), .ZN(n7012) );
  INV_X1 U7626 ( .A(n7844), .ZN(n7013) );
  AOI21_X1 U7627 ( .B1(n7065), .B2(n7067), .A(n11040), .ZN(n7064) );
  INV_X1 U7628 ( .A(n12896), .ZN(n11273) );
  AND2_X1 U7629 ( .A1(n7099), .A2(n7516), .ZN(n6747) );
  INV_X1 U7630 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7516) );
  NAND2_X1 U7631 ( .A1(n7397), .A2(n7402), .ZN(n8005) );
  AOI21_X1 U7632 ( .B1(n13531), .B2(n13530), .A(n13364), .ZN(n13484) );
  AND2_X1 U7633 ( .A1(n6499), .A2(n7160), .ZN(n7157) );
  NAND2_X1 U7634 ( .A1(n13349), .A2(n7159), .ZN(n7158) );
  INV_X1 U7635 ( .A(n7368), .ZN(n7159) );
  AND2_X1 U7636 ( .A1(n8326), .A2(n8065), .ZN(n7163) );
  INV_X1 U7637 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8065) );
  XNOR2_X1 U7638 ( .A(n8645), .B(n13790), .ZN(n13749) );
  INV_X1 U7639 ( .A(n14052), .ZN(n8645) );
  NAND2_X1 U7640 ( .A1(n13806), .A2(n11880), .ZN(n13787) );
  AND2_X1 U7641 ( .A1(n11860), .A2(n11876), .ZN(n7224) );
  AOI21_X1 U7642 ( .B1(n6637), .B2(n14235), .A(n6552), .ZN(n6636) );
  INV_X1 U7643 ( .A(n11758), .ZN(n11764) );
  INV_X1 U7644 ( .A(n6637), .ZN(n6634) );
  XNOR2_X1 U7645 ( .A(n8555), .B(n7503), .ZN(n11845) );
  AND2_X1 U7646 ( .A1(n8066), .A2(n8067), .ZN(n7347) );
  NOR2_X1 U7647 ( .A1(n14143), .A2(n14144), .ZN(n14148) );
  NAND2_X1 U7648 ( .A1(n6666), .A2(n15142), .ZN(n6665) );
  OR2_X1 U7649 ( .A1(n14896), .A2(n14897), .ZN(n7281) );
  XNOR2_X1 U7650 ( .A(n12336), .B(n12351), .ZN(n14896) );
  INV_X1 U7651 ( .A(n12680), .ZN(n12503) );
  INV_X1 U7652 ( .A(n9738), .ZN(n7180) );
  NAND2_X1 U7653 ( .A1(n13307), .A2(n8381), .ZN(n8562) );
  NAND2_X1 U7654 ( .A1(n6884), .A2(n6885), .ZN(n14394) );
  NAND2_X1 U7655 ( .A1(n6881), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6880) );
  NOR2_X1 U7656 ( .A1(n14393), .A2(n6883), .ZN(n6882) );
  INV_X1 U7657 ( .A(n6885), .ZN(n6883) );
  NAND2_X1 U7658 ( .A1(n9323), .A2(n9324), .ZN(n9322) );
  INV_X1 U7659 ( .A(n8136), .ZN(n7313) );
  INV_X1 U7660 ( .A(n7324), .ZN(n7320) );
  NOR2_X1 U7661 ( .A1(n7324), .A2(n7322), .ZN(n7321) );
  NAND2_X1 U7662 ( .A1(n8310), .A2(n7309), .ZN(n7308) );
  INV_X1 U7663 ( .A(n8309), .ZN(n7309) );
  NAND2_X1 U7664 ( .A1(n7317), .A2(n7319), .ZN(n7316) );
  INV_X1 U7665 ( .A(n9388), .ZN(n6954) );
  NOR2_X1 U7666 ( .A1(n9391), .A2(n9388), .ZN(n6955) );
  NAND2_X1 U7667 ( .A1(n6981), .A2(n9400), .ZN(n6980) );
  AND2_X1 U7668 ( .A1(n6964), .A2(n9416), .ZN(n6959) );
  AND2_X1 U7669 ( .A1(n6964), .A2(n9412), .ZN(n6961) );
  INV_X1 U7670 ( .A(n9419), .ZN(n6963) );
  AND2_X1 U7671 ( .A1(n7209), .A2(n6780), .ZN(n6779) );
  NAND2_X1 U7672 ( .A1(n7614), .A2(n7448), .ZN(n6780) );
  NAND2_X1 U7673 ( .A1(n9425), .A2(n6972), .ZN(n6971) );
  OR2_X1 U7674 ( .A1(n12516), .A2(n12032), .ZN(n12262) );
  AND2_X1 U7675 ( .A1(n6515), .A2(n8761), .ZN(n7274) );
  AOI21_X1 U7676 ( .B1(n6652), .B2(n11872), .A(n6544), .ZN(n6651) );
  NAND2_X1 U7677 ( .A1(n6647), .A2(n6650), .ZN(n6642) );
  AOI21_X1 U7678 ( .B1(n6894), .B2(n6891), .A(n6545), .ZN(n6890) );
  INV_X1 U7679 ( .A(n6490), .ZN(n6891) );
  INV_X1 U7680 ( .A(n6894), .ZN(n6892) );
  NOR2_X1 U7681 ( .A1(n6892), .A2(n6645), .ZN(n6644) );
  INV_X1 U7682 ( .A(n6647), .ZN(n6645) );
  NAND2_X1 U7683 ( .A1(n11786), .A2(n7358), .ZN(n6704) );
  AND2_X1 U7684 ( .A1(n11785), .A2(n11850), .ZN(n7358) );
  NOR2_X1 U7685 ( .A1(n7713), .A2(n11581), .ZN(n6803) );
  NAND2_X1 U7686 ( .A1(n6794), .A2(n7495), .ZN(n7496) );
  AND2_X1 U7687 ( .A1(n7495), .A2(n6793), .ZN(n6792) );
  AND2_X1 U7688 ( .A1(n7476), .A2(n7681), .ZN(n7477) );
  NAND2_X1 U7689 ( .A1(n7453), .A2(n15157), .ZN(n7456) );
  INV_X1 U7690 ( .A(n7574), .ZN(n7431) );
  INV_X1 U7691 ( .A(n7430), .ZN(n7213) );
  OAI21_X1 U7692 ( .B1(n14139), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n14094), .ZN(
        n14095) );
  NAND2_X1 U7693 ( .A1(n11926), .A2(n12317), .ZN(n6929) );
  INV_X1 U7694 ( .A(n6923), .ZN(n6917) );
  INV_X1 U7695 ( .A(n6920), .ZN(n6915) );
  INV_X1 U7696 ( .A(n12101), .ZN(n6851) );
  NAND2_X1 U7697 ( .A1(n6620), .A2(n6619), .ZN(n12284) );
  AND2_X1 U7698 ( .A1(n12106), .A2(n7050), .ZN(n12285) );
  NAND2_X1 U7699 ( .A1(n12665), .A2(n12107), .ZN(n7050) );
  NOR2_X1 U7700 ( .A1(n12385), .A2(n12384), .ZN(n12386) );
  AND2_X1 U7701 ( .A1(n12485), .A2(n6509), .ZN(n7239) );
  NAND2_X1 U7702 ( .A1(n12141), .A2(n12145), .ZN(n10151) );
  NOR2_X1 U7703 ( .A1(n10546), .A2(n12334), .ZN(n12141) );
  INV_X1 U7704 ( .A(n7239), .ZN(n7238) );
  INV_X1 U7705 ( .A(n7264), .ZN(n7258) );
  NAND2_X1 U7706 ( .A1(n7263), .A2(n12507), .ZN(n7261) );
  NAND2_X1 U7707 ( .A1(n12262), .A2(n12263), .ZN(n12256) );
  INV_X1 U7708 ( .A(n6838), .ZN(n6834) );
  INV_X1 U7709 ( .A(n12259), .ZN(n6843) );
  NOR2_X1 U7710 ( .A1(n12528), .A2(n12133), .ZN(n6842) );
  OR2_X1 U7711 ( .A1(n12714), .A2(n11971), .ZN(n12243) );
  INV_X1 U7712 ( .A(n12595), .ZN(n7255) );
  OR2_X1 U7713 ( .A1(n12745), .A2(n11778), .ZN(n12216) );
  AOI21_X1 U7714 ( .B1(n11584), .B2(n12205), .A(n9251), .ZN(n11658) );
  INV_X1 U7715 ( .A(n6606), .ZN(n7039) );
  INV_X1 U7716 ( .A(n7031), .ZN(n7030) );
  OAI21_X1 U7717 ( .B1(n8744), .B2(n7032), .A(n8747), .ZN(n7031) );
  INV_X1 U7718 ( .A(n8745), .ZN(n7032) );
  INV_X1 U7719 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8694) );
  NAND2_X1 U7720 ( .A1(n8734), .A2(n10076), .ZN(n8735) );
  AND2_X1 U7721 ( .A1(n9858), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8730) );
  INV_X1 U7722 ( .A(n8894), .ZN(n8721) );
  NAND2_X1 U7723 ( .A1(n10677), .A2(n9615), .ZN(n7195) );
  NOR2_X1 U7724 ( .A1(n7921), .A2(n12822), .ZN(n7930) );
  INV_X1 U7725 ( .A(n7998), .ZN(n7091) );
  NOR2_X1 U7726 ( .A1(n7998), .A2(n6471), .ZN(n7090) );
  INV_X1 U7727 ( .A(n13219), .ZN(n9433) );
  OR2_X1 U7728 ( .A1(n6828), .A2(n13118), .ZN(n6827) );
  INV_X1 U7729 ( .A(n7987), .ZN(n7079) );
  INV_X1 U7730 ( .A(n11268), .ZN(n6996) );
  NAND2_X1 U7731 ( .A1(n14772), .A2(n10893), .ZN(n9596) );
  AOI21_X1 U7732 ( .B1(n7074), .B2(n11238), .A(n6534), .ZN(n7073) );
  OAI21_X1 U7733 ( .B1(n8005), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8029) );
  AND2_X1 U7734 ( .A1(n7197), .A2(n7504), .ZN(n6988) );
  INV_X1 U7735 ( .A(n7151), .ZN(n7150) );
  OAI21_X1 U7736 ( .B1(n13539), .B2(n13540), .A(n13382), .ZN(n7151) );
  INV_X1 U7737 ( .A(n11866), .ZN(n7349) );
  NAND2_X1 U7738 ( .A1(n6707), .A2(n6705), .ZN(n11867) );
  AOI21_X1 U7739 ( .B1(n6708), .B2(n7353), .A(n6706), .ZN(n6705) );
  AND2_X1 U7740 ( .A1(n6648), .A2(n13909), .ZN(n6647) );
  NAND2_X1 U7741 ( .A1(n6651), .A2(n6649), .ZN(n6648) );
  INV_X1 U7742 ( .A(n6652), .ZN(n6649) );
  INV_X1 U7743 ( .A(n6651), .ZN(n6650) );
  AND2_X1 U7744 ( .A1(n8406), .A2(n11855), .ZN(n8403) );
  NAND2_X1 U7745 ( .A1(n6646), .A2(n6651), .ZN(n13907) );
  NAND2_X1 U7746 ( .A1(n13944), .A2(n6652), .ZN(n6646) );
  NAND2_X1 U7747 ( .A1(n14336), .A2(n13330), .ZN(n8340) );
  OR2_X1 U7748 ( .A1(n14336), .A2(n13330), .ZN(n11762) );
  INV_X1 U7749 ( .A(n8566), .ZN(n6769) );
  INV_X1 U7750 ( .A(n8564), .ZN(n6770) );
  INV_X1 U7751 ( .A(n7709), .ZN(n6806) );
  OR2_X1 U7752 ( .A1(n7697), .A2(n6790), .ZN(n6784) );
  INV_X1 U7753 ( .A(n6792), .ZN(n6790) );
  NAND2_X1 U7754 ( .A1(n7697), .A2(n6484), .ZN(n6781) );
  OAI211_X1 U7755 ( .C1(n7676), .C2(n6757), .A(n7483), .B(n6754), .ZN(n7486)
         );
  AND2_X1 U7756 ( .A1(n6759), .A2(n6763), .ZN(n6758) );
  OR2_X1 U7757 ( .A1(n7482), .A2(n10535), .ZN(n6763) );
  NAND2_X1 U7758 ( .A1(n6761), .A2(n6760), .ZN(n6759) );
  INV_X1 U7759 ( .A(n7477), .ZN(n6760) );
  NAND2_X1 U7760 ( .A1(n7464), .A2(n7463), .ZN(n7654) );
  NAND2_X1 U7761 ( .A1(n6773), .A2(n6772), .ZN(n7464) );
  AND2_X1 U7762 ( .A1(n7469), .A2(n7468), .ZN(n7653) );
  NAND2_X1 U7763 ( .A1(n7458), .A2(SI_15_), .ZN(n7645) );
  AOI21_X1 U7764 ( .B1(n7443), .B2(n7217), .A(n6551), .ZN(n7216) );
  NAND2_X1 U7765 ( .A1(n7598), .A2(n7215), .ZN(n7214) );
  INV_X1 U7766 ( .A(n7581), .ZN(n7434) );
  XNOR2_X1 U7767 ( .A(n7432), .B(SI_6_), .ZN(n7574) );
  INV_X1 U7768 ( .A(n7565), .ZN(n7428) );
  XNOR2_X1 U7769 ( .A(n7429), .B(SI_5_), .ZN(n7565) );
  NAND2_X1 U7770 ( .A1(n6701), .A2(n7424), .ZN(n7556) );
  XNOR2_X1 U7771 ( .A(P3_ADDR_REG_4__SCAN_IN), .B(n14095), .ZN(n14130) );
  NOR2_X1 U7772 ( .A1(n14163), .A2(n14162), .ZN(n14108) );
  NAND2_X1 U7773 ( .A1(n6926), .A2(n6929), .ZN(n6925) );
  NAND2_X1 U7774 ( .A1(n12053), .A2(n6927), .ZN(n6926) );
  NAND2_X1 U7775 ( .A1(n12018), .A2(n6928), .ZN(n6927) );
  NAND2_X1 U7776 ( .A1(n10491), .A2(n6930), .ZN(n10896) );
  AND2_X1 U7777 ( .A1(n6931), .A2(n10490), .ZN(n6930) );
  NAND2_X1 U7778 ( .A1(n6936), .A2(n6937), .ZN(n14880) );
  AND2_X1 U7779 ( .A1(n10918), .A2(n10919), .ZN(n6936) );
  OAI21_X1 U7780 ( .B1(n11514), .B2(n6610), .A(n6556), .ZN(n6934) );
  NAND2_X1 U7781 ( .A1(n6510), .A2(n6611), .ZN(n6610) );
  INV_X1 U7782 ( .A(n6904), .ZN(n6903) );
  OAI21_X1 U7783 ( .B1(n6906), .B2(n6905), .A(n12067), .ZN(n6904) );
  NAND2_X1 U7784 ( .A1(n6908), .A2(n6906), .ZN(n11997) );
  NAND2_X1 U7785 ( .A1(n6473), .A2(n12029), .ZN(n6908) );
  AND4_X1 U7786 ( .A1(n9166), .A2(n9165), .A3(n9164), .A4(n9163), .ZN(n11918)
         );
  AND4_X1 U7787 ( .A1(n9149), .A2(n9148), .A3(n9147), .A4(n9146), .ZN(n11955)
         );
  AND3_X1 U7788 ( .A1(n8781), .A2(n8780), .A3(n8779), .ZN(n12047) );
  AND4_X1 U7789 ( .A1(n8940), .A2(n8939), .A3(n8938), .A4(n8937), .ZN(n11385)
         );
  OAI21_X1 U7790 ( .B1(n10143), .B2(n7291), .A(n10124), .ZN(n10125) );
  AND2_X1 U7791 ( .A1(n10204), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7291) );
  OR2_X1 U7792 ( .A1(n10432), .A2(n6480), .ZN(n6808) );
  NAND2_X1 U7793 ( .A1(n10432), .A2(n6810), .ZN(n6807) );
  NAND2_X1 U7794 ( .A1(n6468), .A2(n6810), .ZN(n6809) );
  NAND2_X1 U7795 ( .A1(n7284), .A2(n7283), .ZN(n10432) );
  NAND2_X1 U7796 ( .A1(n10293), .A2(n7288), .ZN(n7283) );
  OR2_X1 U7797 ( .A1(n10276), .A2(n7285), .ZN(n7284) );
  NAND2_X1 U7798 ( .A1(n7288), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7285) );
  OR2_X1 U7799 ( .A1(n10300), .A2(n10299), .ZN(n10511) );
  OR2_X1 U7800 ( .A1(n10516), .A2(n7106), .ZN(n7103) );
  INV_X1 U7801 ( .A(n10649), .ZN(n7105) );
  OR2_X1 U7802 ( .A1(n10516), .A2(n15035), .ZN(n7108) );
  NOR2_X1 U7803 ( .A1(n10759), .A2(n7290), .ZN(n10950) );
  AND2_X1 U7804 ( .A1(n10762), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7290) );
  OR2_X1 U7805 ( .A1(n14899), .A2(n12349), .ZN(n7111) );
  XNOR2_X1 U7806 ( .A(n12386), .B(n12387), .ZN(n14919) );
  NOR2_X1 U7807 ( .A1(n12387), .A2(n12386), .ZN(n12388) );
  OAI21_X1 U7808 ( .B1(n14919), .B2(n7114), .A(n7113), .ZN(n12394) );
  NAND2_X1 U7809 ( .A1(n12374), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7114) );
  NAND2_X1 U7810 ( .A1(n12388), .A2(n12374), .ZN(n7113) );
  OR2_X1 U7811 ( .A1(n14919), .A2(n14920), .ZN(n7116) );
  OAI21_X1 U7812 ( .B1(n14268), .B2(n7118), .A(n7117), .ZN(n14289) );
  NAND2_X1 U7813 ( .A1(n7121), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7118) );
  INV_X1 U7814 ( .A(n14290), .ZN(n7121) );
  OR2_X1 U7815 ( .A1(n14268), .A2(n14269), .ZN(n7120) );
  NOR2_X1 U7816 ( .A1(n12467), .A2(n7128), .ZN(n7127) );
  INV_X1 U7817 ( .A(n12466), .ZN(n7128) );
  AOI21_X1 U7818 ( .B1(n6866), .B2(n12186), .A(n6865), .ZN(n6864) );
  INV_X1 U7819 ( .A(n12199), .ZN(n6865) );
  INV_X1 U7820 ( .A(n6867), .ZN(n6866) );
  OAI21_X1 U7821 ( .B1(n6869), .B2(n12186), .A(n6868), .ZN(n6867) );
  NOR2_X1 U7822 ( .A1(n6871), .A2(n6870), .ZN(n6869) );
  INV_X1 U7823 ( .A(n12189), .ZN(n6871) );
  INV_X1 U7824 ( .A(n9247), .ZN(n6870) );
  NAND2_X1 U7825 ( .A1(n6832), .A2(n12174), .ZN(n11063) );
  INV_X1 U7826 ( .A(n12274), .ZN(n6850) );
  INV_X1 U7827 ( .A(n6848), .ZN(n6847) );
  OAI21_X1 U7828 ( .B1(n12274), .B2(n6849), .A(n12272), .ZN(n6848) );
  NAND2_X1 U7829 ( .A1(n12275), .A2(n12099), .ZN(n12130) );
  AOI21_X1 U7830 ( .B1(n12495), .B2(n12269), .A(n12267), .ZN(n12486) );
  NAND2_X1 U7831 ( .A1(n9273), .A2(n9272), .ZN(n9293) );
  INV_X1 U7832 ( .A(n12276), .ZN(n12108) );
  OR2_X1 U7833 ( .A1(n12032), .A2(n12685), .ZN(n7388) );
  NOR2_X1 U7834 ( .A1(n12267), .A2(n12109), .ZN(n12497) );
  OAI21_X1 U7835 ( .B1(n12506), .B2(n12256), .A(n12263), .ZN(n12495) );
  NOR2_X1 U7836 ( .A1(n12532), .A2(n7264), .ZN(n7262) );
  INV_X1 U7837 ( .A(n12520), .ZN(n7265) );
  OAI21_X1 U7838 ( .B1(n12528), .B2(n6841), .A(n12258), .ZN(n6840) );
  INV_X1 U7839 ( .A(n12134), .ZN(n6841) );
  NOR2_X1 U7840 ( .A1(n7265), .A2(n6840), .ZN(n6838) );
  NAND2_X1 U7841 ( .A1(n12539), .A2(n6842), .ZN(n6839) );
  NOR2_X1 U7842 ( .A1(n12532), .A2(n12531), .ZN(n12530) );
  AND2_X1 U7843 ( .A1(n9090), .A2(n9089), .ZN(n9096) );
  NOR2_X1 U7844 ( .A1(n7249), .A2(n7248), .ZN(n7246) );
  NOR2_X1 U7845 ( .A1(n7252), .A2(n6526), .ZN(n7249) );
  INV_X1 U7846 ( .A(n7251), .ZN(n7248) );
  NAND2_X1 U7847 ( .A1(n7255), .A2(n6491), .ZN(n7247) );
  AND2_X1 U7848 ( .A1(n12243), .A2(n12244), .ZN(n12560) );
  NAND2_X1 U7849 ( .A1(n9064), .A2(n9063), .ZN(n12111) );
  NAND2_X1 U7850 ( .A1(n9253), .A2(n12233), .ZN(n6856) );
  AND2_X1 U7851 ( .A1(n12228), .A2(n12231), .ZN(n12581) );
  NAND2_X1 U7852 ( .A1(n6860), .A2(n12591), .ZN(n6859) );
  INV_X1 U7853 ( .A(n12590), .ZN(n6860) );
  NOR2_X1 U7854 ( .A1(n12579), .A2(n6858), .ZN(n6857) );
  INV_X1 U7855 ( .A(n12233), .ZN(n6858) );
  INV_X1 U7856 ( .A(n12581), .ZN(n12579) );
  OAI21_X1 U7857 ( .B1(n12612), .B2(n12614), .A(n12217), .ZN(n12603) );
  NAND2_X1 U7858 ( .A1(n12216), .A2(n12217), .ZN(n12614) );
  AND2_X1 U7859 ( .A1(n8933), .A2(n8917), .ZN(n7279) );
  AND3_X1 U7860 ( .A1(n8932), .A2(n8931), .A3(n8930), .ZN(n15015) );
  INV_X1 U7861 ( .A(n7035), .ZN(n7034) );
  OAI21_X1 U7862 ( .B1(n7036), .B2(n11910), .A(n11909), .ZN(n7035) );
  AND2_X1 U7863 ( .A1(n6515), .A2(n7276), .ZN(n7275) );
  NOR2_X1 U7864 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), .ZN(
        n7276) );
  XNOR2_X1 U7865 ( .A(n9202), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9217) );
  NAND2_X1 U7866 ( .A1(n9203), .A2(n8762), .ZN(n9201) );
  AOI21_X1 U7867 ( .B1(n7045), .B2(n9083), .A(n6597), .ZN(n7043) );
  INV_X1 U7868 ( .A(n7045), .ZN(n7044) );
  OR2_X1 U7869 ( .A1(n8701), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n9198) );
  XNOR2_X1 U7870 ( .A(n8702), .B(P3_IR_REG_21__SCAN_IN), .ZN(n10145) );
  INV_X1 U7871 ( .A(n8964), .ZN(n7059) );
  OR2_X1 U7872 ( .A1(n8958), .A2(n8730), .ZN(n7060) );
  NAND2_X1 U7873 ( .A1(n9767), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8715) );
  XNOR2_X1 U7874 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8868) );
  INV_X1 U7875 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n8709) );
  AOI21_X1 U7876 ( .B1(n6469), .B2(n6465), .A(n6564), .ZN(n6691) );
  AND2_X1 U7877 ( .A1(n11141), .A2(n9624), .ZN(n7177) );
  AND2_X1 U7878 ( .A1(n7938), .A2(n7937), .ZN(n9697) );
  OR2_X1 U7879 ( .A1(n6439), .A2(n9882), .ZN(n7062) );
  INV_X1 U7880 ( .A(n9543), .ZN(n12959) );
  OR2_X1 U7881 ( .A1(n7940), .A2(n7939), .ZN(n7951) );
  AND2_X1 U7882 ( .A1(n7950), .A2(n7948), .ZN(n13015) );
  NOR2_X1 U7883 ( .A1(n6728), .A2(n7929), .ZN(n6725) );
  INV_X1 U7884 ( .A(n6729), .ZN(n6724) );
  INV_X1 U7885 ( .A(n6725), .ZN(n6723) );
  NAND2_X1 U7886 ( .A1(n6720), .A2(n6717), .ZN(n13032) );
  INV_X1 U7887 ( .A(n6718), .ZN(n6717) );
  OAI21_X1 U7888 ( .B1(n6727), .B2(n6732), .A(n6555), .ZN(n6718) );
  NAND2_X1 U7889 ( .A1(n7093), .A2(n6495), .ZN(n7092) );
  INV_X1 U7890 ( .A(n7095), .ZN(n7093) );
  INV_X1 U7891 ( .A(n9542), .ZN(n13033) );
  NOR2_X1 U7892 ( .A1(n13062), .A2(n13083), .ZN(n6729) );
  XNOR2_X1 U7893 ( .A(n9433), .B(n13036), .ZN(n13052) );
  NOR2_X1 U7894 ( .A1(n13226), .A2(n13080), .ZN(n7096) );
  NOR2_X1 U7895 ( .A1(n13052), .A2(n7096), .ZN(n7095) );
  NAND2_X1 U7896 ( .A1(n7098), .A2(n6470), .ZN(n7097) );
  AND2_X1 U7897 ( .A1(n7928), .A2(n7927), .ZN(n13068) );
  AND2_X1 U7898 ( .A1(n7911), .A2(n7910), .ZN(n13066) );
  INV_X1 U7899 ( .A(n9539), .ZN(n13062) );
  OR2_X1 U7900 ( .A1(n7005), .A2(n7004), .ZN(n7003) );
  INV_X1 U7901 ( .A(n7007), .ZN(n7004) );
  NOR2_X1 U7902 ( .A1(n7888), .A2(n6519), .ZN(n7005) );
  NOR2_X1 U7903 ( .A1(n13172), .A2(n6828), .ZN(n13139) );
  NOR2_X1 U7904 ( .A1(n13172), .A2(n6827), .ZN(n13115) );
  NAND2_X1 U7905 ( .A1(n7083), .A2(n6497), .ZN(n7082) );
  NAND2_X1 U7906 ( .A1(n11745), .A2(n7861), .ZN(n13167) );
  AND2_X1 U7907 ( .A1(n11467), .A2(n7835), .ZN(n7383) );
  NAND2_X1 U7908 ( .A1(n7383), .A2(n7843), .ZN(n11709) );
  OR2_X1 U7909 ( .A1(n11551), .A2(n9534), .ZN(n11552) );
  AND2_X1 U7910 ( .A1(n9534), .A2(n7816), .ZN(n7021) );
  NAND2_X1 U7911 ( .A1(n11152), .A2(n7816), .ZN(n11558) );
  NAND2_X1 U7912 ( .A1(n11220), .A2(n7790), .ZN(n11203) );
  INV_X1 U7913 ( .A(n7075), .ZN(n7074) );
  NAND2_X1 U7914 ( .A1(n11243), .A2(n11242), .ZN(n7077) );
  INV_X1 U7915 ( .A(n7979), .ZN(n7066) );
  INV_X1 U7916 ( .A(n11025), .ZN(n7067) );
  AND2_X1 U7917 ( .A1(n9719), .A2(n9873), .ZN(n13152) );
  AND2_X1 U7918 ( .A1(n11268), .A2(n7747), .ZN(n10814) );
  AND2_X1 U7919 ( .A1(n10820), .A2(n7743), .ZN(n10876) );
  INV_X1 U7920 ( .A(n13069), .ZN(n13153) );
  INV_X1 U7921 ( .A(n6953), .ZN(n9302) );
  NOR2_X1 U7922 ( .A1(n12984), .A2(n12985), .ZN(n7019) );
  NAND2_X1 U7923 ( .A1(n6743), .A2(n6742), .ZN(n6741) );
  NAND2_X1 U7924 ( .A1(n12772), .A2(n14841), .ZN(n6742) );
  INV_X1 U7925 ( .A(n13002), .ZN(n6743) );
  NOR2_X1 U7926 ( .A1(n8033), .A2(n10809), .ZN(n10552) );
  NAND2_X1 U7927 ( .A1(n13297), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6734) );
  OR2_X1 U7928 ( .A1(n7721), .A2(n7718), .ZN(n6738) );
  NOR2_X1 U7929 ( .A1(n6737), .A2(n6736), .ZN(n6735) );
  INV_X1 U7930 ( .A(n7696), .ZN(n7523) );
  AOI21_X1 U7931 ( .B1(n7141), .B2(n7144), .A(n7139), .ZN(n7138) );
  INV_X1 U7932 ( .A(n13496), .ZN(n7139) );
  INV_X1 U7933 ( .A(n13506), .ZN(n7160) );
  NAND2_X1 U7934 ( .A1(n10043), .A2(n7172), .ZN(n10047) );
  NAND2_X1 U7935 ( .A1(n10598), .A2(n14518), .ZN(n7172) );
  NAND2_X1 U7936 ( .A1(n7155), .A2(n7156), .ZN(n7154) );
  AND2_X1 U7937 ( .A1(n8531), .A2(n8530), .ZN(n13755) );
  INV_X1 U7938 ( .A(n8589), .ZN(n8525) );
  OR2_X1 U7939 ( .A1(n6464), .A2(n8121), .ZN(n8122) );
  INV_X1 U7940 ( .A(n8056), .ZN(n7359) );
  INV_X1 U7941 ( .A(n13770), .ZN(n13781) );
  NAND2_X1 U7942 ( .A1(n13756), .A2(n8630), .ZN(n13770) );
  OR2_X1 U7943 ( .A1(n13980), .A2(n13759), .ZN(n8630) );
  NOR2_X1 U7944 ( .A1(n11865), .A2(n7355), .ZN(n7354) );
  INV_X1 U7945 ( .A(n11864), .ZN(n7355) );
  NOR2_X1 U7946 ( .A1(n13821), .A2(n6897), .ZN(n6896) );
  INV_X1 U7947 ( .A(n11877), .ZN(n6897) );
  NAND2_X1 U7948 ( .A1(n13873), .A2(n7357), .ZN(n13852) );
  AND2_X1 U7949 ( .A1(n11858), .A2(n11857), .ZN(n7357) );
  NOR2_X1 U7950 ( .A1(n13870), .A2(n6472), .ZN(n6894) );
  NAND2_X1 U7951 ( .A1(n6639), .A2(n6647), .ZN(n11875) );
  OR2_X1 U7952 ( .A1(n13944), .A2(n6650), .ZN(n6639) );
  NAND2_X1 U7953 ( .A1(n13905), .A2(n11855), .ZN(n13891) );
  NOR2_X1 U7954 ( .A1(n13890), .A2(n7361), .ZN(n7360) );
  INV_X1 U7955 ( .A(n11855), .ZN(n7361) );
  NAND2_X1 U7956 ( .A1(n6944), .A2(n6943), .ZN(n13934) );
  OR2_X1 U7957 ( .A1(n14362), .A2(n14324), .ZN(n11785) );
  INV_X1 U7958 ( .A(n11850), .ZN(n11868) );
  NOR2_X1 U7959 ( .A1(n6633), .A2(n11764), .ZN(n6632) );
  INV_X1 U7960 ( .A(n6636), .ZN(n6633) );
  INV_X1 U7961 ( .A(n6948), .ZN(n6628) );
  NOR2_X1 U7962 ( .A1(n8215), .A2(n8214), .ZN(n8226) );
  AND2_X1 U7963 ( .A1(n11180), .A2(n11190), .ZN(n7356) );
  AND3_X1 U7964 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n8173) );
  AND2_X1 U7965 ( .A1(n8600), .A2(n8599), .ZN(n13970) );
  NAND2_X1 U7966 ( .A1(n11626), .A2(n8381), .ZN(n8519) );
  NAND2_X1 U7967 ( .A1(n8486), .A2(n8485), .ZN(n13827) );
  AND2_X1 U7968 ( .A1(n8423), .A2(n8422), .ZN(n14019) );
  AND2_X1 U7969 ( .A1(n14528), .A2(n10065), .ZN(n14584) );
  XNOR2_X1 U7970 ( .A(n8620), .B(n8619), .ZN(n13295) );
  NAND2_X1 U7971 ( .A1(n8554), .A2(n8553), .ZN(n8557) );
  INV_X1 U7972 ( .A(n6795), .ZN(n8554) );
  OAI21_X1 U7973 ( .B1(n7710), .B2(n6598), .A(n6485), .ZN(n6795) );
  INV_X1 U7974 ( .A(n7366), .ZN(n7364) );
  XNOR2_X1 U7975 ( .A(n7697), .B(n9088), .ZN(n8455) );
  AND2_X1 U7976 ( .A1(n7347), .A2(n7346), .ZN(n7345) );
  INV_X1 U7977 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7346) );
  INV_X1 U7978 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7162) );
  AND2_X1 U7979 ( .A1(n8064), .A2(n8326), .ZN(n8357) );
  XNOR2_X1 U7980 ( .A(n7605), .B(n7606), .ZN(n9851) );
  NAND2_X1 U7981 ( .A1(n7218), .A2(n7442), .ZN(n7605) );
  NAND2_X1 U7982 ( .A1(n6748), .A2(n7370), .ZN(n7544) );
  XNOR2_X1 U7983 ( .A(n14133), .B(n14134), .ZN(n14136) );
  XNOR2_X1 U7984 ( .A(n14093), .B(P3_ADDR_REG_3__SCAN_IN), .ZN(n14139) );
  INV_X1 U7985 ( .A(n6679), .ZN(n14149) );
  OAI21_X1 U7986 ( .B1(n15196), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6538), .ZN(
        n6679) );
  NAND2_X1 U7987 ( .A1(n14100), .A2(n14099), .ZN(n14151) );
  OR2_X1 U7988 ( .A1(n14145), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n14099) );
  NOR2_X1 U7989 ( .A1(n14160), .A2(n14161), .ZN(n14164) );
  INV_X1 U7990 ( .A(n14166), .ZN(n6682) );
  NOR2_X1 U7991 ( .A1(n14401), .A2(n6664), .ZN(n6663) );
  INV_X1 U7992 ( .A(n6667), .ZN(n6664) );
  AND2_X1 U7993 ( .A1(n6672), .A2(n6669), .ZN(n14187) );
  AOI21_X1 U7994 ( .B1(n14177), .B2(n6671), .A(n6670), .ZN(n6669) );
  INV_X1 U7995 ( .A(n6674), .ZN(n6673) );
  NAND2_X1 U7996 ( .A1(n9157), .A2(n9156), .ZN(n12627) );
  INV_X1 U7997 ( .A(n12697), .ZN(n12255) );
  INV_X1 U7998 ( .A(n11955), .ZN(n12309) );
  INV_X1 U7999 ( .A(n12058), .ZN(n12316) );
  AND4_X1 U8000 ( .A1(n9057), .A2(n9056), .A3(n9055), .A4(n9054), .ZN(n12056)
         );
  INV_X1 U8001 ( .A(n11459), .ZN(n12323) );
  NOR2_X1 U8002 ( .A1(n7109), .A2(n10204), .ZN(n10202) );
  INV_X1 U8003 ( .A(n10121), .ZN(n7109) );
  OR2_X1 U8004 ( .A1(n10760), .A2(n10761), .ZN(n7289) );
  XNOR2_X1 U8005 ( .A(n10950), .B(n10957), .ZN(n10760) );
  NAND2_X1 U8006 ( .A1(n7281), .A2(n6514), .ZN(n7280) );
  AND2_X1 U8007 ( .A1(n7280), .A2(n6818), .ZN(n12363) );
  INV_X1 U8008 ( .A(n12338), .ZN(n6818) );
  INV_X1 U8009 ( .A(n7303), .ZN(n7302) );
  AOI211_X1 U8010 ( .C1(n12425), .C2(n12419), .A(n6593), .B(n7304), .ZN(n7303)
         );
  INV_X1 U8011 ( .A(n12406), .ZN(n7304) );
  OAI21_X1 U8012 ( .B1(n12405), .B2(n12429), .A(n12434), .ZN(n7305) );
  AOI21_X1 U8013 ( .B1(n12433), .B2(n12432), .A(n12431), .ZN(n12449) );
  NAND2_X1 U8014 ( .A1(n12763), .A2(n12083), .ZN(n9174) );
  NAND2_X1 U8015 ( .A1(n9050), .A2(n9049), .ZN(n12600) );
  NAND2_X1 U8016 ( .A1(n9009), .A2(n9008), .ZN(n14298) );
  AND2_X1 U8017 ( .A1(n8976), .A2(n8975), .ZN(n11462) );
  AND2_X1 U8018 ( .A1(n14944), .A2(n9292), .ZN(n12621) );
  INV_X1 U8019 ( .A(n12489), .ZN(n12618) );
  INV_X1 U8020 ( .A(n13007), .ZN(n12772) );
  NOR2_X1 U8021 ( .A1(n7186), .A2(n7182), .ZN(n7181) );
  INV_X1 U8022 ( .A(n7187), .ZN(n7186) );
  OAI21_X1 U8023 ( .B1(n9717), .B2(n9721), .A(n7188), .ZN(n7187) );
  NAND2_X1 U8024 ( .A1(n9717), .A2(n7189), .ZN(n7188) );
  OAI21_X1 U8025 ( .B1(n9717), .B2(n9739), .A(n7185), .ZN(n7184) );
  NAND2_X1 U8026 ( .A1(n9717), .A2(n9722), .ZN(n7185) );
  INV_X1 U8027 ( .A(n9715), .ZN(n7182) );
  NOR2_X1 U8028 ( .A1(n12766), .A2(n6694), .ZN(n6693) );
  INV_X1 U8029 ( .A(n9708), .ZN(n6694) );
  NAND2_X1 U8030 ( .A1(n10686), .A2(n10687), .ZN(n10685) );
  NAND2_X1 U8031 ( .A1(n7668), .A2(n7667), .ZN(n13258) );
  NAND2_X1 U8032 ( .A1(n7604), .A2(n7603), .ZN(n14829) );
  NAND2_X1 U8033 ( .A1(n9620), .A2(n9621), .ZN(n11098) );
  AND2_X1 U8034 ( .A1(n9645), .A2(n9639), .ZN(n7199) );
  INV_X1 U8035 ( .A(n12865), .ZN(n12858) );
  NAND2_X1 U8036 ( .A1(n9725), .A2(n13133), .ZN(n12871) );
  NOR2_X1 U8037 ( .A1(n9517), .A2(n9516), .ZN(n9525) );
  INV_X1 U8038 ( .A(n13068), .ZN(n13036) );
  INV_X1 U8039 ( .A(n12846), .ZN(n13080) );
  XNOR2_X1 U8040 ( .A(n7409), .B(P2_IR_REG_19__SCAN_IN), .ZN(n12997) );
  NAND2_X1 U8041 ( .A1(n7198), .A2(n7197), .ZN(n7408) );
  NAND2_X1 U8042 ( .A1(n6744), .A2(n7973), .ZN(n13009) );
  INV_X1 U8043 ( .A(n6745), .ZN(n6744) );
  AND2_X1 U8044 ( .A1(n7006), .A2(n7008), .ZN(n13109) );
  NAND2_X1 U8045 ( .A1(n13147), .A2(n7995), .ZN(n13125) );
  INV_X1 U8046 ( .A(n7684), .ZN(n7537) );
  NOR2_X1 U8047 ( .A1(n13196), .A2(n14852), .ZN(n13197) );
  NAND2_X1 U8048 ( .A1(n8036), .A2(n8035), .ZN(n14763) );
  OAI211_X1 U8049 ( .C1(n8574), .C2(n9754), .A(n8133), .B(n8132), .ZN(n13446)
         );
  INV_X1 U8050 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7410) );
  XNOR2_X1 U8051 ( .A(n7220), .B(n13757), .ZN(n7219) );
  NAND2_X1 U8052 ( .A1(n13780), .A2(n13756), .ZN(n7220) );
  INV_X1 U8053 ( .A(n13970), .ZN(n13764) );
  OAI21_X1 U8054 ( .B1(n6900), .B2(n14549), .A(n11887), .ZN(n11888) );
  NAND2_X1 U8055 ( .A1(n7225), .A2(n11876), .ZN(n13833) );
  AND2_X1 U8056 ( .A1(n14543), .A2(n14536), .ZN(n14511) );
  AND2_X1 U8057 ( .A1(n14543), .A2(n11077), .ZN(n14501) );
  AND2_X1 U8058 ( .A1(n8533), .A2(n8532), .ZN(n14052) );
  INV_X1 U8059 ( .A(n13747), .ZN(n14536) );
  INV_X1 U8060 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14135) );
  XNOR2_X1 U8061 ( .A(n14136), .B(n6685), .ZN(n15207) );
  NOR2_X1 U8062 ( .A1(n14203), .A2(n14202), .ZN(n14201) );
  NOR2_X1 U8063 ( .A1(n14201), .A2(n6658), .ZN(n15203) );
  AOI21_X1 U8064 ( .B1(n14203), .B2(n14202), .A(P2_ADDR_REG_2__SCAN_IN), .ZN(
        n6658) );
  XNOR2_X1 U8065 ( .A(n14164), .B(n6874), .ZN(n14227) );
  INV_X1 U8066 ( .A(n14165), .ZN(n6874) );
  INV_X1 U8067 ( .A(n6656), .ZN(n14388) );
  OAI21_X1 U8068 ( .B1(n14384), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6657), .ZN(
        n6656) );
  AND2_X1 U8069 ( .A1(n6659), .A2(n6665), .ZN(n14400) );
  NAND2_X1 U8070 ( .A1(n6678), .A2(n6677), .ZN(n6676) );
  XNOR2_X1 U8071 ( .A(n14187), .B(n14186), .ZN(n14198) );
  NOR2_X1 U8072 ( .A1(n14198), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n14189) );
  NAND2_X1 U8073 ( .A1(n9329), .A2(n6978), .ZN(n6977) );
  AOI21_X1 U8074 ( .B1(n7312), .B2(n7314), .A(n7311), .ZN(n8166) );
  NOR2_X1 U8075 ( .A1(n8151), .A2(n8150), .ZN(n7311) );
  AOI21_X1 U8076 ( .B1(n8150), .B2(n8151), .A(n7313), .ZN(n7312) );
  OR2_X1 U8077 ( .A1(n8189), .A2(n7344), .ZN(n7343) );
  INV_X1 U8078 ( .A(n8188), .ZN(n7344) );
  NAND2_X1 U8079 ( .A1(n6975), .A2(n9347), .ZN(n6974) );
  NOR2_X1 U8080 ( .A1(n8237), .A2(n8238), .ZN(n7324) );
  NAND2_X1 U8081 ( .A1(n8225), .A2(n7325), .ZN(n7323) );
  AOI21_X1 U8082 ( .B1(n8237), .B2(n8238), .A(n6559), .ZN(n7325) );
  INV_X1 U8083 ( .A(n8274), .ZN(n7332) );
  NAND2_X1 U8084 ( .A1(n6984), .A2(n9366), .ZN(n6983) );
  NAND2_X1 U8085 ( .A1(n6504), .A2(n6475), .ZN(n7306) );
  INV_X1 U8086 ( .A(n9376), .ZN(n6966) );
  NOR2_X1 U8087 ( .A1(n9379), .A2(n9376), .ZN(n6967) );
  OAI21_X1 U8088 ( .B1(n8412), .B2(n8411), .A(n8410), .ZN(n8426) );
  NAND2_X1 U8089 ( .A1(n9394), .A2(n9395), .ZN(n9393) );
  NAND2_X1 U8090 ( .A1(n7335), .A2(n8457), .ZN(n7334) );
  NAND2_X1 U8091 ( .A1(n7338), .A2(n8487), .ZN(n7337) );
  NAND2_X1 U8092 ( .A1(n6963), .A2(n9418), .ZN(n6962) );
  NAND2_X1 U8093 ( .A1(n9417), .A2(n6959), .ZN(n6958) );
  INV_X1 U8094 ( .A(n7210), .ZN(n7209) );
  OAI21_X1 U8095 ( .B1(n7376), .B2(n7211), .A(n7631), .ZN(n7210) );
  INV_X1 U8096 ( .A(n7452), .ZN(n7211) );
  INV_X1 U8097 ( .A(n7456), .ZN(n7207) );
  NAND2_X1 U8098 ( .A1(n7341), .A2(n8520), .ZN(n7340) );
  INV_X1 U8099 ( .A(n12402), .ZN(n7300) );
  NAND2_X1 U8100 ( .A1(n6970), .A2(n9427), .ZN(n6969) );
  INV_X1 U8101 ( .A(n9425), .ZN(n6970) );
  AND2_X1 U8102 ( .A1(n10209), .A2(n10038), .ZN(n10578) );
  INV_X1 U8103 ( .A(n8563), .ZN(n7330) );
  NOR2_X1 U8104 ( .A1(n6548), .A2(n6653), .ZN(n6652) );
  INV_X1 U8105 ( .A(n11873), .ZN(n6653) );
  AOI21_X1 U8106 ( .B1(n6804), .B2(n7713), .A(n6802), .ZN(n6801) );
  NOR2_X1 U8107 ( .A1(n7502), .A2(SI_26_), .ZN(n6802) );
  INV_X1 U8108 ( .A(n7705), .ZN(n6783) );
  NAND2_X1 U8109 ( .A1(n6764), .A2(n7482), .ZN(n7484) );
  NAND2_X1 U8110 ( .A1(n7676), .A2(n7477), .ZN(n6764) );
  NAND2_X1 U8111 ( .A1(n7676), .A2(n6755), .ZN(n6754) );
  NOR2_X1 U8112 ( .A1(n6756), .A2(n6483), .ZN(n6755) );
  INV_X1 U8113 ( .A(n6758), .ZN(n6756) );
  NAND2_X1 U8114 ( .A1(n6758), .A2(n6762), .ZN(n6757) );
  AOI21_X1 U8115 ( .B1(n6774), .B2(n6777), .A(n6560), .ZN(n6772) );
  NOR2_X1 U8116 ( .A1(n7606), .A2(n7599), .ZN(n7215) );
  INV_X1 U8117 ( .A(n7442), .ZN(n7217) );
  AND2_X1 U8118 ( .A1(n6910), .A2(n11936), .ZN(n11938) );
  NOR2_X1 U8119 ( .A1(n11938), .A2(n11937), .ZN(n11940) );
  NAND2_X1 U8120 ( .A1(n11513), .A2(n12323), .ZN(n6611) );
  NAND2_X1 U8121 ( .A1(n11507), .A2(n11516), .ZN(n6935) );
  NOR2_X1 U8122 ( .A1(n12485), .A2(n6616), .ZN(n6615) );
  INV_X1 U8123 ( .A(n12270), .ZN(n6616) );
  CLKBUF_X1 U8124 ( .A(n10274), .Z(n6625) );
  NOR2_X1 U8125 ( .A1(n10344), .A2(n10281), .ZN(n10316) );
  INV_X1 U8126 ( .A(n10433), .ZN(n7288) );
  OR2_X1 U8127 ( .A1(n10649), .A2(n15035), .ZN(n7106) );
  NAND2_X1 U8128 ( .A1(n10515), .A2(n10514), .ZN(n6624) );
  OR2_X1 U8129 ( .A1(n10764), .A2(n10763), .ZN(n10955) );
  INV_X1 U8130 ( .A(n12408), .ZN(n7297) );
  NOR2_X1 U8131 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(n9091), .ZN(n9103) );
  NOR2_X1 U8132 ( .A1(n8996), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9011) );
  OR2_X1 U8133 ( .A1(n12273), .A2(n12297), .ZN(n10171) );
  OR2_X1 U8134 ( .A1(n12477), .A2(n11956), .ZN(n12272) );
  AND2_X1 U8135 ( .A1(n12272), .A2(n9290), .ZN(n12276) );
  INV_X1 U8136 ( .A(n6491), .ZN(n7243) );
  NAND2_X1 U8137 ( .A1(n12720), .A2(n12316), .ZN(n7251) );
  NOR2_X1 U8138 ( .A1(n12581), .A2(n12582), .ZN(n7254) );
  AND2_X1 U8139 ( .A1(n12614), .A2(n7230), .ZN(n7229) );
  NAND2_X1 U8140 ( .A1(n7231), .A2(n9017), .ZN(n7230) );
  NAND2_X1 U8141 ( .A1(n6603), .A2(n9271), .ZN(n7036) );
  NOR2_X1 U8142 ( .A1(n11910), .A2(n7038), .ZN(n7037) );
  INV_X1 U8143 ( .A(n9271), .ZN(n7038) );
  INV_X1 U8144 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7277) );
  INV_X1 U8145 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8762) );
  AND2_X1 U8146 ( .A1(n9206), .A2(n8761), .ZN(n9203) );
  INV_X1 U8147 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8756) );
  INV_X1 U8148 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8755) );
  NOR2_X1 U8149 ( .A1(n9098), .A2(n7046), .ZN(n7045) );
  INV_X1 U8150 ( .A(n9086), .ZN(n7046) );
  AND2_X1 U8151 ( .A1(n8699), .A2(n8756), .ZN(n8703) );
  OR2_X1 U8152 ( .A1(n8928), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n8972) );
  OR2_X1 U8153 ( .A1(n8882), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8896) );
  OR3_X1 U8154 ( .A1(n9718), .A2(n14763), .A3(n14766), .ZN(n9727) );
  INV_X1 U8155 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7395) );
  NOR2_X1 U8156 ( .A1(n12772), .A2(n13209), .ZN(n6825) );
  NOR2_X1 U8157 ( .A1(n7951), .A2(n15074), .ZN(n7961) );
  NAND2_X1 U8158 ( .A1(n7929), .A2(n6731), .ZN(n6719) );
  AND2_X1 U8159 ( .A1(n6729), .A2(n6731), .ZN(n6721) );
  AOI21_X1 U8160 ( .B1(n7003), .B2(n7001), .A(n6546), .ZN(n7000) );
  INV_X1 U8161 ( .A(n6492), .ZN(n7001) );
  INV_X1 U8162 ( .A(n7003), .ZN(n7002) );
  OR2_X1 U8163 ( .A1(n13246), .A2(n13253), .ZN(n6828) );
  NAND2_X1 U8164 ( .A1(n7084), .A2(n7996), .ZN(n7083) );
  INV_X1 U8165 ( .A(n7995), .ZN(n7084) );
  OR2_X1 U8166 ( .A1(n7837), .A2(n7836), .ZN(n7846) );
  NOR2_X1 U8167 ( .A1(n11209), .A2(n14842), .ZN(n6822) );
  AND2_X1 U8168 ( .A1(n9524), .A2(n9548), .ZN(n9719) );
  NAND2_X1 U8169 ( .A1(n13040), .A2(n13028), .ZN(n13022) );
  OR2_X1 U8170 ( .A1(n11723), .A2(n13269), .ZN(n11751) );
  NOR2_X1 U8171 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n6736) );
  INV_X1 U8172 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7514) );
  INV_X1 U8173 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n7102) );
  INV_X1 U8174 ( .A(n7157), .ZN(n7155) );
  AND2_X1 U8175 ( .A1(n8601), .A2(n7328), .ZN(n7327) );
  NAND2_X1 U8176 ( .A1(n7329), .A2(n8563), .ZN(n7328) );
  INV_X1 U8177 ( .A(n8602), .ZN(n7329) );
  NAND2_X1 U8178 ( .A1(n14242), .A2(n14243), .ZN(n6638) );
  NAND2_X1 U8179 ( .A1(n6949), .A2(n14369), .ZN(n6948) );
  XNOR2_X1 U8180 ( .A(n13597), .B(n11318), .ZN(n10708) );
  INV_X1 U8181 ( .A(n6709), .ZN(n6708) );
  OAI21_X1 U8182 ( .B1(n7353), .B2(n11862), .A(n7352), .ZN(n6709) );
  AOI21_X1 U8183 ( .B1(n7354), .B2(n11878), .A(n6550), .ZN(n7352) );
  INV_X1 U8184 ( .A(n7354), .ZN(n7353) );
  INV_X1 U8185 ( .A(n6641), .ZN(n6640) );
  NAND2_X1 U8186 ( .A1(n13944), .A2(n6644), .ZN(n6643) );
  OAI21_X1 U8187 ( .B1(n6892), .B2(n6642), .A(n6890), .ZN(n6641) );
  NAND2_X1 U8188 ( .A1(n6456), .A2(n11851), .ZN(n13946) );
  INV_X1 U8189 ( .A(n11351), .ZN(n11188) );
  NOR2_X1 U8190 ( .A1(n6803), .A2(SI_27_), .ZN(n6799) );
  NAND2_X1 U8191 ( .A1(n7367), .A2(n8048), .ZN(n7366) );
  INV_X1 U8192 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n7367) );
  OR2_X1 U8193 ( .A1(n7495), .A2(n6793), .ZN(n6791) );
  NAND2_X1 U8194 ( .A1(n6792), .A2(n6789), .ZN(n6788) );
  INV_X1 U8195 ( .A(n7492), .ZN(n6789) );
  INV_X1 U8196 ( .A(n7692), .ZN(n7487) );
  NAND2_X1 U8197 ( .A1(n7448), .A2(n7447), .ZN(n7614) );
  INV_X1 U8198 ( .A(n7591), .ZN(n7437) );
  XNOR2_X1 U8199 ( .A(n7438), .B(SI_8_), .ZN(n7591) );
  XNOR2_X1 U8200 ( .A(n7435), .B(SI_7_), .ZN(n7581) );
  NOR2_X1 U8201 ( .A1(n6750), .A2(n7213), .ZN(n6749) );
  OAI21_X1 U8202 ( .B1(n7428), .B2(n7213), .A(n7431), .ZN(n6751) );
  NAND2_X1 U8203 ( .A1(n6496), .A2(n7427), .ZN(n6750) );
  XNOR2_X1 U8204 ( .A(n7426), .B(SI_4_), .ZN(n7557) );
  NAND2_X1 U8205 ( .A1(n7205), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7204) );
  NAND2_X1 U8206 ( .A1(n14092), .A2(n6878), .ZN(n14093) );
  NAND2_X1 U8207 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n6879), .ZN(n6878) );
  NAND2_X1 U8208 ( .A1(n14097), .A2(n14096), .ZN(n14098) );
  OR2_X1 U8209 ( .A1(n14130), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n14096) );
  XNOR2_X1 U8210 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(n14098), .ZN(n14145) );
  AOI22_X1 U8211 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14150), .B1(n14151), .B2(
        n14101), .ZN(n14103) );
  OAI21_X1 U8212 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n14107), .A(n14106), .ZN(
        n14162) );
  OAI21_X1 U8213 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n14110), .A(n14109), .ZN(
        n14125) );
  AND2_X1 U8214 ( .A1(n6438), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n6674) );
  NOR2_X1 U8215 ( .A1(n6674), .A2(n6675), .ZN(n6670) );
  OR2_X1 U8216 ( .A1(n6438), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n6675) );
  NOR2_X1 U8217 ( .A1(n6674), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n6671) );
  AOI21_X1 U8218 ( .B1(n6915), .B2(n12037), .A(n6557), .ZN(n6914) );
  NAND2_X1 U8219 ( .A1(n6917), .A2(n12037), .ZN(n6916) );
  NOR2_X1 U8220 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8862) );
  AOI21_X1 U8221 ( .B1(n12029), .B2(n12028), .A(n12027), .ZN(n12031) );
  NAND2_X1 U8222 ( .A1(n10158), .A2(n10155), .ZN(n10491) );
  NAND2_X1 U8223 ( .A1(n12006), .A2(n10912), .ZN(n6937) );
  NAND2_X1 U8224 ( .A1(n6925), .A2(n6924), .ZN(n6923) );
  INV_X1 U8225 ( .A(n11969), .ZN(n6924) );
  AOI21_X1 U8226 ( .B1(n6925), .B2(n6922), .A(n6921), .ZN(n6920) );
  NOR2_X1 U8227 ( .A1(n11928), .A2(n12058), .ZN(n6921) );
  NOR2_X1 U8228 ( .A1(n11969), .A2(n6489), .ZN(n6922) );
  NAND2_X1 U8229 ( .A1(n9192), .A2(n12277), .ZN(n12057) );
  NAND2_X1 U8230 ( .A1(n10152), .A2(n6502), .ZN(n10238) );
  OR2_X1 U8231 ( .A1(n11924), .A2(n12056), .ZN(n6928) );
  NAND2_X1 U8232 ( .A1(n12007), .A2(n12008), .ZN(n12006) );
  OR3_X1 U8233 ( .A1(n10126), .A2(n9193), .A3(n12273), .ZN(n12055) );
  NAND2_X1 U8234 ( .A1(n6851), .A2(n6513), .ZN(n6844) );
  NAND2_X1 U8235 ( .A1(n6851), .A2(n6549), .ZN(n6845) );
  AND3_X1 U8236 ( .A1(n9081), .A2(n9080), .A3(n9079), .ZN(n11971) );
  AND2_X1 U8237 ( .A1(n8794), .A2(n8793), .ZN(n12020) );
  AND4_X1 U8238 ( .A1(n9029), .A2(n9028), .A3(n9027), .A4(n9026), .ZN(n11778)
         );
  AND4_X1 U8239 ( .A1(n8954), .A2(n8953), .A3(n8952), .A4(n8951), .ZN(n11459)
         );
  AND4_X1 U8240 ( .A1(n8893), .A2(n8892), .A3(n8891), .A4(n8890), .ZN(n11117)
         );
  NOR2_X1 U8241 ( .A1(n10135), .A2(n15026), .ZN(n10277) );
  NOR2_X1 U8242 ( .A1(n10346), .A2(n10345), .ZN(n10344) );
  AOI21_X1 U8243 ( .B1(P3_REG2_REG_0__SCAN_IN), .B2(n6625), .A(n6503), .ZN(
        n10343) );
  INV_X1 U8244 ( .A(n7287), .ZN(n10292) );
  OR2_X1 U8245 ( .A1(n10276), .A2(n10485), .ZN(n7287) );
  NOR2_X1 U8246 ( .A1(n10305), .A2(n10381), .ZN(n10380) );
  OR2_X1 U8247 ( .A1(n10328), .A2(n10327), .ZN(n10515) );
  AOI21_X1 U8248 ( .B1(n10641), .B2(n10640), .A(n10639), .ZN(n10772) );
  XNOR2_X1 U8249 ( .A(n10955), .B(n14207), .ZN(n10765) );
  NOR2_X1 U8250 ( .A1(n12352), .A2(n14900), .ZN(n12355) );
  AND2_X1 U8251 ( .A1(n12383), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n6817) );
  INV_X1 U8252 ( .A(n7116), .ZN(n14918) );
  INV_X1 U8253 ( .A(n7296), .ZN(n12401) );
  AOI21_X1 U8254 ( .B1(n14913), .B2(n12375), .A(n7294), .ZN(n7296) );
  INV_X1 U8255 ( .A(n7295), .ZN(n7294) );
  AOI21_X1 U8256 ( .B1(n12365), .B2(n12375), .A(n7297), .ZN(n7295) );
  NAND2_X1 U8257 ( .A1(n7122), .A2(n7123), .ZN(n12460) );
  AOI21_X1 U8258 ( .B1(n6466), .B2(n12399), .A(n12424), .ZN(n7123) );
  AOI21_X1 U8259 ( .B1(n7235), .B2(n7238), .A(n6562), .ZN(n7233) );
  OR2_X1 U8260 ( .A1(n9133), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9144) );
  NAND2_X1 U8261 ( .A1(n9103), .A2(n15082), .ZN(n9121) );
  OR2_X1 U8262 ( .A1(n9078), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9091) );
  AND2_X1 U8263 ( .A1(n9066), .A2(n9065), .ZN(n9076) );
  NOR2_X1 U8264 ( .A1(n9053), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9066) );
  OR2_X1 U8265 ( .A1(n9051), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9053) );
  AND2_X1 U8266 ( .A1(n9024), .A2(n11679), .ZN(n9037) );
  NAND2_X1 U8267 ( .A1(n6863), .A2(n12201), .ZN(n6862) );
  OR2_X1 U8268 ( .A1(n6864), .A2(n9250), .ZN(n6863) );
  AND2_X1 U8269 ( .A1(n8918), .A2(n8769), .ZN(n8935) );
  INV_X1 U8270 ( .A(n9245), .ZN(n12177) );
  AND3_X1 U8271 ( .A1(n8900), .A2(n8899), .A3(n8898), .ZN(n8914) );
  AOI21_X1 U8272 ( .B1(n7268), .B2(n12160), .A(n6474), .ZN(n7267) );
  INV_X1 U8273 ( .A(n7268), .ZN(n7266) );
  AND2_X1 U8274 ( .A1(n12112), .A2(n8875), .ZN(n7268) );
  AND2_X1 U8275 ( .A1(n10789), .A2(n8875), .ZN(n11133) );
  NAND2_X1 U8276 ( .A1(n10482), .A2(n8846), .ZN(n10802) );
  NAND2_X1 U8277 ( .A1(n14938), .A2(n14935), .ZN(n9241) );
  NAND2_X1 U8278 ( .A1(n10151), .A2(n9240), .ZN(n14935) );
  INV_X1 U8279 ( .A(n7261), .ZN(n7259) );
  OAI21_X1 U8280 ( .B1(n7261), .B2(n7258), .A(n12256), .ZN(n7257) );
  NAND2_X1 U8281 ( .A1(n6843), .A2(n6842), .ZN(n6835) );
  NAND2_X1 U8282 ( .A1(n6834), .A2(n6843), .ZN(n6833) );
  INV_X1 U8283 ( .A(n12250), .ZN(n12540) );
  AND2_X1 U8284 ( .A1(n12247), .A2(n9255), .ZN(n12551) );
  OAI21_X1 U8285 ( .B1(n6855), .B2(n12238), .A(n12232), .ZN(n6852) );
  AND2_X1 U8286 ( .A1(n6857), .A2(n12232), .ZN(n6854) );
  INV_X1 U8287 ( .A(n11462), .ZN(n14308) );
  AND3_X1 U8288 ( .A1(n8946), .A2(n8945), .A3(n8944), .ZN(n11384) );
  INV_X1 U8289 ( .A(n15001), .ZN(n15014) );
  OR2_X1 U8290 ( .A1(n6606), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7042) );
  AOI21_X1 U8291 ( .B1(n7040), .B2(n7039), .A(n6608), .ZN(n7041) );
  NAND2_X1 U8292 ( .A1(n6622), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9129) );
  INV_X1 U8293 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7272) );
  INV_X1 U8294 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8787) );
  AOI21_X1 U8295 ( .B1(n7030), .B2(n7032), .A(n7028), .ZN(n7027) );
  INV_X1 U8296 ( .A(n8748), .ZN(n7028) );
  NAND2_X1 U8297 ( .A1(n8697), .A2(n8695), .ZN(n7270) );
  OR2_X1 U8298 ( .A1(n8992), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n9020) );
  AND2_X1 U8299 ( .A1(n8735), .A2(n6516), .ZN(n8985) );
  AOI21_X1 U8300 ( .B1(n7053), .B2(n7052), .A(n6561), .ZN(n7051) );
  INV_X1 U8301 ( .A(n8720), .ZN(n7052) );
  XNOR2_X1 U8302 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8910) );
  OR2_X1 U8303 ( .A1(n8908), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8928) );
  XNOR2_X1 U8304 ( .A(n9792), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n8894) );
  NOR2_X1 U8305 ( .A1(n8896), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8906) );
  XNOR2_X1 U8306 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8856) );
  XNOR2_X1 U8307 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8838) );
  NAND2_X1 U8308 ( .A1(n8708), .A2(n8707), .ZN(n8826) );
  OR2_X1 U8309 ( .A1(n10274), .A2(n8973), .ZN(n8824) );
  NAND2_X1 U8310 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8802) );
  NAND2_X1 U8311 ( .A1(n7293), .A2(n8973), .ZN(n7292) );
  NAND2_X1 U8312 ( .A1(n8705), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8813) );
  OR2_X1 U8313 ( .A1(n7794), .A2(n7793), .ZN(n7804) );
  INV_X1 U8314 ( .A(n9739), .ZN(n7189) );
  INV_X1 U8315 ( .A(n9615), .ZN(n7193) );
  NAND2_X1 U8316 ( .A1(n7194), .A2(n6689), .ZN(n7191) );
  INV_X1 U8317 ( .A(n10678), .ZN(n6689) );
  INV_X1 U8318 ( .A(n7897), .ZN(n7895) );
  OR2_X1 U8319 ( .A1(n7846), .A2(n7845), .ZN(n7854) );
  NAND2_X1 U8320 ( .A1(n7853), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7864) );
  INV_X1 U8321 ( .A(n7854), .ZN(n7853) );
  OR2_X1 U8322 ( .A1(n7913), .A2(n12779), .ZN(n7921) );
  AOI21_X1 U8323 ( .B1(n10456), .B2(n10458), .A(n10659), .ZN(n9589) );
  OR2_X1 U8324 ( .A1(n9669), .A2(n6465), .ZN(n6692) );
  OR2_X1 U8325 ( .A1(n7820), .A2(n7819), .ZN(n7828) );
  NAND2_X1 U8326 ( .A1(n7827), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7837) );
  INV_X1 U8327 ( .A(n7828), .ZN(n7827) );
  NAND2_X1 U8328 ( .A1(n7862), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7873) );
  INV_X1 U8329 ( .A(n7864), .ZN(n7862) );
  AND2_X1 U8330 ( .A1(n9667), .A2(n9662), .ZN(n7200) );
  AND2_X1 U8331 ( .A1(n7958), .A2(n7957), .ZN(n12958) );
  AND2_X1 U8332 ( .A1(n7920), .A2(n7919), .ZN(n12846) );
  AND2_X1 U8333 ( .A1(n10104), .A2(n10103), .ZN(n12905) );
  OR2_X1 U8334 ( .A1(n10008), .A2(n10009), .ZN(n10097) );
  NOR2_X1 U8335 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7190) );
  NAND2_X1 U8336 ( .A1(n7198), .A2(n7395), .ZN(n7662) );
  NOR2_X1 U8337 ( .A1(n12993), .A2(n12964), .ZN(n12963) );
  AND2_X1 U8338 ( .A1(n7395), .A2(n7396), .ZN(n7197) );
  INV_X1 U8339 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7396) );
  NAND2_X1 U8340 ( .A1(n13040), .A2(n6823), .ZN(n12993) );
  NOR2_X1 U8341 ( .A1(n12995), .A2(n6824), .ZN(n6823) );
  INV_X1 U8342 ( .A(n6825), .ZN(n6824) );
  INV_X1 U8343 ( .A(n7020), .ZN(n12986) );
  AND2_X1 U8344 ( .A1(n7970), .A2(n7969), .ZN(n12977) );
  AOI21_X1 U8345 ( .B1(n7020), .B2(n6746), .A(n13064), .ZN(n6745) );
  NAND2_X1 U8346 ( .A1(n7959), .A2(n9543), .ZN(n6746) );
  AND2_X1 U8347 ( .A1(n13015), .A2(n13016), .ZN(n7949) );
  NAND2_X1 U8348 ( .A1(n7086), .A2(n7088), .ZN(n13013) );
  AOI21_X1 U8349 ( .B1(n7090), .B2(n7092), .A(n7089), .ZN(n7088) );
  NOR2_X1 U8350 ( .A1(n13038), .A2(n9697), .ZN(n7089) );
  INV_X1 U8351 ( .A(n13015), .ZN(n13012) );
  AND2_X1 U8352 ( .A1(n13070), .A2(n13219), .ZN(n13054) );
  AND2_X1 U8353 ( .A1(n13087), .A2(n13074), .ZN(n13070) );
  NAND2_X1 U8354 ( .A1(n13128), .A2(n7889), .ZN(n7006) );
  OR2_X1 U8355 ( .A1(n11730), .A2(n11704), .ZN(n11723) );
  INV_X1 U8356 ( .A(n7081), .ZN(n7080) );
  AOI21_X1 U8357 ( .B1(n7081), .B2(n7079), .A(n6542), .ZN(n7078) );
  AOI21_X1 U8358 ( .B1(n9534), .B2(n7987), .A(n6525), .ZN(n7081) );
  AND2_X1 U8359 ( .A1(n11562), .A2(n11566), .ZN(n11563) );
  INV_X1 U8360 ( .A(n6822), .ZN(n11157) );
  AOI21_X1 U8361 ( .B1(n10978), .B2(n7071), .A(n6528), .ZN(n7070) );
  INV_X1 U8362 ( .A(n7984), .ZN(n7071) );
  NAND2_X1 U8363 ( .A1(n10982), .A2(n7810), .ZN(n11150) );
  NOR2_X1 U8364 ( .A1(n11149), .A2(n6740), .ZN(n6739) );
  INV_X1 U8365 ( .A(n7810), .ZN(n6740) );
  NOR2_X1 U8366 ( .A1(n11244), .A2(n11227), .ZN(n11229) );
  NAND2_X1 U8367 ( .A1(n11229), .A2(n11210), .ZN(n11209) );
  AND2_X1 U8368 ( .A1(n11223), .A2(n7784), .ZN(n7018) );
  NAND2_X1 U8369 ( .A1(n7785), .A2(n7784), .ZN(n11218) );
  OR2_X1 U8370 ( .A1(n11246), .A2(n11247), .ZN(n11244) );
  NAND2_X1 U8371 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n7757) );
  NAND2_X1 U8372 ( .A1(n10819), .A2(n6993), .ZN(n6992) );
  NOR2_X1 U8373 ( .A1(n6995), .A2(n6996), .ZN(n6993) );
  NAND2_X1 U8374 ( .A1(n6994), .A2(n11266), .ZN(n11271) );
  NAND2_X1 U8375 ( .A1(n10819), .A2(n11268), .ZN(n6994) );
  NAND2_X1 U8376 ( .A1(n7748), .A2(n10814), .ZN(n10819) );
  NAND2_X1 U8377 ( .A1(n10874), .A2(n10820), .ZN(n7748) );
  NAND2_X1 U8378 ( .A1(n10875), .A2(n10876), .ZN(n10874) );
  INV_X1 U8379 ( .A(n9580), .ZN(n10557) );
  OR2_X1 U8380 ( .A1(n12995), .A2(n12977), .ZN(n12969) );
  XNOR2_X1 U8381 ( .A(n12964), .B(n12989), .ZN(n12970) );
  INV_X1 U8382 ( .A(n13038), .ZN(n13214) );
  NAND2_X1 U8383 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n6697), .ZN(n6698) );
  NAND2_X1 U8384 ( .A1(n13296), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n6696) );
  NAND2_X1 U8385 ( .A1(n7513), .A2(n6695), .ZN(n8013) );
  AND2_X1 U8386 ( .A1(n7512), .A2(n7101), .ZN(n6695) );
  NAND2_X1 U8387 ( .A1(n6989), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7407) );
  AND2_X1 U8388 ( .A1(n7389), .A2(n7390), .ZN(n7624) );
  AND2_X1 U8389 ( .A1(n6990), .A2(n7568), .ZN(n7623) );
  OR2_X1 U8390 ( .A1(n7600), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n7607) );
  OR2_X1 U8391 ( .A1(n7592), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n7600) );
  OR2_X1 U8392 ( .A1(n7575), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n7582) );
  OR2_X1 U8393 ( .A1(n7559), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n7566) );
  INV_X1 U8394 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8705) );
  AOI21_X1 U8395 ( .B1(n13423), .B2(n13420), .A(n13460), .ZN(n7136) );
  INV_X1 U8396 ( .A(n7136), .ZN(n7134) );
  AND2_X1 U8397 ( .A1(n10227), .A2(n10223), .ZN(n13476) );
  AND2_X1 U8398 ( .A1(n13412), .A2(n13411), .ZN(n13496) );
  OR2_X1 U8399 ( .A1(n8348), .A2(n8347), .ZN(n8377) );
  NAND2_X1 U8400 ( .A1(n8375), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8397) );
  INV_X1 U8401 ( .A(n8377), .ZN(n8375) );
  NAND2_X1 U8402 ( .A1(n7143), .A2(n7148), .ZN(n13430) );
  NAND2_X1 U8403 ( .A1(n13541), .A2(n7150), .ZN(n7143) );
  AND2_X1 U8404 ( .A1(n7150), .A2(n13524), .ZN(n7147) );
  INV_X1 U8405 ( .A(n13523), .ZN(n7145) );
  INV_X1 U8406 ( .A(n13524), .ZN(n7146) );
  AND2_X1 U8407 ( .A1(n11403), .A2(n11400), .ZN(n7171) );
  NAND2_X1 U8408 ( .A1(n11293), .A2(n11292), .ZN(n11401) );
  INV_X1 U8409 ( .A(n10047), .ZN(n10045) );
  AND2_X1 U8410 ( .A1(n11694), .A2(n11687), .ZN(n7167) );
  OR2_X1 U8411 ( .A1(n8241), .A2(n8240), .ZN(n8259) );
  NAND2_X1 U8412 ( .A1(n13476), .A2(n13475), .ZN(n13474) );
  AND2_X1 U8413 ( .A1(n8596), .A2(n8595), .ZN(n8629) );
  INV_X1 U8414 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15174) );
  XNOR2_X1 U8415 ( .A(P3_IR_REG_0__SCAN_IN), .B(keyinput14), .ZN(n15089) );
  OR2_X1 U8416 ( .A1(n6461), .A2(n8109), .ZN(n8110) );
  AND2_X1 U8417 ( .A1(n14409), .A2(n14410), .ZN(n14407) );
  AND2_X1 U8418 ( .A1(n14413), .A2(n14414), .ZN(n14411) );
  NAND2_X1 U8419 ( .A1(n14422), .A2(n6618), .ZN(n13703) );
  OR2_X1 U8420 ( .A1(n13714), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6618) );
  AOI21_X1 U8421 ( .B1(n13749), .B2(n7349), .A(n6547), .ZN(n7348) );
  INV_X1 U8422 ( .A(n13749), .ZN(n7350) );
  NAND2_X1 U8423 ( .A1(n13835), .A2(n11877), .ZN(n13818) );
  NAND2_X1 U8424 ( .A1(n13873), .A2(n11857), .ZN(n13850) );
  NOR2_X1 U8425 ( .A1(n13909), .A2(n7363), .ZN(n7362) );
  INV_X1 U8426 ( .A(n11854), .ZN(n7363) );
  NAND2_X1 U8427 ( .A1(n13925), .A2(n11854), .ZN(n13908) );
  OR2_X1 U8428 ( .A1(n13944), .A2(n11872), .ZN(n6654) );
  NAND2_X1 U8429 ( .A1(n8332), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8348) );
  INV_X1 U8430 ( .A(n8334), .ZN(n8332) );
  AND4_X1 U8431 ( .A1(n8324), .A2(n8323), .A3(n8322), .A4(n8321), .ZN(n13330)
         );
  NAND2_X1 U8432 ( .A1(n6638), .A2(n6637), .ZN(n11759) );
  AND2_X1 U8433 ( .A1(n6638), .A2(n11641), .ZN(n7382) );
  NAND2_X1 U8434 ( .A1(n11636), .A2(n11642), .ZN(n11763) );
  OR2_X1 U8435 ( .A1(n11693), .A2(n8637), .ZN(n14233) );
  NOR2_X1 U8436 ( .A1(n8278), .A2(n8277), .ZN(n8296) );
  NOR2_X1 U8437 ( .A1(n14347), .A2(n6947), .ZN(n14244) );
  INV_X1 U8438 ( .A(n6949), .ZN(n6947) );
  NOR2_X1 U8439 ( .A1(n14347), .A2(n14373), .ZN(n14349) );
  OR2_X1 U8440 ( .A1(n14494), .A2(n14504), .ZN(n14497) );
  AND2_X1 U8441 ( .A1(n11360), .A2(n11359), .ZN(n11362) );
  AND4_X1 U8442 ( .A1(n8231), .A2(n8230), .A3(n8229), .A4(n8228), .ZN(n11528)
         );
  NAND2_X1 U8443 ( .A1(n11190), .A2(n8633), .ZN(n11351) );
  AND2_X1 U8444 ( .A1(n8173), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8192) );
  NAND2_X1 U8445 ( .A1(n8192), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8215) );
  AND4_X1 U8446 ( .A1(n8220), .A2(n8219), .A3(n8218), .A4(n8217), .ZN(n11407)
         );
  NOR2_X2 U8447 ( .A1(n10841), .A2(n11185), .ZN(n11360) );
  INV_X1 U8448 ( .A(n14533), .ZN(n14507) );
  NAND2_X1 U8449 ( .A1(n14535), .A2(n14556), .ZN(n14517) );
  NOR2_X2 U8450 ( .A1(n14517), .A2(n11339), .ZN(n11335) );
  OR2_X1 U8451 ( .A1(n14534), .A2(n13613), .ZN(n14533) );
  NAND2_X1 U8452 ( .A1(n10407), .A2(n14090), .ZN(n14534) );
  NAND2_X1 U8453 ( .A1(n8576), .A2(n8575), .ZN(n13740) );
  OR2_X1 U8454 ( .A1(n13303), .A2(n8574), .ZN(n8576) );
  AND2_X1 U8455 ( .A1(n13809), .A2(n13808), .ZN(n13994) );
  NAND2_X1 U8456 ( .A1(n8438), .A2(n8437), .ZN(n13879) );
  NAND2_X1 U8457 ( .A1(n8597), .A2(n6769), .ZN(n6768) );
  NAND2_X1 U8458 ( .A1(n6767), .A2(n8566), .ZN(n8598) );
  NAND2_X1 U8459 ( .A1(n6805), .A2(n7502), .ZN(n7715) );
  NAND2_X1 U8460 ( .A1(n6800), .A2(n6806), .ZN(n6805) );
  XNOR2_X1 U8461 ( .A(n7706), .B(n7705), .ZN(n11429) );
  NAND2_X1 U8462 ( .A1(n6784), .A2(n6785), .ZN(n7706) );
  AND2_X1 U8463 ( .A1(n6781), .A2(n6787), .ZN(n6785) );
  XNOR2_X1 U8464 ( .A(n8093), .B(n8092), .ZN(n8624) );
  NAND2_X1 U8465 ( .A1(n8669), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8093) );
  OAI211_X1 U8466 ( .C1(n7676), .C2(n6762), .A(n6758), .B(n6753), .ZN(n7688)
         );
  NAND2_X1 U8467 ( .A1(n7676), .A2(n6483), .ZN(n6753) );
  XNOR2_X1 U8468 ( .A(n7683), .B(n7682), .ZN(n10847) );
  XNOR2_X1 U8469 ( .A(n7647), .B(n7646), .ZN(n10452) );
  NAND2_X1 U8470 ( .A1(n7208), .A2(n7452), .ZN(n7630) );
  NAND2_X1 U8471 ( .A1(n7620), .A2(n7376), .ZN(n7208) );
  OR2_X1 U8472 ( .A1(n8268), .A2(n8267), .ZN(n8283) );
  OR2_X1 U8473 ( .A1(n8197), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n8209) );
  NAND2_X1 U8474 ( .A1(n7212), .A2(n7430), .ZN(n7573) );
  INV_X1 U8475 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8181) );
  NAND2_X1 U8476 ( .A1(n7421), .A2(n7420), .ZN(n7552) );
  XNOR2_X1 U8477 ( .A(n7422), .B(SI_3_), .ZN(n7551) );
  NAND2_X1 U8478 ( .A1(n8104), .A2(n8103), .ZN(n8126) );
  NAND2_X1 U8479 ( .A1(n7433), .A2(n7413), .ZN(n8089) );
  NAND2_X1 U8480 ( .A1(n6877), .A2(n6875), .ZN(n14132) );
  NAND2_X1 U8481 ( .A1(n6876), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n6875) );
  NAND2_X1 U8482 ( .A1(n14134), .A2(n14133), .ZN(n6877) );
  XNOR2_X1 U8483 ( .A(n14145), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n14147) );
  NAND2_X1 U8484 ( .A1(n6655), .A2(n14153), .ZN(n14155) );
  AOI21_X1 U8485 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n10190), .A(n14113), .ZN(
        n14123) );
  NAND2_X1 U8486 ( .A1(n14389), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6885) );
  OR2_X1 U8487 ( .A1(n14389), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6886) );
  NAND2_X1 U8488 ( .A1(n14397), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n6667) );
  OAI22_X1 U8489 ( .A1(n6934), .A2(n6933), .B1(n11675), .B2(n11674), .ZN(
        n14251) );
  NOR2_X1 U8490 ( .A1(n11673), .A2(n12321), .ZN(n6933) );
  INV_X1 U8491 ( .A(n6918), .ZN(n11970) );
  AOI21_X1 U8492 ( .B1(n12019), .B2(n6489), .A(n6919), .ZN(n6918) );
  INV_X1 U8493 ( .A(n6925), .ZN(n6919) );
  AND3_X1 U8494 ( .A1(n8873), .A2(n8872), .A3(n8871), .ZN(n12011) );
  NAND2_X1 U8495 ( .A1(n10491), .A2(n10490), .ZN(n10498) );
  NAND2_X1 U8496 ( .A1(n6937), .A2(n10918), .ZN(n10921) );
  OAI21_X1 U8497 ( .B1(n12019), .B2(n6923), .A(n6920), .ZN(n12038) );
  INV_X1 U8498 ( .A(n6934), .ZN(n11672) );
  NAND2_X1 U8499 ( .A1(n11936), .A2(n6911), .ZN(n12045) );
  AND2_X1 U8500 ( .A1(n10163), .A2(n10162), .ZN(n14884) );
  OAI21_X1 U8501 ( .B1(n12019), .B2(n12018), .A(n6928), .ZN(n12054) );
  NAND2_X1 U8502 ( .A1(n11997), .A2(n11948), .ZN(n12066) );
  INV_X1 U8503 ( .A(n14881), .ZN(n14257) );
  AND2_X1 U8504 ( .A1(n10181), .A2(n10180), .ZN(n14893) );
  AOI21_X1 U8505 ( .B1(n14251), .B2(n14252), .A(n6932), .ZN(n11777) );
  AND2_X1 U8506 ( .A1(n11676), .A2(n12320), .ZN(n6932) );
  AND2_X1 U8507 ( .A1(n10165), .A2(n10164), .ZN(n12062) );
  NOR2_X1 U8508 ( .A1(n12131), .A2(n7048), .ZN(n12132) );
  INV_X1 U8509 ( .A(n11385), .ZN(n12324) );
  AOI21_X1 U8510 ( .B1(n10354), .B2(n10353), .A(n10352), .ZN(n10351) );
  INV_X1 U8511 ( .A(n10293), .ZN(n7286) );
  AND2_X1 U8512 ( .A1(n6811), .A2(n10296), .ZN(n10300) );
  NOR2_X1 U8513 ( .A1(n10512), .A2(n10513), .ZN(n10631) );
  INV_X1 U8514 ( .A(n10646), .ZN(n7107) );
  NAND2_X1 U8515 ( .A1(n6814), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n6813) );
  NAND2_X1 U8516 ( .A1(n10632), .A2(n6814), .ZN(n6812) );
  INV_X1 U8517 ( .A(n10634), .ZN(n6814) );
  OR2_X1 U8518 ( .A1(n10953), .A2(n10761), .ZN(n6816) );
  INV_X1 U8519 ( .A(n12388), .ZN(n7115) );
  NOR2_X1 U8520 ( .A1(n14913), .A2(n12365), .ZN(n12366) );
  NOR2_X1 U8521 ( .A1(n12366), .A2(n12373), .ZN(n12400) );
  XNOR2_X1 U8522 ( .A(n12401), .B(n14266), .ZN(n14262) );
  INV_X1 U8523 ( .A(n7120), .ZN(n14267) );
  INV_X1 U8524 ( .A(n12397), .ZN(n7119) );
  NOR2_X1 U8525 ( .A1(n14261), .A2(n12402), .ZN(n14280) );
  NAND2_X1 U8526 ( .A1(n6477), .A2(n12434), .ZN(n6626) );
  INV_X1 U8527 ( .A(n12456), .ZN(n6815) );
  NAND2_X1 U8528 ( .A1(n12465), .A2(n7127), .ZN(n7126) );
  AND2_X1 U8529 ( .A1(n7240), .A2(n6509), .ZN(n12481) );
  NAND2_X1 U8530 ( .A1(n9132), .A2(n9131), .ZN(n12516) );
  NAND2_X1 U8531 ( .A1(n8768), .A2(n8767), .ZN(n12557) );
  NAND2_X1 U8532 ( .A1(n6861), .A2(n6864), .ZN(n11461) );
  NAND2_X1 U8533 ( .A1(n9248), .A2(n6866), .ZN(n6861) );
  AOI21_X1 U8534 ( .B1(n9248), .B2(n6869), .A(n12186), .ZN(n11371) );
  NAND2_X1 U8535 ( .A1(n11056), .A2(n8917), .ZN(n11376) );
  AND2_X1 U8536 ( .A1(n9295), .A2(n11656), .ZN(n14965) );
  NAND2_X1 U8537 ( .A1(n12088), .A2(n12087), .ZN(n12669) );
  NAND2_X1 U8538 ( .A1(n6846), .A2(n6847), .ZN(n12096) );
  INV_X1 U8539 ( .A(n12516), .ZN(n12685) );
  NOR2_X1 U8540 ( .A1(n12530), .A2(n9111), .ZN(n12521) );
  NAND2_X1 U8541 ( .A1(n6839), .A2(n6837), .ZN(n12519) );
  INV_X1 U8542 ( .A(n6840), .ZN(n6837) );
  NAND2_X1 U8543 ( .A1(n9101), .A2(n9100), .ZN(n12697) );
  AOI21_X1 U8544 ( .B1(n12539), .B2(n12110), .A(n12134), .ZN(n12529) );
  INV_X1 U8545 ( .A(n9096), .ZN(n12703) );
  NAND2_X1 U8546 ( .A1(n9074), .A2(n9073), .ZN(n12714) );
  NAND2_X1 U8547 ( .A1(n7247), .A2(n7244), .ZN(n12563) );
  INV_X1 U8548 ( .A(n7246), .ZN(n7244) );
  INV_X1 U8549 ( .A(n12111), .ZN(n12720) );
  AOI21_X1 U8550 ( .B1(n12590), .B2(n6857), .A(n6855), .ZN(n12570) );
  NAND2_X1 U8551 ( .A1(n8790), .A2(n8789), .ZN(n12726) );
  NAND2_X1 U8552 ( .A1(n6859), .A2(n12233), .ZN(n12578) );
  NAND2_X1 U8553 ( .A1(n9035), .A2(n9034), .ZN(n12738) );
  NAND2_X1 U8554 ( .A1(n9023), .A2(n9022), .ZN(n12745) );
  NAND2_X1 U8555 ( .A1(n11652), .A2(n12121), .ZN(n7228) );
  INV_X1 U8556 ( .A(n12730), .ZN(n12744) );
  INV_X1 U8557 ( .A(n11384), .ZN(n14888) );
  AND2_X1 U8558 ( .A1(n9248), .A2(n9247), .ZN(n11412) );
  INV_X1 U8559 ( .A(n15025), .ZN(n15023) );
  AND2_X1 U8560 ( .A1(n9219), .A2(n9218), .ZN(n12750) );
  AND2_X1 U8561 ( .A1(n6939), .A2(n9215), .ZN(n12752) );
  INV_X1 U8562 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8772) );
  INV_X1 U8563 ( .A(n8778), .ZN(n12760) );
  OAI21_X1 U8564 ( .B1(n9270), .B2(n6603), .A(n9271), .ZN(n11911) );
  XNOR2_X1 U8565 ( .A(n9270), .B(n9172), .ZN(n12763) );
  NAND2_X1 U8566 ( .A1(n7047), .A2(n9086), .ZN(n9099) );
  NAND2_X1 U8567 ( .A1(n9085), .A2(n9084), .ZN(n7047) );
  XNOR2_X1 U8568 ( .A(n8698), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12302) );
  INV_X1 U8569 ( .A(n9259), .ZN(n10537) );
  INV_X1 U8570 ( .A(n12454), .ZN(n12459) );
  NAND2_X1 U8571 ( .A1(n7029), .A2(n8745), .ZN(n9046) );
  NAND2_X1 U8572 ( .A1(n9031), .A2(n8744), .ZN(n7029) );
  INV_X1 U8573 ( .A(SI_12_), .ZN(n15162) );
  NAND2_X1 U8574 ( .A1(n7060), .A2(n6586), .ZN(n8967) );
  NAND2_X1 U8575 ( .A1(n7060), .A2(n8731), .ZN(n8965) );
  CLKBUF_X1 U8576 ( .A(n10143), .Z(n6614) );
  NAND2_X1 U8577 ( .A1(n11895), .A2(n9647), .ZN(n11906) );
  AND2_X1 U8578 ( .A1(n11896), .A2(n9646), .ZN(n9647) );
  NAND2_X1 U8579 ( .A1(n7191), .A2(n7192), .ZN(n10726) );
  NAND2_X1 U8580 ( .A1(n12840), .A2(n9675), .ZN(n12802) );
  NAND2_X1 U8581 ( .A1(n11664), .A2(n9655), .ZN(n11835) );
  INV_X1 U8582 ( .A(n10669), .ZN(n9602) );
  OAI21_X1 U8583 ( .B1(n12785), .B2(n6465), .A(n6469), .ZN(n12840) );
  NAND2_X1 U8584 ( .A1(n12785), .A2(n9669), .ZN(n12837) );
  NAND2_X1 U8585 ( .A1(n11442), .A2(n9639), .ZN(n11449) );
  INV_X1 U8586 ( .A(n13085), .ZN(n13231) );
  INV_X1 U8587 ( .A(n7175), .ZN(n7174) );
  OAI21_X1 U8588 ( .B1(n7177), .B2(n7176), .A(n11254), .ZN(n7175) );
  INV_X1 U8589 ( .A(n9629), .ZN(n7176) );
  NAND2_X1 U8590 ( .A1(n11832), .A2(n9662), .ZN(n12860) );
  NAND2_X1 U8591 ( .A1(n10422), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12856) );
  AND2_X1 U8592 ( .A1(n9734), .A2(n9720), .ZN(n12865) );
  AND2_X1 U8593 ( .A1(n12865), .A2(n13190), .ZN(n12841) );
  INV_X1 U8594 ( .A(n9576), .ZN(n9524) );
  INV_X1 U8595 ( .A(n12958), .ZN(n13018) );
  AND2_X1 U8596 ( .A1(n7745), .A2(n7062), .ZN(n7061) );
  OR2_X1 U8597 ( .A1(n6439), .A2(n7739), .ZN(n7741) );
  OR2_X1 U8598 ( .A1(n6439), .A2(n7729), .ZN(n7731) );
  NAND2_X1 U8599 ( .A1(n9455), .A2(n9454), .ZN(n13188) );
  AND2_X1 U8600 ( .A1(n7522), .A2(n7521), .ZN(n13007) );
  AND2_X1 U8601 ( .A1(n7951), .A2(n7941), .ZN(n13025) );
  OAI211_X1 U8602 ( .C1(n13078), .C2(n6723), .A(n6722), .B(n6731), .ZN(n13034)
         );
  NAND2_X1 U8603 ( .A1(n6725), .A2(n6724), .ZN(n6722) );
  NAND2_X1 U8604 ( .A1(n7087), .A2(n7092), .ZN(n13031) );
  NAND2_X1 U8605 ( .A1(n7098), .A2(n6471), .ZN(n7087) );
  NAND2_X1 U8606 ( .A1(n6726), .A2(n6727), .ZN(n13048) );
  NAND2_X1 U8607 ( .A1(n13078), .A2(n6729), .ZN(n6726) );
  NAND2_X1 U8608 ( .A1(n7097), .A2(n7094), .ZN(n13051) );
  INV_X1 U8609 ( .A(n7096), .ZN(n7094) );
  OR3_X1 U8610 ( .A1(n13087), .A2(n13086), .A3(n13190), .ZN(n13229) );
  NAND2_X1 U8611 ( .A1(n6999), .A2(n7003), .ZN(n13095) );
  NAND2_X1 U8612 ( .A1(n13128), .A2(n6492), .ZN(n6999) );
  NAND2_X1 U8613 ( .A1(n7994), .A2(n7993), .ZN(n13149) );
  NAND2_X1 U8614 ( .A1(n7659), .A2(n7658), .ZN(n13262) );
  NAND2_X1 U8615 ( .A1(n11709), .A2(n7844), .ZN(n11719) );
  INV_X1 U8616 ( .A(n9640), .ZN(n11600) );
  NAND2_X1 U8617 ( .A1(n11552), .A2(n7987), .ZN(n11473) );
  NAND2_X1 U8618 ( .A1(n10979), .A2(n10978), .ZN(n10981) );
  NAND2_X1 U8619 ( .A1(n11206), .A2(n7984), .ZN(n10979) );
  NAND2_X1 U8620 ( .A1(n7077), .A2(n7074), .ZN(n11226) );
  NAND2_X1 U8621 ( .A1(n7077), .A2(n7983), .ZN(n11224) );
  OAI21_X1 U8622 ( .B1(n7980), .B2(n7067), .A(n7065), .ZN(n11038) );
  NAND2_X1 U8623 ( .A1(n7980), .A2(n7979), .ZN(n11023) );
  OR2_X1 U8624 ( .A1(n10816), .A2(n12997), .ZN(n13140) );
  NAND2_X1 U8625 ( .A1(n7009), .A2(n8083), .ZN(n7010) );
  NAND2_X1 U8626 ( .A1(n14767), .A2(n9724), .ZN(n13133) );
  INV_X1 U8627 ( .A(n13178), .ZN(n13143) );
  AND2_X2 U8628 ( .A1(n10552), .A2(n10551), .ZN(n14876) );
  INV_X1 U8629 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n7017) );
  OR2_X1 U8630 ( .A1(n13201), .A2(n14798), .ZN(n13204) );
  NAND2_X1 U8631 ( .A1(n8002), .A2(n8001), .ZN(n8003) );
  NOR2_X1 U8632 ( .A1(n13009), .A2(n6741), .ZN(n8004) );
  INV_X1 U8633 ( .A(n13011), .ZN(n8002) );
  OR3_X1 U8634 ( .A1(n13245), .A2(n13244), .A3(n13243), .ZN(n13288) );
  OR2_X1 U8635 ( .A1(n13251), .A2(n13250), .ZN(n13289) );
  NOR2_X1 U8636 ( .A1(n14733), .A2(n14764), .ZN(n14757) );
  AND2_X1 U8637 ( .A1(n9729), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14767) );
  INV_X1 U8638 ( .A(n14767), .ZN(n14764) );
  INV_X1 U8639 ( .A(n7720), .ZN(n7719) );
  XNOR2_X1 U8640 ( .A(n8006), .B(P2_IR_REG_24__SCAN_IN), .ZN(n11432) );
  NAND2_X1 U8641 ( .A1(n7404), .A2(n7403), .ZN(n7405) );
  NAND2_X1 U8642 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n7402), .ZN(n7403) );
  INV_X1 U8643 ( .A(n9723), .ZN(n10893) );
  INV_X1 U8644 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10471) );
  NAND2_X1 U8645 ( .A1(n7513), .A2(n7391), .ZN(n7648) );
  INV_X1 U8646 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10369) );
  INV_X1 U8647 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10078) );
  INV_X1 U8648 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9926) );
  INV_X1 U8649 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9861) );
  INV_X1 U8650 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9781) );
  INV_X1 U8651 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9767) );
  AND2_X1 U8652 ( .A1(n8682), .A2(n11627), .ZN(n10042) );
  NAND2_X1 U8653 ( .A1(n13422), .A2(n13423), .ZN(n13461) );
  OAI21_X1 U8654 ( .B1(n11401), .B2(n7170), .A(n7168), .ZN(n11614) );
  INV_X1 U8655 ( .A(n7169), .ZN(n7168) );
  OAI21_X1 U8656 ( .B1(n7171), .B2(n7170), .A(n11490), .ZN(n7169) );
  INV_X1 U8657 ( .A(n11484), .ZN(n7170) );
  NAND2_X1 U8658 ( .A1(n11485), .A2(n11484), .ZN(n11491) );
  NAND2_X1 U8659 ( .A1(n10577), .A2(n10576), .ZN(n13444) );
  NAND2_X1 U8660 ( .A1(n11688), .A2(n7167), .ZN(n11807) );
  AND2_X1 U8661 ( .A1(n11688), .A2(n11687), .ZN(n11695) );
  NAND2_X1 U8662 ( .A1(n10593), .A2(n10592), .ZN(n10853) );
  NAND2_X1 U8663 ( .A1(n8370), .A2(n8369), .ZN(n14034) );
  NAND2_X1 U8664 ( .A1(n11401), .A2(n7171), .ZN(n11485) );
  AND2_X1 U8665 ( .A1(n11401), .A2(n11400), .ZN(n11404) );
  NAND2_X1 U8666 ( .A1(n13453), .A2(n13359), .ZN(n13531) );
  NAND2_X1 U8667 ( .A1(n13358), .A2(n13357), .ZN(n13359) );
  OAI21_X1 U8668 ( .B1(n11688), .B2(n7166), .A(n7164), .ZN(n13326) );
  AND2_X1 U8669 ( .A1(n7165), .A2(n11812), .ZN(n7164) );
  OR2_X1 U8670 ( .A1(n7167), .A2(n7166), .ZN(n7165) );
  INV_X1 U8671 ( .A(n11806), .ZN(n7166) );
  NAND2_X1 U8672 ( .A1(n11807), .A2(n11806), .ZN(n11813) );
  AND2_X1 U8673 ( .A1(n8389), .A2(n8388), .ZN(n13553) );
  NAND2_X1 U8674 ( .A1(n7153), .A2(n7156), .ZN(n13550) );
  NAND2_X1 U8675 ( .A1(n7161), .A2(n7157), .ZN(n7153) );
  INV_X1 U8676 ( .A(n14339), .ZN(n13562) );
  INV_X1 U8677 ( .A(n14330), .ZN(n13570) );
  AND2_X1 U8678 ( .A1(n10607), .A2(n9800), .ZN(n10541) );
  AND2_X1 U8679 ( .A1(n9833), .A2(n13613), .ZN(n13929) );
  OR2_X1 U8680 ( .A1(n8650), .A2(n8658), .ZN(n8651) );
  INV_X1 U8681 ( .A(n13755), .ZN(n13790) );
  NAND2_X1 U8682 ( .A1(n8517), .A2(n8516), .ZN(n13583) );
  NAND2_X1 U8683 ( .A1(n8498), .A2(n8497), .ZN(n13819) );
  NAND4_X1 U8684 ( .A1(n8162), .A2(n8161), .A3(n8160), .A4(n8159), .ZN(n13596)
         );
  NAND2_X1 U8685 ( .A1(n8525), .A2(n11169), .ZN(n8162) );
  NAND2_X1 U8686 ( .A1(n8124), .A2(n7371), .ZN(n13598) );
  XNOR2_X1 U8687 ( .A(n13703), .B(n6621), .ZN(n14436) );
  NAND2_X1 U8688 ( .A1(n14436), .A2(n14435), .ZN(n14434) );
  NAND2_X1 U8689 ( .A1(n8064), .A2(n7163), .ZN(n8364) );
  NAND2_X1 U8690 ( .A1(n8622), .A2(n8621), .ZN(n13736) );
  AND2_X1 U8691 ( .A1(n6900), .A2(n6501), .ZN(n13782) );
  NAND2_X1 U8692 ( .A1(n13820), .A2(n7354), .ZN(n13801) );
  AND2_X1 U8693 ( .A1(n13806), .A2(n13805), .ZN(n13995) );
  NAND2_X1 U8694 ( .A1(n13816), .A2(n11879), .ZN(n13804) );
  NAND2_X1 U8695 ( .A1(n13886), .A2(n6894), .ZN(n13876) );
  NOR2_X1 U8696 ( .A1(n6893), .A2(n6472), .ZN(n13877) );
  INV_X1 U8697 ( .A(n13886), .ZN(n6893) );
  INV_X1 U8698 ( .A(n14019), .ZN(n13902) );
  NAND2_X1 U8699 ( .A1(n11786), .A2(n11785), .ZN(n11849) );
  NAND2_X1 U8700 ( .A1(n8361), .A2(n8360), .ZN(n13511) );
  NAND2_X1 U8701 ( .A1(n6635), .A2(n6636), .ZN(n11761) );
  NAND2_X1 U8702 ( .A1(n9851), .A2(n8381), .ZN(n6713) );
  INV_X1 U8703 ( .A(n13963), .ZN(n14512) );
  INV_X1 U8704 ( .A(n10867), .ZN(n14537) );
  INV_X1 U8705 ( .A(n11535), .ZN(n11326) );
  OR2_X1 U8706 ( .A1(n11888), .A2(n6711), .ZN(n6710) );
  OR2_X1 U8707 ( .A1(n14006), .A2(n14005), .ZN(n14060) );
  INV_X1 U8708 ( .A(n13863), .ZN(n14064) );
  OR2_X1 U8709 ( .A1(n14024), .A2(n14023), .ZN(n14069) );
  OR2_X1 U8710 ( .A1(n10068), .A2(n9794), .ZN(n14546) );
  INV_X1 U8711 ( .A(n8058), .ZN(n11844) );
  NAND2_X1 U8712 ( .A1(n8557), .A2(n8556), .ZN(n8565) );
  INV_X1 U8713 ( .A(n6630), .ZN(n6629) );
  NAND2_X1 U8714 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n6631) );
  NAND2_X1 U8715 ( .A1(n8080), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8082) );
  INV_X1 U8716 ( .A(n8624), .ZN(n14090) );
  NAND2_X1 U8717 ( .A1(n8094), .A2(n7347), .ZN(n8069) );
  INV_X1 U8718 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10365) );
  OR2_X1 U8719 ( .A1(n8064), .A2(n8325), .ZN(n8327) );
  INV_X1 U8720 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10367) );
  INV_X1 U8721 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10076) );
  INV_X1 U8722 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9858) );
  INV_X1 U8723 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9852) );
  INV_X1 U8724 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9847) );
  INV_X1 U8725 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9839) );
  INV_X1 U8726 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9792) );
  INV_X1 U8727 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9786) );
  AND2_X1 U8728 ( .A1(n8131), .A2(n8143), .ZN(n13631) );
  INV_X1 U8729 ( .A(n7544), .ZN(n7546) );
  NAND2_X1 U8730 ( .A1(n14137), .A2(n14138), .ZN(n14203) );
  NOR2_X1 U8731 ( .A1(n15203), .A2(n15204), .ZN(n14141) );
  XNOR2_X1 U8732 ( .A(n14148), .B(n14147), .ZN(n15196) );
  XNOR2_X1 U8733 ( .A(n14155), .B(n14636), .ZN(n15200) );
  NAND2_X1 U8734 ( .A1(n6683), .A2(n6681), .ZN(n14228) );
  NAND2_X1 U8735 ( .A1(n6682), .A2(n14167), .ZN(n6681) );
  AND2_X1 U8736 ( .A1(n14167), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n6684) );
  NAND2_X1 U8737 ( .A1(n6680), .A2(n14166), .ZN(n14168) );
  OAI21_X1 U8738 ( .B1(n14176), .B2(n14690), .A(n14399), .ZN(n14404) );
  NAND2_X1 U8739 ( .A1(n6662), .A2(n6660), .ZN(n14176) );
  NAND2_X1 U8740 ( .A1(n6668), .A2(n6661), .ZN(n6660) );
  NAND2_X1 U8741 ( .A1(n12419), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10205) );
  INV_X1 U8742 ( .A(n7289), .ZN(n10951) );
  INV_X1 U8743 ( .A(n7281), .ZN(n14895) );
  INV_X1 U8744 ( .A(n7280), .ZN(n12339) );
  NAND2_X1 U8745 ( .A1(n6613), .A2(n6527), .ZN(P3_U3199) );
  OR2_X1 U8746 ( .A1(n12420), .A2(n14927), .ZN(n6613) );
  MUX2_X1 U8747 ( .A(n12501), .B(n12500), .S(n14963), .Z(n12505) );
  OR2_X1 U8748 ( .A1(n12677), .A2(n12676), .ZN(P3_U3455) );
  MUX2_X1 U8749 ( .A(P3_REG0_REG_28__SCAN_IN), .B(n12673), .S(n15025), .Z(
        n12677) );
  AOI21_X1 U8750 ( .B1(n7184), .B2(n7182), .A(n7180), .ZN(n7179) );
  INV_X1 U8751 ( .A(n7184), .ZN(n7183) );
  INV_X1 U8752 ( .A(n7016), .ZN(n7015) );
  OAI21_X1 U8753 ( .B1(n11848), .B2(n6452), .A(n7201), .ZN(P2_U3305) );
  INV_X1 U8754 ( .A(n7202), .ZN(n7201) );
  OAI22_X1 U8755 ( .A1(n9576), .A2(P2_U3088), .B1(n13314), .B2(n15191), .ZN(
        n7202) );
  MUX2_X1 U8756 ( .A(n13727), .B(n13726), .S(n14536), .Z(n13730) );
  OAI21_X1 U8757 ( .B1(n13976), .B2(n13760), .A(n14543), .ZN(n13766) );
  NOR2_X1 U8758 ( .A1(n11888), .A2(n11889), .ZN(n13985) );
  OAI21_X1 U8759 ( .B1(n14038), .B2(n14595), .A(n6950), .ZN(P1_U3559) );
  INV_X1 U8760 ( .A(n6951), .ZN(n6950) );
  OAI22_X1 U8761 ( .A1(n14041), .A2(n14032), .B1(n14597), .B2(n15085), .ZN(
        n6951) );
  NAND2_X1 U8762 ( .A1(n14388), .A2(n14389), .ZN(n14387) );
  NAND2_X1 U8763 ( .A1(n14392), .A2(n6880), .ZN(n14396) );
  INV_X1 U8764 ( .A(n6676), .ZN(n14249) );
  NOR2_X1 U8765 ( .A1(n14189), .A2(n14188), .ZN(n14197) );
  INV_X2 U8766 ( .A(n9304), .ZN(n9357) );
  AND2_X1 U8767 ( .A1(n12834), .A2(n9671), .ZN(n6465) );
  OAI21_X1 U8768 ( .B1(n12579), .B2(n6856), .A(n12228), .ZN(n6855) );
  NAND2_X1 U8769 ( .A1(n12507), .A2(n9127), .ZN(n12520) );
  INV_X1 U8770 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13296) );
  INV_X2 U8771 ( .A(n6439), .ZN(n9488) );
  INV_X1 U8772 ( .A(n10978), .ZN(n7072) );
  INV_X1 U8773 ( .A(n12485), .ZN(n6849) );
  OR2_X1 U8774 ( .A1(n12425), .A2(n12421), .ZN(n6466) );
  INV_X1 U8775 ( .A(n12190), .ZN(n6868) );
  INV_X1 U8776 ( .A(n11865), .ZN(n7223) );
  AND2_X1 U8777 ( .A1(n10321), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6468) );
  AND2_X1 U8778 ( .A1(n6692), .A2(n12832), .ZN(n6469) );
  INV_X1 U8779 ( .A(n13136), .ZN(n9616) );
  OR2_X1 U8780 ( .A1(n13074), .A2(n12846), .ZN(n6470) );
  AND2_X1 U8781 ( .A1(n6495), .A2(n6470), .ZN(n6471) );
  NOR2_X1 U8782 ( .A1(n14019), .A2(n13488), .ZN(n6472) );
  INV_X1 U8783 ( .A(n11641), .ZN(n6901) );
  NOR2_X1 U8784 ( .A1(n13219), .A2(n13036), .ZN(n6732) );
  INV_X1 U8785 ( .A(n12121), .ZN(n7231) );
  AND2_X1 U8786 ( .A1(n12028), .A2(n11944), .ZN(n6473) );
  AND2_X1 U8787 ( .A1(n12328), .A2(n10905), .ZN(n6474) );
  INV_X1 U8788 ( .A(n8255), .ZN(n7322) );
  XNOR2_X1 U8789 ( .A(n7444), .B(SI_10_), .ZN(n7606) );
  AND2_X1 U8790 ( .A1(n8309), .A2(n7310), .ZN(n6475) );
  AND2_X1 U8791 ( .A1(n10582), .A2(n10576), .ZN(n6476) );
  INV_X1 U8792 ( .A(n11269), .ZN(n11266) );
  NAND2_X1 U8793 ( .A1(n7753), .A2(n11024), .ZN(n11269) );
  INV_X1 U8794 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8761) );
  XOR2_X1 U8795 ( .A(n6505), .B(n6815), .Z(n6477) );
  AND2_X1 U8796 ( .A1(n7250), .A2(n7253), .ZN(n6478) );
  OR2_X1 U8797 ( .A1(n6441), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6479) );
  OR2_X1 U8798 ( .A1(n6468), .A2(n6810), .ZN(n6480) );
  NOR2_X1 U8799 ( .A1(n13197), .A2(n12978), .ZN(n6481) );
  AND2_X1 U8800 ( .A1(n7163), .A2(n7162), .ZN(n6482) );
  AND4_X1 U8801 ( .A1(n12095), .A2(n12094), .A3(n12093), .A4(n12092), .ZN(
        n12107) );
  INV_X1 U8802 ( .A(n12107), .ZN(n6619) );
  INV_X1 U8803 ( .A(n7278), .ZN(n10481) );
  INV_X1 U8804 ( .A(n14397), .ZN(n6666) );
  AND2_X1 U8805 ( .A1(n7477), .A2(SI_20_), .ZN(n6483) );
  AND2_X1 U8806 ( .A1(n7492), .A2(SI_24_), .ZN(n6484) );
  NAND2_X1 U8807 ( .A1(n11098), .A2(n7177), .ZN(n11140) );
  OR2_X1 U8808 ( .A1(n6801), .A2(SI_27_), .ZN(n6485) );
  XNOR2_X1 U8809 ( .A(n12898), .B(n10889), .ZN(n9529) );
  INV_X1 U8810 ( .A(n13505), .ZN(n7161) );
  INV_X1 U8811 ( .A(n13061), .ZN(n7098) );
  AND2_X1 U8812 ( .A1(n7746), .A2(n6479), .ZN(n6487) );
  OR2_X1 U8813 ( .A1(n6441), .A2(n7738), .ZN(n6488) );
  NOR2_X1 U8814 ( .A1(n8051), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n8053) );
  INV_X2 U8815 ( .A(n7796), .ZN(n7964) );
  INV_X1 U8816 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7558) );
  AOI21_X1 U8817 ( .B1(n13541), .B2(n13540), .A(n13539), .ZN(n13431) );
  AND2_X1 U8818 ( .A1(n6929), .A2(n6928), .ZN(n6489) );
  AND2_X1 U8819 ( .A1(n13890), .A2(n11874), .ZN(n6490) );
  AND2_X1 U8820 ( .A1(n7254), .A2(n7251), .ZN(n6491) );
  AND2_X1 U8821 ( .A1(n7007), .A2(n7889), .ZN(n6492) );
  OR2_X1 U8822 ( .A1(n10957), .A2(n10950), .ZN(n6493) );
  OAI21_X1 U8823 ( .B1(n7219), .B2(n14549), .A(n13758), .ZN(n13976) );
  AND2_X1 U8824 ( .A1(n7085), .A2(n7993), .ZN(n6494) );
  NAND2_X1 U8825 ( .A1(n9433), .A2(n13036), .ZN(n6495) );
  NAND2_X1 U8826 ( .A1(n7432), .A2(SI_6_), .ZN(n6496) );
  OR2_X1 U8827 ( .A1(n13246), .A2(n13154), .ZN(n6497) );
  INV_X1 U8828 ( .A(n13236), .ZN(n13103) );
  NAND2_X1 U8829 ( .A1(n7695), .A2(n7694), .ZN(n13236) );
  INV_X1 U8830 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6697) );
  NAND2_X1 U8831 ( .A1(n8094), .A2(n8066), .ZN(n6498) );
  OR2_X1 U8832 ( .A1(n13348), .A2(n13514), .ZN(n6499) );
  OR3_X1 U8833 ( .A1(n12323), .A2(n11513), .A3(n12322), .ZN(n6500) );
  NAND2_X1 U8834 ( .A1(n14052), .A2(n13755), .ZN(n6501) );
  AND2_X1 U8835 ( .A1(n10153), .A2(n10149), .ZN(n6502) );
  NOR2_X1 U8836 ( .A1(n10125), .A2(n14962), .ZN(n6503) );
  INV_X1 U8837 ( .A(n13984), .ZN(n6711) );
  AND2_X1 U8838 ( .A1(n11642), .A2(n7308), .ZN(n6504) );
  XNOR2_X1 U8839 ( .A(n13988), .B(n13583), .ZN(n13789) );
  INV_X1 U8840 ( .A(n13789), .ZN(n6706) );
  OR2_X1 U8841 ( .A1(n12449), .A2(n12448), .ZN(n6505) );
  AOI21_X1 U8842 ( .B1(n13541), .B2(n7147), .A(n7144), .ZN(n13495) );
  XNOR2_X1 U8843 ( .A(n6734), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7724) );
  XNOR2_X1 U8844 ( .A(n12627), .B(n11918), .ZN(n12485) );
  OR2_X1 U8845 ( .A1(n9572), .A2(n12621), .ZN(n6506) );
  OR2_X1 U8846 ( .A1(n9576), .A2(n12997), .ZN(n6507) );
  NAND2_X1 U8847 ( .A1(n8064), .A2(n7380), .ZN(n6508) );
  NAND2_X1 U8848 ( .A1(n12503), .A2(n12309), .ZN(n6509) );
  OR2_X1 U8849 ( .A1(n11516), .A2(n11506), .ZN(n6510) );
  INV_X1 U8850 ( .A(n11858), .ZN(n13861) );
  INV_X1 U8851 ( .A(n9330), .ZN(n6978) );
  INV_X1 U8852 ( .A(n13423), .ZN(n7137) );
  AND2_X1 U8853 ( .A1(n13551), .A2(n7154), .ZN(n6511) );
  AND2_X1 U8854 ( .A1(n7161), .A2(n7160), .ZN(n6512) );
  XNOR2_X1 U8855 ( .A(n13231), .B(n13066), .ZN(n13083) );
  AND2_X1 U8856 ( .A1(n7691), .A2(n7690), .ZN(n13242) );
  INV_X1 U8857 ( .A(n13242), .ZN(n13118) );
  AND2_X1 U8858 ( .A1(n12486), .A2(n6850), .ZN(n6513) );
  OR2_X1 U8859 ( .A1(n12351), .A2(n12336), .ZN(n6514) );
  AND2_X1 U8860 ( .A1(n8762), .A2(n7277), .ZN(n6515) );
  OR2_X1 U8861 ( .A1(n8734), .A2(n10076), .ZN(n6516) );
  XNOR2_X1 U8862 ( .A(n13807), .B(n13565), .ZN(n11865) );
  OR2_X1 U8863 ( .A1(n6440), .A2(n8712), .ZN(n6517) );
  AND2_X1 U8864 ( .A1(n9619), .A2(n9618), .ZN(n6518) );
  INV_X1 U8865 ( .A(n6728), .ZN(n6727) );
  OAI22_X1 U8866 ( .A1(n13062), .A2(n6733), .B1(n13226), .B2(n12846), .ZN(
        n6728) );
  AND2_X1 U8867 ( .A1(n13242), .A2(n12881), .ZN(n6519) );
  AND2_X1 U8868 ( .A1(n6494), .A2(n7996), .ZN(n6520) );
  INV_X1 U8869 ( .A(n14516), .ZN(n14518) );
  NAND3_X1 U8870 ( .A1(n8064), .A2(n7380), .A3(n7364), .ZN(n6521) );
  INV_X1 U8871 ( .A(n12160), .ZN(n8874) );
  AND2_X1 U8872 ( .A1(n12165), .A2(n12164), .ZN(n12160) );
  OR2_X1 U8873 ( .A1(n7262), .A2(n7260), .ZN(n6522) );
  NOR2_X1 U8874 ( .A1(n12418), .A2(n7302), .ZN(n6523) );
  INV_X1 U8875 ( .A(n6946), .ZN(n13826) );
  NOR2_X1 U8876 ( .A1(n12350), .A2(n12349), .ZN(n6524) );
  AND2_X1 U8877 ( .A1(n9640), .A2(n12886), .ZN(n6525) );
  AND2_X1 U8878 ( .A1(n12111), .A2(n12058), .ZN(n6526) );
  NAND2_X1 U8879 ( .A1(n7538), .A2(n6459), .ZN(n7543) );
  INV_X1 U8880 ( .A(n7543), .ZN(n7009) );
  NAND2_X1 U8881 ( .A1(n13040), .A2(n6825), .ZN(n6826) );
  AND2_X1 U8882 ( .A1(n7305), .A2(n6523), .ZN(n6527) );
  AND2_X1 U8883 ( .A1(n14842), .A2(n12889), .ZN(n6528) );
  NAND2_X1 U8884 ( .A1(n11875), .A2(n6490), .ZN(n13886) );
  NOR2_X1 U8885 ( .A1(n14280), .A2(n14279), .ZN(n6529) );
  INV_X1 U8886 ( .A(n9348), .ZN(n6975) );
  AND2_X1 U8887 ( .A1(n7717), .A2(n7716), .ZN(n13028) );
  INV_X1 U8888 ( .A(n13028), .ZN(n13209) );
  INV_X1 U8889 ( .A(n9367), .ZN(n6984) );
  INV_X1 U8890 ( .A(n8458), .ZN(n7335) );
  INV_X1 U8891 ( .A(n8488), .ZN(n7338) );
  INV_X1 U8892 ( .A(n8521), .ZN(n7341) );
  NAND2_X1 U8893 ( .A1(n12691), .A2(n12311), .ZN(n12507) );
  NAND3_X1 U8894 ( .A1(n10204), .A2(n15098), .A3(n7293), .ZN(n6530) );
  OR2_X1 U8895 ( .A1(n9571), .A2(n12489), .ZN(n6531) );
  OR2_X1 U8896 ( .A1(n8207), .A2(n8206), .ZN(n6532) );
  AND2_X1 U8897 ( .A1(n7120), .A2(n7119), .ZN(n6533) );
  AND2_X1 U8898 ( .A1(n11227), .A2(n12891), .ZN(n6534) );
  INV_X1 U8899 ( .A(n7599), .ZN(n7440) );
  XNOR2_X1 U8900 ( .A(n7441), .B(SI_9_), .ZN(n7599) );
  AND2_X1 U8901 ( .A1(n13781), .A2(n6501), .ZN(n6535) );
  AND2_X1 U8902 ( .A1(n6839), .A2(n6838), .ZN(n6536) );
  AND2_X1 U8903 ( .A1(n7097), .A2(n7095), .ZN(n6537) );
  OR2_X1 U8904 ( .A1(n14148), .A2(n14147), .ZN(n6538) );
  AND2_X1 U8905 ( .A1(n12745), .A2(n12319), .ZN(n6539) );
  NOR2_X1 U8906 ( .A1(n12894), .A2(n11032), .ZN(n6540) );
  AND2_X1 U8907 ( .A1(n8345), .A2(n7319), .ZN(n6541) );
  NOR2_X1 U8908 ( .A1(n9640), .A2(n12886), .ZN(n6542) );
  NOR2_X1 U8909 ( .A1(n11253), .A2(n12888), .ZN(n6543) );
  NOR2_X1 U8910 ( .A1(n13936), .A2(n13912), .ZN(n6544) );
  NOR2_X1 U8911 ( .A1(n13879), .A2(n13585), .ZN(n6545) );
  NOR2_X1 U8912 ( .A1(n13103), .A2(n13079), .ZN(n6546) );
  NOR2_X1 U8913 ( .A1(n14052), .A2(n13790), .ZN(n6547) );
  OR2_X1 U8914 ( .A1(n9293), .A2(n10787), .ZN(n12275) );
  AND2_X1 U8915 ( .A1(n13936), .A2(n13912), .ZN(n6548) );
  INV_X1 U8916 ( .A(n6438), .ZN(n6873) );
  NAND2_X1 U8917 ( .A1(n6847), .A2(n12275), .ZN(n6549) );
  AND2_X1 U8918 ( .A1(n13807), .A2(n13565), .ZN(n6550) );
  INV_X1 U8919 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7391) );
  AND2_X1 U8920 ( .A1(n7444), .A2(SI_10_), .ZN(n6551) );
  INV_X1 U8921 ( .A(n6733), .ZN(n6730) );
  NAND2_X1 U8922 ( .A1(n13085), .A2(n12880), .ZN(n6733) );
  AND2_X1 U8923 ( .A1(n14336), .A2(n13588), .ZN(n6552) );
  NAND2_X1 U8924 ( .A1(n7323), .A2(n7320), .ZN(n6553) );
  NOR2_X1 U8925 ( .A1(n13236), .A2(n12848), .ZN(n6554) );
  AND2_X1 U8926 ( .A1(n13033), .A2(n6719), .ZN(n6555) );
  INV_X1 U8927 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8765) );
  AND2_X1 U8928 ( .A1(n6500), .A2(n6935), .ZN(n6556) );
  AND2_X1 U8929 ( .A1(n11930), .A2(n12315), .ZN(n6557) );
  AND2_X1 U8930 ( .A1(n6698), .A2(n6696), .ZN(n6558) );
  AND2_X1 U8931 ( .A1(n8224), .A2(n8223), .ZN(n6559) );
  NAND2_X1 U8932 ( .A1(n7457), .A2(n7645), .ZN(n6560) );
  AND2_X1 U8933 ( .A1(n9792), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n6561) );
  OR2_X1 U8934 ( .A1(n12726), .A2(n12020), .ZN(n12228) );
  NOR2_X1 U8935 ( .A1(n12674), .A2(n11956), .ZN(n6562) );
  NOR2_X1 U8936 ( .A1(n9082), .A2(n11971), .ZN(n6563) );
  NAND2_X1 U8937 ( .A1(n9676), .A2(n9675), .ZN(n6564) );
  AND2_X1 U8938 ( .A1(n7195), .A2(n10568), .ZN(n7194) );
  INV_X1 U8939 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n15168) );
  AND2_X1 U8940 ( .A1(n7125), .A2(n6626), .ZN(n6565) );
  AND2_X1 U8941 ( .A1(n13943), .A2(n11851), .ZN(n6566) );
  AND2_X1 U8942 ( .A1(n7433), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6567) );
  INV_X1 U8943 ( .A(n9250), .ZN(n12119) );
  INV_X1 U8944 ( .A(n11948), .ZN(n6905) );
  NAND2_X1 U8945 ( .A1(n11538), .A2(n8632), .ZN(n14504) );
  NOR2_X1 U8946 ( .A1(n12560), .A2(n7246), .ZN(n7245) );
  AND2_X1 U8947 ( .A1(n6866), .A2(n12119), .ZN(n6568) );
  AND2_X1 U8948 ( .A1(n6912), .A2(n11934), .ZN(n6569) );
  INV_X1 U8949 ( .A(n6732), .ZN(n6731) );
  OR2_X1 U8950 ( .A1(n8190), .A2(n8188), .ZN(n6570) );
  OR2_X1 U8951 ( .A1(n6978), .A2(n9329), .ZN(n6571) );
  OR2_X1 U8952 ( .A1(n9366), .A2(n6984), .ZN(n6572) );
  OR2_X1 U8953 ( .A1(n7335), .A2(n8457), .ZN(n6573) );
  OR2_X1 U8954 ( .A1(n7338), .A2(n8487), .ZN(n6574) );
  OR2_X1 U8955 ( .A1(n7341), .A2(n8520), .ZN(n6575) );
  AND2_X1 U8956 ( .A1(n7091), .A2(n7092), .ZN(n6576) );
  AND2_X1 U8957 ( .A1(n6676), .A2(n6873), .ZN(n6577) );
  OR2_X1 U8958 ( .A1(n9347), .A2(n6975), .ZN(n6578) );
  OR2_X1 U8959 ( .A1(n7332), .A2(n8275), .ZN(n6579) );
  OR2_X1 U8960 ( .A1(n8274), .A2(n8276), .ZN(n6580) );
  AND2_X1 U8961 ( .A1(n7124), .A2(n6466), .ZN(n6581) );
  NAND2_X1 U8962 ( .A1(n7158), .A2(n6499), .ZN(n7156) );
  INV_X1 U8963 ( .A(n11024), .ZN(n6995) );
  OR2_X1 U8964 ( .A1(n12895), .A2(n11280), .ZN(n11024) );
  INV_X1 U8965 ( .A(n7101), .ZN(n7100) );
  AND2_X1 U8966 ( .A1(n7514), .A2(n7102), .ZN(n7101) );
  NAND2_X1 U8967 ( .A1(n7330), .A2(n8602), .ZN(n6582) );
  INV_X1 U8968 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7293) );
  OR2_X1 U8969 ( .A1(n7317), .A2(n6541), .ZN(n6583) );
  INV_X1 U8970 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n15098) );
  INV_X1 U8971 ( .A(n7054), .ZN(n7053) );
  NAND2_X1 U8972 ( .A1(n8721), .A2(n7055), .ZN(n7054) );
  OR2_X1 U8973 ( .A1(n7137), .A2(n7135), .ZN(n6584) );
  INV_X1 U8974 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9744) );
  OR2_X1 U8975 ( .A1(n13730), .A2(n13729), .ZN(P1_U3262) );
  CLKBUF_X3 U8976 ( .A(n8147), .Z(n8381) );
  INV_X2 U8977 ( .A(n8142), .ZN(n8125) );
  NAND2_X1 U8978 ( .A1(n11616), .A2(n11615), .ZN(n11688) );
  NAND2_X1 U8979 ( .A1(n8500), .A2(n8499), .ZN(n13807) );
  INV_X1 U8980 ( .A(n13807), .ZN(n6945) );
  AND2_X1 U8981 ( .A1(n7059), .A2(n8731), .ZN(n6586) );
  INV_X1 U8982 ( .A(n6445), .ZN(n7791) );
  XNOR2_X1 U8983 ( .A(n8870), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10385) );
  INV_X1 U8984 ( .A(n10385), .ZN(n6810) );
  XNOR2_X1 U8985 ( .A(n8897), .B(P3_IR_REG_7__SCAN_IN), .ZN(n10645) );
  INV_X1 U8986 ( .A(n10645), .ZN(n6623) );
  INV_X1 U8987 ( .A(n7759), .ZN(n7796) );
  INV_X1 U8988 ( .A(n6762), .ZN(n6761) );
  NAND2_X1 U8989 ( .A1(n7482), .A2(n10535), .ZN(n6762) );
  INV_X1 U8990 ( .A(n6819), .ZN(n7513) );
  NAND2_X1 U8991 ( .A1(n6467), .A2(n6985), .ZN(n6819) );
  NAND2_X1 U8992 ( .A1(n11640), .A2(n11639), .ZN(n14242) );
  NAND2_X1 U8993 ( .A1(n6654), .A2(n11873), .ZN(n13923) );
  NAND2_X1 U8994 ( .A1(n11790), .A2(n11789), .ZN(n11869) );
  NAND2_X1 U8995 ( .A1(n7228), .A2(n9017), .ZN(n12613) );
  OR2_X1 U8996 ( .A1(n6945), .A2(n14032), .ZN(n6587) );
  NAND2_X1 U8997 ( .A1(n12082), .A2(n12081), .ZN(n12665) );
  INV_X1 U8998 ( .A(n12665), .ZN(n6620) );
  NAND2_X1 U8999 ( .A1(n11875), .A2(n11874), .ZN(n13887) );
  OR2_X1 U9000 ( .A1(n7273), .A2(n7270), .ZN(n9047) );
  INV_X1 U9001 ( .A(n6944), .ZN(n13955) );
  NOR2_X1 U9002 ( .A1(n13898), .A2(n13879), .ZN(n6617) );
  INV_X1 U9003 ( .A(n9401), .ZN(n6981) );
  INV_X1 U9004 ( .A(n9418), .ZN(n6965) );
  AND2_X1 U9005 ( .A1(n7116), .A2(n7115), .ZN(n6588) );
  INV_X1 U9006 ( .A(n9427), .ZN(n6972) );
  AND2_X1 U9007 ( .A1(n9460), .A2(n9459), .ZN(n13202) );
  INV_X1 U9008 ( .A(n13202), .ZN(n12995) );
  NAND2_X1 U9009 ( .A1(n7255), .A2(n7254), .ZN(n7250) );
  AND3_X1 U9010 ( .A1(n9095), .A2(n9094), .A3(n9093), .ZN(n11964) );
  INV_X1 U9011 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8712) );
  AND3_X1 U9012 ( .A1(n14392), .A2(n6880), .A3(n6666), .ZN(n6589) );
  AND2_X1 U9013 ( .A1(n6859), .A2(n6857), .ZN(n6590) );
  OR2_X1 U9014 ( .A1(n6981), .A2(n9400), .ZN(n6591) );
  INV_X1 U9015 ( .A(n6787), .ZN(n6786) );
  AND2_X1 U9016 ( .A1(n6788), .A2(n6791), .ZN(n6787) );
  INV_X1 U9017 ( .A(n14589), .ZN(n6712) );
  NAND2_X1 U9018 ( .A1(n8395), .A2(n8394), .ZN(n13936) );
  INV_X1 U9019 ( .A(n13936), .ZN(n6943) );
  AND2_X2 U9020 ( .A1(n10552), .A2(n14763), .ZN(n14858) );
  OR2_X1 U9021 ( .A1(n8008), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n6592) );
  AND2_X1 U9022 ( .A1(n14931), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n6593) );
  NAND2_X1 U9023 ( .A1(n10790), .A2(n8874), .ZN(n10789) );
  NAND2_X1 U9024 ( .A1(n7513), .A2(n7512), .ZN(n8008) );
  NAND2_X1 U9025 ( .A1(n11352), .A2(n11190), .ZN(n11191) );
  OR2_X1 U9026 ( .A1(n14347), .A2(n6948), .ZN(n6594) );
  NAND2_X1 U9027 ( .A1(n10789), .A2(n7268), .ZN(n11132) );
  AND2_X1 U9028 ( .A1(n12229), .A2(n12233), .ZN(n12591) );
  AND2_X1 U9029 ( .A1(n14497), .A2(n11538), .ZN(n6595) );
  INV_X1 U9030 ( .A(n6820), .ZN(n11562) );
  NAND2_X1 U9031 ( .A1(n6822), .A2(n6821), .ZN(n6820) );
  NOR2_X1 U9032 ( .A1(n14858), .A2(n7017), .ZN(n6596) );
  INV_X1 U9033 ( .A(n7253), .ZN(n7252) );
  NAND2_X1 U9034 ( .A1(n9058), .A2(n12020), .ZN(n7253) );
  AND2_X1 U9035 ( .A1(n15191), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6597) );
  NAND2_X1 U9036 ( .A1(n6806), .A2(n6799), .ZN(n6598) );
  NAND2_X1 U9037 ( .A1(n7502), .A2(SI_26_), .ZN(n6804) );
  AND2_X1 U9038 ( .A1(n8752), .A2(n10894), .ZN(n6599) );
  AND2_X1 U9039 ( .A1(n11098), .A2(n9624), .ZN(n6600) );
  AND2_X1 U9040 ( .A1(n7289), .A2(n6493), .ZN(n6601) );
  AND2_X1 U9041 ( .A1(n7108), .A2(n7107), .ZN(n6602) );
  INV_X1 U9042 ( .A(n14588), .ZN(n14549) );
  INV_X1 U9043 ( .A(n12997), .ZN(n11725) );
  NAND2_X1 U9044 ( .A1(n9492), .A2(n7960), .ZN(n13169) );
  INV_X1 U9045 ( .A(n10727), .ZN(n7196) );
  NAND2_X1 U9046 ( .A1(n7619), .A2(n7618), .ZN(n11253) );
  INV_X1 U9047 ( .A(n11253), .ZN(n6821) );
  NAND2_X1 U9048 ( .A1(n10245), .A2(n10246), .ZN(n10158) );
  AND2_X1 U9049 ( .A1(n11917), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6603) );
  INV_X1 U9050 ( .A(SI_24_), .ZN(n6793) );
  OR2_X1 U9051 ( .A1(n14597), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6604) );
  OR2_X1 U9052 ( .A1(n14589), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6605) );
  OR2_X1 U9053 ( .A1(n10041), .A2(n14537), .ZN(n14526) );
  AND2_X1 U9054 ( .A1(n11505), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6606) );
  AND2_X1 U9055 ( .A1(n9561), .A2(n12105), .ZN(n14939) );
  NAND2_X1 U9056 ( .A1(n8831), .A2(n8830), .ZN(n10480) );
  AND2_X1 U9057 ( .A1(n7287), .A2(n7286), .ZN(n6607) );
  AND2_X1 U9058 ( .A1(n11502), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U9059 ( .A1(n8286), .A2(n8285), .ZN(n11693) );
  NOR2_X1 U9060 ( .A1(n10631), .A2(n10632), .ZN(n6609) );
  INV_X1 U9061 ( .A(n14437), .ZN(n6621) );
  INV_X1 U9062 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6876) );
  INV_X1 U9063 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6685) );
  INV_X1 U9064 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6879) );
  INV_X1 U9065 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6686) );
  AOI21_X1 U9066 ( .B1(n13773), .B2(n14519), .A(n13772), .ZN(n13982) );
  INV_X1 U9067 ( .A(n14519), .ZN(n14548) );
  NAND2_X1 U9068 ( .A1(n13997), .A2(n6587), .ZN(P1_U3553) );
  NAND2_X1 U9069 ( .A1(n10836), .A2(n10835), .ZN(n11183) );
  NOR2_X2 U9070 ( .A1(n8080), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n8078) );
  NAND2_X1 U9071 ( .A1(n6940), .A2(n7380), .ZN(n8080) );
  NAND2_X1 U9072 ( .A1(n14529), .A2(n11339), .ZN(n10405) );
  NAND2_X2 U9073 ( .A1(n13927), .A2(n13926), .ZN(n13925) );
  NAND2_X1 U9074 ( .A1(n6612), .A2(n11115), .ZN(n10916) );
  NAND2_X1 U9075 ( .A1(n10930), .A2(n11118), .ZN(n6612) );
  NAND2_X1 U9076 ( .A1(n6909), .A2(n11935), .ZN(n11936) );
  OAI22_X1 U9077 ( .A1(n11777), .A2(n11776), .B1(n11778), .B2(n11775), .ZN(
        n11923) );
  NOR2_X1 U9078 ( .A1(n11939), .A2(n11940), .ZN(n11961) );
  OAI21_X1 U9079 ( .B1(n12019), .B2(n6916), .A(n6914), .ZN(n6913) );
  NOR2_X1 U9080 ( .A1(n15040), .A2(n10765), .ZN(n10958) );
  NOR2_X1 U9081 ( .A1(n10323), .A2(n10380), .ZN(n10328) );
  NAND2_X1 U9082 ( .A1(n10646), .A2(n7105), .ZN(n7104) );
  NOR2_X1 U9083 ( .A1(n10318), .A2(n10319), .ZN(n10436) );
  AOI21_X1 U9084 ( .B1(P3_REG1_REG_4__SCAN_IN), .B2(n10321), .A(n10434), .ZN(
        n10322) );
  AOI22_X1 U9085 ( .A1(n13114), .A2(n7997), .B1(n13118), .B2(n12881), .ZN(
        n13105) );
  NAND2_X1 U9086 ( .A1(n7986), .A2(n7985), .ZN(n11551) );
  OAI21_X1 U9087 ( .B1(n13198), .B2(n14798), .A(n6481), .ZN(n6830) );
  NAND2_X1 U9088 ( .A1(n7140), .A2(n7138), .ZN(n13494) );
  AND4_X2 U9089 ( .A1(n8047), .A2(n8046), .A3(n8045), .A4(n8044), .ZN(n7380)
         );
  INV_X1 U9090 ( .A(n13598), .ZN(n10231) );
  NAND2_X1 U9091 ( .A1(n13558), .A2(n13421), .ZN(n13422) );
  INV_X1 U9092 ( .A(n13443), .ZN(n10582) );
  NAND2_X2 U9093 ( .A1(n13484), .A2(n13483), .ZN(n13541) );
  NAND2_X1 U9094 ( .A1(n13333), .A2(n13332), .ZN(n14332) );
  NAND2_X1 U9095 ( .A1(n8729), .A2(n8728), .ZN(n8958) );
  NAND2_X1 U9096 ( .A1(n8785), .A2(n8750), .ZN(n9060) );
  INV_X1 U9097 ( .A(n9129), .ZN(n7040) );
  NAND2_X1 U9098 ( .A1(n8738), .A2(n8737), .ZN(n9019) );
  INV_X1 U9099 ( .A(n9117), .ZN(n6622) );
  NAND2_X1 U9100 ( .A1(n8723), .A2(n8722), .ZN(n8925) );
  NAND2_X1 U9101 ( .A1(n8726), .A2(n8725), .ZN(n8942) );
  OAI21_X1 U9102 ( .B1(n8885), .B2(n7054), .A(n7051), .ZN(n8911) );
  NAND2_X1 U9103 ( .A1(n8742), .A2(n8741), .ZN(n9031) );
  NAND3_X1 U9104 ( .A1(n12276), .A2(n6615), .A3(n12271), .ZN(n12282) );
  OAI21_X1 U9105 ( .B1(n9128), .B2(n7042), .A(n7041), .ZN(n9151) );
  OAI21_X2 U9106 ( .B1(n9072), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n8753), .ZN(
        n9085) );
  OR2_X2 U9107 ( .A1(n13744), .A2(n13740), .ZN(n13738) );
  NAND2_X1 U9108 ( .A1(n13776), .A2(n13970), .ZN(n13744) );
  INV_X1 U9109 ( .A(n6617), .ZN(n13878) );
  NAND2_X1 U9110 ( .A1(n6628), .A2(n6627), .ZN(n11769) );
  NAND2_X1 U9111 ( .A1(n6952), .A2(n14508), .ZN(n13964) );
  OAI21_X1 U9112 ( .B1(n7129), .B2(n14927), .A(n6565), .ZN(P3_U3201) );
  AOI21_X1 U9113 ( .B1(n12468), .B2(n14924), .A(n7126), .ZN(n7125) );
  NOR2_X2 U9114 ( .A1(n14905), .A2(n14904), .ZN(n14903) );
  NOR2_X1 U9115 ( .A1(n9975), .A2(n9976), .ZN(n9974) );
  NOR2_X1 U9116 ( .A1(n9940), .A2(n9941), .ZN(n10186) );
  NOR2_X1 U9117 ( .A1(n9963), .A2(n9964), .ZN(n9962) );
  AOI21_X1 U9118 ( .B1(n13712), .B2(P1_REG1_REG_13__SCAN_IN), .A(n14407), .ZN(
        n14424) );
  NOR2_X1 U9119 ( .A1(n9987), .A2(n9988), .ZN(n9986) );
  NOR2_X1 U9120 ( .A1(n10188), .A2(n10189), .ZN(n13701) );
  AOI21_X1 U9121 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n14473), .A(n14468), .ZN(
        n13705) );
  AOI21_X1 U9122 ( .B1(n13717), .B2(P1_REG1_REG_16__SCAN_IN), .A(n14454), .ZN(
        n14470) );
  NAND2_X1 U9123 ( .A1(n8985), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8988) );
  NAND2_X1 U9124 ( .A1(n8925), .A2(n8724), .ZN(n8726) );
  NAND2_X1 U9125 ( .A1(n8714), .A2(n8713), .ZN(n8857) );
  NAND2_X1 U9126 ( .A1(n8711), .A2(n8710), .ZN(n8839) );
  NAND2_X1 U9127 ( .A1(n8716), .A2(n8715), .ZN(n8869) );
  NAND2_X1 U9128 ( .A1(n9004), .A2(n9003), .ZN(n8738) );
  NAND2_X1 U9129 ( .A1(n8911), .A2(n8910), .ZN(n8723) );
  NOR2_X1 U9130 ( .A1(n12131), .A2(n12100), .ZN(n12283) );
  XNOR2_X2 U9131 ( .A(n8084), .B(P1_IR_REG_1__SCAN_IN), .ZN(n13602) );
  NAND2_X1 U9132 ( .A1(n12460), .A2(n12461), .ZN(n12464) );
  INV_X1 U9133 ( .A(n6624), .ZN(n10644) );
  NAND2_X1 U9134 ( .A1(n7552), .A2(n7551), .ZN(n6701) );
  NOR2_X2 U9135 ( .A1(n13774), .A2(n13980), .ZN(n13776) );
  NAND2_X1 U9136 ( .A1(n13916), .A2(n14019), .ZN(n13898) );
  NOR2_X2 U9137 ( .A1(n11769), .A2(n14362), .ZN(n11791) );
  NOR2_X2 U9138 ( .A1(n14347), .A2(n14336), .ZN(n6627) );
  XOR2_X1 U9139 ( .A(n13736), .B(n13738), .Z(n6952) );
  XNOR2_X1 U9140 ( .A(n12464), .B(n12463), .ZN(n7129) );
  NOR2_X1 U9141 ( .A1(n10277), .A2(n10278), .ZN(n10346) );
  NAND2_X1 U9142 ( .A1(n12397), .A2(n7121), .ZN(n7117) );
  OAI22_X1 U9143 ( .A1(n8078), .A2(n6631), .B1(P1_IR_REG_31__SCAN_IN), .B2(
        P1_IR_REG_28__SCAN_IN), .ZN(n6630) );
  NAND2_X1 U9144 ( .A1(n6635), .A2(n6632), .ZN(n11790) );
  NAND2_X1 U9145 ( .A1(n15200), .A2(n15201), .ZN(n14156) );
  NAND2_X1 U9146 ( .A1(n14212), .A2(n14211), .ZN(n6655) );
  INV_X1 U9147 ( .A(n14385), .ZN(n6657) );
  AND2_X1 U9148 ( .A1(n14170), .A2(n14171), .ZN(n14384) );
  NOR2_X1 U9149 ( .A1(n14169), .A2(n14229), .ZN(n14170) );
  NAND3_X1 U9150 ( .A1(n14392), .A2(n6880), .A3(n6667), .ZN(n6659) );
  INV_X1 U9151 ( .A(n6665), .ZN(n6661) );
  NAND3_X1 U9152 ( .A1(n14392), .A2(n6880), .A3(n6663), .ZN(n6662) );
  INV_X1 U9153 ( .A(n14401), .ZN(n6668) );
  NAND2_X1 U9154 ( .A1(n14177), .A2(n14702), .ZN(n6677) );
  INV_X1 U9155 ( .A(n14403), .ZN(n6678) );
  NAND2_X1 U9156 ( .A1(n14403), .A2(n6673), .ZN(n6672) );
  NAND2_X1 U9157 ( .A1(n14227), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n6680) );
  NAND2_X1 U9158 ( .A1(n14227), .A2(n6684), .ZN(n6683) );
  NAND2_X1 U9159 ( .A1(n12785), .A2(n6469), .ZN(n6690) );
  NAND2_X1 U9160 ( .A1(n6690), .A2(n6691), .ZN(n12800) );
  NAND2_X1 U9161 ( .A1(n12864), .A2(n9708), .ZN(n12767) );
  OAI21_X2 U9162 ( .B1(n11098), .B2(n7176), .A(n7174), .ZN(n11258) );
  INV_X1 U9163 ( .A(n6440), .ZN(n9485) );
  NAND3_X1 U9164 ( .A1(n6700), .A2(n6699), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n6887) );
  NAND2_X1 U9165 ( .A1(n7415), .A2(n7535), .ZN(n6748) );
  NAND2_X1 U9166 ( .A1(n6458), .A2(n7414), .ZN(n7532) );
  NAND2_X1 U9167 ( .A1(n7590), .A2(n7437), .ZN(n6702) );
  NAND2_X1 U9168 ( .A1(n7580), .A2(n7434), .ZN(n6703) );
  NAND2_X1 U9169 ( .A1(n6704), .A2(n6566), .ZN(n13950) );
  OAI21_X1 U9170 ( .B1(n11863), .B2(n7353), .A(n6708), .ZN(n13788) );
  NAND2_X1 U9171 ( .A1(n11863), .A2(n6708), .ZN(n6707) );
  AND2_X2 U9172 ( .A1(n11863), .A2(n11862), .ZN(n13822) );
  NAND2_X1 U9173 ( .A1(n7351), .A2(n6714), .ZN(n14341) );
  AOI21_X1 U9174 ( .B1(n14504), .B2(n11538), .A(n14346), .ZN(n6714) );
  NAND2_X1 U9175 ( .A1(n11039), .A2(n7774), .ZN(n11239) );
  NAND2_X1 U9176 ( .A1(n6721), .A2(n13078), .ZN(n6720) );
  NOR2_X2 U9177 ( .A1(n7511), .A2(n7510), .ZN(n7512) );
  AND4_X1 U9178 ( .A1(n7512), .A2(n7099), .A3(n6985), .A4(n6467), .ZN(n7518)
         );
  AND2_X1 U9179 ( .A1(n6765), .A2(n6768), .ZN(n8569) );
  NAND3_X1 U9180 ( .A1(n8557), .A2(n6766), .A3(n8556), .ZN(n6765) );
  NAND3_X1 U9181 ( .A1(n8557), .A2(n8556), .A3(n6770), .ZN(n6767) );
  NAND2_X1 U9182 ( .A1(n7613), .A2(n6774), .ZN(n6773) );
  NAND2_X1 U9183 ( .A1(n7697), .A2(n7492), .ZN(n6794) );
  INV_X1 U9184 ( .A(n7710), .ZN(n6800) );
  NOR2_X1 U9185 ( .A1(n10432), .A2(n6468), .ZN(n10295) );
  NAND3_X1 U9186 ( .A1(n6808), .A2(n6809), .A3(n6807), .ZN(n10371) );
  NAND4_X1 U9187 ( .A1(n6808), .A2(n6809), .A3(n6807), .A4(
        P3_REG2_REG_5__SCAN_IN), .ZN(n6811) );
  INV_X1 U9188 ( .A(n6811), .ZN(n10370) );
  OAI21_X1 U9189 ( .B1(n10512), .B2(n6813), .A(n6812), .ZN(n10759) );
  INV_X1 U9190 ( .A(n6826), .ZN(n12992) );
  NOR2_X1 U9191 ( .A1(n13172), .A2(n13253), .ZN(n6829) );
  INV_X1 U9192 ( .A(n6829), .ZN(n13158) );
  NOR2_X2 U9193 ( .A1(n13195), .A2(n6830), .ZN(n7016) );
  NAND2_X1 U9194 ( .A1(n11063), .A2(n12177), .ZN(n6831) );
  NAND2_X1 U9195 ( .A1(n11011), .A2(n12171), .ZN(n6832) );
  INV_X1 U9196 ( .A(n12539), .ZN(n6836) );
  OAI21_X2 U9197 ( .B1(n6836), .B2(n6835), .A(n6833), .ZN(n12506) );
  NAND2_X1 U9198 ( .A1(n12486), .A2(n6850), .ZN(n6846) );
  NAND2_X1 U9199 ( .A1(n6844), .A2(n6845), .ZN(n12102) );
  NOR2_X1 U9200 ( .A1(n12486), .A2(n12485), .ZN(n12484) );
  NAND2_X1 U9201 ( .A1(n12590), .A2(n6854), .ZN(n6853) );
  AOI21_X1 U9202 ( .B1(n9248), .B2(n6568), .A(n6862), .ZN(n11584) );
  AND2_X2 U9203 ( .A1(n8760), .A2(n8759), .ZN(n9206) );
  NAND2_X1 U9204 ( .A1(n14388), .A2(n6886), .ZN(n6884) );
  NAND2_X1 U9205 ( .A1(n6884), .A2(n6882), .ZN(n6881) );
  NAND3_X1 U9206 ( .A1(n12948), .A2(P3_ADDR_REG_19__SCAN_IN), .A3(n6889), .ZN(
        n6888) );
  INV_X1 U9207 ( .A(n11339), .ZN(n14564) );
  OR2_X1 U9208 ( .A1(n8574), .A2(n9747), .ZN(n6895) );
  NAND2_X1 U9209 ( .A1(n13599), .A2(n14564), .ZN(n8116) );
  XNOR2_X1 U9210 ( .A(n7546), .B(n7545), .ZN(n9747) );
  NAND2_X1 U9211 ( .A1(n13786), .A2(n6898), .ZN(n6900) );
  NAND2_X1 U9212 ( .A1(n13786), .A2(n11881), .ZN(n11886) );
  NAND2_X1 U9213 ( .A1(n6902), .A2(n6903), .ZN(n12065) );
  NAND3_X1 U9214 ( .A1(n6473), .A2(n11948), .A3(n12029), .ZN(n6902) );
  NAND3_X1 U9215 ( .A1(n11936), .A2(n6911), .A3(n11964), .ZN(n6910) );
  NAND2_X1 U9216 ( .A1(n11989), .A2(n11934), .ZN(n6909) );
  NAND2_X1 U9217 ( .A1(n11989), .A2(n6569), .ZN(n6911) );
  INV_X1 U9218 ( .A(n6910), .ZN(n12044) );
  INV_X1 U9219 ( .A(n11935), .ZN(n6912) );
  INV_X1 U9220 ( .A(n6913), .ZN(n11990) );
  MUX2_X1 U9221 ( .A(n9240), .B(n10148), .S(n11931), .Z(n10153) );
  INV_X1 U9222 ( .A(n10497), .ZN(n6931) );
  NAND2_X1 U9223 ( .A1(n9212), .A2(n11499), .ZN(n6938) );
  NAND3_X1 U9224 ( .A1(n6938), .A2(n9213), .A3(n9217), .ZN(n6939) );
  AND4_X2 U9225 ( .A1(n8041), .A2(n8040), .A3(n8269), .A4(n8183), .ZN(n6941)
         );
  AND3_X2 U9226 ( .A1(n6941), .A2(n8182), .A3(n6942), .ZN(n8064) );
  AND4_X2 U9227 ( .A1(n6941), .A2(n7365), .A3(n8182), .A4(n6942), .ZN(n6940)
         );
  AND4_X2 U9228 ( .A1(n8303), .A2(n8266), .A3(n8232), .A4(n8311), .ZN(n6942)
         );
  AND2_X1 U9229 ( .A1(n11312), .A2(n14569), .ZN(n11314) );
  AND2_X2 U9230 ( .A1(n11335), .A2(n11079), .ZN(n11312) );
  NOR2_X2 U9231 ( .A1(n13878), .A2(n13863), .ZN(n13860) );
  NOR2_X1 U9232 ( .A1(n11693), .A2(n14373), .ZN(n6949) );
  AND2_X2 U9233 ( .A1(n13964), .A2(n13965), .ZN(n14038) );
  NAND2_X1 U9234 ( .A1(n9303), .A2(n6953), .ZN(n9304) );
  NOR2_X1 U9235 ( .A1(n9302), .A2(n11725), .ZN(n10812) );
  AOI21_X1 U9236 ( .B1(n9576), .B2(n6953), .A(n9518), .ZN(n9519) );
  XNOR2_X1 U9237 ( .A(n9576), .B(n6953), .ZN(n8000) );
  OAI22_X2 U9238 ( .A1(n9389), .A2(n6955), .B1(n9390), .B2(n6954), .ZN(n9394)
         );
  NAND2_X1 U9239 ( .A1(n9413), .A2(n6961), .ZN(n6960) );
  NAND3_X1 U9240 ( .A1(n6960), .A2(n6958), .A3(n6962), .ZN(n9422) );
  NAND2_X1 U9241 ( .A1(n9382), .A2(n9383), .ZN(n9381) );
  NAND2_X1 U9242 ( .A1(n9426), .A2(n6971), .ZN(n6968) );
  NAND2_X1 U9243 ( .A1(n6968), .A2(n6969), .ZN(n9430) );
  NAND2_X1 U9244 ( .A1(n6973), .A2(n6974), .ZN(n9351) );
  NAND3_X1 U9245 ( .A1(n9346), .A2(n6578), .A3(n9345), .ZN(n6973) );
  NAND2_X1 U9246 ( .A1(n6976), .A2(n6977), .ZN(n9333) );
  NAND3_X1 U9247 ( .A1(n9328), .A2(n9327), .A3(n6571), .ZN(n6976) );
  NAND3_X1 U9248 ( .A1(n9399), .A2(n9398), .A3(n6591), .ZN(n6979) );
  NAND2_X1 U9249 ( .A1(n6979), .A2(n6980), .ZN(n9405) );
  NAND2_X1 U9250 ( .A1(n6982), .A2(n6983), .ZN(n9370) );
  NAND3_X1 U9251 ( .A1(n9365), .A2(n9364), .A3(n6572), .ZN(n6982) );
  INV_X1 U9252 ( .A(n7655), .ZN(n7394) );
  NAND3_X1 U9253 ( .A1(n6467), .A2(n6985), .A3(n7190), .ZN(n7655) );
  AND4_X2 U9254 ( .A1(n7540), .A2(n7621), .A3(n6987), .A4(n6986), .ZN(n6985)
         );
  NAND2_X1 U9255 ( .A1(n7198), .A2(n6988), .ZN(n6989) );
  INV_X1 U9256 ( .A(n6989), .ZN(n7406) );
  NAND2_X1 U9257 ( .A1(n7860), .A2(n11741), .ZN(n11745) );
  NAND2_X1 U9258 ( .A1(n11269), .A2(n11024), .ZN(n6991) );
  NAND3_X1 U9259 ( .A1(n7067), .A2(n6992), .A3(n6991), .ZN(n11027) );
  NAND2_X1 U9260 ( .A1(n13128), .A2(n7000), .ZN(n6998) );
  INV_X1 U9261 ( .A(n7888), .ZN(n7008) );
  NAND2_X1 U9262 ( .A1(n7538), .A2(n6567), .ZN(n7011) );
  NAND3_X2 U9263 ( .A1(n7542), .A2(n7011), .A3(n7010), .ZN(n10889) );
  NAND2_X1 U9264 ( .A1(n11709), .A2(n7012), .ZN(n11717) );
  NAND2_X1 U9265 ( .A1(n12980), .A2(n7016), .ZN(n13280) );
  OAI21_X1 U9266 ( .B1(n12980), .B2(n14856), .A(n7014), .ZN(P2_U3496) );
  NAND2_X1 U9267 ( .A1(n12980), .A2(n12979), .ZN(n13194) );
  NAND2_X1 U9268 ( .A1(n11152), .A2(n7021), .ZN(n11556) );
  NAND2_X1 U9269 ( .A1(n11556), .A2(n11468), .ZN(n7834) );
  NAND2_X1 U9270 ( .A1(n7736), .A2(n7735), .ZN(n10875) );
  OAI21_X1 U9271 ( .B1(n9430), .B2(n9429), .A(n9428), .ZN(n9432) );
  NAND2_X1 U9272 ( .A1(n9338), .A2(n9337), .ZN(n9341) );
  NAND2_X1 U9273 ( .A1(n9410), .A2(n9409), .ZN(n9414) );
  NAND2_X1 U9274 ( .A1(n9375), .A2(n9374), .ZN(n9377) );
  NAND2_X1 U9275 ( .A1(n9315), .A2(n9314), .ZN(n9318) );
  NAND2_X1 U9276 ( .A1(n9387), .A2(n9386), .ZN(n9389) );
  NAND2_X1 U9277 ( .A1(n7537), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7550) );
  NAND2_X1 U9278 ( .A1(n9062), .A2(n6599), .ZN(n7022) );
  NAND2_X1 U9279 ( .A1(n9060), .A2(n9059), .ZN(n9062) );
  NAND2_X1 U9280 ( .A1(n8753), .A2(n7022), .ZN(n9072) );
  NAND2_X1 U9281 ( .A1(n9031), .A2(n7030), .ZN(n7026) );
  NAND2_X1 U9282 ( .A1(n7026), .A2(n7027), .ZN(n8783) );
  NAND2_X1 U9283 ( .A1(n9270), .A2(n7037), .ZN(n7033) );
  NAND2_X1 U9284 ( .A1(n7033), .A2(n7034), .ZN(n12078) );
  OAI21_X1 U9285 ( .B1(n9128), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n9129), .ZN(
        n9139) );
  OAI21_X1 U9286 ( .B1(n8885), .B2(n8719), .A(n8720), .ZN(n8895) );
  NAND2_X1 U9287 ( .A1(n8719), .A2(n8720), .ZN(n7055) );
  NAND2_X1 U9288 ( .A1(n8958), .A2(n6586), .ZN(n7058) );
  NAND2_X1 U9289 ( .A1(n7064), .A2(n7063), .ZN(n7982) );
  NAND2_X1 U9290 ( .A1(n7980), .A2(n7065), .ZN(n7063) );
  AOI21_X1 U9291 ( .B1(n11025), .B2(n7066), .A(n6540), .ZN(n7065) );
  OAI21_X1 U9292 ( .B1(n11206), .B2(n7072), .A(n7070), .ZN(n11148) );
  NAND2_X1 U9293 ( .A1(n7069), .A2(n7068), .ZN(n7986) );
  AOI21_X1 U9294 ( .B1(n7070), .B2(n7072), .A(n6543), .ZN(n7068) );
  NAND2_X1 U9295 ( .A1(n11206), .A2(n7070), .ZN(n7069) );
  OAI21_X1 U9296 ( .B1(n11243), .B2(n7075), .A(n7073), .ZN(n11208) );
  AOI21_X2 U9297 ( .B1(n7994), .B2(n6520), .A(n7082), .ZN(n13114) );
  NAND2_X1 U9298 ( .A1(n13061), .A2(n6576), .ZN(n7086) );
  NAND2_X1 U9299 ( .A1(n7104), .A2(n7103), .ZN(n10764) );
  INV_X1 U9300 ( .A(n7108), .ZN(n10647) );
  NAND2_X1 U9301 ( .A1(n7110), .A2(n7112), .ZN(n14901) );
  OAI21_X1 U9302 ( .B1(n12350), .B2(n12349), .A(n14899), .ZN(n7112) );
  NAND2_X1 U9303 ( .A1(n6466), .A2(n12398), .ZN(n7122) );
  INV_X1 U9304 ( .A(n7124), .ZN(n12422) );
  OAI211_X1 U9305 ( .C1(n13558), .C2(n6584), .A(n7132), .B(n7130), .ZN(n13473)
         );
  OAI22_X1 U9306 ( .A1(n7134), .A2(n7131), .B1(n13468), .B2(n7136), .ZN(n7130)
         );
  NOR2_X1 U9307 ( .A1(n13423), .A2(n13468), .ZN(n7131) );
  NAND2_X1 U9308 ( .A1(n13558), .A2(n7133), .ZN(n7132) );
  NOR2_X1 U9309 ( .A1(n7134), .A2(n13468), .ZN(n7133) );
  INV_X1 U9310 ( .A(n13468), .ZN(n7135) );
  NAND2_X1 U9311 ( .A1(n13541), .A2(n7141), .ZN(n7140) );
  NAND2_X1 U9312 ( .A1(n13505), .A2(n7156), .ZN(n7152) );
  NOR2_X1 U9313 ( .A1(n6512), .A2(n7368), .ZN(n13517) );
  NAND2_X1 U9314 ( .A1(n10577), .A2(n6476), .ZN(n10617) );
  NAND2_X1 U9315 ( .A1(n10228), .A2(n10229), .ZN(n10577) );
  NAND2_X1 U9316 ( .A1(n8064), .A2(n6482), .ZN(n8366) );
  INV_X1 U9317 ( .A(n11836), .ZN(n7173) );
  NAND2_X1 U9318 ( .A1(n12769), .A2(n7181), .ZN(n7178) );
  OAI211_X1 U9319 ( .C1(n12769), .C2(n7183), .A(n7178), .B(n7179), .ZN(
        P2_U3192) );
  NAND3_X1 U9320 ( .A1(n7191), .A2(n7192), .A3(n7196), .ZN(n11084) );
  AOI21_X1 U9321 ( .B1(n7194), .B2(n7193), .A(n6518), .ZN(n7192) );
  OAI21_X1 U9322 ( .B1(n10678), .B2(n10677), .A(n9615), .ZN(n10567) );
  NAND2_X1 U9323 ( .A1(n11832), .A2(n7200), .ZN(n12785) );
  NAND2_X2 U9324 ( .A1(n9658), .A2(n11825), .ZN(n11832) );
  OAI211_X1 U9325 ( .C1(n7411), .C2(n9744), .A(n7204), .B(n7203), .ZN(n7416)
         );
  NAND3_X1 U9326 ( .A1(n7411), .A2(n7412), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n7203) );
  INV_X1 U9327 ( .A(n7412), .ZN(n7205) );
  MUX2_X1 U9328 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n7433), .Z(n7419) );
  MUX2_X1 U9329 ( .A(n8712), .B(n9755), .S(n7433), .Z(n7422) );
  MUX2_X1 U9330 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n7433), .Z(n7426) );
  MUX2_X1 U9331 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7433), .Z(n7429) );
  MUX2_X1 U9332 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7433), .Z(n7432) );
  NAND2_X1 U9333 ( .A1(n7564), .A2(n7428), .ZN(n7212) );
  NAND2_X1 U9334 ( .A1(n7598), .A2(n7440), .ZN(n7218) );
  NAND2_X1 U9335 ( .A1(n11652), .A2(n7229), .ZN(n7226) );
  NAND2_X1 U9336 ( .A1(n12496), .A2(n9150), .ZN(n7240) );
  OAI21_X1 U9337 ( .B1(n12496), .B2(n7238), .A(n7235), .ZN(n9269) );
  NAND2_X1 U9338 ( .A1(n7234), .A2(n7233), .ZN(n9274) );
  NAND2_X1 U9339 ( .A1(n12496), .A2(n7235), .ZN(n7234) );
  NAND2_X1 U9340 ( .A1(n7241), .A2(n7242), .ZN(n12550) );
  NAND2_X1 U9341 ( .A1(n12595), .A2(n7245), .ZN(n7241) );
  INV_X1 U9342 ( .A(n7256), .ZN(n12509) );
  INV_X1 U9343 ( .A(n7263), .ZN(n7260) );
  OAI21_X2 U9344 ( .B1(n10790), .B2(n7266), .A(n7267), .ZN(n11013) );
  NAND2_X1 U9345 ( .A1(n8695), .A2(n7269), .ZN(n7271) );
  NAND2_X1 U9346 ( .A1(n7377), .A2(n8851), .ZN(n7273) );
  NOR2_X2 U9347 ( .A1(n7273), .A2(n7271), .ZN(n8760) );
  NAND3_X1 U9348 ( .A1(n7377), .A2(n8851), .A3(n8695), .ZN(n9032) );
  NAND2_X1 U9349 ( .A1(n9206), .A2(n7275), .ZN(n8771) );
  NAND3_X1 U9350 ( .A1(n8831), .A2(n8830), .A3(n7278), .ZN(n10482) );
  NAND2_X1 U9351 ( .A1(n11056), .A2(n7279), .ZN(n11413) );
  NAND2_X1 U9352 ( .A1(n11413), .A2(n12135), .ZN(n8947) );
  XNOR2_X1 U9353 ( .A(n10291), .B(n10317), .ZN(n10276) );
  NAND2_X1 U9354 ( .A1(n14279), .A2(n7301), .ZN(n7298) );
  NAND2_X1 U9355 ( .A1(n14288), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7301) );
  NAND2_X1 U9356 ( .A1(n7307), .A2(n7306), .ZN(n8344) );
  NAND3_X1 U9357 ( .A1(n8294), .A2(n8293), .A3(n6504), .ZN(n7307) );
  INV_X1 U9358 ( .A(n8310), .ZN(n7310) );
  NAND2_X1 U9359 ( .A1(n8134), .A2(n10704), .ZN(n7314) );
  NAND2_X1 U9360 ( .A1(n7315), .A2(n7316), .ZN(n8402) );
  NAND2_X1 U9361 ( .A1(n8346), .A2(n6583), .ZN(n7315) );
  OAI21_X1 U9362 ( .B1(n8345), .B2(n7319), .A(n8362), .ZN(n7318) );
  INV_X1 U9363 ( .A(n8363), .ZN(n7319) );
  NAND2_X1 U9364 ( .A1(n7323), .A2(n7321), .ZN(n8254) );
  NAND2_X1 U9365 ( .A1(n7326), .A2(n7327), .ZN(n8615) );
  NAND3_X1 U9366 ( .A1(n8541), .A2(n6582), .A3(n8540), .ZN(n7326) );
  NAND2_X1 U9367 ( .A1(n7331), .A2(n6579), .ZN(n8289) );
  NAND3_X1 U9368 ( .A1(n8257), .A2(n6580), .A3(n8256), .ZN(n7331) );
  NAND2_X1 U9369 ( .A1(n7333), .A2(n7334), .ZN(n8470) );
  NAND3_X1 U9370 ( .A1(n8446), .A2(n6573), .A3(n8445), .ZN(n7333) );
  NAND2_X1 U9371 ( .A1(n7336), .A2(n7337), .ZN(n8503) );
  NAND3_X1 U9372 ( .A1(n8475), .A2(n6574), .A3(n8474), .ZN(n7336) );
  NAND3_X1 U9373 ( .A1(n8508), .A2(n6575), .A3(n8507), .ZN(n7339) );
  NAND2_X1 U9374 ( .A1(n7339), .A2(n7340), .ZN(n8536) );
  NAND2_X1 U9375 ( .A1(n7342), .A2(n7343), .ZN(n8207) );
  NAND3_X1 U9376 ( .A1(n8170), .A2(n8171), .A3(n6570), .ZN(n7342) );
  NAND2_X1 U9377 ( .A1(n8094), .A2(n7345), .ZN(n8669) );
  NAND2_X1 U9378 ( .A1(n11867), .A2(n11866), .ZN(n13750) );
  OAI21_X2 U9379 ( .B1(n11867), .B2(n7350), .A(n7348), .ZN(n13769) );
  OAI22_X1 U9380 ( .A1(n13769), .A2(n13752), .B1(n13751), .B2(n13980), .ZN(
        n13753) );
  NAND2_X1 U9381 ( .A1(n14494), .A2(n11538), .ZN(n7351) );
  NAND2_X2 U9382 ( .A1(n13822), .A2(n13821), .ZN(n13820) );
  NAND2_X2 U9383 ( .A1(n11765), .A2(n11764), .ZN(n11786) );
  OAI22_X1 U9384 ( .A1(n8462), .A2(n9931), .B1(n8492), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n8120) );
  NAND2_X2 U9385 ( .A1(n13925), .A2(n7362), .ZN(n13905) );
  NAND3_X1 U9386 ( .A1(n8064), .A2(n7380), .A3(n8048), .ZN(n8676) );
  OAI21_X1 U9387 ( .B1(n12499), .B2(n14939), .A(n12498), .ZN(n12679) );
  INV_X1 U9388 ( .A(n7723), .ZN(n13305) );
  NAND2_X1 U9389 ( .A1(n8817), .A2(n12332), .ZN(n12145) );
  NAND2_X1 U9390 ( .A1(n12973), .A2(n13169), .ZN(n12980) );
  AND2_X2 U9391 ( .A1(n10578), .A2(n10041), .ZN(n10598) );
  INV_X1 U9392 ( .A(n7400), .ZN(n7397) );
  NAND2_X2 U9393 ( .A1(n9702), .A2(n12808), .ZN(n12811) );
  OAI21_X2 U9394 ( .B1(n9197), .B2(n9196), .A(n9195), .ZN(n12673) );
  OAI211_X1 U9395 ( .C1(n8402), .C2(n11873), .A(n8403), .B(n13926), .ZN(n8412)
         );
  INV_X1 U9396 ( .A(n10499), .ZN(n8845) );
  OR2_X1 U9397 ( .A1(n10094), .A2(n8968), .ZN(n8790) );
  XNOR2_X1 U9398 ( .A(n9588), .B(n14785), .ZN(n9593) );
  OR2_X1 U9399 ( .A1(n8775), .A2(n8973), .ZN(n8776) );
  NAND4_X1 U9400 ( .A1(n8113), .A2(n8112), .A3(n8111), .A4(n8110), .ZN(n13599)
         );
  INV_X1 U9401 ( .A(n10704), .ZN(n10696) );
  AND2_X1 U9402 ( .A1(n8123), .A2(n8122), .ZN(n7371) );
  AND2_X1 U9403 ( .A1(n12404), .A2(n12403), .ZN(n12405) );
  OR2_X1 U9404 ( .A1(n6461), .A2(n8055), .ZN(n8063) );
  INV_X1 U9405 ( .A(n11149), .ZN(n7815) );
  NOR2_X2 U9406 ( .A1(n8366), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n8094) );
  NAND2_X1 U9407 ( .A1(n8624), .A2(n10945), .ZN(n10041) );
  AND2_X1 U9408 ( .A1(n13346), .A2(n13345), .ZN(n7368) );
  OR2_X1 U9409 ( .A1(n8829), .A2(n6614), .ZN(n7369) );
  INV_X1 U9410 ( .A(n11860), .ZN(n13837) );
  INV_X1 U9411 ( .A(n12387), .ZN(n14916) );
  AND2_X1 U9412 ( .A1(n8993), .A2(n9020), .ZN(n12387) );
  INV_X1 U9413 ( .A(n11708), .ZN(n7843) );
  OR2_X1 U9414 ( .A1(n7417), .A2(n9758), .ZN(n7370) );
  AND2_X1 U9415 ( .A1(n6531), .A2(n9299), .ZN(n7372) );
  NOR2_X1 U9416 ( .A1(n9505), .A2(n9504), .ZN(n7373) );
  AND2_X1 U9417 ( .A1(n9525), .A2(n9519), .ZN(n7374) );
  AND3_X1 U9418 ( .A1(n8667), .A2(n8666), .A3(n8665), .ZN(n7375) );
  AND2_X1 U9419 ( .A1(n7452), .A2(n7451), .ZN(n7376) );
  AND2_X1 U9420 ( .A1(n11629), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7378) );
  INV_X1 U9421 ( .A(n11180), .ZN(n11526) );
  AND2_X1 U9422 ( .A1(n8278), .A2(n8277), .ZN(n7379) );
  INV_X1 U9423 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n8773) );
  AND2_X1 U9424 ( .A1(n13463), .A2(n14534), .ZN(n14588) );
  INV_X1 U9425 ( .A(n8819), .ZN(n8832) );
  AND2_X1 U9426 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7381) );
  INV_X1 U9427 ( .A(n15034), .ZN(n15039) );
  AND2_X1 U9428 ( .A1(n13454), .A2(n13452), .ZN(n7384) );
  INV_X1 U9429 ( .A(n8403), .ZN(n13909) );
  AND2_X1 U9430 ( .A1(n9520), .A2(n12997), .ZN(n7385) );
  INV_X1 U9431 ( .A(n14798), .ZN(n8001) );
  INV_X1 U9432 ( .A(n14852), .ZN(n14841) );
  INV_X1 U9433 ( .A(n11718), .ZN(n7852) );
  INV_X1 U9434 ( .A(n13515), .ZN(n13348) );
  AND2_X1 U9435 ( .A1(n8996), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n7386) );
  AND2_X1 U9436 ( .A1(n12108), .A2(n9185), .ZN(n7387) );
  OR2_X1 U9437 ( .A1(n9530), .A2(n9303), .ZN(n9306) );
  NAND2_X1 U9438 ( .A1(n9304), .A2(n10881), .ZN(n9316) );
  OAI21_X1 U9439 ( .B1(n9304), .B2(n10424), .A(n9316), .ZN(n9319) );
  MUX2_X1 U9440 ( .A(n10706), .B(n8135), .S(n8252), .Z(n8136) );
  INV_X1 U9441 ( .A(n8203), .ZN(n8204) );
  INV_X1 U9442 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8693) );
  INV_X1 U9443 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7393) );
  INV_X1 U9444 ( .A(n10280), .ZN(n10281) );
  AND4_X1 U9445 ( .A1(n8758), .A2(n8757), .A3(n8756), .A4(n8755), .ZN(n8759)
         );
  INV_X1 U9446 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7392) );
  OR2_X1 U9447 ( .A1(n14556), .A2(n10594), .ZN(n10215) );
  AND2_X1 U9448 ( .A1(n10762), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n10763) );
  AND2_X1 U9449 ( .A1(n12383), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12384) );
  INV_X1 U9450 ( .A(n14954), .ZN(n8817) );
  OR2_X1 U9451 ( .A1(n7518), .A2(n13296), .ZN(n7515) );
  INV_X1 U9452 ( .A(n7606), .ZN(n7443) );
  OR2_X1 U9453 ( .A1(n8949), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8977) );
  INV_X1 U9454 ( .A(n12182), .ZN(n8933) );
  NAND2_X1 U9455 ( .A1(n8942), .A2(n8727), .ZN(n8729) );
  INV_X1 U9456 ( .A(n12803), .ZN(n9676) );
  OR2_X1 U9457 ( .A1(n7905), .A2(n12845), .ZN(n7913) );
  INV_X1 U9458 ( .A(n12970), .ZN(n12971) );
  INV_X1 U9459 ( .A(n7883), .ZN(n7881) );
  INV_X1 U9460 ( .A(n8430), .ZN(n8429) );
  OR2_X1 U9461 ( .A1(n8523), .A2(n8522), .ZN(n8544) );
  INV_X1 U9462 ( .A(n8417), .ZN(n8414) );
  INV_X1 U9463 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8214) );
  INV_X1 U9464 ( .A(n7526), .ZN(n7638) );
  AND2_X1 U9465 ( .A1(n11938), .A2(n11937), .ZN(n11939) );
  INV_X1 U9466 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8861) );
  OR2_X1 U9467 ( .A1(n8977), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8996) );
  NOR2_X1 U9468 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(n9144), .ZN(n9158) );
  OR2_X1 U9469 ( .A1(n12691), .A2(n12311), .ZN(n9127) );
  OR2_X1 U9470 ( .A1(n12273), .A2(n12290), .ZN(n10389) );
  NAND2_X1 U9471 ( .A1(n8703), .A2(n8755), .ZN(n8701) );
  NAND2_X1 U9472 ( .A1(n9019), .A2(n8740), .ZN(n8742) );
  NAND2_X1 U9473 ( .A1(n8712), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8713) );
  AND2_X1 U9474 ( .A1(n9703), .A2(n9701), .ZN(n12808) );
  INV_X1 U9475 ( .A(n12859), .ZN(n9667) );
  INV_X1 U9476 ( .A(n7804), .ZN(n7803) );
  AND2_X1 U9477 ( .A1(n9509), .A2(n9508), .ZN(n9510) );
  NAND2_X1 U9478 ( .A1(n7895), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n7905) );
  OAI22_X1 U9479 ( .A1(n12977), .A2(n13069), .B1(n13067), .B2(n12814), .ZN(
        n7972) );
  NAND2_X1 U9480 ( .A1(n7881), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n7890) );
  INV_X1 U9481 ( .A(n10814), .ZN(n10821) );
  OAI211_X1 U9482 ( .C1(n9754), .C2(n7543), .A(n6517), .B(n7555), .ZN(n14785)
         );
  INV_X1 U9483 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7402) );
  INV_X1 U9484 ( .A(n14328), .ZN(n13332) );
  AND2_X1 U9485 ( .A1(n13363), .A2(n13362), .ZN(n13364) );
  INV_X1 U9486 ( .A(n11296), .ZN(n11292) );
  INV_X1 U9487 ( .A(n11619), .ZN(n11615) );
  OR2_X1 U9488 ( .A1(n8478), .A2(n8476), .ZN(n8490) );
  NAND2_X1 U9489 ( .A1(n8429), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8447) );
  AND2_X1 U9490 ( .A1(n8544), .A2(n8524), .ZN(n13425) );
  OR2_X1 U9491 ( .A1(n8447), .A2(n13543), .ZN(n8478) );
  NAND2_X1 U9492 ( .A1(n8414), .A2(n8413), .ZN(n8430) );
  OR2_X1 U9493 ( .A1(n8259), .A2(n8258), .ZN(n8278) );
  NAND2_X1 U9494 ( .A1(n7445), .A2(n8956), .ZN(n7448) );
  NOR2_X1 U9495 ( .A1(n14173), .A2(n14172), .ZN(n14113) );
  NOR2_X1 U9496 ( .A1(n8888), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8918) );
  AND2_X1 U9497 ( .A1(n9011), .A2(n9010), .ZN(n9024) );
  INV_X1 U9498 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n8934) );
  NAND2_X1 U9499 ( .A1(n12334), .A2(n10252), .ZN(n14947) );
  NAND2_X1 U9500 ( .A1(n11961), .A2(n12046), .ZN(n12029) );
  INV_X1 U9501 ( .A(n12055), .ZN(n12300) );
  OR2_X1 U9502 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(n9121), .ZN(n9133) );
  NAND2_X1 U9503 ( .A1(n9076), .A2(n9075), .ZN(n9078) );
  NAND2_X1 U9504 ( .A1(n9037), .A2(n9036), .ZN(n9051) );
  INV_X1 U9505 ( .A(n11983), .ZN(n9195) );
  OR2_X1 U9506 ( .A1(n12302), .A2(n10145), .ZN(n15001) );
  OR2_X1 U9507 ( .A1(n12751), .A2(n9743), .ZN(n10177) );
  NAND2_X1 U9508 ( .A1(n7775), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7794) );
  BUF_X4 U9509 ( .A(n9588), .Z(n9716) );
  OR2_X1 U9510 ( .A1(n7890), .A2(n12827), .ZN(n7897) );
  NAND2_X1 U9511 ( .A1(n7803), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7820) );
  INV_X1 U9512 ( .A(n12841), .ZN(n12872) );
  OR2_X1 U9513 ( .A1(n12996), .A2(n6441), .ZN(n7970) );
  OR2_X1 U9514 ( .A1(n7873), .A2(n7872), .ZN(n7883) );
  OR2_X1 U9515 ( .A1(n10023), .A2(n10024), .ZN(n10104) );
  OR2_X1 U9516 ( .A1(n10100), .A2(n10101), .ZN(n12930) );
  OAI21_X1 U9517 ( .B1(n11716), .B2(n7852), .A(n7990), .ZN(n11738) );
  INV_X1 U9518 ( .A(n13152), .ZN(n13067) );
  NAND2_X1 U9519 ( .A1(n13135), .A2(n10824), .ZN(n13178) );
  AND2_X1 U9520 ( .A1(n13524), .A2(n13391), .ZN(n13432) );
  INV_X1 U9521 ( .A(n13819), .ZN(n13565) );
  OR2_X1 U9522 ( .A1(n8397), .A2(n8396), .ZN(n8417) );
  INV_X1 U9523 ( .A(n13511), .ZN(n14355) );
  NAND2_X1 U9524 ( .A1(n8617), .A2(n8616), .ZN(n8620) );
  XNOR2_X1 U9525 ( .A(n8598), .B(n8597), .ZN(n9470) );
  AND2_X1 U9526 ( .A1(n7456), .A2(n7455), .ZN(n7631) );
  OAI21_X1 U9527 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n14112), .A(n14111), .ZN(
        n14172) );
  NAND2_X1 U9528 ( .A1(n8935), .A2(n8934), .ZN(n8949) );
  INV_X1 U9529 ( .A(n14893), .ZN(n12073) );
  AND4_X1 U9530 ( .A1(n9182), .A2(n9181), .A3(n9180), .A4(n9179), .ZN(n11956)
         );
  INV_X1 U9531 ( .A(n14939), .ZN(n14948) );
  INV_X1 U9532 ( .A(n11656), .ZN(n14959) );
  INV_X1 U9533 ( .A(n12655), .ZN(n12661) );
  AND2_X1 U9534 ( .A1(n6619), .A2(n12469), .ZN(n12666) );
  INV_X1 U9535 ( .A(n10177), .ZN(n12298) );
  NAND2_X1 U9536 ( .A1(n8783), .A2(n8782), .ZN(n8785) );
  AND2_X1 U9537 ( .A1(n8929), .A2(n8972), .ZN(n10957) );
  XNOR2_X1 U9538 ( .A(n8840), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10317) );
  INV_X1 U9539 ( .A(n9721), .ZN(n9722) );
  AND2_X1 U9540 ( .A1(n7932), .A2(n7922), .ZN(n13055) );
  INV_X1 U9541 ( .A(n11346), .ZN(n9521) );
  AND3_X1 U9542 ( .A1(n7894), .A2(n7893), .A3(n7892), .ZN(n12797) );
  OR2_X1 U9543 ( .A1(n6439), .A2(n7722), .ZN(n7728) );
  AND2_X1 U9544 ( .A1(n9887), .A2(n9874), .ZN(n14724) );
  AND2_X1 U9545 ( .A1(n9887), .A2(n9867), .ZN(n14728) );
  INV_X1 U9546 ( .A(n13140), .ZN(n13185) );
  NAND2_X2 U9547 ( .A1(n10816), .A2(n13133), .ZN(n13135) );
  INV_X1 U9548 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8037) );
  AND2_X1 U9549 ( .A1(n14839), .A2(n14838), .ZN(n14798) );
  AND2_X1 U9550 ( .A1(n8015), .A2(n8034), .ZN(n14733) );
  OR2_X1 U9551 ( .A1(n8319), .A2(n8318), .ZN(n8334) );
  INV_X1 U9552 ( .A(n14556), .ZN(n13479) );
  OAI21_X1 U9553 ( .B1(n10853), .B2(n10852), .A(n10851), .ZN(n10859) );
  OR2_X1 U9554 ( .A1(n13469), .A2(n8589), .ZN(n8551) );
  AND3_X1 U9555 ( .A1(n8421), .A2(n8420), .A3(n8419), .ZN(n13488) );
  AND4_X1 U9556 ( .A1(n8339), .A2(n8338), .A3(n8337), .A4(n8336), .ZN(n14324)
         );
  INV_X1 U9557 ( .A(n14478), .ZN(n14440) );
  INV_X1 U9558 ( .A(n14482), .ZN(n14442) );
  INV_X1 U9559 ( .A(n14526), .ZN(n14508) );
  OR2_X1 U9560 ( .A1(n10540), .A2(n10068), .ZN(n13952) );
  INV_X1 U9561 ( .A(n14584), .ZN(n14574) );
  AND2_X1 U9562 ( .A1(n10541), .A2(n10417), .ZN(n11075) );
  INV_X1 U9563 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8326) );
  AND2_X1 U9564 ( .A1(n10129), .A2(n10128), .ZN(n14931) );
  INV_X1 U9565 ( .A(n12557), .ZN(n12708) );
  AND4_X1 U9566 ( .A1(n12095), .A2(n9189), .A3(n9188), .A4(n9187), .ZN(n10787)
         );
  INV_X1 U9567 ( .A(n11964), .ZN(n12313) );
  OR2_X1 U9568 ( .A1(n9295), .A2(n9294), .ZN(n12489) );
  OR2_X1 U9569 ( .A1(n14965), .A2(n9291), .ZN(n14944) );
  AND2_X2 U9570 ( .A1(n9568), .A2(n12298), .ZN(n15025) );
  CLKBUF_X1 U9571 ( .A(n9807), .Z(n9830) );
  INV_X1 U9572 ( .A(SI_13_), .ZN(n15157) );
  INV_X1 U9573 ( .A(n12351), .ZN(n14899) );
  OR2_X1 U9574 ( .A1(n12828), .A2(n13069), .ZN(n12869) );
  INV_X1 U9575 ( .A(n12871), .ZN(n12829) );
  INV_X1 U9576 ( .A(n9735), .ZN(n12989) );
  INV_X1 U9577 ( .A(n9697), .ZN(n13017) );
  INV_X1 U9578 ( .A(n14657), .ZN(n14716) );
  OR2_X1 U9579 ( .A1(n9887), .A2(P2_U3088), .ZN(n14731) );
  AND2_X1 U9580 ( .A1(n13163), .A2(n10813), .ZN(n13182) );
  INV_X1 U9581 ( .A(n14876), .ZN(n14873) );
  OR2_X1 U9582 ( .A1(n14858), .A2(n8037), .ZN(n8038) );
  OR2_X1 U9583 ( .A1(n13267), .A2(n13266), .ZN(n13292) );
  INV_X1 U9584 ( .A(n14858), .ZN(n14856) );
  INV_X1 U9585 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10363) );
  AND2_X1 U9586 ( .A1(n10610), .A2(n11344), .ZN(n14339) );
  INV_X1 U9587 ( .A(n14335), .ZN(n13580) );
  NAND2_X1 U9588 ( .A1(n8551), .A2(n8550), .ZN(n13759) );
  INV_X1 U9589 ( .A(n13488), .ZN(n13913) );
  INV_X1 U9590 ( .A(n10709), .ZN(n13597) );
  OR2_X1 U9591 ( .A1(n9956), .A2(n9942), .ZN(n14482) );
  INV_X1 U9592 ( .A(n14501), .ZN(n13958) );
  INV_X1 U9593 ( .A(n14511), .ZN(n13899) );
  INV_X1 U9594 ( .A(n14597), .ZN(n14595) );
  AND2_X1 U9595 ( .A1(n9832), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9800) );
  INV_X1 U9596 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10468) );
  INV_X1 U9597 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9927) );
  NAND2_X1 U9598 ( .A1(n9268), .A2(n9267), .ZN(P3_U3487) );
  NAND2_X1 U9599 ( .A1(n8039), .A2(n8038), .ZN(P2_U3494) );
  NAND2_X1 U9600 ( .A1(n7394), .A2(n7393), .ZN(n7663) );
  NAND2_X1 U9601 ( .A1(n7406), .A2(n7509), .ZN(n7400) );
  INV_X1 U9602 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n7398) );
  XNOR2_X2 U9603 ( .A(n7399), .B(n7398), .ZN(n9576) );
  NAND2_X1 U9604 ( .A1(n7400), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7401) );
  NAND2_X1 U9605 ( .A1(n7401), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n7404) );
  NAND2_X1 U9606 ( .A1(n7408), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7409) );
  NAND2_X1 U9607 ( .A1(n10893), .A2(n11725), .ZN(n9522) );
  NAND2_X1 U9608 ( .A1(n14772), .A2(n9522), .ZN(n14852) );
  XNOR2_X1 U9609 ( .A(n7416), .B(SI_1_), .ZN(n7536) );
  INV_X1 U9610 ( .A(n7536), .ZN(n7415) );
  AND2_X1 U9611 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n7413) );
  AND2_X1 U9612 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7414) );
  INV_X1 U9613 ( .A(n7416), .ZN(n7417) );
  INV_X1 U9614 ( .A(SI_1_), .ZN(n9758) );
  XNOR2_X2 U9615 ( .A(n7419), .B(SI_2_), .ZN(n7545) );
  INV_X1 U9616 ( .A(n7545), .ZN(n7418) );
  NAND2_X1 U9617 ( .A1(n7544), .A2(n7418), .ZN(n7421) );
  NAND2_X1 U9618 ( .A1(n7419), .A2(SI_2_), .ZN(n7420) );
  INV_X1 U9619 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9755) );
  INV_X1 U9620 ( .A(n7422), .ZN(n7423) );
  NAND2_X1 U9621 ( .A1(n7423), .A2(SI_3_), .ZN(n7424) );
  NAND2_X1 U9622 ( .A1(n7426), .A2(SI_4_), .ZN(n7427) );
  NAND2_X1 U9623 ( .A1(n7429), .A2(SI_5_), .ZN(n7430) );
  MUX2_X1 U9624 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6459), .Z(n7435) );
  NAND2_X1 U9625 ( .A1(n7435), .A2(SI_7_), .ZN(n7436) );
  MUX2_X1 U9626 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6459), .Z(n7438) );
  NAND2_X1 U9627 ( .A1(n7438), .A2(SI_8_), .ZN(n7439) );
  MUX2_X1 U9628 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n6459), .Z(n7441) );
  NAND2_X1 U9629 ( .A1(n7441), .A2(SI_9_), .ZN(n7442) );
  MUX2_X1 U9630 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n6459), .Z(n7444) );
  MUX2_X1 U9631 ( .A(n9858), .B(n9861), .S(n6459), .Z(n7445) );
  INV_X1 U9632 ( .A(SI_11_), .ZN(n8956) );
  INV_X1 U9633 ( .A(n7445), .ZN(n7446) );
  NAND2_X1 U9634 ( .A1(n7446), .A2(SI_11_), .ZN(n7447) );
  MUX2_X1 U9635 ( .A(n9927), .B(n9926), .S(n6459), .Z(n7449) );
  NAND2_X1 U9636 ( .A1(n7449), .A2(n15162), .ZN(n7452) );
  INV_X1 U9637 ( .A(n7449), .ZN(n7450) );
  NAND2_X1 U9638 ( .A1(n7450), .A2(SI_12_), .ZN(n7451) );
  MUX2_X1 U9639 ( .A(n10076), .B(n10078), .S(n6459), .Z(n7453) );
  INV_X1 U9640 ( .A(n7453), .ZN(n7454) );
  NAND2_X1 U9641 ( .A1(n7454), .A2(SI_13_), .ZN(n7455) );
  MUX2_X1 U9642 ( .A(n10367), .B(n10369), .S(n6458), .Z(n7526) );
  NAND2_X1 U9643 ( .A1(n7638), .A2(SI_14_), .ZN(n7457) );
  MUX2_X1 U9644 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n6459), .Z(n7458) );
  NOR2_X1 U9645 ( .A1(n7638), .A2(SI_14_), .ZN(n7462) );
  INV_X1 U9646 ( .A(n7458), .ZN(n7460) );
  INV_X1 U9647 ( .A(SI_15_), .ZN(n7459) );
  NAND2_X1 U9648 ( .A1(n7460), .A2(n7459), .ZN(n7644) );
  INV_X1 U9649 ( .A(n7644), .ZN(n7461) );
  AOI21_X1 U9650 ( .B1(n7462), .B2(n7645), .A(n7461), .ZN(n7463) );
  MUX2_X1 U9651 ( .A(n10365), .B(n10363), .S(n6459), .Z(n7466) );
  INV_X1 U9652 ( .A(SI_16_), .ZN(n7465) );
  NAND2_X1 U9653 ( .A1(n7466), .A2(n7465), .ZN(n7469) );
  INV_X1 U9654 ( .A(n7466), .ZN(n7467) );
  NAND2_X1 U9655 ( .A1(n7467), .A2(SI_16_), .ZN(n7468) );
  NAND2_X1 U9656 ( .A1(n7654), .A2(n7653), .ZN(n7470) );
  MUX2_X1 U9657 ( .A(n10468), .B(n10471), .S(n6459), .Z(n7471) );
  INV_X1 U9658 ( .A(SI_17_), .ZN(n10031) );
  INV_X1 U9659 ( .A(n7471), .ZN(n7472) );
  NAND2_X1 U9660 ( .A1(n7472), .A2(SI_17_), .ZN(n7473) );
  MUX2_X1 U9661 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n6459), .Z(n7674) );
  NAND2_X1 U9662 ( .A1(n7674), .A2(SI_18_), .ZN(n7476) );
  MUX2_X1 U9663 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n6459), .Z(n7478) );
  NAND2_X1 U9664 ( .A1(n7478), .A2(SI_19_), .ZN(n7681) );
  NOR2_X1 U9665 ( .A1(n7674), .A2(SI_18_), .ZN(n7481) );
  INV_X1 U9666 ( .A(n7478), .ZN(n7479) );
  INV_X1 U9667 ( .A(SI_19_), .ZN(n10113) );
  NAND2_X1 U9668 ( .A1(n7479), .A2(n10113), .ZN(n7680) );
  INV_X1 U9669 ( .A(n7680), .ZN(n7480) );
  AOI21_X1 U9670 ( .B1(n7481), .B2(n7681), .A(n7480), .ZN(n7482) );
  INV_X1 U9671 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10868) );
  INV_X1 U9672 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10894) );
  MUX2_X1 U9673 ( .A(n10868), .B(n10894), .S(n6459), .Z(n7689) );
  INV_X1 U9674 ( .A(n7689), .ZN(n7483) );
  INV_X1 U9675 ( .A(SI_20_), .ZN(n10535) );
  MUX2_X1 U9676 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6458), .Z(n7488) );
  XNOR2_X1 U9677 ( .A(n7488), .B(SI_21_), .ZN(n7692) );
  NAND2_X1 U9678 ( .A1(n7488), .A2(SI_21_), .ZN(n7489) );
  MUX2_X1 U9679 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n6458), .Z(n7696) );
  INV_X1 U9680 ( .A(SI_22_), .ZN(n9088) );
  MUX2_X1 U9681 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n6459), .Z(n7700) );
  INV_X1 U9682 ( .A(n7700), .ZN(n7491) );
  INV_X1 U9683 ( .A(SI_23_), .ZN(n10943) );
  AOI22_X1 U9684 ( .A1(n7523), .A2(n9088), .B1(n7491), .B2(n10943), .ZN(n7492)
         );
  OAI21_X1 U9685 ( .B1(n7523), .B2(n9088), .A(n10943), .ZN(n7494) );
  AND2_X1 U9686 ( .A1(SI_22_), .A2(SI_23_), .ZN(n7493) );
  AOI22_X1 U9687 ( .A1(n7494), .A2(n7700), .B1(n7696), .B2(n7493), .ZN(n7495)
         );
  MUX2_X1 U9688 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n6458), .Z(n7705) );
  NAND2_X1 U9689 ( .A1(n7496), .A2(SI_24_), .ZN(n7497) );
  INV_X1 U9690 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11502) );
  INV_X1 U9691 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11505) );
  MUX2_X1 U9692 ( .A(n11502), .B(n11505), .S(n6459), .Z(n7499) );
  INV_X1 U9693 ( .A(SI_25_), .ZN(n11498) );
  NAND2_X1 U9694 ( .A1(n7499), .A2(n11498), .ZN(n7502) );
  INV_X1 U9695 ( .A(n7499), .ZN(n7500) );
  NAND2_X1 U9696 ( .A1(n7500), .A2(SI_25_), .ZN(n7501) );
  NAND2_X1 U9697 ( .A1(n7502), .A2(n7501), .ZN(n7709) );
  INV_X1 U9698 ( .A(SI_26_), .ZN(n11581) );
  INV_X1 U9699 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n11629) );
  INV_X1 U9700 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n11630) );
  MUX2_X1 U9701 ( .A(n11629), .B(n11630), .S(n6459), .Z(n7713) );
  INV_X1 U9702 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n11846) );
  INV_X1 U9703 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13313) );
  MUX2_X1 U9704 ( .A(n11846), .B(n13313), .S(n6459), .Z(n8552) );
  XNOR2_X1 U9705 ( .A(n8552), .B(SI_27_), .ZN(n7503) );
  NOR2_X1 U9706 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n7507) );
  NOR2_X1 U9707 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7506) );
  INV_X1 U9708 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7504) );
  NAND4_X1 U9709 ( .A1(n7507), .A2(n7506), .A3(n7505), .A4(n7504), .ZN(n7511)
         );
  INV_X1 U9710 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n7508) );
  NAND4_X1 U9711 ( .A1(n8028), .A2(n7402), .A3(n7509), .A4(n7508), .ZN(n7510)
         );
  INV_X1 U9712 ( .A(n7518), .ZN(n7519) );
  NAND2_X1 U9713 ( .A1(n11845), .A2(n9469), .ZN(n7522) );
  NAND2_X1 U9714 ( .A1(n9485), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7521) );
  XNOR2_X1 U9715 ( .A(n8455), .B(n7523), .ZN(n11847) );
  NAND2_X1 U9716 ( .A1(n11847), .A2(n9469), .ZN(n7525) );
  NAND2_X1 U9717 ( .A1(n9485), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n7524) );
  XNOR2_X1 U9718 ( .A(n7640), .B(SI_14_), .ZN(n7639) );
  XNOR2_X1 U9719 ( .A(n7639), .B(n7526), .ZN(n10366) );
  NAND2_X1 U9720 ( .A1(n10366), .A2(n9469), .ZN(n7530) );
  NAND2_X1 U9721 ( .A1(n6819), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7527) );
  XNOR2_X1 U9722 ( .A(n7527), .B(P2_IR_REG_14__SCAN_IN), .ZN(n14675) );
  INV_X1 U9723 ( .A(n14675), .ZN(n12919) );
  OAI22_X1 U9724 ( .A1(n6440), .A2(n10369), .B1(n9862), .B2(n12919), .ZN(n7528) );
  INV_X1 U9725 ( .A(n7528), .ZN(n7529) );
  INV_X1 U9726 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7534) );
  NAND2_X1 U9727 ( .A1(n6459), .A2(SI_0_), .ZN(n7531) );
  NAND2_X1 U9728 ( .A1(n7531), .A2(n8705), .ZN(n7533) );
  NAND2_X1 U9729 ( .A1(n7533), .A2(n7532), .ZN(n13315) );
  MUX2_X1 U9730 ( .A(n7534), .B(n13315), .S(n7538), .Z(n10561) );
  INV_X1 U9731 ( .A(n10561), .ZN(n14773) );
  XNOR2_X1 U9732 ( .A(n7535), .B(n7536), .ZN(n8083) );
  INV_X1 U9733 ( .A(n8083), .ZN(n9751) );
  INV_X1 U9734 ( .A(n7538), .ZN(n7617) );
  NAND2_X1 U9735 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7539) );
  MUX2_X1 U9736 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7539), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n7541) );
  INV_X1 U9737 ( .A(n7540), .ZN(n7547) );
  NAND2_X1 U9738 ( .A1(n7541), .A2(n7547), .ZN(n9879) );
  INV_X1 U9739 ( .A(n9879), .ZN(n9908) );
  NAND2_X1 U9740 ( .A1(n7617), .A2(n9908), .ZN(n7542) );
  NOR2_X1 U9741 ( .A1(n14773), .A2(n10889), .ZN(n10872) );
  NAND2_X1 U9742 ( .A1(n7547), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7548) );
  XNOR2_X1 U9743 ( .A(n7548), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9919) );
  NAND2_X1 U9744 ( .A1(n7617), .A2(n9919), .ZN(n7549) );
  OAI211_X2 U9745 ( .C1(n9747), .C2(n7543), .A(n7550), .B(n7549), .ZN(n10881)
         );
  INV_X1 U9746 ( .A(n10881), .ZN(n14779) );
  AND2_X1 U9747 ( .A1(n10872), .A2(n14779), .ZN(n10870) );
  XNOR2_X1 U9748 ( .A(n7552), .B(n7551), .ZN(n9754) );
  INV_X1 U9749 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7553) );
  AND2_X1 U9750 ( .A1(n7540), .A2(n7553), .ZN(n7622) );
  INV_X1 U9751 ( .A(n7622), .ZN(n7559) );
  NAND2_X1 U9752 ( .A1(n7559), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7554) );
  XNOR2_X1 U9753 ( .A(n7554), .B(P2_IR_REG_3__SCAN_IN), .ZN(n14608) );
  NAND2_X1 U9754 ( .A1(n7617), .A2(n14608), .ZN(n7555) );
  NAND2_X1 U9755 ( .A1(n10870), .A2(n10825), .ZN(n11277) );
  XNOR2_X1 U9756 ( .A(n7556), .B(n7557), .ZN(n9764) );
  NAND2_X1 U9757 ( .A1(n9764), .A2(n7009), .ZN(n7563) );
  NAND2_X1 U9758 ( .A1(n7566), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7560) );
  XNOR2_X1 U9759 ( .A(n7558), .B(n7560), .ZN(n9902) );
  OAI22_X1 U9760 ( .A1(n6440), .A2(n9767), .B1(n9862), .B2(n9902), .ZN(n7561)
         );
  INV_X1 U9761 ( .A(n7561), .ZN(n7562) );
  NAND2_X1 U9762 ( .A1(n7563), .A2(n7562), .ZN(n14793) );
  XNOR2_X1 U9763 ( .A(n7564), .B(n7565), .ZN(n9780) );
  NAND2_X1 U9764 ( .A1(n9780), .A2(n9469), .ZN(n7572) );
  INV_X1 U9765 ( .A(n7566), .ZN(n7567) );
  NAND2_X1 U9766 ( .A1(n7567), .A2(n7558), .ZN(n7575) );
  NAND2_X1 U9767 ( .A1(n7575), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7569) );
  XNOR2_X1 U9768 ( .A(n7569), .B(n7568), .ZN(n10011) );
  OAI22_X1 U9769 ( .A1(n6440), .A2(n9781), .B1(n9862), .B2(n10011), .ZN(n7570)
         );
  INV_X1 U9770 ( .A(n7570), .ZN(n7571) );
  NAND2_X1 U9771 ( .A1(n7572), .A2(n7571), .ZN(n11032) );
  INV_X1 U9772 ( .A(n11032), .ZN(n14801) );
  NAND2_X1 U9773 ( .A1(n11276), .A2(n14801), .ZN(n11045) );
  XNOR2_X1 U9774 ( .A(n7573), .B(n7574), .ZN(n9785) );
  NAND2_X1 U9775 ( .A1(n9785), .A2(n9469), .ZN(n7579) );
  INV_X1 U9776 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9788) );
  NAND2_X1 U9777 ( .A1(n7582), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7576) );
  INV_X1 U9778 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7583) );
  XNOR2_X1 U9779 ( .A(n7576), .B(n7583), .ZN(n14619) );
  OAI22_X1 U9780 ( .A1(n6440), .A2(n9788), .B1(n9862), .B2(n14619), .ZN(n7577)
         );
  INV_X1 U9781 ( .A(n7577), .ZN(n7578) );
  NAND2_X1 U9782 ( .A1(n7579), .A2(n7578), .ZN(n11048) );
  OR2_X1 U9783 ( .A1(n11045), .A2(n11048), .ZN(n11246) );
  XNOR2_X1 U9784 ( .A(n7580), .B(n7581), .ZN(n9789) );
  NAND2_X1 U9785 ( .A1(n9789), .A2(n9469), .ZN(n7589) );
  INV_X1 U9786 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9790) );
  INV_X1 U9787 ( .A(n7582), .ZN(n7584) );
  NAND2_X1 U9788 ( .A1(n7584), .A2(n7583), .ZN(n7592) );
  NAND2_X1 U9789 ( .A1(n7592), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7586) );
  INV_X1 U9790 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n7585) );
  XNOR2_X1 U9791 ( .A(n7586), .B(n7585), .ZN(n14632) );
  OAI22_X1 U9792 ( .A1(n6440), .A2(n9790), .B1(n9862), .B2(n14632), .ZN(n7587)
         );
  INV_X1 U9793 ( .A(n7587), .ZN(n7588) );
  NAND2_X1 U9794 ( .A1(n7589), .A2(n7588), .ZN(n11247) );
  XNOR2_X1 U9795 ( .A(n7590), .B(n7591), .ZN(n9836) );
  NAND2_X1 U9796 ( .A1(n9836), .A2(n9469), .ZN(n7597) );
  INV_X1 U9797 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9837) );
  NAND2_X1 U9798 ( .A1(n7600), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7594) );
  INV_X1 U9799 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7593) );
  XNOR2_X1 U9800 ( .A(n7594), .B(n7593), .ZN(n14645) );
  OAI22_X1 U9801 ( .A1(n6440), .A2(n9837), .B1(n9862), .B2(n14645), .ZN(n7595)
         );
  INV_X1 U9802 ( .A(n7595), .ZN(n7596) );
  XNOR2_X1 U9803 ( .A(n7598), .B(n7599), .ZN(n9846) );
  NAND2_X1 U9804 ( .A1(n9846), .A2(n9469), .ZN(n7604) );
  INV_X1 U9805 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9849) );
  NAND2_X1 U9806 ( .A1(n7607), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7601) );
  INV_X1 U9807 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7608) );
  XNOR2_X1 U9808 ( .A(n7601), .B(n7608), .ZN(n10083) );
  OAI22_X1 U9809 ( .A1(n6440), .A2(n9849), .B1(n9862), .B2(n10083), .ZN(n7602)
         );
  INV_X1 U9810 ( .A(n7602), .ZN(n7603) );
  INV_X1 U9811 ( .A(n14829), .ZN(n11210) );
  NAND2_X1 U9812 ( .A1(n9851), .A2(n9469), .ZN(n7612) );
  INV_X1 U9813 ( .A(n7607), .ZN(n7609) );
  NAND2_X1 U9814 ( .A1(n7609), .A2(n7608), .ZN(n7615) );
  NAND2_X1 U9815 ( .A1(n7615), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7610) );
  XNOR2_X1 U9816 ( .A(n7610), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10102) );
  AOI22_X1 U9817 ( .A1(n9485), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n10102), 
        .B2(n7617), .ZN(n7611) );
  XNOR2_X1 U9818 ( .A(n7613), .B(n7614), .ZN(n9857) );
  NAND2_X1 U9819 ( .A1(n9857), .A2(n9469), .ZN(n7619) );
  OAI21_X1 U9820 ( .B1(n7615), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7616) );
  XNOR2_X1 U9821 ( .A(n7616), .B(P2_IR_REG_11__SCAN_IN), .ZN(n12903) );
  AOI22_X1 U9822 ( .A1(n12903), .A2(n7617), .B1(n9485), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n7618) );
  XNOR2_X1 U9823 ( .A(n7620), .B(n7376), .ZN(n9925) );
  NAND2_X1 U9824 ( .A1(n9925), .A2(n9469), .ZN(n7629) );
  NAND4_X1 U9825 ( .A1(n7624), .A2(n7623), .A3(n7622), .A4(n7621), .ZN(n7632)
         );
  NAND2_X1 U9826 ( .A1(n7632), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7626) );
  INV_X1 U9827 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7625) );
  XNOR2_X1 U9828 ( .A(n7626), .B(n7625), .ZN(n12928) );
  OAI22_X1 U9829 ( .A1(n6440), .A2(n9926), .B1(n9862), .B2(n12928), .ZN(n7627)
         );
  INV_X1 U9830 ( .A(n7627), .ZN(n7628) );
  INV_X1 U9831 ( .A(n13273), .ZN(n11566) );
  XNOR2_X1 U9832 ( .A(n7630), .B(n7631), .ZN(n10075) );
  NAND2_X1 U9833 ( .A1(n10075), .A2(n9469), .ZN(n7637) );
  OAI21_X1 U9834 ( .B1(n7632), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7633) );
  MUX2_X1 U9835 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7633), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n7634) );
  AND2_X1 U9836 ( .A1(n7634), .A2(n6819), .ZN(n12931) );
  INV_X1 U9837 ( .A(n12931), .ZN(n14660) );
  OAI22_X1 U9838 ( .A1(n6440), .A2(n10078), .B1(n9862), .B2(n14660), .ZN(n7635) );
  INV_X1 U9839 ( .A(n7635), .ZN(n7636) );
  NAND2_X1 U9840 ( .A1(n11563), .A2(n11600), .ZN(n11704) );
  NAND2_X1 U9841 ( .A1(n7639), .A2(n7638), .ZN(n7643) );
  INV_X1 U9842 ( .A(n7640), .ZN(n7641) );
  NAND2_X1 U9843 ( .A1(n7641), .A2(SI_14_), .ZN(n7642) );
  NAND2_X1 U9844 ( .A1(n7643), .A2(n7642), .ZN(n7647) );
  NAND2_X1 U9845 ( .A1(n7645), .A2(n7644), .ZN(n7646) );
  NAND2_X1 U9846 ( .A1(n10452), .A2(n9469), .ZN(n7652) );
  INV_X1 U9847 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10455) );
  NAND2_X1 U9848 ( .A1(n7648), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7649) );
  XNOR2_X1 U9849 ( .A(n7649), .B(n7392), .ZN(n14678) );
  OAI22_X1 U9850 ( .A1(n6440), .A2(n10455), .B1(n9862), .B2(n14678), .ZN(n7650) );
  INV_X1 U9851 ( .A(n7650), .ZN(n7651) );
  XNOR2_X1 U9852 ( .A(n7654), .B(n7653), .ZN(n10361) );
  NAND2_X1 U9853 ( .A1(n10361), .A2(n9469), .ZN(n7659) );
  NAND2_X1 U9854 ( .A1(n7655), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7656) );
  XNOR2_X1 U9855 ( .A(n7656), .B(P2_IR_REG_16__SCAN_IN), .ZN(n14699) );
  INV_X1 U9856 ( .A(n14699), .ZN(n10362) );
  OAI22_X1 U9857 ( .A1(n6440), .A2(n10363), .B1(n9862), .B2(n10362), .ZN(n7657) );
  INV_X1 U9858 ( .A(n7657), .ZN(n7658) );
  XNOR2_X1 U9859 ( .A(n7661), .B(n7660), .ZN(n10466) );
  NAND2_X1 U9860 ( .A1(n10466), .A2(n9469), .ZN(n7668) );
  NAND2_X1 U9861 ( .A1(n7663), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7664) );
  MUX2_X1 U9862 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7664), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n7665) );
  AND2_X1 U9863 ( .A1(n7662), .A2(n7665), .ZN(n14712) );
  INV_X1 U9864 ( .A(n14712), .ZN(n10469) );
  OAI22_X1 U9865 ( .A1(n6440), .A2(n10471), .B1(n9862), .B2(n10469), .ZN(n7666) );
  INV_X1 U9866 ( .A(n7666), .ZN(n7667) );
  INV_X1 U9867 ( .A(n13258), .ZN(n13179) );
  XNOR2_X1 U9868 ( .A(n7676), .B(SI_18_), .ZN(n7675) );
  INV_X1 U9869 ( .A(n7674), .ZN(n7669) );
  XNOR2_X1 U9870 ( .A(n7675), .B(n7669), .ZN(n10755) );
  NAND2_X1 U9871 ( .A1(n10755), .A2(n9469), .ZN(n7673) );
  INV_X1 U9872 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10758) );
  NAND2_X1 U9873 ( .A1(n7662), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7670) );
  XNOR2_X1 U9874 ( .A(n7670), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14727) );
  INV_X1 U9875 ( .A(n14727), .ZN(n12935) );
  OAI22_X1 U9876 ( .A1(n6440), .A2(n10758), .B1(n12935), .B2(n9862), .ZN(n7671) );
  INV_X1 U9877 ( .A(n7671), .ZN(n7672) );
  NAND2_X1 U9878 ( .A1(n7675), .A2(n7674), .ZN(n7679) );
  INV_X1 U9879 ( .A(n7676), .ZN(n7677) );
  NAND2_X1 U9880 ( .A1(n7677), .A2(SI_18_), .ZN(n7678) );
  NAND2_X1 U9881 ( .A1(n7679), .A2(n7678), .ZN(n7683) );
  NAND2_X1 U9882 ( .A1(n7681), .A2(n7680), .ZN(n7682) );
  NAND2_X1 U9883 ( .A1(n10847), .A2(n9469), .ZN(n7687) );
  INV_X1 U9884 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10850) );
  OAI22_X1 U9885 ( .A1(n6440), .A2(n10850), .B1(n11725), .B2(n9862), .ZN(n7685) );
  INV_X1 U9886 ( .A(n7685), .ZN(n7686) );
  XNOR2_X1 U9887 ( .A(n7688), .B(n7689), .ZN(n10866) );
  NAND2_X1 U9888 ( .A1(n10866), .A2(n9469), .ZN(n7691) );
  NAND2_X1 U9889 ( .A1(n9485), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7690) );
  XNOR2_X1 U9890 ( .A(n7693), .B(n7692), .ZN(n10944) );
  NAND2_X1 U9891 ( .A1(n10944), .A2(n9469), .ZN(n7695) );
  NAND2_X1 U9892 ( .A1(n9485), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7694) );
  NAND2_X1 U9893 ( .A1(n8455), .A2(n7696), .ZN(n7699) );
  NAND2_X1 U9894 ( .A1(n7697), .A2(SI_22_), .ZN(n7698) );
  XNOR2_X1 U9895 ( .A(n7700), .B(SI_23_), .ZN(n7701) );
  NAND2_X1 U9896 ( .A1(n11343), .A2(n9469), .ZN(n7704) );
  NAND2_X1 U9897 ( .A1(n9485), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7703) );
  NAND2_X1 U9898 ( .A1(n11429), .A2(n9469), .ZN(n7708) );
  NAND2_X1 U9899 ( .A1(n9485), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7707) );
  AND2_X2 U9900 ( .A1(n7708), .A2(n7707), .ZN(n13219) );
  XNOR2_X1 U9901 ( .A(n7710), .B(n7709), .ZN(n11500) );
  NAND2_X1 U9902 ( .A1(n11500), .A2(n9469), .ZN(n7712) );
  NAND2_X1 U9903 ( .A1(n9485), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7711) );
  AND2_X2 U9904 ( .A1(n13054), .A2(n13038), .ZN(n13040) );
  XNOR2_X1 U9905 ( .A(n7713), .B(SI_26_), .ZN(n7714) );
  NAND2_X1 U9906 ( .A1(n11626), .A2(n9469), .ZN(n7717) );
  NAND2_X1 U9907 ( .A1(n9485), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7716) );
  INV_X2 U9908 ( .A(n9596), .ZN(n9578) );
  AOI211_X1 U9909 ( .C1(n12772), .C2(n13022), .A(n13190), .B(n12992), .ZN(
        n13002) );
  INV_X1 U9910 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7718) );
  NAND2_X1 U9911 ( .A1(n7719), .A2(n7718), .ZN(n13297) );
  NAND2_X1 U9912 ( .A1(n7720), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7721) );
  INV_X1 U9913 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7722) );
  NAND2_X1 U9914 ( .A1(n7737), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7727) );
  AND2_X2 U9915 ( .A1(n13302), .A2(n13305), .ZN(n7754) );
  NAND2_X1 U9916 ( .A1(n6446), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7726) );
  AND2_X2 U9917 ( .A1(n7724), .A2(n13305), .ZN(n7759) );
  NAND2_X1 U9918 ( .A1(n7759), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7725) );
  NAND2_X1 U9919 ( .A1(n6446), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7733) );
  NAND2_X1 U9920 ( .A1(n7737), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7732) );
  INV_X1 U9921 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7729) );
  NAND2_X1 U9922 ( .A1(n7759), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7730) );
  INV_X1 U9923 ( .A(n12899), .ZN(n7734) );
  NAND2_X1 U9924 ( .A1(n7734), .A2(n14773), .ZN(n9580) );
  NAND2_X1 U9925 ( .A1(n9529), .A2(n10557), .ZN(n7736) );
  INV_X1 U9926 ( .A(n12898), .ZN(n10478) );
  NAND2_X1 U9927 ( .A1(n10478), .A2(n10889), .ZN(n7735) );
  NAND2_X1 U9928 ( .A1(n7759), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7742) );
  INV_X1 U9929 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7738) );
  INV_X1 U9930 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7739) );
  NAND2_X1 U9931 ( .A1(n10424), .A2(n10881), .ZN(n10820) );
  NAND2_X1 U9932 ( .A1(n12897), .A2(n14779), .ZN(n7743) );
  NAND2_X1 U9933 ( .A1(n7759), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7746) );
  INV_X1 U9934 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7744) );
  NAND2_X1 U9935 ( .A1(n6446), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7745) );
  NAND2_X1 U9936 ( .A1(n11273), .A2(n14785), .ZN(n11268) );
  NAND2_X1 U9937 ( .A1(n12896), .A2(n10825), .ZN(n7747) );
  NAND2_X1 U9938 ( .A1(n6446), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7752) );
  OAI21_X1 U9939 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n7757), .ZN(n10672) );
  INV_X1 U9940 ( .A(n10672), .ZN(n11275) );
  NAND2_X1 U9941 ( .A1(n7737), .A2(n11275), .ZN(n7751) );
  NAND2_X1 U9942 ( .A1(n9488), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7750) );
  NAND2_X1 U9943 ( .A1(n7759), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7749) );
  NAND4_X1 U9944 ( .A1(n7752), .A2(n7751), .A3(n7750), .A4(n7749), .ZN(n12895)
         );
  INV_X1 U9945 ( .A(n14793), .ZN(n11280) );
  NAND2_X1 U9946 ( .A1(n12895), .A2(n11280), .ZN(n7753) );
  NAND2_X1 U9947 ( .A1(n6445), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7763) );
  INV_X1 U9948 ( .A(n7757), .ZN(n7755) );
  NAND2_X1 U9949 ( .A1(n7755), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7768) );
  INV_X1 U9950 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U9951 ( .A1(n7757), .A2(n7756), .ZN(n7758) );
  AND2_X1 U9952 ( .A1(n7768), .A2(n7758), .ZN(n11031) );
  NAND2_X1 U9953 ( .A1(n7737), .A2(n11031), .ZN(n7762) );
  NAND2_X1 U9954 ( .A1(n9488), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7761) );
  NAND2_X1 U9955 ( .A1(n7964), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7760) );
  NAND4_X1 U9956 ( .A1(n7763), .A2(n7762), .A3(n7761), .A4(n7760), .ZN(n12894)
         );
  INV_X1 U9957 ( .A(n12894), .ZN(n11274) );
  NAND2_X1 U9958 ( .A1(n11274), .A2(n11032), .ZN(n7765) );
  NAND2_X1 U9959 ( .A1(n14801), .A2(n12894), .ZN(n7764) );
  NAND2_X1 U9960 ( .A1(n7765), .A2(n7764), .ZN(n11025) );
  NAND2_X1 U9961 ( .A1(n11027), .A2(n7765), .ZN(n11041) );
  NAND2_X1 U9962 ( .A1(n7964), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7773) );
  NAND2_X1 U9963 ( .A1(n9488), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7772) );
  INV_X1 U9964 ( .A(n7768), .ZN(n7766) );
  NAND2_X1 U9965 ( .A1(n7766), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7777) );
  INV_X1 U9966 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7767) );
  NAND2_X1 U9967 ( .A1(n7768), .A2(n7767), .ZN(n7769) );
  AND2_X1 U9968 ( .A1(n7777), .A2(n7769), .ZN(n11047) );
  NAND2_X1 U9969 ( .A1(n7737), .A2(n11047), .ZN(n7771) );
  NAND2_X1 U9970 ( .A1(n6445), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7770) );
  NAND4_X1 U9971 ( .A1(n7773), .A2(n7772), .A3(n7771), .A4(n7770), .ZN(n12893)
         );
  XNOR2_X1 U9972 ( .A(n11048), .B(n12893), .ZN(n11040) );
  NAND2_X1 U9973 ( .A1(n11041), .A2(n11040), .ZN(n11039) );
  INV_X1 U9974 ( .A(n12893), .ZN(n10691) );
  NAND2_X1 U9975 ( .A1(n11048), .A2(n10691), .ZN(n7774) );
  NAND2_X1 U9976 ( .A1(n7964), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7782) );
  NAND2_X1 U9977 ( .A1(n9488), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7781) );
  INV_X1 U9978 ( .A(n7777), .ZN(n7775) );
  INV_X1 U9979 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7776) );
  NAND2_X1 U9980 ( .A1(n7777), .A2(n7776), .ZN(n7778) );
  AND2_X1 U9981 ( .A1(n7794), .A2(n7778), .ZN(n11248) );
  NAND2_X1 U9982 ( .A1(n7737), .A2(n11248), .ZN(n7780) );
  NAND2_X1 U9983 ( .A1(n6445), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7779) );
  NAND4_X1 U9984 ( .A1(n7782), .A2(n7781), .A3(n7780), .A4(n7779), .ZN(n12892)
         );
  INV_X1 U9985 ( .A(n12892), .ZN(n10680) );
  OR2_X1 U9986 ( .A1(n11247), .A2(n10680), .ZN(n7783) );
  NAND2_X1 U9987 ( .A1(n11247), .A2(n10680), .ZN(n7784) );
  NAND2_X1 U9988 ( .A1(n7964), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7789) );
  XNOR2_X1 U9989 ( .A(n7794), .B(P2_REG3_REG_8__SCAN_IN), .ZN(n11231) );
  NAND2_X1 U9990 ( .A1(n7737), .A2(n11231), .ZN(n7788) );
  NAND2_X1 U9991 ( .A1(n9488), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U9992 ( .A1(n6445), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7786) );
  NAND4_X1 U9993 ( .A1(n7789), .A2(n7788), .A3(n7787), .A4(n7786), .ZN(n12891)
         );
  INV_X1 U9994 ( .A(n11223), .ZN(n11217) );
  INV_X1 U9995 ( .A(n12891), .ZN(n11085) );
  OR2_X1 U9996 ( .A1(n11227), .A2(n11085), .ZN(n7790) );
  NAND2_X1 U9997 ( .A1(n6446), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7800) );
  INV_X1 U9998 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10732) );
  INV_X1 U9999 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7792) );
  OAI21_X1 U10000 ( .B1(n7794), .B2(n10732), .A(n7792), .ZN(n7795) );
  NAND2_X1 U10001 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n7793) );
  AND2_X1 U10002 ( .A1(n7795), .A2(n7804), .ZN(n11211) );
  NAND2_X1 U10003 ( .A1(n7737), .A2(n11211), .ZN(n7799) );
  NAND2_X1 U10004 ( .A1(n9488), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7798) );
  NAND2_X1 U10005 ( .A1(n7964), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7797) );
  NAND4_X1 U10006 ( .A1(n7800), .A2(n7799), .A3(n7798), .A4(n7797), .ZN(n12890) );
  INV_X1 U10007 ( .A(n12890), .ZN(n7801) );
  XNOR2_X1 U10008 ( .A(n14829), .B(n7801), .ZN(n11207) );
  INV_X1 U10009 ( .A(n11207), .ZN(n11202) );
  NAND2_X1 U10010 ( .A1(n11203), .A2(n11202), .ZN(n11201) );
  OR2_X1 U10011 ( .A1(n14829), .A2(n7801), .ZN(n7802) );
  NAND2_X1 U10012 ( .A1(n11201), .A2(n7802), .ZN(n10983) );
  NAND2_X1 U10013 ( .A1(n7964), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7809) );
  INV_X1 U10014 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n15072) );
  NAND2_X1 U10015 ( .A1(n7804), .A2(n15072), .ZN(n7805) );
  AND2_X1 U10016 ( .A1(n7820), .A2(n7805), .ZN(n11144) );
  NAND2_X1 U10017 ( .A1(n7737), .A2(n11144), .ZN(n7808) );
  NAND2_X1 U10018 ( .A1(n9488), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7807) );
  NAND2_X1 U10019 ( .A1(n6445), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7806) );
  NAND4_X1 U10020 ( .A1(n7809), .A2(n7808), .A3(n7807), .A4(n7806), .ZN(n12889) );
  INV_X1 U10021 ( .A(n12889), .ZN(n11256) );
  XNOR2_X1 U10022 ( .A(n14842), .B(n11256), .ZN(n10978) );
  OR2_X1 U10023 ( .A1(n14842), .A2(n11256), .ZN(n7810) );
  NAND2_X1 U10024 ( .A1(n6446), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7814) );
  XNOR2_X1 U10025 ( .A(n7820), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n11263) );
  NAND2_X1 U10026 ( .A1(n7737), .A2(n11263), .ZN(n7813) );
  NAND2_X1 U10027 ( .A1(n9488), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7812) );
  NAND2_X1 U10028 ( .A1(n7964), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7811) );
  NAND4_X1 U10029 ( .A1(n7814), .A2(n7813), .A3(n7812), .A4(n7811), .ZN(n12888) );
  INV_X1 U10030 ( .A(n12888), .ZN(n11555) );
  XNOR2_X1 U10031 ( .A(n11253), .B(n11555), .ZN(n11149) );
  NAND2_X1 U10032 ( .A1(n11253), .A2(n11555), .ZN(n7816) );
  NAND2_X1 U10033 ( .A1(n7964), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7825) );
  NAND2_X1 U10034 ( .A1(n9488), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7824) );
  INV_X1 U10035 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7818) );
  INV_X1 U10036 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7817) );
  OAI21_X1 U10037 ( .B1(n7820), .B2(n7818), .A(n7817), .ZN(n7821) );
  NAND2_X1 U10038 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n7819) );
  AND2_X1 U10039 ( .A1(n7821), .A2(n7828), .ZN(n11564) );
  NAND2_X1 U10040 ( .A1(n7737), .A2(n11564), .ZN(n7823) );
  NAND2_X1 U10041 ( .A1(n6445), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7822) );
  NAND4_X1 U10042 ( .A1(n7825), .A2(n7824), .A3(n7823), .A4(n7822), .ZN(n12887) );
  XNOR2_X1 U10043 ( .A(n13273), .B(n12887), .ZN(n9534) );
  INV_X1 U10044 ( .A(n9534), .ZN(n11559) );
  INV_X1 U10045 ( .A(n12887), .ZN(n7826) );
  OR2_X1 U10046 ( .A1(n13273), .A2(n7826), .ZN(n11468) );
  NAND2_X1 U10047 ( .A1(n6446), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7833) );
  INV_X1 U10048 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n15172) );
  NAND2_X1 U10049 ( .A1(n7828), .A2(n15172), .ZN(n7829) );
  AND2_X1 U10050 ( .A1(n7837), .A2(n7829), .ZN(n11475) );
  NAND2_X1 U10051 ( .A1(n7737), .A2(n11475), .ZN(n7832) );
  NAND2_X1 U10052 ( .A1(n9488), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7831) );
  NAND2_X1 U10053 ( .A1(n7964), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7830) );
  NAND4_X1 U10054 ( .A1(n7833), .A2(n7832), .A3(n7831), .A4(n7830), .ZN(n12886) );
  XNOR2_X1 U10055 ( .A(n9640), .B(n12886), .ZN(n11474) );
  NAND2_X1 U10056 ( .A1(n7834), .A2(n11474), .ZN(n11467) );
  INV_X1 U10057 ( .A(n12886), .ZN(n11554) );
  OR2_X1 U10058 ( .A1(n9640), .A2(n11554), .ZN(n7835) );
  NAND2_X1 U10059 ( .A1(n6445), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7842) );
  INV_X1 U10060 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7836) );
  NAND2_X1 U10061 ( .A1(n7837), .A2(n7836), .ZN(n7838) );
  AND2_X1 U10062 ( .A1(n7846), .A2(n7838), .ZN(n11898) );
  NAND2_X1 U10063 ( .A1(n7737), .A2(n11898), .ZN(n7841) );
  NAND2_X1 U10064 ( .A1(n9488), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7840) );
  NAND2_X1 U10065 ( .A1(n7759), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7839) );
  NAND4_X1 U10066 ( .A1(n7842), .A2(n7841), .A3(n7840), .A4(n7839), .ZN(n12885) );
  INV_X1 U10067 ( .A(n12885), .ZN(n11452) );
  XNOR2_X1 U10068 ( .A(n11730), .B(n11452), .ZN(n11708) );
  NAND2_X1 U10069 ( .A1(n11730), .A2(n11452), .ZN(n7844) );
  NAND2_X1 U10070 ( .A1(n6446), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7851) );
  INV_X1 U10071 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7845) );
  NAND2_X1 U10072 ( .A1(n7846), .A2(n7845), .ZN(n7847) );
  AND2_X1 U10073 ( .A1(n7854), .A2(n7847), .ZN(n11724) );
  NAND2_X1 U10074 ( .A1(n7737), .A2(n11724), .ZN(n7850) );
  NAND2_X1 U10075 ( .A1(n9488), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7849) );
  NAND2_X1 U10076 ( .A1(n7964), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7848) );
  NAND4_X1 U10077 ( .A1(n7851), .A2(n7850), .A3(n7849), .A4(n7848), .ZN(n12884) );
  INV_X1 U10078 ( .A(n12884), .ZN(n11711) );
  XNOR2_X1 U10079 ( .A(n13269), .B(n11711), .ZN(n11718) );
  OR2_X1 U10080 ( .A1(n13269), .A2(n11711), .ZN(n11742) );
  NAND2_X1 U10081 ( .A1(n11717), .A2(n11742), .ZN(n7860) );
  NAND2_X1 U10082 ( .A1(n7759), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7859) );
  NAND2_X1 U10083 ( .A1(n9488), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7858) );
  INV_X1 U10084 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n11837) );
  NAND2_X1 U10085 ( .A1(n7854), .A2(n11837), .ZN(n7855) );
  AND2_X1 U10086 ( .A1(n7864), .A2(n7855), .ZN(n11840) );
  NAND2_X1 U10087 ( .A1(n7737), .A2(n11840), .ZN(n7857) );
  NAND2_X1 U10088 ( .A1(n6446), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7856) );
  NAND4_X1 U10089 ( .A1(n7859), .A2(n7858), .A3(n7857), .A4(n7856), .ZN(n12883) );
  XNOR2_X1 U10090 ( .A(n13262), .B(n12883), .ZN(n11741) );
  INV_X1 U10091 ( .A(n12883), .ZN(n11826) );
  OR2_X1 U10092 ( .A1(n13262), .A2(n11826), .ZN(n7861) );
  INV_X1 U10093 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7863) );
  NAND2_X1 U10094 ( .A1(n7864), .A2(n7863), .ZN(n7865) );
  AND2_X1 U10095 ( .A1(n7873), .A2(n7865), .ZN(n13176) );
  NAND2_X1 U10096 ( .A1(n13176), .A2(n7737), .ZN(n7869) );
  NAND2_X1 U10097 ( .A1(n7759), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7868) );
  NAND2_X1 U10098 ( .A1(n9488), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7867) );
  NAND2_X1 U10099 ( .A1(n6445), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7866) );
  NAND4_X1 U10100 ( .A1(n7869), .A2(n7868), .A3(n7867), .A4(n7866), .ZN(n13151) );
  INV_X1 U10101 ( .A(n13151), .ZN(n7992) );
  NAND2_X1 U10102 ( .A1(n13258), .A2(n7992), .ZN(n7870) );
  OR2_X1 U10103 ( .A1(n13258), .A2(n7992), .ZN(n7871) );
  INV_X1 U10104 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7872) );
  NAND2_X1 U10105 ( .A1(n7873), .A2(n7872), .ZN(n7874) );
  NAND2_X1 U10106 ( .A1(n7883), .A2(n7874), .ZN(n13159) );
  NAND2_X1 U10107 ( .A1(n6445), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7876) );
  NAND2_X1 U10108 ( .A1(n7759), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7875) );
  AND2_X1 U10109 ( .A1(n7876), .A2(n7875), .ZN(n7878) );
  NAND2_X1 U10110 ( .A1(n9488), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7877) );
  OAI211_X1 U10111 ( .C1(n13159), .C2(n6441), .A(n7878), .B(n7877), .ZN(n12882) );
  INV_X1 U10112 ( .A(n12882), .ZN(n12786) );
  NAND2_X1 U10113 ( .A1(n13253), .A2(n12786), .ZN(n7879) );
  OR2_X1 U10114 ( .A1(n13253), .A2(n12786), .ZN(n7880) );
  INV_X1 U10115 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n7887) );
  INV_X1 U10116 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7882) );
  NAND2_X1 U10117 ( .A1(n7883), .A2(n7882), .ZN(n7884) );
  NAND2_X1 U10118 ( .A1(n7890), .A2(n7884), .ZN(n13134) );
  OR2_X1 U10119 ( .A1(n13134), .A2(n6441), .ZN(n7886) );
  AOI22_X1 U10120 ( .A1(n9488), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n7759), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n7885) );
  OAI211_X1 U10121 ( .C1(n7791), .C2(n7887), .A(n7886), .B(n7885), .ZN(n13154)
         );
  INV_X1 U10122 ( .A(n13154), .ZN(n12833) );
  NAND2_X1 U10123 ( .A1(n13246), .A2(n12833), .ZN(n7889) );
  NOR2_X1 U10124 ( .A1(n13246), .A2(n12833), .ZN(n7888) );
  INV_X1 U10125 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n12827) );
  NAND2_X1 U10126 ( .A1(n7890), .A2(n12827), .ZN(n7891) );
  AND2_X1 U10127 ( .A1(n7897), .A2(n7891), .ZN(n13117) );
  NAND2_X1 U10128 ( .A1(n13117), .A2(n7737), .ZN(n7894) );
  AOI22_X1 U10129 ( .A1(n7759), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n6446), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n7893) );
  NAND2_X1 U10130 ( .A1(n9488), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n7892) );
  INV_X1 U10131 ( .A(n12797), .ZN(n12881) );
  INV_X1 U10132 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7896) );
  NAND2_X1 U10133 ( .A1(n7897), .A2(n7896), .ZN(n7898) );
  NAND2_X1 U10134 ( .A1(n7905), .A2(n7898), .ZN(n13100) );
  OR2_X1 U10135 ( .A1(n13100), .A2(n6441), .ZN(n7904) );
  INV_X1 U10136 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n7901) );
  NAND2_X1 U10137 ( .A1(n9488), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U10138 ( .A1(n6446), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7899) );
  OAI211_X1 U10139 ( .C1(n7796), .C2(n7901), .A(n7900), .B(n7899), .ZN(n7902)
         );
  INV_X1 U10140 ( .A(n7902), .ZN(n7903) );
  NAND2_X1 U10141 ( .A1(n7904), .A2(n7903), .ZN(n13079) );
  INV_X1 U10142 ( .A(n13079), .ZN(n12848) );
  INV_X1 U10143 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n12845) );
  NAND2_X1 U10144 ( .A1(n7905), .A2(n12845), .ZN(n7906) );
  AND2_X1 U10145 ( .A1(n7913), .A2(n7906), .ZN(n12844) );
  NAND2_X1 U10146 ( .A1(n12844), .A2(n7737), .ZN(n7911) );
  INV_X1 U10147 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n15140) );
  NAND2_X1 U10148 ( .A1(n6446), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n7908) );
  NAND2_X1 U10149 ( .A1(n7964), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n7907) );
  OAI211_X1 U10150 ( .C1(n15140), .C2(n6439), .A(n7908), .B(n7907), .ZN(n7909)
         );
  INV_X1 U10151 ( .A(n7909), .ZN(n7910) );
  INV_X1 U10152 ( .A(n13083), .ZN(n7912) );
  INV_X1 U10153 ( .A(n13066), .ZN(n12880) );
  INV_X1 U10154 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n12779) );
  NAND2_X1 U10155 ( .A1(n7913), .A2(n12779), .ZN(n7914) );
  NAND2_X1 U10156 ( .A1(n7921), .A2(n7914), .ZN(n12780) );
  INV_X1 U10157 ( .A(n12780), .ZN(n13072) );
  NAND2_X1 U10158 ( .A1(n13072), .A2(n7737), .ZN(n7920) );
  INV_X1 U10159 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n7917) );
  NAND2_X1 U10160 ( .A1(n7759), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n7916) );
  NAND2_X1 U10161 ( .A1(n6446), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n7915) );
  OAI211_X1 U10162 ( .C1(n6439), .C2(n7917), .A(n7916), .B(n7915), .ZN(n7918)
         );
  INV_X1 U10163 ( .A(n7918), .ZN(n7919) );
  XNOR2_X1 U10164 ( .A(n13226), .B(n13080), .ZN(n9539) );
  INV_X1 U10165 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n12822) );
  INV_X1 U10166 ( .A(n7930), .ZN(n7932) );
  NAND2_X1 U10167 ( .A1(n7921), .A2(n12822), .ZN(n7922) );
  NAND2_X1 U10168 ( .A1(n13055), .A2(n7737), .ZN(n7928) );
  INV_X1 U10169 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n7925) );
  NAND2_X1 U10170 ( .A1(n6446), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n7924) );
  NAND2_X1 U10171 ( .A1(n7759), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n7923) );
  OAI211_X1 U10172 ( .C1(n7925), .C2(n6439), .A(n7924), .B(n7923), .ZN(n7926)
         );
  INV_X1 U10173 ( .A(n7926), .ZN(n7927) );
  INV_X1 U10174 ( .A(n13052), .ZN(n7929) );
  NAND2_X1 U10175 ( .A1(n7930), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n7940) );
  INV_X1 U10176 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n7931) );
  NAND2_X1 U10177 ( .A1(n7932), .A2(n7931), .ZN(n7933) );
  NAND2_X1 U10178 ( .A1(n7940), .A2(n7933), .ZN(n13041) );
  OR2_X1 U10179 ( .A1(n13041), .A2(n6441), .ZN(n7938) );
  INV_X1 U10180 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n15110) );
  NAND2_X1 U10181 ( .A1(n9488), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n7935) );
  NAND2_X1 U10182 ( .A1(n7759), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n7934) );
  OAI211_X1 U10183 ( .C1(n7791), .C2(n15110), .A(n7935), .B(n7934), .ZN(n7936)
         );
  INV_X1 U10184 ( .A(n7936), .ZN(n7937) );
  XNOR2_X1 U10185 ( .A(n13214), .B(n9697), .ZN(n9542) );
  INV_X1 U10186 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7939) );
  NAND2_X1 U10187 ( .A1(n7940), .A2(n7939), .ZN(n7941) );
  NAND2_X1 U10188 ( .A1(n13025), .A2(n7737), .ZN(n7947) );
  INV_X1 U10189 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n7944) );
  NAND2_X1 U10190 ( .A1(n6446), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7943) );
  NAND2_X1 U10191 ( .A1(n7759), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n7942) );
  OAI211_X1 U10192 ( .C1(n7944), .C2(n6439), .A(n7943), .B(n7942), .ZN(n7945)
         );
  INV_X1 U10193 ( .A(n7945), .ZN(n7946) );
  NAND2_X1 U10194 ( .A1(n13209), .A2(n12814), .ZN(n7948) );
  OR2_X1 U10195 ( .A1(n13038), .A2(n13017), .ZN(n13016) );
  INV_X1 U10196 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n15074) );
  INV_X1 U10197 ( .A(n7961), .ZN(n7962) );
  NAND2_X1 U10198 ( .A1(n7951), .A2(n15074), .ZN(n7952) );
  NAND2_X1 U10199 ( .A1(n7962), .A2(n7952), .ZN(n13003) );
  OR2_X1 U10200 ( .A1(n13003), .A2(n6441), .ZN(n7958) );
  INV_X1 U10201 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n7955) );
  NAND2_X1 U10202 ( .A1(n7759), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n7954) );
  NAND2_X1 U10203 ( .A1(n6446), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7953) );
  OAI211_X1 U10204 ( .C1(n7955), .C2(n6439), .A(n7954), .B(n7953), .ZN(n7956)
         );
  INV_X1 U10205 ( .A(n7956), .ZN(n7957) );
  NAND2_X1 U10206 ( .A1(n9524), .A2(n12997), .ZN(n9492) );
  INV_X1 U10207 ( .A(n10947), .ZN(n9548) );
  NAND2_X1 U10208 ( .A1(n9548), .A2(n9723), .ZN(n7960) );
  INV_X1 U10209 ( .A(n13169), .ZN(n13064) );
  NAND2_X1 U10210 ( .A1(n7961), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n12965) );
  INV_X1 U10211 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9732) );
  NAND2_X1 U10212 ( .A1(n7962), .A2(n9732), .ZN(n7963) );
  NAND2_X1 U10213 ( .A1(n12965), .A2(n7963), .ZN(n12996) );
  INV_X1 U10214 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n7967) );
  NAND2_X1 U10215 ( .A1(n9488), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7966) );
  NAND2_X1 U10216 ( .A1(n6446), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7965) );
  OAI211_X1 U10217 ( .C1(n7796), .C2(n7967), .A(n7966), .B(n7965), .ZN(n7968)
         );
  INV_X1 U10218 ( .A(n7968), .ZN(n7969) );
  NAND2_X1 U10219 ( .A1(n9719), .A2(n7971), .ZN(n13069) );
  INV_X1 U10220 ( .A(n7971), .ZN(n9873) );
  INV_X1 U10221 ( .A(n7972), .ZN(n7973) );
  AND2_X1 U10222 ( .A1(n12899), .A2(n14773), .ZN(n10553) );
  OAI22_X1 U10223 ( .A1(n9529), .A2(n10553), .B1(n12898), .B2(n10889), .ZN(
        n10869) );
  INV_X1 U10224 ( .A(n10876), .ZN(n7974) );
  NAND2_X1 U10225 ( .A1(n10869), .A2(n7974), .ZN(n7976) );
  NAND2_X1 U10226 ( .A1(n10424), .A2(n14779), .ZN(n7975) );
  NAND2_X1 U10227 ( .A1(n7976), .A2(n7975), .ZN(n10815) );
  NAND2_X1 U10228 ( .A1(n10815), .A2(n10821), .ZN(n7978) );
  NAND2_X1 U10229 ( .A1(n11273), .A2(n10825), .ZN(n7977) );
  NAND2_X1 U10230 ( .A1(n7978), .A2(n7977), .ZN(n11267) );
  NAND2_X1 U10231 ( .A1(n11267), .A2(n11269), .ZN(n7980) );
  NAND2_X1 U10232 ( .A1(n10690), .A2(n11280), .ZN(n7979) );
  INV_X1 U10233 ( .A(n11040), .ZN(n11037) );
  OR2_X1 U10234 ( .A1(n11048), .A2(n12893), .ZN(n7981) );
  NAND2_X1 U10235 ( .A1(n7982), .A2(n7981), .ZN(n11243) );
  XNOR2_X1 U10236 ( .A(n11247), .B(n12892), .ZN(n11238) );
  INV_X1 U10237 ( .A(n11238), .ZN(n11242) );
  OR2_X1 U10238 ( .A1(n11247), .A2(n12892), .ZN(n7983) );
  NAND2_X1 U10239 ( .A1(n11208), .A2(n11207), .ZN(n11206) );
  NAND2_X1 U10240 ( .A1(n14829), .A2(n12890), .ZN(n7984) );
  NAND2_X1 U10241 ( .A1(n11253), .A2(n12888), .ZN(n7985) );
  OR2_X1 U10242 ( .A1(n13273), .A2(n12887), .ZN(n7987) );
  NOR2_X1 U10243 ( .A1(n11730), .A2(n12885), .ZN(n7989) );
  NAND2_X1 U10244 ( .A1(n11730), .A2(n12885), .ZN(n7988) );
  OR2_X1 U10245 ( .A1(n13269), .A2(n12884), .ZN(n7990) );
  NAND2_X1 U10246 ( .A1(n13262), .A2(n12883), .ZN(n7991) );
  XNOR2_X1 U10247 ( .A(n13258), .B(n7992), .ZN(n13180) );
  NAND2_X1 U10248 ( .A1(n13181), .A2(n13180), .ZN(n7994) );
  NAND2_X1 U10249 ( .A1(n13258), .A2(n13151), .ZN(n7993) );
  XNOR2_X1 U10250 ( .A(n13253), .B(n12882), .ZN(n13150) );
  OR2_X1 U10251 ( .A1(n13253), .A2(n12882), .ZN(n7995) );
  NAND2_X1 U10252 ( .A1(n13246), .A2(n13154), .ZN(n7996) );
  NAND2_X1 U10253 ( .A1(n13242), .A2(n12797), .ZN(n7997) );
  XOR2_X1 U10254 ( .A(n13079), .B(n13236), .Z(n13104) );
  AOI22_X1 U10255 ( .A1(n13105), .A2(n13104), .B1(n12848), .B2(n13103), .ZN(
        n13084) );
  NAND2_X1 U10256 ( .A1(n13084), .A2(n13083), .ZN(n13082) );
  NOR2_X1 U10257 ( .A1(n13214), .A2(n13017), .ZN(n7998) );
  INV_X1 U10258 ( .A(n12814), .ZN(n13035) );
  XNOR2_X1 U10259 ( .A(n12960), .B(n12959), .ZN(n13011) );
  NAND2_X1 U10260 ( .A1(n8000), .A2(n11725), .ZN(n14839) );
  NAND2_X1 U10261 ( .A1(n9303), .A2(n10893), .ZN(n14838) );
  NAND2_X1 U10262 ( .A1(n8004), .A2(n8003), .ZN(n13206) );
  NAND2_X1 U10263 ( .A1(n8029), .A2(n8028), .ZN(n8031) );
  NAND2_X1 U10264 ( .A1(n8031), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8006) );
  INV_X1 U10265 ( .A(P2_B_REG_SCAN_IN), .ZN(n8007) );
  XNOR2_X1 U10266 ( .A(n11432), .B(n8007), .ZN(n8011) );
  NAND2_X1 U10267 ( .A1(n8008), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8009) );
  MUX2_X1 U10268 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8009), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8010) );
  NAND2_X1 U10269 ( .A1(n8010), .A2(n6592), .ZN(n11503) );
  NAND2_X1 U10270 ( .A1(n8011), .A2(n11503), .ZN(n8015) );
  NAND2_X1 U10271 ( .A1(n6592), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8012) );
  MUX2_X1 U10272 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8012), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8014) );
  NAND2_X1 U10273 ( .A1(n8014), .A2(n8013), .ZN(n11632) );
  INV_X1 U10274 ( .A(n11632), .ZN(n8034) );
  INV_X1 U10275 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14765) );
  NAND2_X1 U10276 ( .A1(n14733), .A2(n14765), .ZN(n8017) );
  NAND2_X1 U10277 ( .A1(n11632), .A2(n11503), .ZN(n8016) );
  NAND2_X1 U10278 ( .A1(n8017), .A2(n8016), .ZN(n14766) );
  NAND2_X1 U10279 ( .A1(n13136), .A2(n12997), .ZN(n9726) );
  NAND2_X1 U10280 ( .A1(n14766), .A2(n9726), .ZN(n8033) );
  NOR4_X1 U10281 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8026) );
  INV_X1 U10282 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n15141) );
  INV_X1 U10283 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n15126) );
  INV_X1 U10284 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15169) );
  INV_X1 U10285 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n15159) );
  NAND4_X1 U10286 ( .A1(n15141), .A2(n15126), .A3(n15169), .A4(n15159), .ZN(
        n8023) );
  NOR4_X1 U10287 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n8021) );
  NOR4_X1 U10288 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n8020) );
  NOR4_X1 U10289 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n8019) );
  NOR4_X1 U10290 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n8018) );
  NAND4_X1 U10291 ( .A1(n8021), .A2(n8020), .A3(n8019), .A4(n8018), .ZN(n8022)
         );
  NOR4_X1 U10292 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        n8023), .A4(n8022), .ZN(n8025) );
  NOR4_X1 U10293 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8024) );
  NAND3_X1 U10294 ( .A1(n8026), .A2(n8025), .A3(n8024), .ZN(n8027) );
  AND2_X1 U10295 ( .A1(n14733), .A2(n8027), .ZN(n9718) );
  NAND2_X1 U10296 ( .A1(n9719), .A2(n9522), .ZN(n9728) );
  INV_X1 U10297 ( .A(n9728), .ZN(n8032) );
  NOR2_X1 U10298 ( .A1(n11632), .A2(n11503), .ZN(n9740) );
  OR2_X1 U10299 ( .A1(n8029), .A2(n8028), .ZN(n8030) );
  AND2_X1 U10300 ( .A1(n8031), .A2(n8030), .ZN(n9863) );
  AOI21_X1 U10301 ( .B1(n11432), .B2(n9740), .A(n9863), .ZN(n9729) );
  INV_X1 U10302 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14762) );
  NAND2_X1 U10303 ( .A1(n14733), .A2(n14762), .ZN(n8036) );
  OR2_X1 U10304 ( .A1(n11432), .A2(n8034), .ZN(n8035) );
  NAND2_X1 U10305 ( .A1(n13206), .A2(n14858), .ZN(n8039) );
  NOR2_X1 U10306 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n8041) );
  NOR2_X2 U10307 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .ZN(n8040) );
  INV_X2 U10308 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8232) );
  INV_X2 U10309 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8266) );
  INV_X2 U10310 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8311) );
  NOR2_X2 U10311 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n8043) );
  NOR2_X2 U10312 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n8042) );
  AND3_X2 U10313 ( .A1(n8043), .A2(n8042), .A3(n8144), .ZN(n8182) );
  NOR3_X1 U10314 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .A3(P1_IR_REG_23__SCAN_IN), .ZN(n8047) );
  NOR2_X1 U10315 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n8046) );
  NOR2_X1 U10316 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), 
        .ZN(n8045) );
  NOR2_X1 U10317 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), 
        .ZN(n8044) );
  INV_X1 U10318 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U10319 ( .A1(n8078), .A2(n8049), .ZN(n8051) );
  NAND2_X1 U10320 ( .A1(n8079), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8052) );
  INV_X1 U10321 ( .A(n8053), .ZN(n14079) );
  INV_X1 U10322 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n8055) );
  AND2_X2 U10323 ( .A1(n8056), .A2(n11844), .ZN(n8172) );
  NAND2_X1 U10324 ( .A1(n8172), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8062) );
  INV_X1 U10325 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8057) );
  OR2_X1 U10326 ( .A1(n8119), .A2(n8057), .ZN(n8061) );
  INV_X1 U10327 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n8059) );
  OR2_X1 U10328 ( .A1(n8492), .A2(n8059), .ZN(n8060) );
  INV_X1 U10329 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8066) );
  INV_X1 U10330 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8067) );
  NAND2_X1 U10331 ( .A1(n8069), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8068) );
  INV_X1 U10332 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n8072) );
  OR2_X1 U10333 ( .A1(n6461), .A2(n8072), .ZN(n8077) );
  INV_X1 U10334 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n13600) );
  OR2_X1 U10335 ( .A1(n8492), .A2(n13600), .ZN(n8076) );
  INV_X1 U10336 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n8073) );
  OR2_X1 U10337 ( .A1(n8119), .A2(n8073), .ZN(n8074) );
  INV_X1 U10338 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8081) );
  XNOR2_X2 U10339 ( .A(n8082), .B(n8081), .ZN(n8684) );
  NAND2_X4 U10340 ( .A1(n8685), .A2(n8684), .ZN(n9834) );
  NAND2_X2 U10341 ( .A1(n6463), .A2(n7433), .ZN(n8574) );
  NAND2_X1 U10342 ( .A1(n8147), .A2(n8083), .ZN(n8087) );
  NAND2_X1 U10343 ( .A1(n8125), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8086) );
  INV_X1 U10344 ( .A(n9834), .ZN(n8315) );
  NAND2_X1 U10345 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8084) );
  NAND2_X1 U10346 ( .A1(n8315), .A2(n13602), .ZN(n8085) );
  NAND2_X1 U10347 ( .A1(n14518), .A2(n10209), .ZN(n8090) );
  INV_X1 U10348 ( .A(SI_0_), .ZN(n9762) );
  INV_X1 U10349 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8811) );
  OAI21_X1 U10350 ( .B1(n6459), .B2(n9762), .A(n8811), .ZN(n8088) );
  AND2_X1 U10351 ( .A1(n8089), .A2(n8088), .ZN(n14091) );
  MUX2_X1 U10352 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14091), .S(n6463), .Z(n10396)
         );
  NAND2_X1 U10353 ( .A1(n8090), .A2(n10396), .ZN(n8091) );
  OAI211_X1 U10354 ( .C1(n14518), .C2(n10209), .A(n10403), .B(n8091), .ZN(
        n8115) );
  INV_X1 U10355 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8092) );
  NAND2_X1 U10356 ( .A1(n14090), .A2(n10945), .ZN(n8097) );
  INV_X1 U10357 ( .A(n8094), .ZN(n8095) );
  NAND2_X1 U10358 ( .A1(n8095), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8096) );
  MUX2_X1 U10359 ( .A(n8097), .B(n10041), .S(n13747), .Z(n8584) );
  XNOR2_X1 U10360 ( .A(n14090), .B(n13747), .ZN(n8098) );
  NAND2_X1 U10361 ( .A1(n8098), .A2(n14537), .ZN(n8099) );
  NAND2_X1 U10362 ( .A1(n14516), .A2(n10396), .ZN(n10404) );
  OAI21_X1 U10363 ( .B1(n10404), .B2(n8100), .A(n8252), .ZN(n8102) );
  AOI21_X1 U10364 ( .B1(n10404), .B2(n8100), .A(n14556), .ZN(n8101) );
  OAI22_X1 U10365 ( .A1(n8102), .A2(n8101), .B1(n6435), .B2(n8252), .ZN(n8114)
         );
  NAND2_X1 U10366 ( .A1(n8125), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8107) );
  INV_X1 U10367 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n8104) );
  INV_X1 U10368 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n8103) );
  NAND2_X1 U10369 ( .A1(n8126), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8105) );
  NAND2_X1 U10370 ( .A1(n8315), .A2(n13619), .ZN(n8106) );
  NAND2_X1 U10371 ( .A1(n8172), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8113) );
  INV_X1 U10372 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n13617) );
  OR2_X1 U10373 ( .A1(n8492), .A2(n13617), .ZN(n8112) );
  INV_X1 U10374 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n8108) );
  OR2_X1 U10375 ( .A1(n8119), .A2(n8108), .ZN(n8111) );
  INV_X1 U10376 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n8109) );
  OAI211_X1 U10377 ( .C1(n8115), .C2(n8252), .A(n8114), .B(n11330), .ZN(n8118)
         );
  MUX2_X1 U10378 ( .A(n10405), .B(n8116), .S(n8252), .Z(n8117) );
  NAND2_X1 U10379 ( .A1(n8118), .A2(n8117), .ZN(n8134) );
  NAND2_X1 U10380 ( .A1(n8590), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8124) );
  INV_X1 U10381 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9931) );
  INV_X1 U10382 ( .A(n8120), .ZN(n8123) );
  INV_X1 U10383 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n8121) );
  NAND2_X1 U10384 ( .A1(n8125), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8133) );
  INV_X1 U10385 ( .A(n8126), .ZN(n8128) );
  INV_X1 U10386 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8127) );
  NAND2_X1 U10387 ( .A1(n8128), .A2(n8127), .ZN(n8130) );
  NAND2_X1 U10388 ( .A1(n8130), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8129) );
  MUX2_X1 U10389 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8129), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n8131) );
  OR2_X1 U10390 ( .A1(n8130), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n8143) );
  NAND2_X1 U10391 ( .A1(n8315), .A2(n13631), .ZN(n8132) );
  INV_X2 U10392 ( .A(n13446), .ZN(n11079) );
  NAND2_X1 U10393 ( .A1(n13598), .A2(n11079), .ZN(n8135) );
  AND2_X1 U10394 ( .A1(n10706), .A2(n8135), .ZN(n10704) );
  NAND2_X1 U10395 ( .A1(n8493), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8141) );
  INV_X1 U10396 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n8137) );
  OR2_X1 U10397 ( .A1(n8157), .A2(n8137), .ZN(n8140) );
  XNOR2_X1 U10398 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n11315) );
  OR2_X1 U10399 ( .A1(n8492), .A2(n11315), .ZN(n8139) );
  INV_X1 U10400 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11316) );
  OR2_X1 U10401 ( .A1(n8577), .A2(n11316), .ZN(n8138) );
  AND4_X2 U10402 ( .A1(n8141), .A2(n8140), .A3(n8139), .A4(n8138), .ZN(n10709)
         );
  INV_X1 U10403 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9765) );
  NAND2_X1 U10404 ( .A1(n8143), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8145) );
  XNOR2_X1 U10405 ( .A(n8145), .B(n8144), .ZN(n13643) );
  OAI22_X1 U10406 ( .A1(n8392), .A2(n9765), .B1(n6463), .B2(n13643), .ZN(n8146) );
  INV_X1 U10407 ( .A(n8146), .ZN(n8149) );
  NAND2_X1 U10408 ( .A1(n8381), .A2(n9764), .ZN(n8148) );
  MUX2_X1 U10409 ( .A(n10709), .B(n14569), .S(n8252), .Z(n8151) );
  INV_X1 U10410 ( .A(n14569), .ZN(n11318) );
  MUX2_X1 U10411 ( .A(n11318), .B(n13597), .S(n8252), .Z(n8150) );
  INV_X1 U10412 ( .A(n8166), .ZN(n8164) );
  NAND2_X1 U10413 ( .A1(n9780), .A2(n8381), .ZN(n8155) );
  INV_X1 U10414 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9783) );
  OR2_X1 U10415 ( .A1(n8182), .A2(n8325), .ZN(n8152) );
  XNOR2_X1 U10416 ( .A(n8152), .B(n8181), .ZN(n9977) );
  OAI22_X1 U10417 ( .A1(n8392), .A2(n9783), .B1(n9834), .B2(n9977), .ZN(n8153)
         );
  INV_X1 U10418 ( .A(n8153), .ZN(n8154) );
  NAND2_X1 U10419 ( .A1(n8155), .A2(n8154), .ZN(n11170) );
  AOI21_X1 U10420 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8156) );
  NOR2_X1 U10421 ( .A1(n8156), .A2(n8173), .ZN(n11169) );
  INV_X1 U10422 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9934) );
  OR2_X1 U10423 ( .A1(n8462), .A2(n9934), .ZN(n8161) );
  INV_X1 U10424 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n8158) );
  OR2_X1 U10425 ( .A1(n8157), .A2(n8158), .ZN(n8160) );
  INV_X1 U10426 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9951) );
  OR2_X1 U10427 ( .A1(n8577), .A2(n9951), .ZN(n8159) );
  MUX2_X1 U10428 ( .A(n11170), .B(n13596), .S(n8252), .Z(n8165) );
  INV_X1 U10429 ( .A(n8165), .ZN(n8163) );
  NAND2_X1 U10430 ( .A1(n8164), .A2(n8163), .ZN(n8171) );
  NAND2_X1 U10431 ( .A1(n8166), .A2(n8165), .ZN(n8169) );
  MUX2_X1 U10432 ( .A(n13596), .B(n11170), .S(n8252), .Z(n8168) );
  NAND2_X1 U10433 ( .A1(n8169), .A2(n8168), .ZN(n8170) );
  NAND2_X1 U10434 ( .A1(n8591), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8180) );
  INV_X1 U10435 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9952) );
  OR2_X1 U10436 ( .A1(n8577), .A2(n9952), .ZN(n8179) );
  INV_X1 U10437 ( .A(n8192), .ZN(n8176) );
  INV_X1 U10438 ( .A(n8173), .ZN(n8174) );
  INV_X1 U10439 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n15125) );
  NAND2_X1 U10440 ( .A1(n8174), .A2(n15125), .ZN(n8175) );
  NAND2_X1 U10441 ( .A1(n8176), .A2(n8175), .ZN(n10860) );
  OR2_X1 U10442 ( .A1(n8589), .A2(n10860), .ZN(n8178) );
  INV_X1 U10443 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9935) );
  OR2_X1 U10444 ( .A1(n8462), .A2(n9935), .ZN(n8177) );
  NAND4_X1 U10445 ( .A1(n8180), .A2(n8179), .A3(n8178), .A4(n8177), .ZN(n13595) );
  NAND2_X1 U10446 ( .A1(n9785), .A2(n8381), .ZN(n8187) );
  NAND2_X1 U10447 ( .A1(n8182), .A2(n8181), .ZN(n8197) );
  NAND2_X1 U10448 ( .A1(n8197), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8184) );
  XNOR2_X1 U10449 ( .A(n8184), .B(n8183), .ZN(n13658) );
  OAI22_X1 U10450 ( .A1(n8392), .A2(n9786), .B1(n9834), .B2(n13658), .ZN(n8185) );
  INV_X1 U10451 ( .A(n8185), .ZN(n8186) );
  NAND2_X1 U10452 ( .A1(n8187), .A2(n8186), .ZN(n10857) );
  MUX2_X1 U10453 ( .A(n13595), .B(n10857), .S(n8252), .Z(n8189) );
  MUX2_X1 U10454 ( .A(n10857), .B(n13595), .S(n8252), .Z(n8188) );
  INV_X1 U10455 ( .A(n8189), .ZN(n8190) );
  NAND2_X1 U10456 ( .A1(n8493), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8196) );
  INV_X1 U10457 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n8191) );
  OR2_X1 U10458 ( .A1(n8157), .A2(n8191), .ZN(n8195) );
  OAI21_X1 U10459 ( .B1(n8192), .B2(P1_REG3_REG_7__SCAN_IN), .A(n8215), .ZN(
        n11109) );
  OR2_X1 U10460 ( .A1(n8589), .A2(n11109), .ZN(n8194) );
  INV_X1 U10461 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9953) );
  OR2_X1 U10462 ( .A1(n8577), .A2(n9953), .ZN(n8193) );
  NAND4_X1 U10463 ( .A1(n8196), .A2(n8195), .A3(n8194), .A4(n8193), .ZN(n13594) );
  NAND2_X1 U10464 ( .A1(n9789), .A2(n8381), .ZN(n8202) );
  NAND2_X1 U10465 ( .A1(n8209), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8199) );
  INV_X1 U10466 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8198) );
  XNOR2_X1 U10467 ( .A(n8199), .B(n8198), .ZN(n13671) );
  OAI22_X1 U10468 ( .A1(n8392), .A2(n9792), .B1(n9834), .B2(n13671), .ZN(n8200) );
  INV_X1 U10469 ( .A(n8200), .ZN(n8201) );
  NAND2_X1 U10470 ( .A1(n8202), .A2(n8201), .ZN(n11185) );
  MUX2_X1 U10471 ( .A(n13594), .B(n11185), .S(n8167), .Z(n8206) );
  MUX2_X1 U10472 ( .A(n13594), .B(n11185), .S(n8252), .Z(n8203) );
  AOI21_X1 U10473 ( .B1(n8207), .B2(n8206), .A(n8204), .ZN(n8205) );
  INV_X1 U10474 ( .A(n8205), .ZN(n8208) );
  NAND2_X1 U10475 ( .A1(n8208), .A2(n6532), .ZN(n8222) );
  NAND2_X1 U10476 ( .A1(n9836), .A2(n8381), .ZN(n8213) );
  NOR2_X1 U10477 ( .A1(n8209), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8233) );
  OR2_X1 U10478 ( .A1(n8233), .A2(n8325), .ZN(n8210) );
  XNOR2_X1 U10479 ( .A(n8210), .B(n8232), .ZN(n9965) );
  OAI22_X1 U10480 ( .A1(n8392), .A2(n9839), .B1(n9834), .B2(n9965), .ZN(n8211)
         );
  INV_X1 U10481 ( .A(n8211), .ZN(n8212) );
  NAND2_X1 U10482 ( .A1(n8213), .A2(n8212), .ZN(n14575) );
  NAND2_X1 U10483 ( .A1(n8591), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8220) );
  INV_X1 U10484 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9937) );
  OR2_X1 U10485 ( .A1(n8462), .A2(n9937), .ZN(n8219) );
  AND2_X1 U10486 ( .A1(n8215), .A2(n8214), .ZN(n8216) );
  OR2_X1 U10487 ( .A1(n8216), .A2(n8226), .ZN(n11357) );
  OR2_X1 U10488 ( .A1(n8589), .A2(n11357), .ZN(n8218) );
  INV_X1 U10489 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11358) );
  OR2_X1 U10490 ( .A1(n8577), .A2(n11358), .ZN(n8217) );
  NAND2_X1 U10491 ( .A1(n14575), .A2(n11407), .ZN(n8633) );
  OR2_X1 U10492 ( .A1(n14575), .A2(n11407), .ZN(n11190) );
  MUX2_X1 U10493 ( .A(n8633), .B(n11190), .S(n8252), .Z(n8221) );
  NAND2_X1 U10494 ( .A1(n8222), .A2(n8221), .ZN(n8225) );
  INV_X1 U10495 ( .A(n11407), .ZN(n13593) );
  MUX2_X1 U10496 ( .A(n13593), .B(n14575), .S(n8252), .Z(n8224) );
  NAND2_X1 U10497 ( .A1(n14575), .A2(n13593), .ZN(n8223) );
  NAND2_X1 U10498 ( .A1(n8591), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8231) );
  INV_X1 U10499 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9938) );
  OR2_X1 U10500 ( .A1(n8462), .A2(n9938), .ZN(n8230) );
  NAND2_X1 U10501 ( .A1(n8226), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8241) );
  OR2_X1 U10502 ( .A1(n8226), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8227) );
  NAND2_X1 U10503 ( .A1(n8241), .A2(n8227), .ZN(n11405) );
  OR2_X1 U10504 ( .A1(n8589), .A2(n11405), .ZN(n8229) );
  INV_X1 U10505 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9954) );
  OR2_X1 U10506 ( .A1(n8577), .A2(n9954), .ZN(n8228) );
  NAND2_X1 U10507 ( .A1(n9846), .A2(n8381), .ZN(n8236) );
  NAND2_X1 U10508 ( .A1(n8233), .A2(n8232), .ZN(n8268) );
  NAND2_X1 U10509 ( .A1(n8268), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8247) );
  XNOR2_X1 U10510 ( .A(n8247), .B(n8266), .ZN(n9989) );
  OAI22_X1 U10511 ( .A1(n8392), .A2(n9847), .B1(n9834), .B2(n9989), .ZN(n8234)
         );
  INV_X1 U10512 ( .A(n8234), .ZN(n8235) );
  MUX2_X1 U10513 ( .A(n11528), .B(n11535), .S(n8167), .Z(n8238) );
  INV_X1 U10514 ( .A(n11528), .ZN(n13592) );
  MUX2_X1 U10515 ( .A(n13592), .B(n11326), .S(n8252), .Z(n8237) );
  NAND2_X1 U10516 ( .A1(n8493), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8246) );
  INV_X1 U10517 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n8239) );
  OR2_X1 U10518 ( .A1(n8157), .A2(n8239), .ZN(n8245) );
  INV_X1 U10519 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8240) );
  NAND2_X1 U10520 ( .A1(n8241), .A2(n8240), .ZN(n8242) );
  NAND2_X1 U10521 ( .A1(n8259), .A2(n8242), .ZN(n14499) );
  OR2_X1 U10522 ( .A1(n8589), .A2(n14499), .ZN(n8244) );
  INV_X1 U10523 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9955) );
  OR2_X1 U10524 ( .A1(n8577), .A2(n9955), .ZN(n8243) );
  NAND4_X1 U10525 ( .A1(n8246), .A2(n8245), .A3(n8244), .A4(n8243), .ZN(n13591) );
  NAND2_X1 U10526 ( .A1(n8247), .A2(n8266), .ZN(n8248) );
  NAND2_X1 U10527 ( .A1(n8248), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8249) );
  INV_X1 U10528 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n8265) );
  XNOR2_X1 U10529 ( .A(n8249), .B(n8265), .ZN(n13688) );
  OAI22_X1 U10530 ( .A1(n8392), .A2(n9852), .B1(n9834), .B2(n13688), .ZN(n8250) );
  INV_X1 U10531 ( .A(n8250), .ZN(n8251) );
  MUX2_X1 U10532 ( .A(n13591), .B(n14502), .S(n8252), .Z(n8255) );
  MUX2_X1 U10533 ( .A(n13591), .B(n14502), .S(n8167), .Z(n8253) );
  NAND2_X1 U10534 ( .A1(n8254), .A2(n8253), .ZN(n8257) );
  NAND2_X1 U10535 ( .A1(n6553), .A2(n7322), .ZN(n8256) );
  NAND2_X1 U10536 ( .A1(n8591), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8264) );
  INV_X1 U10537 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10193) );
  OR2_X1 U10538 ( .A1(n8577), .A2(n10193), .ZN(n8263) );
  INV_X1 U10539 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8258) );
  NAND2_X1 U10540 ( .A1(n8259), .A2(n8258), .ZN(n8260) );
  NAND2_X1 U10541 ( .A1(n8278), .A2(n8260), .ZN(n14343) );
  OR2_X1 U10542 ( .A1(n8589), .A2(n14343), .ZN(n8262) );
  INV_X1 U10543 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10187) );
  OR2_X1 U10544 ( .A1(n8462), .A2(n10187), .ZN(n8261) );
  NAND4_X1 U10545 ( .A1(n8264), .A2(n8263), .A3(n8262), .A4(n8261), .ZN(n14506) );
  NAND2_X1 U10546 ( .A1(n9857), .A2(n8381), .ZN(n8273) );
  NAND2_X1 U10547 ( .A1(n8266), .A2(n8265), .ZN(n8267) );
  NAND2_X1 U10548 ( .A1(n8283), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8270) );
  XNOR2_X1 U10549 ( .A(n8270), .B(n8269), .ZN(n10192) );
  OAI22_X1 U10550 ( .A1(n8392), .A2(n9858), .B1(n9834), .B2(n10192), .ZN(n8271) );
  INV_X1 U10551 ( .A(n8271), .ZN(n8272) );
  MUX2_X1 U10552 ( .A(n14506), .B(n14373), .S(n8167), .Z(n8275) );
  MUX2_X1 U10553 ( .A(n14506), .B(n14373), .S(n8252), .Z(n8274) );
  INV_X1 U10554 ( .A(n8275), .ZN(n8276) );
  NAND2_X1 U10555 ( .A1(n8591), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8282) );
  INV_X1 U10556 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8277) );
  OR2_X1 U10557 ( .A1(n7379), .A2(n8296), .ZN(n11697) );
  OR2_X1 U10558 ( .A1(n8589), .A2(n11697), .ZN(n8281) );
  INV_X1 U10559 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n13711) );
  OR2_X1 U10560 ( .A1(n8577), .A2(n13711), .ZN(n8280) );
  INV_X1 U10561 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n13702) );
  OR2_X1 U10562 ( .A1(n8462), .A2(n13702), .ZN(n8279) );
  NAND4_X1 U10563 ( .A1(n8282), .A2(n8281), .A3(n8280), .A4(n8279), .ZN(n13590) );
  NAND2_X1 U10564 ( .A1(n9925), .A2(n8147), .ZN(n8286) );
  OAI21_X1 U10565 ( .B1(n8283), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8304) );
  XNOR2_X1 U10566 ( .A(n8304), .B(n8303), .ZN(n13710) );
  OAI22_X1 U10567 ( .A1(n8392), .A2(n9927), .B1(n9834), .B2(n13710), .ZN(n8284) );
  INV_X1 U10568 ( .A(n8284), .ZN(n8285) );
  MUX2_X1 U10569 ( .A(n13590), .B(n11693), .S(n8252), .Z(n8290) );
  NAND2_X1 U10570 ( .A1(n8289), .A2(n8290), .ZN(n8288) );
  MUX2_X1 U10571 ( .A(n13590), .B(n11693), .S(n8167), .Z(n8287) );
  NAND2_X1 U10572 ( .A1(n8288), .A2(n8287), .ZN(n8294) );
  INV_X1 U10573 ( .A(n8289), .ZN(n8292) );
  INV_X1 U10574 ( .A(n8290), .ZN(n8291) );
  NAND2_X1 U10575 ( .A1(n8292), .A2(n8291), .ZN(n8293) );
  NAND2_X1 U10576 ( .A1(n8493), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8302) );
  INV_X1 U10577 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8295) );
  OR2_X1 U10578 ( .A1(n8157), .A2(n8295), .ZN(n8301) );
  NAND2_X1 U10579 ( .A1(n8296), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8319) );
  OR2_X1 U10580 ( .A1(n8296), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8297) );
  NAND2_X1 U10581 ( .A1(n8319), .A2(n8297), .ZN(n14239) );
  OR2_X1 U10582 ( .A1(n8589), .A2(n14239), .ZN(n8300) );
  INV_X1 U10583 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n8298) );
  OR2_X1 U10584 ( .A1(n8577), .A2(n8298), .ZN(n8299) );
  NAND4_X1 U10585 ( .A1(n8302), .A2(n8301), .A3(n8300), .A4(n8299), .ZN(n13589) );
  NAND2_X1 U10586 ( .A1(n10075), .A2(n8381), .ZN(n8308) );
  NAND2_X1 U10587 ( .A1(n8304), .A2(n8303), .ZN(n8305) );
  NAND2_X1 U10588 ( .A1(n8305), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8312) );
  XNOR2_X1 U10589 ( .A(n8312), .B(n8311), .ZN(n14417) );
  OAI22_X1 U10590 ( .A1(n8392), .A2(n10076), .B1(n14417), .B2(n9834), .ZN(
        n8306) );
  INV_X1 U10591 ( .A(n8306), .ZN(n8307) );
  MUX2_X1 U10592 ( .A(n13589), .B(n14241), .S(n8167), .Z(n8310) );
  MUX2_X1 U10593 ( .A(n13589), .B(n14241), .S(n8252), .Z(n8309) );
  NAND2_X1 U10594 ( .A1(n10366), .A2(n8381), .ZN(n8317) );
  NAND2_X1 U10595 ( .A1(n8312), .A2(n8311), .ZN(n8313) );
  NAND2_X1 U10596 ( .A1(n8313), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8314) );
  XNOR2_X1 U10597 ( .A(n8314), .B(P1_IR_REG_14__SCAN_IN), .ZN(n13714) );
  AOI22_X1 U10598 ( .A1(n8315), .A2(n13714), .B1(n8125), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8316) );
  NAND2_X1 U10599 ( .A1(n8591), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8324) );
  INV_X1 U10600 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U10601 ( .A1(n8319), .A2(n8318), .ZN(n8320) );
  NAND2_X1 U10602 ( .A1(n8334), .A2(n8320), .ZN(n14338) );
  OR2_X1 U10603 ( .A1(n8589), .A2(n14338), .ZN(n8323) );
  INV_X1 U10604 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n13713) );
  OR2_X1 U10605 ( .A1(n8577), .A2(n13713), .ZN(n8322) );
  INV_X1 U10606 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n13700) );
  OR2_X1 U10607 ( .A1(n8462), .A2(n13700), .ZN(n8321) );
  NAND2_X1 U10608 ( .A1(n11762), .A2(n8340), .ZN(n11643) );
  NAND2_X1 U10609 ( .A1(n10452), .A2(n8381), .ZN(n8330) );
  INV_X1 U10610 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10453) );
  INV_X1 U10611 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8325) );
  XNOR2_X1 U10612 ( .A(n8327), .B(n8326), .ZN(n14437) );
  OAI22_X1 U10613 ( .A1(n8392), .A2(n10453), .B1(n9834), .B2(n14437), .ZN(
        n8328) );
  INV_X1 U10614 ( .A(n8328), .ZN(n8329) );
  NAND2_X1 U10615 ( .A1(n8493), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n8339) );
  INV_X1 U10616 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n8331) );
  OR2_X1 U10617 ( .A1(n8157), .A2(n8331), .ZN(n8338) );
  INV_X1 U10618 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8333) );
  NAND2_X1 U10619 ( .A1(n8334), .A2(n8333), .ZN(n8335) );
  NAND2_X1 U10620 ( .A1(n8348), .A2(n8335), .ZN(n13574) );
  OR2_X1 U10621 ( .A1(n8589), .A2(n13574), .ZN(n8337) );
  INV_X1 U10622 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11770) );
  OR2_X1 U10623 ( .A1(n8577), .A2(n11770), .ZN(n8336) );
  NAND2_X1 U10624 ( .A1(n14362), .A2(n14324), .ZN(n8631) );
  NAND2_X1 U10625 ( .A1(n8631), .A2(n8340), .ZN(n8342) );
  NAND2_X1 U10626 ( .A1(n11785), .A2(n11762), .ZN(n8341) );
  MUX2_X1 U10627 ( .A(n8342), .B(n8341), .S(n8167), .Z(n8343) );
  OR2_X1 U10628 ( .A1(n8344), .A2(n8343), .ZN(n8346) );
  MUX2_X1 U10629 ( .A(n8631), .B(n11785), .S(n8252), .Z(n8345) );
  INV_X1 U10630 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8347) );
  NAND2_X1 U10631 ( .A1(n8348), .A2(n8347), .ZN(n8349) );
  AND2_X1 U10632 ( .A1(n8377), .A2(n8349), .ZN(n13507) );
  NAND2_X1 U10633 ( .A1(n8525), .A2(n13507), .ZN(n8356) );
  INV_X1 U10634 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8350) );
  OR2_X1 U10635 ( .A1(n8462), .A2(n8350), .ZN(n8355) );
  INV_X1 U10636 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n8351) );
  OR2_X1 U10637 ( .A1(n8157), .A2(n8351), .ZN(n8354) );
  INV_X1 U10638 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n8352) );
  OR2_X1 U10639 ( .A1(n8577), .A2(n8352), .ZN(n8353) );
  NAND4_X1 U10640 ( .A1(n8356), .A2(n8355), .A3(n8354), .A4(n8353), .ZN(n13586) );
  NAND2_X1 U10641 ( .A1(n10361), .A2(n8381), .ZN(n8361) );
  OR2_X1 U10642 ( .A1(n8357), .A2(n8325), .ZN(n8358) );
  XNOR2_X1 U10643 ( .A(n8358), .B(P1_IR_REG_16__SCAN_IN), .ZN(n13717) );
  INV_X1 U10644 ( .A(n13717), .ZN(n14459) );
  OAI22_X1 U10645 ( .A1(n8392), .A2(n10365), .B1(n9834), .B2(n14459), .ZN(
        n8359) );
  INV_X1 U10646 ( .A(n8359), .ZN(n8360) );
  MUX2_X1 U10647 ( .A(n13586), .B(n13511), .S(n8167), .Z(n8363) );
  MUX2_X1 U10648 ( .A(n13586), .B(n13511), .S(n8252), .Z(n8362) );
  NAND2_X1 U10649 ( .A1(n10466), .A2(n8381), .ZN(n8370) );
  NAND2_X1 U10650 ( .A1(n8364), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8365) );
  MUX2_X1 U10651 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8365), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n8367) );
  AND2_X1 U10652 ( .A1(n8367), .A2(n8366), .ZN(n14473) );
  INV_X1 U10653 ( .A(n14473), .ZN(n10467) );
  OAI22_X1 U10654 ( .A1(n8392), .A2(n10468), .B1(n9834), .B2(n10467), .ZN(
        n8368) );
  INV_X1 U10655 ( .A(n8368), .ZN(n8369) );
  INV_X1 U10656 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n13957) );
  INV_X1 U10657 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n8371) );
  OR2_X1 U10658 ( .A1(n8157), .A2(n8371), .ZN(n8374) );
  INV_X1 U10659 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8372) );
  OR2_X1 U10660 ( .A1(n8462), .A2(n8372), .ZN(n8373) );
  AND2_X1 U10661 ( .A1(n8374), .A2(n8373), .ZN(n8380) );
  INV_X1 U10662 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8376) );
  NAND2_X1 U10663 ( .A1(n8377), .A2(n8376), .ZN(n8378) );
  NAND2_X1 U10664 ( .A1(n8397), .A2(n8378), .ZN(n13953) );
  OR2_X1 U10665 ( .A1(n13953), .A2(n8589), .ZN(n8379) );
  OAI211_X1 U10666 ( .C1(n8577), .C2(n13957), .A(n8380), .B(n8379), .ZN(n13928) );
  NAND2_X1 U10667 ( .A1(n14034), .A2(n13928), .ZN(n11873) );
  NAND2_X1 U10668 ( .A1(n10847), .A2(n8147), .ZN(n8384) );
  INV_X1 U10669 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10848) );
  OAI22_X1 U10670 ( .A1(n8392), .A2(n10848), .B1(n14536), .B2(n9834), .ZN(
        n8382) );
  INV_X1 U10671 ( .A(n8382), .ZN(n8383) );
  INV_X1 U10672 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8396) );
  XNOR2_X1 U10673 ( .A(n8417), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n13918) );
  NAND2_X1 U10674 ( .A1(n13918), .A2(n8525), .ZN(n8389) );
  INV_X1 U10675 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14027) );
  NAND2_X1 U10676 ( .A1(n8591), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8386) );
  NAND2_X1 U10677 ( .A1(n8590), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8385) );
  OAI211_X1 U10678 ( .C1(n8462), .C2(n14027), .A(n8386), .B(n8385), .ZN(n8387)
         );
  INV_X1 U10679 ( .A(n8387), .ZN(n8388) );
  OR2_X1 U10680 ( .A1(n13917), .A2(n13553), .ZN(n8406) );
  NAND2_X1 U10681 ( .A1(n13917), .A2(n13553), .ZN(n11855) );
  NAND2_X1 U10682 ( .A1(n10755), .A2(n8381), .ZN(n8395) );
  INV_X1 U10683 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10756) );
  NAND2_X1 U10684 ( .A1(n8366), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8391) );
  INV_X1 U10685 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8390) );
  XNOR2_X1 U10686 ( .A(n8391), .B(n8390), .ZN(n14477) );
  OAI22_X1 U10687 ( .A1(n8392), .A2(n10756), .B1(n9834), .B2(n14477), .ZN(
        n8393) );
  INV_X1 U10688 ( .A(n8393), .ZN(n8394) );
  NAND2_X1 U10689 ( .A1(n8397), .A2(n8396), .ZN(n8398) );
  NAND2_X1 U10690 ( .A1(n8417), .A2(n8398), .ZN(n13937) );
  AOI22_X1 U10691 ( .A1(n8493), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n8591), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n8400) );
  INV_X1 U10692 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14480) );
  OR2_X1 U10693 ( .A1(n8577), .A2(n14480), .ZN(n8399) );
  OAI211_X1 U10694 ( .C1(n13937), .C2(n8589), .A(n8400), .B(n8399), .ZN(n13912) );
  XNOR2_X1 U10695 ( .A(n13936), .B(n13912), .ZN(n13926) );
  NOR2_X1 U10696 ( .A1(n14034), .A2(n13928), .ZN(n11872) );
  MUX2_X1 U10697 ( .A(n13928), .B(n14034), .S(n8252), .Z(n8401) );
  AOI21_X1 U10698 ( .B1(n8402), .B2(n11872), .A(n8401), .ZN(n8411) );
  INV_X1 U10699 ( .A(n13912), .ZN(n13948) );
  OR3_X1 U10700 ( .A1(n13936), .A2(n13948), .A3(n8252), .ZN(n8405) );
  NAND3_X1 U10701 ( .A1(n13936), .A2(n13948), .A3(n8252), .ZN(n8404) );
  AND2_X1 U10702 ( .A1(n8405), .A2(n8404), .ZN(n8408) );
  MUX2_X1 U10703 ( .A(n11855), .B(n8406), .S(n8167), .Z(n8407) );
  OAI21_X1 U10704 ( .B1(n13909), .B2(n8408), .A(n8407), .ZN(n8409) );
  INV_X1 U10705 ( .A(n8409), .ZN(n8410) );
  AND2_X1 U10706 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n8413) );
  INV_X1 U10707 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8416) );
  INV_X1 U10708 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8415) );
  OAI21_X1 U10709 ( .B1(n8417), .B2(n8416), .A(n8415), .ZN(n8418) );
  NAND2_X1 U10710 ( .A1(n8430), .A2(n8418), .ZN(n13896) );
  OR2_X1 U10711 ( .A1(n13896), .A2(n8589), .ZN(n8421) );
  AOI22_X1 U10712 ( .A1(n8591), .A2(P1_REG0_REG_20__SCAN_IN), .B1(n8590), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n8420) );
  NAND2_X1 U10713 ( .A1(n8493), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8419) );
  NAND2_X1 U10714 ( .A1(n10866), .A2(n8381), .ZN(n8423) );
  NAND2_X1 U10715 ( .A1(n8125), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8422) );
  MUX2_X1 U10716 ( .A(n13488), .B(n14019), .S(n8167), .Z(n8425) );
  MUX2_X1 U10717 ( .A(n13913), .B(n13902), .S(n8252), .Z(n8424) );
  OAI21_X1 U10718 ( .B1(n8426), .B2(n8425), .A(n8424), .ZN(n8428) );
  NAND2_X1 U10719 ( .A1(n8426), .A2(n8425), .ZN(n8427) );
  NAND2_X1 U10720 ( .A1(n8428), .A2(n8427), .ZN(n8441) );
  INV_X1 U10721 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n15112) );
  NAND2_X1 U10722 ( .A1(n8430), .A2(n15112), .ZN(n8431) );
  NAND2_X1 U10723 ( .A1(n8447), .A2(n8431), .ZN(n13486) );
  OR2_X1 U10724 ( .A1(n13486), .A2(n8589), .ZN(n8436) );
  INV_X1 U10725 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n14017) );
  NAND2_X1 U10726 ( .A1(n8591), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8433) );
  NAND2_X1 U10727 ( .A1(n8590), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8432) );
  OAI211_X1 U10728 ( .C1(n8462), .C2(n14017), .A(n8433), .B(n8432), .ZN(n8434)
         );
  INV_X1 U10729 ( .A(n8434), .ZN(n8435) );
  NAND2_X1 U10730 ( .A1(n8436), .A2(n8435), .ZN(n13585) );
  NAND2_X1 U10731 ( .A1(n10944), .A2(n8381), .ZN(n8438) );
  NAND2_X1 U10732 ( .A1(n8125), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8437) );
  MUX2_X1 U10733 ( .A(n13585), .B(n13879), .S(n8252), .Z(n8442) );
  NAND2_X1 U10734 ( .A1(n8441), .A2(n8442), .ZN(n8440) );
  MUX2_X1 U10735 ( .A(n13585), .B(n13879), .S(n8167), .Z(n8439) );
  NAND2_X1 U10736 ( .A1(n8440), .A2(n8439), .ZN(n8446) );
  INV_X1 U10737 ( .A(n8441), .ZN(n8444) );
  INV_X1 U10738 ( .A(n8442), .ZN(n8443) );
  NAND2_X1 U10739 ( .A1(n8444), .A2(n8443), .ZN(n8445) );
  INV_X1 U10740 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13543) );
  NAND2_X1 U10741 ( .A1(n8447), .A2(n13543), .ZN(n8448) );
  NAND2_X1 U10742 ( .A1(n8478), .A2(n8448), .ZN(n13857) );
  OR2_X1 U10743 ( .A1(n13857), .A2(n8589), .ZN(n8454) );
  INV_X1 U10744 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8451) );
  NAND2_X1 U10745 ( .A1(n8590), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8450) );
  NAND2_X1 U10746 ( .A1(n8591), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8449) );
  OAI211_X1 U10747 ( .C1(n8462), .C2(n8451), .A(n8450), .B(n8449), .ZN(n8452)
         );
  INV_X1 U10748 ( .A(n8452), .ZN(n8453) );
  NAND2_X1 U10749 ( .A1(n8454), .A2(n8453), .ZN(n13487) );
  NAND2_X1 U10750 ( .A1(n8455), .A2(n7433), .ZN(n8456) );
  XNOR2_X1 U10751 ( .A(n8456), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14089) );
  MUX2_X1 U10752 ( .A(n13487), .B(n13863), .S(n8167), .Z(n8458) );
  MUX2_X1 U10753 ( .A(n13487), .B(n13863), .S(n8252), .Z(n8457) );
  XNOR2_X1 U10754 ( .A(n8478), .B(P1_REG3_REG_23__SCAN_IN), .ZN(n13843) );
  NAND2_X1 U10755 ( .A1(n13843), .A2(n8525), .ZN(n8465) );
  INV_X1 U10756 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n8461) );
  NAND2_X1 U10757 ( .A1(n8591), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8460) );
  NAND2_X1 U10758 ( .A1(n8590), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8459) );
  OAI211_X1 U10759 ( .C1(n8462), .C2(n8461), .A(n8460), .B(n8459), .ZN(n8463)
         );
  INV_X1 U10760 ( .A(n8463), .ZN(n8464) );
  NAND2_X1 U10761 ( .A1(n8465), .A2(n8464), .ZN(n13856) );
  NAND2_X1 U10762 ( .A1(n11343), .A2(n8381), .ZN(n8467) );
  NAND2_X1 U10763 ( .A1(n8125), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8466) );
  MUX2_X1 U10764 ( .A(n13856), .B(n14001), .S(n8252), .Z(n8471) );
  NAND2_X1 U10765 ( .A1(n8470), .A2(n8471), .ZN(n8469) );
  MUX2_X1 U10766 ( .A(n13856), .B(n14001), .S(n8167), .Z(n8468) );
  NAND2_X1 U10767 ( .A1(n8469), .A2(n8468), .ZN(n8475) );
  INV_X1 U10768 ( .A(n8470), .ZN(n8473) );
  INV_X1 U10769 ( .A(n8471), .ZN(n8472) );
  NAND2_X1 U10770 ( .A1(n8473), .A2(n8472), .ZN(n8474) );
  NAND2_X1 U10771 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n8476) );
  INV_X1 U10772 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13438) );
  INV_X1 U10773 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8477) );
  OAI21_X1 U10774 ( .B1(n8478), .B2(n13438), .A(n8477), .ZN(n8479) );
  AND2_X1 U10775 ( .A1(n8490), .A2(n8479), .ZN(n13828) );
  NAND2_X1 U10776 ( .A1(n13828), .A2(n8525), .ZN(n8484) );
  INV_X1 U10777 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n15108) );
  NAND2_X1 U10778 ( .A1(n8591), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8481) );
  NAND2_X1 U10779 ( .A1(n8590), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8480) );
  OAI211_X1 U10780 ( .C1(n15108), .C2(n8462), .A(n8481), .B(n8480), .ZN(n8482)
         );
  INV_X1 U10781 ( .A(n8482), .ZN(n8483) );
  NAND2_X1 U10782 ( .A1(n8484), .A2(n8483), .ZN(n13584) );
  NAND2_X1 U10783 ( .A1(n11429), .A2(n8381), .ZN(n8486) );
  NAND2_X1 U10784 ( .A1(n8125), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8485) );
  MUX2_X1 U10785 ( .A(n13584), .B(n13827), .S(n8167), .Z(n8488) );
  MUX2_X1 U10786 ( .A(n13584), .B(n13827), .S(n8252), .Z(n8487) );
  INV_X1 U10787 ( .A(n8490), .ZN(n8489) );
  NAND2_X1 U10788 ( .A1(n8489), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8511) );
  INV_X1 U10789 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n15171) );
  NAND2_X1 U10790 ( .A1(n8490), .A2(n15171), .ZN(n8491) );
  NAND2_X1 U10791 ( .A1(n8511), .A2(n8491), .ZN(n13810) );
  OR2_X1 U10792 ( .A1(n13810), .A2(n8492), .ZN(n8498) );
  INV_X1 U10793 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n15135) );
  NAND2_X1 U10794 ( .A1(n8493), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8495) );
  NAND2_X1 U10795 ( .A1(n8590), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8494) );
  OAI211_X1 U10796 ( .C1(n8157), .C2(n15135), .A(n8495), .B(n8494), .ZN(n8496)
         );
  INV_X1 U10797 ( .A(n8496), .ZN(n8497) );
  NAND2_X1 U10798 ( .A1(n11500), .A2(n8381), .ZN(n8500) );
  NAND2_X1 U10799 ( .A1(n8125), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8499) );
  MUX2_X1 U10800 ( .A(n13819), .B(n13807), .S(n8252), .Z(n8504) );
  NAND2_X1 U10801 ( .A1(n8503), .A2(n8504), .ZN(n8502) );
  MUX2_X1 U10802 ( .A(n13819), .B(n13807), .S(n8167), .Z(n8501) );
  NAND2_X1 U10803 ( .A1(n8502), .A2(n8501), .ZN(n8508) );
  INV_X1 U10804 ( .A(n8503), .ZN(n8506) );
  INV_X1 U10805 ( .A(n8504), .ZN(n8505) );
  NAND2_X1 U10806 ( .A1(n8506), .A2(n8505), .ZN(n8507) );
  INV_X1 U10807 ( .A(n8511), .ZN(n8509) );
  NAND2_X1 U10808 ( .A1(n8509), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8523) );
  INV_X1 U10809 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8510) );
  NAND2_X1 U10810 ( .A1(n8511), .A2(n8510), .ZN(n8512) );
  NAND2_X1 U10811 ( .A1(n8523), .A2(n8512), .ZN(n13792) );
  OR2_X1 U10812 ( .A1(n13792), .A2(n8589), .ZN(n8517) );
  INV_X1 U10813 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n15113) );
  NAND2_X1 U10814 ( .A1(n8590), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8514) );
  NAND2_X1 U10815 ( .A1(n8591), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8513) );
  OAI211_X1 U10816 ( .C1(n8462), .C2(n15113), .A(n8514), .B(n8513), .ZN(n8515)
         );
  INV_X1 U10817 ( .A(n8515), .ZN(n8516) );
  NAND2_X1 U10818 ( .A1(n8125), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8518) );
  MUX2_X1 U10819 ( .A(n13583), .B(n13988), .S(n8167), .Z(n8521) );
  MUX2_X1 U10820 ( .A(n13583), .B(n13988), .S(n8252), .Z(n8520) );
  INV_X1 U10821 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8522) );
  NAND2_X1 U10822 ( .A1(n8523), .A2(n8522), .ZN(n8524) );
  NAND2_X1 U10823 ( .A1(n13425), .A2(n8525), .ZN(n8531) );
  INV_X1 U10824 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U10825 ( .A1(n8591), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8527) );
  NAND2_X1 U10826 ( .A1(n8590), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8526) );
  OAI211_X1 U10827 ( .C1(n8528), .C2(n8462), .A(n8527), .B(n8526), .ZN(n8529)
         );
  INV_X1 U10828 ( .A(n8529), .ZN(n8530) );
  NAND2_X1 U10829 ( .A1(n11845), .A2(n8381), .ZN(n8533) );
  NAND2_X1 U10830 ( .A1(n8125), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8532) );
  MUX2_X1 U10831 ( .A(n13755), .B(n14052), .S(n8167), .Z(n8537) );
  NAND2_X1 U10832 ( .A1(n8536), .A2(n8537), .ZN(n8535) );
  MUX2_X1 U10833 ( .A(n13755), .B(n14052), .S(n8252), .Z(n8534) );
  NAND2_X1 U10834 ( .A1(n8535), .A2(n8534), .ZN(n8541) );
  INV_X1 U10835 ( .A(n8536), .ZN(n8539) );
  INV_X1 U10836 ( .A(n8537), .ZN(n8538) );
  NAND2_X1 U10837 ( .A1(n8539), .A2(n8538), .ZN(n8540) );
  INV_X1 U10838 ( .A(n8544), .ZN(n8542) );
  NAND2_X1 U10839 ( .A1(n8542), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n13762) );
  INV_X1 U10840 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8543) );
  NAND2_X1 U10841 ( .A1(n8544), .A2(n8543), .ZN(n8545) );
  NAND2_X1 U10842 ( .A1(n13762), .A2(n8545), .ZN(n13469) );
  INV_X1 U10843 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U10844 ( .A1(n8590), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U10845 ( .A1(n8591), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8546) );
  OAI211_X1 U10846 ( .C1(n8462), .C2(n8548), .A(n8547), .B(n8546), .ZN(n8549)
         );
  INV_X1 U10847 ( .A(n8549), .ZN(n8550) );
  INV_X1 U10848 ( .A(SI_27_), .ZN(n11596) );
  INV_X1 U10849 ( .A(n8552), .ZN(n8553) );
  INV_X1 U10850 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11917) );
  INV_X1 U10851 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13310) );
  MUX2_X1 U10852 ( .A(n11917), .B(n13310), .S(n6459), .Z(n8558) );
  INV_X1 U10853 ( .A(SI_28_), .ZN(n12764) );
  NAND2_X1 U10854 ( .A1(n8558), .A2(n12764), .ZN(n8566) );
  INV_X1 U10855 ( .A(n8558), .ZN(n8559) );
  NAND2_X1 U10856 ( .A1(n8559), .A2(SI_28_), .ZN(n8560) );
  NAND2_X1 U10857 ( .A1(n8566), .A2(n8560), .ZN(n8564) );
  NAND2_X1 U10858 ( .A1(n8125), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8561) );
  MUX2_X1 U10859 ( .A(n13759), .B(n13980), .S(n8167), .Z(n8602) );
  MUX2_X1 U10860 ( .A(n13759), .B(n13980), .S(n8252), .Z(n8563) );
  INV_X1 U10861 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14086) );
  INV_X1 U10862 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13304) );
  MUX2_X1 U10863 ( .A(n14086), .B(n13304), .S(n6459), .Z(n8567) );
  XNOR2_X1 U10864 ( .A(n8567), .B(SI_29_), .ZN(n8597) );
  INV_X1 U10865 ( .A(SI_29_), .ZN(n12762) );
  NAND2_X1 U10866 ( .A1(n8567), .A2(n12762), .ZN(n8568) );
  NAND2_X1 U10867 ( .A1(n8569), .A2(n8568), .ZN(n8572) );
  MUX2_X1 U10868 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6458), .Z(n8570) );
  NAND2_X1 U10869 ( .A1(n8570), .A2(SI_30_), .ZN(n8616) );
  OAI21_X1 U10870 ( .B1(n8570), .B2(SI_30_), .A(n8616), .ZN(n8571) );
  NAND2_X1 U10871 ( .A1(n8572), .A2(n8571), .ZN(n8573) );
  NAND2_X1 U10872 ( .A1(n8125), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8575) );
  INV_X1 U10873 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n15085) );
  NOR2_X1 U10874 ( .A1(n8462), .A2(n15085), .ZN(n8580) );
  INV_X1 U10875 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n13731) );
  NOR2_X1 U10876 ( .A1(n8577), .A2(n13731), .ZN(n8579) );
  INV_X1 U10877 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14039) );
  NOR2_X1 U10878 ( .A1(n8157), .A2(n14039), .ZN(n8578) );
  OR3_X1 U10879 ( .A1(n8580), .A2(n8579), .A3(n8578), .ZN(n13734) );
  NAND2_X1 U10880 ( .A1(n8252), .A2(n13734), .ZN(n8585) );
  INV_X1 U10881 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n13968) );
  NAND2_X1 U10882 ( .A1(n8590), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8582) );
  NAND2_X1 U10883 ( .A1(n8591), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8581) );
  OAI211_X1 U10884 ( .C1(n8462), .C2(n13968), .A(n8582), .B(n8581), .ZN(n13745) );
  INV_X1 U10885 ( .A(n13745), .ZN(n8583) );
  AOI21_X1 U10886 ( .B1(n8585), .B2(n8584), .A(n8583), .ZN(n8586) );
  AOI21_X1 U10887 ( .B1(n13740), .B2(n8167), .A(n8586), .ZN(n8609) );
  OAI21_X1 U10888 ( .B1(n13734), .B2(n10867), .A(n13745), .ZN(n8587) );
  INV_X1 U10889 ( .A(n8587), .ZN(n8588) );
  MUX2_X1 U10890 ( .A(n8588), .B(n13740), .S(n8252), .Z(n8607) );
  OR2_X1 U10891 ( .A1(n13762), .A2(n8589), .ZN(n8596) );
  INV_X1 U10892 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n13977) );
  NAND2_X1 U10893 ( .A1(n8590), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8593) );
  NAND2_X1 U10894 ( .A1(n8591), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8592) );
  OAI211_X1 U10895 ( .C1(n8462), .C2(n13977), .A(n8593), .B(n8592), .ZN(n8594)
         );
  INV_X1 U10896 ( .A(n8594), .ZN(n8595) );
  NAND2_X1 U10897 ( .A1(n9470), .A2(n8381), .ZN(n8600) );
  NAND2_X1 U10898 ( .A1(n8125), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8599) );
  MUX2_X1 U10899 ( .A(n8629), .B(n13970), .S(n8167), .Z(n8604) );
  INV_X1 U10900 ( .A(n8629), .ZN(n13582) );
  MUX2_X1 U10901 ( .A(n13582), .B(n13764), .S(n8252), .Z(n8603) );
  AOI22_X1 U10902 ( .A1(n8609), .A2(n8607), .B1(n8604), .B2(n8603), .ZN(n8601)
         );
  INV_X1 U10903 ( .A(n8603), .ZN(n8606) );
  INV_X1 U10904 ( .A(n8604), .ZN(n8605) );
  NAND2_X1 U10905 ( .A1(n8606), .A2(n8605), .ZN(n8608) );
  NAND2_X1 U10906 ( .A1(n8609), .A2(n8608), .ZN(n8613) );
  INV_X1 U10907 ( .A(n8607), .ZN(n8612) );
  INV_X1 U10908 ( .A(n8608), .ZN(n8611) );
  INV_X1 U10909 ( .A(n8609), .ZN(n8610) );
  AOI22_X1 U10910 ( .A1(n8613), .A2(n8612), .B1(n8611), .B2(n8610), .ZN(n8614)
         );
  NAND2_X1 U10911 ( .A1(n8615), .A2(n8614), .ZN(n8655) );
  MUX2_X1 U10912 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6459), .Z(n8618) );
  XNOR2_X1 U10913 ( .A(n8618), .B(SI_31_), .ZN(n8619) );
  NAND2_X1 U10914 ( .A1(n13295), .A2(n8147), .ZN(n8622) );
  NAND2_X1 U10915 ( .A1(n8125), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8621) );
  NAND2_X1 U10916 ( .A1(n13736), .A2(n8252), .ZN(n8664) );
  NOR2_X1 U10917 ( .A1(n13736), .A2(n8252), .ZN(n8656) );
  INV_X1 U10918 ( .A(n10209), .ZN(n8623) );
  NAND2_X1 U10919 ( .A1(n8623), .A2(n13747), .ZN(n8627) );
  NAND2_X1 U10920 ( .A1(n8624), .A2(n10867), .ZN(n8625) );
  NAND2_X1 U10921 ( .A1(n14534), .A2(n8625), .ZN(n8626) );
  NAND2_X1 U10922 ( .A1(n8627), .A2(n8626), .ZN(n8660) );
  NAND2_X1 U10923 ( .A1(n10945), .A2(n14537), .ZN(n8658) );
  NAND2_X1 U10924 ( .A1(n8660), .A2(n8658), .ZN(n8661) );
  AOI21_X1 U10925 ( .B1(n8656), .B2(n13734), .A(n8661), .ZN(n8628) );
  OAI21_X1 U10926 ( .B1(n13734), .B2(n8664), .A(n8628), .ZN(n8652) );
  XOR2_X1 U10927 ( .A(n13734), .B(n13736), .Z(n8653) );
  XNOR2_X1 U10928 ( .A(n13764), .B(n8629), .ZN(n13757) );
  XOR2_X1 U10929 ( .A(n13745), .B(n13740), .Z(n8648) );
  NAND2_X1 U10930 ( .A1(n13980), .A2(n13759), .ZN(n13756) );
  INV_X1 U10931 ( .A(n13584), .ZN(n13500) );
  XNOR2_X1 U10932 ( .A(n13827), .B(n13500), .ZN(n11878) );
  INV_X1 U10933 ( .A(n13856), .ZN(n11861) );
  XNOR2_X1 U10934 ( .A(n14001), .B(n11861), .ZN(n11860) );
  INV_X1 U10935 ( .A(n13487), .ZN(n15190) );
  XNOR2_X1 U10936 ( .A(n14064), .B(n15190), .ZN(n11858) );
  INV_X1 U10937 ( .A(n13926), .ZN(n13924) );
  NAND2_X1 U10938 ( .A1(n11785), .A2(n8631), .ZN(n11758) );
  INV_X1 U10939 ( .A(n11643), .ZN(n11642) );
  INV_X1 U10940 ( .A(n13589), .ZN(n14327) );
  XNOR2_X1 U10941 ( .A(n14241), .B(n14327), .ZN(n14243) );
  INV_X1 U10942 ( .A(n13591), .ZN(n11181) );
  OR2_X1 U10943 ( .A1(n14502), .A2(n11181), .ZN(n11538) );
  NAND2_X1 U10944 ( .A1(n14502), .A2(n11181), .ZN(n8632) );
  INV_X1 U10945 ( .A(n13594), .ZN(n11184) );
  XNOR2_X1 U10946 ( .A(n11185), .B(n11184), .ZN(n11174) );
  XNOR2_X1 U10947 ( .A(n14518), .B(n14535), .ZN(n14553) );
  INV_X1 U10948 ( .A(n11330), .ZN(n11334) );
  NAND2_X1 U10949 ( .A1(n10403), .A2(n6457), .ZN(n10397) );
  NOR4_X1 U10950 ( .A1(n14553), .A2(n10696), .A3(n11334), .A4(n10397), .ZN(
        n8634) );
  XNOR2_X1 U10951 ( .A(n10857), .B(n13595), .ZN(n10833) );
  XNOR2_X1 U10952 ( .A(n13596), .B(n11170), .ZN(n10712) );
  NAND4_X1 U10953 ( .A1(n8634), .A2(n10833), .A3(n10712), .A4(n10708), .ZN(
        n8635) );
  NOR4_X1 U10954 ( .A1(n14504), .A2(n11174), .A3(n11351), .A4(n8635), .ZN(
        n8636) );
  XNOR2_X1 U10955 ( .A(n11326), .B(n13592), .ZN(n11180) );
  NAND2_X1 U10956 ( .A1(n8636), .A2(n11180), .ZN(n8639) );
  INV_X1 U10957 ( .A(n14506), .ZN(n11539) );
  XNOR2_X1 U10958 ( .A(n14373), .B(n11539), .ZN(n14346) );
  INV_X1 U10959 ( .A(n13590), .ZN(n8637) );
  NAND2_X1 U10960 ( .A1(n11693), .A2(n8637), .ZN(n8638) );
  NAND2_X1 U10961 ( .A1(n14233), .A2(n8638), .ZN(n11637) );
  NOR4_X1 U10962 ( .A1(n14243), .A2(n8639), .A3(n14346), .A4(n11637), .ZN(
        n8641) );
  INV_X1 U10963 ( .A(n11872), .ZN(n8640) );
  NAND2_X1 U10964 ( .A1(n8640), .A2(n11873), .ZN(n13943) );
  XNOR2_X1 U10965 ( .A(n13511), .B(n13586), .ZN(n11850) );
  NAND4_X1 U10966 ( .A1(n11642), .A2(n8641), .A3(n13943), .A4(n11850), .ZN(
        n8642) );
  NOR4_X1 U10967 ( .A1(n13909), .A2(n13924), .A3(n11758), .A4(n8642), .ZN(
        n8643) );
  XNOR2_X1 U10968 ( .A(n13902), .B(n13913), .ZN(n13888) );
  XNOR2_X1 U10969 ( .A(n13879), .B(n13585), .ZN(n13870) );
  NAND4_X1 U10970 ( .A1(n11858), .A2(n8643), .A3(n13888), .A4(n13870), .ZN(
        n8644) );
  NOR4_X1 U10971 ( .A1(n11865), .A2(n11878), .A3(n11860), .A4(n8644), .ZN(
        n8646) );
  NAND4_X1 U10972 ( .A1(n13770), .A2(n8646), .A3(n13749), .A4(n13789), .ZN(
        n8647) );
  NOR4_X1 U10973 ( .A1(n8653), .A2(n13757), .A3(n8648), .A4(n8647), .ZN(n8649)
         );
  XNOR2_X1 U10974 ( .A(n8649), .B(n13747), .ZN(n8650) );
  OAI21_X1 U10975 ( .B1(n8655), .B2(n8652), .A(n8651), .ZN(n8675) );
  NOR2_X1 U10976 ( .A1(n8653), .A2(n8660), .ZN(n8654) );
  NAND2_X1 U10977 ( .A1(n8655), .A2(n8654), .ZN(n8668) );
  INV_X1 U10978 ( .A(n8656), .ZN(n8657) );
  XNOR2_X1 U10979 ( .A(n8657), .B(n8660), .ZN(n8659) );
  INV_X1 U10980 ( .A(n13736), .ZN(n14041) );
  NAND4_X1 U10981 ( .A1(n8659), .A2(n14041), .A3(n13734), .A4(n8658), .ZN(
        n8667) );
  OR3_X1 U10982 ( .A1(n8664), .A2(n13734), .A3(n8660), .ZN(n8666) );
  INV_X1 U10983 ( .A(n13734), .ZN(n8663) );
  INV_X1 U10984 ( .A(n8661), .ZN(n8662) );
  NAND4_X1 U10985 ( .A1(n8664), .A2(n8663), .A3(n8662), .A4(n13736), .ZN(n8665) );
  NAND2_X1 U10986 ( .A1(n8668), .A2(n7375), .ZN(n8674) );
  OAI21_X1 U10987 ( .B1(n8669), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8671) );
  INV_X1 U10988 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8670) );
  XNOR2_X1 U10989 ( .A(n8671), .B(n8670), .ZN(n9832) );
  INV_X1 U10990 ( .A(n9832), .ZN(n8672) );
  NAND2_X1 U10991 ( .A1(n8672), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11344) );
  INV_X1 U10992 ( .A(n11344), .ZN(n8673) );
  OAI21_X1 U10993 ( .B1(n8675), .B2(n8674), .A(n8673), .ZN(n8688) );
  INV_X1 U10994 ( .A(n14534), .ZN(n9833) );
  NAND2_X1 U10995 ( .A1(n10867), .A2(n14536), .ZN(n8683) );
  NAND2_X1 U10996 ( .A1(n8676), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8677) );
  MUX2_X1 U10997 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8677), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n8678) );
  NAND2_X1 U10998 ( .A1(n8678), .A2(n6521), .ZN(n11501) );
  NAND2_X1 U10999 ( .A1(n6508), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8679) );
  MUX2_X1 U11000 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8679), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n8680) );
  NAND2_X1 U11001 ( .A1(n8680), .A2(n8676), .ZN(n11430) );
  NOR2_X1 U11002 ( .A1(n11501), .A2(n11430), .ZN(n8682) );
  NAND2_X1 U11003 ( .A1(n6521), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8681) );
  XNOR2_X1 U11004 ( .A(n8681), .B(P1_IR_REG_26__SCAN_IN), .ZN(n11627) );
  AOI21_X1 U11005 ( .B1(n9833), .B2(n8683), .A(n10042), .ZN(n10607) );
  INV_X1 U11006 ( .A(n8684), .ZN(n9942) );
  INV_X1 U11007 ( .A(n8685), .ZN(n13613) );
  NAND3_X1 U11008 ( .A1(n10541), .A2(n9942), .A3(n13929), .ZN(n8686) );
  OAI211_X1 U11009 ( .C1(n14090), .C2(n11344), .A(n8686), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8687) );
  NAND2_X1 U11010 ( .A1(n8688), .A2(n8687), .ZN(P1_U3242) );
  AND2_X1 U11011 ( .A1(n8760), .A2(n8787), .ZN(n8699) );
  NAND2_X1 U11012 ( .A1(n9198), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8698) );
  OR2_X1 U11013 ( .A1(n8699), .A2(n8973), .ZN(n8700) );
  XNOR2_X1 U11014 ( .A(n8700), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12454) );
  NAND2_X1 U11015 ( .A1(n12302), .A2(n12454), .ZN(n9561) );
  NAND2_X1 U11016 ( .A1(n8701), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8702) );
  OR2_X1 U11017 ( .A1(n8703), .A2(n8973), .ZN(n8704) );
  XNOR2_X1 U11018 ( .A(n8704), .B(P3_IR_REG_20__SCAN_IN), .ZN(n9259) );
  NAND2_X1 U11019 ( .A1(n10145), .A2(n9259), .ZN(n12105) );
  INV_X1 U11020 ( .A(n8813), .ZN(n8706) );
  NAND2_X1 U11021 ( .A1(n8801), .A2(n8706), .ZN(n8708) );
  NAND2_X1 U11022 ( .A1(n9744), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8707) );
  XNOR2_X1 U11023 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8825) );
  NAND2_X1 U11024 ( .A1(n8826), .A2(n8825), .ZN(n8711) );
  NAND2_X1 U11025 ( .A1(n8709), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8710) );
  NAND2_X1 U11026 ( .A1(n8839), .A2(n8838), .ZN(n8714) );
  NAND2_X1 U11027 ( .A1(n8857), .A2(n8856), .ZN(n8716) );
  NAND2_X1 U11028 ( .A1(n8869), .A2(n8868), .ZN(n8718) );
  NAND2_X1 U11029 ( .A1(n9781), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8717) );
  NOR2_X1 U11030 ( .A1(n9786), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8719) );
  NAND2_X1 U11031 ( .A1(n9786), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8720) );
  NAND2_X1 U11032 ( .A1(n9839), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8722) );
  XNOR2_X1 U11033 ( .A(n9847), .B(P1_DATAO_REG_9__SCAN_IN), .ZN(n8924) );
  INV_X1 U11034 ( .A(n8924), .ZN(n8724) );
  NAND2_X1 U11035 ( .A1(n9847), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8725) );
  XNOR2_X1 U11036 ( .A(n9852), .B(P1_DATAO_REG_10__SCAN_IN), .ZN(n8941) );
  INV_X1 U11037 ( .A(n8941), .ZN(n8727) );
  NAND2_X1 U11038 ( .A1(n9852), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8728) );
  NAND2_X1 U11039 ( .A1(n9861), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U11040 ( .A1(n9927), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8733) );
  NAND2_X1 U11041 ( .A1(n9926), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8732) );
  NAND2_X1 U11042 ( .A1(n8733), .A2(n8732), .ZN(n8964) );
  NAND2_X1 U11043 ( .A1(n8988), .A2(n8735), .ZN(n9004) );
  NAND2_X1 U11044 ( .A1(n10367), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8737) );
  NAND2_X1 U11045 ( .A1(n10369), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8736) );
  AND2_X1 U11046 ( .A1(n8737), .A2(n8736), .ZN(n9003) );
  NAND2_X1 U11047 ( .A1(n10453), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8741) );
  NAND2_X1 U11048 ( .A1(n10455), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8739) );
  NAND2_X1 U11049 ( .A1(n8741), .A2(n8739), .ZN(n9018) );
  INV_X1 U11050 ( .A(n9018), .ZN(n8740) );
  NAND2_X1 U11051 ( .A1(n10365), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U11052 ( .A1(n10363), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U11053 ( .A1(n8745), .A2(n8743), .ZN(n9030) );
  INV_X1 U11054 ( .A(n9030), .ZN(n8744) );
  NAND2_X1 U11055 ( .A1(n10468), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8748) );
  NAND2_X1 U11056 ( .A1(n10471), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8746) );
  NAND2_X1 U11057 ( .A1(n8748), .A2(n8746), .ZN(n9045) );
  INV_X1 U11058 ( .A(n9045), .ZN(n8747) );
  NAND2_X1 U11059 ( .A1(n10756), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8750) );
  NAND2_X1 U11060 ( .A1(n10758), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8749) );
  AND2_X1 U11061 ( .A1(n8750), .A2(n8749), .ZN(n8782) );
  NAND2_X1 U11062 ( .A1(n10848), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U11063 ( .A1(n10850), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8751) );
  AND2_X1 U11064 ( .A1(n8752), .A2(n8751), .ZN(n9059) );
  INV_X1 U11065 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10946) );
  NAND2_X1 U11066 ( .A1(n10946), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9086) );
  INV_X1 U11067 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10949) );
  NAND2_X1 U11068 ( .A1(n10949), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8754) );
  NAND2_X1 U11069 ( .A1(n9086), .A2(n8754), .ZN(n9083) );
  XNOR2_X1 U11070 ( .A(n9085), .B(n9083), .ZN(n10748) );
  NOR2_X1 U11071 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_22__SCAN_IN), 
        .ZN(n8758) );
  NOR2_X1 U11072 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n8757) );
  INV_X1 U11073 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8763) );
  NAND2_X2 U11074 ( .A1(n8829), .A2(n7433), .ZN(n8968) );
  NAND2_X1 U11075 ( .A1(n10748), .A2(n12083), .ZN(n8768) );
  NAND2_X2 U11076 ( .A1(n8829), .A2(n6459), .ZN(n9155) );
  INV_X2 U11077 ( .A(n9007), .ZN(n12086) );
  INV_X1 U11078 ( .A(SI_21_), .ZN(n10749) );
  OR2_X1 U11079 ( .A1(n12086), .A2(n10749), .ZN(n8767) );
  NAND2_X1 U11080 ( .A1(n8862), .A2(n8861), .ZN(n8876) );
  OR2_X1 U11081 ( .A1(n8876), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8888) );
  NOR2_X1 U11082 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_REG3_REG_9__SCAN_IN), 
        .ZN(n8769) );
  INV_X1 U11083 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n9010) );
  INV_X1 U11084 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n11679) );
  INV_X1 U11085 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n9036) );
  INV_X1 U11086 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n9065) );
  INV_X1 U11087 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n9075) );
  NAND2_X1 U11088 ( .A1(n9078), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8770) );
  NAND2_X1 U11089 ( .A1(n9091), .A2(n8770), .ZN(n12556) );
  NOR2_X2 U11090 ( .A1(n8771), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n8775) );
  NAND2_X1 U11091 ( .A1(n8775), .A2(n8772), .ZN(n12753) );
  INV_X1 U11092 ( .A(n11907), .ZN(n8777) );
  AND2_X2 U11093 ( .A1(n8777), .A2(n8778), .ZN(n8819) );
  INV_X2 U11094 ( .A(n8832), .ZN(n9162) );
  NAND2_X1 U11095 ( .A1(n12556), .A2(n9162), .ZN(n8781) );
  AOI22_X1 U11096 ( .A1(n6443), .A2(P3_REG1_REG_21__SCAN_IN), .B1(n12089), 
        .B2(P3_REG0_REG_21__SCAN_IN), .ZN(n8780) );
  BUF_X4 U11097 ( .A(n6460), .Z(n12091) );
  NAND2_X1 U11098 ( .A1(n12091), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8779) );
  OR2_X1 U11099 ( .A1(n8783), .A2(n8782), .ZN(n8784) );
  NAND2_X1 U11100 ( .A1(n8785), .A2(n8784), .ZN(n10094) );
  INV_X1 U11101 ( .A(n8760), .ZN(n8786) );
  NAND2_X1 U11102 ( .A1(n8786), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8788) );
  XNOR2_X1 U11103 ( .A(n8788), .B(n8787), .ZN(n12452) );
  INV_X1 U11104 ( .A(n12452), .ZN(n12427) );
  AOI22_X1 U11105 ( .A1(n9007), .A2(SI_18_), .B1(n9193), .B2(n12427), .ZN(
        n8789) );
  INV_X1 U11106 ( .A(n12726), .ZN(n9058) );
  INV_X1 U11107 ( .A(n9066), .ZN(n8792) );
  NAND2_X1 U11108 ( .A1(n9053), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8791) );
  NAND2_X1 U11109 ( .A1(n8792), .A2(n8791), .ZN(n12587) );
  AOI22_X1 U11110 ( .A1(n12587), .A2(n9162), .B1(n12091), .B2(
        P3_REG2_REG_18__SCAN_IN), .ZN(n8794) );
  AOI22_X1 U11111 ( .A1(n6444), .A2(P3_REG1_REG_18__SCAN_IN), .B1(n12089), 
        .B2(P3_REG0_REG_18__SCAN_IN), .ZN(n8793) );
  NAND2_X1 U11112 ( .A1(n8795), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8797) );
  NAND2_X1 U11113 ( .A1(n8806), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8796) );
  AND2_X1 U11114 ( .A1(n8797), .A2(n8796), .ZN(n8800) );
  NAND2_X1 U11115 ( .A1(n8833), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8799) );
  NAND2_X1 U11116 ( .A1(n8819), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8798) );
  NAND3_X2 U11117 ( .A1(n8800), .A2(n8799), .A3(n8798), .ZN(n12332) );
  INV_X1 U11118 ( .A(n12332), .ZN(n8816) );
  XNOR2_X1 U11119 ( .A(n8801), .B(n8813), .ZN(n9759) );
  OR2_X1 U11120 ( .A1(n8968), .A2(n9759), .ZN(n8805) );
  INV_X1 U11121 ( .A(n10274), .ZN(n8803) );
  NAND2_X1 U11122 ( .A1(n8819), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8810) );
  NAND2_X1 U11123 ( .A1(n8795), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8809) );
  NAND2_X1 U11124 ( .A1(n6460), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8808) );
  NAND2_X1 U11125 ( .A1(n8833), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8807) );
  NAND4_X1 U11126 ( .A1(n8810), .A2(n8809), .A3(n8808), .A4(n8807), .ZN(n12334) );
  OR2_X1 U11127 ( .A1(n9155), .A2(n9762), .ZN(n8815) );
  NAND2_X1 U11128 ( .A1(n8811), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8812) );
  AND2_X1 U11129 ( .A1(n8813), .A2(n8812), .ZN(n9763) );
  OR2_X1 U11130 ( .A1(n8968), .A2(n9763), .ZN(n8814) );
  OAI211_X1 U11131 ( .C1(n10204), .C2(n8829), .A(n8815), .B(n8814), .ZN(n10252) );
  NAND2_X1 U11132 ( .A1(n10236), .A2(n14947), .ZN(n8818) );
  NAND2_X1 U11133 ( .A1(n8816), .A2(n8817), .ZN(n10148) );
  NAND2_X1 U11134 ( .A1(n8818), .A2(n10148), .ZN(n14937) );
  NAND2_X1 U11135 ( .A1(n8819), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8823) );
  NAND2_X1 U11136 ( .A1(n6442), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8822) );
  NAND2_X1 U11137 ( .A1(n6460), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8821) );
  NAND2_X1 U11138 ( .A1(n8833), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8820) );
  INV_X1 U11139 ( .A(n6448), .ZN(n10359) );
  XNOR2_X1 U11140 ( .A(n8826), .B(n8825), .ZN(n9776) );
  OR2_X1 U11141 ( .A1(n8968), .A2(n9776), .ZN(n8828) );
  OR2_X1 U11142 ( .A1(n9155), .A2(SI_2_), .ZN(n8827) );
  OAI211_X1 U11143 ( .C1(n10359), .C2(n8829), .A(n8828), .B(n8827), .ZN(n14943) );
  XNOR2_X1 U11144 ( .A(n12331), .B(n14943), .ZN(n12116) );
  NAND2_X1 U11145 ( .A1(n14937), .A2(n12116), .ZN(n8831) );
  INV_X1 U11146 ( .A(n12331), .ZN(n10161) );
  NAND2_X1 U11147 ( .A1(n10161), .A2(n14943), .ZN(n8830) );
  INV_X1 U11148 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10486) );
  NAND2_X1 U11149 ( .A1(n8819), .A2(n10486), .ZN(n8837) );
  NAND2_X1 U11150 ( .A1(n6443), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8836) );
  NAND2_X1 U11151 ( .A1(n6460), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8835) );
  NAND2_X1 U11152 ( .A1(n8833), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8834) );
  OR2_X1 U11153 ( .A1(n9155), .A2(SI_3_), .ZN(n8843) );
  XNOR2_X1 U11154 ( .A(n8839), .B(n8838), .ZN(n9778) );
  OR2_X1 U11155 ( .A1(n8968), .A2(n9778), .ZN(n8842) );
  NAND2_X1 U11156 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6530), .ZN(n8840) );
  OR2_X1 U11157 ( .A1(n8829), .A2(n10317), .ZN(n8841) );
  NAND2_X1 U11158 ( .A1(n10499), .A2(n14976), .ZN(n12153) );
  INV_X1 U11159 ( .A(n14976), .ZN(n8844) );
  NAND2_X1 U11160 ( .A1(n8845), .A2(n14976), .ZN(n8846) );
  NAND2_X1 U11161 ( .A1(n12089), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8850) );
  NAND2_X1 U11162 ( .A1(n6437), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8849) );
  OR2_X1 U11163 ( .A1(n7381), .A2(n8862), .ZN(n10503) );
  NAND2_X1 U11164 ( .A1(n9162), .A2(n10503), .ZN(n8848) );
  NAND2_X1 U11165 ( .A1(n12091), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8847) );
  NAND4_X1 U11166 ( .A1(n8850), .A2(n8849), .A3(n8848), .A4(n8847), .ZN(n12330) );
  NOR2_X1 U11167 ( .A1(n8851), .A2(n8973), .ZN(n8852) );
  MUX2_X1 U11168 ( .A(n8973), .B(n8852), .S(P3_IR_REG_4__SCAN_IN), .Z(n8853)
         );
  INV_X1 U11169 ( .A(n8853), .ZN(n8855) );
  NAND2_X1 U11170 ( .A1(n8851), .A2(n8854), .ZN(n8882) );
  NAND2_X1 U11171 ( .A1(n8855), .A2(n8882), .ZN(n10321) );
  INV_X1 U11172 ( .A(n10321), .ZN(n10450) );
  XNOR2_X1 U11173 ( .A(n8857), .B(n8856), .ZN(n9772) );
  OR2_X1 U11174 ( .A1(n8968), .A2(n9772), .ZN(n8859) );
  OR2_X1 U11175 ( .A1(n12086), .A2(SI_4_), .ZN(n8858) );
  OAI211_X1 U11176 ( .C1(n10450), .C2(n8829), .A(n8859), .B(n8858), .ZN(n12156) );
  NAND2_X1 U11177 ( .A1(n10802), .A2(n12115), .ZN(n10801) );
  INV_X1 U11178 ( .A(n12156), .ZN(n14984) );
  NAND2_X1 U11179 ( .A1(n12330), .A2(n14984), .ZN(n8860) );
  NAND2_X1 U11180 ( .A1(n12089), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8867) );
  NAND2_X1 U11181 ( .A1(n12090), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8866) );
  OR2_X1 U11182 ( .A1(n8862), .A2(n8861), .ZN(n8863) );
  NAND2_X1 U11183 ( .A1(n8876), .A2(n8863), .ZN(n12012) );
  NAND2_X1 U11184 ( .A1(n9162), .A2(n12012), .ZN(n8865) );
  NAND2_X1 U11185 ( .A1(n12091), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8864) );
  OR2_X1 U11186 ( .A1(n9155), .A2(SI_5_), .ZN(n8873) );
  XNOR2_X1 U11187 ( .A(n8869), .B(n8868), .ZN(n9774) );
  OR2_X1 U11188 ( .A1(n8968), .A2(n9774), .ZN(n8872) );
  NAND2_X1 U11189 ( .A1(n8882), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8870) );
  OR2_X1 U11190 ( .A1(n8829), .A2(n10385), .ZN(n8871) );
  NAND2_X1 U11191 ( .A1(n10902), .A2(n12011), .ZN(n12165) );
  INV_X1 U11192 ( .A(n10902), .ZN(n12329) );
  INV_X1 U11193 ( .A(n12011), .ZN(n14990) );
  NAND2_X1 U11194 ( .A1(n12329), .A2(n14990), .ZN(n12164) );
  NAND2_X1 U11195 ( .A1(n10902), .A2(n14990), .ZN(n8875) );
  NAND2_X1 U11196 ( .A1(n12089), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8881) );
  NAND2_X1 U11197 ( .A1(n6444), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8880) );
  NAND2_X1 U11198 ( .A1(n8876), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8877) );
  NAND2_X1 U11199 ( .A1(n8888), .A2(n8877), .ZN(n10901) );
  NAND2_X1 U11200 ( .A1(n9162), .A2(n10901), .ZN(n8879) );
  NAND2_X1 U11201 ( .A1(n12091), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8878) );
  NAND2_X1 U11202 ( .A1(n8896), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8883) );
  XNOR2_X1 U11203 ( .A(n8883), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10325) );
  INV_X1 U11204 ( .A(n10325), .ZN(n10334) );
  INV_X1 U11205 ( .A(SI_6_), .ZN(n9760) );
  OR2_X1 U11206 ( .A1(n9155), .A2(n9760), .ZN(n8887) );
  XNOR2_X1 U11207 ( .A(n9788), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8884) );
  XNOR2_X1 U11208 ( .A(n8885), .B(n8884), .ZN(n9761) );
  OR2_X1 U11209 ( .A1(n8968), .A2(n9761), .ZN(n8886) );
  OAI211_X1 U11210 ( .C1(n8829), .C2(n10334), .A(n8887), .B(n8886), .ZN(n10905) );
  NAND2_X1 U11211 ( .A1(n10933), .A2(n10905), .ZN(n12168) );
  INV_X1 U11212 ( .A(n10933), .ZN(n12328) );
  INV_X1 U11213 ( .A(n10905), .ZN(n14995) );
  NAND2_X1 U11214 ( .A1(n12328), .A2(n14995), .ZN(n12169) );
  NAND2_X1 U11215 ( .A1(n12168), .A2(n12169), .ZN(n12112) );
  NAND2_X1 U11216 ( .A1(n12089), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8893) );
  NAND2_X1 U11217 ( .A1(n6444), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8892) );
  AND2_X1 U11218 ( .A1(n8888), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8889) );
  OR2_X1 U11219 ( .A1(n8889), .A2(n8918), .ZN(n11018) );
  NAND2_X1 U11220 ( .A1(n9162), .A2(n11018), .ZN(n8891) );
  NAND2_X1 U11221 ( .A1(n12091), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8890) );
  XNOR2_X1 U11222 ( .A(n8895), .B(n8894), .ZN(n9770) );
  OR2_X1 U11223 ( .A1(n8968), .A2(n9770), .ZN(n8900) );
  OR2_X1 U11224 ( .A1(n12086), .A2(SI_7_), .ZN(n8899) );
  OR2_X1 U11225 ( .A1(n8906), .A2(n8973), .ZN(n8897) );
  OR2_X1 U11226 ( .A1(n8829), .A2(n10645), .ZN(n8898) );
  NAND2_X1 U11227 ( .A1(n11117), .A2(n8914), .ZN(n12174) );
  INV_X1 U11228 ( .A(n11117), .ZN(n12327) );
  INV_X1 U11229 ( .A(n8914), .ZN(n15002) );
  NAND2_X1 U11230 ( .A1(n12327), .A2(n15002), .ZN(n12175) );
  NAND2_X1 U11231 ( .A1(n12174), .A2(n12175), .ZN(n11014) );
  NAND2_X1 U11232 ( .A1(n11013), .A2(n11014), .ZN(n11012) );
  NAND2_X1 U11233 ( .A1(n12089), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8904) );
  NAND2_X1 U11234 ( .A1(n12090), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8903) );
  INV_X1 U11235 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10651) );
  XNOR2_X1 U11236 ( .A(n8918), .B(n10651), .ZN(n11120) );
  NAND2_X1 U11237 ( .A1(n9162), .A2(n11120), .ZN(n8902) );
  NAND2_X1 U11238 ( .A1(n12091), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8901) );
  INV_X1 U11239 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8905) );
  NAND2_X1 U11240 ( .A1(n8906), .A2(n8905), .ZN(n8908) );
  NAND2_X1 U11241 ( .A1(n8908), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8907) );
  MUX2_X1 U11242 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8907), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n8909) );
  NAND2_X1 U11243 ( .A1(n8909), .A2(n8928), .ZN(n10762) );
  XNOR2_X1 U11244 ( .A(n8911), .B(n8910), .ZN(n9756) );
  OR2_X1 U11245 ( .A1(n8968), .A2(n9756), .ZN(n8913) );
  INV_X1 U11246 ( .A(SI_8_), .ZN(n9757) );
  OR2_X1 U11247 ( .A1(n12086), .A2(n9757), .ZN(n8912) );
  OAI211_X1 U11248 ( .C1(n8829), .C2(n10762), .A(n8913), .B(n8912), .ZN(n15009) );
  NAND2_X1 U11249 ( .A1(n10935), .A2(n15009), .ZN(n12179) );
  INV_X1 U11250 ( .A(n10935), .ZN(n12326) );
  INV_X1 U11251 ( .A(n15009), .ZN(n8916) );
  NAND2_X1 U11252 ( .A1(n12326), .A2(n8916), .ZN(n12180) );
  NAND2_X1 U11253 ( .A1(n12179), .A2(n12180), .ZN(n9245) );
  NAND2_X1 U11254 ( .A1(n12327), .A2(n8914), .ZN(n11054) );
  AND2_X1 U11255 ( .A1(n9245), .A2(n11054), .ZN(n8915) );
  NAND2_X1 U11256 ( .A1(n11012), .A2(n8915), .ZN(n11056) );
  NAND2_X1 U11257 ( .A1(n10935), .A2(n8916), .ZN(n8917) );
  NAND2_X1 U11258 ( .A1(n12090), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8923) );
  NAND2_X1 U11259 ( .A1(n12089), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8922) );
  INV_X1 U11260 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n10926) );
  AOI21_X1 U11261 ( .B1(n8918), .B2(n10651), .A(n10926), .ZN(n8919) );
  OR2_X1 U11262 ( .A1(n8935), .A2(n8919), .ZN(n11379) );
  NAND2_X1 U11263 ( .A1(n9162), .A2(n11379), .ZN(n8921) );
  NAND2_X1 U11264 ( .A1(n12091), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8920) );
  NAND4_X1 U11265 ( .A1(n8923), .A2(n8922), .A3(n8921), .A4(n8920), .ZN(n12325) );
  XNOR2_X1 U11266 ( .A(n8925), .B(n8924), .ZN(n14205) );
  OR2_X1 U11267 ( .A1(n8968), .A2(n14205), .ZN(n8932) );
  OR2_X1 U11268 ( .A1(n12086), .A2(SI_9_), .ZN(n8931) );
  NAND2_X1 U11269 ( .A1(n8928), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8927) );
  MUX2_X1 U11270 ( .A(n8927), .B(P3_IR_REG_31__SCAN_IN), .S(n8926), .Z(n8929)
         );
  OR2_X1 U11271 ( .A1(n8829), .A2(n10957), .ZN(n8930) );
  NAND2_X1 U11272 ( .A1(n12325), .A2(n15015), .ZN(n12135) );
  OAI21_X1 U11273 ( .B1(n12325), .B2(n15015), .A(n12135), .ZN(n12182) );
  OR2_X1 U11274 ( .A1(n8935), .A2(n8934), .ZN(n8936) );
  AND2_X1 U11275 ( .A1(n8949), .A2(n8936), .ZN(n14894) );
  INV_X1 U11276 ( .A(n14894), .ZN(n11418) );
  NAND2_X1 U11277 ( .A1(n9162), .A2(n11418), .ZN(n8940) );
  NAND2_X1 U11278 ( .A1(n12090), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8939) );
  NAND2_X1 U11279 ( .A1(n12091), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8938) );
  NAND2_X1 U11280 ( .A1(n12089), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8937) );
  XNOR2_X1 U11281 ( .A(n8942), .B(n8941), .ZN(n9768) );
  OR2_X1 U11282 ( .A1(n8968), .A2(n9768), .ZN(n8946) );
  OR2_X1 U11283 ( .A1(n9155), .A2(SI_10_), .ZN(n8945) );
  NAND2_X1 U11284 ( .A1(n8972), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8943) );
  INV_X1 U11285 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8970) );
  XNOR2_X1 U11286 ( .A(n8943), .B(n8970), .ZN(n12348) );
  INV_X1 U11287 ( .A(n12348), .ZN(n10965) );
  OR2_X1 U11288 ( .A1(n8829), .A2(n10965), .ZN(n8944) );
  NAND2_X1 U11289 ( .A1(n11385), .A2(n11384), .ZN(n9249) );
  NAND2_X1 U11290 ( .A1(n12324), .A2(n14888), .ZN(n12189) );
  NAND2_X1 U11291 ( .A1(n9249), .A2(n12189), .ZN(n12184) );
  NAND2_X1 U11292 ( .A1(n8947), .A2(n12184), .ZN(n11415) );
  NAND2_X1 U11293 ( .A1(n12324), .A2(n11384), .ZN(n8948) );
  NAND2_X1 U11294 ( .A1(n11415), .A2(n8948), .ZN(n11368) );
  NAND2_X1 U11295 ( .A1(n12090), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8954) );
  NAND2_X1 U11296 ( .A1(n12089), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8953) );
  NAND2_X1 U11297 ( .A1(n8949), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8950) );
  NAND2_X1 U11298 ( .A1(n8977), .A2(n8950), .ZN(n11391) );
  NAND2_X1 U11299 ( .A1(n9162), .A2(n11391), .ZN(n8952) );
  NAND2_X1 U11300 ( .A1(n12091), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8951) );
  OAI21_X1 U11301 ( .B1(n8972), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8955) );
  XNOR2_X1 U11302 ( .A(n8955), .B(P3_IR_REG_11__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U11303 ( .A1(n9007), .A2(n8956), .B1(n9193), .B2(n14899), .ZN(n8960) );
  XNOR2_X1 U11304 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8957) );
  XNOR2_X1 U11305 ( .A(n8958), .B(n8957), .ZN(n14208) );
  NAND2_X1 U11306 ( .A1(n14208), .A2(n12083), .ZN(n8959) );
  NAND2_X1 U11307 ( .A1(n8960), .A2(n8959), .ZN(n12187) );
  NAND2_X1 U11308 ( .A1(n11459), .A2(n12187), .ZN(n8961) );
  NAND2_X1 U11309 ( .A1(n11368), .A2(n8961), .ZN(n8963) );
  INV_X1 U11310 ( .A(n12187), .ZN(n14312) );
  NAND2_X1 U11311 ( .A1(n12323), .A2(n14312), .ZN(n8962) );
  NAND2_X1 U11312 ( .A1(n8963), .A2(n8962), .ZN(n11457) );
  NAND2_X1 U11313 ( .A1(n8965), .A2(n8964), .ZN(n8966) );
  NAND2_X1 U11314 ( .A1(n8967), .A2(n8966), .ZN(n9784) );
  OR2_X1 U11315 ( .A1(n9784), .A2(n8968), .ZN(n8976) );
  INV_X1 U11316 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8969) );
  NAND2_X1 U11317 ( .A1(n8970), .A2(n8969), .ZN(n8971) );
  NOR2_X1 U11318 ( .A1(n8972), .A2(n8971), .ZN(n8990) );
  OR2_X1 U11319 ( .A1(n8990), .A2(n8973), .ZN(n8974) );
  INV_X1 U11320 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8989) );
  XNOR2_X1 U11321 ( .A(n8974), .B(n8989), .ZN(n12383) );
  INV_X1 U11322 ( .A(n12383), .ZN(n12353) );
  AOI22_X1 U11323 ( .A1(n9007), .A2(SI_12_), .B1(n9193), .B2(n12353), .ZN(
        n8975) );
  NAND2_X1 U11324 ( .A1(n6444), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8982) );
  NAND2_X1 U11325 ( .A1(n12089), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8981) );
  NAND2_X1 U11326 ( .A1(n8977), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8978) );
  NAND2_X1 U11327 ( .A1(n8996), .A2(n8978), .ZN(n11463) );
  NAND2_X1 U11328 ( .A1(n9162), .A2(n11463), .ZN(n8980) );
  NAND2_X1 U11329 ( .A1(n12091), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8979) );
  NAND4_X1 U11330 ( .A1(n8982), .A2(n8981), .A3(n8980), .A4(n8979), .ZN(n12322) );
  NAND2_X1 U11331 ( .A1(n11462), .A2(n12322), .ZN(n12204) );
  INV_X1 U11332 ( .A(n12322), .ZN(n11506) );
  NAND2_X1 U11333 ( .A1(n11506), .A2(n14308), .ZN(n12201) );
  NAND2_X1 U11334 ( .A1(n12204), .A2(n12201), .ZN(n9250) );
  NAND2_X1 U11335 ( .A1(n11457), .A2(n9250), .ZN(n8984) );
  NAND2_X1 U11336 ( .A1(n14308), .A2(n12322), .ZN(n8983) );
  NAND2_X1 U11337 ( .A1(n8984), .A2(n8983), .ZN(n11585) );
  INV_X1 U11338 ( .A(n8985), .ZN(n8986) );
  NAND2_X1 U11339 ( .A1(n8986), .A2(n10078), .ZN(n8987) );
  NAND2_X1 U11340 ( .A1(n8988), .A2(n8987), .ZN(n9850) );
  NAND2_X1 U11341 ( .A1(n9850), .A2(n12083), .ZN(n8995) );
  NAND2_X1 U11342 ( .A1(n8990), .A2(n8989), .ZN(n8992) );
  NAND2_X1 U11343 ( .A1(n8992), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8991) );
  MUX2_X1 U11344 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8991), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n8993) );
  AOI22_X1 U11345 ( .A1(n9007), .A2(n15157), .B1(n9193), .B2(n14916), .ZN(
        n8994) );
  NAND2_X1 U11346 ( .A1(n8995), .A2(n8994), .ZN(n14303) );
  NAND2_X1 U11347 ( .A1(n6444), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9000) );
  NAND2_X1 U11348 ( .A1(n12089), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8999) );
  OR2_X1 U11349 ( .A1(n7386), .A2(n9011), .ZN(n11588) );
  NAND2_X1 U11350 ( .A1(n9162), .A2(n11588), .ZN(n8998) );
  NAND2_X1 U11351 ( .A1(n12091), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8997) );
  NAND4_X1 U11352 ( .A1(n9000), .A2(n8999), .A3(n8998), .A4(n8997), .ZN(n12321) );
  OR2_X1 U11353 ( .A1(n14303), .A2(n12321), .ZN(n12205) );
  NAND2_X1 U11354 ( .A1(n14303), .A2(n12321), .ZN(n12206) );
  NAND2_X1 U11355 ( .A1(n12205), .A2(n12206), .ZN(n12122) );
  NAND2_X1 U11356 ( .A1(n11585), .A2(n12122), .ZN(n9002) );
  INV_X1 U11357 ( .A(n12321), .ZN(n11675) );
  OR2_X1 U11358 ( .A1(n14303), .A2(n11675), .ZN(n9001) );
  NAND2_X1 U11359 ( .A1(n9002), .A2(n9001), .ZN(n11652) );
  XNOR2_X1 U11360 ( .A(n9004), .B(n9003), .ZN(n14216) );
  NAND2_X1 U11361 ( .A1(n14216), .A2(n12083), .ZN(n9009) );
  INV_X1 U11362 ( .A(SI_14_), .ZN(n14214) );
  NAND2_X1 U11363 ( .A1(n9020), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9006) );
  INV_X1 U11364 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9005) );
  XNOR2_X1 U11365 ( .A(n9006), .B(n9005), .ZN(n14219) );
  AOI22_X1 U11366 ( .A1(n9007), .A2(n14214), .B1(n9193), .B2(n14219), .ZN(
        n9008) );
  NAND2_X1 U11367 ( .A1(n6444), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9016) );
  NAND2_X1 U11368 ( .A1(n12089), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9015) );
  NAND2_X1 U11369 ( .A1(n12091), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9014) );
  NOR2_X1 U11370 ( .A1(n9011), .A2(n9010), .ZN(n9012) );
  OR2_X1 U11371 ( .A1(n9024), .A2(n9012), .ZN(n11655) );
  NAND2_X1 U11372 ( .A1(n9162), .A2(n11655), .ZN(n9013) );
  NAND4_X1 U11373 ( .A1(n9016), .A2(n9015), .A3(n9014), .A4(n9013), .ZN(n12320) );
  OR2_X1 U11374 ( .A1(n14298), .A2(n12320), .ZN(n9252) );
  NAND2_X1 U11375 ( .A1(n14298), .A2(n12320), .ZN(n12210) );
  NAND2_X1 U11376 ( .A1(n9252), .A2(n12210), .ZN(n12121) );
  INV_X1 U11377 ( .A(n12320), .ZN(n11678) );
  OR2_X1 U11378 ( .A1(n14298), .A2(n11678), .ZN(n9017) );
  XNOR2_X1 U11379 ( .A(n9019), .B(n9018), .ZN(n14220) );
  NAND2_X1 U11380 ( .A1(n14220), .A2(n12083), .ZN(n9023) );
  OAI21_X1 U11381 ( .B1(n9020), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9021) );
  XNOR2_X1 U11382 ( .A(n9021), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12412) );
  AOI22_X1 U11383 ( .A1(n9007), .A2(SI_15_), .B1(n9193), .B2(n12412), .ZN(
        n9022) );
  NOR2_X1 U11384 ( .A1(n9024), .A2(n11679), .ZN(n9025) );
  OR2_X1 U11385 ( .A1(n9037), .A2(n9025), .ZN(n12617) );
  NAND2_X1 U11386 ( .A1(n9162), .A2(n12617), .ZN(n9029) );
  NAND2_X1 U11387 ( .A1(n6444), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U11388 ( .A1(n12091), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n9027) );
  NAND2_X1 U11389 ( .A1(n12089), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9026) );
  NAND2_X1 U11390 ( .A1(n12745), .A2(n11778), .ZN(n12217) );
  INV_X1 U11391 ( .A(n11778), .ZN(n12319) );
  XNOR2_X1 U11392 ( .A(n9031), .B(n9030), .ZN(n14224) );
  NAND2_X1 U11393 ( .A1(n14224), .A2(n12083), .ZN(n9035) );
  NAND2_X1 U11394 ( .A1(n9032), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9033) );
  XNOR2_X1 U11395 ( .A(n9033), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U11396 ( .A1(n9007), .A2(SI_16_), .B1(n9193), .B2(n12414), .ZN(
        n9034) );
  NAND2_X1 U11397 ( .A1(n6444), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n9042) );
  NAND2_X1 U11398 ( .A1(n12091), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n9041) );
  OR2_X1 U11399 ( .A1(n9037), .A2(n9036), .ZN(n9038) );
  NAND2_X1 U11400 ( .A1(n9051), .A2(n9038), .ZN(n12604) );
  NAND2_X1 U11401 ( .A1(n9162), .A2(n12604), .ZN(n9040) );
  NAND2_X1 U11402 ( .A1(n12089), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9039) );
  NAND4_X1 U11403 ( .A1(n9042), .A2(n9041), .A3(n9040), .A4(n9039), .ZN(n12318) );
  AND2_X1 U11404 ( .A1(n12738), .A2(n12318), .ZN(n9044) );
  OR2_X1 U11405 ( .A1(n12738), .A2(n12318), .ZN(n9043) );
  XNOR2_X1 U11406 ( .A(n9046), .B(n9045), .ZN(n10030) );
  NAND2_X1 U11407 ( .A1(n10030), .A2(n12083), .ZN(n9050) );
  NAND2_X1 U11408 ( .A1(n9047), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9048) );
  XNOR2_X1 U11409 ( .A(n9048), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12425) );
  AOI22_X1 U11410 ( .A1(n9007), .A2(SI_17_), .B1(n9193), .B2(n12425), .ZN(
        n9049) );
  NAND2_X1 U11411 ( .A1(n12089), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U11412 ( .A1(n6443), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9056) );
  NAND2_X1 U11413 ( .A1(n9051), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9052) );
  NAND2_X1 U11414 ( .A1(n9053), .A2(n9052), .ZN(n12599) );
  NAND2_X1 U11415 ( .A1(n9162), .A2(n12599), .ZN(n9055) );
  NAND2_X1 U11416 ( .A1(n12091), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n9054) );
  OR2_X1 U11417 ( .A1(n12600), .A2(n12056), .ZN(n12229) );
  NAND2_X1 U11418 ( .A1(n12600), .A2(n12056), .ZN(n12233) );
  INV_X1 U11419 ( .A(n12600), .ZN(n12731) );
  NOR2_X1 U11420 ( .A1(n12731), .A2(n12056), .ZN(n12582) );
  NAND2_X1 U11421 ( .A1(n12726), .A2(n12020), .ZN(n12231) );
  OR2_X1 U11422 ( .A1(n9060), .A2(n9059), .ZN(n9061) );
  NAND2_X1 U11423 ( .A1(n9062), .A2(n9061), .ZN(n10114) );
  NAND2_X1 U11424 ( .A1(n10114), .A2(n12083), .ZN(n9064) );
  AOI22_X1 U11425 ( .A1(n9007), .A2(n10113), .B1(n9193), .B2(n12459), .ZN(
        n9063) );
  XNOR2_X1 U11426 ( .A(n9066), .B(n9065), .ZN(n12575) );
  NAND2_X1 U11427 ( .A1(n12575), .A2(n9162), .ZN(n9071) );
  NAND2_X1 U11428 ( .A1(n12089), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9068) );
  NAND2_X1 U11429 ( .A1(n6443), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9067) );
  AND2_X1 U11430 ( .A1(n9068), .A2(n9067), .ZN(n9070) );
  NAND2_X1 U11431 ( .A1(n12091), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n9069) );
  XNOR2_X1 U11432 ( .A(n9072), .B(n10868), .ZN(n10534) );
  NAND2_X1 U11433 ( .A1(n10534), .A2(n12083), .ZN(n9074) );
  OR2_X1 U11434 ( .A1(n12086), .A2(n10535), .ZN(n9073) );
  OR2_X1 U11435 ( .A1(n9076), .A2(n9075), .ZN(n9077) );
  NAND2_X1 U11436 ( .A1(n9078), .A2(n9077), .ZN(n12567) );
  NAND2_X1 U11437 ( .A1(n12567), .A2(n9162), .ZN(n9081) );
  AOI22_X1 U11438 ( .A1(n6444), .A2(P3_REG1_REG_20__SCAN_IN), .B1(n12091), 
        .B2(P3_REG2_REG_20__SCAN_IN), .ZN(n9080) );
  NAND2_X1 U11439 ( .A1(n12089), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9079) );
  NAND2_X1 U11440 ( .A1(n12714), .A2(n11971), .ZN(n12244) );
  INV_X1 U11441 ( .A(n12714), .ZN(n9082) );
  NAND2_X1 U11442 ( .A1(n12557), .A2(n12047), .ZN(n9255) );
  NOR2_X1 U11443 ( .A1(n12550), .A2(n12551), .ZN(n12549) );
  INV_X1 U11444 ( .A(n9083), .ZN(n9084) );
  INV_X1 U11445 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9087) );
  XNOR2_X1 U11446 ( .A(n9087), .B(P1_DATAO_REG_22__SCAN_IN), .ZN(n9098) );
  XNOR2_X1 U11447 ( .A(n9099), .B(n9098), .ZN(n10783) );
  NAND2_X1 U11448 ( .A1(n10783), .A2(n12083), .ZN(n9090) );
  OR2_X1 U11449 ( .A1(n9155), .A2(n9088), .ZN(n9089) );
  NAND2_X1 U11450 ( .A1(n9091), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9092) );
  INV_X1 U11451 ( .A(n9103), .ZN(n9102) );
  NAND2_X1 U11452 ( .A1(n9092), .A2(n9102), .ZN(n12545) );
  NAND2_X1 U11453 ( .A1(n12545), .A2(n9162), .ZN(n9095) );
  AOI22_X1 U11454 ( .A1(n6444), .A2(P3_REG1_REG_22__SCAN_IN), .B1(n12089), 
        .B2(P3_REG0_REG_22__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U11455 ( .A1(n12091), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n9093) );
  NOR2_X1 U11456 ( .A1(n9096), .A2(n11964), .ZN(n9097) );
  OAI22_X2 U11457 ( .A1(n12541), .A2(n9097), .B1(n12313), .B2(n12703), .ZN(
        n12532) );
  INV_X1 U11458 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n15191) );
  XNOR2_X1 U11459 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n9112) );
  XNOR2_X1 U11460 ( .A(n9113), .B(n9112), .ZN(n10941) );
  NAND2_X1 U11461 ( .A1(n10941), .A2(n12083), .ZN(n9101) );
  OR2_X1 U11462 ( .A1(n9155), .A2(n10943), .ZN(n9100) );
  NAND2_X1 U11463 ( .A1(n12089), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U11464 ( .A1(n6443), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9107) );
  NAND2_X1 U11465 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(n9102), .ZN(n9104) );
  INV_X1 U11466 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n15082) );
  NAND2_X1 U11467 ( .A1(n9104), .A2(n9121), .ZN(n12536) );
  NAND2_X1 U11468 ( .A1(n9162), .A2(n12536), .ZN(n9106) );
  NAND2_X1 U11469 ( .A1(n6460), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9105) );
  NAND4_X1 U11470 ( .A1(n9108), .A2(n9107), .A3(n9106), .A4(n9105), .ZN(n12312) );
  NAND2_X1 U11471 ( .A1(n12697), .A2(n12312), .ZN(n9110) );
  OR2_X1 U11472 ( .A1(n12697), .A2(n12312), .ZN(n9109) );
  NAND2_X1 U11473 ( .A1(n9110), .A2(n9109), .ZN(n12531) );
  INV_X1 U11474 ( .A(n9110), .ZN(n9111) );
  INV_X1 U11475 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9114) );
  NAND2_X1 U11476 ( .A1(n9114), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9115) );
  INV_X1 U11477 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11435) );
  NAND2_X1 U11478 ( .A1(n9117), .A2(n11435), .ZN(n9118) );
  NAND2_X1 U11479 ( .A1(n9129), .A2(n9118), .ZN(n9128) );
  INV_X1 U11480 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11431) );
  XNOR2_X1 U11481 ( .A(n9128), .B(n11431), .ZN(n11303) );
  NAND2_X1 U11482 ( .A1(n11303), .A2(n12083), .ZN(n9120) );
  OR2_X1 U11483 ( .A1(n12086), .A2(n6793), .ZN(n9119) );
  NAND2_X1 U11484 ( .A1(n6444), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9126) );
  NAND2_X1 U11485 ( .A1(n12091), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9125) );
  NAND2_X1 U11486 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(n9121), .ZN(n9122) );
  NAND2_X1 U11487 ( .A1(n9122), .A2(n9133), .ZN(n12525) );
  NAND2_X1 U11488 ( .A1(n9162), .A2(n12525), .ZN(n9124) );
  NAND2_X1 U11489 ( .A1(n12089), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9123) );
  NAND4_X1 U11490 ( .A1(n9126), .A2(n9125), .A3(n9124), .A4(n9123), .ZN(n12311) );
  AOI22_X1 U11491 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n11505), .B2(n11502), .ZN(n9130) );
  XNOR2_X1 U11492 ( .A(n9139), .B(n9130), .ZN(n11496) );
  NAND2_X1 U11493 ( .A1(n11496), .A2(n12083), .ZN(n9132) );
  OR2_X1 U11494 ( .A1(n9155), .A2(n11498), .ZN(n9131) );
  NAND2_X1 U11495 ( .A1(n12089), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n9138) );
  NAND2_X1 U11496 ( .A1(n6444), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9137) );
  NAND2_X1 U11497 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(n9133), .ZN(n9134) );
  NAND2_X1 U11498 ( .A1(n9134), .A2(n9144), .ZN(n12515) );
  NAND2_X1 U11499 ( .A1(n9162), .A2(n12515), .ZN(n9136) );
  NAND2_X1 U11500 ( .A1(n6460), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9135) );
  NAND2_X1 U11501 ( .A1(n12516), .A2(n12032), .ZN(n12263) );
  AOI22_X1 U11502 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n11630), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n11629), .ZN(n9140) );
  INV_X1 U11503 ( .A(n9140), .ZN(n9141) );
  XNOR2_X1 U11504 ( .A(n9151), .B(n9141), .ZN(n11580) );
  NAND2_X1 U11505 ( .A1(n11580), .A2(n12083), .ZN(n9143) );
  OR2_X1 U11506 ( .A1(n12086), .A2(n11581), .ZN(n9142) );
  NAND2_X1 U11507 ( .A1(n12089), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9149) );
  NAND2_X1 U11508 ( .A1(n6443), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9148) );
  NAND2_X1 U11509 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(n9144), .ZN(n9145) );
  INV_X1 U11510 ( .A(n9158), .ZN(n9160) );
  NAND2_X1 U11511 ( .A1(n9145), .A2(n9160), .ZN(n12502) );
  NAND2_X1 U11512 ( .A1(n9162), .A2(n12502), .ZN(n9147) );
  NAND2_X1 U11513 ( .A1(n12091), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9146) );
  NAND2_X1 U11514 ( .A1(n12680), .A2(n11955), .ZN(n9150) );
  NAND2_X1 U11515 ( .A1(n11630), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9152) );
  AOI22_X1 U11516 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n13313), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n11846), .ZN(n9154) );
  XNOR2_X1 U11517 ( .A(n9168), .B(n9154), .ZN(n11595) );
  NAND2_X1 U11518 ( .A1(n11595), .A2(n12083), .ZN(n9157) );
  OR2_X1 U11519 ( .A1(n9155), .A2(n11596), .ZN(n9156) );
  NAND2_X1 U11520 ( .A1(n6443), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9166) );
  NAND2_X1 U11521 ( .A1(n12091), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9165) );
  INV_X1 U11522 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9159) );
  NAND2_X1 U11523 ( .A1(n9159), .A2(n9158), .ZN(n9177) );
  NAND2_X1 U11524 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(n9160), .ZN(n9161) );
  NAND2_X1 U11525 ( .A1(n9177), .A2(n9161), .ZN(n12487) );
  NAND2_X1 U11526 ( .A1(n9162), .A2(n12487), .ZN(n9164) );
  NAND2_X1 U11527 ( .A1(n12089), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9163) );
  INV_X1 U11528 ( .A(n12627), .ZN(n12490) );
  NAND2_X1 U11529 ( .A1(n12490), .A2(n11918), .ZN(n9185) );
  AND2_X1 U11530 ( .A1(n13313), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9167) );
  NAND2_X1 U11531 ( .A1(n11846), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9169) );
  AOI22_X1 U11532 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n13310), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n11917), .ZN(n9171) );
  INV_X1 U11533 ( .A(n9171), .ZN(n9172) );
  OR2_X1 U11534 ( .A1(n12086), .A2(n12764), .ZN(n9173) );
  NAND2_X2 U11535 ( .A1(n9174), .A2(n9173), .ZN(n12477) );
  NAND2_X1 U11536 ( .A1(n6444), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9182) );
  NAND2_X1 U11537 ( .A1(n12089), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9181) );
  INV_X1 U11538 ( .A(n9177), .ZN(n9176) );
  INV_X1 U11539 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n9175) );
  NAND2_X1 U11540 ( .A1(n9176), .A2(n9175), .ZN(n9296) );
  NAND2_X1 U11541 ( .A1(n9177), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9178) );
  NAND2_X1 U11542 ( .A1(n9296), .A2(n9178), .ZN(n12476) );
  NAND2_X1 U11543 ( .A1(n9162), .A2(n12476), .ZN(n9180) );
  NAND2_X1 U11544 ( .A1(n12091), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9179) );
  NAND2_X1 U11545 ( .A1(n12477), .A2(n11956), .ZN(n9290) );
  AOI21_X1 U11546 ( .B1(n12480), .B2(n9185), .A(n12108), .ZN(n9183) );
  INV_X1 U11547 ( .A(n9183), .ZN(n9184) );
  NAND2_X1 U11548 ( .A1(n14948), .A2(n9184), .ZN(n9197) );
  INV_X1 U11549 ( .A(n9269), .ZN(n9196) );
  INV_X1 U11550 ( .A(n9296), .ZN(n9186) );
  NAND2_X1 U11551 ( .A1(n8819), .A2(n9186), .ZN(n12095) );
  NAND2_X1 U11552 ( .A1(n6444), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9189) );
  NAND2_X1 U11553 ( .A1(n6460), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9188) );
  NAND2_X1 U11554 ( .A1(n12089), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9187) );
  INV_X1 U11555 ( .A(n9190), .ZN(n12299) );
  AND2_X1 U11556 ( .A1(n12299), .A2(n10118), .ZN(n10126) );
  OR2_X1 U11557 ( .A1(n9193), .A2(n10126), .ZN(n9192) );
  NAND2_X2 U11558 ( .A1(n12302), .A2(n10145), .ZN(n12273) );
  OR2_X1 U11559 ( .A1(n11918), .A2(n12055), .ZN(n9194) );
  OAI21_X1 U11560 ( .B1(n10787), .B2(n12057), .A(n9194), .ZN(n11983) );
  OAI21_X1 U11561 ( .B1(n9198), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9200) );
  INV_X1 U11562 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9199) );
  XNOR2_X1 U11563 ( .A(n9200), .B(n9199), .ZN(n10169) );
  NAND2_X1 U11564 ( .A1(n10169), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12751) );
  NAND2_X1 U11565 ( .A1(n9201), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9202) );
  INV_X1 U11566 ( .A(n9203), .ZN(n9209) );
  NAND2_X1 U11567 ( .A1(n9209), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9204) );
  MUX2_X1 U11568 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9204), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9205) );
  NAND2_X1 U11569 ( .A1(n9205), .A2(n9201), .ZN(n11499) );
  INV_X1 U11570 ( .A(n9206), .ZN(n9207) );
  NAND2_X1 U11571 ( .A1(n9207), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9208) );
  MUX2_X1 U11572 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9208), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n9210) );
  NAND2_X1 U11573 ( .A1(n9210), .A2(n9209), .ZN(n11305) );
  NOR2_X1 U11574 ( .A1(n11499), .A2(n11305), .ZN(n9211) );
  AND2_X1 U11575 ( .A1(n9217), .A2(n9211), .ZN(n9743) );
  XNOR2_X1 U11576 ( .A(n11305), .B(P3_B_REG_SCAN_IN), .ZN(n9212) );
  INV_X1 U11577 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9213) );
  INV_X1 U11578 ( .A(n11305), .ZN(n9214) );
  OR2_X1 U11579 ( .A1(n9217), .A2(n9214), .ZN(n9215) );
  INV_X1 U11580 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9216) );
  NAND2_X1 U11581 ( .A1(n9802), .A2(n9216), .ZN(n9219) );
  INV_X1 U11582 ( .A(n9217), .ZN(n11583) );
  NAND2_X1 U11583 ( .A1(n11583), .A2(n11499), .ZN(n9218) );
  NAND2_X1 U11584 ( .A1(n12752), .A2(n12750), .ZN(n9559) );
  INV_X1 U11585 ( .A(n12752), .ZN(n9220) );
  INV_X1 U11586 ( .A(n12750), .ZN(n9282) );
  NAND2_X1 U11587 ( .A1(n9220), .A2(n9282), .ZN(n9565) );
  NOR2_X1 U11588 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .ZN(
        n9224) );
  NOR4_X1 U11589 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n9223) );
  NOR4_X1 U11590 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n9222) );
  NOR4_X1 U11591 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n9221) );
  NAND4_X1 U11592 ( .A1(n9224), .A2(n9223), .A3(n9222), .A4(n9221), .ZN(n9230)
         );
  NOR4_X1 U11593 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9228) );
  NOR4_X1 U11594 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n9227) );
  NOR4_X1 U11595 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9226) );
  NOR4_X1 U11596 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9225) );
  NAND4_X1 U11597 ( .A1(n9228), .A2(n9227), .A3(n9226), .A4(n9225), .ZN(n9229)
         );
  OAI21_X1 U11598 ( .B1(n9230), .B2(n9229), .A(n9802), .ZN(n9563) );
  NAND4_X1 U11599 ( .A1(n12298), .A2(n9559), .A3(n9565), .A4(n9563), .ZN(n9280) );
  NAND2_X1 U11600 ( .A1(n12302), .A2(n12459), .ZN(n9231) );
  OAI21_X1 U11601 ( .B1(n15001), .B2(n9259), .A(n9231), .ZN(n9232) );
  NAND2_X1 U11602 ( .A1(n10537), .A2(n12459), .ZN(n12290) );
  NAND2_X1 U11603 ( .A1(n9232), .A2(n12290), .ZN(n9233) );
  NAND2_X1 U11604 ( .A1(n9233), .A2(n12273), .ZN(n9234) );
  NAND2_X1 U11605 ( .A1(n9234), .A2(n9282), .ZN(n9237) );
  INV_X1 U11606 ( .A(n12290), .ZN(n12297) );
  AND2_X1 U11607 ( .A1(n9259), .A2(n12459), .ZN(n9235) );
  NAND2_X1 U11608 ( .A1(n12302), .A2(n9235), .ZN(n9263) );
  NAND2_X1 U11609 ( .A1(n12273), .A2(n9263), .ZN(n9283) );
  NAND2_X1 U11610 ( .A1(n10171), .A2(n9283), .ZN(n9281) );
  NAND2_X1 U11611 ( .A1(n9281), .A2(n12750), .ZN(n9236) );
  NAND2_X1 U11612 ( .A1(n9237), .A2(n9236), .ZN(n9238) );
  NOR2_X4 U11613 ( .A1(n9280), .A2(n9238), .ZN(n15034) );
  MUX2_X1 U11614 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n12673), .S(n15034), .Z(
        n9239) );
  INV_X1 U11615 ( .A(n9239), .ZN(n9268) );
  INV_X1 U11616 ( .A(n10252), .ZN(n10546) );
  INV_X1 U11617 ( .A(n12116), .ZN(n14938) );
  INV_X1 U11618 ( .A(n14943), .ZN(n10248) );
  NAND2_X1 U11619 ( .A1(n10161), .A2(n10248), .ZN(n12151) );
  NAND2_X1 U11620 ( .A1(n9241), .A2(n12151), .ZN(n10479) );
  NAND2_X1 U11621 ( .A1(n10479), .A2(n10481), .ZN(n9242) );
  NAND2_X1 U11622 ( .A1(n9242), .A2(n12153), .ZN(n10799) );
  INV_X1 U11623 ( .A(n12115), .ZN(n12155) );
  NAND2_X1 U11624 ( .A1(n10799), .A2(n12155), .ZN(n9243) );
  INV_X1 U11625 ( .A(n12330), .ZN(n10492) );
  NAND2_X1 U11626 ( .A1(n10492), .A2(n14984), .ZN(n12157) );
  NAND2_X1 U11627 ( .A1(n9243), .A2(n12157), .ZN(n10788) );
  NAND2_X1 U11628 ( .A1(n10788), .A2(n12160), .ZN(n9244) );
  NAND2_X1 U11629 ( .A1(n9244), .A2(n12165), .ZN(n11130) );
  INV_X1 U11630 ( .A(n12112), .ZN(n11129) );
  NAND2_X1 U11631 ( .A1(n11130), .A2(n11129), .ZN(n11128) );
  NAND2_X1 U11632 ( .A1(n11128), .A2(n12168), .ZN(n11011) );
  INV_X1 U11633 ( .A(n11014), .ZN(n12171) );
  INV_X1 U11634 ( .A(n15015), .ZN(n12192) );
  NOR2_X1 U11635 ( .A1(n12325), .A2(n12192), .ZN(n9246) );
  OR2_X2 U11636 ( .A1(n11375), .A2(n9246), .ZN(n9248) );
  NAND2_X1 U11637 ( .A1(n12325), .A2(n12192), .ZN(n9247) );
  INV_X1 U11638 ( .A(n9249), .ZN(n12186) );
  XNOR2_X1 U11639 ( .A(n12323), .B(n12187), .ZN(n12190) );
  NAND2_X1 U11640 ( .A1(n11459), .A2(n14312), .ZN(n12199) );
  INV_X1 U11641 ( .A(n12206), .ZN(n9251) );
  INV_X1 U11642 ( .A(n9252), .ZN(n12211) );
  AOI21_X2 U11643 ( .B1(n11658), .B2(n12210), .A(n12211), .ZN(n12612) );
  XNOR2_X1 U11644 ( .A(n12738), .B(n12318), .ZN(n12606) );
  INV_X1 U11645 ( .A(n12738), .ZN(n12215) );
  NOR2_X1 U11646 ( .A1(n12215), .A2(n12318), .ZN(n12224) );
  INV_X1 U11647 ( .A(n12591), .ZN(n9253) );
  NAND2_X1 U11648 ( .A1(n12111), .A2(n12316), .ZN(n12237) );
  NOR2_X1 U11649 ( .A1(n12111), .A2(n12316), .ZN(n12239) );
  INV_X1 U11650 ( .A(n12243), .ZN(n9254) );
  AOI21_X1 U11651 ( .B1(n12561), .B2(n12560), .A(n9254), .ZN(n12548) );
  INV_X1 U11652 ( .A(n9255), .ZN(n12249) );
  OAI21_X1 U11653 ( .B1(n12548), .B2(n12249), .A(n12247), .ZN(n12539) );
  NAND2_X1 U11654 ( .A1(n12703), .A2(n11964), .ZN(n12110) );
  NOR2_X1 U11655 ( .A1(n12703), .A2(n11964), .ZN(n12134) );
  INV_X1 U11656 ( .A(n12531), .ZN(n12528) );
  NAND2_X1 U11657 ( .A1(n12255), .A2(n12312), .ZN(n12258) );
  INV_X1 U11658 ( .A(n12691), .ZN(n9256) );
  NOR2_X1 U11659 ( .A1(n9256), .A2(n12311), .ZN(n12259) );
  NAND2_X1 U11660 ( .A1(n12680), .A2(n12309), .ZN(n12269) );
  INV_X1 U11661 ( .A(n12484), .ZN(n9257) );
  NAND2_X1 U11662 ( .A1(n12627), .A2(n11918), .ZN(n9289) );
  NAND2_X1 U11663 ( .A1(n9257), .A2(n9289), .ZN(n9258) );
  XNOR2_X2 U11664 ( .A(n9258), .B(n12108), .ZN(n12675) );
  OR2_X1 U11665 ( .A1(n9259), .A2(n10145), .ZN(n9260) );
  XNOR2_X1 U11666 ( .A(n12302), .B(n9260), .ZN(n9262) );
  OR2_X1 U11667 ( .A1(n10145), .A2(n12454), .ZN(n9261) );
  NAND2_X1 U11668 ( .A1(n9262), .A2(n9261), .ZN(n10166) );
  AND2_X1 U11669 ( .A1(n15001), .A2(n12297), .ZN(n9265) );
  INV_X1 U11670 ( .A(n9263), .ZN(n9264) );
  AOI21_X1 U11671 ( .B1(n10166), .B2(n9265), .A(n9264), .ZN(n14936) );
  NAND2_X1 U11672 ( .A1(n10537), .A2(n12454), .ZN(n14955) );
  OR2_X1 U11673 ( .A1(n12302), .A2(n14955), .ZN(n15018) );
  NAND2_X1 U11674 ( .A1(n14936), .A2(n15018), .ZN(n15007) );
  NAND2_X1 U11675 ( .A1(n15034), .A2(n15007), .ZN(n12664) );
  INV_X1 U11676 ( .A(n12477), .ZN(n12674) );
  NAND2_X1 U11677 ( .A1(n15034), .A2(n15014), .ZN(n12655) );
  OAI22_X1 U11678 ( .A1(n12675), .A2(n12664), .B1(n12674), .B2(n12655), .ZN(
        n9266) );
  INV_X1 U11679 ( .A(n9266), .ZN(n9267) );
  NAND2_X1 U11680 ( .A1(n13310), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9271) );
  XNOR2_X1 U11681 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n11908) );
  XNOR2_X1 U11682 ( .A(n11911), .B(n11908), .ZN(n12759) );
  NAND2_X1 U11683 ( .A1(n12759), .A2(n12083), .ZN(n9273) );
  OR2_X1 U11684 ( .A1(n12086), .A2(n12762), .ZN(n9272) );
  NAND2_X1 U11685 ( .A1(n9293), .A2(n10787), .ZN(n12099) );
  XNOR2_X1 U11686 ( .A(n9274), .B(n12130), .ZN(n9279) );
  AOI21_X1 U11687 ( .B1(n12299), .B2(P3_B_REG_SCAN_IN), .A(n12057), .ZN(n12469) );
  NAND2_X1 U11688 ( .A1(n12089), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9277) );
  NAND2_X1 U11689 ( .A1(n6443), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9276) );
  NAND2_X1 U11690 ( .A1(n6460), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9275) );
  NAND4_X1 U11691 ( .A1(n12095), .A2(n9277), .A3(n9276), .A4(n9275), .ZN(
        n12306) );
  INV_X1 U11692 ( .A(n11956), .ZN(n12307) );
  AOI22_X1 U11693 ( .A1(n12469), .A2(n12306), .B1(n12307), .B2(n12300), .ZN(
        n9278) );
  OAI21_X1 U11694 ( .B1(n9279), .B2(n14939), .A(n9278), .ZN(n9569) );
  INV_X1 U11695 ( .A(n9280), .ZN(n9287) );
  NAND2_X1 U11696 ( .A1(n9282), .A2(n9281), .ZN(n9285) );
  NAND2_X1 U11697 ( .A1(n12750), .A2(n9283), .ZN(n9284) );
  AND2_X1 U11698 ( .A1(n9285), .A2(n9284), .ZN(n9286) );
  NAND2_X1 U11699 ( .A1(n9287), .A2(n9286), .ZN(n9295) );
  NOR2_X1 U11700 ( .A1(n15001), .A2(n14955), .ZN(n9288) );
  NAND2_X1 U11701 ( .A1(n12298), .A2(n9288), .ZN(n11656) );
  INV_X2 U11702 ( .A(n14965), .ZN(n14963) );
  NAND2_X1 U11703 ( .A1(n9569), .A2(n14963), .ZN(n9301) );
  NAND2_X1 U11704 ( .A1(n9290), .A2(n9289), .ZN(n12274) );
  XOR2_X1 U11705 ( .A(n12130), .B(n12096), .Z(n9572) );
  INV_X1 U11706 ( .A(n10145), .ZN(n12140) );
  OR2_X1 U11707 ( .A1(n14955), .A2(n12140), .ZN(n9291) );
  OR2_X1 U11708 ( .A1(n14965), .A2(n14936), .ZN(n9292) );
  INV_X1 U11709 ( .A(n9293), .ZN(n9571) );
  NAND2_X1 U11710 ( .A1(n15014), .A2(n14955), .ZN(n9294) );
  NOR2_X1 U11711 ( .A1(n11656), .A2(n9296), .ZN(n12470) );
  INV_X1 U11712 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n9297) );
  NOR2_X1 U11713 ( .A1(n14963), .A2(n9297), .ZN(n9298) );
  NOR2_X1 U11714 ( .A1(n12470), .A2(n9298), .ZN(n9299) );
  NAND2_X1 U11715 ( .A1(n9301), .A2(n9300), .ZN(P3_U3204) );
  MUX2_X1 U11716 ( .A(n12846), .B(n13074), .S(n9513), .Z(n9446) );
  MUX2_X1 U11717 ( .A(n13226), .B(n13080), .S(n9513), .Z(n9445) );
  NAND2_X1 U11718 ( .A1(n9580), .A2(n9302), .ZN(n9307) );
  NAND2_X1 U11719 ( .A1(n12899), .A2(n10561), .ZN(n9530) );
  NAND2_X1 U11720 ( .A1(n9530), .A2(n9357), .ZN(n9305) );
  NAND3_X1 U11721 ( .A1(n9307), .A2(n9306), .A3(n9305), .ZN(n9310) );
  MUX2_X1 U11722 ( .A(n10889), .B(n12898), .S(n9304), .Z(n9311) );
  NAND2_X1 U11723 ( .A1(n9310), .A2(n9311), .ZN(n9309) );
  MUX2_X1 U11724 ( .A(n12898), .B(n10889), .S(n9304), .Z(n9308) );
  NAND2_X1 U11725 ( .A1(n9309), .A2(n9308), .ZN(n9315) );
  INV_X1 U11726 ( .A(n9310), .ZN(n9313) );
  INV_X1 U11727 ( .A(n9311), .ZN(n9312) );
  NAND2_X1 U11728 ( .A1(n9313), .A2(n9312), .ZN(n9314) );
  MUX2_X1 U11729 ( .A(n10881), .B(n12897), .S(n9304), .Z(n9317) );
  INV_X1 U11730 ( .A(n9319), .ZN(n9320) );
  MUX2_X1 U11731 ( .A(n14785), .B(n12896), .S(n9473), .Z(n9324) );
  INV_X1 U11732 ( .A(n9357), .ZN(n9473) );
  MUX2_X1 U11733 ( .A(n12896), .B(n14785), .S(n9473), .Z(n9321) );
  NAND2_X1 U11734 ( .A1(n9322), .A2(n9321), .ZN(n9328) );
  INV_X1 U11735 ( .A(n9323), .ZN(n9326) );
  INV_X1 U11736 ( .A(n9324), .ZN(n9325) );
  NAND2_X1 U11737 ( .A1(n9326), .A2(n9325), .ZN(n9327) );
  MUX2_X1 U11738 ( .A(n12895), .B(n14793), .S(n9473), .Z(n9330) );
  MUX2_X1 U11739 ( .A(n14793), .B(n12895), .S(n9473), .Z(n9329) );
  MUX2_X1 U11740 ( .A(n11032), .B(n12894), .S(n9402), .Z(n9334) );
  NAND2_X1 U11741 ( .A1(n9333), .A2(n9334), .ZN(n9332) );
  MUX2_X1 U11742 ( .A(n12894), .B(n11032), .S(n9402), .Z(n9331) );
  NAND2_X1 U11743 ( .A1(n9332), .A2(n9331), .ZN(n9338) );
  INV_X1 U11744 ( .A(n9333), .ZN(n9336) );
  INV_X1 U11745 ( .A(n9334), .ZN(n9335) );
  NAND2_X1 U11746 ( .A1(n9336), .A2(n9335), .ZN(n9337) );
  MUX2_X1 U11747 ( .A(n12893), .B(n11048), .S(n9402), .Z(n9342) );
  NAND2_X1 U11748 ( .A1(n9341), .A2(n9342), .ZN(n9340) );
  MUX2_X1 U11749 ( .A(n11048), .B(n12893), .S(n9402), .Z(n9339) );
  NAND2_X1 U11750 ( .A1(n9340), .A2(n9339), .ZN(n9346) );
  INV_X1 U11751 ( .A(n9341), .ZN(n9344) );
  INV_X1 U11752 ( .A(n9342), .ZN(n9343) );
  NAND2_X1 U11753 ( .A1(n9344), .A2(n9343), .ZN(n9345) );
  MUX2_X1 U11754 ( .A(n12892), .B(n11247), .S(n9357), .Z(n9348) );
  MUX2_X1 U11755 ( .A(n12892), .B(n11247), .S(n9402), .Z(n9347) );
  MUX2_X1 U11756 ( .A(n12891), .B(n11227), .S(n9513), .Z(n9352) );
  NAND2_X1 U11757 ( .A1(n9351), .A2(n9352), .ZN(n9350) );
  MUX2_X1 U11758 ( .A(n12891), .B(n11227), .S(n9357), .Z(n9349) );
  NAND2_X1 U11759 ( .A1(n9350), .A2(n9349), .ZN(n9356) );
  INV_X1 U11760 ( .A(n9351), .ZN(n9354) );
  INV_X1 U11761 ( .A(n9352), .ZN(n9353) );
  NAND2_X1 U11762 ( .A1(n9354), .A2(n9353), .ZN(n9355) );
  NAND2_X1 U11763 ( .A1(n9356), .A2(n9355), .ZN(n9360) );
  MUX2_X1 U11764 ( .A(n12890), .B(n14829), .S(n9357), .Z(n9361) );
  NAND2_X1 U11765 ( .A1(n9360), .A2(n9361), .ZN(n9359) );
  MUX2_X1 U11766 ( .A(n12890), .B(n14829), .S(n9513), .Z(n9358) );
  NAND2_X1 U11767 ( .A1(n9359), .A2(n9358), .ZN(n9365) );
  INV_X1 U11768 ( .A(n9360), .ZN(n9363) );
  INV_X1 U11769 ( .A(n9361), .ZN(n9362) );
  NAND2_X1 U11770 ( .A1(n9363), .A2(n9362), .ZN(n9364) );
  MUX2_X1 U11771 ( .A(n12889), .B(n14842), .S(n9513), .Z(n9367) );
  MUX2_X1 U11772 ( .A(n12889), .B(n14842), .S(n9357), .Z(n9366) );
  MUX2_X1 U11773 ( .A(n12888), .B(n11253), .S(n9357), .Z(n9371) );
  NAND2_X1 U11774 ( .A1(n9370), .A2(n9371), .ZN(n9369) );
  MUX2_X1 U11775 ( .A(n12888), .B(n11253), .S(n9402), .Z(n9368) );
  NAND2_X1 U11776 ( .A1(n9369), .A2(n9368), .ZN(n9375) );
  INV_X1 U11777 ( .A(n9370), .ZN(n9373) );
  INV_X1 U11778 ( .A(n9371), .ZN(n9372) );
  NAND2_X1 U11779 ( .A1(n9373), .A2(n9372), .ZN(n9374) );
  INV_X1 U11780 ( .A(n9357), .ZN(n9513) );
  MUX2_X1 U11781 ( .A(n12887), .B(n13273), .S(n9513), .Z(n9378) );
  MUX2_X1 U11782 ( .A(n12887), .B(n13273), .S(n9411), .Z(n9376) );
  INV_X1 U11783 ( .A(n9378), .ZN(n9379) );
  MUX2_X1 U11784 ( .A(n12886), .B(n9640), .S(n9411), .Z(n9383) );
  MUX2_X1 U11785 ( .A(n12886), .B(n9640), .S(n9513), .Z(n9380) );
  NAND2_X1 U11786 ( .A1(n9381), .A2(n9380), .ZN(n9387) );
  INV_X1 U11787 ( .A(n9382), .ZN(n9385) );
  INV_X1 U11788 ( .A(n9383), .ZN(n9384) );
  NAND2_X1 U11789 ( .A1(n9385), .A2(n9384), .ZN(n9386) );
  MUX2_X1 U11790 ( .A(n12885), .B(n11730), .S(n9513), .Z(n9390) );
  MUX2_X1 U11791 ( .A(n12885), .B(n11730), .S(n9411), .Z(n9388) );
  INV_X1 U11792 ( .A(n9390), .ZN(n9391) );
  INV_X1 U11793 ( .A(n9357), .ZN(n9402) );
  INV_X1 U11794 ( .A(n9402), .ZN(n9411) );
  MUX2_X1 U11795 ( .A(n12884), .B(n13269), .S(n9411), .Z(n9395) );
  MUX2_X1 U11796 ( .A(n12884), .B(n13269), .S(n9402), .Z(n9392) );
  NAND2_X1 U11797 ( .A1(n9393), .A2(n9392), .ZN(n9399) );
  INV_X1 U11798 ( .A(n9394), .ZN(n9397) );
  INV_X1 U11799 ( .A(n9395), .ZN(n9396) );
  NAND2_X1 U11800 ( .A1(n9397), .A2(n9396), .ZN(n9398) );
  MUX2_X1 U11801 ( .A(n12883), .B(n13262), .S(n9402), .Z(n9401) );
  MUX2_X1 U11802 ( .A(n12883), .B(n13262), .S(n9411), .Z(n9400) );
  MUX2_X1 U11803 ( .A(n13151), .B(n13258), .S(n9411), .Z(n9406) );
  NAND2_X1 U11804 ( .A1(n9405), .A2(n9406), .ZN(n9404) );
  MUX2_X1 U11805 ( .A(n13151), .B(n13258), .S(n9402), .Z(n9403) );
  NAND2_X1 U11806 ( .A1(n9404), .A2(n9403), .ZN(n9410) );
  INV_X1 U11807 ( .A(n9405), .ZN(n9408) );
  INV_X1 U11808 ( .A(n9406), .ZN(n9407) );
  NAND2_X1 U11809 ( .A1(n9408), .A2(n9407), .ZN(n9409) );
  MUX2_X1 U11810 ( .A(n12882), .B(n13253), .S(n9513), .Z(n9415) );
  NAND2_X1 U11811 ( .A1(n9414), .A2(n9415), .ZN(n9413) );
  MUX2_X1 U11812 ( .A(n12882), .B(n13253), .S(n9411), .Z(n9412) );
  INV_X1 U11813 ( .A(n9414), .ZN(n9417) );
  INV_X1 U11814 ( .A(n9415), .ZN(n9416) );
  MUX2_X1 U11815 ( .A(n13154), .B(n13246), .S(n9411), .Z(n9418) );
  MUX2_X1 U11816 ( .A(n13154), .B(n13246), .S(n9513), .Z(n9419) );
  MUX2_X1 U11817 ( .A(n12797), .B(n13242), .S(n9513), .Z(n9421) );
  MUX2_X1 U11818 ( .A(n13118), .B(n12881), .S(n9513), .Z(n9420) );
  OAI21_X1 U11819 ( .B1(n9422), .B2(n9421), .A(n9420), .ZN(n9424) );
  NAND2_X1 U11820 ( .A1(n9422), .A2(n9421), .ZN(n9423) );
  NAND2_X1 U11821 ( .A1(n9424), .A2(n9423), .ZN(n9426) );
  MUX2_X1 U11822 ( .A(n13236), .B(n13079), .S(n9473), .Z(n9427) );
  MUX2_X1 U11823 ( .A(n13079), .B(n13236), .S(n9473), .Z(n9425) );
  MUX2_X1 U11824 ( .A(n13066), .B(n13085), .S(n9513), .Z(n9429) );
  MUX2_X1 U11825 ( .A(n13231), .B(n12880), .S(n9513), .Z(n9428) );
  NAND2_X1 U11826 ( .A1(n9430), .A2(n9429), .ZN(n9431) );
  NAND2_X1 U11827 ( .A1(n9432), .A2(n9431), .ZN(n9435) );
  MUX2_X1 U11828 ( .A(n9697), .B(n13038), .S(n9357), .Z(n9443) );
  MUX2_X1 U11829 ( .A(n13017), .B(n13214), .S(n9513), .Z(n9442) );
  NAND2_X1 U11830 ( .A1(n9443), .A2(n9442), .ZN(n9440) );
  MUX2_X1 U11831 ( .A(n13068), .B(n13219), .S(n9411), .Z(n9437) );
  MUX2_X1 U11832 ( .A(n13036), .B(n9433), .S(n9513), .Z(n9436) );
  NAND2_X1 U11833 ( .A1(n9437), .A2(n9436), .ZN(n9434) );
  AND2_X1 U11834 ( .A1(n9440), .A2(n9434), .ZN(n9444) );
  OAI211_X1 U11835 ( .C1(n9446), .C2(n9445), .A(n9435), .B(n9444), .ZN(n9453)
         );
  MUX2_X1 U11836 ( .A(n12814), .B(n13028), .S(n9402), .Z(n9476) );
  MUX2_X1 U11837 ( .A(n13035), .B(n13209), .S(n9411), .Z(n9475) );
  INV_X1 U11838 ( .A(n9436), .ZN(n9439) );
  INV_X1 U11839 ( .A(n9437), .ZN(n9438) );
  NAND3_X1 U11840 ( .A1(n9440), .A2(n9439), .A3(n9438), .ZN(n9441) );
  OAI21_X1 U11841 ( .B1(n9443), .B2(n9442), .A(n9441), .ZN(n9451) );
  INV_X1 U11842 ( .A(n9444), .ZN(n9449) );
  INV_X1 U11843 ( .A(n9445), .ZN(n9448) );
  INV_X1 U11844 ( .A(n9446), .ZN(n9447) );
  NOR3_X1 U11845 ( .A1(n9449), .A2(n9448), .A3(n9447), .ZN(n9450) );
  AOI211_X1 U11846 ( .C1(n9476), .C2(n9475), .A(n9451), .B(n9450), .ZN(n9452)
         );
  NAND2_X1 U11847 ( .A1(n9453), .A2(n9452), .ZN(n9479) );
  NAND2_X1 U11848 ( .A1(n13295), .A2(n9469), .ZN(n9455) );
  NAND2_X1 U11849 ( .A1(n9485), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9454) );
  NAND2_X1 U11850 ( .A1(n9488), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9458) );
  NAND2_X1 U11851 ( .A1(n7964), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9457) );
  NAND2_X1 U11852 ( .A1(n6445), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9456) );
  AND3_X1 U11853 ( .A1(n9458), .A2(n9457), .A3(n9456), .ZN(n9512) );
  XNOR2_X1 U11854 ( .A(n13188), .B(n9512), .ZN(n9526) );
  NAND2_X1 U11855 ( .A1(n13307), .A2(n9469), .ZN(n9460) );
  NAND2_X1 U11856 ( .A1(n9485), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9459) );
  MUX2_X1 U11857 ( .A(n12977), .B(n13202), .S(n9513), .Z(n9500) );
  INV_X1 U11858 ( .A(n12977), .ZN(n12961) );
  MUX2_X1 U11859 ( .A(n12961), .B(n12995), .S(n9411), .Z(n9499) );
  OR2_X1 U11860 ( .A1(n12965), .A2(n6441), .ZN(n9468) );
  INV_X1 U11861 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9464) );
  NAND2_X1 U11862 ( .A1(n7759), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9463) );
  NAND2_X1 U11863 ( .A1(n6446), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9462) );
  OAI211_X1 U11864 ( .C1(n6439), .C2(n9464), .A(n9463), .B(n9462), .ZN(n9466)
         );
  INV_X1 U11865 ( .A(n9466), .ZN(n9467) );
  AND2_X1 U11866 ( .A1(n9468), .A2(n9467), .ZN(n9735) );
  NAND2_X1 U11867 ( .A1(n9470), .A2(n9469), .ZN(n9472) );
  NAND2_X1 U11868 ( .A1(n9485), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9471) );
  MUX2_X1 U11869 ( .A(n9735), .B(n13196), .S(n9411), .Z(n9496) );
  INV_X1 U11870 ( .A(n13196), .ZN(n12964) );
  MUX2_X1 U11871 ( .A(n12989), .B(n12964), .S(n9473), .Z(n9495) );
  NAND2_X1 U11872 ( .A1(n9496), .A2(n9495), .ZN(n9501) );
  OAI21_X1 U11873 ( .B1(n9500), .B2(n9499), .A(n9501), .ZN(n9474) );
  MUX2_X1 U11874 ( .A(n12958), .B(n13007), .S(n9513), .Z(n9481) );
  MUX2_X1 U11875 ( .A(n12772), .B(n13018), .S(n9402), .Z(n9480) );
  OAI22_X1 U11876 ( .A1(n9481), .A2(n9480), .B1(n9476), .B2(n9475), .ZN(n9477)
         );
  NAND2_X1 U11877 ( .A1(n9479), .A2(n9478), .ZN(n9511) );
  INV_X1 U11878 ( .A(n9480), .ZN(n9483) );
  INV_X1 U11879 ( .A(n9481), .ZN(n9482) );
  NOR3_X1 U11880 ( .A1(n9484), .A2(n9483), .A3(n9482), .ZN(n9505) );
  INV_X1 U11881 ( .A(n13303), .ZN(n9486) );
  AOI22_X1 U11882 ( .A1(n9486), .A2(n9469), .B1(n9485), .B2(
        P1_DATAO_REG_30__SCAN_IN), .ZN(n9487) );
  NAND2_X1 U11883 ( .A1(n9488), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9491) );
  NAND2_X1 U11884 ( .A1(n7759), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9490) );
  NAND2_X1 U11885 ( .A1(n6446), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9489) );
  AND3_X1 U11886 ( .A1(n9491), .A2(n9490), .A3(n9489), .ZN(n9527) );
  INV_X1 U11887 ( .A(n9512), .ZN(n12950) );
  OAI211_X1 U11888 ( .C1(n9492), .C2(n9723), .A(n9548), .B(n9522), .ZN(n9493)
         );
  AOI21_X1 U11889 ( .B1(n12950), .B2(n9402), .A(n9493), .ZN(n9494) );
  OAI22_X1 U11890 ( .A1(n9487), .A2(n9513), .B1(n9527), .B2(n9494), .ZN(n9507)
         );
  MUX2_X1 U11891 ( .A(n9527), .B(n9487), .S(n9513), .Z(n9506) );
  INV_X1 U11892 ( .A(n9495), .ZN(n9498) );
  INV_X1 U11893 ( .A(n9496), .ZN(n9497) );
  AOI22_X1 U11894 ( .A1(n9507), .A2(n9506), .B1(n9498), .B2(n9497), .ZN(n9503)
         );
  NAND3_X1 U11895 ( .A1(n9501), .A2(n9500), .A3(n9499), .ZN(n9502) );
  AOI21_X1 U11896 ( .B1(n9503), .B2(n9502), .A(n9526), .ZN(n9504) );
  INV_X1 U11897 ( .A(n9506), .ZN(n9509) );
  INV_X1 U11898 ( .A(n9507), .ZN(n9508) );
  AOI21_X1 U11899 ( .B1(n9511), .B2(n7373), .A(n9510), .ZN(n9517) );
  NOR2_X1 U11900 ( .A1(n9513), .A2(n9512), .ZN(n9515) );
  NOR2_X1 U11901 ( .A1(n9411), .A2(n12950), .ZN(n9514) );
  MUX2_X1 U11902 ( .A(n9515), .B(n9514), .S(n13188), .Z(n9516) );
  OAI21_X1 U11903 ( .B1(n10947), .B2(n12997), .A(n9522), .ZN(n9518) );
  MUX2_X1 U11904 ( .A(n9524), .B(n9548), .S(n9723), .Z(n9520) );
  NAND2_X1 U11905 ( .A1(n9863), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11346) );
  OAI21_X1 U11906 ( .B1(n9525), .B2(n7385), .A(n9521), .ZN(n9554) );
  INV_X1 U11907 ( .A(n13311), .ZN(n12949) );
  INV_X1 U11908 ( .A(n9522), .ZN(n9733) );
  NAND4_X1 U11909 ( .A1(n14767), .A2(n12949), .A3(n9733), .A4(n13152), .ZN(
        n9523) );
  OAI211_X1 U11910 ( .C1(n9524), .C2(n11346), .A(n9523), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9553) );
  INV_X1 U11911 ( .A(n9525), .ZN(n9551) );
  INV_X1 U11912 ( .A(n9526), .ZN(n9546) );
  INV_X1 U11913 ( .A(n9527), .ZN(n12975) );
  XOR2_X1 U11914 ( .A(n12975), .B(n9487), .Z(n9545) );
  NAND2_X1 U11915 ( .A1(n12995), .A2(n12977), .ZN(n9528) );
  XNOR2_X1 U11916 ( .A(n13118), .B(n12881), .ZN(n13113) );
  INV_X1 U11917 ( .A(n9530), .ZN(n10472) );
  NOR2_X1 U11918 ( .A1(n10472), .A2(n10557), .ZN(n14768) );
  NAND4_X1 U11919 ( .A1(n9529), .A2(n10876), .A3(n9723), .A4(n14768), .ZN(
        n9531) );
  NOR4_X1 U11920 ( .A1(n11025), .A2(n11269), .A3(n9531), .A4(n10821), .ZN(
        n9532) );
  NAND4_X1 U11921 ( .A1(n9532), .A2(n11223), .A3(n11238), .A4(n11040), .ZN(
        n9533) );
  NOR4_X1 U11922 ( .A1(n11149), .A2(n10978), .A3(n11207), .A4(n9533), .ZN(
        n9535) );
  NAND4_X1 U11923 ( .A1(n11741), .A2(n9535), .A3(n11474), .A4(n9534), .ZN(
        n9536) );
  NOR4_X1 U11924 ( .A1(n11718), .A2(n11708), .A3(n9536), .A4(n13180), .ZN(
        n9537) );
  XNOR2_X1 U11925 ( .A(n13246), .B(n13154), .ZN(n13126) );
  NAND4_X1 U11926 ( .A1(n13113), .A2(n9537), .A3(n13126), .A4(n13150), .ZN(
        n9538) );
  NOR3_X1 U11927 ( .A1(n13083), .A2(n13104), .A3(n9538), .ZN(n9540) );
  NAND4_X1 U11928 ( .A1(n13015), .A2(n9540), .A3(n9539), .A4(n13052), .ZN(
        n9541) );
  NOR4_X1 U11929 ( .A1(n12984), .A2(n9543), .A3(n9542), .A4(n9541), .ZN(n9544)
         );
  NAND4_X1 U11930 ( .A1(n9546), .A2(n9545), .A3(n9544), .A4(n12970), .ZN(n9547) );
  XOR2_X1 U11931 ( .A(n12997), .B(n9547), .Z(n9549) );
  NOR3_X1 U11932 ( .A1(n9549), .A2(n9548), .A3(n11346), .ZN(n9550) );
  OAI21_X1 U11933 ( .B1(n9551), .B2(n9723), .A(n9550), .ZN(n9552) );
  OAI211_X1 U11934 ( .C1(n7374), .C2(n9554), .A(n9553), .B(n9552), .ZN(
        P2_U3328) );
  MUX2_X1 U11935 ( .A(P3_REG1_REG_29__SCAN_IN), .B(n9569), .S(n15034), .Z(
        n9555) );
  INV_X1 U11936 ( .A(n9555), .ZN(n9558) );
  OAI22_X1 U11937 ( .A1(n9572), .A2(n12664), .B1(n9571), .B2(n12655), .ZN(
        n9556) );
  INV_X1 U11938 ( .A(n9556), .ZN(n9557) );
  NAND2_X1 U11939 ( .A1(n9558), .A2(n9557), .ZN(P3_U3488) );
  INV_X1 U11940 ( .A(n9559), .ZN(n9560) );
  NAND2_X1 U11941 ( .A1(n9560), .A2(n9563), .ZN(n10167) );
  INV_X1 U11942 ( .A(n9561), .ZN(n9562) );
  OR2_X1 U11943 ( .A1(n10537), .A2(n10145), .ZN(n12293) );
  INV_X1 U11944 ( .A(n12293), .ZN(n10144) );
  NAND2_X1 U11945 ( .A1(n9562), .A2(n10144), .ZN(n10168) );
  AND2_X1 U11946 ( .A1(n10168), .A2(n10389), .ZN(n9567) );
  INV_X1 U11947 ( .A(n10166), .ZN(n9566) );
  INV_X1 U11948 ( .A(n9563), .ZN(n9564) );
  OR2_X1 U11949 ( .A1(n9565), .A2(n9564), .ZN(n10178) );
  OAI22_X1 U11950 ( .A1(n10167), .A2(n9567), .B1(n9566), .B2(n10178), .ZN(
        n9568) );
  MUX2_X1 U11951 ( .A(P3_REG0_REG_29__SCAN_IN), .B(n9569), .S(n15025), .Z(
        n9570) );
  INV_X1 U11952 ( .A(n9570), .ZN(n9575) );
  NAND2_X1 U11953 ( .A1(n15025), .A2(n15007), .ZN(n12748) );
  NAND2_X1 U11954 ( .A1(n15025), .A2(n15014), .ZN(n12730) );
  OAI22_X1 U11955 ( .A1(n9572), .A2(n12748), .B1(n9571), .B2(n12730), .ZN(
        n9573) );
  INV_X1 U11956 ( .A(n9573), .ZN(n9574) );
  NAND2_X1 U11957 ( .A1(n9575), .A2(n9574), .ZN(P3_U3456) );
  INV_X1 U11958 ( .A(n10889), .ZN(n10562) );
  XNOR2_X1 U11959 ( .A(n10562), .B(n9588), .ZN(n9585) );
  INV_X1 U11960 ( .A(n9585), .ZN(n9577) );
  NAND2_X1 U11961 ( .A1(n9596), .A2(n12898), .ZN(n9584) );
  XNOR2_X1 U11962 ( .A(n9577), .B(n9584), .ZN(n10427) );
  NAND2_X1 U11963 ( .A1(n9578), .A2(n14773), .ZN(n9579) );
  AND2_X1 U11964 ( .A1(n9580), .A2(n9579), .ZN(n10473) );
  NAND2_X1 U11965 ( .A1(n9716), .A2(n10561), .ZN(n9581) );
  NAND2_X1 U11966 ( .A1(n10473), .A2(n9581), .ZN(n10426) );
  NAND2_X1 U11967 ( .A1(n10427), .A2(n10426), .ZN(n10425) );
  XNOR2_X1 U11968 ( .A(n9588), .B(n14779), .ZN(n9587) );
  INV_X1 U11969 ( .A(n9587), .ZN(n9583) );
  NAND2_X1 U11970 ( .A1(n9596), .A2(n12897), .ZN(n9586) );
  INV_X1 U11971 ( .A(n9586), .ZN(n9582) );
  NAND2_X1 U11972 ( .A1(n9583), .A2(n9582), .ZN(n10458) );
  INV_X1 U11973 ( .A(n10458), .ZN(n9590) );
  AND2_X1 U11974 ( .A1(n9585), .A2(n9584), .ZN(n10456) );
  AND2_X1 U11975 ( .A1(n9587), .A2(n9586), .ZN(n10659) );
  NAND2_X1 U11976 ( .A1(n9596), .A2(n12896), .ZN(n9591) );
  XNOR2_X1 U11977 ( .A(n9593), .B(n9591), .ZN(n10662) );
  OAI211_X1 U11978 ( .C1(n10425), .C2(n9590), .A(n9589), .B(n10662), .ZN(n9595) );
  INV_X1 U11979 ( .A(n9591), .ZN(n9592) );
  NAND2_X1 U11980 ( .A1(n9593), .A2(n9592), .ZN(n9594) );
  NAND2_X1 U11981 ( .A1(n9595), .A2(n9594), .ZN(n10670) );
  INV_X1 U11982 ( .A(n10670), .ZN(n9603) );
  XNOR2_X1 U11983 ( .A(n9716), .B(n11280), .ZN(n9597) );
  NAND2_X1 U11984 ( .A1(n9596), .A2(n12895), .ZN(n9598) );
  NAND2_X1 U11985 ( .A1(n9597), .A2(n9598), .ZN(n9604) );
  INV_X1 U11986 ( .A(n9597), .ZN(n9600) );
  INV_X1 U11987 ( .A(n9598), .ZN(n9599) );
  NAND2_X1 U11988 ( .A1(n9600), .A2(n9599), .ZN(n9601) );
  NAND2_X1 U11989 ( .A1(n9604), .A2(n9601), .ZN(n10669) );
  NAND2_X1 U11990 ( .A1(n9603), .A2(n9602), .ZN(n10667) );
  NAND2_X1 U11991 ( .A1(n10667), .A2(n9604), .ZN(n10686) );
  XNOR2_X1 U11992 ( .A(n14801), .B(n9716), .ZN(n9605) );
  NAND2_X1 U11993 ( .A1(n9616), .A2(n12894), .ZN(n9606) );
  NAND2_X1 U11994 ( .A1(n9605), .A2(n9606), .ZN(n9610) );
  INV_X1 U11995 ( .A(n9605), .ZN(n9608) );
  INV_X1 U11996 ( .A(n9606), .ZN(n9607) );
  NAND2_X1 U11997 ( .A1(n9608), .A2(n9607), .ZN(n9609) );
  AND2_X1 U11998 ( .A1(n9610), .A2(n9609), .ZN(n10687) );
  XNOR2_X1 U11999 ( .A(n11048), .B(n9709), .ZN(n9611) );
  NAND2_X1 U12000 ( .A1(n9616), .A2(n12893), .ZN(n9612) );
  XNOR2_X1 U12001 ( .A(n9611), .B(n9612), .ZN(n10677) );
  INV_X1 U12002 ( .A(n9611), .ZN(n9614) );
  INV_X1 U12003 ( .A(n9612), .ZN(n9613) );
  NAND2_X1 U12004 ( .A1(n9614), .A2(n9613), .ZN(n9615) );
  XNOR2_X1 U12005 ( .A(n11247), .B(n9716), .ZN(n9619) );
  NAND2_X1 U12006 ( .A1(n9616), .A2(n12892), .ZN(n9617) );
  XNOR2_X1 U12007 ( .A(n9619), .B(n9617), .ZN(n10568) );
  INV_X1 U12008 ( .A(n9617), .ZN(n9618) );
  XNOR2_X1 U12009 ( .A(n11227), .B(n9716), .ZN(n10727) );
  AND2_X1 U12010 ( .A1(n13190), .A2(n12891), .ZN(n10728) );
  NAND2_X1 U12011 ( .A1(n11084), .A2(n10728), .ZN(n9621) );
  XNOR2_X1 U12012 ( .A(n14829), .B(n9709), .ZN(n9623) );
  NAND2_X1 U12013 ( .A1(n13190), .A2(n12890), .ZN(n9622) );
  XNOR2_X1 U12014 ( .A(n9623), .B(n9622), .ZN(n11095) );
  AOI21_X1 U12015 ( .B1(n10726), .B2(n10727), .A(n11095), .ZN(n9620) );
  NAND2_X1 U12016 ( .A1(n9623), .A2(n9622), .ZN(n9624) );
  XNOR2_X1 U12017 ( .A(n14842), .B(n9716), .ZN(n9625) );
  AND2_X1 U12018 ( .A1(n13190), .A2(n12889), .ZN(n9626) );
  NAND2_X1 U12019 ( .A1(n9625), .A2(n9626), .ZN(n9629) );
  INV_X1 U12020 ( .A(n9625), .ZN(n11257) );
  INV_X1 U12021 ( .A(n9626), .ZN(n9627) );
  NAND2_X1 U12022 ( .A1(n11257), .A2(n9627), .ZN(n9628) );
  AND2_X1 U12023 ( .A1(n9629), .A2(n9628), .ZN(n11141) );
  XNOR2_X1 U12024 ( .A(n11253), .B(n9716), .ZN(n9630) );
  AND2_X1 U12025 ( .A1(n13190), .A2(n12888), .ZN(n9631) );
  NAND2_X1 U12026 ( .A1(n9630), .A2(n9631), .ZN(n9634) );
  INV_X1 U12027 ( .A(n9630), .ZN(n11436) );
  INV_X1 U12028 ( .A(n9631), .ZN(n9632) );
  NAND2_X1 U12029 ( .A1(n11436), .A2(n9632), .ZN(n9633) );
  AND2_X1 U12030 ( .A1(n9634), .A2(n9633), .ZN(n11254) );
  XNOR2_X1 U12031 ( .A(n13273), .B(n9716), .ZN(n9636) );
  NAND2_X1 U12032 ( .A1(n13190), .A2(n12887), .ZN(n9637) );
  XNOR2_X1 U12033 ( .A(n9636), .B(n9637), .ZN(n11446) );
  AND2_X1 U12034 ( .A1(n11446), .A2(n9634), .ZN(n9635) );
  INV_X1 U12035 ( .A(n9636), .ZN(n9638) );
  NAND2_X1 U12036 ( .A1(n9638), .A2(n9637), .ZN(n9639) );
  XNOR2_X1 U12037 ( .A(n9640), .B(n9716), .ZN(n11893) );
  AND2_X1 U12038 ( .A1(n13190), .A2(n12886), .ZN(n9641) );
  NAND2_X1 U12039 ( .A1(n11893), .A2(n9641), .ZN(n9646) );
  INV_X1 U12040 ( .A(n11893), .ZN(n9643) );
  INV_X1 U12041 ( .A(n9641), .ZN(n9642) );
  NAND2_X1 U12042 ( .A1(n9643), .A2(n9642), .ZN(n9644) );
  NAND2_X1 U12043 ( .A1(n9646), .A2(n9644), .ZN(n11448) );
  INV_X1 U12044 ( .A(n11448), .ZN(n9645) );
  XNOR2_X1 U12045 ( .A(n11730), .B(n9716), .ZN(n9648) );
  NAND2_X1 U12046 ( .A1(n13190), .A2(n12885), .ZN(n9649) );
  XNOR2_X1 U12047 ( .A(n9648), .B(n9649), .ZN(n11896) );
  INV_X1 U12048 ( .A(n9648), .ZN(n9650) );
  NAND2_X1 U12049 ( .A1(n9650), .A2(n9649), .ZN(n9651) );
  XNOR2_X1 U12050 ( .A(n13269), .B(n9716), .ZN(n9653) );
  AND2_X1 U12051 ( .A1(n13190), .A2(n12884), .ZN(n9652) );
  INV_X1 U12052 ( .A(n9653), .ZN(n9654) );
  XNOR2_X1 U12053 ( .A(n13262), .B(n9709), .ZN(n11827) );
  NAND2_X1 U12054 ( .A1(n13190), .A2(n12883), .ZN(n9656) );
  XNOR2_X1 U12055 ( .A(n11827), .B(n9656), .ZN(n11836) );
  NAND2_X1 U12056 ( .A1(n11827), .A2(n9656), .ZN(n9657) );
  NAND2_X1 U12057 ( .A1(n11833), .A2(n9657), .ZN(n9658) );
  XNOR2_X1 U12058 ( .A(n13258), .B(n9716), .ZN(n9659) );
  NAND2_X1 U12059 ( .A1(n13190), .A2(n13151), .ZN(n9660) );
  XNOR2_X1 U12060 ( .A(n9659), .B(n9660), .ZN(n11825) );
  INV_X1 U12061 ( .A(n9659), .ZN(n9661) );
  NAND2_X1 U12062 ( .A1(n9661), .A2(n9660), .ZN(n9662) );
  XNOR2_X1 U12063 ( .A(n13253), .B(n9716), .ZN(n9663) );
  AND2_X1 U12064 ( .A1(n13190), .A2(n12882), .ZN(n9664) );
  NAND2_X1 U12065 ( .A1(n9663), .A2(n9664), .ZN(n9668) );
  INV_X1 U12066 ( .A(n9663), .ZN(n12787) );
  INV_X1 U12067 ( .A(n9664), .ZN(n9665) );
  NAND2_X1 U12068 ( .A1(n12787), .A2(n9665), .ZN(n9666) );
  NAND2_X1 U12069 ( .A1(n9668), .A2(n9666), .ZN(n12859) );
  XNOR2_X1 U12070 ( .A(n13246), .B(n9716), .ZN(n9670) );
  NAND2_X1 U12071 ( .A1(n13154), .A2(n13190), .ZN(n9671) );
  XNOR2_X1 U12072 ( .A(n9670), .B(n9671), .ZN(n12795) );
  AND2_X1 U12073 ( .A1(n12795), .A2(n9668), .ZN(n9669) );
  INV_X1 U12074 ( .A(n9670), .ZN(n12834) );
  XNOR2_X1 U12075 ( .A(n13242), .B(n9716), .ZN(n9674) );
  NOR2_X1 U12076 ( .A1(n12797), .A2(n13136), .ZN(n9672) );
  XNOR2_X1 U12077 ( .A(n9674), .B(n9672), .ZN(n12832) );
  INV_X1 U12078 ( .A(n9672), .ZN(n9673) );
  NAND2_X1 U12079 ( .A1(n9674), .A2(n9673), .ZN(n9675) );
  XNOR2_X1 U12080 ( .A(n13236), .B(n9709), .ZN(n9677) );
  NAND2_X1 U12081 ( .A1(n13079), .A2(n13190), .ZN(n9678) );
  XNOR2_X1 U12082 ( .A(n9677), .B(n9678), .ZN(n12803) );
  INV_X1 U12083 ( .A(n9677), .ZN(n9680) );
  INV_X1 U12084 ( .A(n9678), .ZN(n9679) );
  NAND2_X1 U12085 ( .A1(n9680), .A2(n9679), .ZN(n9681) );
  NAND2_X1 U12086 ( .A1(n12800), .A2(n9681), .ZN(n9685) );
  XNOR2_X1 U12087 ( .A(n13085), .B(n9716), .ZN(n9683) );
  XNOR2_X1 U12088 ( .A(n9685), .B(n9683), .ZN(n12842) );
  NOR2_X1 U12089 ( .A1(n13066), .A2(n13136), .ZN(n9682) );
  NAND2_X1 U12090 ( .A1(n12842), .A2(n9682), .ZN(n12843) );
  INV_X1 U12091 ( .A(n9683), .ZN(n9684) );
  NAND2_X1 U12092 ( .A1(n9685), .A2(n9684), .ZN(n9686) );
  XNOR2_X1 U12093 ( .A(n13074), .B(n9716), .ZN(n9687) );
  XNOR2_X1 U12094 ( .A(n9689), .B(n9687), .ZN(n12776) );
  NAND2_X1 U12095 ( .A1(n13080), .A2(n13190), .ZN(n12775) );
  NAND2_X1 U12096 ( .A1(n12776), .A2(n12775), .ZN(n9691) );
  INV_X1 U12097 ( .A(n9687), .ZN(n9688) );
  OR2_X1 U12098 ( .A1(n9689), .A2(n9688), .ZN(n9690) );
  NAND2_X1 U12099 ( .A1(n9691), .A2(n9690), .ZN(n12820) );
  XNOR2_X1 U12100 ( .A(n13219), .B(n9709), .ZN(n9692) );
  NOR2_X1 U12101 ( .A1(n13068), .A2(n13136), .ZN(n9693) );
  NAND2_X1 U12102 ( .A1(n9692), .A2(n9693), .ZN(n9696) );
  INV_X1 U12103 ( .A(n9692), .ZN(n12810) );
  INV_X1 U12104 ( .A(n9693), .ZN(n9694) );
  NAND2_X1 U12105 ( .A1(n12810), .A2(n9694), .ZN(n9695) );
  NAND2_X1 U12106 ( .A1(n9696), .A2(n9695), .ZN(n12819) );
  OR2_X2 U12107 ( .A1(n12820), .A2(n12819), .ZN(n12807) );
  NAND2_X1 U12108 ( .A1(n12807), .A2(n9696), .ZN(n9702) );
  XNOR2_X1 U12109 ( .A(n13038), .B(n9709), .ZN(n9698) );
  NOR2_X1 U12110 ( .A1(n9697), .A2(n13136), .ZN(n9699) );
  NAND2_X1 U12111 ( .A1(n9698), .A2(n9699), .ZN(n9703) );
  INV_X1 U12112 ( .A(n9698), .ZN(n12873) );
  INV_X1 U12113 ( .A(n9699), .ZN(n9700) );
  NAND2_X1 U12114 ( .A1(n12873), .A2(n9700), .ZN(n9701) );
  XNOR2_X1 U12115 ( .A(n13028), .B(n9716), .ZN(n9707) );
  NOR2_X1 U12116 ( .A1(n12814), .A2(n13136), .ZN(n9705) );
  XNOR2_X1 U12117 ( .A(n9707), .B(n9705), .ZN(n12874) );
  AND2_X1 U12118 ( .A1(n12874), .A2(n9703), .ZN(n9704) );
  INV_X1 U12119 ( .A(n9705), .ZN(n9706) );
  NAND2_X1 U12120 ( .A1(n9707), .A2(n9706), .ZN(n9708) );
  XNOR2_X1 U12121 ( .A(n13007), .B(n9709), .ZN(n9710) );
  NOR2_X1 U12122 ( .A1(n12958), .A2(n13136), .ZN(n9711) );
  NAND2_X1 U12123 ( .A1(n9710), .A2(n9711), .ZN(n9715) );
  INV_X1 U12124 ( .A(n9710), .ZN(n9713) );
  INV_X1 U12125 ( .A(n9711), .ZN(n9712) );
  NAND2_X1 U12126 ( .A1(n9713), .A2(n9712), .ZN(n9714) );
  NAND2_X1 U12127 ( .A1(n9715), .A2(n9714), .ZN(n12766) );
  XNOR2_X1 U12128 ( .A(n13202), .B(n9716), .ZN(n9717) );
  INV_X1 U12129 ( .A(n9719), .ZN(n9864) );
  AND2_X1 U12130 ( .A1(n14852), .A2(n9864), .ZN(n9720) );
  NAND2_X1 U12131 ( .A1(n12961), .A2(n12841), .ZN(n9739) );
  OAI21_X1 U12132 ( .B1(n12977), .B2(n13136), .A(n12865), .ZN(n9721) );
  AND2_X1 U12133 ( .A1(n14772), .A2(n9723), .ZN(n10824) );
  NAND2_X1 U12134 ( .A1(n9734), .A2(n10824), .ZN(n9725) );
  INV_X1 U12135 ( .A(n9726), .ZN(n9724) );
  NAND2_X1 U12136 ( .A1(n9727), .A2(n9726), .ZN(n9731) );
  AND2_X1 U12137 ( .A1(n9729), .A2(n9728), .ZN(n9730) );
  NAND2_X1 U12138 ( .A1(n9731), .A2(n9730), .ZN(n10422) );
  OAI22_X1 U12139 ( .A1(n12996), .A2(n12856), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9732), .ZN(n9737) );
  NAND2_X1 U12140 ( .A1(n9734), .A2(n9733), .ZN(n12828) );
  OR2_X1 U12141 ( .A1(n12828), .A2(n13067), .ZN(n12847) );
  OAI22_X1 U12142 ( .A1(n9735), .A2(n12869), .B1(n12958), .B2(n12847), .ZN(
        n9736) );
  AOI211_X1 U12143 ( .C1(n12995), .C2(n12871), .A(n9737), .B(n9736), .ZN(n9738) );
  INV_X1 U12144 ( .A(n9740), .ZN(n9741) );
  NOR2_X1 U12145 ( .A1(n9863), .A2(n9741), .ZN(n9742) );
  NAND2_X1 U12146 ( .A1(n11432), .A2(n9742), .ZN(n9866) );
  NOR2_X1 U12147 ( .A1(P2_U3088), .A2(n9866), .ZN(P2_U3947) );
  INV_X1 U12148 ( .A(n9743), .ZN(n10170) );
  OR2_X2 U12149 ( .A1(n10170), .A2(n12751), .ZN(n12333) );
  INV_X1 U12150 ( .A(n12333), .ZN(P3_U3897) );
  AND2_X2 U12151 ( .A1(n9800), .A2(n10042), .ZN(P1_U4016) );
  NOR2_X1 U12152 ( .A1(n6459), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13299) );
  INV_X2 U12153 ( .A(n13299), .ZN(n13314) );
  AND2_X1 U12154 ( .A1(n6459), .A2(P2_U3088), .ZN(n13306) );
  OAI222_X1 U12155 ( .A1(n13314), .A2(n9744), .B1(n6452), .B2(n9751), .C1(
        P2_U3088), .C2(n9879), .ZN(P2_U3326) );
  AOI22_X1 U12156 ( .A1(n13299), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n9919), 
        .B2(P2_STATE_REG_SCAN_IN), .ZN(n9745) );
  OAI21_X1 U12157 ( .B1(n9747), .B2(n6452), .A(n9745), .ZN(P2_U3325) );
  AND2_X1 U12158 ( .A1(n6459), .A2(P1_U3086), .ZN(n14081) );
  INV_X2 U12159 ( .A(n14081), .ZN(n14085) );
  INV_X1 U12160 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9748) );
  NAND2_X1 U12161 ( .A1(n7433), .A2(P1_U3086), .ZN(n14083) );
  INV_X1 U12162 ( .A(n13619), .ZN(n9746) );
  OAI222_X1 U12163 ( .A1(n14085), .A2(n9748), .B1(n14083), .B2(n9747), .C1(
        P1_U3086), .C2(n9746), .ZN(P1_U3353) );
  AOI22_X1 U12164 ( .A1(n14608), .A2(P2_STATE_REG_SCAN_IN), .B1(n13299), .B2(
        P1_DATAO_REG_3__SCAN_IN), .ZN(n9749) );
  OAI21_X1 U12165 ( .B1(n9754), .B2(n6452), .A(n9749), .ZN(P2_U3324) );
  INV_X1 U12166 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9752) );
  CLKBUF_X1 U12167 ( .A(n14083), .Z(n14088) );
  INV_X1 U12168 ( .A(n13602), .ZN(n9750) );
  OAI222_X1 U12169 ( .A1(n14085), .A2(n9752), .B1(n14088), .B2(n9751), .C1(
        P1_U3086), .C2(n9750), .ZN(P1_U3354) );
  INV_X1 U12170 ( .A(n13631), .ZN(n9753) );
  OAI222_X1 U12171 ( .A1(n14085), .A2(n9755), .B1(n14083), .B2(n9754), .C1(
        P1_U3086), .C2(n9753), .ZN(P1_U3352) );
  NAND2_X1 U12172 ( .A1(n6459), .A2(P3_U3151), .ZN(n14213) );
  NOR2_X2 U12173 ( .A1(n6459), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14223) );
  INV_X1 U12174 ( .A(n14223), .ZN(n14215) );
  OAI222_X1 U12175 ( .A1(P3_U3151), .A2(n10762), .B1(n14213), .B2(n9757), .C1(
        n14215), .C2(n9756), .ZN(P3_U3287) );
  OAI222_X1 U12176 ( .A1(n14215), .A2(n9759), .B1(n14213), .B2(n9758), .C1(
        P3_U3151), .C2(n6614), .ZN(P3_U3294) );
  OAI222_X1 U12177 ( .A1(P3_U3151), .A2(n10334), .B1(n14215), .B2(n9761), .C1(
        n9760), .C2(n14213), .ZN(P3_U3289) );
  OAI222_X1 U12178 ( .A1(P3_U3151), .A2(n10204), .B1(n14215), .B2(n9763), .C1(
        n9762), .C2(n14213), .ZN(P3_U3295) );
  INV_X1 U12179 ( .A(n9764), .ZN(n9766) );
  OAI222_X1 U12180 ( .A1(n14085), .A2(n9765), .B1(n14083), .B2(n9766), .C1(
        P1_U3086), .C2(n13643), .ZN(P1_U3351) );
  OAI222_X1 U12181 ( .A1(n13314), .A2(n9767), .B1(n6452), .B2(n9766), .C1(
        P2_U3088), .C2(n9902), .ZN(P2_U3323) );
  INV_X1 U12182 ( .A(n14213), .ZN(n14222) );
  AOI222_X1 U12183 ( .A1(n9768), .A2(n14223), .B1(SI_10_), .B2(n14222), .C1(
        n10965), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9769) );
  INV_X1 U12184 ( .A(n9769), .ZN(P3_U3285) );
  AOI222_X1 U12185 ( .A1(n9770), .A2(n14223), .B1(SI_7_), .B2(n14222), .C1(
        n10645), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9771) );
  INV_X1 U12186 ( .A(n9771), .ZN(P3_U3288) );
  AOI222_X1 U12187 ( .A1(n9772), .A2(n14223), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10450), .C1(SI_4_), .C2(n14222), .ZN(n9773) );
  INV_X1 U12188 ( .A(n9773), .ZN(P3_U3291) );
  AOI222_X1 U12189 ( .A1(n9774), .A2(n14223), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10385), .C1(SI_5_), .C2(n14222), .ZN(n9775) );
  INV_X1 U12190 ( .A(n9775), .ZN(P3_U3290) );
  AOI222_X1 U12191 ( .A1(n9776), .A2(n14223), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10359), .C1(SI_2_), .C2(n14222), .ZN(n9777) );
  INV_X1 U12192 ( .A(n9777), .ZN(P3_U3293) );
  AOI222_X1 U12193 ( .A1(n9778), .A2(n14223), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10317), .C1(SI_3_), .C2(n14222), .ZN(n9779) );
  INV_X1 U12194 ( .A(n9779), .ZN(P3_U3292) );
  INV_X1 U12195 ( .A(n9780), .ZN(n9782) );
  OAI222_X1 U12196 ( .A1(n13314), .A2(n9781), .B1(n6452), .B2(n9782), .C1(
        P2_U3088), .C2(n10011), .ZN(P2_U3322) );
  OAI222_X1 U12197 ( .A1(n14085), .A2(n9783), .B1(n14083), .B2(n9782), .C1(
        P1_U3086), .C2(n9977), .ZN(P1_U3350) );
  OAI222_X1 U12198 ( .A1(P3_U3151), .A2(n12383), .B1(n14213), .B2(n15162), 
        .C1(n14215), .C2(n9784), .ZN(P3_U3283) );
  INV_X1 U12199 ( .A(n9785), .ZN(n9787) );
  OAI222_X1 U12200 ( .A1(n14085), .A2(n9786), .B1(n14083), .B2(n9787), .C1(
        P1_U3086), .C2(n13658), .ZN(P1_U3349) );
  OAI222_X1 U12201 ( .A1(n13314), .A2(n9788), .B1(n6452), .B2(n9787), .C1(
        P2_U3088), .C2(n14619), .ZN(P2_U3321) );
  INV_X1 U12202 ( .A(n9789), .ZN(n9791) );
  OAI222_X1 U12203 ( .A1(n13314), .A2(n9790), .B1(n6452), .B2(n9791), .C1(
        P2_U3088), .C2(n14632), .ZN(P2_U3320) );
  OAI222_X1 U12204 ( .A1(n14085), .A2(n9792), .B1(n14083), .B2(n9791), .C1(
        P1_U3086), .C2(n13671), .ZN(P1_U3348) );
  INV_X1 U12205 ( .A(n10042), .ZN(n10038) );
  NAND2_X1 U12206 ( .A1(n9800), .A2(n10038), .ZN(n10068) );
  NAND3_X1 U12207 ( .A1(n11501), .A2(P1_B_REG_SCAN_IN), .A3(n11430), .ZN(n9793) );
  OAI211_X1 U12208 ( .C1(P1_B_REG_SCAN_IN), .C2(n11430), .A(n11627), .B(n9793), 
        .ZN(n10061) );
  INV_X1 U12209 ( .A(n10061), .ZN(n9794) );
  INV_X1 U12210 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9797) );
  INV_X1 U12211 ( .A(n11501), .ZN(n9795) );
  OR2_X1 U12212 ( .A1(n9795), .A2(n11627), .ZN(n10062) );
  INV_X1 U12213 ( .A(n10062), .ZN(n9796) );
  AOI22_X1 U12214 ( .A1(n14546), .A2(n9797), .B1(n9800), .B2(n9796), .ZN(
        P1_U3446) );
  INV_X1 U12215 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9801) );
  INV_X1 U12216 ( .A(n11430), .ZN(n9798) );
  OR2_X1 U12217 ( .A1(n9798), .A2(n11627), .ZN(n10048) );
  INV_X1 U12218 ( .A(n10048), .ZN(n9799) );
  AOI22_X1 U12219 ( .A1(n14546), .A2(n9801), .B1(n9800), .B2(n9799), .ZN(
        P1_U3445) );
  NOR2_X1 U12220 ( .A1(n12751), .A2(n9802), .ZN(n9807) );
  INV_X1 U12221 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9803) );
  NOR2_X1 U12222 ( .A1(n9830), .A2(n9803), .ZN(P3_U3238) );
  INV_X1 U12223 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9804) );
  NOR2_X1 U12224 ( .A1(n9807), .A2(n9804), .ZN(P3_U3239) );
  INV_X1 U12225 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9805) );
  NOR2_X1 U12226 ( .A1(n9807), .A2(n9805), .ZN(P3_U3244) );
  INV_X1 U12227 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9806) );
  NOR2_X1 U12228 ( .A1(n9807), .A2(n9806), .ZN(P3_U3245) );
  INV_X1 U12229 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9808) );
  NOR2_X1 U12230 ( .A1(n9830), .A2(n9808), .ZN(P3_U3246) );
  INV_X1 U12231 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9809) );
  NOR2_X1 U12232 ( .A1(n9830), .A2(n9809), .ZN(P3_U3247) );
  INV_X1 U12233 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9810) );
  NOR2_X1 U12234 ( .A1(n9807), .A2(n9810), .ZN(P3_U3240) );
  INV_X1 U12235 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9811) );
  NOR2_X1 U12236 ( .A1(n9807), .A2(n9811), .ZN(P3_U3241) );
  INV_X1 U12237 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9812) );
  NOR2_X1 U12238 ( .A1(n9807), .A2(n9812), .ZN(P3_U3242) );
  INV_X1 U12239 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9813) );
  NOR2_X1 U12240 ( .A1(n9807), .A2(n9813), .ZN(P3_U3234) );
  INV_X1 U12241 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9814) );
  NOR2_X1 U12242 ( .A1(n9807), .A2(n9814), .ZN(P3_U3235) );
  INV_X1 U12243 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9815) );
  NOR2_X1 U12244 ( .A1(n9807), .A2(n9815), .ZN(P3_U3236) );
  INV_X1 U12245 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9816) );
  NOR2_X1 U12246 ( .A1(n9807), .A2(n9816), .ZN(P3_U3237) );
  INV_X1 U12247 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9817) );
  NOR2_X1 U12248 ( .A1(n9830), .A2(n9817), .ZN(P3_U3254) );
  INV_X1 U12249 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n15161) );
  NOR2_X1 U12250 ( .A1(n9830), .A2(n15161), .ZN(P3_U3255) );
  INV_X1 U12251 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n15084) );
  NOR2_X1 U12252 ( .A1(n9830), .A2(n15084), .ZN(P3_U3256) );
  INV_X1 U12253 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9818) );
  NOR2_X1 U12254 ( .A1(n9830), .A2(n9818), .ZN(P3_U3257) );
  INV_X1 U12255 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9819) );
  NOR2_X1 U12256 ( .A1(n9807), .A2(n9819), .ZN(P3_U3258) );
  INV_X1 U12257 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9820) );
  NOR2_X1 U12258 ( .A1(n9830), .A2(n9820), .ZN(P3_U3259) );
  INV_X1 U12259 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9821) );
  NOR2_X1 U12260 ( .A1(n9830), .A2(n9821), .ZN(P3_U3260) );
  INV_X1 U12261 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9822) );
  NOR2_X1 U12262 ( .A1(n9830), .A2(n9822), .ZN(P3_U3261) );
  INV_X1 U12263 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9823) );
  NOR2_X1 U12264 ( .A1(n9830), .A2(n9823), .ZN(P3_U3262) );
  INV_X1 U12265 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n15096) );
  NOR2_X1 U12266 ( .A1(n9830), .A2(n15096), .ZN(P3_U3248) );
  INV_X1 U12267 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9824) );
  NOR2_X1 U12268 ( .A1(n9830), .A2(n9824), .ZN(P3_U3249) );
  INV_X1 U12269 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9825) );
  NOR2_X1 U12270 ( .A1(n9830), .A2(n9825), .ZN(P3_U3250) );
  INV_X1 U12271 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9826) );
  NOR2_X1 U12272 ( .A1(n9830), .A2(n9826), .ZN(P3_U3251) );
  INV_X1 U12273 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9827) );
  NOR2_X1 U12274 ( .A1(n9830), .A2(n9827), .ZN(P3_U3263) );
  INV_X1 U12275 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9828) );
  NOR2_X1 U12276 ( .A1(n9830), .A2(n9828), .ZN(P3_U3252) );
  INV_X1 U12277 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9829) );
  NOR2_X1 U12278 ( .A1(n9830), .A2(n9829), .ZN(P3_U3253) );
  INV_X1 U12279 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9831) );
  NOR2_X1 U12280 ( .A1(n9830), .A2(n9831), .ZN(P3_U3243) );
  NAND2_X1 U12281 ( .A1(n10068), .A2(n11344), .ZN(n9842) );
  NAND2_X1 U12282 ( .A1(n9833), .A2(n9832), .ZN(n9835) );
  NAND2_X1 U12283 ( .A1(n9835), .A2(n9834), .ZN(n9840) );
  NAND2_X1 U12284 ( .A1(n9842), .A2(n9840), .ZN(n14492) );
  INV_X1 U12285 ( .A(n14492), .ZN(n13642) );
  NOR2_X1 U12286 ( .A1(n13642), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12287 ( .A(n9836), .ZN(n9838) );
  OAI222_X1 U12288 ( .A1(n13314), .A2(n9837), .B1(n6452), .B2(n9838), .C1(
        P2_U3088), .C2(n14645), .ZN(P2_U3319) );
  OAI222_X1 U12289 ( .A1(n14085), .A2(n9839), .B1(n14083), .B2(n9838), .C1(
        P1_U3086), .C2(n9965), .ZN(P1_U3347) );
  INV_X1 U12290 ( .A(n9840), .ZN(n9841) );
  NAND2_X1 U12291 ( .A1(n9842), .A2(n9841), .ZN(n9956) );
  INV_X1 U12292 ( .A(n9956), .ZN(n9943) );
  AOI21_X1 U12293 ( .B1(n9942), .B2(n8057), .A(n8685), .ZN(n13616) );
  OAI21_X1 U12294 ( .B1(n9942), .B2(P1_REG1_REG_0__SCAN_IN), .A(n13616), .ZN(
        n9843) );
  XNOR2_X1 U12295 ( .A(n9843), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9844) );
  AOI22_X1 U12296 ( .A1(n9943), .A2(n9844), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9845) );
  OAI21_X1 U12297 ( .B1(n14492), .B2(n6686), .A(n9845), .ZN(P1_U3243) );
  INV_X1 U12298 ( .A(n9846), .ZN(n9848) );
  OAI222_X1 U12299 ( .A1(n14085), .A2(n9847), .B1(n14083), .B2(n9848), .C1(
        P1_U3086), .C2(n9989), .ZN(P1_U3346) );
  OAI222_X1 U12300 ( .A1(n13314), .A2(n9849), .B1(n6452), .B2(n9848), .C1(
        P2_U3088), .C2(n10083), .ZN(P2_U3318) );
  OAI222_X1 U12301 ( .A1(P3_U3151), .A2(n14916), .B1(n14213), .B2(n15157), 
        .C1(n14215), .C2(n9850), .ZN(P3_U3282) );
  INV_X1 U12302 ( .A(n9851), .ZN(n9854) );
  OAI222_X1 U12303 ( .A1(n14085), .A2(n9852), .B1(n14083), .B2(n9854), .C1(
        P1_U3086), .C2(n13688), .ZN(P1_U3345) );
  INV_X1 U12304 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9855) );
  INV_X1 U12305 ( .A(n10102), .ZN(n9853) );
  OAI222_X1 U12306 ( .A1(n13314), .A2(n9855), .B1(n6452), .B2(n9854), .C1(
        P2_U3088), .C2(n9853), .ZN(P2_U3317) );
  NAND2_X1 U12307 ( .A1(n12333), .A2(P3_DATAO_REG_17__SCAN_IN), .ZN(n9856) );
  OAI21_X1 U12308 ( .B1(n12056), .B2(n12333), .A(n9856), .ZN(P3_U3508) );
  INV_X1 U12309 ( .A(n9857), .ZN(n9860) );
  OAI222_X1 U12310 ( .A1(n14085), .A2(n9858), .B1(n14083), .B2(n9860), .C1(
        P1_U3086), .C2(n10192), .ZN(P1_U3344) );
  INV_X1 U12311 ( .A(n12903), .ZN(n9859) );
  OAI222_X1 U12312 ( .A1(n13314), .A2(n9861), .B1(n6452), .B2(n9860), .C1(
        P2_U3088), .C2(n9859), .ZN(P2_U3316) );
  OAI21_X1 U12313 ( .B1(n9864), .B2(n9863), .A(n9862), .ZN(n9865) );
  NAND2_X1 U12314 ( .A1(n9866), .A2(n9865), .ZN(n9887) );
  NOR2_X1 U12315 ( .A1(n9873), .A2(P2_U3088), .ZN(n9867) );
  INV_X1 U12316 ( .A(n14728), .ZN(n14659) );
  INV_X1 U12317 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15197) );
  XNOR2_X1 U12318 ( .A(n10011), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n9876) );
  XNOR2_X1 U12319 ( .A(n9879), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n9911) );
  AND2_X1 U12320 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9910) );
  NAND2_X1 U12321 ( .A1(n9911), .A2(n9910), .ZN(n9909) );
  NAND2_X1 U12322 ( .A1(n9908), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9868) );
  NAND2_X1 U12323 ( .A1(n9909), .A2(n9868), .ZN(n9921) );
  INV_X1 U12324 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10873) );
  XNOR2_X1 U12325 ( .A(n9919), .B(n10873), .ZN(n9922) );
  NAND2_X1 U12326 ( .A1(n9921), .A2(n9922), .ZN(n9920) );
  NAND2_X1 U12327 ( .A1(n9919), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9869) );
  NAND2_X1 U12328 ( .A1(n9920), .A2(n9869), .ZN(n14600) );
  INV_X1 U12329 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10818) );
  XNOR2_X1 U12330 ( .A(n14608), .B(n10818), .ZN(n14601) );
  NAND2_X1 U12331 ( .A1(n14600), .A2(n14601), .ZN(n14599) );
  NAND2_X1 U12332 ( .A1(n14608), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9870) );
  NAND2_X1 U12333 ( .A1(n14599), .A2(n9870), .ZN(n9893) );
  XNOR2_X1 U12334 ( .A(n9902), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n9894) );
  NAND2_X1 U12335 ( .A1(n9893), .A2(n9894), .ZN(n9892) );
  INV_X1 U12336 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9871) );
  OR2_X1 U12337 ( .A1(n9902), .A2(n9871), .ZN(n9872) );
  NAND2_X1 U12338 ( .A1(n9892), .A2(n9872), .ZN(n9875) );
  NAND2_X1 U12339 ( .A1(n9873), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13308) );
  NOR2_X1 U12340 ( .A1(n13308), .A2(n13311), .ZN(n9874) );
  NAND2_X1 U12341 ( .A1(n9875), .A2(n9876), .ZN(n10013) );
  OAI211_X1 U12342 ( .C1(n9876), .C2(n9875), .A(n14724), .B(n10013), .ZN(n9877) );
  NAND2_X1 U12343 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10689) );
  OAI211_X1 U12344 ( .C1(n15197), .C2(n14731), .A(n9877), .B(n10689), .ZN(
        n9878) );
  INV_X1 U12345 ( .A(n9878), .ZN(n9891) );
  XNOR2_X1 U12346 ( .A(n10011), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n9889) );
  XNOR2_X1 U12347 ( .A(n9879), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n9905) );
  AND2_X1 U12348 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9904) );
  NAND2_X1 U12349 ( .A1(n9905), .A2(n9904), .ZN(n9903) );
  NAND2_X1 U12350 ( .A1(n9908), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9880) );
  NAND2_X1 U12351 ( .A1(n9903), .A2(n9880), .ZN(n9915) );
  XNOR2_X1 U12352 ( .A(n9919), .B(n7739), .ZN(n9916) );
  NAND2_X1 U12353 ( .A1(n9915), .A2(n9916), .ZN(n9914) );
  NAND2_X1 U12354 ( .A1(n9919), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9881) );
  NAND2_X1 U12355 ( .A1(n9914), .A2(n9881), .ZN(n14603) );
  INV_X1 U12356 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9882) );
  XNOR2_X1 U12357 ( .A(n14608), .B(n9882), .ZN(n14604) );
  NAND2_X1 U12358 ( .A1(n14603), .A2(n14604), .ZN(n14602) );
  NAND2_X1 U12359 ( .A1(n14608), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9883) );
  NAND2_X1 U12360 ( .A1(n14602), .A2(n9883), .ZN(n9898) );
  XNOR2_X1 U12361 ( .A(n9902), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n9899) );
  NAND2_X1 U12362 ( .A1(n9898), .A2(n9899), .ZN(n9897) );
  INV_X1 U12363 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9884) );
  OR2_X1 U12364 ( .A1(n9902), .A2(n9884), .ZN(n9885) );
  NAND2_X1 U12365 ( .A1(n9897), .A2(n9885), .ZN(n9888) );
  NOR2_X1 U12366 ( .A1(n13308), .A2(n12949), .ZN(n9886) );
  AND2_X1 U12367 ( .A1(n9887), .A2(n9886), .ZN(n14657) );
  NAND2_X1 U12368 ( .A1(n9888), .A2(n9889), .ZN(n10002) );
  OAI211_X1 U12369 ( .C1(n9889), .C2(n9888), .A(n14657), .B(n10002), .ZN(n9890) );
  OAI211_X1 U12370 ( .C1(n14659), .C2(n10011), .A(n9891), .B(n9890), .ZN(
        P2_U3219) );
  INV_X1 U12371 ( .A(n14731), .ZN(n14598) );
  OAI211_X1 U12372 ( .C1(n9894), .C2(n9893), .A(n14724), .B(n9892), .ZN(n9895)
         );
  NAND2_X1 U12373 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10671) );
  NAND2_X1 U12374 ( .A1(n9895), .A2(n10671), .ZN(n9896) );
  AOI21_X1 U12375 ( .B1(n14598), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n9896), .ZN(
        n9901) );
  OAI211_X1 U12376 ( .C1(n9899), .C2(n9898), .A(n14657), .B(n9897), .ZN(n9900)
         );
  OAI211_X1 U12377 ( .C1(n14659), .C2(n9902), .A(n9901), .B(n9900), .ZN(
        P2_U3218) );
  INV_X1 U12378 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10885) );
  OAI211_X1 U12379 ( .C1(n9905), .C2(n9904), .A(n14657), .B(n9903), .ZN(n9906)
         );
  OAI21_X1 U12380 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n10885), .A(n9906), .ZN(
        n9907) );
  AOI21_X1 U12381 ( .B1(n9908), .B2(n14728), .A(n9907), .ZN(n9913) );
  OAI211_X1 U12382 ( .C1(n9911), .C2(n9910), .A(n14724), .B(n9909), .ZN(n9912)
         );
  OAI211_X1 U12383 ( .C1(n6685), .C2(n14731), .A(n9913), .B(n9912), .ZN(
        P2_U3215) );
  INV_X1 U12384 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15154) );
  OAI211_X1 U12385 ( .C1(n9916), .C2(n9915), .A(n14657), .B(n9914), .ZN(n9917)
         );
  OAI21_X1 U12386 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7738), .A(n9917), .ZN(
        n9918) );
  AOI21_X1 U12387 ( .B1(n9919), .B2(n14728), .A(n9918), .ZN(n9924) );
  OAI211_X1 U12388 ( .C1(n9922), .C2(n9921), .A(n14724), .B(n9920), .ZN(n9923)
         );
  OAI211_X1 U12389 ( .C1(n15154), .C2(n14731), .A(n9924), .B(n9923), .ZN(
        P2_U3216) );
  INV_X1 U12390 ( .A(n9925), .ZN(n9928) );
  OAI222_X1 U12391 ( .A1(n13314), .A2(n9926), .B1(n6452), .B2(n9928), .C1(
        n12928), .C2(P2_U3088), .ZN(P2_U3315) );
  OAI222_X1 U12392 ( .A1(P1_U3086), .A2(n13710), .B1(n14088), .B2(n9928), .C1(
        n9927), .C2(n14085), .ZN(P1_U3343) );
  MUX2_X1 U12393 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10187), .S(n10192), .Z(
        n9941) );
  INV_X1 U12394 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9939) );
  INV_X1 U12395 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9936) );
  INV_X1 U12396 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9933) );
  MUX2_X1 U12397 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n8072), .S(n13602), .Z(
        n13605) );
  AND2_X1 U12398 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n13604) );
  NAND2_X1 U12399 ( .A1(n13605), .A2(n13604), .ZN(n13603) );
  NAND2_X1 U12400 ( .A1(n13602), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9929) );
  NAND2_X1 U12401 ( .A1(n13603), .A2(n9929), .ZN(n13624) );
  MUX2_X1 U12402 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n8109), .S(n13619), .Z(
        n13625) );
  NAND2_X1 U12403 ( .A1(n13624), .A2(n13625), .ZN(n13623) );
  NAND2_X1 U12404 ( .A1(n13619), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9930) );
  NAND2_X1 U12405 ( .A1(n13623), .A2(n9930), .ZN(n13636) );
  XNOR2_X1 U12406 ( .A(n13631), .B(n9931), .ZN(n13637) );
  NAND2_X1 U12407 ( .A1(n13636), .A2(n13637), .ZN(n13635) );
  NAND2_X1 U12408 ( .A1(n13631), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9932) );
  NAND2_X1 U12409 ( .A1(n13635), .A2(n9932), .ZN(n13646) );
  XNOR2_X1 U12410 ( .A(n13643), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n13647) );
  NAND2_X1 U12411 ( .A1(n13646), .A2(n13647), .ZN(n13645) );
  OAI21_X1 U12412 ( .B1(n9933), .B2(n13643), .A(n13645), .ZN(n9975) );
  MUX2_X1 U12413 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9934), .S(n9977), .Z(n9976)
         );
  AOI21_X1 U12414 ( .B1(n9977), .B2(n9934), .A(n9974), .ZN(n13663) );
  XNOR2_X1 U12415 ( .A(n13658), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n13664) );
  NAND2_X1 U12416 ( .A1(n13663), .A2(n13664), .ZN(n13662) );
  OAI21_X1 U12417 ( .B1(n13658), .B2(n9935), .A(n13662), .ZN(n13680) );
  MUX2_X1 U12418 ( .A(n9936), .B(P1_REG1_REG_7__SCAN_IN), .S(n13671), .Z(
        n13681) );
  NAND2_X1 U12419 ( .A1(n13680), .A2(n13681), .ZN(n13679) );
  OAI21_X1 U12420 ( .B1(n13671), .B2(n9936), .A(n13679), .ZN(n9963) );
  MUX2_X1 U12421 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9937), .S(n9965), .Z(n9964)
         );
  AOI21_X1 U12422 ( .B1(n9965), .B2(n9937), .A(n9962), .ZN(n9987) );
  MUX2_X1 U12423 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9938), .S(n9989), .Z(n9988)
         );
  AOI21_X1 U12424 ( .B1(n9938), .B2(n9989), .A(n9986), .ZN(n13687) );
  MUX2_X1 U12425 ( .A(n9939), .B(P1_REG1_REG_10__SCAN_IN), .S(n13688), .Z(
        n13686) );
  NAND2_X1 U12426 ( .A1(n13687), .A2(n13686), .ZN(n13685) );
  OAI21_X1 U12427 ( .B1(n13688), .B2(n9939), .A(n13685), .ZN(n9940) );
  AOI21_X1 U12428 ( .B1(n9941), .B2(n9940), .A(n10186), .ZN(n9961) );
  INV_X1 U12429 ( .A(n10192), .ZN(n9946) );
  AND2_X1 U12430 ( .A1(n9943), .A2(n8685), .ZN(n14489) );
  INV_X1 U12431 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14112) );
  NAND2_X1 U12432 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9944) );
  OAI21_X1 U12433 ( .B1(n14492), .B2(n14112), .A(n9944), .ZN(n9945) );
  AOI21_X1 U12434 ( .B1(n9946), .B2(n14489), .A(n9945), .ZN(n9960) );
  MUX2_X1 U12435 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n8073), .S(n13602), .Z(
        n13607) );
  AND2_X1 U12436 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13612) );
  NAND2_X1 U12437 ( .A1(n13607), .A2(n13612), .ZN(n13606) );
  NAND2_X1 U12438 ( .A1(n13602), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9947) );
  NAND2_X1 U12439 ( .A1(n13606), .A2(n9947), .ZN(n13621) );
  MUX2_X1 U12440 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n8108), .S(n13619), .Z(
        n13622) );
  NAND2_X1 U12441 ( .A1(n13621), .A2(n13622), .ZN(n13620) );
  NAND2_X1 U12442 ( .A1(n13619), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U12443 ( .A1(n13620), .A2(n9948), .ZN(n13633) );
  INV_X1 U12444 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9949) );
  XNOR2_X1 U12445 ( .A(n13631), .B(n9949), .ZN(n13634) );
  NAND2_X1 U12446 ( .A1(n13633), .A2(n13634), .ZN(n13632) );
  NAND2_X1 U12447 ( .A1(n13631), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9950) );
  NAND2_X1 U12448 ( .A1(n13632), .A2(n9950), .ZN(n13652) );
  XNOR2_X1 U12449 ( .A(n13643), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n13653) );
  NAND2_X1 U12450 ( .A1(n13652), .A2(n13653), .ZN(n13651) );
  OAI21_X1 U12451 ( .B1(n11316), .B2(n13643), .A(n13651), .ZN(n9981) );
  MUX2_X1 U12452 ( .A(n9951), .B(P1_REG2_REG_5__SCAN_IN), .S(n9977), .Z(n9982)
         );
  NAND2_X1 U12453 ( .A1(n9981), .A2(n9982), .ZN(n9980) );
  OAI21_X1 U12454 ( .B1(n9951), .B2(n9977), .A(n9980), .ZN(n13666) );
  XNOR2_X1 U12455 ( .A(n13658), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n13667) );
  NAND2_X1 U12456 ( .A1(n13666), .A2(n13667), .ZN(n13665) );
  OAI21_X1 U12457 ( .B1(n13658), .B2(n9952), .A(n13665), .ZN(n13677) );
  MUX2_X1 U12458 ( .A(n9953), .B(P1_REG2_REG_7__SCAN_IN), .S(n13671), .Z(
        n13678) );
  NAND2_X1 U12459 ( .A1(n13677), .A2(n13678), .ZN(n13676) );
  OAI21_X1 U12460 ( .B1(n13671), .B2(n9953), .A(n13676), .ZN(n9969) );
  XNOR2_X1 U12461 ( .A(n9965), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n9970) );
  NAND2_X1 U12462 ( .A1(n9969), .A2(n9970), .ZN(n9968) );
  OAI21_X1 U12463 ( .B1(n11358), .B2(n9965), .A(n9968), .ZN(n9994) );
  MUX2_X1 U12464 ( .A(n9954), .B(P1_REG2_REG_9__SCAN_IN), .S(n9989), .Z(n9995)
         );
  NAND2_X1 U12465 ( .A1(n9994), .A2(n9995), .ZN(n9993) );
  OAI21_X1 U12466 ( .B1(n9989), .B2(n9954), .A(n9993), .ZN(n13694) );
  MUX2_X1 U12467 ( .A(n9955), .B(P1_REG2_REG_10__SCAN_IN), .S(n13688), .Z(
        n13693) );
  NAND2_X1 U12468 ( .A1(n13694), .A2(n13693), .ZN(n13692) );
  OAI21_X1 U12469 ( .B1(n13688), .B2(n9955), .A(n13692), .ZN(n9958) );
  XNOR2_X1 U12470 ( .A(n10192), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n9957) );
  NAND2_X1 U12471 ( .A1(n9958), .A2(n9957), .ZN(n10191) );
  OR3_X1 U12472 ( .A1(n9956), .A2(n8684), .A3(n8685), .ZN(n14478) );
  OAI211_X1 U12473 ( .C1(n9958), .C2(n9957), .A(n10191), .B(n14440), .ZN(n9959) );
  OAI211_X1 U12474 ( .C1(n9961), .C2(n14482), .A(n9960), .B(n9959), .ZN(
        P1_U3254) );
  AOI21_X1 U12475 ( .B1(n9964), .B2(n9963), .A(n9962), .ZN(n9973) );
  INV_X1 U12476 ( .A(n9965), .ZN(n9967) );
  INV_X1 U12477 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14107) );
  NAND2_X1 U12478 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11297) );
  OAI21_X1 U12479 ( .B1(n14492), .B2(n14107), .A(n11297), .ZN(n9966) );
  AOI21_X1 U12480 ( .B1(n9967), .B2(n14489), .A(n9966), .ZN(n9972) );
  OAI211_X1 U12481 ( .C1(n9970), .C2(n9969), .A(n14440), .B(n9968), .ZN(n9971)
         );
  OAI211_X1 U12482 ( .C1(n9973), .C2(n14482), .A(n9972), .B(n9971), .ZN(
        P1_U3251) );
  AOI21_X1 U12483 ( .B1(n9976), .B2(n9975), .A(n9974), .ZN(n9985) );
  INV_X1 U12484 ( .A(n9977), .ZN(n9979) );
  INV_X1 U12485 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14146) );
  NAND2_X1 U12486 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10611) );
  OAI21_X1 U12487 ( .B1(n14492), .B2(n14146), .A(n10611), .ZN(n9978) );
  AOI21_X1 U12488 ( .B1(n9979), .B2(n14489), .A(n9978), .ZN(n9984) );
  OAI211_X1 U12489 ( .C1(n9982), .C2(n9981), .A(n14440), .B(n9980), .ZN(n9983)
         );
  OAI211_X1 U12490 ( .C1(n9985), .C2(n14482), .A(n9984), .B(n9983), .ZN(
        P1_U3248) );
  AOI21_X1 U12491 ( .B1(n9988), .B2(n9987), .A(n9986), .ZN(n9998) );
  INV_X1 U12492 ( .A(n9989), .ZN(n9992) );
  INV_X1 U12493 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n15155) );
  NAND2_X1 U12494 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n9990) );
  OAI21_X1 U12495 ( .B1(n14492), .B2(n15155), .A(n9990), .ZN(n9991) );
  AOI21_X1 U12496 ( .B1(n9992), .B2(n14489), .A(n9991), .ZN(n9997) );
  OAI211_X1 U12497 ( .C1(n9995), .C2(n9994), .A(n14440), .B(n9993), .ZN(n9996)
         );
  OAI211_X1 U12498 ( .C1(n9998), .C2(n14482), .A(n9997), .B(n9996), .ZN(
        P1_U3252) );
  INV_X1 U12499 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9999) );
  MUX2_X1 U12500 ( .A(n9999), .B(P2_REG1_REG_10__SCAN_IN), .S(n10102), .Z(
        n10009) );
  INV_X1 U12501 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10000) );
  OR2_X1 U12502 ( .A1(n10011), .A2(n10000), .ZN(n10001) );
  NAND2_X1 U12503 ( .A1(n10002), .A2(n10001), .ZN(n14612) );
  INV_X1 U12504 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n14864) );
  MUX2_X1 U12505 ( .A(n14864), .B(P2_REG1_REG_6__SCAN_IN), .S(n14619), .Z(
        n14613) );
  NAND2_X1 U12506 ( .A1(n14612), .A2(n14613), .ZN(n14611) );
  OR2_X1 U12507 ( .A1(n14619), .A2(n14864), .ZN(n10003) );
  NAND2_X1 U12508 ( .A1(n14611), .A2(n10003), .ZN(n14625) );
  INV_X1 U12509 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n14866) );
  MUX2_X1 U12510 ( .A(n14866), .B(P2_REG1_REG_7__SCAN_IN), .S(n14632), .Z(
        n14626) );
  NAND2_X1 U12511 ( .A1(n14625), .A2(n14626), .ZN(n14624) );
  OR2_X1 U12512 ( .A1(n14632), .A2(n14866), .ZN(n10004) );
  NAND2_X1 U12513 ( .A1(n14624), .A2(n10004), .ZN(n14641) );
  INV_X1 U12514 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n14868) );
  MUX2_X1 U12515 ( .A(n14868), .B(P2_REG1_REG_8__SCAN_IN), .S(n14645), .Z(
        n14642) );
  NAND2_X1 U12516 ( .A1(n14641), .A2(n14642), .ZN(n14640) );
  OR2_X1 U12517 ( .A1(n14645), .A2(n14868), .ZN(n10005) );
  NAND2_X1 U12518 ( .A1(n14640), .A2(n10005), .ZN(n10081) );
  INV_X1 U12519 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n14870) );
  MUX2_X1 U12520 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n14870), .S(n10083), .Z(
        n10082) );
  OR2_X1 U12521 ( .A1(n10081), .A2(n10082), .ZN(n10079) );
  NAND2_X1 U12522 ( .A1(n10083), .A2(n14870), .ZN(n10006) );
  NAND2_X1 U12523 ( .A1(n10079), .A2(n10006), .ZN(n10008) );
  INV_X1 U12524 ( .A(n10097), .ZN(n10007) );
  AOI211_X1 U12525 ( .C1(n10009), .C2(n10008), .A(n10007), .B(n14716), .ZN(
        n10029) );
  XNOR2_X1 U12526 ( .A(n10102), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n10024) );
  INV_X1 U12527 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10010) );
  OR2_X1 U12528 ( .A1(n10011), .A2(n10010), .ZN(n10012) );
  NAND2_X1 U12529 ( .A1(n10013), .A2(n10012), .ZN(n14615) );
  XNOR2_X1 U12530 ( .A(n14619), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n14616) );
  NAND2_X1 U12531 ( .A1(n14615), .A2(n14616), .ZN(n14614) );
  INV_X1 U12532 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10014) );
  OR2_X1 U12533 ( .A1(n14619), .A2(n10014), .ZN(n10015) );
  NAND2_X1 U12534 ( .A1(n14614), .A2(n10015), .ZN(n14628) );
  XNOR2_X1 U12535 ( .A(n14632), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n14629) );
  NAND2_X1 U12536 ( .A1(n14628), .A2(n14629), .ZN(n14627) );
  INV_X1 U12537 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10016) );
  OR2_X1 U12538 ( .A1(n14632), .A2(n10016), .ZN(n10017) );
  NAND2_X1 U12539 ( .A1(n14627), .A2(n10017), .ZN(n14638) );
  XNOR2_X1 U12540 ( .A(n14645), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n14639) );
  NAND2_X1 U12541 ( .A1(n14638), .A2(n14639), .ZN(n14637) );
  INV_X1 U12542 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10018) );
  OR2_X1 U12543 ( .A1(n14645), .A2(n10018), .ZN(n10019) );
  NAND2_X1 U12544 ( .A1(n14637), .A2(n10019), .ZN(n10086) );
  INV_X1 U12545 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10020) );
  MUX2_X1 U12546 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n10020), .S(n10083), .Z(
        n10085) );
  OR2_X1 U12547 ( .A1(n10086), .A2(n10085), .ZN(n10088) );
  NAND2_X1 U12548 ( .A1(n10083), .A2(n10020), .ZN(n10021) );
  NAND2_X1 U12549 ( .A1(n10088), .A2(n10021), .ZN(n10023) );
  INV_X1 U12550 ( .A(n10104), .ZN(n10022) );
  INV_X1 U12551 ( .A(n14724), .ZN(n14706) );
  AOI211_X1 U12552 ( .C1(n10024), .C2(n10023), .A(n10022), .B(n14706), .ZN(
        n10028) );
  INV_X1 U12553 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14231) );
  NAND2_X1 U12554 ( .A1(n14728), .A2(n10102), .ZN(n10026) );
  NAND2_X1 U12555 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n10025)
         );
  OAI211_X1 U12556 ( .C1(n14231), .C2(n14731), .A(n10026), .B(n10025), .ZN(
        n10027) );
  OR3_X1 U12557 ( .A1(n10029), .A2(n10028), .A3(n10027), .ZN(P2_U3224) );
  INV_X1 U12558 ( .A(n12425), .ZN(n12437) );
  INV_X1 U12559 ( .A(n10030), .ZN(n10032) );
  OAI222_X1 U12560 ( .A1(n12437), .A2(P3_U3151), .B1(n14215), .B2(n10032), 
        .C1(n10031), .C2(n14213), .ZN(P3_U3278) );
  OAI211_X1 U12561 ( .C1(n14706), .C2(P2_REG2_REG_0__SCAN_IN), .A(
        P2_IR_REG_0__SCAN_IN), .B(n14659), .ZN(n10033) );
  AOI21_X1 U12562 ( .B1(n14657), .B2(n7729), .A(n10033), .ZN(n10037) );
  AOI21_X1 U12563 ( .B1(n14724), .B2(P2_REG2_REG_0__SCAN_IN), .A(
        P2_IR_REG_0__SCAN_IN), .ZN(n10036) );
  AOI22_X1 U12564 ( .A1(n14598), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n10035) );
  NAND3_X1 U12565 ( .A1(n10033), .A2(n14657), .A3(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10034) );
  OAI211_X1 U12566 ( .C1(n10037), .C2(n10036), .A(n10035), .B(n10034), .ZN(
        P2_U3214) );
  OR2_X1 U12567 ( .A1(n14516), .A2(n6486), .ZN(n10040) );
  INV_X2 U12568 ( .A(n10578), .ZN(n10594) );
  INV_X2 U12569 ( .A(n10594), .ZN(n13465) );
  AOI22_X1 U12570 ( .A1(n13465), .A2(n10396), .B1(n10042), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n10039) );
  NAND2_X1 U12571 ( .A1(n10040), .A2(n10039), .ZN(n10044) );
  INV_X1 U12572 ( .A(n10044), .ZN(n10224) );
  AOI22_X1 U12573 ( .A1(n6449), .A2(n10396), .B1(n10042), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n10043) );
  NAND2_X1 U12574 ( .A1(n10045), .A2(n10044), .ZN(n10226) );
  INV_X1 U12575 ( .A(n10226), .ZN(n10046) );
  AOI21_X1 U12576 ( .B1(n10224), .B2(n10047), .A(n10046), .ZN(n13611) );
  OR2_X1 U12577 ( .A1(n10061), .A2(P1_D_REG_0__SCAN_IN), .ZN(n10049) );
  NAND2_X1 U12578 ( .A1(n10049), .A2(n10048), .ZN(n10416) );
  INV_X1 U12579 ( .A(n10416), .ZN(n10060) );
  NOR4_X1 U12580 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n10058) );
  NOR4_X1 U12581 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n10057) );
  OR4_X1 U12582 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n10055) );
  NOR4_X1 U12583 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n10053) );
  NOR4_X1 U12584 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n10052) );
  NOR4_X1 U12585 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n10051) );
  NOR4_X1 U12586 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n10050) );
  NAND4_X1 U12587 ( .A1(n10053), .A2(n10052), .A3(n10051), .A4(n10050), .ZN(
        n10054) );
  NOR4_X1 U12588 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n10055), .A4(n10054), .ZN(n10056) );
  AND3_X1 U12589 ( .A1(n10058), .A2(n10057), .A3(n10056), .ZN(n10059) );
  OR2_X1 U12590 ( .A1(n10061), .A2(n10059), .ZN(n10415) );
  NAND2_X1 U12591 ( .A1(n10060), .A2(n10415), .ZN(n10538) );
  INV_X1 U12592 ( .A(n10538), .ZN(n10064) );
  OR2_X1 U12593 ( .A1(n10061), .A2(P1_D_REG_1__SCAN_IN), .ZN(n10063) );
  NAND2_X1 U12594 ( .A1(n10063), .A2(n10062), .ZN(n10418) );
  INV_X1 U12595 ( .A(n10418), .ZN(n11074) );
  NAND2_X1 U12596 ( .A1(n10064), .A2(n11074), .ZN(n10071) );
  OR2_X1 U12597 ( .A1(n10068), .A2(n10071), .ZN(n10069) );
  INV_X1 U12598 ( .A(n10069), .ZN(n10067) );
  OR2_X1 U12599 ( .A1(n10041), .A2(n10867), .ZN(n14528) );
  OR2_X1 U12600 ( .A1(n10041), .A2(n14536), .ZN(n10065) );
  AND2_X1 U12601 ( .A1(n14584), .A2(n14534), .ZN(n10066) );
  NAND2_X1 U12602 ( .A1(n10067), .A2(n10066), .ZN(n14330) );
  NAND2_X1 U12603 ( .A1(n14508), .A2(n13747), .ZN(n10540) );
  OR2_X1 U12604 ( .A1(n10069), .A2(n14528), .ZN(n10070) );
  NAND2_X1 U12605 ( .A1(n13952), .A2(n10070), .ZN(n14335) );
  NAND2_X1 U12606 ( .A1(n10540), .A2(n10071), .ZN(n10608) );
  NAND2_X1 U12607 ( .A1(n10608), .A2(n10541), .ZN(n13478) );
  AOI22_X1 U12608 ( .A1(n14335), .A2(n10396), .B1(n13478), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n10074) );
  INV_X1 U12609 ( .A(n10071), .ZN(n10072) );
  NAND2_X1 U12610 ( .A1(n10541), .A2(n10072), .ZN(n13544) );
  OR2_X1 U12611 ( .A1(n13544), .A2(n14533), .ZN(n14325) );
  INV_X1 U12612 ( .A(n14325), .ZN(n13567) );
  NAND2_X1 U12613 ( .A1(n13567), .A2(n8100), .ZN(n10073) );
  OAI211_X1 U12614 ( .C1(n13611), .C2(n14330), .A(n10074), .B(n10073), .ZN(
        P1_U3232) );
  INV_X1 U12615 ( .A(n10075), .ZN(n10077) );
  OAI222_X1 U12616 ( .A1(n14085), .A2(n10076), .B1(n14088), .B2(n10077), .C1(
        n14417), .C2(P1_U3086), .ZN(P1_U3342) );
  OAI222_X1 U12617 ( .A1(n13314), .A2(n10078), .B1(n6452), .B2(n10077), .C1(
        n14660), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U12618 ( .A(n10079), .ZN(n10080) );
  AOI21_X1 U12619 ( .B1(n10082), .B2(n10081), .A(n10080), .ZN(n10093) );
  INV_X1 U12620 ( .A(n10083), .ZN(n10091) );
  INV_X1 U12621 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10084) );
  NAND2_X1 U12622 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n11091) );
  OAI21_X1 U12623 ( .B1(n14731), .B2(n10084), .A(n11091), .ZN(n10090) );
  NAND2_X1 U12624 ( .A1(n10086), .A2(n10085), .ZN(n10087) );
  AOI21_X1 U12625 ( .B1(n10088), .B2(n10087), .A(n14706), .ZN(n10089) );
  AOI211_X1 U12626 ( .C1(n14728), .C2(n10091), .A(n10090), .B(n10089), .ZN(
        n10092) );
  OAI21_X1 U12627 ( .B1(n10093), .B2(n14716), .A(n10092), .ZN(P2_U3223) );
  INV_X1 U12628 ( .A(SI_18_), .ZN(n10095) );
  OAI222_X1 U12629 ( .A1(P3_U3151), .A2(n12452), .B1(n14213), .B2(n10095), 
        .C1(n14215), .C2(n10094), .ZN(P3_U3277) );
  INV_X1 U12630 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n15147) );
  XNOR2_X1 U12631 ( .A(n12928), .B(n15147), .ZN(n10101) );
  NAND2_X1 U12632 ( .A1(n10102), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10096) );
  NAND2_X1 U12633 ( .A1(n10097), .A2(n10096), .ZN(n12910) );
  INV_X1 U12634 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n14874) );
  MUX2_X1 U12635 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n14874), .S(n12903), .Z(
        n12909) );
  NAND2_X1 U12636 ( .A1(n12910), .A2(n12909), .ZN(n12908) );
  NAND2_X1 U12637 ( .A1(n12903), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10098) );
  NAND2_X1 U12638 ( .A1(n12908), .A2(n10098), .ZN(n10100) );
  INV_X1 U12639 ( .A(n12930), .ZN(n10099) );
  AOI21_X1 U12640 ( .B1(n10101), .B2(n10100), .A(n10099), .ZN(n10112) );
  XNOR2_X1 U12641 ( .A(n12928), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n10107) );
  NAND2_X1 U12642 ( .A1(n10102), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10103) );
  INV_X1 U12643 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11161) );
  XNOR2_X1 U12644 ( .A(n12903), .B(n11161), .ZN(n12906) );
  NAND2_X1 U12645 ( .A1(n12905), .A2(n12906), .ZN(n12904) );
  OR2_X1 U12646 ( .A1(n12903), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10105) );
  NAND2_X1 U12647 ( .A1(n12904), .A2(n10105), .ZN(n10106) );
  NAND2_X1 U12648 ( .A1(n10106), .A2(n10107), .ZN(n12916) );
  OAI21_X1 U12649 ( .B1(n10107), .B2(n10106), .A(n12916), .ZN(n10110) );
  AND2_X1 U12650 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n11439) );
  AOI21_X1 U12651 ( .B1(n14598), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n11439), 
        .ZN(n10108) );
  OAI21_X1 U12652 ( .B1(n12928), .B2(n14659), .A(n10108), .ZN(n10109) );
  AOI21_X1 U12653 ( .B1(n10110), .B2(n14724), .A(n10109), .ZN(n10111) );
  OAI21_X1 U12654 ( .B1(n10112), .B2(n14716), .A(n10111), .ZN(P2_U3226) );
  OAI222_X1 U12655 ( .A1(n14215), .A2(n10114), .B1(n14213), .B2(n10113), .C1(
        P3_U3151), .C2(n12459), .ZN(P3_U3276) );
  INV_X1 U12656 ( .A(n10169), .ZN(n10115) );
  NAND2_X1 U12657 ( .A1(n10115), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12304) );
  NAND2_X1 U12658 ( .A1(n10177), .A2(n12304), .ZN(n10128) );
  OR2_X1 U12659 ( .A1(n12273), .A2(n10115), .ZN(n10116) );
  AND2_X1 U12660 ( .A1(n8829), .A2(n10116), .ZN(n10127) );
  AND2_X1 U12661 ( .A1(n10128), .A2(n10127), .ZN(n10130) );
  INV_X1 U12662 ( .A(n10130), .ZN(n10117) );
  MUX2_X1 U12663 ( .A(n10117), .B(n12333), .S(n12299), .Z(n14917) );
  INV_X1 U12664 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10120) );
  INV_X1 U12665 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10119) );
  INV_X4 U12666 ( .A(n10118), .ZN(n12455) );
  MUX2_X1 U12667 ( .A(n10120), .B(n10119), .S(n12455), .Z(n10121) );
  MUX2_X1 U12668 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n9191), .Z(n10122) );
  NOR2_X1 U12669 ( .A1(n10122), .A2(n6614), .ZN(n10258) );
  AOI21_X1 U12670 ( .B1(n10122), .B2(n6614), .A(n10258), .ZN(n10123) );
  NAND2_X1 U12671 ( .A1(n10123), .A2(n10202), .ZN(n10354) );
  OAI21_X1 U12672 ( .B1(n10202), .B2(n10123), .A(n10354), .ZN(n10141) );
  NOR2_X2 U12673 ( .A1(n12333), .A2(n12299), .ZN(n14924) );
  INV_X1 U12674 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n14962) );
  NAND2_X1 U12675 ( .A1(n6625), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10124) );
  AOI21_X1 U12676 ( .B1(n14962), .B2(n10125), .A(n6503), .ZN(n10139) );
  NAND2_X1 U12677 ( .A1(n10130), .A2(n10126), .ZN(n14933) );
  INV_X1 U12678 ( .A(n10127), .ZN(n10129) );
  AOI22_X1 U12679 ( .A1(n14931), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10138) );
  NAND2_X1 U12680 ( .A1(n10130), .A2(n12455), .ZN(n14927) );
  INV_X1 U12681 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15026) );
  INV_X1 U12682 ( .A(n10143), .ZN(n10131) );
  NAND2_X1 U12683 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10204), .ZN(n10132) );
  NAND2_X1 U12684 ( .A1(n10131), .A2(n10132), .ZN(n10134) );
  NOR2_X1 U12685 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10132), .ZN(n10278) );
  INV_X1 U12686 ( .A(n10278), .ZN(n10133) );
  NAND2_X1 U12687 ( .A1(n10134), .A2(n10133), .ZN(n10135) );
  AOI21_X1 U12688 ( .B1(n15026), .B2(n10135), .A(n10277), .ZN(n10136) );
  OR2_X1 U12689 ( .A1(n14927), .A2(n10136), .ZN(n10137) );
  OAI211_X1 U12690 ( .C1(n10139), .C2(n14933), .A(n10138), .B(n10137), .ZN(
        n10140) );
  AOI21_X1 U12691 ( .B1(n10141), .B2(n14924), .A(n10140), .ZN(n10142) );
  OAI21_X1 U12692 ( .B1(n6614), .B2(n14917), .A(n10142), .ZN(P3_U3183) );
  NAND2_X1 U12693 ( .A1(n12752), .A2(n10144), .ZN(n10147) );
  OAI21_X1 U12694 ( .B1(n10145), .B2(n12459), .A(n10537), .ZN(n10146) );
  NAND3_X1 U12695 ( .A1(n12332), .A2(n11931), .A3(n14954), .ZN(n10149) );
  NAND2_X1 U12696 ( .A1(n14947), .A2(n11931), .ZN(n10150) );
  NAND2_X1 U12697 ( .A1(n10151), .A2(n10150), .ZN(n10152) );
  NAND2_X1 U12698 ( .A1(n10238), .A2(n10153), .ZN(n10245) );
  XNOR2_X1 U12699 ( .A(n14943), .B(n11931), .ZN(n10154) );
  XNOR2_X1 U12700 ( .A(n10154), .B(n12331), .ZN(n10246) );
  XNOR2_X1 U12701 ( .A(n14976), .B(n11931), .ZN(n10489) );
  XNOR2_X1 U12702 ( .A(n10489), .B(n10499), .ZN(n10159) );
  NAND2_X1 U12703 ( .A1(n10161), .A2(n10154), .ZN(n10160) );
  AND2_X1 U12704 ( .A1(n10159), .A2(n10160), .ZN(n10155) );
  NAND2_X1 U12705 ( .A1(n10166), .A2(n15001), .ZN(n10156) );
  OAI22_X1 U12706 ( .A1(n10167), .A2(n10156), .B1(n10168), .B2(n10178), .ZN(
        n10157) );
  NAND2_X1 U12707 ( .A1(n10157), .A2(n12298), .ZN(n14881) );
  NAND2_X1 U12708 ( .A1(n10491), .A2(n14257), .ZN(n10185) );
  AOI21_X1 U12709 ( .B1(n10158), .B2(n10160), .A(n10159), .ZN(n10184) );
  OAI22_X1 U12710 ( .A1(n10161), .A2(n12055), .B1(n10492), .B2(n12057), .ZN(
        n10483) );
  INV_X1 U12711 ( .A(n10178), .ZN(n10163) );
  NOR2_X1 U12712 ( .A1(n10177), .A2(n12290), .ZN(n10162) );
  NAND2_X1 U12713 ( .A1(n10167), .A2(n14955), .ZN(n10165) );
  NOR2_X1 U12714 ( .A1(n10177), .A2(n15001), .ZN(n10164) );
  AOI22_X1 U12715 ( .A1(n10483), .A2(n14884), .B1(n14976), .B2(n12062), .ZN(
        n10183) );
  NAND2_X1 U12716 ( .A1(n10167), .A2(n10166), .ZN(n10175) );
  INV_X1 U12717 ( .A(n10168), .ZN(n10173) );
  NAND3_X1 U12718 ( .A1(n10171), .A2(n10170), .A3(n10169), .ZN(n10172) );
  AOI21_X1 U12719 ( .B1(n10178), .B2(n10173), .A(n10172), .ZN(n10174) );
  NAND2_X1 U12720 ( .A1(n10175), .A2(n10174), .ZN(n10176) );
  NAND2_X1 U12721 ( .A1(n10176), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10181) );
  NOR2_X1 U12722 ( .A1(n10177), .A2(n10389), .ZN(n10179) );
  NAND2_X1 U12723 ( .A1(n10179), .A2(n10178), .ZN(n10180) );
  MUX2_X1 U12724 ( .A(n14893), .B(P3_STATE_REG_SCAN_IN), .S(
        P3_REG3_REG_3__SCAN_IN), .Z(n10182) );
  OAI211_X1 U12725 ( .C1(n10185), .C2(n10184), .A(n10183), .B(n10182), .ZN(
        P3_U3158) );
  MUX2_X1 U12726 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n13702), .S(n13710), .Z(
        n10189) );
  AOI21_X1 U12727 ( .B1(n10192), .B2(n10187), .A(n10186), .ZN(n10188) );
  AOI21_X1 U12728 ( .B1(n10189), .B2(n10188), .A(n13701), .ZN(n10201) );
  INV_X1 U12729 ( .A(n13710), .ZN(n10199) );
  INV_X1 U12730 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10190) );
  NAND2_X1 U12731 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n11696)
         );
  OAI21_X1 U12732 ( .B1(n14492), .B2(n10190), .A(n11696), .ZN(n10198) );
  MUX2_X1 U12733 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n13711), .S(n13710), .Z(
        n10195) );
  OAI21_X1 U12734 ( .B1(n10193), .B2(n10192), .A(n10191), .ZN(n10194) );
  NOR2_X1 U12735 ( .A1(n10194), .A2(n10195), .ZN(n13709) );
  AOI21_X1 U12736 ( .B1(n10195), .B2(n10194), .A(n13709), .ZN(n10196) );
  NOR2_X1 U12737 ( .A1(n10196), .A2(n14478), .ZN(n10197) );
  AOI211_X1 U12738 ( .C1(n14489), .C2(n10199), .A(n10198), .B(n10197), .ZN(
        n10200) );
  OAI21_X1 U12739 ( .B1(n10201), .B2(n14482), .A(n10200), .ZN(P1_U3255) );
  INV_X1 U12740 ( .A(n14933), .ZN(n12434) );
  INV_X1 U12741 ( .A(n14927), .ZN(n10336) );
  NOR3_X1 U12742 ( .A1(n12434), .A2(n10336), .A3(n14924), .ZN(n10208) );
  MUX2_X1 U12743 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n12455), .Z(n10203) );
  AOI21_X1 U12744 ( .B1(n10204), .B2(n10203), .A(n10202), .ZN(n10207) );
  AOI22_X1 U12745 ( .A1(n14931), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n10206) );
  INV_X1 U12746 ( .A(n14917), .ZN(n12419) );
  OAI211_X1 U12747 ( .C1(n10208), .C2(n10207), .A(n10206), .B(n10205), .ZN(
        P3_U3182) );
  OAI22_X1 U12748 ( .A1(n14529), .A2(n6486), .B1(n14564), .B2(n10594), .ZN(
        n10211) );
  OR2_X1 U12749 ( .A1(n8624), .A2(n13747), .ZN(n10210) );
  XNOR2_X1 U12750 ( .A(n10211), .B(n13404), .ZN(n10575) );
  OR2_X1 U12751 ( .A1(n14529), .A2(n13360), .ZN(n10213) );
  NAND2_X1 U12752 ( .A1(n13462), .A2(n11339), .ZN(n10212) );
  NAND2_X1 U12753 ( .A1(n10213), .A2(n10212), .ZN(n10573) );
  XNOR2_X1 U12754 ( .A(n10575), .B(n10573), .ZN(n10229) );
  NAND2_X1 U12755 ( .A1(n8100), .A2(n6449), .ZN(n10214) );
  NAND2_X1 U12756 ( .A1(n10215), .A2(n10214), .ZN(n10216) );
  XNOR2_X1 U12757 ( .A(n10216), .B(n13404), .ZN(n10219) );
  NAND2_X1 U12758 ( .A1(n13479), .A2(n13462), .ZN(n10218) );
  NAND2_X1 U12759 ( .A1(n8100), .A2(n10598), .ZN(n10217) );
  AND2_X1 U12760 ( .A1(n10218), .A2(n10217), .ZN(n10220) );
  NAND2_X1 U12761 ( .A1(n10219), .A2(n10220), .ZN(n10227) );
  INV_X1 U12762 ( .A(n10219), .ZN(n10222) );
  INV_X1 U12763 ( .A(n10220), .ZN(n10221) );
  NAND2_X1 U12764 ( .A1(n10222), .A2(n10221), .ZN(n10223) );
  NAND2_X1 U12765 ( .A1(n10224), .A2(n13463), .ZN(n10225) );
  NAND2_X1 U12766 ( .A1(n10226), .A2(n10225), .ZN(n13475) );
  NAND2_X1 U12767 ( .A1(n13474), .A2(n10227), .ZN(n10228) );
  OAI21_X1 U12768 ( .B1(n10229), .B2(n10228), .A(n10577), .ZN(n10230) );
  NAND2_X1 U12769 ( .A1(n10230), .A2(n13570), .ZN(n10235) );
  INV_X1 U12770 ( .A(n13544), .ZN(n13534) );
  OR2_X1 U12771 ( .A1(n10231), .A2(n14533), .ZN(n10233) );
  NAND2_X1 U12772 ( .A1(n8100), .A2(n13929), .ZN(n10232) );
  NAND2_X1 U12773 ( .A1(n10233), .A2(n10232), .ZN(n11331) );
  AOI22_X1 U12774 ( .A1(n13534), .A2(n11331), .B1(n13478), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10234) );
  OAI211_X1 U12775 ( .C1(n14564), .C2(n13580), .A(n10235), .B(n10234), .ZN(
        P1_U3237) );
  NOR2_X1 U12776 ( .A1(n12073), .A2(P3_U3151), .ZN(n10257) );
  INV_X1 U12777 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10244) );
  INV_X1 U12778 ( .A(n12141), .ZN(n14953) );
  NAND3_X1 U12779 ( .A1(n14953), .A2(n10236), .A3(n11980), .ZN(n10237) );
  OAI211_X1 U12780 ( .C1(n6502), .C2(n14947), .A(n10238), .B(n10237), .ZN(
        n10239) );
  NAND2_X1 U12781 ( .A1(n10239), .A2(n14257), .ZN(n10243) );
  NAND2_X1 U12782 ( .A1(n12334), .A2(n12300), .ZN(n10241) );
  INV_X1 U12783 ( .A(n12057), .ZN(n12069) );
  NAND2_X1 U12784 ( .A1(n12331), .A2(n12069), .ZN(n10240) );
  NAND2_X1 U12785 ( .A1(n10241), .A2(n10240), .ZN(n14950) );
  AOI22_X1 U12786 ( .A1(n14950), .A2(n14884), .B1(n12062), .B2(n14954), .ZN(
        n10242) );
  OAI211_X1 U12787 ( .C1(n10257), .C2(n10244), .A(n10243), .B(n10242), .ZN(
        P3_U3162) );
  INV_X1 U12788 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10251) );
  OAI21_X1 U12789 ( .B1(n10246), .B2(n10245), .A(n10158), .ZN(n10247) );
  NAND2_X1 U12790 ( .A1(n10247), .A2(n14257), .ZN(n10250) );
  OAI22_X1 U12791 ( .A1(n8816), .A2(n12055), .B1(n10499), .B2(n12057), .ZN(
        n14942) );
  AOI22_X1 U12792 ( .A1(n14942), .A2(n14884), .B1(n10248), .B2(n12062), .ZN(
        n10249) );
  OAI211_X1 U12793 ( .C1(n10257), .C2(n10251), .A(n10250), .B(n10249), .ZN(
        P3_U3177) );
  INV_X1 U12794 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10256) );
  NOR2_X1 U12795 ( .A1(n8816), .A2(n12057), .ZN(n10391) );
  AOI22_X1 U12796 ( .A1(n10391), .A2(n14884), .B1(n12062), .B2(n10252), .ZN(
        n10255) );
  INV_X1 U12797 ( .A(n12334), .ZN(n10253) );
  NOR2_X1 U12798 ( .A1(n10253), .A2(n10252), .ZN(n12138) );
  INV_X1 U12799 ( .A(n12138), .ZN(n12139) );
  NAND2_X1 U12800 ( .A1(n14953), .A2(n12139), .ZN(n12113) );
  NAND2_X1 U12801 ( .A1(n12113), .A2(n14257), .ZN(n10254) );
  OAI211_X1 U12802 ( .C1(n10257), .C2(n10256), .A(n10255), .B(n10254), .ZN(
        P3_U3172) );
  INV_X1 U12803 ( .A(n10258), .ZN(n10353) );
  INV_X1 U12804 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10260) );
  INV_X1 U12805 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10259) );
  MUX2_X1 U12806 ( .A(n10260), .B(n10259), .S(n12455), .Z(n10261) );
  NAND2_X1 U12807 ( .A1(n10261), .A2(n10359), .ZN(n10264) );
  INV_X1 U12808 ( .A(n10261), .ZN(n10262) );
  NAND2_X1 U12809 ( .A1(n10262), .A2(n6448), .ZN(n10263) );
  NAND2_X1 U12810 ( .A1(n10264), .A2(n10263), .ZN(n10352) );
  INV_X1 U12811 ( .A(n10264), .ZN(n10271) );
  INV_X1 U12812 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10485) );
  INV_X1 U12813 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10265) );
  MUX2_X1 U12814 ( .A(n10485), .B(n10265), .S(n12455), .Z(n10266) );
  NAND2_X1 U12815 ( .A1(n10266), .A2(n10317), .ZN(n10444) );
  INV_X1 U12816 ( .A(n10266), .ZN(n10268) );
  INV_X1 U12817 ( .A(n10317), .ZN(n10267) );
  NAND2_X1 U12818 ( .A1(n10268), .A2(n10267), .ZN(n10269) );
  AND2_X1 U12819 ( .A1(n10444), .A2(n10269), .ZN(n10270) );
  OAI21_X1 U12820 ( .B1(n10351), .B2(n10271), .A(n10270), .ZN(n10445) );
  INV_X1 U12821 ( .A(n10445), .ZN(n10273) );
  NOR3_X1 U12822 ( .A1(n10351), .A2(n10271), .A3(n10270), .ZN(n10272) );
  OAI21_X1 U12823 ( .B1(n10273), .B2(n10272), .A(n14924), .ZN(n10290) );
  NAND2_X1 U12824 ( .A1(P3_REG2_REG_2__SCAN_IN), .A2(n6448), .ZN(n10275) );
  OAI21_X1 U12825 ( .B1(P3_REG2_REG_2__SCAN_IN), .B2(n6448), .A(n10275), .ZN(
        n10342) );
  NOR2_X1 U12826 ( .A1(n10343), .A2(n10342), .ZN(n10341) );
  AOI21_X1 U12827 ( .B1(P3_REG2_REG_2__SCAN_IN), .B2(n6448), .A(n10341), .ZN(
        n10291) );
  AOI21_X1 U12828 ( .B1(n10485), .B2(n10276), .A(n10292), .ZN(n10287) );
  NAND2_X1 U12829 ( .A1(P3_REG1_REG_2__SCAN_IN), .A2(n6447), .ZN(n10280) );
  OAI21_X1 U12830 ( .B1(P3_REG1_REG_2__SCAN_IN), .B2(n6448), .A(n10280), .ZN(
        n10345) );
  XNOR2_X1 U12831 ( .A(n10316), .B(n10317), .ZN(n10282) );
  NOR2_X1 U12832 ( .A1(n10265), .A2(n10282), .ZN(n10318) );
  AOI21_X1 U12833 ( .B1(n10265), .B2(n10282), .A(n10318), .ZN(n10283) );
  OR2_X1 U12834 ( .A1(n14927), .A2(n10283), .ZN(n10286) );
  NOR2_X1 U12835 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10486), .ZN(n10284) );
  AOI21_X1 U12836 ( .B1(n14931), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10284), .ZN(
        n10285) );
  OAI211_X1 U12837 ( .C1(n10287), .C2(n14933), .A(n10286), .B(n10285), .ZN(
        n10288) );
  AOI21_X1 U12838 ( .B1(n12419), .B2(n10317), .A(n10288), .ZN(n10289) );
  NAND2_X1 U12839 ( .A1(n10290), .A2(n10289), .ZN(P3_U3185) );
  NOR2_X1 U12840 ( .A1(n10317), .A2(n10291), .ZN(n10293) );
  NAND2_X1 U12841 ( .A1(P3_REG2_REG_4__SCAN_IN), .A2(n10321), .ZN(n10294) );
  OAI21_X1 U12842 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n10321), .A(n10294), .ZN(
        n10433) );
  INV_X1 U12843 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10372) );
  INV_X1 U12844 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10309) );
  OR2_X1 U12845 ( .A1(n10325), .A2(n10309), .ZN(n10510) );
  NAND2_X1 U12846 ( .A1(n10325), .A2(n10309), .ZN(n10297) );
  NAND2_X1 U12847 ( .A1(n10510), .A2(n10297), .ZN(n10299) );
  INV_X1 U12848 ( .A(n10511), .ZN(n10298) );
  AOI21_X1 U12849 ( .B1(n10300), .B2(n10299), .A(n10298), .ZN(n10340) );
  INV_X1 U12850 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n15087) );
  INV_X1 U12851 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15030) );
  MUX2_X1 U12852 ( .A(n15087), .B(n15030), .S(n12455), .Z(n10301) );
  NAND2_X1 U12853 ( .A1(n10301), .A2(n10450), .ZN(n10304) );
  INV_X1 U12854 ( .A(n10301), .ZN(n10302) );
  NAND2_X1 U12855 ( .A1(n10302), .A2(n10321), .ZN(n10303) );
  NAND2_X1 U12856 ( .A1(n10304), .A2(n10303), .ZN(n10443) );
  INV_X1 U12857 ( .A(n10304), .ZN(n10375) );
  INV_X1 U12858 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10305) );
  MUX2_X1 U12859 ( .A(n10372), .B(n10305), .S(n12455), .Z(n10306) );
  NAND2_X1 U12860 ( .A1(n10306), .A2(n10385), .ZN(n10314) );
  INV_X1 U12861 ( .A(n10306), .ZN(n10307) );
  NAND2_X1 U12862 ( .A1(n10307), .A2(n6810), .ZN(n10308) );
  AND2_X1 U12863 ( .A1(n10314), .A2(n10308), .ZN(n10374) );
  INV_X1 U12864 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10324) );
  MUX2_X1 U12865 ( .A(n10309), .B(n10324), .S(n12455), .Z(n10310) );
  NAND2_X1 U12866 ( .A1(n10310), .A2(n10325), .ZN(n10517) );
  INV_X1 U12867 ( .A(n10310), .ZN(n10311) );
  NAND2_X1 U12868 ( .A1(n10311), .A2(n10334), .ZN(n10312) );
  NAND2_X1 U12869 ( .A1(n10517), .A2(n10312), .ZN(n10313) );
  AOI21_X1 U12870 ( .B1(n10373), .B2(n10314), .A(n10313), .ZN(n10523) );
  AND3_X1 U12871 ( .A1(n10373), .A2(n10314), .A3(n10313), .ZN(n10315) );
  OAI21_X1 U12872 ( .B1(n10523), .B2(n10315), .A(n14924), .ZN(n10339) );
  NOR2_X1 U12873 ( .A1(n10317), .A2(n10316), .ZN(n10319) );
  NAND2_X1 U12874 ( .A1(P3_REG1_REG_4__SCAN_IN), .A2(n10321), .ZN(n10320) );
  OAI21_X1 U12875 ( .B1(P3_REG1_REG_4__SCAN_IN), .B2(n10321), .A(n10320), .ZN(
        n10435) );
  NOR2_X1 U12876 ( .A1(n10436), .A2(n10435), .ZN(n10434) );
  NOR2_X1 U12877 ( .A1(n10385), .A2(n10322), .ZN(n10323) );
  XNOR2_X1 U12878 ( .A(n10322), .B(n10385), .ZN(n10381) );
  INV_X1 U12879 ( .A(n10328), .ZN(n10330) );
  OR2_X1 U12880 ( .A1(n10325), .A2(n10324), .ZN(n10514) );
  NAND2_X1 U12881 ( .A1(n10325), .A2(n10324), .ZN(n10326) );
  NAND2_X1 U12882 ( .A1(n10514), .A2(n10326), .ZN(n10327) );
  INV_X1 U12883 ( .A(n10327), .ZN(n10329) );
  OAI21_X1 U12884 ( .B1(n10330), .B2(n10329), .A(n10515), .ZN(n10337) );
  INV_X1 U12885 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10331) );
  NOR2_X1 U12886 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10331), .ZN(n10332) );
  AOI21_X1 U12887 ( .B1(n14931), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n10332), .ZN(
        n10333) );
  OAI21_X1 U12888 ( .B1(n14917), .B2(n10334), .A(n10333), .ZN(n10335) );
  AOI21_X1 U12889 ( .B1(n10337), .B2(n10336), .A(n10335), .ZN(n10338) );
  OAI211_X1 U12890 ( .C1(n10340), .C2(n14933), .A(n10339), .B(n10338), .ZN(
        P3_U3188) );
  AOI21_X1 U12891 ( .B1(n10343), .B2(n10342), .A(n10341), .ZN(n10350) );
  AOI22_X1 U12892 ( .A1(n14931), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10349) );
  AOI21_X1 U12893 ( .B1(n10346), .B2(n10345), .A(n10344), .ZN(n10347) );
  OR2_X1 U12894 ( .A1(n14927), .A2(n10347), .ZN(n10348) );
  OAI211_X1 U12895 ( .C1(n10350), .C2(n14933), .A(n10349), .B(n10348), .ZN(
        n10358) );
  INV_X1 U12896 ( .A(n10351), .ZN(n10356) );
  NAND3_X1 U12897 ( .A1(n10354), .A2(n10353), .A3(n10352), .ZN(n10355) );
  INV_X1 U12898 ( .A(n14924), .ZN(n14906) );
  AOI21_X1 U12899 ( .B1(n10356), .B2(n10355), .A(n14906), .ZN(n10357) );
  AOI211_X1 U12900 ( .C1(n12419), .C2(n10359), .A(n10358), .B(n10357), .ZN(
        n10360) );
  INV_X1 U12901 ( .A(n10360), .ZN(P3_U3184) );
  INV_X1 U12902 ( .A(n10361), .ZN(n10364) );
  OAI222_X1 U12903 ( .A1(n13314), .A2(n10363), .B1(n6452), .B2(n10364), .C1(
        n10362), .C2(P2_U3088), .ZN(P2_U3311) );
  OAI222_X1 U12904 ( .A1(n14085), .A2(n10365), .B1(n14088), .B2(n10364), .C1(
        n14459), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U12905 ( .A(n10366), .ZN(n10368) );
  INV_X1 U12906 ( .A(n13714), .ZN(n14425) );
  OAI222_X1 U12907 ( .A1(n14085), .A2(n10367), .B1(n14088), .B2(n10368), .C1(
        n14425), .C2(P1_U3086), .ZN(P1_U3341) );
  OAI222_X1 U12908 ( .A1(n13314), .A2(n10369), .B1(n6452), .B2(n10368), .C1(
        n12919), .C2(P2_U3088), .ZN(P2_U3313) );
  AOI21_X1 U12909 ( .B1(n10372), .B2(n10371), .A(n10370), .ZN(n10388) );
  INV_X1 U12910 ( .A(n10373), .ZN(n10377) );
  NOR3_X1 U12911 ( .A1(n10442), .A2(n10375), .A3(n10374), .ZN(n10376) );
  OAI21_X1 U12912 ( .B1(n10377), .B2(n10376), .A(n14924), .ZN(n10387) );
  INV_X1 U12913 ( .A(n14931), .ZN(n12368) );
  INV_X1 U12914 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n10379) );
  AND2_X1 U12915 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n12010) );
  INV_X1 U12916 ( .A(n12010), .ZN(n10378) );
  OAI21_X1 U12917 ( .B1(n12368), .B2(n10379), .A(n10378), .ZN(n10384) );
  AOI21_X1 U12918 ( .B1(n10305), .B2(n10381), .A(n10380), .ZN(n10382) );
  NOR2_X1 U12919 ( .A1(n10382), .A2(n14927), .ZN(n10383) );
  AOI211_X1 U12920 ( .C1(n12419), .C2(n10385), .A(n10384), .B(n10383), .ZN(
        n10386) );
  OAI211_X1 U12921 ( .C1(n10388), .C2(n14933), .A(n10387), .B(n10386), .ZN(
        P3_U3187) );
  INV_X1 U12922 ( .A(n10389), .ZN(n10390) );
  NOR2_X1 U12923 ( .A1(n10390), .A2(n15014), .ZN(n10392) );
  AOI21_X1 U12924 ( .B1(n12113), .B2(n10392), .A(n10391), .ZN(n10550) );
  INV_X1 U12925 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10393) );
  OAI22_X1 U12926 ( .A1(n12730), .A2(n10546), .B1(n15025), .B2(n10393), .ZN(
        n10394) );
  INV_X1 U12927 ( .A(n10394), .ZN(n10395) );
  OAI21_X1 U12928 ( .B1(n10550), .B2(n15023), .A(n10395), .ZN(P3_U3390) );
  NAND2_X1 U12929 ( .A1(n14518), .A2(n10396), .ZN(n14515) );
  NAND2_X1 U12930 ( .A1(n10397), .A2(n14515), .ZN(n10400) );
  NAND2_X1 U12931 ( .A1(n10398), .A2(n14556), .ZN(n10399) );
  NAND2_X1 U12932 ( .A1(n10400), .A2(n10399), .ZN(n11333) );
  NAND2_X1 U12933 ( .A1(n11333), .A2(n11334), .ZN(n10402) );
  NAND2_X1 U12934 ( .A1(n14529), .A2(n14564), .ZN(n10401) );
  NAND2_X1 U12935 ( .A1(n10402), .A2(n10401), .ZN(n10697) );
  XNOR2_X1 U12936 ( .A(n10696), .B(n10697), .ZN(n10413) );
  OAI21_X1 U12937 ( .B1(n6435), .B2(n10404), .A(n10403), .ZN(n11329) );
  NAND2_X1 U12938 ( .A1(n11329), .A2(n11330), .ZN(n10406) );
  NAND2_X1 U12939 ( .A1(n10406), .A2(n10405), .ZN(n10705) );
  XNOR2_X1 U12940 ( .A(n10696), .B(n10705), .ZN(n10411) );
  OR2_X1 U12941 ( .A1(n8624), .A2(n14536), .ZN(n10409) );
  NAND2_X1 U12942 ( .A1(n10407), .A2(n14537), .ZN(n10408) );
  NAND2_X1 U12943 ( .A1(n10409), .A2(n10408), .ZN(n14519) );
  AOI22_X1 U12944 ( .A1(n13929), .A2(n13599), .B1(n13597), .B2(n14507), .ZN(
        n10410) );
  OAI21_X1 U12945 ( .B1(n10411), .B2(n14548), .A(n10410), .ZN(n10412) );
  AOI21_X1 U12946 ( .B1(n14588), .B2(n10413), .A(n10412), .ZN(n11083) );
  INV_X1 U12947 ( .A(n11312), .ZN(n10414) );
  OAI211_X1 U12948 ( .C1(n11079), .C2(n11335), .A(n10414), .B(n14508), .ZN(
        n11076) );
  NAND2_X1 U12949 ( .A1(n11083), .A2(n11076), .ZN(n10544) );
  AND2_X1 U12950 ( .A1(n10416), .A2(n10415), .ZN(n10417) );
  AND2_X1 U12951 ( .A1(n10540), .A2(n10418), .ZN(n10419) );
  AND2_X2 U12952 ( .A1(n11075), .A2(n10419), .ZN(n14589) );
  NAND2_X1 U12953 ( .A1(n14589), .A2(n14574), .ZN(n14077) );
  OAI22_X1 U12954 ( .A1(n14077), .A2(n11079), .B1(n14589), .B2(n8121), .ZN(
        n10420) );
  AOI21_X1 U12955 ( .B1(n10544), .B2(n14589), .A(n10420), .ZN(n10421) );
  INV_X1 U12956 ( .A(n10421), .ZN(P1_U3468) );
  OR2_X1 U12957 ( .A1(n10422), .A2(P2_U3088), .ZN(n10474) );
  INV_X1 U12958 ( .A(n10474), .ZN(n10431) );
  INV_X1 U12959 ( .A(n12828), .ZN(n12798) );
  NAND2_X1 U12960 ( .A1(n13152), .A2(n12899), .ZN(n10423) );
  OAI21_X1 U12961 ( .B1(n10424), .B2(n13069), .A(n10423), .ZN(n10558) );
  OAI21_X1 U12962 ( .B1(n10427), .B2(n10426), .A(n10425), .ZN(n10428) );
  AOI22_X1 U12963 ( .A1(n12798), .A2(n10558), .B1(n12865), .B2(n10428), .ZN(
        n10430) );
  NAND2_X1 U12964 ( .A1(n12871), .A2(n10889), .ZN(n10429) );
  OAI211_X1 U12965 ( .C1(n10431), .C2(n10885), .A(n10430), .B(n10429), .ZN(
        P2_U3194) );
  AOI21_X1 U12966 ( .B1(n6607), .B2(n10433), .A(n10432), .ZN(n10441) );
  INV_X1 U12967 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10502) );
  NOR2_X1 U12968 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10502), .ZN(n10439) );
  AOI21_X1 U12969 ( .B1(n10436), .B2(n10435), .A(n10434), .ZN(n10437) );
  NOR2_X1 U12970 ( .A1(n10437), .A2(n14927), .ZN(n10438) );
  AOI211_X1 U12971 ( .C1(n14931), .C2(P3_ADDR_REG_4__SCAN_IN), .A(n10439), .B(
        n10438), .ZN(n10440) );
  OAI21_X1 U12972 ( .B1(n10441), .B2(n14933), .A(n10440), .ZN(n10449) );
  INV_X1 U12973 ( .A(n10442), .ZN(n10447) );
  NAND3_X1 U12974 ( .A1(n10445), .A2(n10444), .A3(n10443), .ZN(n10446) );
  AOI21_X1 U12975 ( .B1(n10447), .B2(n10446), .A(n14906), .ZN(n10448) );
  AOI211_X1 U12976 ( .C1(n12419), .C2(n10450), .A(n10449), .B(n10448), .ZN(
        n10451) );
  INV_X1 U12977 ( .A(n10451), .ZN(P3_U3186) );
  INV_X1 U12978 ( .A(n10452), .ZN(n10454) );
  OAI222_X1 U12979 ( .A1(n14085), .A2(n10453), .B1(n14088), .B2(n10454), .C1(
        P1_U3086), .C2(n14437), .ZN(P1_U3340) );
  OAI222_X1 U12980 ( .A1(n13314), .A2(n10455), .B1(n6452), .B2(n10454), .C1(
        P2_U3088), .C2(n14678), .ZN(P2_U3312) );
  INV_X1 U12981 ( .A(n10425), .ZN(n10457) );
  NOR2_X1 U12982 ( .A1(n10457), .A2(n10456), .ZN(n10461) );
  INV_X1 U12983 ( .A(n10659), .ZN(n10459) );
  NAND2_X1 U12984 ( .A1(n10459), .A2(n10458), .ZN(n10460) );
  NOR2_X1 U12985 ( .A1(n10461), .A2(n10460), .ZN(n10660) );
  AOI21_X1 U12986 ( .B1(n10461), .B2(n10460), .A(n10660), .ZN(n10465) );
  NAND2_X1 U12987 ( .A1(n13152), .A2(n12898), .ZN(n10462) );
  OAI21_X1 U12988 ( .B1(n11273), .B2(n13069), .A(n10462), .ZN(n10877) );
  AOI22_X1 U12989 ( .A1(n12798), .A2(n10877), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n10474), .ZN(n10464) );
  NAND2_X1 U12990 ( .A1(n12871), .A2(n10881), .ZN(n10463) );
  OAI211_X1 U12991 ( .C1(n10465), .C2(n12858), .A(n10464), .B(n10463), .ZN(
        P2_U3209) );
  INV_X1 U12992 ( .A(n10466), .ZN(n10470) );
  OAI222_X1 U12993 ( .A1(n14085), .A2(n10468), .B1(n14088), .B2(n10470), .C1(
        n10467), .C2(P1_U3086), .ZN(P1_U3338) );
  OAI222_X1 U12994 ( .A1(n13314), .A2(n10471), .B1(n6452), .B2(n10470), .C1(
        n10469), .C2(P2_U3088), .ZN(P2_U3310) );
  AOI22_X1 U12995 ( .A1(n12841), .A2(n10472), .B1(n14773), .B2(n12871), .ZN(
        n10477) );
  INV_X1 U12996 ( .A(n10473), .ZN(n10475) );
  AOI22_X1 U12997 ( .A1(n12865), .A2(n10475), .B1(n10474), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n10476) );
  OAI211_X1 U12998 ( .C1(n10478), .C2(n12869), .A(n10477), .B(n10476), .ZN(
        P2_U3204) );
  XNOR2_X1 U12999 ( .A(n10479), .B(n7278), .ZN(n14979) );
  AOI21_X1 U13000 ( .B1(n10480), .B2(n10481), .A(n14939), .ZN(n10484) );
  AOI21_X1 U13001 ( .B1(n10484), .B2(n10482), .A(n10483), .ZN(n14978) );
  MUX2_X1 U13002 ( .A(n10485), .B(n14978), .S(n14963), .Z(n10488) );
  AOI22_X1 U13003 ( .A1(n12618), .A2(n14976), .B1(n14959), .B2(n10486), .ZN(
        n10487) );
  OAI211_X1 U13004 ( .C1(n12621), .C2(n14979), .A(n10488), .B(n10487), .ZN(
        P3_U3230) );
  NAND2_X1 U13005 ( .A1(n8845), .A2(n10489), .ZN(n10490) );
  XNOR2_X1 U13006 ( .A(n12156), .B(n11931), .ZN(n10493) );
  NAND2_X1 U13007 ( .A1(n10492), .A2(n10493), .ZN(n10895) );
  INV_X1 U13008 ( .A(n10493), .ZN(n10494) );
  NAND2_X1 U13009 ( .A1(n10494), .A2(n12330), .ZN(n10495) );
  NAND2_X1 U13010 ( .A1(n10895), .A2(n10495), .ZN(n10497) );
  INV_X1 U13011 ( .A(n10896), .ZN(n10496) );
  AOI21_X1 U13012 ( .B1(n10498), .B2(n10497), .A(n10496), .ZN(n10507) );
  OR2_X1 U13013 ( .A1(n10499), .A2(n12055), .ZN(n10500) );
  OAI21_X1 U13014 ( .B1(n10902), .B2(n12057), .A(n10500), .ZN(n10803) );
  NAND2_X1 U13015 ( .A1(n12062), .A2(n14984), .ZN(n10501) );
  OAI21_X1 U13016 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n10502), .A(n10501), .ZN(
        n10505) );
  INV_X1 U13017 ( .A(n10503), .ZN(n10800) );
  NOR2_X1 U13018 ( .A1(n14893), .A2(n10800), .ZN(n10504) );
  AOI211_X1 U13019 ( .C1(n14884), .C2(n10803), .A(n10505), .B(n10504), .ZN(
        n10506) );
  OAI21_X1 U13020 ( .B1(n10507), .B2(n14881), .A(n10506), .ZN(P3_U3170) );
  OAI22_X1 U13021 ( .A1(n12655), .A2(n10546), .B1(n15034), .B2(n10119), .ZN(
        n10508) );
  INV_X1 U13022 ( .A(n10508), .ZN(n10509) );
  OAI21_X1 U13023 ( .B1(n10550), .B2(n15039), .A(n10509), .ZN(P3_U3459) );
  INV_X1 U13024 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10513) );
  AOI21_X1 U13025 ( .B1(n10513), .B2(n10512), .A(n10631), .ZN(n10533) );
  INV_X1 U13026 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15035) );
  AOI21_X1 U13027 ( .B1(n15035), .B2(n10516), .A(n10647), .ZN(n10530) );
  INV_X1 U13028 ( .A(n10517), .ZN(n10522) );
  MUX2_X1 U13029 ( .A(n10513), .B(n15035), .S(n12455), .Z(n10518) );
  NAND2_X1 U13030 ( .A1(n10518), .A2(n10645), .ZN(n10640) );
  INV_X1 U13031 ( .A(n10518), .ZN(n10519) );
  NAND2_X1 U13032 ( .A1(n10519), .A2(n6623), .ZN(n10520) );
  AND2_X1 U13033 ( .A1(n10640), .A2(n10520), .ZN(n10521) );
  OAI21_X1 U13034 ( .B1(n10523), .B2(n10522), .A(n10521), .ZN(n10641) );
  INV_X1 U13035 ( .A(n10641), .ZN(n10525) );
  NOR3_X1 U13036 ( .A1(n10523), .A2(n10522), .A3(n10521), .ZN(n10524) );
  OAI21_X1 U13037 ( .B1(n10525), .B2(n10524), .A(n14924), .ZN(n10529) );
  INV_X1 U13038 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n10936) );
  NOR2_X1 U13039 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10936), .ZN(n10527) );
  NOR2_X1 U13040 ( .A1(n14917), .A2(n6623), .ZN(n10526) );
  AOI211_X1 U13041 ( .C1(n14931), .C2(P3_ADDR_REG_7__SCAN_IN), .A(n10527), .B(
        n10526), .ZN(n10528) );
  OAI211_X1 U13042 ( .C1(n10530), .C2(n14927), .A(n10529), .B(n10528), .ZN(
        n10531) );
  INV_X1 U13043 ( .A(n10531), .ZN(n10532) );
  OAI21_X1 U13044 ( .B1(n10533), .B2(n14933), .A(n10532), .ZN(P3_U3189) );
  INV_X1 U13045 ( .A(n10534), .ZN(n10536) );
  OAI222_X1 U13046 ( .A1(P3_U3151), .A2(n10537), .B1(n14215), .B2(n10536), 
        .C1(n10535), .C2(n14213), .ZN(P3_U3275) );
  NOR2_X1 U13047 ( .A1(n10538), .A2(n11074), .ZN(n10539) );
  AND2_X1 U13048 ( .A1(n10540), .A2(n10539), .ZN(n10542) );
  AND2_X2 U13049 ( .A1(n10542), .A2(n10541), .ZN(n14597) );
  NAND2_X1 U13050 ( .A1(n14597), .A2(n14574), .ZN(n14032) );
  OAI22_X1 U13051 ( .A1(n14032), .A2(n11079), .B1(n14597), .B2(n9931), .ZN(
        n10543) );
  AOI21_X1 U13052 ( .B1(n10544), .B2(n14597), .A(n10543), .ZN(n10545) );
  INV_X1 U13053 ( .A(n10545), .ZN(P1_U3531) );
  NOR2_X1 U13054 ( .A1(n12489), .A2(n10546), .ZN(n10548) );
  NOR2_X1 U13055 ( .A1(n14963), .A2(n10120), .ZN(n10547) );
  AOI211_X1 U13056 ( .C1(n14959), .C2(P3_REG3_REG_0__SCAN_IN), .A(n10548), .B(
        n10547), .ZN(n10549) );
  OAI21_X1 U13057 ( .B1(n14965), .B2(n10550), .A(n10549), .ZN(P3_U3233) );
  INV_X1 U13058 ( .A(n14763), .ZN(n10551) );
  INV_X1 U13059 ( .A(n14839), .ZN(n14836) );
  INV_X1 U13060 ( .A(n14838), .ZN(n10556) );
  INV_X1 U13061 ( .A(n10553), .ZN(n10554) );
  XNOR2_X1 U13062 ( .A(n9529), .B(n10554), .ZN(n10891) );
  INV_X1 U13063 ( .A(n10891), .ZN(n10555) );
  OAI21_X1 U13064 ( .B1(n14836), .B2(n10556), .A(n10555), .ZN(n10565) );
  XNOR2_X1 U13065 ( .A(n10557), .B(n9529), .ZN(n10559) );
  AOI21_X1 U13066 ( .B1(n10559), .B2(n13169), .A(n10558), .ZN(n10886) );
  INV_X1 U13067 ( .A(n10872), .ZN(n10560) );
  OAI211_X1 U13068 ( .C1(n10562), .C2(n10561), .A(n9578), .B(n10560), .ZN(
        n10884) );
  NAND2_X1 U13069 ( .A1(n14841), .A2(n10889), .ZN(n10563) );
  AND2_X1 U13070 ( .A1(n10884), .A2(n10563), .ZN(n10564) );
  AND3_X1 U13071 ( .A1(n10565), .A2(n10886), .A3(n10564), .ZN(n14775) );
  NAND2_X1 U13072 ( .A1(n14873), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10566) );
  OAI21_X1 U13073 ( .B1(n14873), .B2(n14775), .A(n10566), .ZN(P2_U3500) );
  XNOR2_X1 U13074 ( .A(n10567), .B(n10568), .ZN(n10572) );
  OAI22_X1 U13075 ( .A1(n13067), .A2(n10691), .B1(n11085), .B2(n13069), .ZN(
        n11240) );
  NAND2_X1 U13076 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n14634) );
  INV_X1 U13077 ( .A(n14634), .ZN(n10569) );
  AOI21_X1 U13078 ( .B1(n12798), .B2(n11240), .A(n10569), .ZN(n10571) );
  INV_X1 U13079 ( .A(n12856), .ZN(n12867) );
  AOI22_X1 U13080 ( .A1(n11247), .A2(n12871), .B1(n12867), .B2(n11248), .ZN(
        n10570) );
  OAI211_X1 U13081 ( .C1(n10572), .C2(n12858), .A(n10571), .B(n10570), .ZN(
        P2_U3185) );
  INV_X1 U13082 ( .A(n10573), .ZN(n10574) );
  NAND2_X1 U13083 ( .A1(n10575), .A2(n10574), .ZN(n10576) );
  OAI22_X1 U13084 ( .A1(n10231), .A2(n6486), .B1(n11079), .B2(n10594), .ZN(
        n10579) );
  XNOR2_X1 U13085 ( .A(n10579), .B(n13463), .ZN(n10584) );
  OR2_X1 U13086 ( .A1(n10231), .A2(n13360), .ZN(n10581) );
  NAND2_X1 U13087 ( .A1(n6449), .A2(n13446), .ZN(n10580) );
  NAND2_X1 U13088 ( .A1(n10581), .A2(n10580), .ZN(n10583) );
  XNOR2_X1 U13089 ( .A(n10584), .B(n10583), .ZN(n13443) );
  NAND2_X1 U13090 ( .A1(n10584), .A2(n10583), .ZN(n10618) );
  OAI22_X1 U13091 ( .A1(n10709), .A2(n6486), .B1(n14569), .B2(n10594), .ZN(
        n10585) );
  XNOR2_X1 U13092 ( .A(n10585), .B(n13463), .ZN(n10620) );
  OR2_X1 U13093 ( .A1(n10709), .A2(n13360), .ZN(n10587) );
  NAND2_X1 U13094 ( .A1(n11318), .A2(n13462), .ZN(n10586) );
  NAND2_X1 U13095 ( .A1(n10587), .A2(n10586), .ZN(n10619) );
  NAND2_X1 U13096 ( .A1(n10620), .A2(n10619), .ZN(n10588) );
  AND2_X1 U13097 ( .A1(n10618), .A2(n10588), .ZN(n10589) );
  NAND2_X1 U13098 ( .A1(n10617), .A2(n10589), .ZN(n10593) );
  INV_X1 U13099 ( .A(n10620), .ZN(n10591) );
  INV_X1 U13100 ( .A(n10619), .ZN(n10590) );
  NAND2_X1 U13101 ( .A1(n10591), .A2(n10590), .ZN(n10592) );
  NAND2_X1 U13102 ( .A1(n13596), .A2(n6449), .ZN(n10596) );
  NAND2_X1 U13103 ( .A1(n11170), .A2(n13465), .ZN(n10595) );
  NAND2_X1 U13104 ( .A1(n10596), .A2(n10595), .ZN(n10597) );
  XNOR2_X1 U13105 ( .A(n10597), .B(n13404), .ZN(n10601) );
  NAND2_X1 U13106 ( .A1(n13596), .A2(n10598), .ZN(n10600) );
  NAND2_X1 U13107 ( .A1(n11170), .A2(n6449), .ZN(n10599) );
  AND2_X1 U13108 ( .A1(n10600), .A2(n10599), .ZN(n10602) );
  AND2_X1 U13109 ( .A1(n10601), .A2(n10602), .ZN(n10852) );
  INV_X1 U13110 ( .A(n10852), .ZN(n10605) );
  INV_X1 U13111 ( .A(n10601), .ZN(n10604) );
  INV_X1 U13112 ( .A(n10602), .ZN(n10603) );
  NAND2_X1 U13113 ( .A1(n10604), .A2(n10603), .ZN(n10851) );
  NAND2_X1 U13114 ( .A1(n10605), .A2(n10851), .ZN(n10606) );
  XNOR2_X1 U13115 ( .A(n10853), .B(n10606), .ZN(n10616) );
  NAND2_X1 U13116 ( .A1(n10608), .A2(n10607), .ZN(n10609) );
  NAND2_X1 U13117 ( .A1(n10609), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10610) );
  INV_X1 U13118 ( .A(n11170), .ZN(n10751) );
  NOR2_X1 U13119 ( .A1(n13580), .A2(n10751), .ZN(n10614) );
  INV_X1 U13120 ( .A(n13595), .ZN(n11006) );
  INV_X1 U13121 ( .A(n13929), .ZN(n14523) );
  OR2_X1 U13122 ( .A1(n13544), .A2(n14523), .ZN(n14326) );
  OR2_X1 U13123 ( .A1(n14326), .A2(n10709), .ZN(n10612) );
  OAI211_X1 U13124 ( .C1(n11006), .C2(n14325), .A(n10612), .B(n10611), .ZN(
        n10613) );
  AOI211_X1 U13125 ( .C1(n11169), .C2(n13562), .A(n10614), .B(n10613), .ZN(
        n10615) );
  OAI21_X1 U13126 ( .B1(n10616), .B2(n14330), .A(n10615), .ZN(P1_U3227) );
  NAND2_X1 U13127 ( .A1(n10617), .A2(n10618), .ZN(n10622) );
  XNOR2_X1 U13128 ( .A(n10620), .B(n10619), .ZN(n10621) );
  XNOR2_X1 U13129 ( .A(n10622), .B(n10621), .ZN(n10628) );
  OR2_X1 U13130 ( .A1(n10231), .A2(n14523), .ZN(n10624) );
  NAND2_X1 U13131 ( .A1(n13596), .A2(n14507), .ZN(n10623) );
  NAND2_X1 U13132 ( .A1(n10624), .A2(n10623), .ZN(n11307) );
  AND2_X1 U13133 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n13641) );
  AOI21_X1 U13134 ( .B1(n13534), .B2(n11307), .A(n13641), .ZN(n10626) );
  NAND2_X1 U13135 ( .A1(n14335), .A2(n11318), .ZN(n10625) );
  OAI211_X1 U13136 ( .C1(n14339), .C2(n11315), .A(n10626), .B(n10625), .ZN(
        n10627) );
  AOI21_X1 U13137 ( .B1(n10628), .B2(n13570), .A(n10627), .ZN(n10629) );
  INV_X1 U13138 ( .A(n10629), .ZN(P1_U3230) );
  NOR2_X1 U13139 ( .A1(n10645), .A2(n10630), .ZN(n10632) );
  NAND2_X1 U13140 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n10762), .ZN(n10633) );
  OAI21_X1 U13141 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n10762), .A(n10633), .ZN(
        n10634) );
  AOI21_X1 U13142 ( .B1(n6609), .B2(n10634), .A(n10759), .ZN(n10658) );
  INV_X1 U13143 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11065) );
  MUX2_X1 U13144 ( .A(n11065), .B(n15037), .S(n12455), .Z(n10636) );
  INV_X1 U13145 ( .A(n10762), .ZN(n10635) );
  NAND2_X1 U13146 ( .A1(n10636), .A2(n10635), .ZN(n10766) );
  INV_X1 U13147 ( .A(n10636), .ZN(n10637) );
  NAND2_X1 U13148 ( .A1(n10637), .A2(n10762), .ZN(n10638) );
  NAND2_X1 U13149 ( .A1(n10766), .A2(n10638), .ZN(n10639) );
  INV_X1 U13150 ( .A(n10772), .ZN(n10643) );
  NAND3_X1 U13151 ( .A1(n10641), .A2(n10640), .A3(n10639), .ZN(n10642) );
  AOI21_X1 U13152 ( .B1(n10643), .B2(n10642), .A(n14906), .ZN(n10656) );
  NOR2_X1 U13153 ( .A1(n10645), .A2(n10644), .ZN(n10646) );
  NAND2_X1 U13154 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n10762), .ZN(n10648) );
  OAI21_X1 U13155 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n10762), .A(n10648), .ZN(
        n10649) );
  AOI21_X1 U13156 ( .B1(n6602), .B2(n10649), .A(n10764), .ZN(n10650) );
  NOR2_X1 U13157 ( .A1(n10650), .A2(n14927), .ZN(n10655) );
  NOR2_X1 U13158 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10651), .ZN(n10652) );
  AOI21_X1 U13159 ( .B1(n14931), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n10652), .ZN(
        n10653) );
  OAI21_X1 U13160 ( .B1(n14917), .B2(n10762), .A(n10653), .ZN(n10654) );
  NOR3_X1 U13161 ( .A1(n10656), .A2(n10655), .A3(n10654), .ZN(n10657) );
  OAI21_X1 U13162 ( .B1(n10658), .B2(n14933), .A(n10657), .ZN(P3_U3190) );
  NOR2_X1 U13163 ( .A1(n10660), .A2(n10659), .ZN(n10661) );
  XNOR2_X1 U13164 ( .A(n10662), .B(n10661), .ZN(n10666) );
  INV_X1 U13165 ( .A(n12847), .ZN(n12875) );
  OAI22_X1 U13166 ( .A1(n12856), .A2(P2_REG3_REG_3__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n7744), .ZN(n10664) );
  OAI22_X1 U13167 ( .A1(n12829), .A2(n10825), .B1(n12869), .B2(n10690), .ZN(
        n10663) );
  AOI211_X1 U13168 ( .C1(n12875), .C2(n12897), .A(n10664), .B(n10663), .ZN(
        n10665) );
  OAI21_X1 U13169 ( .B1(n10666), .B2(n12858), .A(n10665), .ZN(P2_U3190) );
  INV_X1 U13170 ( .A(n10667), .ZN(n10668) );
  AOI21_X1 U13171 ( .B1(n10670), .B2(n10669), .A(n10668), .ZN(n10676) );
  OAI21_X1 U13172 ( .B1(n12856), .B2(n10672), .A(n10671), .ZN(n10674) );
  OAI22_X1 U13173 ( .A1(n12829), .A2(n11280), .B1(n12869), .B2(n11274), .ZN(
        n10673) );
  AOI211_X1 U13174 ( .C1(n12875), .C2(n12896), .A(n10674), .B(n10673), .ZN(
        n10675) );
  OAI21_X1 U13175 ( .B1(n10676), .B2(n12858), .A(n10675), .ZN(P2_U3202) );
  XNOR2_X1 U13176 ( .A(n10678), .B(n10677), .ZN(n10684) );
  INV_X1 U13177 ( .A(n11047), .ZN(n10679) );
  NAND2_X1 U13178 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n14621) );
  OAI21_X1 U13179 ( .B1(n12856), .B2(n10679), .A(n14621), .ZN(n10682) );
  INV_X1 U13180 ( .A(n11048), .ZN(n14808) );
  OAI22_X1 U13181 ( .A1(n12829), .A2(n14808), .B1(n12869), .B2(n10680), .ZN(
        n10681) );
  AOI211_X1 U13182 ( .C1(n12875), .C2(n12894), .A(n10682), .B(n10681), .ZN(
        n10683) );
  OAI21_X1 U13183 ( .B1(n10684), .B2(n12858), .A(n10683), .ZN(P2_U3211) );
  OAI21_X1 U13184 ( .B1(n10687), .B2(n10686), .A(n10685), .ZN(n10694) );
  NAND2_X1 U13185 ( .A1(n12867), .A2(n11031), .ZN(n10688) );
  OAI211_X1 U13186 ( .C1(n12847), .C2(n10690), .A(n10689), .B(n10688), .ZN(
        n10693) );
  OAI22_X1 U13187 ( .A1(n12829), .A2(n14801), .B1(n12869), .B2(n10691), .ZN(
        n10692) );
  AOI211_X1 U13188 ( .C1(n12865), .C2(n10694), .A(n10693), .B(n10692), .ZN(
        n10695) );
  INV_X1 U13189 ( .A(n10695), .ZN(P2_U3199) );
  NAND2_X1 U13190 ( .A1(n10697), .A2(n10696), .ZN(n10699) );
  NAND2_X1 U13191 ( .A1(n10231), .A2(n11079), .ZN(n10698) );
  NAND2_X1 U13192 ( .A1(n10699), .A2(n10698), .ZN(n11310) );
  INV_X1 U13193 ( .A(n10708), .ZN(n11311) );
  NAND2_X1 U13194 ( .A1(n11310), .A2(n11311), .ZN(n10701) );
  NAND2_X1 U13195 ( .A1(n10709), .A2(n14569), .ZN(n10700) );
  NAND2_X1 U13196 ( .A1(n10701), .A2(n10700), .ZN(n10738) );
  INV_X1 U13197 ( .A(n10712), .ZN(n10739) );
  NAND2_X1 U13198 ( .A1(n10738), .A2(n10739), .ZN(n10703) );
  INV_X1 U13199 ( .A(n13596), .ZN(n10862) );
  NAND2_X1 U13200 ( .A1(n10862), .A2(n10751), .ZN(n10702) );
  NAND2_X1 U13201 ( .A1(n10703), .A2(n10702), .ZN(n10830) );
  XNOR2_X1 U13202 ( .A(n10830), .B(n10833), .ZN(n10718) );
  NAND2_X1 U13203 ( .A1(n10705), .A2(n10704), .ZN(n10707) );
  NAND2_X1 U13204 ( .A1(n10707), .A2(n10706), .ZN(n11306) );
  NAND2_X1 U13205 ( .A1(n11306), .A2(n10708), .ZN(n10711) );
  NAND2_X1 U13206 ( .A1(n10709), .A2(n11318), .ZN(n10710) );
  NAND2_X1 U13207 ( .A1(n10711), .A2(n10710), .ZN(n10737) );
  NAND2_X1 U13208 ( .A1(n10737), .A2(n10712), .ZN(n10714) );
  NAND2_X1 U13209 ( .A1(n10862), .A2(n11170), .ZN(n10713) );
  NAND2_X1 U13210 ( .A1(n10714), .A2(n10713), .ZN(n10834) );
  XNOR2_X1 U13211 ( .A(n10834), .B(n10833), .ZN(n10716) );
  OAI22_X1 U13212 ( .A1(n10862), .A2(n14523), .B1(n11184), .B2(n14533), .ZN(
        n10715) );
  AOI21_X1 U13213 ( .B1(n10716), .B2(n14519), .A(n10715), .ZN(n10717) );
  OAI21_X1 U13214 ( .B1(n10718), .B2(n14549), .A(n10717), .ZN(n11099) );
  NAND2_X1 U13215 ( .A1(n11314), .A2(n10751), .ZN(n10744) );
  OR2_X1 U13216 ( .A1(n10744), .A2(n10857), .ZN(n10841) );
  INV_X1 U13217 ( .A(n10841), .ZN(n10719) );
  AOI211_X1 U13218 ( .C1(n10857), .C2(n10744), .A(n14526), .B(n10719), .ZN(
        n11104) );
  NOR2_X1 U13219 ( .A1(n11099), .A2(n11104), .ZN(n10725) );
  INV_X1 U13220 ( .A(n10857), .ZN(n11102) );
  INV_X1 U13221 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10720) );
  OAI22_X1 U13222 ( .A1(n14077), .A2(n11102), .B1(n14589), .B2(n10720), .ZN(
        n10721) );
  INV_X1 U13223 ( .A(n10721), .ZN(n10722) );
  OAI21_X1 U13224 ( .B1(n10725), .B2(n6712), .A(n10722), .ZN(P1_U3477) );
  OAI22_X1 U13225 ( .A1(n14032), .A2(n11102), .B1(n14597), .B2(n9935), .ZN(
        n10723) );
  INV_X1 U13226 ( .A(n10723), .ZN(n10724) );
  OAI21_X1 U13227 ( .B1(n10725), .B2(n14595), .A(n10724), .ZN(P1_U3534) );
  XNOR2_X1 U13228 ( .A(n7196), .B(n10728), .ZN(n10729) );
  XNOR2_X1 U13229 ( .A(n10726), .B(n10729), .ZN(n10736) );
  NAND2_X1 U13230 ( .A1(n13153), .A2(n12890), .ZN(n10731) );
  NAND2_X1 U13231 ( .A1(n13152), .A2(n12892), .ZN(n10730) );
  AND2_X1 U13232 ( .A1(n10731), .A2(n10730), .ZN(n11221) );
  OAI22_X1 U13233 ( .A1(n12828), .A2(n11221), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10732), .ZN(n10734) );
  INV_X1 U13234 ( .A(n11227), .ZN(n14822) );
  NOR2_X1 U13235 ( .A1(n12829), .A2(n14822), .ZN(n10733) );
  AOI211_X1 U13236 ( .C1(n12867), .C2(n11231), .A(n10734), .B(n10733), .ZN(
        n10735) );
  OAI21_X1 U13237 ( .B1(n10736), .B2(n12858), .A(n10735), .ZN(P2_U3193) );
  XNOR2_X1 U13238 ( .A(n10737), .B(n10739), .ZN(n10743) );
  XNOR2_X1 U13239 ( .A(n10738), .B(n10739), .ZN(n10740) );
  NAND2_X1 U13240 ( .A1(n10740), .A2(n14588), .ZN(n10742) );
  AOI22_X1 U13241 ( .A1(n13597), .A2(n13929), .B1(n14507), .B2(n13595), .ZN(
        n10741) );
  OAI211_X1 U13242 ( .C1(n10743), .C2(n14548), .A(n10742), .B(n10741), .ZN(
        n11167) );
  INV_X1 U13243 ( .A(n11167), .ZN(n10745) );
  OAI211_X1 U13244 ( .C1(n11314), .C2(n10751), .A(n14508), .B(n10744), .ZN(
        n11173) );
  NAND2_X1 U13245 ( .A1(n10745), .A2(n11173), .ZN(n10753) );
  OAI22_X1 U13246 ( .A1(n14077), .A2(n10751), .B1(n14589), .B2(n8158), .ZN(
        n10746) );
  AOI21_X1 U13247 ( .B1(n10753), .B2(n14589), .A(n10746), .ZN(n10747) );
  INV_X1 U13248 ( .A(n10747), .ZN(P1_U3474) );
  INV_X1 U13249 ( .A(n10748), .ZN(n10750) );
  OAI222_X1 U13250 ( .A1(P3_U3151), .A2(n12140), .B1(n14215), .B2(n10750), 
        .C1(n10749), .C2(n14213), .ZN(P3_U3274) );
  OAI22_X1 U13251 ( .A1(n14032), .A2(n10751), .B1(n14597), .B2(n9934), .ZN(
        n10752) );
  AOI21_X1 U13252 ( .B1(n10753), .B2(n14597), .A(n10752), .ZN(n10754) );
  INV_X1 U13253 ( .A(n10754), .ZN(P1_U3533) );
  INV_X1 U13254 ( .A(n10755), .ZN(n10757) );
  OAI222_X1 U13255 ( .A1(n14085), .A2(n10756), .B1(n14088), .B2(n10757), .C1(
        n14477), .C2(P1_U3086), .ZN(P1_U3337) );
  OAI222_X1 U13256 ( .A1(n13314), .A2(n10758), .B1(n6452), .B2(n10757), .C1(
        n12935), .C2(P2_U3088), .ZN(P2_U3309) );
  INV_X1 U13257 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10761) );
  INV_X1 U13258 ( .A(n10957), .ZN(n14207) );
  AOI21_X1 U13259 ( .B1(n10761), .B2(n10760), .A(n10951), .ZN(n10782) );
  INV_X1 U13260 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15040) );
  AOI21_X1 U13261 ( .B1(n15040), .B2(n10765), .A(n10958), .ZN(n10779) );
  INV_X1 U13262 ( .A(n10766), .ZN(n10771) );
  MUX2_X1 U13263 ( .A(n10761), .B(n15040), .S(n12455), .Z(n10767) );
  NAND2_X1 U13264 ( .A1(n10767), .A2(n10957), .ZN(n10970) );
  INV_X1 U13265 ( .A(n10767), .ZN(n10768) );
  NAND2_X1 U13266 ( .A1(n10768), .A2(n14207), .ZN(n10769) );
  AND2_X1 U13267 ( .A1(n10970), .A2(n10769), .ZN(n10770) );
  OAI21_X1 U13268 ( .B1(n10772), .B2(n10771), .A(n10770), .ZN(n10971) );
  INV_X1 U13269 ( .A(n10971), .ZN(n10774) );
  NOR3_X1 U13270 ( .A1(n10772), .A2(n10771), .A3(n10770), .ZN(n10773) );
  OAI21_X1 U13271 ( .B1(n10774), .B2(n10773), .A(n14924), .ZN(n10778) );
  NOR2_X1 U13272 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10926), .ZN(n10776) );
  NOR2_X1 U13273 ( .A1(n14917), .A2(n14207), .ZN(n10775) );
  AOI211_X1 U13274 ( .C1(n14931), .C2(P3_ADDR_REG_9__SCAN_IN), .A(n10776), .B(
        n10775), .ZN(n10777) );
  OAI211_X1 U13275 ( .C1(n10779), .C2(n14927), .A(n10778), .B(n10777), .ZN(
        n10780) );
  INV_X1 U13276 ( .A(n10780), .ZN(n10781) );
  OAI21_X1 U13277 ( .B1(n10782), .B2(n14933), .A(n10781), .ZN(P3_U3191) );
  INV_X1 U13278 ( .A(n10783), .ZN(n10785) );
  OAI22_X1 U13279 ( .A1(n12302), .A2(P3_U3151), .B1(SI_22_), .B2(n14213), .ZN(
        n10784) );
  AOI21_X1 U13280 ( .B1(n10785), .B2(n14223), .A(n10784), .ZN(P3_U3273) );
  NAND2_X1 U13281 ( .A1(n12333), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n10786) );
  OAI21_X1 U13282 ( .B1(n10787), .B2(n12333), .A(n10786), .ZN(P3_U3520) );
  XOR2_X1 U13283 ( .A(n12160), .B(n10788), .Z(n14991) );
  OAI21_X1 U13284 ( .B1(n10790), .B2(n8874), .A(n10789), .ZN(n10793) );
  OR2_X1 U13285 ( .A1(n10933), .A2(n12057), .ZN(n10792) );
  NAND2_X1 U13286 ( .A1(n12330), .A2(n12300), .ZN(n10791) );
  NAND2_X1 U13287 ( .A1(n10792), .A2(n10791), .ZN(n12013) );
  AOI21_X1 U13288 ( .B1(n10793), .B2(n14948), .A(n12013), .ZN(n10794) );
  OAI21_X1 U13289 ( .B1(n14991), .B2(n14936), .A(n10794), .ZN(n14993) );
  NAND2_X1 U13290 ( .A1(n14993), .A2(n14963), .ZN(n10798) );
  INV_X1 U13291 ( .A(n12012), .ZN(n10795) );
  OAI22_X1 U13292 ( .A1(n12489), .A2(n14990), .B1(n10795), .B2(n11656), .ZN(
        n10796) );
  AOI21_X1 U13293 ( .B1(n14965), .B2(P3_REG2_REG_5__SCAN_IN), .A(n10796), .ZN(
        n10797) );
  OAI211_X1 U13294 ( .C1(n14991), .C2(n14944), .A(n10798), .B(n10797), .ZN(
        P3_U3228) );
  XNOR2_X1 U13295 ( .A(n10799), .B(n12115), .ZN(n14986) );
  INV_X1 U13296 ( .A(n14986), .ZN(n14988) );
  INV_X1 U13297 ( .A(n12621), .ZN(n12492) );
  OAI22_X1 U13298 ( .A1(n12489), .A2(n12156), .B1(n10800), .B2(n11656), .ZN(
        n10807) );
  OAI211_X1 U13299 ( .C1(n10802), .C2(n12115), .A(n10801), .B(n14948), .ZN(
        n10805) );
  INV_X1 U13300 ( .A(n10803), .ZN(n10804) );
  NAND2_X1 U13301 ( .A1(n10805), .A2(n10804), .ZN(n14983) );
  MUX2_X1 U13302 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n14983), .S(n14963), .Z(
        n10806) );
  AOI211_X1 U13303 ( .C1(n14988), .C2(n12492), .A(n10807), .B(n10806), .ZN(
        n10808) );
  INV_X1 U13304 ( .A(n10808), .ZN(P3_U3229) );
  INV_X1 U13305 ( .A(n10809), .ZN(n10811) );
  INV_X1 U13306 ( .A(n14766), .ZN(n10810) );
  NAND3_X1 U13307 ( .A1(n10811), .A2(n10810), .A3(n14763), .ZN(n10816) );
  NAND2_X1 U13308 ( .A1(n13135), .A2(n10812), .ZN(n13163) );
  NAND2_X1 U13309 ( .A1(n13135), .A2(n14836), .ZN(n10813) );
  XNOR2_X1 U13310 ( .A(n10815), .B(n10814), .ZN(n14788) );
  XNOR2_X1 U13311 ( .A(n10870), .B(n10825), .ZN(n10817) );
  NOR2_X1 U13312 ( .A1(n10817), .A2(n13190), .ZN(n14784) );
  OAI22_X1 U13313 ( .A1(n13135), .A2(n10818), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13133), .ZN(n10827) );
  INV_X2 U13314 ( .A(n13135), .ZN(n13187) );
  NAND3_X1 U13315 ( .A1(n10874), .A2(n10821), .A3(n10820), .ZN(n10822) );
  NAND2_X1 U13316 ( .A1(n10819), .A2(n10822), .ZN(n10823) );
  AOI222_X1 U13317 ( .A1(n13169), .A2(n10823), .B1(n12895), .B2(n13153), .C1(
        n12897), .C2(n13152), .ZN(n14787) );
  OAI22_X1 U13318 ( .A1(n13187), .A2(n14787), .B1(n13178), .B2(n10825), .ZN(
        n10826) );
  AOI211_X1 U13319 ( .C1(n13185), .C2(n14784), .A(n10827), .B(n10826), .ZN(
        n10828) );
  OAI21_X1 U13320 ( .B1(n13182), .B2(n14788), .A(n10828), .ZN(P2_U3262) );
  INV_X1 U13321 ( .A(n10833), .ZN(n10829) );
  NAND2_X1 U13322 ( .A1(n10830), .A2(n10829), .ZN(n10832) );
  OR2_X1 U13323 ( .A1(n13595), .A2(n10857), .ZN(n10831) );
  NAND2_X1 U13324 ( .A1(n10832), .A2(n10831), .ZN(n11175) );
  INV_X1 U13325 ( .A(n11174), .ZN(n11182) );
  XNOR2_X1 U13326 ( .A(n11175), .B(n11182), .ZN(n10840) );
  NAND2_X1 U13327 ( .A1(n10834), .A2(n10833), .ZN(n10836) );
  NAND2_X1 U13328 ( .A1(n10857), .A2(n11006), .ZN(n10835) );
  XNOR2_X1 U13329 ( .A(n11183), .B(n11182), .ZN(n10838) );
  OAI22_X1 U13330 ( .A1(n11006), .A2(n14523), .B1(n11407), .B2(n14533), .ZN(
        n10837) );
  AOI21_X1 U13331 ( .B1(n10838), .B2(n14519), .A(n10837), .ZN(n10839) );
  OAI21_X1 U13332 ( .B1(n10840), .B2(n14549), .A(n10839), .ZN(n11107) );
  AOI211_X1 U13333 ( .C1(n11185), .C2(n10841), .A(n14526), .B(n11360), .ZN(
        n11112) );
  NOR2_X1 U13334 ( .A1(n11107), .A2(n11112), .ZN(n10846) );
  INV_X1 U13335 ( .A(n11185), .ZN(n11108) );
  OAI22_X1 U13336 ( .A1(n14032), .A2(n11108), .B1(n14597), .B2(n9936), .ZN(
        n10842) );
  INV_X1 U13337 ( .A(n10842), .ZN(n10843) );
  OAI21_X1 U13338 ( .B1(n10846), .B2(n14595), .A(n10843), .ZN(P1_U3535) );
  OAI22_X1 U13339 ( .A1(n14077), .A2(n11108), .B1(n14589), .B2(n8191), .ZN(
        n10844) );
  INV_X1 U13340 ( .A(n10844), .ZN(n10845) );
  OAI21_X1 U13341 ( .B1(n10846), .B2(n6712), .A(n10845), .ZN(P1_U3480) );
  INV_X1 U13342 ( .A(n10847), .ZN(n10849) );
  OAI222_X1 U13343 ( .A1(n14085), .A2(n10848), .B1(n14088), .B2(n10849), .C1(
        P1_U3086), .C2(n14536), .ZN(P1_U3336) );
  OAI222_X1 U13344 ( .A1(n13314), .A2(n10850), .B1(n6452), .B2(n10849), .C1(
        n11725), .C2(P2_U3088), .ZN(P2_U3308) );
  NAND2_X1 U13345 ( .A1(n10857), .A2(n13465), .ZN(n10855) );
  NAND2_X1 U13346 ( .A1(n13595), .A2(n13462), .ZN(n10854) );
  NAND2_X1 U13347 ( .A1(n10855), .A2(n10854), .ZN(n10856) );
  XNOR2_X1 U13348 ( .A(n10856), .B(n13463), .ZN(n10994) );
  AOI22_X1 U13349 ( .A1(n10857), .A2(n13462), .B1(n10598), .B2(n13595), .ZN(
        n10995) );
  XNOR2_X1 U13350 ( .A(n10994), .B(n10995), .ZN(n10858) );
  NAND2_X1 U13351 ( .A1(n10859), .A2(n10858), .ZN(n10998) );
  OAI211_X1 U13352 ( .C1(n10859), .C2(n10858), .A(n10998), .B(n13570), .ZN(
        n10865) );
  INV_X1 U13353 ( .A(n10860), .ZN(n11100) );
  AOI22_X1 U13354 ( .A1(n13567), .A2(n13594), .B1(P1_REG3_REG_6__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10861) );
  OAI21_X1 U13355 ( .B1(n10862), .B2(n14326), .A(n10861), .ZN(n10863) );
  AOI21_X1 U13356 ( .B1(n11100), .B2(n13562), .A(n10863), .ZN(n10864) );
  OAI211_X1 U13357 ( .C1(n11102), .C2(n13580), .A(n10865), .B(n10864), .ZN(
        P1_U3239) );
  INV_X1 U13358 ( .A(n10866), .ZN(n10892) );
  OAI222_X1 U13359 ( .A1(n14085), .A2(n10868), .B1(n14088), .B2(n10892), .C1(
        n10867), .C2(P1_U3086), .ZN(P1_U3335) );
  XNOR2_X1 U13360 ( .A(n10869), .B(n10876), .ZN(n14776) );
  INV_X1 U13361 ( .A(n10870), .ZN(n10871) );
  OAI211_X1 U13362 ( .C1(n14779), .C2(n10872), .A(n10871), .B(n13136), .ZN(
        n14777) );
  OAI22_X1 U13363 ( .A1(n13140), .A2(n14777), .B1(n13135), .B2(n10873), .ZN(
        n10880) );
  OAI21_X1 U13364 ( .B1(n10876), .B2(n10875), .A(n10874), .ZN(n10878) );
  AOI21_X1 U13365 ( .B1(n10878), .B2(n13169), .A(n10877), .ZN(n14778) );
  OAI22_X1 U13366 ( .A1(n13187), .A2(n14778), .B1(n7738), .B2(n13133), .ZN(
        n10879) );
  AOI211_X1 U13367 ( .C1(n13143), .C2(n10881), .A(n10880), .B(n10879), .ZN(
        n10882) );
  OAI21_X1 U13368 ( .B1(n13182), .B2(n14776), .A(n10882), .ZN(P2_U3263) );
  INV_X1 U13369 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10883) );
  OAI22_X1 U13370 ( .A1(n13140), .A2(n10884), .B1(n13135), .B2(n10883), .ZN(
        n10888) );
  OAI22_X1 U13371 ( .A1(n13187), .A2(n10886), .B1(n10885), .B2(n13133), .ZN(
        n10887) );
  AOI211_X1 U13372 ( .C1(n13143), .C2(n10889), .A(n10888), .B(n10887), .ZN(
        n10890) );
  OAI21_X1 U13373 ( .B1(n13182), .B2(n10891), .A(n10890), .ZN(P2_U3264) );
  OAI222_X1 U13374 ( .A1(n13314), .A2(n10894), .B1(P2_U3088), .B2(n10893), 
        .C1(n6452), .C2(n10892), .ZN(P2_U3307) );
  XNOR2_X1 U13375 ( .A(n10905), .B(n11980), .ZN(n10914) );
  XNOR2_X1 U13376 ( .A(n10933), .B(n10914), .ZN(n10900) );
  XNOR2_X1 U13377 ( .A(n12011), .B(n11931), .ZN(n10897) );
  XNOR2_X1 U13378 ( .A(n10897), .B(n10902), .ZN(n12008) );
  INV_X1 U13379 ( .A(n10897), .ZN(n10898) );
  NAND2_X1 U13380 ( .A1(n10898), .A2(n10902), .ZN(n10911) );
  NAND2_X1 U13381 ( .A1(n12006), .A2(n10911), .ZN(n10899) );
  NOR2_X1 U13382 ( .A1(n10899), .A2(n10900), .ZN(n10931) );
  AOI211_X1 U13383 ( .C1(n10900), .C2(n10899), .A(n14881), .B(n10931), .ZN(
        n10909) );
  INV_X1 U13384 ( .A(n10901), .ZN(n11131) );
  OR2_X1 U13385 ( .A1(n10902), .A2(n12055), .ZN(n10904) );
  OR2_X1 U13386 ( .A1(n11117), .A2(n12057), .ZN(n10903) );
  NAND2_X1 U13387 ( .A1(n10904), .A2(n10903), .ZN(n11134) );
  NAND2_X1 U13388 ( .A1(n11134), .A2(n14884), .ZN(n10907) );
  AOI22_X1 U13389 ( .A1(n12062), .A2(n10905), .B1(P3_REG3_REG_6__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10906) );
  OAI211_X1 U13390 ( .C1(n11131), .C2(n14893), .A(n10907), .B(n10906), .ZN(
        n10908) );
  OR2_X1 U13391 ( .A1(n10909), .A2(n10908), .ZN(P3_U3179) );
  XNOR2_X1 U13392 ( .A(n15015), .B(n11931), .ZN(n11386) );
  XNOR2_X1 U13393 ( .A(n11386), .B(n12325), .ZN(n10922) );
  XNOR2_X1 U13394 ( .A(n11014), .B(n11931), .ZN(n11115) );
  XNOR2_X1 U13395 ( .A(n15009), .B(n11931), .ZN(n10915) );
  XNOR2_X1 U13396 ( .A(n10935), .B(n10915), .ZN(n11118) );
  NAND2_X1 U13397 ( .A1(n10933), .A2(n10914), .ZN(n10910) );
  AND4_X1 U13398 ( .A1(n11115), .A2(n11118), .A3(n10911), .A4(n10910), .ZN(
        n10912) );
  INV_X1 U13399 ( .A(n11118), .ZN(n10913) );
  INV_X1 U13400 ( .A(n11115), .ZN(n10932) );
  OAI21_X1 U13401 ( .B1(n11117), .B2(n10913), .A(n10932), .ZN(n10917) );
  NOR2_X1 U13402 ( .A1(n10933), .A2(n10914), .ZN(n10930) );
  AOI22_X1 U13403 ( .A1(n10917), .A2(n10916), .B1(n10915), .B2(n12326), .ZN(
        n10918) );
  INV_X1 U13404 ( .A(n10922), .ZN(n10919) );
  INV_X1 U13405 ( .A(n14880), .ZN(n10920) );
  AOI21_X1 U13406 ( .B1(n10922), .B2(n10921), .A(n10920), .ZN(n10929) );
  OR2_X1 U13407 ( .A1(n10935), .A2(n12055), .ZN(n10923) );
  OAI21_X1 U13408 ( .B1(n11385), .B2(n12057), .A(n10923), .ZN(n11377) );
  NAND2_X1 U13409 ( .A1(n11377), .A2(n14884), .ZN(n10925) );
  NAND2_X1 U13410 ( .A1(n12062), .A2(n15015), .ZN(n10924) );
  OAI211_X1 U13411 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n10926), .A(n10925), .B(
        n10924), .ZN(n10927) );
  AOI21_X1 U13412 ( .B1(n11379), .B2(n12073), .A(n10927), .ZN(n10928) );
  OAI21_X1 U13413 ( .B1(n10929), .B2(n14881), .A(n10928), .ZN(P3_U3171) );
  NOR2_X1 U13414 ( .A1(n10931), .A2(n10930), .ZN(n11116) );
  XNOR2_X1 U13415 ( .A(n11116), .B(n10932), .ZN(n10940) );
  OR2_X1 U13416 ( .A1(n10933), .A2(n12055), .ZN(n10934) );
  OAI21_X1 U13417 ( .B1(n10935), .B2(n12057), .A(n10934), .ZN(n11015) );
  INV_X1 U13418 ( .A(n12062), .ZN(n14889) );
  OAI22_X1 U13419 ( .A1(n14889), .A2(n15002), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10936), .ZN(n10937) );
  AOI21_X1 U13420 ( .B1(n11015), .B2(n14884), .A(n10937), .ZN(n10939) );
  NAND2_X1 U13421 ( .A1(n12073), .A2(n11018), .ZN(n10938) );
  OAI211_X1 U13422 ( .C1(n10940), .C2(n14881), .A(n10939), .B(n10938), .ZN(
        P3_U3153) );
  NAND2_X1 U13423 ( .A1(n10941), .A2(n14223), .ZN(n10942) );
  OAI211_X1 U13424 ( .C1(n10943), .C2(n14213), .A(n10942), .B(n12304), .ZN(
        P3_U3272) );
  INV_X1 U13425 ( .A(n10944), .ZN(n10948) );
  OAI222_X1 U13426 ( .A1(n14085), .A2(n10946), .B1(n14088), .B2(n10948), .C1(
        P1_U3086), .C2(n10945), .ZN(P1_U3334) );
  OAI222_X1 U13427 ( .A1(n13314), .A2(n10949), .B1(n6452), .B2(n10948), .C1(
        n10947), .C2(P2_U3088), .ZN(P2_U3306) );
  NAND2_X1 U13428 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n12348), .ZN(n10952) );
  OAI21_X1 U13429 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n12348), .A(n10952), 
        .ZN(n10953) );
  AOI21_X1 U13430 ( .B1(n6601), .B2(n10953), .A(n12335), .ZN(n10954) );
  NAND2_X1 U13431 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n14886)
         );
  OAI21_X1 U13432 ( .B1(n10954), .B2(n14933), .A(n14886), .ZN(n10977) );
  NOR2_X1 U13433 ( .A1(n10957), .A2(n10956), .ZN(n10959) );
  NAND2_X1 U13434 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n12348), .ZN(n10960) );
  OAI21_X1 U13435 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(n12348), .A(n10960), 
        .ZN(n10961) );
  AOI21_X1 U13436 ( .B1(n10962), .B2(n10961), .A(n12350), .ZN(n10975) );
  AOI22_X1 U13437 ( .A1(n12419), .A2(n10965), .B1(n14931), .B2(
        P3_ADDR_REG_10__SCAN_IN), .ZN(n10974) );
  INV_X1 U13438 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10964) );
  INV_X1 U13439 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n10963) );
  MUX2_X1 U13440 ( .A(n10964), .B(n10963), .S(n12455), .Z(n10966) );
  NAND2_X1 U13441 ( .A1(n10966), .A2(n10965), .ZN(n12340) );
  INV_X1 U13442 ( .A(n10966), .ZN(n10967) );
  NAND2_X1 U13443 ( .A1(n10967), .A2(n12348), .ZN(n10968) );
  NAND2_X1 U13444 ( .A1(n12340), .A2(n10968), .ZN(n10969) );
  AOI21_X1 U13445 ( .B1(n10971), .B2(n10970), .A(n10969), .ZN(n12342) );
  AND3_X1 U13446 ( .A1(n10971), .A2(n10970), .A3(n10969), .ZN(n10972) );
  OAI21_X1 U13447 ( .B1(n12342), .B2(n10972), .A(n14924), .ZN(n10973) );
  OAI211_X1 U13448 ( .C1(n10975), .C2(n14927), .A(n10974), .B(n10973), .ZN(
        n10976) );
  OR2_X1 U13449 ( .A1(n10977), .A2(n10976), .ZN(P3_U3192) );
  OR2_X1 U13450 ( .A1(n10979), .A2(n10978), .ZN(n10980) );
  NAND2_X1 U13451 ( .A1(n10981), .A2(n10980), .ZN(n14840) );
  OAI211_X1 U13452 ( .C1(n10983), .C2(n7072), .A(n10982), .B(n13169), .ZN(
        n10986) );
  NAND2_X1 U13453 ( .A1(n13153), .A2(n12888), .ZN(n10985) );
  NAND2_X1 U13454 ( .A1(n13152), .A2(n12890), .ZN(n10984) );
  AND2_X1 U13455 ( .A1(n10985), .A2(n10984), .ZN(n11142) );
  NAND2_X1 U13456 ( .A1(n10986), .A2(n11142), .ZN(n14846) );
  NAND2_X1 U13457 ( .A1(n14846), .A2(n13135), .ZN(n10993) );
  INV_X1 U13458 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10988) );
  INV_X1 U13459 ( .A(n11144), .ZN(n10987) );
  OAI22_X1 U13460 ( .A1(n13135), .A2(n10988), .B1(n10987), .B2(n13133), .ZN(
        n10991) );
  AOI21_X1 U13461 ( .B1(n11209), .B2(n14842), .A(n13190), .ZN(n10989) );
  NAND2_X1 U13462 ( .A1(n10989), .A2(n11157), .ZN(n14844) );
  NOR2_X1 U13463 ( .A1(n14844), .A2(n13140), .ZN(n10990) );
  AOI211_X1 U13464 ( .C1(n13143), .C2(n14842), .A(n10991), .B(n10990), .ZN(
        n10992) );
  OAI211_X1 U13465 ( .C1(n13182), .C2(n14840), .A(n10993), .B(n10992), .ZN(
        P2_U3255) );
  INV_X1 U13466 ( .A(n10994), .ZN(n10996) );
  OR2_X1 U13467 ( .A1(n10996), .A2(n10995), .ZN(n10997) );
  NAND2_X1 U13468 ( .A1(n10998), .A2(n10997), .ZN(n11004) );
  NAND2_X1 U13469 ( .A1(n11185), .A2(n13465), .ZN(n11000) );
  NAND2_X1 U13470 ( .A1(n13594), .A2(n13462), .ZN(n10999) );
  NAND2_X1 U13471 ( .A1(n11000), .A2(n10999), .ZN(n11001) );
  XNOR2_X1 U13472 ( .A(n11001), .B(n13463), .ZN(n11289) );
  AND2_X1 U13473 ( .A1(n13594), .A2(n10598), .ZN(n11002) );
  AOI21_X1 U13474 ( .B1(n11185), .B2(n6449), .A(n11002), .ZN(n11287) );
  XNOR2_X1 U13475 ( .A(n11289), .B(n11287), .ZN(n11003) );
  NAND2_X1 U13476 ( .A1(n11004), .A2(n11003), .ZN(n11291) );
  OAI211_X1 U13477 ( .C1(n11004), .C2(n11003), .A(n11291), .B(n13570), .ZN(
        n11010) );
  INV_X1 U13478 ( .A(n11109), .ZN(n11008) );
  AOI22_X1 U13479 ( .A1(n13567), .A2(n13593), .B1(P1_REG3_REG_7__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11005) );
  OAI21_X1 U13480 ( .B1(n11006), .B2(n14326), .A(n11005), .ZN(n11007) );
  AOI21_X1 U13481 ( .B1(n11008), .B2(n13562), .A(n11007), .ZN(n11009) );
  OAI211_X1 U13482 ( .C1(n11108), .C2(n13580), .A(n11010), .B(n11009), .ZN(
        P1_U3213) );
  XNOR2_X1 U13483 ( .A(n11011), .B(n11014), .ZN(n15003) );
  OAI211_X1 U13484 ( .C1(n11014), .C2(n11013), .A(n11012), .B(n14948), .ZN(
        n11017) );
  INV_X1 U13485 ( .A(n11015), .ZN(n11016) );
  OAI211_X1 U13486 ( .C1(n14936), .C2(n15003), .A(n11017), .B(n11016), .ZN(
        n15005) );
  NAND2_X1 U13487 ( .A1(n15005), .A2(n14963), .ZN(n11022) );
  INV_X1 U13488 ( .A(n11018), .ZN(n11019) );
  OAI22_X1 U13489 ( .A1(n12489), .A2(n15002), .B1(n11019), .B2(n11656), .ZN(
        n11020) );
  AOI21_X1 U13490 ( .B1(n14965), .B2(P3_REG2_REG_7__SCAN_IN), .A(n11020), .ZN(
        n11021) );
  OAI211_X1 U13491 ( .C1(n15003), .C2(n14944), .A(n11022), .B(n11021), .ZN(
        P3_U3226) );
  XNOR2_X1 U13492 ( .A(n11023), .B(n7067), .ZN(n14799) );
  NAND3_X1 U13493 ( .A1(n11271), .A2(n11025), .A3(n11024), .ZN(n11026) );
  NAND2_X1 U13494 ( .A1(n11027), .A2(n11026), .ZN(n11028) );
  NAND2_X1 U13495 ( .A1(n11028), .A2(n13169), .ZN(n11030) );
  AOI22_X1 U13496 ( .A1(n13153), .A2(n12893), .B1(n13152), .B2(n12895), .ZN(
        n11029) );
  NAND2_X1 U13497 ( .A1(n11030), .A2(n11029), .ZN(n14803) );
  OAI211_X1 U13498 ( .C1(n11276), .C2(n14801), .A(n9578), .B(n11045), .ZN(
        n14800) );
  INV_X1 U13499 ( .A(n13133), .ZN(n13175) );
  AOI22_X1 U13500 ( .A1(n13187), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n11031), 
        .B2(n13175), .ZN(n11034) );
  NAND2_X1 U13501 ( .A1(n13143), .A2(n11032), .ZN(n11033) );
  OAI211_X1 U13502 ( .C1(n13140), .C2(n14800), .A(n11034), .B(n11033), .ZN(
        n11035) );
  AOI21_X1 U13503 ( .B1(n13135), .B2(n14803), .A(n11035), .ZN(n11036) );
  OAI21_X1 U13504 ( .B1(n13182), .B2(n14799), .A(n11036), .ZN(P2_U3260) );
  XNOR2_X1 U13505 ( .A(n11038), .B(n11037), .ZN(n14806) );
  INV_X1 U13506 ( .A(n14806), .ZN(n11053) );
  OAI21_X1 U13507 ( .B1(n11041), .B2(n11040), .A(n11039), .ZN(n11042) );
  NAND2_X1 U13508 ( .A1(n11042), .A2(n13169), .ZN(n11044) );
  AOI22_X1 U13509 ( .A1(n13153), .A2(n12892), .B1(n13152), .B2(n12894), .ZN(
        n11043) );
  NAND2_X1 U13510 ( .A1(n11044), .A2(n11043), .ZN(n14811) );
  XNOR2_X1 U13511 ( .A(n11045), .B(n14808), .ZN(n11046) );
  NAND2_X1 U13512 ( .A1(n11046), .A2(n9578), .ZN(n14807) );
  AOI22_X1 U13513 ( .A1(n13187), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n11047), 
        .B2(n13175), .ZN(n11050) );
  NAND2_X1 U13514 ( .A1(n13143), .A2(n11048), .ZN(n11049) );
  OAI211_X1 U13515 ( .C1(n14807), .C2(n13140), .A(n11050), .B(n11049), .ZN(
        n11051) );
  AOI21_X1 U13516 ( .B1(n13135), .B2(n14811), .A(n11051), .ZN(n11052) );
  OAI21_X1 U13517 ( .B1(n13182), .B2(n11053), .A(n11052), .ZN(P2_U3259) );
  NAND2_X1 U13518 ( .A1(n11012), .A2(n11054), .ZN(n11055) );
  NAND2_X1 U13519 ( .A1(n11055), .A2(n12177), .ZN(n11057) );
  NAND2_X1 U13520 ( .A1(n11057), .A2(n11056), .ZN(n11058) );
  NAND2_X1 U13521 ( .A1(n11058), .A2(n14948), .ZN(n11062) );
  OR2_X1 U13522 ( .A1(n11117), .A2(n12055), .ZN(n11060) );
  NAND2_X1 U13523 ( .A1(n12325), .A2(n12069), .ZN(n11059) );
  NAND2_X1 U13524 ( .A1(n11060), .A2(n11059), .ZN(n11121) );
  INV_X1 U13525 ( .A(n11121), .ZN(n11061) );
  NAND2_X1 U13526 ( .A1(n11062), .A2(n11061), .ZN(n15012) );
  INV_X1 U13527 ( .A(n15012), .ZN(n11068) );
  XNOR2_X1 U13528 ( .A(n11063), .B(n12177), .ZN(n15008) );
  AOI22_X1 U13529 ( .A1(n12618), .A2(n15009), .B1(n11120), .B2(n14959), .ZN(
        n11064) );
  OAI21_X1 U13530 ( .B1(n11065), .B2(n14963), .A(n11064), .ZN(n11066) );
  AOI21_X1 U13531 ( .B1(n15008), .B2(n12492), .A(n11066), .ZN(n11067) );
  OAI21_X1 U13532 ( .B1(n11068), .B2(n14965), .A(n11067), .ZN(P3_U3225) );
  AOI21_X1 U13533 ( .B1(n13064), .B2(n14839), .A(n14768), .ZN(n11069) );
  AOI21_X1 U13534 ( .B1(n13153), .B2(n12898), .A(n11069), .ZN(n14769) );
  INV_X1 U13535 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11070) );
  OAI22_X1 U13536 ( .A1(n13187), .A2(n14769), .B1(n11070), .B2(n13133), .ZN(
        n11071) );
  AOI21_X1 U13537 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n13187), .A(n11071), .ZN(
        n11073) );
  NAND2_X1 U13538 ( .A1(n13185), .A2(n9578), .ZN(n12953) );
  INV_X1 U13539 ( .A(n12953), .ZN(n11570) );
  OAI21_X1 U13540 ( .B1(n11570), .B2(n13143), .A(n14773), .ZN(n11072) );
  OAI211_X1 U13541 ( .C1(n14768), .C2(n13163), .A(n11073), .B(n11072), .ZN(
        P2_U3265) );
  NAND2_X1 U13542 ( .A1(n11075), .A2(n11074), .ZN(n13767) );
  INV_X2 U13543 ( .A(n14543), .ZN(n14545) );
  INV_X1 U13544 ( .A(n11076), .ZN(n11081) );
  INV_X1 U13545 ( .A(n14528), .ZN(n11077) );
  INV_X1 U13546 ( .A(n13952), .ZN(n14542) );
  INV_X1 U13547 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n13447) );
  AOI22_X1 U13548 ( .A1(n14545), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n14542), 
        .B2(n13447), .ZN(n11078) );
  OAI21_X1 U13549 ( .B1(n13958), .B2(n11079), .A(n11078), .ZN(n11080) );
  AOI21_X1 U13550 ( .B1(n14511), .B2(n11081), .A(n11080), .ZN(n11082) );
  OAI21_X1 U13551 ( .B1(n11083), .B2(n14545), .A(n11082), .ZN(P1_U3290) );
  INV_X1 U13552 ( .A(n10726), .ZN(n11087) );
  INV_X1 U13553 ( .A(n11084), .ZN(n11086) );
  OAI33_X1 U13554 ( .A1(n12858), .A2(n11087), .A3(n7196), .B1(n12872), .B2(
        n11086), .B3(n11085), .ZN(n11096) );
  AND2_X1 U13555 ( .A1(n12871), .A2(n14829), .ZN(n11094) );
  NAND2_X1 U13556 ( .A1(n13153), .A2(n12889), .ZN(n11089) );
  NAND2_X1 U13557 ( .A1(n13152), .A2(n12891), .ZN(n11088) );
  AND2_X1 U13558 ( .A1(n11089), .A2(n11088), .ZN(n11204) );
  INV_X1 U13559 ( .A(n11211), .ZN(n11090) );
  OR2_X1 U13560 ( .A1(n12856), .A2(n11090), .ZN(n11092) );
  OAI211_X1 U13561 ( .C1(n12828), .C2(n11204), .A(n11092), .B(n11091), .ZN(
        n11093) );
  AOI211_X1 U13562 ( .C1(n11096), .C2(n11095), .A(n11094), .B(n11093), .ZN(
        n11097) );
  OAI21_X1 U13563 ( .B1(n11098), .B2(n12858), .A(n11097), .ZN(P2_U3203) );
  INV_X1 U13564 ( .A(n11099), .ZN(n11106) );
  AOI22_X1 U13565 ( .A1(n14545), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n11100), 
        .B2(n14542), .ZN(n11101) );
  OAI21_X1 U13566 ( .B1(n13958), .B2(n11102), .A(n11101), .ZN(n11103) );
  AOI21_X1 U13567 ( .B1(n11104), .B2(n14511), .A(n11103), .ZN(n11105) );
  OAI21_X1 U13568 ( .B1(n11106), .B2(n14545), .A(n11105), .ZN(P1_U3287) );
  INV_X1 U13569 ( .A(n11107), .ZN(n11114) );
  NOR2_X1 U13570 ( .A1(n13958), .A2(n11108), .ZN(n11111) );
  OAI22_X1 U13571 ( .A1(n14543), .A2(n9953), .B1(n11109), .B2(n13952), .ZN(
        n11110) );
  AOI211_X1 U13572 ( .C1(n11112), .C2(n14511), .A(n11111), .B(n11110), .ZN(
        n11113) );
  OAI21_X1 U13573 ( .B1(n11114), .B2(n14545), .A(n11113), .ZN(P1_U3286) );
  MUX2_X1 U13574 ( .A(n11117), .B(n11116), .S(n11115), .Z(n11119) );
  XNOR2_X1 U13575 ( .A(n11119), .B(n11118), .ZN(n11126) );
  INV_X1 U13576 ( .A(n11120), .ZN(n11124) );
  NAND2_X1 U13577 ( .A1(n11121), .A2(n14884), .ZN(n11123) );
  AOI22_X1 U13578 ( .A1(n12062), .A2(n15009), .B1(P3_REG3_REG_8__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11122) );
  OAI211_X1 U13579 ( .C1(n14893), .C2(n11124), .A(n11123), .B(n11122), .ZN(
        n11125) );
  AOI21_X1 U13580 ( .B1(n11126), .B2(n14257), .A(n11125), .ZN(n11127) );
  INV_X1 U13581 ( .A(n11127), .ZN(P3_U3161) );
  OAI21_X1 U13582 ( .B1(n11130), .B2(n11129), .A(n11128), .ZN(n14999) );
  OAI22_X1 U13583 ( .A1(n12489), .A2(n14995), .B1(n11131), .B2(n11656), .ZN(
        n11138) );
  OAI211_X1 U13584 ( .C1(n11133), .C2(n12112), .A(n11132), .B(n14948), .ZN(
        n11136) );
  INV_X1 U13585 ( .A(n11134), .ZN(n11135) );
  NAND2_X1 U13586 ( .A1(n11136), .A2(n11135), .ZN(n14997) );
  MUX2_X1 U13587 ( .A(n14997), .B(P3_REG2_REG_6__SCAN_IN), .S(n14965), .Z(
        n11137) );
  AOI211_X1 U13588 ( .C1(n12492), .C2(n14999), .A(n11138), .B(n11137), .ZN(
        n11139) );
  INV_X1 U13589 ( .A(n11139), .ZN(P3_U3227) );
  INV_X1 U13590 ( .A(n14842), .ZN(n11147) );
  OAI211_X1 U13591 ( .C1(n11141), .C2(n6600), .A(n11140), .B(n12865), .ZN(
        n11146) );
  OAI22_X1 U13592 ( .A1(n12828), .A2(n11142), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15072), .ZN(n11143) );
  AOI21_X1 U13593 ( .B1(n11144), .B2(n12867), .A(n11143), .ZN(n11145) );
  OAI211_X1 U13594 ( .C1(n11147), .C2(n12829), .A(n11146), .B(n11145), .ZN(
        P2_U3189) );
  XNOR2_X1 U13595 ( .A(n11148), .B(n7815), .ZN(n14850) );
  INV_X1 U13596 ( .A(n14850), .ZN(n11166) );
  NAND2_X1 U13597 ( .A1(n11150), .A2(n11149), .ZN(n11151) );
  NAND2_X1 U13598 ( .A1(n11152), .A2(n11151), .ZN(n11153) );
  NAND2_X1 U13599 ( .A1(n11153), .A2(n13169), .ZN(n11156) );
  NAND2_X1 U13600 ( .A1(n13153), .A2(n12887), .ZN(n11155) );
  NAND2_X1 U13601 ( .A1(n13152), .A2(n12889), .ZN(n11154) );
  AND2_X1 U13602 ( .A1(n11155), .A2(n11154), .ZN(n11261) );
  NAND2_X1 U13603 ( .A1(n11156), .A2(n11261), .ZN(n14855) );
  NAND2_X1 U13604 ( .A1(n11157), .A2(n11253), .ZN(n11158) );
  NAND2_X1 U13605 ( .A1(n11158), .A2(n9578), .ZN(n11159) );
  OR2_X1 U13606 ( .A1(n11159), .A2(n11562), .ZN(n14851) );
  INV_X1 U13607 ( .A(n11263), .ZN(n11160) );
  OAI22_X1 U13608 ( .A1(n13135), .A2(n11161), .B1(n11160), .B2(n13133), .ZN(
        n11162) );
  AOI21_X1 U13609 ( .B1(n13143), .B2(n11253), .A(n11162), .ZN(n11163) );
  OAI21_X1 U13610 ( .B1(n14851), .B2(n13140), .A(n11163), .ZN(n11164) );
  AOI21_X1 U13611 ( .B1(n14855), .B2(n13135), .A(n11164), .ZN(n11165) );
  OAI21_X1 U13612 ( .B1(n13182), .B2(n11166), .A(n11165), .ZN(P2_U3254) );
  MUX2_X1 U13613 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n11167), .S(n14543), .Z(
        n11168) );
  INV_X1 U13614 ( .A(n11168), .ZN(n11172) );
  AOI22_X1 U13615 ( .A1(n14501), .A2(n11170), .B1(n14542), .B2(n11169), .ZN(
        n11171) );
  OAI211_X1 U13616 ( .C1(n13899), .C2(n11173), .A(n11172), .B(n11171), .ZN(
        P1_U3288) );
  NAND2_X1 U13617 ( .A1(n11175), .A2(n11174), .ZN(n11177) );
  OR2_X1 U13618 ( .A1(n11185), .A2(n13594), .ZN(n11176) );
  NAND2_X1 U13619 ( .A1(n11177), .A2(n11176), .ZN(n11349) );
  NAND2_X1 U13620 ( .A1(n11349), .A2(n11351), .ZN(n11179) );
  OR2_X1 U13621 ( .A1(n14575), .A2(n13593), .ZN(n11178) );
  NAND2_X1 U13622 ( .A1(n11179), .A2(n11178), .ZN(n11527) );
  XNOR2_X1 U13623 ( .A(n11527), .B(n11526), .ZN(n11195) );
  OAI22_X1 U13624 ( .A1(n11181), .A2(n14533), .B1(n11407), .B2(n14523), .ZN(
        n11194) );
  NAND2_X1 U13625 ( .A1(n11183), .A2(n11182), .ZN(n11187) );
  NAND2_X1 U13626 ( .A1(n11185), .A2(n11184), .ZN(n11186) );
  NAND2_X1 U13627 ( .A1(n11187), .A2(n11186), .ZN(n11350) );
  INV_X1 U13628 ( .A(n11350), .ZN(n11189) );
  NAND2_X1 U13629 ( .A1(n11191), .A2(n11526), .ZN(n11192) );
  AOI21_X1 U13630 ( .B1(n11537), .B2(n11192), .A(n14548), .ZN(n11193) );
  AOI211_X1 U13631 ( .C1(n11195), .C2(n14588), .A(n11194), .B(n11193), .ZN(
        n11328) );
  INV_X1 U13632 ( .A(n14575), .ZN(n11359) );
  NAND2_X1 U13633 ( .A1(n11362), .A2(n11535), .ZN(n14505) );
  OAI211_X1 U13634 ( .C1(n11362), .C2(n11535), .A(n14508), .B(n14505), .ZN(
        n11323) );
  AND2_X1 U13635 ( .A1(n11328), .A2(n11323), .ZN(n11200) );
  INV_X1 U13636 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11196) );
  OAI22_X1 U13637 ( .A1(n11535), .A2(n14077), .B1(n14589), .B2(n11196), .ZN(
        n11197) );
  INV_X1 U13638 ( .A(n11197), .ZN(n11198) );
  OAI21_X1 U13639 ( .B1(n11200), .B2(n6712), .A(n11198), .ZN(P1_U3486) );
  INV_X1 U13640 ( .A(n14032), .ZN(n11574) );
  AOI22_X1 U13641 ( .A1(n11326), .A2(n11574), .B1(n14595), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n11199) );
  OAI21_X1 U13642 ( .B1(n11200), .B2(n14595), .A(n11199), .ZN(P1_U3537) );
  OAI211_X1 U13643 ( .C1(n11203), .C2(n11202), .A(n11201), .B(n13169), .ZN(
        n11205) );
  NAND2_X1 U13644 ( .A1(n11205), .A2(n11204), .ZN(n14834) );
  INV_X1 U13645 ( .A(n14834), .ZN(n11216) );
  OAI21_X1 U13646 ( .B1(n11208), .B2(n11207), .A(n11206), .ZN(n14832) );
  INV_X1 U13647 ( .A(n14832), .ZN(n14835) );
  INV_X1 U13648 ( .A(n13182), .ZN(n13122) );
  OAI211_X1 U13649 ( .C1(n11229), .C2(n11210), .A(n11209), .B(n13136), .ZN(
        n14830) );
  AOI22_X1 U13650 ( .A1(n13187), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n11211), 
        .B2(n13175), .ZN(n11213) );
  NAND2_X1 U13651 ( .A1(n13143), .A2(n14829), .ZN(n11212) );
  OAI211_X1 U13652 ( .C1(n14830), .C2(n13140), .A(n11213), .B(n11212), .ZN(
        n11214) );
  AOI21_X1 U13653 ( .B1(n14835), .B2(n13122), .A(n11214), .ZN(n11215) );
  OAI21_X1 U13654 ( .B1(n11216), .B2(n13187), .A(n11215), .ZN(P2_U3256) );
  NAND2_X1 U13655 ( .A1(n11218), .A2(n11217), .ZN(n11219) );
  NAND3_X1 U13656 ( .A1(n11220), .A2(n13169), .A3(n11219), .ZN(n11222) );
  NAND2_X1 U13657 ( .A1(n11222), .A2(n11221), .ZN(n14827) );
  INV_X1 U13658 ( .A(n14827), .ZN(n11237) );
  NAND2_X1 U13659 ( .A1(n11224), .A2(n11223), .ZN(n11225) );
  NAND2_X1 U13660 ( .A1(n11226), .A2(n11225), .ZN(n14823) );
  INV_X1 U13661 ( .A(n14823), .ZN(n11235) );
  NAND2_X1 U13662 ( .A1(n11244), .A2(n11227), .ZN(n11228) );
  NAND2_X1 U13663 ( .A1(n11228), .A2(n13136), .ZN(n11230) );
  OR2_X1 U13664 ( .A1(n11230), .A2(n11229), .ZN(n14821) );
  AOI22_X1 U13665 ( .A1(n13187), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n11231), 
        .B2(n13175), .ZN(n11233) );
  OR2_X1 U13666 ( .A1(n13178), .A2(n14822), .ZN(n11232) );
  OAI211_X1 U13667 ( .C1(n14821), .C2(n13140), .A(n11233), .B(n11232), .ZN(
        n11234) );
  AOI21_X1 U13668 ( .B1(n11235), .B2(n13122), .A(n11234), .ZN(n11236) );
  OAI21_X1 U13669 ( .B1(n11237), .B2(n13187), .A(n11236), .ZN(P2_U3257) );
  XNOR2_X1 U13670 ( .A(n11239), .B(n11238), .ZN(n11241) );
  AOI21_X1 U13671 ( .B1(n11241), .B2(n13169), .A(n11240), .ZN(n14816) );
  XNOR2_X1 U13672 ( .A(n11243), .B(n11242), .ZN(n14819) );
  INV_X1 U13673 ( .A(n11247), .ZN(n14815) );
  INV_X1 U13674 ( .A(n11244), .ZN(n11245) );
  AOI211_X1 U13675 ( .C1(n11247), .C2(n11246), .A(n13190), .B(n11245), .ZN(
        n14813) );
  NAND2_X1 U13676 ( .A1(n14813), .A2(n13185), .ZN(n11250) );
  AOI22_X1 U13677 ( .A1(n13187), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n11248), 
        .B2(n13175), .ZN(n11249) );
  OAI211_X1 U13678 ( .C1(n14815), .C2(n13178), .A(n11250), .B(n11249), .ZN(
        n11251) );
  AOI21_X1 U13679 ( .B1(n14819), .B2(n13122), .A(n11251), .ZN(n11252) );
  OAI21_X1 U13680 ( .B1(n13187), .B2(n14816), .A(n11252), .ZN(P2_U3258) );
  INV_X1 U13681 ( .A(n11254), .ZN(n11255) );
  AOI21_X1 U13682 ( .B1(n11140), .B2(n11255), .A(n12858), .ZN(n11260) );
  NOR3_X1 U13683 ( .A1(n12872), .A2(n11257), .A3(n11256), .ZN(n11259) );
  OAI21_X1 U13684 ( .B1(n11260), .B2(n11259), .A(n11258), .ZN(n11265) );
  NAND2_X1 U13685 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n12900)
         );
  OAI21_X1 U13686 ( .B1(n12828), .B2(n11261), .A(n12900), .ZN(n11262) );
  AOI21_X1 U13687 ( .B1(n11263), .B2(n12867), .A(n11262), .ZN(n11264) );
  OAI211_X1 U13688 ( .C1(n6821), .C2(n12829), .A(n11265), .B(n11264), .ZN(
        P2_U3208) );
  XNOR2_X1 U13689 ( .A(n11267), .B(n11266), .ZN(n14795) );
  NAND3_X1 U13690 ( .A1(n10819), .A2(n11269), .A3(n11268), .ZN(n11270) );
  AND2_X1 U13691 ( .A1(n11271), .A2(n11270), .ZN(n11272) );
  OAI222_X1 U13692 ( .A1(n13069), .A2(n11274), .B1(n13067), .B2(n11273), .C1(
        n13064), .C2(n11272), .ZN(n14791) );
  AOI22_X1 U13693 ( .A1(n13187), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n11275), 
        .B2(n13175), .ZN(n11279) );
  AOI211_X1 U13694 ( .C1(n14793), .C2(n11277), .A(n13190), .B(n11276), .ZN(
        n14792) );
  NAND2_X1 U13695 ( .A1(n13185), .A2(n14792), .ZN(n11278) );
  OAI211_X1 U13696 ( .C1(n11280), .C2(n13178), .A(n11279), .B(n11278), .ZN(
        n11281) );
  AOI21_X1 U13697 ( .B1(n13135), .B2(n14791), .A(n11281), .ZN(n11282) );
  OAI21_X1 U13698 ( .B1(n13182), .B2(n14795), .A(n11282), .ZN(P2_U3261) );
  NAND2_X1 U13699 ( .A1(n14575), .A2(n13465), .ZN(n11284) );
  OR2_X1 U13700 ( .A1(n11407), .A2(n6486), .ZN(n11283) );
  NAND2_X1 U13701 ( .A1(n11284), .A2(n11283), .ZN(n11285) );
  XNOR2_X1 U13702 ( .A(n11285), .B(n13404), .ZN(n11399) );
  NOR2_X1 U13703 ( .A1(n11407), .A2(n13360), .ZN(n11286) );
  AOI21_X1 U13704 ( .B1(n14575), .B2(n13462), .A(n11286), .ZN(n11398) );
  XNOR2_X1 U13705 ( .A(n11399), .B(n11398), .ZN(n11296) );
  INV_X1 U13706 ( .A(n11287), .ZN(n11288) );
  NAND2_X1 U13707 ( .A1(n11289), .A2(n11288), .ZN(n11290) );
  NAND2_X1 U13708 ( .A1(n11291), .A2(n11290), .ZN(n11295) );
  INV_X1 U13709 ( .A(n11295), .ZN(n11293) );
  INV_X1 U13710 ( .A(n11401), .ZN(n11294) );
  AOI21_X1 U13711 ( .B1(n11296), .B2(n11295), .A(n11294), .ZN(n11302) );
  INV_X1 U13712 ( .A(n14326), .ZN(n13577) );
  OAI21_X1 U13713 ( .B1(n14325), .B2(n11528), .A(n11297), .ZN(n11298) );
  AOI21_X1 U13714 ( .B1(n13577), .B2(n13594), .A(n11298), .ZN(n11299) );
  OAI21_X1 U13715 ( .B1(n14339), .B2(n11357), .A(n11299), .ZN(n11300) );
  AOI21_X1 U13716 ( .B1(n14575), .B2(n14335), .A(n11300), .ZN(n11301) );
  OAI21_X1 U13717 ( .B1(n11302), .B2(n14330), .A(n11301), .ZN(P1_U3221) );
  INV_X1 U13718 ( .A(n11303), .ZN(n11304) );
  OAI222_X1 U13719 ( .A1(n11305), .A2(P3_U3151), .B1(n14215), .B2(n11304), 
        .C1(n6793), .C2(n14213), .ZN(P3_U3271) );
  XNOR2_X1 U13720 ( .A(n11306), .B(n11311), .ZN(n11309) );
  INV_X1 U13721 ( .A(n11307), .ZN(n11308) );
  OAI21_X1 U13722 ( .B1(n11309), .B2(n14548), .A(n11308), .ZN(n14570) );
  INV_X1 U13723 ( .A(n14570), .ZN(n11322) );
  XNOR2_X1 U13724 ( .A(n11310), .B(n11311), .ZN(n14572) );
  NAND2_X1 U13725 ( .A1(n14543), .A2(n14588), .ZN(n13963) );
  OAI21_X1 U13726 ( .B1(n11312), .B2(n14569), .A(n14508), .ZN(n11313) );
  OR2_X1 U13727 ( .A1(n11314), .A2(n11313), .ZN(n14568) );
  OAI22_X1 U13728 ( .A1(n14543), .A2(n11316), .B1(n11315), .B2(n13952), .ZN(
        n11317) );
  AOI21_X1 U13729 ( .B1(n14501), .B2(n11318), .A(n11317), .ZN(n11319) );
  OAI21_X1 U13730 ( .B1(n13899), .B2(n14568), .A(n11319), .ZN(n11320) );
  AOI21_X1 U13731 ( .B1(n14572), .B2(n14512), .A(n11320), .ZN(n11321) );
  OAI21_X1 U13732 ( .B1(n11322), .B2(n14545), .A(n11321), .ZN(P1_U3289) );
  OAI22_X1 U13733 ( .A1(n14543), .A2(n9954), .B1(n11405), .B2(n13952), .ZN(
        n11325) );
  NOR2_X1 U13734 ( .A1(n11323), .A2(n13899), .ZN(n11324) );
  AOI211_X1 U13735 ( .C1(n14501), .C2(n11326), .A(n11325), .B(n11324), .ZN(
        n11327) );
  OAI21_X1 U13736 ( .B1(n11328), .B2(n14545), .A(n11327), .ZN(P1_U3284) );
  XNOR2_X1 U13737 ( .A(n11330), .B(n11329), .ZN(n11332) );
  AOI21_X1 U13738 ( .B1(n11332), .B2(n14519), .A(n11331), .ZN(n14563) );
  XNOR2_X1 U13739 ( .A(n11334), .B(n11333), .ZN(n14566) );
  INV_X1 U13740 ( .A(n14517), .ZN(n11337) );
  INV_X1 U13741 ( .A(n11335), .ZN(n11336) );
  OAI211_X1 U13742 ( .C1(n14564), .C2(n11337), .A(n11336), .B(n14508), .ZN(
        n14562) );
  OAI22_X1 U13743 ( .A1(n14543), .A2(n8108), .B1(n13617), .B2(n13952), .ZN(
        n11338) );
  AOI21_X1 U13744 ( .B1(n14501), .B2(n11339), .A(n11338), .ZN(n11340) );
  OAI21_X1 U13745 ( .B1(n13899), .B2(n14562), .A(n11340), .ZN(n11341) );
  AOI21_X1 U13746 ( .B1(n14512), .B2(n14566), .A(n11341), .ZN(n11342) );
  OAI21_X1 U13747 ( .B1(n14545), .B2(n14563), .A(n11342), .ZN(P1_U3291) );
  INV_X1 U13748 ( .A(n11343), .ZN(n11348) );
  NAND2_X1 U13749 ( .A1(n14081), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11345) );
  OAI211_X1 U13750 ( .C1(n11348), .C2(n14083), .A(n11345), .B(n11344), .ZN(
        P1_U3332) );
  NAND2_X1 U13751 ( .A1(n13299), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n11347) );
  OAI211_X1 U13752 ( .C1(n11348), .C2(n6452), .A(n11347), .B(n11346), .ZN(
        P2_U3304) );
  XNOR2_X1 U13753 ( .A(n11349), .B(n11351), .ZN(n14580) );
  INV_X1 U13754 ( .A(n14580), .ZN(n11367) );
  AOI21_X1 U13755 ( .B1(n11350), .B2(n11351), .A(n14548), .ZN(n11353) );
  NAND2_X1 U13756 ( .A1(n11353), .A2(n11352), .ZN(n14578) );
  INV_X1 U13757 ( .A(n14578), .ZN(n11356) );
  OR2_X1 U13758 ( .A1(n11528), .A2(n14533), .ZN(n11355) );
  NAND2_X1 U13759 ( .A1(n13594), .A2(n13929), .ZN(n11354) );
  NAND2_X1 U13760 ( .A1(n11355), .A2(n11354), .ZN(n14573) );
  OAI21_X1 U13761 ( .B1(n11356), .B2(n14573), .A(n14543), .ZN(n11366) );
  OAI22_X1 U13762 ( .A1(n14543), .A2(n11358), .B1(n11357), .B2(n13952), .ZN(
        n11364) );
  OAI21_X1 U13763 ( .B1(n11360), .B2(n11359), .A(n14508), .ZN(n11361) );
  OR2_X1 U13764 ( .A1(n11362), .A2(n11361), .ZN(n14576) );
  NOR2_X1 U13765 ( .A1(n14576), .A2(n13899), .ZN(n11363) );
  AOI211_X1 U13766 ( .C1(n14501), .C2(n14575), .A(n11364), .B(n11363), .ZN(
        n11365) );
  OAI211_X1 U13767 ( .C1(n11367), .C2(n13963), .A(n11366), .B(n11365), .ZN(
        P1_U3285) );
  XNOR2_X1 U13768 ( .A(n11368), .B(n6868), .ZN(n11370) );
  NAND2_X1 U13769 ( .A1(n12322), .A2(n12069), .ZN(n11369) );
  OAI21_X1 U13770 ( .B1(n11385), .B2(n12055), .A(n11369), .ZN(n11392) );
  AOI21_X1 U13771 ( .B1(n11370), .B2(n14948), .A(n11392), .ZN(n14315) );
  XNOR2_X1 U13772 ( .A(n11371), .B(n12190), .ZN(n14313) );
  AOI22_X1 U13773 ( .A1(n14965), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n14959), 
        .B2(n11391), .ZN(n11372) );
  OAI21_X1 U13774 ( .B1(n12187), .B2(n12489), .A(n11372), .ZN(n11373) );
  AOI21_X1 U13775 ( .B1(n14313), .B2(n12492), .A(n11373), .ZN(n11374) );
  OAI21_X1 U13776 ( .B1(n14315), .B2(n14965), .A(n11374), .ZN(P3_U3222) );
  XNOR2_X1 U13777 ( .A(n11375), .B(n8933), .ZN(n15019) );
  INV_X1 U13778 ( .A(n15019), .ZN(n15021) );
  AOI21_X1 U13779 ( .B1(n11376), .B2(n12182), .A(n14939), .ZN(n11378) );
  AOI21_X1 U13780 ( .B1(n11378), .B2(n11413), .A(n11377), .ZN(n15017) );
  AOI22_X1 U13781 ( .A1(n14965), .A2(P3_REG2_REG_9__SCAN_IN), .B1(n14959), 
        .B2(n11379), .ZN(n11381) );
  NAND2_X1 U13782 ( .A1(n12618), .A2(n15015), .ZN(n11380) );
  OAI211_X1 U13783 ( .C1(n15017), .C2(n14965), .A(n11381), .B(n11380), .ZN(
        n11382) );
  AOI21_X1 U13784 ( .B1(n12492), .B2(n15021), .A(n11382), .ZN(n11383) );
  INV_X1 U13785 ( .A(n11383), .ZN(P3_U3224) );
  XNOR2_X1 U13786 ( .A(n12187), .B(n11980), .ZN(n11513) );
  XNOR2_X1 U13787 ( .A(n11384), .B(n11931), .ZN(n11389) );
  XNOR2_X1 U13788 ( .A(n11389), .B(n11385), .ZN(n14878) );
  INV_X1 U13789 ( .A(n11386), .ZN(n11387) );
  INV_X1 U13790 ( .A(n12325), .ZN(n12137) );
  NAND2_X1 U13791 ( .A1(n11387), .A2(n12137), .ZN(n14879) );
  AND2_X1 U13792 ( .A1(n14878), .A2(n14879), .ZN(n11388) );
  NAND2_X1 U13793 ( .A1(n14880), .A2(n11388), .ZN(n14877) );
  NAND2_X1 U13794 ( .A1(n12324), .A2(n11389), .ZN(n11390) );
  NAND2_X1 U13795 ( .A1(n14877), .A2(n11390), .ZN(n11514) );
  XOR2_X1 U13796 ( .A(n11513), .B(n11514), .Z(n11515) );
  XNOR2_X1 U13797 ( .A(n11515), .B(n12323), .ZN(n11397) );
  INV_X1 U13798 ( .A(n11391), .ZN(n11394) );
  NAND2_X1 U13799 ( .A1(n11392), .A2(n14884), .ZN(n11393) );
  NAND2_X1 U13800 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n14898)
         );
  OAI211_X1 U13801 ( .C1(n11394), .C2(n14893), .A(n11393), .B(n14898), .ZN(
        n11395) );
  AOI21_X1 U13802 ( .B1(n14312), .B2(n12062), .A(n11395), .ZN(n11396) );
  OAI21_X1 U13803 ( .B1(n11397), .B2(n14881), .A(n11396), .ZN(P3_U3176) );
  NAND2_X1 U13804 ( .A1(n11399), .A2(n11398), .ZN(n11400) );
  OAI22_X1 U13805 ( .A1(n11535), .A2(n10594), .B1(n11528), .B2(n6486), .ZN(
        n11402) );
  XNOR2_X1 U13806 ( .A(n11402), .B(n13404), .ZN(n11481) );
  OAI22_X1 U13807 ( .A1(n11535), .A2(n6486), .B1(n11528), .B2(n13360), .ZN(
        n11482) );
  XNOR2_X1 U13808 ( .A(n11481), .B(n11482), .ZN(n11403) );
  OAI211_X1 U13809 ( .C1(n11404), .C2(n11403), .A(n11485), .B(n13570), .ZN(
        n11411) );
  INV_X1 U13810 ( .A(n11405), .ZN(n11409) );
  AOI22_X1 U13811 ( .A1(n13567), .A2(n13591), .B1(P1_REG3_REG_9__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11406) );
  OAI21_X1 U13812 ( .B1(n11407), .B2(n14326), .A(n11406), .ZN(n11408) );
  AOI21_X1 U13813 ( .B1(n11409), .B2(n13562), .A(n11408), .ZN(n11410) );
  OAI211_X1 U13814 ( .C1(n11535), .C2(n13580), .A(n11411), .B(n11410), .ZN(
        P1_U3231) );
  XNOR2_X1 U13815 ( .A(n11412), .B(n12184), .ZN(n11428) );
  INV_X1 U13816 ( .A(n12184), .ZN(n12118) );
  NAND3_X1 U13817 ( .A1(n11413), .A2(n12118), .A3(n12135), .ZN(n11414) );
  AND3_X1 U13818 ( .A1(n11415), .A2(n14948), .A3(n11414), .ZN(n11417) );
  NAND2_X1 U13819 ( .A1(n12325), .A2(n12300), .ZN(n11416) );
  OAI21_X1 U13820 ( .B1(n11459), .B2(n12057), .A(n11416), .ZN(n14885) );
  OR2_X1 U13821 ( .A1(n11417), .A2(n14885), .ZN(n11426) );
  AOI22_X1 U13822 ( .A1(n14965), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n14959), 
        .B2(n11418), .ZN(n11419) );
  OAI21_X1 U13823 ( .B1(n14888), .B2(n12489), .A(n11419), .ZN(n11420) );
  AOI21_X1 U13824 ( .B1(n11426), .B2(n14963), .A(n11420), .ZN(n11421) );
  OAI21_X1 U13825 ( .B1(n12621), .B2(n11428), .A(n11421), .ZN(P3_U3223) );
  INV_X1 U13826 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n11422) );
  OAI22_X1 U13827 ( .A1(n12730), .A2(n14888), .B1(n15025), .B2(n11422), .ZN(
        n11423) );
  AOI21_X1 U13828 ( .B1(n11426), .B2(n15025), .A(n11423), .ZN(n11424) );
  OAI21_X1 U13829 ( .B1(n11428), .B2(n12748), .A(n11424), .ZN(P3_U3420) );
  OAI22_X1 U13830 ( .A1(n12655), .A2(n14888), .B1(n15034), .B2(n10963), .ZN(
        n11425) );
  AOI21_X1 U13831 ( .B1(n11426), .B2(n15034), .A(n11425), .ZN(n11427) );
  OAI21_X1 U13832 ( .B1(n11428), .B2(n12664), .A(n11427), .ZN(P3_U3469) );
  INV_X1 U13833 ( .A(n11429), .ZN(n11434) );
  OAI222_X1 U13834 ( .A1(n14085), .A2(n11431), .B1(n14088), .B2(n11434), .C1(
        P1_U3086), .C2(n11430), .ZN(P1_U3331) );
  INV_X1 U13835 ( .A(n11432), .ZN(n11433) );
  OAI222_X1 U13836 ( .A1(n13314), .A2(n11435), .B1(n6452), .B2(n11434), .C1(
        n11433), .C2(P2_U3088), .ZN(P2_U3303) );
  INV_X1 U13837 ( .A(n11258), .ZN(n11438) );
  NOR3_X1 U13838 ( .A1(n12872), .A2(n11436), .A3(n11555), .ZN(n11437) );
  AOI21_X1 U13839 ( .B1(n11438), .B2(n12865), .A(n11437), .ZN(n11447) );
  NAND2_X1 U13840 ( .A1(n12875), .A2(n12888), .ZN(n11441) );
  AOI21_X1 U13841 ( .B1(n12867), .B2(n11564), .A(n11439), .ZN(n11440) );
  OAI211_X1 U13842 ( .C1(n11554), .C2(n12869), .A(n11441), .B(n11440), .ZN(
        n11444) );
  NOR2_X1 U13843 ( .A1(n11442), .A2(n12858), .ZN(n11443) );
  AOI211_X1 U13844 ( .C1(n13273), .C2(n12871), .A(n11444), .B(n11443), .ZN(
        n11445) );
  OAI21_X1 U13845 ( .B1(n11447), .B2(n11446), .A(n11445), .ZN(P2_U3196) );
  AOI21_X1 U13846 ( .B1(n11449), .B2(n11448), .A(n12858), .ZN(n11450) );
  NAND2_X1 U13847 ( .A1(n11450), .A2(n11895), .ZN(n11456) );
  NAND2_X1 U13848 ( .A1(n13152), .A2(n12887), .ZN(n11451) );
  OAI21_X1 U13849 ( .B1(n11452), .B2(n13069), .A(n11451), .ZN(n11471) );
  INV_X1 U13850 ( .A(n11471), .ZN(n11453) );
  OAI22_X1 U13851 ( .A1(n12828), .A2(n11453), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15172), .ZN(n11454) );
  AOI21_X1 U13852 ( .B1(n11475), .B2(n12867), .A(n11454), .ZN(n11455) );
  OAI211_X1 U13853 ( .C1(n11600), .C2(n12829), .A(n11456), .B(n11455), .ZN(
        P2_U3206) );
  XNOR2_X1 U13854 ( .A(n11457), .B(n12119), .ZN(n11460) );
  NAND2_X1 U13855 ( .A1(n12321), .A2(n12069), .ZN(n11458) );
  OAI21_X1 U13856 ( .B1(n11459), .B2(n12055), .A(n11458), .ZN(n11519) );
  AOI21_X1 U13857 ( .B1(n11460), .B2(n14948), .A(n11519), .ZN(n14311) );
  XNOR2_X1 U13858 ( .A(n11461), .B(n12119), .ZN(n14309) );
  NOR2_X1 U13859 ( .A1(n11462), .A2(n12489), .ZN(n11465) );
  INV_X1 U13860 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12337) );
  INV_X1 U13861 ( .A(n11463), .ZN(n11522) );
  OAI22_X1 U13862 ( .A1(n14963), .A2(n12337), .B1(n11522), .B2(n11656), .ZN(
        n11464) );
  AOI211_X1 U13863 ( .C1(n14309), .C2(n12492), .A(n11465), .B(n11464), .ZN(
        n11466) );
  OAI21_X1 U13864 ( .B1(n14311), .B2(n14965), .A(n11466), .ZN(P3_U3221) );
  INV_X1 U13865 ( .A(n11468), .ZN(n11469) );
  NOR2_X1 U13866 ( .A1(n11474), .A2(n11469), .ZN(n11470) );
  AOI21_X1 U13867 ( .B1(n11556), .B2(n11470), .A(n13064), .ZN(n11472) );
  AOI21_X1 U13868 ( .B1(n11467), .B2(n11472), .A(n11471), .ZN(n11599) );
  XOR2_X1 U13869 ( .A(n11474), .B(n11473), .Z(n11602) );
  NAND2_X1 U13870 ( .A1(n11602), .A2(n13122), .ZN(n11480) );
  OAI211_X1 U13871 ( .C1(n11563), .C2(n11600), .A(n9578), .B(n11704), .ZN(
        n11598) );
  INV_X1 U13872 ( .A(n11598), .ZN(n11478) );
  AOI22_X1 U13873 ( .A1(n13187), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11475), 
        .B2(n13175), .ZN(n11476) );
  OAI21_X1 U13874 ( .B1(n11600), .B2(n13178), .A(n11476), .ZN(n11477) );
  AOI21_X1 U13875 ( .B1(n11478), .B2(n13185), .A(n11477), .ZN(n11479) );
  OAI211_X1 U13876 ( .C1(n11599), .C2(n13187), .A(n11480), .B(n11479), .ZN(
        P2_U3252) );
  INV_X1 U13877 ( .A(n14502), .ZN(n14585) );
  INV_X1 U13878 ( .A(n11481), .ZN(n11483) );
  NAND2_X1 U13879 ( .A1(n11483), .A2(n11482), .ZN(n11484) );
  NAND2_X1 U13880 ( .A1(n14502), .A2(n13465), .ZN(n11487) );
  NAND2_X1 U13881 ( .A1(n13591), .A2(n13462), .ZN(n11486) );
  NAND2_X1 U13882 ( .A1(n11487), .A2(n11486), .ZN(n11488) );
  XNOR2_X1 U13883 ( .A(n11488), .B(n13463), .ZN(n11612) );
  AND2_X1 U13884 ( .A1(n13591), .A2(n10598), .ZN(n11489) );
  AOI21_X1 U13885 ( .B1(n14502), .B2(n6449), .A(n11489), .ZN(n11610) );
  XNOR2_X1 U13886 ( .A(n11612), .B(n11610), .ZN(n11490) );
  OAI211_X1 U13887 ( .C1(n11491), .C2(n11490), .A(n11614), .B(n13570), .ZN(
        n11495) );
  OR2_X1 U13888 ( .A1(n11528), .A2(n14523), .ZN(n14495) );
  NAND2_X1 U13889 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n13689)
         );
  OAI21_X1 U13890 ( .B1(n13544), .B2(n14495), .A(n13689), .ZN(n11493) );
  NOR2_X1 U13891 ( .A1(n14339), .A2(n14499), .ZN(n11492) );
  AOI211_X1 U13892 ( .C1(n13567), .C2(n14506), .A(n11493), .B(n11492), .ZN(
        n11494) );
  OAI211_X1 U13893 ( .C1(n14585), .C2(n13580), .A(n11495), .B(n11494), .ZN(
        P1_U3217) );
  INV_X1 U13894 ( .A(n11496), .ZN(n11497) );
  OAI222_X1 U13895 ( .A1(P3_U3151), .A2(n11499), .B1(n14213), .B2(n11498), 
        .C1(n14215), .C2(n11497), .ZN(P3_U3270) );
  INV_X1 U13896 ( .A(n11500), .ZN(n11504) );
  OAI222_X1 U13897 ( .A1(n14085), .A2(n11502), .B1(n14088), .B2(n11504), .C1(
        P1_U3086), .C2(n11501), .ZN(P1_U3330) );
  OAI222_X1 U13898 ( .A1(n13314), .A2(n11505), .B1(n6452), .B2(n11504), .C1(
        n11503), .C2(P2_U3088), .ZN(P2_U3302) );
  XNOR2_X1 U13899 ( .A(n14308), .B(n11980), .ZN(n11516) );
  OAI21_X1 U13900 ( .B1(n12323), .B2(n11513), .A(n12322), .ZN(n11507) );
  XNOR2_X1 U13901 ( .A(n14303), .B(n11980), .ZN(n11673) );
  XNOR2_X1 U13902 ( .A(n11673), .B(n11675), .ZN(n11508) );
  XNOR2_X1 U13903 ( .A(n11672), .B(n11508), .ZN(n11512) );
  INV_X1 U13904 ( .A(n14303), .ZN(n11592) );
  AOI22_X1 U13905 ( .A1(n12069), .A2(n12320), .B1(n12322), .B2(n12300), .ZN(
        n11586) );
  INV_X1 U13906 ( .A(n14884), .ZN(n12071) );
  NAND2_X1 U13907 ( .A1(n12073), .A2(n11588), .ZN(n11509) );
  NAND2_X1 U13908 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n14915)
         );
  OAI211_X1 U13909 ( .C1(n11586), .C2(n12071), .A(n11509), .B(n14915), .ZN(
        n11510) );
  AOI21_X1 U13910 ( .B1(n11592), .B2(n12062), .A(n11510), .ZN(n11511) );
  OAI21_X1 U13911 ( .B1(n11512), .B2(n14881), .A(n11511), .ZN(P3_U3174) );
  AOI22_X1 U13912 ( .A1(n11515), .A2(n12323), .B1(n11514), .B2(n11513), .ZN(
        n11518) );
  XNOR2_X1 U13913 ( .A(n11516), .B(n12322), .ZN(n11517) );
  XNOR2_X1 U13914 ( .A(n11518), .B(n11517), .ZN(n11524) );
  AOI22_X1 U13915 ( .A1(n11519), .A2(n14884), .B1(P3_REG3_REG_12__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11521) );
  NAND2_X1 U13916 ( .A1(n14308), .A2(n12062), .ZN(n11520) );
  OAI211_X1 U13917 ( .C1(n11522), .C2(n14893), .A(n11521), .B(n11520), .ZN(
        n11523) );
  AOI21_X1 U13918 ( .B1(n11524), .B2(n14257), .A(n11523), .ZN(n11525) );
  INV_X1 U13919 ( .A(n11525), .ZN(P3_U3164) );
  NAND2_X1 U13920 ( .A1(n11527), .A2(n11526), .ZN(n11530) );
  NAND2_X1 U13921 ( .A1(n11535), .A2(n11528), .ZN(n11529) );
  NAND2_X1 U13922 ( .A1(n11530), .A2(n11529), .ZN(n14503) );
  NAND2_X1 U13923 ( .A1(n14503), .A2(n14504), .ZN(n11532) );
  OR2_X1 U13924 ( .A1(n14502), .A2(n13591), .ZN(n11531) );
  NAND2_X1 U13925 ( .A1(n11532), .A2(n11531), .ZN(n14345) );
  NAND2_X1 U13926 ( .A1(n14345), .A2(n14346), .ZN(n11534) );
  OR2_X1 U13927 ( .A1(n14373), .A2(n14506), .ZN(n11533) );
  NAND2_X1 U13928 ( .A1(n11534), .A2(n11533), .ZN(n11638) );
  INV_X1 U13929 ( .A(n11637), .ZN(n11542) );
  XNOR2_X1 U13930 ( .A(n11638), .B(n11542), .ZN(n11545) );
  OR2_X1 U13931 ( .A1(n11535), .A2(n13592), .ZN(n11536) );
  OR2_X1 U13932 ( .A1(n14373), .A2(n11539), .ZN(n11540) );
  NAND2_X1 U13933 ( .A1(n14341), .A2(n11540), .ZN(n11541) );
  NAND2_X1 U13934 ( .A1(n11541), .A2(n11542), .ZN(n11633) );
  OAI211_X1 U13935 ( .C1(n11542), .C2(n11541), .A(n11633), .B(n14519), .ZN(
        n11544) );
  AOI22_X1 U13936 ( .A1(n13929), .A2(n14506), .B1(n13589), .B2(n14507), .ZN(
        n11543) );
  OAI211_X1 U13937 ( .C1(n11545), .C2(n14549), .A(n11544), .B(n11543), .ZN(
        n11573) );
  INV_X1 U13938 ( .A(n11573), .ZN(n11550) );
  OR2_X2 U13939 ( .A1(n14505), .A2(n14502), .ZN(n14347) );
  INV_X1 U13940 ( .A(n14349), .ZN(n11546) );
  INV_X1 U13941 ( .A(n11693), .ZN(n11702) );
  AOI211_X1 U13942 ( .C1(n11693), .C2(n11546), .A(n14526), .B(n14244), .ZN(
        n11572) );
  NOR2_X1 U13943 ( .A1(n11702), .A2(n13958), .ZN(n11548) );
  OAI22_X1 U13944 ( .A1(n14543), .A2(n13711), .B1(n11697), .B2(n13952), .ZN(
        n11547) );
  AOI211_X1 U13945 ( .C1(n11572), .C2(n14511), .A(n11548), .B(n11547), .ZN(
        n11549) );
  OAI21_X1 U13946 ( .B1(n11550), .B2(n14545), .A(n11549), .ZN(P1_U3281) );
  INV_X1 U13947 ( .A(n11551), .ZN(n11553) );
  OAI21_X1 U13948 ( .B1(n11553), .B2(n11559), .A(n11552), .ZN(n11567) );
  OAI22_X1 U13949 ( .A1(n13067), .A2(n11555), .B1(n11554), .B2(n13069), .ZN(
        n11561) );
  INV_X1 U13950 ( .A(n11556), .ZN(n11557) );
  AOI211_X1 U13951 ( .C1(n11559), .C2(n11558), .A(n13064), .B(n11557), .ZN(
        n11560) );
  AOI211_X1 U13952 ( .C1(n14836), .C2(n11567), .A(n11561), .B(n11560), .ZN(
        n13276) );
  AOI21_X1 U13953 ( .B1(n13273), .B2(n6820), .A(n11563), .ZN(n13274) );
  AOI22_X1 U13954 ( .A1(n13187), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11564), 
        .B2(n13175), .ZN(n11565) );
  OAI21_X1 U13955 ( .B1(n11566), .B2(n13178), .A(n11565), .ZN(n11569) );
  INV_X1 U13956 ( .A(n11567), .ZN(n13277) );
  NOR2_X1 U13957 ( .A1(n13277), .A2(n13163), .ZN(n11568) );
  AOI211_X1 U13958 ( .C1(n13274), .C2(n11570), .A(n11569), .B(n11568), .ZN(
        n11571) );
  OAI21_X1 U13959 ( .B1(n13276), .B2(n13187), .A(n11571), .ZN(P2_U3253) );
  NOR2_X1 U13960 ( .A1(n11573), .A2(n11572), .ZN(n11579) );
  AOI22_X1 U13961 ( .A1(n11693), .A2(n11574), .B1(n14595), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n11575) );
  OAI21_X1 U13962 ( .B1(n11579), .B2(n14595), .A(n11575), .ZN(P1_U3540) );
  INV_X1 U13963 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11576) );
  OAI22_X1 U13964 ( .A1(n11702), .A2(n14077), .B1(n14589), .B2(n11576), .ZN(
        n11577) );
  INV_X1 U13965 ( .A(n11577), .ZN(n11578) );
  OAI21_X1 U13966 ( .B1(n11579), .B2(n6712), .A(n11578), .ZN(P1_U3495) );
  INV_X1 U13967 ( .A(n11580), .ZN(n11582) );
  OAI222_X1 U13968 ( .A1(n11583), .A2(P3_U3151), .B1(n14215), .B2(n11582), 
        .C1(n11581), .C2(n14213), .ZN(P3_U3269) );
  INV_X1 U13969 ( .A(n12122), .ZN(n12203) );
  XNOR2_X1 U13970 ( .A(n11584), .B(n12203), .ZN(n14305) );
  XNOR2_X1 U13971 ( .A(n11585), .B(n12122), .ZN(n11587) );
  OAI21_X1 U13972 ( .B1(n11587), .B2(n14939), .A(n11586), .ZN(n14306) );
  NAND2_X1 U13973 ( .A1(n14306), .A2(n14963), .ZN(n11594) );
  INV_X1 U13974 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n11590) );
  INV_X1 U13975 ( .A(n11588), .ZN(n11589) );
  OAI22_X1 U13976 ( .A1(n14963), .A2(n11590), .B1(n11589), .B2(n11656), .ZN(
        n11591) );
  AOI21_X1 U13977 ( .B1(n11592), .B2(n12618), .A(n11591), .ZN(n11593) );
  OAI211_X1 U13978 ( .C1(n12621), .C2(n14305), .A(n11594), .B(n11593), .ZN(
        P3_U3220) );
  INV_X1 U13979 ( .A(n11595), .ZN(n11597) );
  OAI222_X1 U13980 ( .A1(n14215), .A2(n11597), .B1(n14213), .B2(n11596), .C1(
        P3_U3151), .C2(n12455), .ZN(P3_U3268) );
  OAI211_X1 U13981 ( .C1(n11600), .C2(n14852), .A(n11599), .B(n11598), .ZN(
        n11601) );
  AOI21_X1 U13982 ( .B1(n11602), .B2(n8001), .A(n11601), .ZN(n11605) );
  NAND2_X1 U13983 ( .A1(n14873), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11603) );
  OAI21_X1 U13984 ( .B1(n11605), .B2(n14873), .A(n11603), .ZN(P2_U3512) );
  NAND2_X1 U13985 ( .A1(n14856), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n11604) );
  OAI21_X1 U13986 ( .B1(n11605), .B2(n14856), .A(n11604), .ZN(P2_U3469) );
  NAND2_X1 U13987 ( .A1(n14373), .A2(n13465), .ZN(n11607) );
  NAND2_X1 U13988 ( .A1(n14506), .A2(n13462), .ZN(n11606) );
  NAND2_X1 U13989 ( .A1(n11607), .A2(n11606), .ZN(n11608) );
  XNOR2_X1 U13990 ( .A(n11608), .B(n13404), .ZN(n11686) );
  AND2_X1 U13991 ( .A1(n14506), .A2(n10598), .ZN(n11609) );
  AOI21_X1 U13992 ( .B1(n14373), .B2(n6449), .A(n11609), .ZN(n11685) );
  XNOR2_X1 U13993 ( .A(n11686), .B(n11685), .ZN(n11619) );
  INV_X1 U13994 ( .A(n11610), .ZN(n11611) );
  NAND2_X1 U13995 ( .A1(n11612), .A2(n11611), .ZN(n11613) );
  NAND2_X1 U13996 ( .A1(n11614), .A2(n11613), .ZN(n11618) );
  INV_X1 U13997 ( .A(n11618), .ZN(n11616) );
  INV_X1 U13998 ( .A(n11688), .ZN(n11617) );
  AOI21_X1 U13999 ( .B1(n11619), .B2(n11618), .A(n11617), .ZN(n11625) );
  NAND2_X1 U14000 ( .A1(n13591), .A2(n13929), .ZN(n11621) );
  NAND2_X1 U14001 ( .A1(n13590), .A2(n14507), .ZN(n11620) );
  NAND2_X1 U14002 ( .A1(n11621), .A2(n11620), .ZN(n14340) );
  AOI22_X1 U14003 ( .A1(n13534), .A2(n14340), .B1(P1_REG3_REG_11__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11622) );
  OAI21_X1 U14004 ( .B1(n14339), .B2(n14343), .A(n11622), .ZN(n11623) );
  AOI21_X1 U14005 ( .B1(n14373), .B2(n14335), .A(n11623), .ZN(n11624) );
  OAI21_X1 U14006 ( .B1(n11625), .B2(n14330), .A(n11624), .ZN(P1_U3236) );
  INV_X1 U14007 ( .A(n11626), .ZN(n11631) );
  INV_X1 U14008 ( .A(n11627), .ZN(n11628) );
  OAI222_X1 U14009 ( .A1(n14085), .A2(n11629), .B1(n14083), .B2(n11631), .C1(
        n11628), .C2(P1_U3086), .ZN(P1_U3329) );
  OAI222_X1 U14010 ( .A1(n11632), .A2(P2_U3088), .B1(n6452), .B2(n11631), .C1(
        n11630), .C2(n13314), .ZN(P2_U3301) );
  NAND2_X1 U14011 ( .A1(n11633), .A2(n14233), .ZN(n11634) );
  INV_X1 U14012 ( .A(n14243), .ZN(n14235) );
  NAND2_X1 U14013 ( .A1(n11634), .A2(n14235), .ZN(n14232) );
  OR2_X1 U14014 ( .A1(n14241), .A2(n14327), .ZN(n11635) );
  NAND2_X1 U14015 ( .A1(n14232), .A2(n11635), .ZN(n11636) );
  OAI211_X1 U14016 ( .C1(n11636), .C2(n11642), .A(n11763), .B(n14519), .ZN(
        n11646) );
  INV_X1 U14017 ( .A(n14324), .ZN(n13587) );
  AOI22_X1 U14018 ( .A1(n13587), .A2(n14507), .B1(n13929), .B2(n13589), .ZN(
        n11645) );
  NAND2_X1 U14019 ( .A1(n11638), .A2(n11637), .ZN(n11640) );
  OR2_X1 U14020 ( .A1(n11693), .A2(n13590), .ZN(n11639) );
  OR2_X1 U14021 ( .A1(n14241), .A2(n13589), .ZN(n11641) );
  OAI211_X1 U14022 ( .C1(n7382), .C2(n11643), .A(n14588), .B(n11759), .ZN(
        n11644) );
  NAND3_X1 U14023 ( .A1(n11646), .A2(n11645), .A3(n11644), .ZN(n11797) );
  INV_X1 U14024 ( .A(n11797), .ZN(n11651) );
  INV_X1 U14025 ( .A(n14241), .ZN(n14369) );
  INV_X1 U14026 ( .A(n11769), .ZN(n11647) );
  AOI211_X1 U14027 ( .C1(n14336), .C2(n6594), .A(n14526), .B(n11647), .ZN(
        n11796) );
  INV_X1 U14028 ( .A(n14336), .ZN(n11802) );
  NOR2_X1 U14029 ( .A1(n11802), .A2(n13958), .ZN(n11649) );
  OAI22_X1 U14030 ( .A1(n14543), .A2(n13713), .B1(n14338), .B2(n13952), .ZN(
        n11648) );
  AOI211_X1 U14031 ( .C1(n11796), .C2(n14511), .A(n11649), .B(n11648), .ZN(
        n11650) );
  OAI21_X1 U14032 ( .B1(n11651), .B2(n14545), .A(n11650), .ZN(P1_U3279) );
  XNOR2_X1 U14033 ( .A(n11652), .B(n7231), .ZN(n11654) );
  NAND2_X1 U14034 ( .A1(n12321), .A2(n12300), .ZN(n11653) );
  OAI21_X1 U14035 ( .B1(n11778), .B2(n12057), .A(n11653), .ZN(n14253) );
  AOI21_X1 U14036 ( .B1(n11654), .B2(n14948), .A(n14253), .ZN(n14297) );
  INV_X1 U14037 ( .A(n14298), .ZN(n11661) );
  INV_X1 U14038 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n11657) );
  INV_X1 U14039 ( .A(n11655), .ZN(n14260) );
  OAI22_X1 U14040 ( .A1(n14963), .A2(n11657), .B1(n14260), .B2(n11656), .ZN(
        n11660) );
  XNOR2_X1 U14041 ( .A(n11658), .B(n12121), .ZN(n14299) );
  NOR2_X1 U14042 ( .A1(n14299), .A2(n12621), .ZN(n11659) );
  AOI211_X1 U14043 ( .C1(n12618), .C2(n11661), .A(n11660), .B(n11659), .ZN(
        n11662) );
  OAI21_X1 U14044 ( .B1(n14965), .B2(n14297), .A(n11662), .ZN(P3_U3219) );
  AOI22_X1 U14045 ( .A1(n11663), .A2(n12865), .B1(n12841), .B2(n12884), .ZN(
        n11671) );
  INV_X1 U14046 ( .A(n11664), .ZN(n11670) );
  INV_X1 U14047 ( .A(n11724), .ZN(n11667) );
  NAND2_X1 U14048 ( .A1(n13152), .A2(n12885), .ZN(n11665) );
  OAI21_X1 U14049 ( .B1(n11826), .B2(n13069), .A(n11665), .ZN(n11720) );
  AOI22_X1 U14050 ( .A1(n12798), .A2(n11720), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11666) );
  OAI21_X1 U14051 ( .B1(n11667), .B2(n12856), .A(n11666), .ZN(n11668) );
  AOI21_X1 U14052 ( .B1(n13269), .B2(n12871), .A(n11668), .ZN(n11669) );
  OAI21_X1 U14053 ( .B1(n11671), .B2(n11670), .A(n11669), .ZN(P2_U3213) );
  INV_X1 U14054 ( .A(n11673), .ZN(n11674) );
  XNOR2_X1 U14055 ( .A(n14298), .B(n11980), .ZN(n11676) );
  XNOR2_X1 U14056 ( .A(n11676), .B(n11678), .ZN(n14252) );
  XNOR2_X1 U14057 ( .A(n12745), .B(n11980), .ZN(n11775) );
  XNOR2_X1 U14058 ( .A(n11775), .B(n11778), .ZN(n11776) );
  XNOR2_X1 U14059 ( .A(n11777), .B(n11776), .ZN(n11684) );
  INV_X1 U14060 ( .A(n12617), .ZN(n11681) );
  INV_X1 U14061 ( .A(n12318), .ZN(n11677) );
  OAI22_X1 U14062 ( .A1(n11678), .A2(n12055), .B1(n11677), .B2(n12057), .ZN(
        n12615) );
  NOR2_X1 U14063 ( .A1(n11679), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14264) );
  AOI21_X1 U14064 ( .B1(n12615), .B2(n14884), .A(n14264), .ZN(n11680) );
  OAI21_X1 U14065 ( .B1(n11681), .B2(n14893), .A(n11680), .ZN(n11682) );
  AOI21_X1 U14066 ( .B1(n12745), .B2(n12062), .A(n11682), .ZN(n11683) );
  OAI21_X1 U14067 ( .B1(n11684), .B2(n14881), .A(n11683), .ZN(P3_U3181) );
  NAND2_X1 U14068 ( .A1(n11686), .A2(n11685), .ZN(n11687) );
  NAND2_X1 U14069 ( .A1(n11693), .A2(n13465), .ZN(n11690) );
  NAND2_X1 U14070 ( .A1(n13590), .A2(n13462), .ZN(n11689) );
  NAND2_X1 U14071 ( .A1(n11690), .A2(n11689), .ZN(n11691) );
  XNOR2_X1 U14072 ( .A(n11691), .B(n13463), .ZN(n11805) );
  AND2_X1 U14073 ( .A1(n13590), .A2(n10598), .ZN(n11692) );
  AOI21_X1 U14074 ( .B1(n11693), .B2(n13462), .A(n11692), .ZN(n11803) );
  XNOR2_X1 U14075 ( .A(n11805), .B(n11803), .ZN(n11694) );
  OAI211_X1 U14076 ( .C1(n11695), .C2(n11694), .A(n11807), .B(n13570), .ZN(
        n11701) );
  OAI21_X1 U14077 ( .B1(n14325), .B2(n14327), .A(n11696), .ZN(n11699) );
  NOR2_X1 U14078 ( .A1(n14339), .A2(n11697), .ZN(n11698) );
  AOI211_X1 U14079 ( .C1(n13577), .C2(n14506), .A(n11699), .B(n11698), .ZN(
        n11700) );
  OAI211_X1 U14080 ( .C1(n11702), .C2(n13580), .A(n11701), .B(n11700), .ZN(
        P1_U3224) );
  XNOR2_X1 U14081 ( .A(n11703), .B(n11708), .ZN(n11734) );
  AOI21_X1 U14082 ( .B1(n11730), .B2(n11704), .A(n13190), .ZN(n11705) );
  NAND2_X1 U14083 ( .A1(n11705), .A2(n11723), .ZN(n11731) );
  AOI22_X1 U14084 ( .A1(n13187), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11898), 
        .B2(n13175), .ZN(n11707) );
  NAND2_X1 U14085 ( .A1(n11730), .A2(n13143), .ZN(n11706) );
  OAI211_X1 U14086 ( .C1(n11731), .C2(n13140), .A(n11707), .B(n11706), .ZN(
        n11714) );
  OAI21_X1 U14087 ( .B1(n7383), .B2(n7843), .A(n11709), .ZN(n11712) );
  NAND2_X1 U14088 ( .A1(n13152), .A2(n12886), .ZN(n11710) );
  OAI21_X1 U14089 ( .B1(n11711), .B2(n13069), .A(n11710), .ZN(n11897) );
  AOI21_X1 U14090 ( .B1(n11712), .B2(n13169), .A(n11897), .ZN(n11732) );
  NOR2_X1 U14091 ( .A1(n11732), .A2(n13187), .ZN(n11713) );
  AOI211_X1 U14092 ( .C1(n11734), .C2(n13122), .A(n11714), .B(n11713), .ZN(
        n11715) );
  INV_X1 U14093 ( .A(n11715), .ZN(P2_U3251) );
  XNOR2_X1 U14094 ( .A(n11716), .B(n11718), .ZN(n13272) );
  AOI21_X1 U14095 ( .B1(n11719), .B2(n11718), .A(n13064), .ZN(n11721) );
  AOI21_X1 U14096 ( .B1(n11717), .B2(n11721), .A(n11720), .ZN(n13271) );
  INV_X1 U14097 ( .A(n11751), .ZN(n11722) );
  AOI211_X1 U14098 ( .C1(n13269), .C2(n11723), .A(n13190), .B(n11722), .ZN(
        n13268) );
  AOI22_X1 U14099 ( .A1(n13268), .A2(n11725), .B1(n13175), .B2(n11724), .ZN(
        n11726) );
  AOI21_X1 U14100 ( .B1(n13271), .B2(n11726), .A(n13187), .ZN(n11727) );
  INV_X1 U14101 ( .A(n11727), .ZN(n11729) );
  AOI22_X1 U14102 ( .A1(n13269), .A2(n13143), .B1(n13187), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n11728) );
  OAI211_X1 U14103 ( .C1(n13182), .C2(n13272), .A(n11729), .B(n11728), .ZN(
        P2_U3250) );
  INV_X1 U14104 ( .A(n11730), .ZN(n11901) );
  OAI211_X1 U14105 ( .C1(n11901), .C2(n14852), .A(n11732), .B(n11731), .ZN(
        n11733) );
  AOI21_X1 U14106 ( .B1(n11734), .B2(n8001), .A(n11733), .ZN(n11737) );
  NAND2_X1 U14107 ( .A1(n14873), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n11735) );
  OAI21_X1 U14108 ( .B1(n11737), .B2(n14873), .A(n11735), .ZN(P2_U3513) );
  NAND2_X1 U14109 ( .A1(n14856), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n11736) );
  OAI21_X1 U14110 ( .B1(n11737), .B2(n14856), .A(n11736), .ZN(P2_U3472) );
  NAND2_X1 U14111 ( .A1(n11738), .A2(n11741), .ZN(n11739) );
  NAND2_X1 U14112 ( .A1(n11740), .A2(n11739), .ZN(n13265) );
  INV_X1 U14113 ( .A(n11741), .ZN(n11743) );
  NAND3_X1 U14114 ( .A1(n11717), .A2(n11743), .A3(n11742), .ZN(n11744) );
  NAND3_X1 U14115 ( .A1(n11745), .A2(n13169), .A3(n11744), .ZN(n11748) );
  NAND2_X1 U14116 ( .A1(n13153), .A2(n13151), .ZN(n11747) );
  NAND2_X1 U14117 ( .A1(n13152), .A2(n12884), .ZN(n11746) );
  AND2_X1 U14118 ( .A1(n11747), .A2(n11746), .ZN(n11838) );
  NAND2_X1 U14119 ( .A1(n11748), .A2(n11838), .ZN(n13267) );
  NAND2_X1 U14120 ( .A1(n13267), .A2(n13135), .ZN(n11757) );
  INV_X1 U14121 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11750) );
  INV_X1 U14122 ( .A(n11840), .ZN(n11749) );
  OAI22_X1 U14123 ( .A1(n13135), .A2(n11750), .B1(n11749), .B2(n13133), .ZN(
        n11755) );
  NAND2_X1 U14124 ( .A1(n11751), .A2(n13262), .ZN(n11752) );
  NAND2_X1 U14125 ( .A1(n11752), .A2(n13136), .ZN(n11753) );
  OR2_X1 U14126 ( .A1(n11753), .A2(n13171), .ZN(n13264) );
  NOR2_X1 U14127 ( .A1(n13264), .A2(n13140), .ZN(n11754) );
  AOI211_X1 U14128 ( .C1(n13143), .C2(n13262), .A(n11755), .B(n11754), .ZN(
        n11756) );
  OAI211_X1 U14129 ( .C1(n13182), .C2(n13265), .A(n11757), .B(n11756), .ZN(
        P2_U3249) );
  INV_X1 U14130 ( .A(n13330), .ZN(n13588) );
  INV_X1 U14131 ( .A(n11790), .ZN(n11760) );
  AOI21_X1 U14132 ( .B1(n11764), .B2(n11761), .A(n11760), .ZN(n14365) );
  NAND2_X1 U14133 ( .A1(n11763), .A2(n11762), .ZN(n11765) );
  OAI211_X1 U14134 ( .C1(n11765), .C2(n11764), .A(n11786), .B(n14519), .ZN(
        n14363) );
  INV_X1 U14135 ( .A(n14363), .ZN(n11768) );
  OR2_X1 U14136 ( .A1(n13330), .A2(n14523), .ZN(n11767) );
  NAND2_X1 U14137 ( .A1(n13586), .A2(n14507), .ZN(n11766) );
  NAND2_X1 U14138 ( .A1(n11767), .A2(n11766), .ZN(n14361) );
  OAI21_X1 U14139 ( .B1(n11768), .B2(n14361), .A(n14543), .ZN(n11774) );
  AOI211_X1 U14140 ( .C1(n14362), .C2(n11769), .A(n14526), .B(n11791), .ZN(
        n14360) );
  INV_X1 U14141 ( .A(n14362), .ZN(n13581) );
  NOR2_X1 U14142 ( .A1(n13581), .A2(n13958), .ZN(n11772) );
  OAI22_X1 U14143 ( .A1(n14543), .A2(n11770), .B1(n13574), .B2(n13952), .ZN(
        n11771) );
  AOI211_X1 U14144 ( .C1(n14360), .C2(n14511), .A(n11772), .B(n11771), .ZN(
        n11773) );
  OAI211_X1 U14145 ( .C1(n14365), .C2(n13963), .A(n11774), .B(n11773), .ZN(
        P1_U3278) );
  XNOR2_X1 U14146 ( .A(n12738), .B(n11980), .ZN(n11920) );
  XNOR2_X1 U14147 ( .A(n11920), .B(n12318), .ZN(n11922) );
  XNOR2_X1 U14148 ( .A(n11923), .B(n11922), .ZN(n11784) );
  INV_X1 U14149 ( .A(n12604), .ZN(n11781) );
  OR2_X1 U14150 ( .A1(n11778), .A2(n12055), .ZN(n11779) );
  OAI21_X1 U14151 ( .B1(n12056), .B2(n12057), .A(n11779), .ZN(n12607) );
  NAND2_X1 U14152 ( .A1(n12607), .A2(n14884), .ZN(n11780) );
  NAND2_X1 U14153 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n14287)
         );
  OAI211_X1 U14154 ( .C1(n11781), .C2(n14893), .A(n11780), .B(n14287), .ZN(
        n11782) );
  AOI21_X1 U14155 ( .B1(n12738), .B2(n12062), .A(n11782), .ZN(n11783) );
  OAI21_X1 U14156 ( .B1(n11784), .B2(n14881), .A(n11783), .ZN(P3_U3166) );
  XNOR2_X1 U14157 ( .A(n11849), .B(n11868), .ZN(n11788) );
  AOI22_X1 U14158 ( .A1(n13587), .A2(n13929), .B1(n14507), .B2(n13928), .ZN(
        n13509) );
  INV_X1 U14159 ( .A(n13509), .ZN(n11787) );
  AOI21_X1 U14160 ( .B1(n11788), .B2(n14519), .A(n11787), .ZN(n14356) );
  OR2_X1 U14161 ( .A1(n14362), .A2(n13587), .ZN(n11789) );
  XNOR2_X1 U14162 ( .A(n11869), .B(n11868), .ZN(n14359) );
  NAND2_X1 U14163 ( .A1(n11791), .A2(n14355), .ZN(n13956) );
  OAI211_X1 U14164 ( .C1(n11791), .C2(n14355), .A(n13956), .B(n14508), .ZN(
        n14354) );
  AOI22_X1 U14165 ( .A1(n14545), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n13507), 
        .B2(n14542), .ZN(n11793) );
  NAND2_X1 U14166 ( .A1(n13511), .A2(n14501), .ZN(n11792) );
  OAI211_X1 U14167 ( .C1(n14354), .C2(n13899), .A(n11793), .B(n11792), .ZN(
        n11794) );
  AOI21_X1 U14168 ( .B1(n14359), .B2(n14512), .A(n11794), .ZN(n11795) );
  OAI21_X1 U14169 ( .B1(n14356), .B2(n14545), .A(n11795), .ZN(P1_U3277) );
  INV_X1 U14170 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n11798) );
  NOR2_X1 U14171 ( .A1(n11797), .A2(n11796), .ZN(n11800) );
  MUX2_X1 U14172 ( .A(n11798), .B(n11800), .S(n14589), .Z(n11799) );
  OAI21_X1 U14173 ( .B1(n11802), .B2(n14077), .A(n11799), .ZN(P1_U3501) );
  MUX2_X1 U14174 ( .A(n13700), .B(n11800), .S(n14597), .Z(n11801) );
  OAI21_X1 U14175 ( .B1(n11802), .B2(n14032), .A(n11801), .ZN(P1_U3542) );
  INV_X1 U14176 ( .A(n11803), .ZN(n11804) );
  NAND2_X1 U14177 ( .A1(n11805), .A2(n11804), .ZN(n11806) );
  NAND2_X1 U14178 ( .A1(n14241), .A2(n13465), .ZN(n11809) );
  NAND2_X1 U14179 ( .A1(n13589), .A2(n13462), .ZN(n11808) );
  NAND2_X1 U14180 ( .A1(n11809), .A2(n11808), .ZN(n11810) );
  XNOR2_X1 U14181 ( .A(n11810), .B(n13463), .ZN(n13324) );
  AND2_X1 U14182 ( .A1(n13589), .A2(n10598), .ZN(n11811) );
  AOI21_X1 U14183 ( .B1(n14241), .B2(n6449), .A(n11811), .ZN(n13322) );
  XNOR2_X1 U14184 ( .A(n13324), .B(n13322), .ZN(n11812) );
  OAI211_X1 U14185 ( .C1(n11813), .C2(n11812), .A(n13326), .B(n13570), .ZN(
        n11819) );
  OR2_X1 U14186 ( .A1(n13330), .A2(n14533), .ZN(n11815) );
  NAND2_X1 U14187 ( .A1(n13590), .A2(n13929), .ZN(n11814) );
  NAND2_X1 U14188 ( .A1(n11815), .A2(n11814), .ZN(n14237) );
  NAND2_X1 U14189 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14419)
         );
  INV_X1 U14190 ( .A(n14419), .ZN(n11817) );
  NOR2_X1 U14191 ( .A1(n14339), .A2(n14239), .ZN(n11816) );
  AOI211_X1 U14192 ( .C1(n13534), .C2(n14237), .A(n11817), .B(n11816), .ZN(
        n11818) );
  OAI211_X1 U14193 ( .C1(n14369), .C2(n13580), .A(n11819), .B(n11818), .ZN(
        P1_U3234) );
  INV_X1 U14194 ( .A(n13176), .ZN(n11823) );
  NAND2_X1 U14195 ( .A1(n13153), .A2(n12882), .ZN(n11821) );
  NAND2_X1 U14196 ( .A1(n13152), .A2(n12883), .ZN(n11820) );
  NAND2_X1 U14197 ( .A1(n11821), .A2(n11820), .ZN(n13168) );
  AOI22_X1 U14198 ( .A1(n12798), .A2(n13168), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11822) );
  OAI21_X1 U14199 ( .B1(n11823), .B2(n12856), .A(n11822), .ZN(n11824) );
  AOI21_X1 U14200 ( .B1(n13258), .B2(n12871), .A(n11824), .ZN(n11831) );
  INV_X1 U14201 ( .A(n11825), .ZN(n11829) );
  OAI22_X1 U14202 ( .A1(n11827), .A2(n12858), .B1(n11826), .B2(n12872), .ZN(
        n11828) );
  NAND3_X1 U14203 ( .A1(n11833), .A2(n11829), .A3(n11828), .ZN(n11830) );
  OAI211_X1 U14204 ( .C1(n11832), .C2(n12858), .A(n11831), .B(n11830), .ZN(
        P2_U3200) );
  INV_X1 U14205 ( .A(n11833), .ZN(n11834) );
  AOI21_X1 U14206 ( .B1(n11836), .B2(n11835), .A(n11834), .ZN(n11843) );
  OAI22_X1 U14207 ( .A1(n12828), .A2(n11838), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11837), .ZN(n11839) );
  AOI21_X1 U14208 ( .B1(n11840), .B2(n12867), .A(n11839), .ZN(n11842) );
  NAND2_X1 U14209 ( .A1(n13262), .A2(n12871), .ZN(n11841) );
  OAI211_X1 U14210 ( .C1(n11843), .C2(n12858), .A(n11842), .B(n11841), .ZN(
        P2_U3198) );
  INV_X1 U14211 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n11912) );
  OAI222_X1 U14212 ( .A1(n11844), .A2(P1_U3086), .B1(n14083), .B2(n13303), 
        .C1(n11912), .C2(n14085), .ZN(P1_U3325) );
  INV_X1 U14213 ( .A(n11845), .ZN(n13312) );
  OAI222_X1 U14214 ( .A1(n14085), .A2(n11846), .B1(n14088), .B2(n13312), .C1(
        n8684), .C2(P1_U3086), .ZN(P1_U3328) );
  INV_X1 U14215 ( .A(n11847), .ZN(n11848) );
  INV_X1 U14216 ( .A(n13586), .ZN(n13947) );
  NAND2_X1 U14217 ( .A1(n13511), .A2(n13947), .ZN(n11851) );
  INV_X1 U14218 ( .A(n13943), .ZN(n13945) );
  INV_X1 U14219 ( .A(n13928), .ZN(n11852) );
  OR2_X1 U14220 ( .A1(n14034), .A2(n11852), .ZN(n11853) );
  NAND2_X1 U14221 ( .A1(n13950), .A2(n11853), .ZN(n13927) );
  OR2_X1 U14222 ( .A1(n13936), .A2(n13948), .ZN(n11854) );
  INV_X1 U14223 ( .A(n13888), .ZN(n13890) );
  NAND2_X1 U14224 ( .A1(n14019), .A2(n13913), .ZN(n13871) );
  INV_X1 U14225 ( .A(n13585), .ZN(n11856) );
  OR2_X1 U14226 ( .A1(n13879), .A2(n11856), .ZN(n11857) );
  NAND2_X1 U14227 ( .A1(n13863), .A2(n15190), .ZN(n11859) );
  NAND2_X1 U14228 ( .A1(n13836), .A2(n13837), .ZN(n11863) );
  NAND2_X1 U14229 ( .A1(n14001), .A2(n11861), .ZN(n11862) );
  OR2_X1 U14230 ( .A1(n13827), .A2(n13500), .ZN(n11864) );
  INV_X1 U14231 ( .A(n13583), .ZN(n13501) );
  NAND2_X1 U14232 ( .A1(n13988), .A2(n13501), .ZN(n11866) );
  NOR2_X1 U14233 ( .A1(n13750), .A2(n14548), .ZN(n11885) );
  NAND2_X1 U14234 ( .A1(n13750), .A2(n14519), .ZN(n11883) );
  NAND2_X1 U14235 ( .A1(n11869), .A2(n11868), .ZN(n11871) );
  OR2_X1 U14236 ( .A1(n13511), .A2(n13586), .ZN(n11870) );
  INV_X1 U14237 ( .A(n13553), .ZN(n13930) );
  OR2_X1 U14238 ( .A1(n13917), .A2(n13930), .ZN(n11874) );
  OR2_X1 U14239 ( .A1(n13863), .A2(n13487), .ZN(n11876) );
  NAND2_X1 U14240 ( .A1(n14001), .A2(n13856), .ZN(n11877) );
  INV_X1 U14241 ( .A(n11878), .ZN(n13821) );
  OR2_X1 U14242 ( .A1(n13827), .A2(n13584), .ZN(n11879) );
  NAND2_X1 U14243 ( .A1(n13807), .A2(n13819), .ZN(n11880) );
  NAND2_X1 U14244 ( .A1(n13988), .A2(n13583), .ZN(n11881) );
  NAND2_X1 U14245 ( .A1(n11886), .A2(n14588), .ZN(n11882) );
  NAND2_X1 U14246 ( .A1(n11883), .A2(n11882), .ZN(n11884) );
  MUX2_X1 U14247 ( .A(n11885), .B(n11884), .S(n13749), .Z(n11889) );
  AOI22_X1 U14248 ( .A1(n13759), .A2(n14507), .B1(n13929), .B2(n13583), .ZN(
        n11887) );
  INV_X1 U14249 ( .A(n14001), .ZN(n13845) );
  OAI211_X1 U14250 ( .C1(n14052), .C2(n13794), .A(n14508), .B(n13774), .ZN(
        n13984) );
  AOI22_X1 U14251 ( .A1(n13425), .A2(n14542), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n14545), .ZN(n11890) );
  OAI21_X1 U14252 ( .B1(n14052), .B2(n13958), .A(n11890), .ZN(n11891) );
  AOI21_X1 U14253 ( .B1(n6711), .B2(n14511), .A(n11891), .ZN(n11892) );
  OAI21_X1 U14254 ( .B1(n13985), .B2(n14545), .A(n11892), .ZN(P1_U3266) );
  NAND3_X1 U14255 ( .A1(n11893), .A2(n12841), .A3(n12886), .ZN(n11894) );
  OAI21_X1 U14256 ( .B1(n11895), .B2(n12858), .A(n11894), .ZN(n11904) );
  INV_X1 U14257 ( .A(n11896), .ZN(n11903) );
  AOI22_X1 U14258 ( .A1(n12798), .A2(n11897), .B1(P2_REG3_REG_14__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11900) );
  NAND2_X1 U14259 ( .A1(n12867), .A2(n11898), .ZN(n11899) );
  OAI211_X1 U14260 ( .C1(n11901), .C2(n12829), .A(n11900), .B(n11899), .ZN(
        n11902) );
  AOI21_X1 U14261 ( .B1(n11904), .B2(n11903), .A(n11902), .ZN(n11905) );
  OAI21_X1 U14262 ( .B1(n11906), .B2(n12858), .A(n11905), .ZN(P2_U3187) );
  INV_X1 U14263 ( .A(n11908), .ZN(n11910) );
  NAND2_X1 U14264 ( .A1(n14086), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11909) );
  INV_X1 U14265 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13301) );
  NAND2_X1 U14266 ( .A1(n13301), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12076) );
  NAND2_X1 U14267 ( .A1(n11912), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n11913) );
  NAND2_X1 U14268 ( .A1(n12076), .A2(n11913), .ZN(n12077) );
  XNOR2_X1 U14269 ( .A(n12078), .B(n12077), .ZN(n12084) );
  INV_X1 U14270 ( .A(n12084), .ZN(n11914) );
  INV_X1 U14271 ( .A(SI_30_), .ZN(n12085) );
  INV_X1 U14272 ( .A(n13307), .ZN(n11916) );
  OAI222_X1 U14273 ( .A1(n14085), .A2(n11917), .B1(n14083), .B2(n11916), .C1(
        P1_U3086), .C2(n8685), .ZN(P1_U3327) );
  XNOR2_X1 U14274 ( .A(n12627), .B(n11931), .ZN(n11919) );
  INV_X1 U14275 ( .A(n11918), .ZN(n12308) );
  NOR2_X1 U14276 ( .A1(n11919), .A2(n12308), .ZN(n11977) );
  AOI21_X1 U14277 ( .B1(n11919), .B2(n12308), .A(n11977), .ZN(n11953) );
  INV_X1 U14278 ( .A(n11920), .ZN(n11921) );
  XNOR2_X1 U14279 ( .A(n12600), .B(n11980), .ZN(n11924) );
  XNOR2_X1 U14280 ( .A(n11924), .B(n12056), .ZN(n12018) );
  XNOR2_X1 U14281 ( .A(n12726), .B(n11980), .ZN(n11925) );
  XOR2_X1 U14282 ( .A(n12020), .B(n11925), .Z(n12053) );
  INV_X1 U14283 ( .A(n11925), .ZN(n11926) );
  INV_X1 U14284 ( .A(n12020), .ZN(n12317) );
  XNOR2_X1 U14285 ( .A(n12111), .B(n11980), .ZN(n11927) );
  XNOR2_X1 U14286 ( .A(n11927), .B(n12316), .ZN(n11969) );
  INV_X1 U14287 ( .A(n11927), .ZN(n11928) );
  XNOR2_X1 U14288 ( .A(n12714), .B(n11980), .ZN(n11929) );
  XOR2_X1 U14289 ( .A(n11971), .B(n11929), .Z(n12037) );
  INV_X1 U14290 ( .A(n11929), .ZN(n11930) );
  INV_X1 U14291 ( .A(n11971), .ZN(n12315) );
  XNOR2_X1 U14292 ( .A(n12557), .B(n11931), .ZN(n11932) );
  INV_X1 U14293 ( .A(n12047), .ZN(n12314) );
  NOR2_X1 U14294 ( .A1(n11932), .A2(n12314), .ZN(n11933) );
  AOI21_X1 U14295 ( .B1(n11932), .B2(n12314), .A(n11933), .ZN(n11991) );
  NAND2_X1 U14296 ( .A1(n11990), .A2(n11991), .ZN(n11989) );
  INV_X1 U14297 ( .A(n11933), .ZN(n11934) );
  XNOR2_X1 U14298 ( .A(n12703), .B(n11980), .ZN(n11935) );
  XNOR2_X1 U14299 ( .A(n12255), .B(n11980), .ZN(n11937) );
  INV_X1 U14300 ( .A(n12312), .ZN(n12046) );
  INV_X1 U14301 ( .A(n11940), .ZN(n12028) );
  XNOR2_X1 U14302 ( .A(n12691), .B(n11980), .ZN(n11941) );
  INV_X1 U14303 ( .A(n12311), .ZN(n11963) );
  NAND2_X1 U14304 ( .A1(n11941), .A2(n11963), .ZN(n11944) );
  INV_X1 U14305 ( .A(n11941), .ZN(n11942) );
  NAND2_X1 U14306 ( .A1(n11942), .A2(n12311), .ZN(n11943) );
  NAND2_X1 U14307 ( .A1(n11944), .A2(n11943), .ZN(n12027) );
  INV_X1 U14308 ( .A(n11944), .ZN(n11999) );
  XNOR2_X1 U14309 ( .A(n12516), .B(n11980), .ZN(n11945) );
  NAND2_X1 U14310 ( .A1(n11945), .A2(n12032), .ZN(n11948) );
  INV_X1 U14311 ( .A(n11945), .ZN(n11946) );
  INV_X1 U14312 ( .A(n12032), .ZN(n12310) );
  NAND2_X1 U14313 ( .A1(n11946), .A2(n12310), .ZN(n11947) );
  AND2_X1 U14314 ( .A1(n11948), .A2(n11947), .ZN(n11998) );
  XNOR2_X1 U14315 ( .A(n12680), .B(n11980), .ZN(n11949) );
  NOR2_X1 U14316 ( .A1(n11949), .A2(n12309), .ZN(n11950) );
  AOI21_X1 U14317 ( .B1(n11949), .B2(n12309), .A(n11950), .ZN(n12067) );
  INV_X1 U14318 ( .A(n11950), .ZN(n11951) );
  NAND2_X1 U14319 ( .A1(n12065), .A2(n11951), .ZN(n11952) );
  NAND2_X1 U14320 ( .A1(n11952), .A2(n11953), .ZN(n11979) );
  OAI21_X1 U14321 ( .B1(n11953), .B2(n11952), .A(n11979), .ZN(n11954) );
  NAND2_X1 U14322 ( .A1(n11954), .A2(n14257), .ZN(n11960) );
  OAI22_X1 U14323 ( .A1(n11956), .A2(n12057), .B1(n11955), .B2(n12055), .ZN(
        n12482) );
  AOI22_X1 U14324 ( .A1(n12482), .A2(n14884), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11959) );
  NAND2_X1 U14325 ( .A1(n12627), .A2(n12062), .ZN(n11958) );
  NAND2_X1 U14326 ( .A1(n12073), .A2(n12487), .ZN(n11957) );
  NAND4_X1 U14327 ( .A1(n11960), .A2(n11959), .A3(n11958), .A4(n11957), .ZN(
        P3_U3154) );
  OAI21_X1 U14328 ( .B1(n12046), .B2(n11961), .A(n12029), .ZN(n11962) );
  NAND2_X1 U14329 ( .A1(n11962), .A2(n14257), .ZN(n11968) );
  OAI22_X1 U14330 ( .A1(n11964), .A2(n12055), .B1(n11963), .B2(n12057), .ZN(
        n12533) );
  INV_X1 U14331 ( .A(n12533), .ZN(n11965) );
  OAI22_X1 U14332 ( .A1(n11965), .A2(n12071), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15082), .ZN(n11966) );
  AOI21_X1 U14333 ( .B1(n12536), .B2(n12073), .A(n11966), .ZN(n11967) );
  OAI211_X1 U14334 ( .C1(n12255), .C2(n14889), .A(n11968), .B(n11967), .ZN(
        P3_U3156) );
  XNOR2_X1 U14335 ( .A(n11970), .B(n11969), .ZN(n11976) );
  INV_X1 U14336 ( .A(n12575), .ZN(n11973) );
  OAI22_X1 U14337 ( .A1(n11971), .A2(n12057), .B1(n12020), .B2(n12055), .ZN(
        n12572) );
  NAND2_X1 U14338 ( .A1(n12572), .A2(n14884), .ZN(n11972) );
  NAND2_X1 U14339 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12466)
         );
  OAI211_X1 U14340 ( .C1(n14893), .C2(n11973), .A(n11972), .B(n12466), .ZN(
        n11974) );
  AOI21_X1 U14341 ( .B1(n12720), .B2(n12062), .A(n11974), .ZN(n11975) );
  OAI21_X1 U14342 ( .B1(n11976), .B2(n14881), .A(n11975), .ZN(P3_U3159) );
  INV_X1 U14343 ( .A(n11977), .ZN(n11978) );
  NAND2_X1 U14344 ( .A1(n11979), .A2(n11978), .ZN(n11982) );
  XNOR2_X1 U14345 ( .A(n12108), .B(n11980), .ZN(n11981) );
  XNOR2_X1 U14346 ( .A(n11982), .B(n11981), .ZN(n11988) );
  INV_X1 U14347 ( .A(n12476), .ZN(n11985) );
  AOI22_X1 U14348 ( .A1(n11983), .A2(n14884), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11984) );
  OAI21_X1 U14349 ( .B1(n11985), .B2(n14893), .A(n11984), .ZN(n11986) );
  AOI21_X1 U14350 ( .B1(n12477), .B2(n12062), .A(n11986), .ZN(n11987) );
  OAI21_X1 U14351 ( .B1(n11988), .B2(n14881), .A(n11987), .ZN(P3_U3160) );
  OAI21_X1 U14352 ( .B1(n11991), .B2(n11990), .A(n11989), .ZN(n11992) );
  NAND2_X1 U14353 ( .A1(n11992), .A2(n14257), .ZN(n11996) );
  AOI22_X1 U14354 ( .A1(n12313), .A2(n12069), .B1(n12300), .B2(n12315), .ZN(
        n12552) );
  INV_X1 U14355 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n11993) );
  OAI22_X1 U14356 ( .A1(n12552), .A2(n12071), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11993), .ZN(n11994) );
  AOI21_X1 U14357 ( .B1(n12556), .B2(n12073), .A(n11994), .ZN(n11995) );
  OAI211_X1 U14358 ( .C1(n12708), .C2(n14889), .A(n11996), .B(n11995), .ZN(
        P3_U3163) );
  INV_X1 U14359 ( .A(n11997), .ZN(n12001) );
  NOR3_X1 U14360 ( .A1(n12031), .A2(n11999), .A3(n11998), .ZN(n12000) );
  OAI21_X1 U14361 ( .B1(n12001), .B2(n12000), .A(n14257), .ZN(n12005) );
  AOI22_X1 U14362 ( .A1(n12309), .A2(n12069), .B1(n12300), .B2(n12311), .ZN(
        n12511) );
  INV_X1 U14363 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n12002) );
  OAI22_X1 U14364 ( .A1(n12511), .A2(n12071), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12002), .ZN(n12003) );
  AOI21_X1 U14365 ( .B1(n12515), .B2(n12073), .A(n12003), .ZN(n12004) );
  OAI211_X1 U14366 ( .C1(n12685), .C2(n14889), .A(n12005), .B(n12004), .ZN(
        P3_U3165) );
  OAI21_X1 U14367 ( .B1(n12008), .B2(n12007), .A(n12006), .ZN(n12009) );
  NAND2_X1 U14368 ( .A1(n12009), .A2(n14257), .ZN(n12017) );
  AOI21_X1 U14369 ( .B1(n12062), .B2(n12011), .A(n12010), .ZN(n12016) );
  NAND2_X1 U14370 ( .A1(n12073), .A2(n12012), .ZN(n12015) );
  NAND2_X1 U14371 ( .A1(n12013), .A2(n14884), .ZN(n12014) );
  NAND4_X1 U14372 ( .A1(n12017), .A2(n12016), .A3(n12015), .A4(n12014), .ZN(
        P3_U3167) );
  XNOR2_X1 U14373 ( .A(n12019), .B(n12018), .ZN(n12026) );
  OR2_X1 U14374 ( .A1(n12020), .A2(n12057), .ZN(n12022) );
  NAND2_X1 U14375 ( .A1(n12318), .A2(n12300), .ZN(n12021) );
  AND2_X1 U14376 ( .A1(n12022), .A2(n12021), .ZN(n12596) );
  NAND2_X1 U14377 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12406)
         );
  NAND2_X1 U14378 ( .A1(n12073), .A2(n12599), .ZN(n12023) );
  OAI211_X1 U14379 ( .C1(n12596), .C2(n12071), .A(n12406), .B(n12023), .ZN(
        n12024) );
  AOI21_X1 U14380 ( .B1(n12600), .B2(n12062), .A(n12024), .ZN(n12025) );
  OAI21_X1 U14381 ( .B1(n12026), .B2(n14881), .A(n12025), .ZN(P3_U3168) );
  AND3_X1 U14382 ( .A1(n12029), .A2(n12028), .A3(n12027), .ZN(n12030) );
  OAI21_X1 U14383 ( .B1(n12031), .B2(n12030), .A(n14257), .ZN(n12036) );
  OAI22_X1 U14384 ( .A1(n12046), .A2(n12055), .B1(n12032), .B2(n12057), .ZN(
        n12522) );
  AOI22_X1 U14385 ( .A1(n12522), .A2(n14884), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12035) );
  NAND2_X1 U14386 ( .A1(n12691), .A2(n12062), .ZN(n12034) );
  NAND2_X1 U14387 ( .A1(n12073), .A2(n12525), .ZN(n12033) );
  NAND4_X1 U14388 ( .A1(n12036), .A2(n12035), .A3(n12034), .A4(n12033), .ZN(
        P3_U3169) );
  XNOR2_X1 U14389 ( .A(n12038), .B(n12037), .ZN(n12043) );
  INV_X1 U14390 ( .A(n12567), .ZN(n12040) );
  OAI22_X1 U14391 ( .A1(n12047), .A2(n12057), .B1(n12058), .B2(n12055), .ZN(
        n12564) );
  AOI22_X1 U14392 ( .A1(n12564), .A2(n14884), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12039) );
  OAI21_X1 U14393 ( .B1(n12040), .B2(n14893), .A(n12039), .ZN(n12041) );
  AOI21_X1 U14394 ( .B1(n12714), .B2(n12062), .A(n12041), .ZN(n12042) );
  OAI21_X1 U14395 ( .B1(n12043), .B2(n14881), .A(n12042), .ZN(P3_U3173) );
  AOI21_X1 U14396 ( .B1(n12313), .B2(n12045), .A(n12044), .ZN(n12052) );
  INV_X1 U14397 ( .A(n12545), .ZN(n12049) );
  OAI22_X1 U14398 ( .A1(n12047), .A2(n12055), .B1(n12046), .B2(n12057), .ZN(
        n12542) );
  AOI22_X1 U14399 ( .A1(n12542), .A2(n14884), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12048) );
  OAI21_X1 U14400 ( .B1(n12049), .B2(n14893), .A(n12048), .ZN(n12050) );
  AOI21_X1 U14401 ( .B1(n12703), .B2(n12062), .A(n12050), .ZN(n12051) );
  OAI21_X1 U14402 ( .B1(n12052), .B2(n14881), .A(n12051), .ZN(P3_U3175) );
  XNOR2_X1 U14403 ( .A(n12054), .B(n12053), .ZN(n12064) );
  INV_X1 U14404 ( .A(n12587), .ZN(n12060) );
  OAI22_X1 U14405 ( .A1(n12058), .A2(n12057), .B1(n12056), .B2(n12055), .ZN(
        n12584) );
  NAND2_X1 U14406 ( .A1(n12584), .A2(n14884), .ZN(n12059) );
  NAND2_X1 U14407 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12442)
         );
  OAI211_X1 U14408 ( .C1(n12060), .C2(n14893), .A(n12059), .B(n12442), .ZN(
        n12061) );
  AOI21_X1 U14409 ( .B1(n12726), .B2(n12062), .A(n12061), .ZN(n12063) );
  OAI21_X1 U14410 ( .B1(n12064), .B2(n14881), .A(n12063), .ZN(P3_U3178) );
  OAI21_X1 U14411 ( .B1(n12067), .B2(n12066), .A(n12065), .ZN(n12068) );
  NAND2_X1 U14412 ( .A1(n12068), .A2(n14257), .ZN(n12075) );
  AOI22_X1 U14413 ( .A1(n12300), .A2(n12310), .B1(n12308), .B2(n12069), .ZN(
        n12498) );
  INV_X1 U14414 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n12070) );
  OAI22_X1 U14415 ( .A1(n12498), .A2(n12071), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12070), .ZN(n12072) );
  AOI21_X1 U14416 ( .B1(n12502), .B2(n12073), .A(n12072), .ZN(n12074) );
  OAI211_X1 U14417 ( .C1(n12680), .C2(n14889), .A(n12075), .B(n12074), .ZN(
        P3_U3180) );
  OAI21_X1 U14418 ( .B1(n12078), .B2(n12077), .A(n12076), .ZN(n12080) );
  XNOR2_X1 U14419 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12079) );
  XNOR2_X1 U14420 ( .A(n12080), .B(n12079), .ZN(n12757) );
  NAND2_X1 U14421 ( .A1(n12757), .A2(n12083), .ZN(n12082) );
  INV_X1 U14422 ( .A(SI_31_), .ZN(n12754) );
  OR2_X1 U14423 ( .A1(n12086), .A2(n12754), .ZN(n12081) );
  NAND2_X1 U14424 ( .A1(n12084), .A2(n12083), .ZN(n12088) );
  OR2_X1 U14425 ( .A1(n12086), .A2(n12085), .ZN(n12087) );
  INV_X1 U14426 ( .A(n12669), .ZN(n12626) );
  NAND2_X1 U14427 ( .A1(n12626), .A2(n12306), .ZN(n12106) );
  NAND2_X1 U14428 ( .A1(n12089), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12094) );
  NAND2_X1 U14429 ( .A1(n6443), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12093) );
  NAND2_X1 U14430 ( .A1(n12091), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12092) );
  NAND2_X1 U14431 ( .A1(n12106), .A2(n6619), .ZN(n12103) );
  INV_X1 U14432 ( .A(n12306), .ZN(n12097) );
  NAND2_X1 U14433 ( .A1(n12669), .A2(n12097), .ZN(n12098) );
  NAND2_X1 U14434 ( .A1(n12284), .A2(n12098), .ZN(n12131) );
  INV_X1 U14435 ( .A(n12099), .ZN(n12100) );
  OAI21_X1 U14436 ( .B1(n12626), .B2(n6619), .A(n12283), .ZN(n12101) );
  AOI21_X1 U14437 ( .B1(n12665), .B2(n12103), .A(n12102), .ZN(n12104) );
  XNOR2_X1 U14438 ( .A(n12104), .B(n12459), .ZN(n12296) );
  INV_X1 U14439 ( .A(n12105), .ZN(n12295) );
  INV_X1 U14440 ( .A(n12269), .ZN(n12109) );
  INV_X1 U14441 ( .A(n12110), .ZN(n12133) );
  OR2_X1 U14442 ( .A1(n12134), .A2(n12133), .ZN(n12250) );
  XNOR2_X1 U14443 ( .A(n12111), .B(n12316), .ZN(n12571) );
  NOR4_X1 U14444 ( .A1(n7278), .A2(n12113), .A3(n12112), .A4(n10236), .ZN(
        n12114) );
  NAND4_X1 U14445 ( .A1(n12114), .A2(n12171), .A3(n12160), .A4(n12177), .ZN(
        n12117) );
  NOR4_X1 U14446 ( .A1(n12117), .A2(n8933), .A3(n12116), .A4(n12115), .ZN(
        n12120) );
  NAND4_X1 U14447 ( .A1(n12120), .A2(n12119), .A3(n12118), .A4(n6868), .ZN(
        n12123) );
  NOR4_X1 U14448 ( .A1(n12123), .A2(n12614), .A3(n12122), .A4(n12121), .ZN(
        n12124) );
  NAND4_X1 U14449 ( .A1(n12581), .A2(n12591), .A3(n12124), .A4(n12606), .ZN(
        n12125) );
  NOR2_X1 U14450 ( .A1(n12571), .A2(n12125), .ZN(n12126) );
  NAND4_X1 U14451 ( .A1(n12540), .A2(n12551), .A3(n12560), .A4(n12126), .ZN(
        n12127) );
  NOR4_X1 U14452 ( .A1(n12256), .A2(n7265), .A3(n12528), .A4(n12127), .ZN(
        n12128) );
  NAND4_X1 U14453 ( .A1(n12276), .A2(n12497), .A3(n12128), .A4(n6849), .ZN(
        n12129) );
  XNOR2_X1 U14454 ( .A(n12132), .B(n12454), .ZN(n12292) );
  MUX2_X1 U14455 ( .A(n12134), .B(n12133), .S(n12273), .Z(n12254) );
  INV_X1 U14456 ( .A(n12135), .ZN(n12136) );
  AOI21_X1 U14457 ( .B1(n12137), .B2(n12273), .A(n12136), .ZN(n12198) );
  OAI21_X1 U14458 ( .B1(n12138), .B2(n12140), .A(n12273), .ZN(n12143) );
  NAND3_X1 U14459 ( .A1(n12145), .A2(n12139), .A3(n12302), .ZN(n12142) );
  AOI22_X1 U14460 ( .A1(n12143), .A2(n12142), .B1(n12141), .B2(n12140), .ZN(
        n12144) );
  MUX2_X1 U14461 ( .A(n12277), .B(n12144), .S(n9240), .Z(n12150) );
  OAI21_X1 U14462 ( .B1(n12277), .B2(n12145), .A(n14938), .ZN(n12149) );
  INV_X1 U14463 ( .A(n12146), .ZN(n12147) );
  AOI21_X1 U14464 ( .B1(n12331), .B2(n14943), .A(n12147), .ZN(n12148) );
  OAI22_X1 U14465 ( .A1(n12150), .A2(n12149), .B1(n12148), .B2(n12273), .ZN(
        n12154) );
  AOI21_X1 U14466 ( .B1(n12153), .B2(n12151), .A(n12277), .ZN(n12152) );
  AOI21_X1 U14467 ( .B1(n12154), .B2(n12153), .A(n12152), .ZN(n12162) );
  OAI21_X1 U14468 ( .B1(n12277), .B2(n12146), .A(n12155), .ZN(n12161) );
  NAND2_X1 U14469 ( .A1(n12330), .A2(n12156), .ZN(n12158) );
  MUX2_X1 U14470 ( .A(n12158), .B(n12157), .S(n12273), .Z(n12159) );
  OAI211_X1 U14471 ( .C1(n12162), .C2(n12161), .A(n12160), .B(n12159), .ZN(
        n12163) );
  INV_X1 U14472 ( .A(n12163), .ZN(n12173) );
  NAND2_X1 U14473 ( .A1(n12169), .A2(n12164), .ZN(n12167) );
  NAND2_X1 U14474 ( .A1(n12168), .A2(n12165), .ZN(n12166) );
  MUX2_X1 U14475 ( .A(n12167), .B(n12166), .S(n12277), .Z(n12172) );
  MUX2_X1 U14476 ( .A(n12169), .B(n12168), .S(n12273), .Z(n12170) );
  OAI211_X1 U14477 ( .C1(n12173), .C2(n12172), .A(n12171), .B(n12170), .ZN(
        n12178) );
  MUX2_X1 U14478 ( .A(n12175), .B(n12174), .S(n12277), .Z(n12176) );
  NAND3_X1 U14479 ( .A1(n12178), .A2(n12177), .A3(n12176), .ZN(n12183) );
  MUX2_X1 U14480 ( .A(n12180), .B(n12179), .S(n12273), .Z(n12181) );
  AND3_X1 U14481 ( .A1(n12183), .A2(n12182), .A3(n12181), .ZN(n12185) );
  NOR3_X1 U14482 ( .A1(n12185), .A2(n12190), .A3(n12184), .ZN(n12193) );
  INV_X1 U14483 ( .A(n12193), .ZN(n12197) );
  NAND2_X1 U14484 ( .A1(n6868), .A2(n12186), .ZN(n12195) );
  NAND2_X1 U14485 ( .A1(n12323), .A2(n12187), .ZN(n12188) );
  OAI211_X1 U14486 ( .C1(n12190), .C2(n12189), .A(n12204), .B(n12188), .ZN(
        n12191) );
  AOI21_X1 U14487 ( .B1(n12193), .B2(n12192), .A(n12191), .ZN(n12194) );
  MUX2_X1 U14488 ( .A(n12195), .B(n12194), .S(n12277), .Z(n12196) );
  OAI21_X1 U14489 ( .B1(n12198), .B2(n12197), .A(n12196), .ZN(n12202) );
  AOI21_X1 U14490 ( .B1(n12201), .B2(n12199), .A(n12277), .ZN(n12200) );
  AOI21_X1 U14491 ( .B1(n12202), .B2(n12201), .A(n12200), .ZN(n12209) );
  OAI21_X1 U14492 ( .B1(n12277), .B2(n12204), .A(n12203), .ZN(n12208) );
  MUX2_X1 U14493 ( .A(n12206), .B(n12205), .S(n12273), .Z(n12207) );
  OAI21_X1 U14494 ( .B1(n12209), .B2(n12208), .A(n12207), .ZN(n12214) );
  INV_X1 U14495 ( .A(n12210), .ZN(n12212) );
  MUX2_X1 U14496 ( .A(n12212), .B(n12211), .S(n12273), .Z(n12213) );
  AOI211_X1 U14497 ( .C1(n12214), .C2(n7231), .A(n12213), .B(n12614), .ZN(
        n12222) );
  NAND2_X1 U14498 ( .A1(n12215), .A2(n12318), .ZN(n12223) );
  NAND2_X1 U14499 ( .A1(n12223), .A2(n12216), .ZN(n12220) );
  INV_X1 U14500 ( .A(n12224), .ZN(n12218) );
  NAND2_X1 U14501 ( .A1(n12218), .A2(n12217), .ZN(n12219) );
  MUX2_X1 U14502 ( .A(n12220), .B(n12219), .S(n12277), .Z(n12221) );
  NOR2_X1 U14503 ( .A1(n12222), .A2(n12221), .ZN(n12227) );
  INV_X1 U14504 ( .A(n12223), .ZN(n12225) );
  MUX2_X1 U14505 ( .A(n12225), .B(n12224), .S(n12273), .Z(n12226) );
  OAI211_X1 U14506 ( .C1(n12227), .C2(n12226), .A(n12581), .B(n12591), .ZN(
        n12242) );
  INV_X1 U14507 ( .A(n12231), .ZN(n12230) );
  OAI211_X1 U14508 ( .C1(n12230), .C2(n12229), .A(n12237), .B(n12228), .ZN(
        n12235) );
  INV_X1 U14509 ( .A(n12239), .ZN(n12232) );
  OAI211_X1 U14510 ( .C1(n12233), .C2(n12579), .A(n12232), .B(n12231), .ZN(
        n12234) );
  MUX2_X1 U14511 ( .A(n12235), .B(n12234), .S(n12273), .Z(n12236) );
  INV_X1 U14512 ( .A(n12236), .ZN(n12241) );
  INV_X1 U14513 ( .A(n12237), .ZN(n12238) );
  MUX2_X1 U14514 ( .A(n12239), .B(n12238), .S(n12273), .Z(n12240) );
  AOI21_X1 U14515 ( .B1(n12242), .B2(n12241), .A(n12240), .ZN(n12246) );
  INV_X1 U14516 ( .A(n12560), .ZN(n12562) );
  MUX2_X1 U14517 ( .A(n12244), .B(n12243), .S(n12273), .Z(n12245) );
  OAI21_X1 U14518 ( .B1(n12246), .B2(n12562), .A(n12245), .ZN(n12252) );
  INV_X1 U14519 ( .A(n12247), .ZN(n12248) );
  MUX2_X1 U14520 ( .A(n12249), .B(n12248), .S(n12273), .Z(n12251) );
  AOI211_X1 U14521 ( .C1(n12252), .C2(n12551), .A(n12251), .B(n12250), .ZN(
        n12253) );
  OAI33_X1 U14522 ( .A1(n12312), .A2(n12255), .A3(n12273), .B1(n12528), .B2(
        n12254), .B3(n12253), .ZN(n12257) );
  INV_X1 U14523 ( .A(n12256), .ZN(n12508) );
  NAND3_X1 U14524 ( .A1(n12257), .A2(n12508), .A3(n12520), .ZN(n12266) );
  INV_X1 U14525 ( .A(n12258), .ZN(n12261) );
  XNOR2_X1 U14526 ( .A(n12259), .B(n12277), .ZN(n12260) );
  OAI211_X1 U14527 ( .C1(n7265), .C2(n12261), .A(n12508), .B(n12260), .ZN(
        n12265) );
  MUX2_X1 U14528 ( .A(n12263), .B(n12262), .S(n12273), .Z(n12264) );
  NAND4_X1 U14529 ( .A1(n12266), .A2(n12497), .A3(n12265), .A4(n12264), .ZN(
        n12271) );
  INV_X1 U14530 ( .A(n12267), .ZN(n12268) );
  MUX2_X1 U14531 ( .A(n12269), .B(n12268), .S(n12273), .Z(n12270) );
  OAI21_X1 U14532 ( .B1(n12274), .B2(n12273), .A(n12272), .ZN(n12281) );
  INV_X1 U14533 ( .A(n12275), .ZN(n12280) );
  NAND3_X1 U14534 ( .A1(n12276), .A2(n12490), .A3(n12308), .ZN(n12278) );
  AOI21_X1 U14535 ( .B1(n12282), .B2(n12278), .A(n12277), .ZN(n12279) );
  AOI211_X1 U14536 ( .C1(n12282), .C2(n12281), .A(n12280), .B(n12279), .ZN(
        n12288) );
  INV_X1 U14537 ( .A(n12283), .ZN(n12287) );
  INV_X1 U14538 ( .A(n12284), .ZN(n12286) );
  OAI22_X1 U14539 ( .A1(n12288), .A2(n12287), .B1(n12286), .B2(n12285), .ZN(
        n12289) );
  MUX2_X1 U14540 ( .A(n12290), .B(n14955), .S(n12289), .Z(n12291) );
  OAI21_X1 U14541 ( .B1(n12293), .B2(n12292), .A(n12291), .ZN(n12294) );
  AOI21_X1 U14542 ( .B1(n12296), .B2(n12295), .A(n12294), .ZN(n12305) );
  NAND4_X1 U14543 ( .A1(n12300), .A2(n12299), .A3(n12298), .A4(n12297), .ZN(
        n12301) );
  OAI211_X1 U14544 ( .C1(n12302), .C2(n12304), .A(n12301), .B(P3_B_REG_SCAN_IN), .ZN(n12303) );
  OAI21_X1 U14545 ( .B1(n12305), .B2(n12304), .A(n12303), .ZN(P3_U3296) );
  MUX2_X1 U14546 ( .A(n6619), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12333), .Z(
        P3_U3522) );
  MUX2_X1 U14547 ( .A(n12306), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12333), .Z(
        P3_U3521) );
  MUX2_X1 U14548 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12307), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14549 ( .A(n12308), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12333), .Z(
        P3_U3518) );
  MUX2_X1 U14550 ( .A(n12309), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12333), .Z(
        P3_U3517) );
  MUX2_X1 U14551 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12310), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14552 ( .A(n12311), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12333), .Z(
        P3_U3515) );
  MUX2_X1 U14553 ( .A(n12312), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12333), .Z(
        P3_U3514) );
  MUX2_X1 U14554 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12313), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14555 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12314), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14556 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12315), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14557 ( .A(n12316), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12333), .Z(
        P3_U3510) );
  MUX2_X1 U14558 ( .A(n12317), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12333), .Z(
        P3_U3509) );
  MUX2_X1 U14559 ( .A(n12318), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12333), .Z(
        P3_U3507) );
  MUX2_X1 U14560 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12319), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14561 ( .A(n12320), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12333), .Z(
        P3_U3505) );
  MUX2_X1 U14562 ( .A(n12321), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12333), .Z(
        P3_U3504) );
  MUX2_X1 U14563 ( .A(n12322), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12333), .Z(
        P3_U3503) );
  MUX2_X1 U14564 ( .A(n12323), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12333), .Z(
        P3_U3502) );
  MUX2_X1 U14565 ( .A(n12324), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12333), .Z(
        P3_U3501) );
  MUX2_X1 U14566 ( .A(n12325), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12333), .Z(
        P3_U3500) );
  MUX2_X1 U14567 ( .A(n12326), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12333), .Z(
        P3_U3499) );
  MUX2_X1 U14568 ( .A(n12327), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12333), .Z(
        P3_U3498) );
  MUX2_X1 U14569 ( .A(n12328), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12333), .Z(
        P3_U3497) );
  MUX2_X1 U14570 ( .A(n12329), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12333), .Z(
        P3_U3496) );
  MUX2_X1 U14571 ( .A(n12330), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12333), .Z(
        P3_U3495) );
  MUX2_X1 U14572 ( .A(n8845), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12333), .Z(
        P3_U3494) );
  MUX2_X1 U14573 ( .A(n12331), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12333), .Z(
        P3_U3493) );
  MUX2_X1 U14574 ( .A(n12332), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12333), .Z(
        P3_U3492) );
  MUX2_X1 U14575 ( .A(n12334), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12333), .Z(
        P3_U3491) );
  INV_X1 U14576 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n14897) );
  AOI22_X1 U14577 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n12353), .B1(n12383), 
        .B2(n12337), .ZN(n12338) );
  AOI21_X1 U14578 ( .B1(n12339), .B2(n12338), .A(n12363), .ZN(n12362) );
  INV_X1 U14579 ( .A(n12340), .ZN(n12341) );
  NOR2_X1 U14580 ( .A1(n12342), .A2(n12341), .ZN(n14905) );
  MUX2_X1 U14581 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12455), .Z(n12343) );
  XNOR2_X1 U14582 ( .A(n12343), .B(n14899), .ZN(n14904) );
  NOR2_X1 U14583 ( .A1(n12343), .A2(n14899), .ZN(n12345) );
  MUX2_X1 U14584 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12455), .Z(n12370) );
  XNOR2_X1 U14585 ( .A(n12370), .B(n12383), .ZN(n12344) );
  NOR3_X1 U14586 ( .A1(n14903), .A2(n12345), .A3(n12344), .ZN(n12369) );
  NOR2_X1 U14587 ( .A1(n12369), .A2(n14906), .ZN(n12360) );
  OAI21_X1 U14588 ( .B1(n14903), .B2(n12345), .A(n12344), .ZN(n12359) );
  NAND2_X1 U14589 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P3_U3151), .ZN(n12347)
         );
  NAND2_X1 U14590 ( .A1(n14931), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n12346) );
  OAI211_X1 U14591 ( .C1(n14917), .C2(n12383), .A(n12347), .B(n12346), .ZN(
        n12358) );
  INV_X1 U14592 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14902) );
  NOR2_X1 U14593 ( .A1(n12351), .A2(n6524), .ZN(n12352) );
  INV_X1 U14594 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n15132) );
  AOI22_X1 U14595 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n12353), .B1(n12383), 
        .B2(n15132), .ZN(n12354) );
  NOR2_X1 U14596 ( .A1(n12355), .A2(n12354), .ZN(n12385) );
  AOI21_X1 U14597 ( .B1(n12355), .B2(n12354), .A(n12385), .ZN(n12356) );
  NOR2_X1 U14598 ( .A1(n12356), .A2(n14927), .ZN(n12357) );
  AOI211_X1 U14599 ( .C1(n12360), .C2(n12359), .A(n12358), .B(n12357), .ZN(
        n12361) );
  OAI21_X1 U14600 ( .B1(n12362), .B2(n14933), .A(n12361), .ZN(P3_U3194) );
  NOR2_X1 U14601 ( .A1(n12387), .A2(n12364), .ZN(n12365) );
  NOR2_X1 U14602 ( .A1(n11590), .A2(n14914), .ZN(n14913) );
  NAND2_X1 U14603 ( .A1(n14219), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12408) );
  OAI21_X1 U14604 ( .B1(n14219), .B2(P3_REG2_REG_14__SCAN_IN), .A(n12408), 
        .ZN(n12373) );
  AOI21_X1 U14605 ( .B1(n12366), .B2(n12373), .A(n12400), .ZN(n12393) );
  INV_X1 U14606 ( .A(n14219), .ZN(n12382) );
  INV_X1 U14607 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n12367) );
  NAND2_X1 U14608 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(P3_U3151), .ZN(n14255)
         );
  OAI21_X1 U14609 ( .B1(n12368), .B2(n12367), .A(n14255), .ZN(n12381) );
  MUX2_X1 U14610 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12455), .Z(n12371) );
  XNOR2_X1 U14611 ( .A(n12371), .B(n12387), .ZN(n14922) );
  NAND2_X1 U14612 ( .A1(n14923), .A2(n14922), .ZN(n14921) );
  INV_X1 U14613 ( .A(n12371), .ZN(n12372) );
  NAND2_X1 U14614 ( .A1(n12372), .A2(n12387), .ZN(n12377) );
  INV_X1 U14615 ( .A(n12373), .ZN(n12375) );
  AND2_X1 U14616 ( .A1(n14219), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12395) );
  INV_X1 U14617 ( .A(n12395), .ZN(n12407) );
  OAI21_X1 U14618 ( .B1(P3_REG1_REG_14__SCAN_IN), .B2(n14219), .A(n12407), 
        .ZN(n12389) );
  INV_X1 U14619 ( .A(n12389), .ZN(n12374) );
  MUX2_X1 U14620 ( .A(n12375), .B(n12374), .S(n12455), .Z(n12376) );
  NAND3_X1 U14621 ( .A1(n14921), .A2(n12377), .A3(n12376), .ZN(n12410) );
  INV_X1 U14622 ( .A(n12410), .ZN(n12379) );
  AOI21_X1 U14623 ( .B1(n14921), .B2(n12377), .A(n12376), .ZN(n12378) );
  NOR3_X1 U14624 ( .A1(n12379), .A2(n12378), .A3(n14906), .ZN(n12380) );
  AOI211_X1 U14625 ( .C1(n12419), .C2(n12382), .A(n12381), .B(n12380), .ZN(
        n12392) );
  INV_X1 U14626 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14920) );
  AOI21_X1 U14627 ( .B1(n6588), .B2(n12389), .A(n12394), .ZN(n12390) );
  OR2_X1 U14628 ( .A1(n12390), .A2(n14927), .ZN(n12391) );
  OAI211_X1 U14629 ( .C1(n12393), .C2(n14933), .A(n12392), .B(n12391), .ZN(
        P3_U3196) );
  INV_X1 U14630 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12399) );
  INV_X1 U14631 ( .A(n12414), .ZN(n14288) );
  NOR2_X1 U14632 ( .A1(n12412), .A2(n12396), .ZN(n12397) );
  INV_X1 U14633 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14269) );
  INV_X1 U14634 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12658) );
  AOI22_X1 U14635 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12414), .B1(n14288), 
        .B2(n12658), .ZN(n14290) );
  XNOR2_X1 U14636 ( .A(n12421), .B(n12425), .ZN(n12398) );
  AOI21_X1 U14637 ( .B1(n12399), .B2(n12398), .A(n12422), .ZN(n12420) );
  INV_X1 U14638 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12403) );
  INV_X1 U14639 ( .A(n12412), .ZN(n14266) );
  AND2_X1 U14640 ( .A1(n14266), .A2(n12401), .ZN(n12402) );
  INV_X1 U14641 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14263) );
  INV_X1 U14642 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12609) );
  AOI22_X1 U14643 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12414), .B1(n14288), 
        .B2(n12609), .ZN(n14279) );
  MUX2_X1 U14644 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12455), .Z(n12438) );
  XOR2_X1 U14645 ( .A(n12425), .B(n12438), .Z(n12417) );
  MUX2_X1 U14646 ( .A(n12408), .B(n12407), .S(n12455), .Z(n12409) );
  NAND2_X1 U14647 ( .A1(n12410), .A2(n12409), .ZN(n12411) );
  INV_X1 U14648 ( .A(n12411), .ZN(n12413) );
  XNOR2_X1 U14649 ( .A(n12411), .B(n14266), .ZN(n14271) );
  MUX2_X1 U14650 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12455), .Z(n14272) );
  AOI21_X1 U14651 ( .B1(n12413), .B2(n12412), .A(n14270), .ZN(n14285) );
  MUX2_X1 U14652 ( .A(n12609), .B(n12658), .S(n12455), .Z(n12415) );
  NOR2_X1 U14653 ( .A1(n12415), .A2(n12414), .ZN(n14281) );
  NAND2_X1 U14654 ( .A1(n12415), .A2(n12414), .ZN(n14282) );
  OAI21_X1 U14655 ( .B1(n14285), .B2(n14281), .A(n14282), .ZN(n12416) );
  NOR2_X1 U14656 ( .A1(n12416), .A2(n12417), .ZN(n12436) );
  AOI211_X1 U14657 ( .C1(n12417), .C2(n12416), .A(n14906), .B(n12436), .ZN(
        n12418) );
  NAND2_X1 U14658 ( .A1(n12452), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12461) );
  OAI21_X1 U14659 ( .B1(n12452), .B2(P3_REG1_REG_18__SCAN_IN), .A(n12461), 
        .ZN(n12424) );
  INV_X1 U14660 ( .A(n12460), .ZN(n12423) );
  AOI21_X1 U14661 ( .B1(n6581), .B2(n12424), .A(n12423), .ZN(n12447) );
  NOR2_X1 U14662 ( .A1(n12426), .A2(n12425), .ZN(n12428) );
  INV_X1 U14663 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12586) );
  AND2_X1 U14664 ( .A1(n12452), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12448) );
  AOI21_X1 U14665 ( .B1(n12427), .B2(n12586), .A(n12448), .ZN(n12430) );
  NOR3_X1 U14666 ( .A1(n12428), .A2(n12429), .A3(n12430), .ZN(n12435) );
  INV_X1 U14667 ( .A(n12428), .ZN(n12433) );
  INV_X1 U14668 ( .A(n12429), .ZN(n12432) );
  INV_X1 U14669 ( .A(n12430), .ZN(n12431) );
  OAI21_X1 U14670 ( .B1(n12435), .B2(n12449), .A(n12434), .ZN(n12446) );
  AOI21_X1 U14671 ( .B1(n12438), .B2(n12437), .A(n12436), .ZN(n12450) );
  XNOR2_X1 U14672 ( .A(n12450), .B(n12452), .ZN(n12440) );
  INV_X1 U14673 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12652) );
  MUX2_X1 U14674 ( .A(n12586), .B(n12652), .S(n12455), .Z(n12439) );
  NAND2_X1 U14675 ( .A1(n12440), .A2(n12439), .ZN(n12451) );
  OAI21_X1 U14676 ( .B1(n12440), .B2(n12439), .A(n12451), .ZN(n12444) );
  NAND2_X1 U14677 ( .A1(n14931), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n12441) );
  OAI211_X1 U14678 ( .C1(n14917), .C2(n12452), .A(n12442), .B(n12441), .ZN(
        n12443) );
  AOI21_X1 U14679 ( .B1(n12444), .B2(n14924), .A(n12443), .ZN(n12445) );
  OAI211_X1 U14680 ( .C1(n12447), .C2(n14927), .A(n12446), .B(n12445), .ZN(
        P3_U3200) );
  XNOR2_X1 U14681 ( .A(n12454), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12456) );
  INV_X1 U14682 ( .A(n12450), .ZN(n12453) );
  OAI21_X1 U14683 ( .B1(n12453), .B2(n12452), .A(n12451), .ZN(n12458) );
  XNOR2_X1 U14684 ( .A(n12454), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12462) );
  MUX2_X1 U14685 ( .A(n12456), .B(n12462), .S(n12455), .Z(n12457) );
  XNOR2_X1 U14686 ( .A(n12458), .B(n12457), .ZN(n12468) );
  NOR2_X1 U14687 ( .A1(n14917), .A2(n12459), .ZN(n12467) );
  INV_X1 U14688 ( .A(n12462), .ZN(n12463) );
  NAND2_X1 U14689 ( .A1(n14931), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12465) );
  AOI21_X1 U14690 ( .B1(n12666), .B2(n14963), .A(n12470), .ZN(n12473) );
  NAND2_X1 U14691 ( .A1(n14965), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12471) );
  OAI211_X1 U14692 ( .C1(n6620), .C2(n12489), .A(n12473), .B(n12471), .ZN(
        P3_U3202) );
  NAND2_X1 U14693 ( .A1(n14965), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n12472) );
  OAI211_X1 U14694 ( .C1(n12626), .C2(n12489), .A(n12473), .B(n12472), .ZN(
        P3_U3203) );
  INV_X1 U14695 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12475) );
  INV_X1 U14696 ( .A(n12673), .ZN(n12474) );
  AOI22_X1 U14697 ( .A1(n12477), .A2(n12618), .B1(n14959), .B2(n12476), .ZN(
        n12478) );
  OAI211_X1 U14698 ( .C1(n12621), .C2(n12675), .A(n12479), .B(n12478), .ZN(
        P3_U3205) );
  OAI21_X1 U14699 ( .B1(n12485), .B2(n12481), .A(n12480), .ZN(n12483) );
  AOI21_X1 U14700 ( .B1(n12483), .B2(n14948), .A(n12482), .ZN(n12629) );
  AOI21_X1 U14701 ( .B1(n12486), .B2(n12485), .A(n12484), .ZN(n12630) );
  INV_X1 U14702 ( .A(n12630), .ZN(n12493) );
  AOI22_X1 U14703 ( .A1(n14965), .A2(P3_REG2_REG_27__SCAN_IN), .B1(n14959), 
        .B2(n12487), .ZN(n12488) );
  OAI21_X1 U14704 ( .B1(n12490), .B2(n12489), .A(n12488), .ZN(n12491) );
  AOI21_X1 U14705 ( .B1(n12493), .B2(n12492), .A(n12491), .ZN(n12494) );
  OAI21_X1 U14706 ( .B1(n12629), .B2(n14965), .A(n12494), .ZN(P3_U3206) );
  XOR2_X1 U14707 ( .A(n12497), .B(n12495), .Z(n12681) );
  INV_X1 U14708 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12501) );
  XOR2_X1 U14709 ( .A(n12497), .B(n12496), .Z(n12499) );
  INV_X1 U14710 ( .A(n12679), .ZN(n12500) );
  AOI22_X1 U14711 ( .A1(n12503), .A2(n12618), .B1(n14959), .B2(n12502), .ZN(
        n12504) );
  OAI211_X1 U14712 ( .C1(n12621), .C2(n12681), .A(n12505), .B(n12504), .ZN(
        P3_U3207) );
  XNOR2_X1 U14713 ( .A(n12506), .B(n12508), .ZN(n12686) );
  INV_X1 U14714 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n12514) );
  NAND2_X1 U14715 ( .A1(n12508), .A2(n12507), .ZN(n12510) );
  OAI211_X1 U14716 ( .C1(n6522), .C2(n12510), .A(n12509), .B(n14948), .ZN(
        n12512) );
  NAND2_X1 U14717 ( .A1(n12512), .A2(n12511), .ZN(n12684) );
  INV_X1 U14718 ( .A(n12684), .ZN(n12513) );
  MUX2_X1 U14719 ( .A(n12514), .B(n12513), .S(n14963), .Z(n12518) );
  AOI22_X1 U14720 ( .A1(n12516), .A2(n12618), .B1(n14959), .B2(n12515), .ZN(
        n12517) );
  OAI211_X1 U14721 ( .C1(n12621), .C2(n12686), .A(n12518), .B(n12517), .ZN(
        P3_U3208) );
  AOI21_X1 U14722 ( .B1(n7265), .B2(n12519), .A(n6536), .ZN(n12694) );
  INV_X1 U14723 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12524) );
  AOI211_X1 U14724 ( .C1(n12521), .C2(n12520), .A(n14939), .B(n6522), .ZN(
        n12523) );
  NOR2_X1 U14725 ( .A1(n12523), .A2(n12522), .ZN(n12689) );
  MUX2_X1 U14726 ( .A(n12524), .B(n12689), .S(n14963), .Z(n12527) );
  AOI22_X1 U14727 ( .A1(n12691), .A2(n12618), .B1(n14959), .B2(n12525), .ZN(
        n12526) );
  OAI211_X1 U14728 ( .C1(n12621), .C2(n12694), .A(n12527), .B(n12526), .ZN(
        P3_U3209) );
  XNOR2_X1 U14729 ( .A(n12529), .B(n12528), .ZN(n12700) );
  INV_X1 U14730 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12535) );
  NOR2_X1 U14731 ( .A1(n12534), .A2(n12533), .ZN(n12695) );
  MUX2_X1 U14732 ( .A(n12535), .B(n12695), .S(n14963), .Z(n12538) );
  AOI22_X1 U14733 ( .A1(n12697), .A2(n12618), .B1(n14959), .B2(n12536), .ZN(
        n12537) );
  OAI211_X1 U14734 ( .C1(n12621), .C2(n12700), .A(n12538), .B(n12537), .ZN(
        P3_U3210) );
  XNOR2_X1 U14735 ( .A(n12539), .B(n12540), .ZN(n12706) );
  INV_X1 U14736 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12544) );
  XNOR2_X1 U14737 ( .A(n12541), .B(n12540), .ZN(n12543) );
  AOI21_X1 U14738 ( .B1(n12543), .B2(n14948), .A(n12542), .ZN(n12701) );
  MUX2_X1 U14739 ( .A(n12544), .B(n12701), .S(n14963), .Z(n12547) );
  AOI22_X1 U14740 ( .A1(n12703), .A2(n12618), .B1(n14959), .B2(n12545), .ZN(
        n12546) );
  OAI211_X1 U14741 ( .C1(n12621), .C2(n12706), .A(n12547), .B(n12546), .ZN(
        P3_U3211) );
  XOR2_X1 U14742 ( .A(n12551), .B(n12548), .Z(n12709) );
  INV_X1 U14743 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12555) );
  AOI21_X1 U14744 ( .B1(n12551), .B2(n12550), .A(n12549), .ZN(n12553) );
  OAI21_X1 U14745 ( .B1(n12553), .B2(n14939), .A(n12552), .ZN(n12707) );
  INV_X1 U14746 ( .A(n12707), .ZN(n12554) );
  MUX2_X1 U14747 ( .A(n12555), .B(n12554), .S(n14963), .Z(n12559) );
  AOI22_X1 U14748 ( .A1(n12557), .A2(n12618), .B1(n14959), .B2(n12556), .ZN(
        n12558) );
  OAI211_X1 U14749 ( .C1(n12621), .C2(n12709), .A(n12559), .B(n12558), .ZN(
        P3_U3212) );
  XNOR2_X1 U14750 ( .A(n12561), .B(n12560), .ZN(n12717) );
  INV_X1 U14751 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12566) );
  XNOR2_X1 U14752 ( .A(n12563), .B(n12562), .ZN(n12565) );
  AOI21_X1 U14753 ( .B1(n12565), .B2(n14948), .A(n12564), .ZN(n12712) );
  MUX2_X1 U14754 ( .A(n12566), .B(n12712), .S(n14963), .Z(n12569) );
  AOI22_X1 U14755 ( .A1(n12714), .A2(n12618), .B1(n14959), .B2(n12567), .ZN(
        n12568) );
  OAI211_X1 U14756 ( .C1(n12621), .C2(n12717), .A(n12569), .B(n12568), .ZN(
        P3_U3213) );
  XNOR2_X1 U14757 ( .A(n12570), .B(n12571), .ZN(n12723) );
  INV_X1 U14758 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12574) );
  XOR2_X1 U14759 ( .A(n12571), .B(n6478), .Z(n12573) );
  AOI21_X1 U14760 ( .B1(n12573), .B2(n14948), .A(n12572), .ZN(n12718) );
  MUX2_X1 U14761 ( .A(n12574), .B(n12718), .S(n14963), .Z(n12577) );
  AOI22_X1 U14762 ( .A1(n12720), .A2(n12618), .B1(n12575), .B2(n14959), .ZN(
        n12576) );
  OAI211_X1 U14763 ( .C1(n12621), .C2(n12723), .A(n12577), .B(n12576), .ZN(
        P3_U3214) );
  AOI21_X1 U14764 ( .B1(n12579), .B2(n12578), .A(n6590), .ZN(n12580) );
  INV_X1 U14765 ( .A(n12580), .ZN(n12729) );
  OAI21_X1 U14766 ( .B1(n12595), .B2(n12582), .A(n12581), .ZN(n12583) );
  AOI21_X1 U14767 ( .B1(n7250), .B2(n12583), .A(n14939), .ZN(n12585) );
  NOR2_X1 U14768 ( .A1(n12585), .A2(n12584), .ZN(n12724) );
  MUX2_X1 U14769 ( .A(n12586), .B(n12724), .S(n14963), .Z(n12589) );
  AOI22_X1 U14770 ( .A1(n12726), .A2(n12618), .B1(n14959), .B2(n12587), .ZN(
        n12588) );
  OAI211_X1 U14771 ( .C1(n12621), .C2(n12729), .A(n12589), .B(n12588), .ZN(
        P3_U3215) );
  XNOR2_X1 U14772 ( .A(n12590), .B(n12591), .ZN(n12732) );
  NAND2_X1 U14773 ( .A1(n12592), .A2(n12591), .ZN(n12593) );
  NAND2_X1 U14774 ( .A1(n12593), .A2(n14948), .ZN(n12594) );
  OR2_X1 U14775 ( .A1(n12595), .A2(n12594), .ZN(n12597) );
  NAND2_X1 U14776 ( .A1(n12597), .A2(n12596), .ZN(n12733) );
  MUX2_X1 U14777 ( .A(P3_REG2_REG_17__SCAN_IN), .B(n12733), .S(n14963), .Z(
        n12598) );
  INV_X1 U14778 ( .A(n12598), .ZN(n12602) );
  AOI22_X1 U14779 ( .A1(n12600), .A2(n12618), .B1(n14959), .B2(n12599), .ZN(
        n12601) );
  OAI211_X1 U14780 ( .C1(n12621), .C2(n12732), .A(n12602), .B(n12601), .ZN(
        P3_U3216) );
  XOR2_X1 U14781 ( .A(n12606), .B(n12603), .Z(n12741) );
  AOI22_X1 U14782 ( .A1(n12738), .A2(n12618), .B1(n14959), .B2(n12604), .ZN(
        n12611) );
  XNOR2_X1 U14783 ( .A(n12605), .B(n12606), .ZN(n12608) );
  AOI21_X1 U14784 ( .B1(n12608), .B2(n14948), .A(n12607), .ZN(n12736) );
  MUX2_X1 U14785 ( .A(n12609), .B(n12736), .S(n14963), .Z(n12610) );
  OAI211_X1 U14786 ( .C1(n12741), .C2(n12621), .A(n12611), .B(n12610), .ZN(
        P3_U3217) );
  XOR2_X1 U14787 ( .A(n12614), .B(n12612), .Z(n12749) );
  XOR2_X1 U14788 ( .A(n12613), .B(n12614), .Z(n12616) );
  AOI21_X1 U14789 ( .B1(n12616), .B2(n14948), .A(n12615), .ZN(n12742) );
  MUX2_X1 U14790 ( .A(n14263), .B(n12742), .S(n14963), .Z(n12620) );
  AOI22_X1 U14791 ( .A1(n12745), .A2(n12618), .B1(n14959), .B2(n12617), .ZN(
        n12619) );
  OAI211_X1 U14792 ( .C1(n12621), .C2(n12749), .A(n12620), .B(n12619), .ZN(
        P3_U3218) );
  INV_X1 U14793 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12623) );
  NAND2_X1 U14794 ( .A1(n12665), .A2(n12661), .ZN(n12622) );
  NAND2_X1 U14795 ( .A1(n12666), .A2(n15034), .ZN(n12625) );
  OAI211_X1 U14796 ( .C1(n15034), .C2(n12623), .A(n12622), .B(n12625), .ZN(
        P3_U3490) );
  NAND2_X1 U14797 ( .A1(n15039), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n12624) );
  OAI211_X1 U14798 ( .C1(n12626), .C2(n12655), .A(n12625), .B(n12624), .ZN(
        P3_U3489) );
  INV_X1 U14799 ( .A(n15007), .ZN(n14304) );
  NAND2_X1 U14800 ( .A1(n12627), .A2(n15014), .ZN(n12628) );
  OAI211_X1 U14801 ( .C1(n14304), .C2(n12630), .A(n12629), .B(n12628), .ZN(
        n12678) );
  MUX2_X1 U14802 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n12678), .S(n15034), .Z(
        P3_U3486) );
  MUX2_X1 U14803 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n12679), .S(n15034), .Z(
        n12632) );
  OAI22_X1 U14804 ( .A1(n12681), .A2(n12664), .B1(n12680), .B2(n12655), .ZN(
        n12631) );
  OR2_X1 U14805 ( .A1(n12632), .A2(n12631), .ZN(P3_U3485) );
  MUX2_X1 U14806 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n12684), .S(n15034), .Z(
        n12634) );
  OAI22_X1 U14807 ( .A1(n12686), .A2(n12664), .B1(n12685), .B2(n12655), .ZN(
        n12633) );
  OR2_X1 U14808 ( .A1(n12634), .A2(n12633), .ZN(P3_U3484) );
  INV_X1 U14809 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12635) );
  MUX2_X1 U14810 ( .A(n12635), .B(n12689), .S(n15034), .Z(n12637) );
  NAND2_X1 U14811 ( .A1(n12691), .A2(n12661), .ZN(n12636) );
  OAI211_X1 U14812 ( .C1(n12694), .C2(n12664), .A(n12637), .B(n12636), .ZN(
        P3_U3483) );
  INV_X1 U14813 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12638) );
  MUX2_X1 U14814 ( .A(n12638), .B(n12695), .S(n15034), .Z(n12640) );
  NAND2_X1 U14815 ( .A1(n12697), .A2(n12661), .ZN(n12639) );
  OAI211_X1 U14816 ( .C1(n12664), .C2(n12700), .A(n12640), .B(n12639), .ZN(
        P3_U3482) );
  INV_X1 U14817 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12641) );
  MUX2_X1 U14818 ( .A(n12641), .B(n12701), .S(n15034), .Z(n12643) );
  NAND2_X1 U14819 ( .A1(n12703), .A2(n12661), .ZN(n12642) );
  OAI211_X1 U14820 ( .C1(n12706), .C2(n12664), .A(n12643), .B(n12642), .ZN(
        P3_U3481) );
  MUX2_X1 U14821 ( .A(P3_REG1_REG_21__SCAN_IN), .B(n12707), .S(n15034), .Z(
        n12645) );
  OAI22_X1 U14822 ( .A1(n12709), .A2(n12664), .B1(n12708), .B2(n12655), .ZN(
        n12644) );
  OR2_X1 U14823 ( .A1(n12645), .A2(n12644), .ZN(P3_U3480) );
  INV_X1 U14824 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12646) );
  MUX2_X1 U14825 ( .A(n12646), .B(n12712), .S(n15034), .Z(n12648) );
  NAND2_X1 U14826 ( .A1(n12714), .A2(n12661), .ZN(n12647) );
  OAI211_X1 U14827 ( .C1(n12664), .C2(n12717), .A(n12648), .B(n12647), .ZN(
        P3_U3479) );
  INV_X1 U14828 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12649) );
  MUX2_X1 U14829 ( .A(n12649), .B(n12718), .S(n15034), .Z(n12651) );
  NAND2_X1 U14830 ( .A1(n12720), .A2(n12661), .ZN(n12650) );
  OAI211_X1 U14831 ( .C1(n12723), .C2(n12664), .A(n12651), .B(n12650), .ZN(
        P3_U3478) );
  MUX2_X1 U14832 ( .A(n12652), .B(n12724), .S(n15034), .Z(n12654) );
  NAND2_X1 U14833 ( .A1(n12726), .A2(n12661), .ZN(n12653) );
  OAI211_X1 U14834 ( .C1(n12664), .C2(n12729), .A(n12654), .B(n12653), .ZN(
        P3_U3477) );
  OAI22_X1 U14835 ( .A1(n12732), .A2(n12664), .B1(n12731), .B2(n12655), .ZN(
        n12657) );
  MUX2_X1 U14836 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12733), .S(n15034), .Z(
        n12656) );
  OR2_X1 U14837 ( .A1(n12657), .A2(n12656), .ZN(P3_U3476) );
  MUX2_X1 U14838 ( .A(n12658), .B(n12736), .S(n15034), .Z(n12660) );
  NAND2_X1 U14839 ( .A1(n12738), .A2(n12661), .ZN(n12659) );
  OAI211_X1 U14840 ( .C1(n12741), .C2(n12664), .A(n12660), .B(n12659), .ZN(
        P3_U3475) );
  MUX2_X1 U14841 ( .A(n14269), .B(n12742), .S(n15034), .Z(n12663) );
  NAND2_X1 U14842 ( .A1(n12745), .A2(n12661), .ZN(n12662) );
  OAI211_X1 U14843 ( .C1(n12664), .C2(n12749), .A(n12663), .B(n12662), .ZN(
        P3_U3474) );
  INV_X1 U14844 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12668) );
  NAND2_X1 U14845 ( .A1(n12665), .A2(n12744), .ZN(n12667) );
  NAND2_X1 U14846 ( .A1(n12666), .A2(n15025), .ZN(n12670) );
  OAI211_X1 U14847 ( .C1(n15025), .C2(n12668), .A(n12667), .B(n12670), .ZN(
        P3_U3458) );
  INV_X1 U14848 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n12672) );
  NAND2_X1 U14849 ( .A1(n12669), .A2(n12744), .ZN(n12671) );
  OAI211_X1 U14850 ( .C1(n15025), .C2(n12672), .A(n12671), .B(n12670), .ZN(
        P3_U3457) );
  OAI22_X1 U14851 ( .A1(n12675), .A2(n12748), .B1(n12674), .B2(n12730), .ZN(
        n12676) );
  MUX2_X1 U14852 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n12678), .S(n15025), .Z(
        P3_U3454) );
  MUX2_X1 U14853 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n12679), .S(n15025), .Z(
        n12683) );
  OAI22_X1 U14854 ( .A1(n12681), .A2(n12748), .B1(n12680), .B2(n12730), .ZN(
        n12682) );
  OR2_X1 U14855 ( .A1(n12683), .A2(n12682), .ZN(P3_U3453) );
  MUX2_X1 U14856 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n12684), .S(n15025), .Z(
        n12688) );
  OAI22_X1 U14857 ( .A1(n12686), .A2(n12748), .B1(n12685), .B2(n12730), .ZN(
        n12687) );
  OR2_X1 U14858 ( .A1(n12688), .A2(n12687), .ZN(P3_U3452) );
  INV_X1 U14859 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12690) );
  MUX2_X1 U14860 ( .A(n12690), .B(n12689), .S(n15025), .Z(n12693) );
  NAND2_X1 U14861 ( .A1(n12691), .A2(n12744), .ZN(n12692) );
  OAI211_X1 U14862 ( .C1(n12694), .C2(n12748), .A(n12693), .B(n12692), .ZN(
        P3_U3451) );
  INV_X1 U14863 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12696) );
  MUX2_X1 U14864 ( .A(n12696), .B(n12695), .S(n15025), .Z(n12699) );
  NAND2_X1 U14865 ( .A1(n12697), .A2(n12744), .ZN(n12698) );
  OAI211_X1 U14866 ( .C1(n12700), .C2(n12748), .A(n12699), .B(n12698), .ZN(
        P3_U3450) );
  INV_X1 U14867 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12702) );
  MUX2_X1 U14868 ( .A(n12702), .B(n12701), .S(n15025), .Z(n12705) );
  NAND2_X1 U14869 ( .A1(n12703), .A2(n12744), .ZN(n12704) );
  OAI211_X1 U14870 ( .C1(n12706), .C2(n12748), .A(n12705), .B(n12704), .ZN(
        P3_U3449) );
  MUX2_X1 U14871 ( .A(P3_REG0_REG_21__SCAN_IN), .B(n12707), .S(n15025), .Z(
        n12711) );
  OAI22_X1 U14872 ( .A1(n12709), .A2(n12748), .B1(n12708), .B2(n12730), .ZN(
        n12710) );
  OR2_X1 U14873 ( .A1(n12711), .A2(n12710), .ZN(P3_U3448) );
  INV_X1 U14874 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12713) );
  MUX2_X1 U14875 ( .A(n12713), .B(n12712), .S(n15025), .Z(n12716) );
  NAND2_X1 U14876 ( .A1(n12714), .A2(n12744), .ZN(n12715) );
  OAI211_X1 U14877 ( .C1(n12717), .C2(n12748), .A(n12716), .B(n12715), .ZN(
        P3_U3447) );
  INV_X1 U14878 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12719) );
  MUX2_X1 U14879 ( .A(n12719), .B(n12718), .S(n15025), .Z(n12722) );
  NAND2_X1 U14880 ( .A1(n12720), .A2(n12744), .ZN(n12721) );
  OAI211_X1 U14881 ( .C1(n12723), .C2(n12748), .A(n12722), .B(n12721), .ZN(
        P3_U3446) );
  INV_X1 U14882 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12725) );
  MUX2_X1 U14883 ( .A(n12725), .B(n12724), .S(n15025), .Z(n12728) );
  NAND2_X1 U14884 ( .A1(n12726), .A2(n12744), .ZN(n12727) );
  OAI211_X1 U14885 ( .C1(n12729), .C2(n12748), .A(n12728), .B(n12727), .ZN(
        P3_U3444) );
  OAI22_X1 U14886 ( .A1(n12732), .A2(n12748), .B1(n12731), .B2(n12730), .ZN(
        n12735) );
  MUX2_X1 U14887 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n12733), .S(n15025), .Z(
        n12734) );
  OR2_X1 U14888 ( .A1(n12735), .A2(n12734), .ZN(P3_U3441) );
  INV_X1 U14889 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12737) );
  MUX2_X1 U14890 ( .A(n12737), .B(n12736), .S(n15025), .Z(n12740) );
  NAND2_X1 U14891 ( .A1(n12738), .A2(n12744), .ZN(n12739) );
  OAI211_X1 U14892 ( .C1(n12741), .C2(n12748), .A(n12740), .B(n12739), .ZN(
        P3_U3438) );
  INV_X1 U14893 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12743) );
  MUX2_X1 U14894 ( .A(n12743), .B(n12742), .S(n15025), .Z(n12747) );
  NAND2_X1 U14895 ( .A1(n12745), .A2(n12744), .ZN(n12746) );
  OAI211_X1 U14896 ( .C1(n12749), .C2(n12748), .A(n12747), .B(n12746), .ZN(
        P3_U3435) );
  MUX2_X1 U14897 ( .A(n12750), .B(P3_D_REG_1__SCAN_IN), .S(n12751), .Z(
        P3_U3377) );
  MUX2_X1 U14898 ( .A(n12752), .B(P3_D_REG_0__SCAN_IN), .S(n12751), .Z(
        P3_U3376) );
  NAND3_X1 U14899 ( .A1(n8773), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n12755) );
  OAI22_X1 U14900 ( .A1(n12753), .A2(n12755), .B1(n12754), .B2(n14213), .ZN(
        n12756) );
  AOI21_X1 U14901 ( .B1(n12757), .B2(n14223), .A(n12756), .ZN(n12758) );
  INV_X1 U14902 ( .A(n12758), .ZN(P3_U3264) );
  INV_X1 U14903 ( .A(n12759), .ZN(n12761) );
  OAI222_X1 U14904 ( .A1(n14213), .A2(n12762), .B1(n14215), .B2(n12761), .C1(
        n12760), .C2(P3_U3151), .ZN(P3_U3266) );
  INV_X1 U14905 ( .A(n12763), .ZN(n12765) );
  NAND2_X1 U14906 ( .A1(n12767), .A2(n12766), .ZN(n12768) );
  NAND3_X1 U14907 ( .A1(n12769), .A2(n12865), .A3(n12768), .ZN(n12774) );
  OAI22_X1 U14908 ( .A1(n12856), .A2(n13003), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15074), .ZN(n12771) );
  OAI22_X1 U14909 ( .A1(n12977), .A2(n12869), .B1(n12814), .B2(n12847), .ZN(
        n12770) );
  AOI211_X1 U14910 ( .C1(n12772), .C2(n12871), .A(n12771), .B(n12770), .ZN(
        n12773) );
  NAND2_X1 U14911 ( .A1(n12774), .A2(n12773), .ZN(P2_U3186) );
  NAND2_X1 U14912 ( .A1(n12841), .A2(n13080), .ZN(n12778) );
  NAND2_X1 U14913 ( .A1(n12865), .A2(n12775), .ZN(n12777) );
  MUX2_X1 U14914 ( .A(n12778), .B(n12777), .S(n12776), .Z(n12784) );
  OAI22_X1 U14915 ( .A1(n12856), .A2(n12780), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12779), .ZN(n12782) );
  OAI22_X1 U14916 ( .A1(n13066), .A2(n12847), .B1(n12869), .B2(n13068), .ZN(
        n12781) );
  AOI211_X1 U14917 ( .C1(n13226), .C2(n12871), .A(n12782), .B(n12781), .ZN(
        n12783) );
  NAND2_X1 U14918 ( .A1(n12784), .A2(n12783), .ZN(P2_U3188) );
  INV_X1 U14919 ( .A(n12785), .ZN(n12857) );
  NOR3_X1 U14920 ( .A1(n12787), .A2(n12786), .A3(n12872), .ZN(n12788) );
  AOI21_X1 U14921 ( .B1(n12857), .B2(n12865), .A(n12788), .ZN(n12796) );
  OR2_X1 U14922 ( .A1(n12797), .A2(n13069), .ZN(n12790) );
  NAND2_X1 U14923 ( .A1(n13152), .A2(n12882), .ZN(n12789) );
  NAND2_X1 U14924 ( .A1(n12790), .A2(n12789), .ZN(n13130) );
  NAND2_X1 U14925 ( .A1(n12798), .A2(n13130), .ZN(n12791) );
  NAND2_X1 U14926 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n12946)
         );
  OAI211_X1 U14927 ( .C1(n12856), .C2(n13134), .A(n12791), .B(n12946), .ZN(
        n12793) );
  NOR2_X1 U14928 ( .A1(n12837), .A2(n12858), .ZN(n12792) );
  AOI211_X1 U14929 ( .C1(n13246), .C2(n12871), .A(n12793), .B(n12792), .ZN(
        n12794) );
  OAI21_X1 U14930 ( .B1(n12796), .B2(n12795), .A(n12794), .ZN(P2_U3191) );
  OAI22_X1 U14931 ( .A1(n13066), .A2(n13069), .B1(n12797), .B2(n13067), .ZN(
        n13096) );
  AOI22_X1 U14932 ( .A1(n12798), .A2(n13096), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12799) );
  OAI21_X1 U14933 ( .B1(n13100), .B2(n12856), .A(n12799), .ZN(n12805) );
  INV_X1 U14934 ( .A(n12800), .ZN(n12801) );
  AOI211_X1 U14935 ( .C1(n12803), .C2(n12802), .A(n12858), .B(n12801), .ZN(
        n12804) );
  AOI211_X1 U14936 ( .C1(n13236), .C2(n12871), .A(n12805), .B(n12804), .ZN(
        n12806) );
  INV_X1 U14937 ( .A(n12806), .ZN(P2_U3195) );
  INV_X1 U14938 ( .A(n12808), .ZN(n12809) );
  AOI21_X1 U14939 ( .B1(n12807), .B2(n12809), .A(n12858), .ZN(n12813) );
  NOR3_X1 U14940 ( .A1(n12810), .A2(n13068), .A3(n12872), .ZN(n12812) );
  OAI21_X1 U14941 ( .B1(n12813), .B2(n12812), .A(n12811), .ZN(n12818) );
  NOR2_X1 U14942 ( .A1(n12856), .A2(n13041), .ZN(n12816) );
  OAI22_X1 U14943 ( .A1(n12814), .A2(n12869), .B1(n12847), .B2(n13068), .ZN(
        n12815) );
  AOI211_X1 U14944 ( .C1(P2_REG3_REG_25__SCAN_IN), .C2(P2_U3088), .A(n12816), 
        .B(n12815), .ZN(n12817) );
  OAI211_X1 U14945 ( .C1(n13038), .C2(n12829), .A(n12818), .B(n12817), .ZN(
        P2_U3197) );
  AOI21_X1 U14946 ( .B1(n12820), .B2(n12819), .A(n12858), .ZN(n12821) );
  NAND2_X1 U14947 ( .A1(n12821), .A2(n12807), .ZN(n12825) );
  AOI22_X1 U14948 ( .A1(n13017), .A2(n13153), .B1(n13152), .B2(n13080), .ZN(
        n13049) );
  OAI22_X1 U14949 ( .A1(n13049), .A2(n12828), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12822), .ZN(n12823) );
  AOI21_X1 U14950 ( .B1(n13055), .B2(n12867), .A(n12823), .ZN(n12824) );
  OAI211_X1 U14951 ( .C1(n13219), .C2(n12829), .A(n12825), .B(n12824), .ZN(
        P2_U3201) );
  AND2_X1 U14952 ( .A1(n13154), .A2(n13152), .ZN(n12826) );
  AOI21_X1 U14953 ( .B1(n13079), .B2(n13153), .A(n12826), .ZN(n13111) );
  OAI22_X1 U14954 ( .A1(n12828), .A2(n13111), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12827), .ZN(n12831) );
  NOR2_X1 U14955 ( .A1(n13242), .A2(n12829), .ZN(n12830) );
  AOI211_X1 U14956 ( .C1(n12867), .C2(n13117), .A(n12831), .B(n12830), .ZN(
        n12839) );
  INV_X1 U14957 ( .A(n12832), .ZN(n12836) );
  OAI22_X1 U14958 ( .A1(n12834), .A2(n12858), .B1(n12833), .B2(n12872), .ZN(
        n12835) );
  NAND3_X1 U14959 ( .A1(n12837), .A2(n12836), .A3(n12835), .ZN(n12838) );
  OAI211_X1 U14960 ( .C1(n12840), .C2(n12858), .A(n12839), .B(n12838), .ZN(
        P2_U3205) );
  AOI22_X1 U14961 ( .A1(n12842), .A2(n12865), .B1(n12841), .B2(n12880), .ZN(
        n12853) );
  INV_X1 U14962 ( .A(n12843), .ZN(n12852) );
  INV_X1 U14963 ( .A(n12844), .ZN(n13088) );
  OAI22_X1 U14964 ( .A1(n12856), .A2(n13088), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12845), .ZN(n12850) );
  OAI22_X1 U14965 ( .A1(n12848), .A2(n12847), .B1(n12869), .B2(n12846), .ZN(
        n12849) );
  AOI211_X1 U14966 ( .C1(n13231), .C2(n12871), .A(n12850), .B(n12849), .ZN(
        n12851) );
  OAI21_X1 U14967 ( .B1(n12853), .B2(n12852), .A(n12851), .ZN(P2_U3207) );
  INV_X1 U14968 ( .A(n12869), .ZN(n12854) );
  AOI22_X1 U14969 ( .A1(n12854), .A2(n13154), .B1(n12875), .B2(n13151), .ZN(
        n12855) );
  NAND2_X1 U14970 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14729)
         );
  OAI211_X1 U14971 ( .C1(n12856), .C2(n13159), .A(n12855), .B(n14729), .ZN(
        n12862) );
  AOI211_X1 U14972 ( .C1(n12860), .C2(n12859), .A(n12858), .B(n12857), .ZN(
        n12861) );
  AOI211_X1 U14973 ( .C1(n13253), .C2(n12871), .A(n12862), .B(n12861), .ZN(
        n12863) );
  INV_X1 U14974 ( .A(n12863), .ZN(P2_U3210) );
  OAI21_X1 U14975 ( .B1(n12874), .B2(n12811), .A(n12864), .ZN(n12866) );
  NAND2_X1 U14976 ( .A1(n12866), .A2(n12865), .ZN(n12879) );
  AOI22_X1 U14977 ( .A1(n12867), .A2(n13025), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12868) );
  OAI21_X1 U14978 ( .B1(n12958), .B2(n12869), .A(n12868), .ZN(n12870) );
  AOI21_X1 U14979 ( .B1(n13209), .B2(n12871), .A(n12870), .ZN(n12878) );
  NOR3_X1 U14980 ( .A1(n12874), .A2(n12873), .A3(n12872), .ZN(n12876) );
  OAI21_X1 U14981 ( .B1(n12876), .B2(n12875), .A(n13017), .ZN(n12877) );
  NAND3_X1 U14982 ( .A1(n12879), .A2(n12878), .A3(n12877), .ZN(P2_U3212) );
  MUX2_X1 U14983 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n12950), .S(n6451), .Z(
        P2_U3562) );
  MUX2_X1 U14984 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n12975), .S(n6451), .Z(
        P2_U3561) );
  MUX2_X1 U14985 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n12989), .S(n6451), .Z(
        P2_U3560) );
  MUX2_X1 U14986 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n12961), .S(n6451), .Z(
        P2_U3559) );
  MUX2_X1 U14987 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13018), .S(n6451), .Z(
        P2_U3558) );
  MUX2_X1 U14988 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13035), .S(n6451), .Z(
        P2_U3557) );
  MUX2_X1 U14989 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13017), .S(n6451), .Z(
        P2_U3556) );
  MUX2_X1 U14990 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13036), .S(n6451), .Z(
        P2_U3555) );
  MUX2_X1 U14991 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13080), .S(n6451), .Z(
        P2_U3554) );
  MUX2_X1 U14992 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n12880), .S(n6451), .Z(
        P2_U3553) );
  MUX2_X1 U14993 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13079), .S(n6451), .Z(
        P2_U3552) );
  MUX2_X1 U14994 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n12881), .S(n6451), .Z(
        P2_U3551) );
  MUX2_X1 U14995 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13154), .S(n6451), .Z(
        P2_U3550) );
  MUX2_X1 U14996 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n12882), .S(n6451), .Z(
        P2_U3549) );
  MUX2_X1 U14997 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13151), .S(n6451), .Z(
        P2_U3548) );
  MUX2_X1 U14998 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n12883), .S(n6451), .Z(
        P2_U3547) );
  MUX2_X1 U14999 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n12884), .S(n6451), .Z(
        P2_U3546) );
  MUX2_X1 U15000 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n12885), .S(n6451), .Z(
        P2_U3545) );
  MUX2_X1 U15001 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n12886), .S(n6451), .Z(
        P2_U3544) );
  MUX2_X1 U15002 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n12887), .S(n6451), .Z(
        P2_U3543) );
  MUX2_X1 U15003 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n12888), .S(n6451), .Z(
        P2_U3542) );
  MUX2_X1 U15004 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n12889), .S(n6451), .Z(
        P2_U3541) );
  MUX2_X1 U15005 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n12890), .S(n6451), .Z(
        P2_U3540) );
  MUX2_X1 U15006 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n12891), .S(n6451), .Z(
        P2_U3539) );
  MUX2_X1 U15007 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n12892), .S(n6451), .Z(
        P2_U3538) );
  MUX2_X1 U15008 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n12893), .S(n6451), .Z(
        P2_U3537) );
  MUX2_X1 U15009 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n12894), .S(n6451), .Z(
        P2_U3536) );
  MUX2_X1 U15010 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n12895), .S(n6451), .Z(
        P2_U3535) );
  MUX2_X1 U15011 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n12896), .S(n6451), .Z(
        P2_U3534) );
  MUX2_X1 U15012 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n12897), .S(n6451), .Z(
        P2_U3533) );
  MUX2_X1 U15013 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n12898), .S(n6451), .Z(
        P2_U3532) );
  MUX2_X1 U15014 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n12899), .S(n6451), .Z(
        P2_U3531) );
  INV_X1 U15015 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n12901) );
  OAI21_X1 U15016 ( .B1(n14731), .B2(n12901), .A(n12900), .ZN(n12902) );
  AOI21_X1 U15017 ( .B1(n12903), .B2(n14728), .A(n12902), .ZN(n12913) );
  OAI21_X1 U15018 ( .B1(n12906), .B2(n12905), .A(n12904), .ZN(n12907) );
  NAND2_X1 U15019 ( .A1(n12907), .A2(n14724), .ZN(n12912) );
  OAI211_X1 U15020 ( .C1(n12910), .C2(n12909), .A(n12908), .B(n14657), .ZN(
        n12911) );
  NAND3_X1 U15021 ( .A1(n12913), .A2(n12912), .A3(n12911), .ZN(P2_U3225) );
  INV_X1 U15022 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n12914) );
  NAND2_X1 U15023 ( .A1(n12928), .A2(n12914), .ZN(n12915) );
  NAND2_X1 U15024 ( .A1(n12916), .A2(n12915), .ZN(n14651) );
  NAND2_X1 U15025 ( .A1(n12931), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n12917) );
  OAI21_X1 U15026 ( .B1(n12931), .B2(P2_REG2_REG_13__SCAN_IN), .A(n12917), 
        .ZN(n14650) );
  NOR2_X1 U15027 ( .A1(n14651), .A2(n14650), .ZN(n14654) );
  AOI21_X1 U15028 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n12931), .A(n14654), 
        .ZN(n12918) );
  NOR2_X1 U15029 ( .A1(n12918), .A2(n12919), .ZN(n12920) );
  INV_X1 U15030 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n15134) );
  XNOR2_X1 U15031 ( .A(n12919), .B(n12918), .ZN(n14669) );
  NOR2_X1 U15032 ( .A1(n15134), .A2(n14669), .ZN(n14668) );
  NOR2_X1 U15033 ( .A1(n12920), .A2(n14668), .ZN(n12921) );
  NOR2_X1 U15034 ( .A1(n12921), .A2(n14678), .ZN(n12922) );
  INV_X1 U15035 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n14683) );
  XNOR2_X1 U15036 ( .A(n12921), .B(n14678), .ZN(n14684) );
  NOR2_X1 U15037 ( .A1(n14683), .A2(n14684), .ZN(n14682) );
  NOR2_X1 U15038 ( .A1(n12922), .A2(n14682), .ZN(n14696) );
  NAND2_X1 U15039 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n14699), .ZN(n12923) );
  OAI21_X1 U15040 ( .B1(n14699), .B2(P2_REG2_REG_16__SCAN_IN), .A(n12923), 
        .ZN(n14695) );
  NOR2_X1 U15041 ( .A1(n14696), .A2(n14695), .ZN(n14694) );
  AOI21_X1 U15042 ( .B1(n14699), .B2(P2_REG2_REG_16__SCAN_IN), .A(n14694), 
        .ZN(n14709) );
  NAND2_X1 U15043 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n14712), .ZN(n12924) );
  OAI21_X1 U15044 ( .B1(n14712), .B2(P2_REG2_REG_17__SCAN_IN), .A(n12924), 
        .ZN(n14708) );
  NOR2_X1 U15045 ( .A1(n14709), .A2(n14708), .ZN(n14707) );
  AOI21_X1 U15046 ( .B1(n14712), .B2(P2_REG2_REG_17__SCAN_IN), .A(n14707), 
        .ZN(n12925) );
  XNOR2_X1 U15047 ( .A(n14727), .B(n12925), .ZN(n14722) );
  INV_X1 U15048 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n14721) );
  NAND2_X1 U15049 ( .A1(n14722), .A2(n14721), .ZN(n14720) );
  NAND2_X1 U15050 ( .A1(n12925), .A2(n12935), .ZN(n12926) );
  NAND2_X1 U15051 ( .A1(n14720), .A2(n12926), .ZN(n12927) );
  INV_X1 U15052 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n15070) );
  XOR2_X1 U15053 ( .A(n12927), .B(n15070), .Z(n12939) );
  INV_X1 U15054 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n12938) );
  NAND2_X1 U15055 ( .A1(n12928), .A2(n15147), .ZN(n12929) );
  NAND2_X1 U15056 ( .A1(n12930), .A2(n12929), .ZN(n14656) );
  XNOR2_X1 U15057 ( .A(n12931), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n14655) );
  NOR2_X1 U15058 ( .A1(n14656), .A2(n14655), .ZN(n14662) );
  AOI21_X1 U15059 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n12931), .A(n14662), 
        .ZN(n14672) );
  XNOR2_X1 U15060 ( .A(n14675), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n14671) );
  NOR2_X1 U15061 ( .A1(n14672), .A2(n14671), .ZN(n14670) );
  AOI21_X1 U15062 ( .B1(n14675), .B2(P2_REG1_REG_14__SCAN_IN), .A(n14670), 
        .ZN(n12932) );
  NOR2_X1 U15063 ( .A1(n12932), .A2(n14678), .ZN(n12933) );
  INV_X1 U15064 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14680) );
  XNOR2_X1 U15065 ( .A(n14678), .B(n12932), .ZN(n14681) );
  NOR2_X1 U15066 ( .A1(n14680), .A2(n14681), .ZN(n14679) );
  NOR2_X1 U15067 ( .A1(n12933), .A2(n14679), .ZN(n14693) );
  XNOR2_X1 U15068 ( .A(n14699), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14692) );
  NOR2_X1 U15069 ( .A1(n14693), .A2(n14692), .ZN(n14691) );
  AOI21_X1 U15070 ( .B1(n14699), .B2(P2_REG1_REG_16__SCAN_IN), .A(n14691), 
        .ZN(n14705) );
  XNOR2_X1 U15071 ( .A(n14712), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14704) );
  NOR2_X1 U15072 ( .A1(n14705), .A2(n14704), .ZN(n14703) );
  AOI21_X1 U15073 ( .B1(n14712), .B2(P2_REG1_REG_17__SCAN_IN), .A(n14703), 
        .ZN(n12934) );
  NOR2_X1 U15074 ( .A1(n12934), .A2(n12935), .ZN(n12936) );
  INV_X1 U15075 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14718) );
  XNOR2_X1 U15076 ( .A(n12935), .B(n12934), .ZN(n14719) );
  NOR2_X1 U15077 ( .A1(n14718), .A2(n14719), .ZN(n14717) );
  NOR2_X1 U15078 ( .A1(n12936), .A2(n14717), .ZN(n12937) );
  XOR2_X1 U15079 ( .A(n12938), .B(n12937), .Z(n12942) );
  AOI22_X1 U15080 ( .A1(n12939), .A2(n14724), .B1(n14657), .B2(n12942), .ZN(
        n12945) );
  INV_X1 U15081 ( .A(n12939), .ZN(n12940) );
  AOI21_X1 U15082 ( .B1(n14724), .B2(n12940), .A(n14728), .ZN(n12941) );
  OAI21_X1 U15083 ( .B1(n12942), .B2(n14716), .A(n12941), .ZN(n12943) );
  INV_X1 U15084 ( .A(n12943), .ZN(n12944) );
  MUX2_X1 U15085 ( .A(n12945), .B(n12944), .S(n12997), .Z(n12947) );
  OAI211_X1 U15086 ( .C1(n12948), .C2(n14731), .A(n12947), .B(n12946), .ZN(
        P2_U3233) );
  NAND2_X1 U15087 ( .A1(n12963), .A2(n9487), .ZN(n12954) );
  XNOR2_X1 U15088 ( .A(n12954), .B(n13188), .ZN(n13191) );
  NAND2_X1 U15089 ( .A1(n12949), .A2(P2_B_REG_SCAN_IN), .ZN(n12974) );
  NAND3_X1 U15090 ( .A1(n13153), .A2(n12950), .A3(n12974), .ZN(n13192) );
  NOR2_X1 U15091 ( .A1(n13187), .A2(n13192), .ZN(n12956) );
  AOI21_X1 U15092 ( .B1(n13187), .B2(P2_REG2_REG_31__SCAN_IN), .A(n12956), 
        .ZN(n12952) );
  NAND2_X1 U15093 ( .A1(n13188), .A2(n13143), .ZN(n12951) );
  OAI211_X1 U15094 ( .C1(n13191), .C2(n12953), .A(n12952), .B(n12951), .ZN(
        P2_U3234) );
  OAI211_X1 U15095 ( .C1(n12963), .C2(n9487), .A(n13136), .B(n12954), .ZN(
        n13193) );
  NOR2_X1 U15096 ( .A1(n9487), .A2(n13178), .ZN(n12955) );
  AOI211_X1 U15097 ( .C1(n13187), .C2(P2_REG2_REG_30__SCAN_IN), .A(n12956), 
        .B(n12955), .ZN(n12957) );
  OAI21_X1 U15098 ( .B1(n13140), .B2(n13193), .A(n12957), .ZN(P2_U3235) );
  OAI22_X2 U15099 ( .A1(n12960), .A2(n12959), .B1(n13007), .B2(n12958), .ZN(
        n12983) );
  AOI22_X1 U15100 ( .A1(n12983), .A2(n12984), .B1(n12995), .B2(n12961), .ZN(
        n12962) );
  XNOR2_X1 U15101 ( .A(n12962), .B(n12970), .ZN(n13198) );
  AOI211_X1 U15102 ( .C1(n12964), .C2(n12993), .A(n13190), .B(n12963), .ZN(
        n13195) );
  INV_X1 U15103 ( .A(n12965), .ZN(n12966) );
  AOI22_X1 U15104 ( .A1(n12966), .A2(n13175), .B1(n13187), .B2(
        P2_REG2_REG_29__SCAN_IN), .ZN(n12967) );
  OAI21_X1 U15105 ( .B1(n13196), .B2(n13178), .A(n12967), .ZN(n12968) );
  AOI21_X1 U15106 ( .B1(n13195), .B2(n13185), .A(n12968), .ZN(n12982) );
  NOR2_X1 U15107 ( .A1(n13007), .A2(n13018), .ZN(n12985) );
  NAND2_X1 U15108 ( .A1(n12987), .A2(n12969), .ZN(n12972) );
  XNOR2_X1 U15109 ( .A(n12972), .B(n12971), .ZN(n12973) );
  NAND3_X1 U15110 ( .A1(n13153), .A2(n12975), .A3(n12974), .ZN(n12976) );
  OAI21_X1 U15111 ( .B1(n12977), .B2(n13067), .A(n12976), .ZN(n12978) );
  INV_X1 U15112 ( .A(n12978), .ZN(n12979) );
  NAND2_X1 U15113 ( .A1(n13194), .A2(n13135), .ZN(n12981) );
  OAI211_X1 U15114 ( .C1(n13198), .C2(n13182), .A(n12982), .B(n12981), .ZN(
        P2_U3236) );
  XNOR2_X1 U15115 ( .A(n12983), .B(n12984), .ZN(n13201) );
  AOI22_X1 U15116 ( .A1(n12995), .A2(n13143), .B1(n13187), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n13001) );
  OAI21_X1 U15117 ( .B1(n12986), .B2(n12985), .A(n12984), .ZN(n12988) );
  NAND3_X1 U15118 ( .A1(n12988), .A2(n13169), .A3(n12987), .ZN(n12991) );
  AOI22_X1 U15119 ( .A1(n13153), .A2(n12989), .B1(n13018), .B2(n13152), .ZN(
        n12990) );
  NAND2_X1 U15120 ( .A1(n12991), .A2(n12990), .ZN(n13199) );
  INV_X1 U15121 ( .A(n12993), .ZN(n12994) );
  AOI211_X1 U15122 ( .C1(n12995), .C2(n6826), .A(n13190), .B(n12994), .ZN(
        n13200) );
  INV_X1 U15123 ( .A(n13200), .ZN(n12998) );
  OAI22_X1 U15124 ( .A1(n12998), .A2(n12997), .B1(n13133), .B2(n12996), .ZN(
        n12999) );
  OAI21_X1 U15125 ( .B1(n13199), .B2(n12999), .A(n13135), .ZN(n13000) );
  OAI211_X1 U15126 ( .C1(n13201), .C2(n13182), .A(n13001), .B(n13000), .ZN(
        P2_U3237) );
  NAND2_X1 U15127 ( .A1(n13002), .A2(n13185), .ZN(n13006) );
  INV_X1 U15128 ( .A(n13003), .ZN(n13004) );
  AOI22_X1 U15129 ( .A1(n13187), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n13004), 
        .B2(n13175), .ZN(n13005) );
  OAI211_X1 U15130 ( .C1(n13007), .C2(n13178), .A(n13006), .B(n13005), .ZN(
        n13008) );
  AOI21_X1 U15131 ( .B1(n13009), .B2(n13135), .A(n13008), .ZN(n13010) );
  OAI21_X1 U15132 ( .B1(n13182), .B2(n13011), .A(n13010), .ZN(P2_U3238) );
  XNOR2_X1 U15133 ( .A(n13013), .B(n13012), .ZN(n13211) );
  NAND2_X1 U15134 ( .A1(n13014), .A2(n13169), .ZN(n13021) );
  AOI21_X1 U15135 ( .B1(n13032), .B2(n13016), .A(n13015), .ZN(n13020) );
  AOI22_X1 U15136 ( .A1(n13018), .A2(n13153), .B1(n13152), .B2(n13017), .ZN(
        n13019) );
  OAI21_X1 U15137 ( .B1(n13021), .B2(n13020), .A(n13019), .ZN(n13207) );
  INV_X1 U15138 ( .A(n13040), .ZN(n13024) );
  INV_X1 U15139 ( .A(n13022), .ZN(n13023) );
  AOI211_X1 U15140 ( .C1(n13209), .C2(n13024), .A(n13190), .B(n13023), .ZN(
        n13208) );
  NAND2_X1 U15141 ( .A1(n13208), .A2(n13185), .ZN(n13027) );
  AOI22_X1 U15142 ( .A1(n13187), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n13025), 
        .B2(n13175), .ZN(n13026) );
  OAI211_X1 U15143 ( .C1(n13028), .C2(n13178), .A(n13027), .B(n13026), .ZN(
        n13029) );
  AOI21_X1 U15144 ( .B1(n13207), .B2(n13135), .A(n13029), .ZN(n13030) );
  OAI21_X1 U15145 ( .B1(n13211), .B2(n13182), .A(n13030), .ZN(P2_U3239) );
  XNOR2_X1 U15146 ( .A(n13031), .B(n13033), .ZN(n13217) );
  OAI21_X1 U15147 ( .B1(n13034), .B2(n13033), .A(n13032), .ZN(n13037) );
  AOI222_X1 U15148 ( .A1(n13169), .A2(n13037), .B1(n13036), .B2(n13152), .C1(
        n13035), .C2(n13153), .ZN(n13216) );
  INV_X1 U15149 ( .A(n13216), .ZN(n13046) );
  NOR2_X1 U15150 ( .A1(n13054), .A2(n13038), .ZN(n13039) );
  OR3_X1 U15151 ( .A1(n13040), .A2(n13039), .A3(n13190), .ZN(n13212) );
  INV_X1 U15152 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13042) );
  OAI22_X1 U15153 ( .A1(n13135), .A2(n13042), .B1(n13041), .B2(n13133), .ZN(
        n13043) );
  AOI21_X1 U15154 ( .B1(n13214), .B2(n13143), .A(n13043), .ZN(n13044) );
  OAI21_X1 U15155 ( .B1(n13212), .B2(n13140), .A(n13044), .ZN(n13045) );
  AOI21_X1 U15156 ( .B1(n13046), .B2(n13135), .A(n13045), .ZN(n13047) );
  OAI21_X1 U15157 ( .B1(n13182), .B2(n13217), .A(n13047), .ZN(P2_U3240) );
  XNOR2_X1 U15158 ( .A(n13048), .B(n13052), .ZN(n13050) );
  OAI21_X1 U15159 ( .B1(n13050), .B2(n13064), .A(n13049), .ZN(n13220) );
  INV_X1 U15160 ( .A(n13220), .ZN(n13060) );
  AOI21_X1 U15161 ( .B1(n13052), .B2(n13051), .A(n6537), .ZN(n13222) );
  NOR2_X1 U15162 ( .A1(n13070), .A2(n13219), .ZN(n13053) );
  OR3_X1 U15163 ( .A1(n13054), .A2(n13053), .A3(n13190), .ZN(n13218) );
  NOR2_X1 U15164 ( .A1(n13218), .A2(n13140), .ZN(n13058) );
  AOI22_X1 U15165 ( .A1(n13187), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13055), 
        .B2(n13175), .ZN(n13056) );
  OAI21_X1 U15166 ( .B1(n13219), .B2(n13178), .A(n13056), .ZN(n13057) );
  AOI211_X1 U15167 ( .C1(n13222), .C2(n13122), .A(n13058), .B(n13057), .ZN(
        n13059) );
  OAI21_X1 U15168 ( .B1(n13187), .B2(n13060), .A(n13059), .ZN(P2_U3241) );
  XNOR2_X1 U15169 ( .A(n13061), .B(n13062), .ZN(n13228) );
  XNOR2_X1 U15170 ( .A(n13063), .B(n13062), .ZN(n13065) );
  OAI222_X1 U15171 ( .A1(n13069), .A2(n13068), .B1(n13067), .B2(n13066), .C1(
        n13065), .C2(n13064), .ZN(n13224) );
  NAND2_X1 U15172 ( .A1(n13224), .A2(n13135), .ZN(n13077) );
  INV_X1 U15173 ( .A(n13087), .ZN(n13071) );
  AOI211_X1 U15174 ( .C1(n13226), .C2(n13071), .A(n13190), .B(n13070), .ZN(
        n13225) );
  AOI22_X1 U15175 ( .A1(n13187), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n13072), 
        .B2(n13175), .ZN(n13073) );
  OAI21_X1 U15176 ( .B1(n13074), .B2(n13178), .A(n13073), .ZN(n13075) );
  AOI21_X1 U15177 ( .B1(n13225), .B2(n13185), .A(n13075), .ZN(n13076) );
  OAI211_X1 U15178 ( .C1(n13182), .C2(n13228), .A(n13077), .B(n13076), .ZN(
        P2_U3242) );
  XNOR2_X1 U15179 ( .A(n13078), .B(n13083), .ZN(n13081) );
  AOI222_X1 U15180 ( .A1(n13169), .A2(n13081), .B1(n13080), .B2(n13153), .C1(
        n13079), .C2(n13152), .ZN(n13233) );
  OAI21_X1 U15181 ( .B1(n13084), .B2(n13083), .A(n13082), .ZN(n13234) );
  INV_X1 U15182 ( .A(n13234), .ZN(n13093) );
  NOR2_X1 U15183 ( .A1(n13085), .A2(n13098), .ZN(n13086) );
  INV_X1 U15184 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13089) );
  OAI22_X1 U15185 ( .A1(n13135), .A2(n13089), .B1(n13088), .B2(n13133), .ZN(
        n13090) );
  AOI21_X1 U15186 ( .B1(n13231), .B2(n13143), .A(n13090), .ZN(n13091) );
  OAI21_X1 U15187 ( .B1(n13229), .B2(n13140), .A(n13091), .ZN(n13092) );
  AOI21_X1 U15188 ( .B1(n13093), .B2(n13122), .A(n13092), .ZN(n13094) );
  OAI21_X1 U15189 ( .B1(n13233), .B2(n13187), .A(n13094), .ZN(P2_U3243) );
  XNOR2_X1 U15190 ( .A(n13095), .B(n13104), .ZN(n13097) );
  AOI21_X1 U15191 ( .B1(n13097), .B2(n13169), .A(n13096), .ZN(n13238) );
  INV_X1 U15192 ( .A(n13115), .ZN(n13099) );
  AOI211_X1 U15193 ( .C1(n13236), .C2(n13099), .A(n13190), .B(n13098), .ZN(
        n13235) );
  INV_X1 U15194 ( .A(n13100), .ZN(n13101) );
  AOI22_X1 U15195 ( .A1(n13187), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13101), 
        .B2(n13175), .ZN(n13102) );
  OAI21_X1 U15196 ( .B1(n13103), .B2(n13178), .A(n13102), .ZN(n13107) );
  XOR2_X1 U15197 ( .A(n13105), .B(n13104), .Z(n13239) );
  NOR2_X1 U15198 ( .A1(n13239), .A2(n13182), .ZN(n13106) );
  AOI211_X1 U15199 ( .C1(n13235), .C2(n13185), .A(n13107), .B(n13106), .ZN(
        n13108) );
  OAI21_X1 U15200 ( .B1(n13187), .B2(n13238), .A(n13108), .ZN(P2_U3244) );
  XNOR2_X1 U15201 ( .A(n13109), .B(n13113), .ZN(n13110) );
  NAND2_X1 U15202 ( .A1(n13110), .A2(n13169), .ZN(n13112) );
  NAND2_X1 U15203 ( .A1(n13112), .A2(n13111), .ZN(n13245) );
  INV_X1 U15204 ( .A(n13245), .ZN(n13124) );
  XNOR2_X1 U15205 ( .A(n13114), .B(n13113), .ZN(n13240) );
  OAI21_X1 U15206 ( .B1(n13139), .B2(n13242), .A(n13136), .ZN(n13116) );
  OR2_X1 U15207 ( .A1(n13116), .A2(n13115), .ZN(n13241) );
  AOI22_X1 U15208 ( .A1(n13187), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13117), 
        .B2(n13175), .ZN(n13120) );
  NAND2_X1 U15209 ( .A1(n13118), .A2(n13143), .ZN(n13119) );
  OAI211_X1 U15210 ( .C1(n13241), .C2(n13140), .A(n13120), .B(n13119), .ZN(
        n13121) );
  AOI21_X1 U15211 ( .B1(n13240), .B2(n13122), .A(n13121), .ZN(n13123) );
  OAI21_X1 U15212 ( .B1(n13124), .B2(n13187), .A(n13123), .ZN(P2_U3245) );
  XNOR2_X1 U15213 ( .A(n13125), .B(n13126), .ZN(n13249) );
  INV_X1 U15214 ( .A(n13126), .ZN(n13127) );
  XNOR2_X1 U15215 ( .A(n13128), .B(n13127), .ZN(n13129) );
  NAND2_X1 U15216 ( .A1(n13129), .A2(n13169), .ZN(n13132) );
  INV_X1 U15217 ( .A(n13130), .ZN(n13131) );
  NAND2_X1 U15218 ( .A1(n13132), .A2(n13131), .ZN(n13250) );
  NAND2_X1 U15219 ( .A1(n13250), .A2(n13135), .ZN(n13145) );
  OAI22_X1 U15220 ( .A1(n13135), .A2(n15070), .B1(n13134), .B2(n13133), .ZN(
        n13142) );
  NAND2_X1 U15221 ( .A1(n13158), .A2(n13246), .ZN(n13137) );
  NAND2_X1 U15222 ( .A1(n13137), .A2(n13136), .ZN(n13138) );
  OR2_X1 U15223 ( .A1(n13139), .A2(n13138), .ZN(n13248) );
  NOR2_X1 U15224 ( .A1(n13248), .A2(n13140), .ZN(n13141) );
  AOI211_X1 U15225 ( .C1(n13143), .C2(n13246), .A(n13142), .B(n13141), .ZN(
        n13144) );
  OAI211_X1 U15226 ( .C1(n13182), .C2(n13249), .A(n13145), .B(n13144), .ZN(
        P2_U3246) );
  XOR2_X1 U15227 ( .A(n13146), .B(n13150), .Z(n13157) );
  INV_X1 U15228 ( .A(n13147), .ZN(n13148) );
  AOI21_X1 U15229 ( .B1(n13150), .B2(n13149), .A(n13148), .ZN(n13256) );
  AOI22_X1 U15230 ( .A1(n13154), .A2(n13153), .B1(n13152), .B2(n13151), .ZN(
        n13155) );
  OAI21_X1 U15231 ( .B1(n13256), .B2(n14839), .A(n13155), .ZN(n13156) );
  AOI21_X1 U15232 ( .B1(n13157), .B2(n13169), .A(n13156), .ZN(n13255) );
  AOI211_X1 U15233 ( .C1(n13253), .C2(n13172), .A(n13190), .B(n6829), .ZN(
        n13252) );
  INV_X1 U15234 ( .A(n13253), .ZN(n13162) );
  INV_X1 U15235 ( .A(n13159), .ZN(n13160) );
  AOI22_X1 U15236 ( .A1(n13187), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13160), 
        .B2(n13175), .ZN(n13161) );
  OAI21_X1 U15237 ( .B1(n13162), .B2(n13178), .A(n13161), .ZN(n13165) );
  NOR2_X1 U15238 ( .A1(n13256), .A2(n13163), .ZN(n13164) );
  AOI211_X1 U15239 ( .C1(n13252), .C2(n13185), .A(n13165), .B(n13164), .ZN(
        n13166) );
  OAI21_X1 U15240 ( .B1(n13187), .B2(n13255), .A(n13166), .ZN(P2_U3247) );
  XNOR2_X1 U15241 ( .A(n13167), .B(n13180), .ZN(n13170) );
  AOI21_X1 U15242 ( .B1(n13170), .B2(n13169), .A(n13168), .ZN(n13260) );
  INV_X1 U15243 ( .A(n13171), .ZN(n13174) );
  INV_X1 U15244 ( .A(n13172), .ZN(n13173) );
  AOI211_X1 U15245 ( .C1(n13258), .C2(n13174), .A(n13190), .B(n13173), .ZN(
        n13257) );
  AOI22_X1 U15246 ( .A1(n13187), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13176), 
        .B2(n13175), .ZN(n13177) );
  OAI21_X1 U15247 ( .B1(n13179), .B2(n13178), .A(n13177), .ZN(n13184) );
  XNOR2_X1 U15248 ( .A(n13181), .B(n13180), .ZN(n13261) );
  NOR2_X1 U15249 ( .A1(n13261), .A2(n13182), .ZN(n13183) );
  AOI211_X1 U15250 ( .C1(n13257), .C2(n13185), .A(n13184), .B(n13183), .ZN(
        n13186) );
  OAI21_X1 U15251 ( .B1(n13187), .B2(n13260), .A(n13186), .ZN(P2_U3248) );
  NAND2_X1 U15252 ( .A1(n13188), .A2(n14841), .ZN(n13189) );
  OAI211_X1 U15253 ( .C1(n13191), .C2(n13190), .A(n13192), .B(n13189), .ZN(
        n13278) );
  MUX2_X1 U15254 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13278), .S(n14876), .Z(
        P2_U3530) );
  OAI211_X1 U15255 ( .C1(n9487), .C2(n14852), .A(n13193), .B(n13192), .ZN(
        n13279) );
  MUX2_X1 U15256 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13279), .S(n14876), .Z(
        P2_U3529) );
  MUX2_X1 U15257 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13280), .S(n14876), .Z(
        P2_U3528) );
  INV_X1 U15258 ( .A(n13199), .ZN(n13205) );
  NAND2_X1 U15259 ( .A1(n12995), .A2(n14841), .ZN(n13203) );
  NAND4_X1 U15260 ( .A1(n13205), .A2(n12998), .A3(n13204), .A4(n13203), .ZN(
        n13281) );
  MUX2_X1 U15261 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13281), .S(n14876), .Z(
        P2_U3527) );
  MUX2_X1 U15262 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13206), .S(n14876), .Z(
        P2_U3526) );
  AOI211_X1 U15263 ( .C1(n14841), .C2(n13209), .A(n13208), .B(n13207), .ZN(
        n13210) );
  OAI21_X1 U15264 ( .B1(n14798), .B2(n13211), .A(n13210), .ZN(n13282) );
  MUX2_X1 U15265 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13282), .S(n14876), .Z(
        P2_U3525) );
  INV_X1 U15266 ( .A(n13212), .ZN(n13213) );
  AOI21_X1 U15267 ( .B1(n14841), .B2(n13214), .A(n13213), .ZN(n13215) );
  OAI211_X1 U15268 ( .C1(n14798), .C2(n13217), .A(n13216), .B(n13215), .ZN(
        n13283) );
  MUX2_X1 U15269 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13283), .S(n14876), .Z(
        P2_U3524) );
  OAI21_X1 U15270 ( .B1(n13219), .B2(n14852), .A(n13218), .ZN(n13221) );
  AOI211_X1 U15271 ( .C1(n13222), .C2(n8001), .A(n13221), .B(n13220), .ZN(
        n13223) );
  INV_X1 U15272 ( .A(n13223), .ZN(n13284) );
  MUX2_X1 U15273 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13284), .S(n14876), .Z(
        P2_U3523) );
  AOI211_X1 U15274 ( .C1(n14841), .C2(n13226), .A(n13225), .B(n13224), .ZN(
        n13227) );
  OAI21_X1 U15275 ( .B1(n14798), .B2(n13228), .A(n13227), .ZN(n13285) );
  MUX2_X1 U15276 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13285), .S(n14876), .Z(
        P2_U3522) );
  INV_X1 U15277 ( .A(n13229), .ZN(n13230) );
  AOI21_X1 U15278 ( .B1(n14841), .B2(n13231), .A(n13230), .ZN(n13232) );
  OAI211_X1 U15279 ( .C1(n14798), .C2(n13234), .A(n13233), .B(n13232), .ZN(
        n13286) );
  MUX2_X1 U15280 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13286), .S(n14876), .Z(
        P2_U3521) );
  AOI21_X1 U15281 ( .B1(n14841), .B2(n13236), .A(n13235), .ZN(n13237) );
  OAI211_X1 U15282 ( .C1(n13239), .C2(n14798), .A(n13238), .B(n13237), .ZN(
        n13287) );
  MUX2_X1 U15283 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13287), .S(n14876), .Z(
        P2_U3520) );
  AND2_X1 U15284 ( .A1(n13240), .A2(n8001), .ZN(n13244) );
  OAI21_X1 U15285 ( .B1(n13242), .B2(n14852), .A(n13241), .ZN(n13243) );
  MUX2_X1 U15286 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13288), .S(n14876), .Z(
        P2_U3519) );
  NAND2_X1 U15287 ( .A1(n13246), .A2(n14841), .ZN(n13247) );
  OAI211_X1 U15288 ( .C1(n13249), .C2(n14798), .A(n13248), .B(n13247), .ZN(
        n13251) );
  MUX2_X1 U15289 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13289), .S(n14876), .Z(
        P2_U3518) );
  AOI21_X1 U15290 ( .B1(n14841), .B2(n13253), .A(n13252), .ZN(n13254) );
  OAI211_X1 U15291 ( .C1(n13256), .C2(n14838), .A(n13255), .B(n13254), .ZN(
        n13290) );
  MUX2_X1 U15292 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13290), .S(n14876), .Z(
        P2_U3517) );
  AOI21_X1 U15293 ( .B1(n14841), .B2(n13258), .A(n13257), .ZN(n13259) );
  OAI211_X1 U15294 ( .C1(n14798), .C2(n13261), .A(n13260), .B(n13259), .ZN(
        n13291) );
  MUX2_X1 U15295 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13291), .S(n14876), .Z(
        P2_U3516) );
  NAND2_X1 U15296 ( .A1(n13262), .A2(n14841), .ZN(n13263) );
  OAI211_X1 U15297 ( .C1(n13265), .C2(n14798), .A(n13264), .B(n13263), .ZN(
        n13266) );
  MUX2_X1 U15298 ( .A(n13292), .B(P2_REG1_REG_16__SCAN_IN), .S(n14873), .Z(
        P2_U3515) );
  AOI21_X1 U15299 ( .B1(n14841), .B2(n13269), .A(n13268), .ZN(n13270) );
  OAI211_X1 U15300 ( .C1(n14798), .C2(n13272), .A(n13271), .B(n13270), .ZN(
        n13293) );
  MUX2_X1 U15301 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13293), .S(n14876), .Z(
        P2_U3514) );
  AOI22_X1 U15302 ( .A1(n13274), .A2(n9578), .B1(n14841), .B2(n13273), .ZN(
        n13275) );
  OAI211_X1 U15303 ( .C1(n13277), .C2(n14838), .A(n13276), .B(n13275), .ZN(
        n13294) );
  MUX2_X1 U15304 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n13294), .S(n14876), .Z(
        P2_U3511) );
  MUX2_X1 U15305 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13278), .S(n14858), .Z(
        P2_U3498) );
  MUX2_X1 U15306 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13279), .S(n14858), .Z(
        P2_U3497) );
  MUX2_X1 U15307 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13281), .S(n14858), .Z(
        P2_U3495) );
  MUX2_X1 U15308 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13282), .S(n14858), .Z(
        P2_U3493) );
  MUX2_X1 U15309 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13283), .S(n14858), .Z(
        P2_U3492) );
  MUX2_X1 U15310 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13284), .S(n14858), .Z(
        P2_U3491) );
  MUX2_X1 U15311 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13285), .S(n14858), .Z(
        P2_U3490) );
  MUX2_X1 U15312 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13286), .S(n14858), .Z(
        P2_U3489) );
  MUX2_X1 U15313 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13287), .S(n14858), .Z(
        P2_U3488) );
  MUX2_X1 U15314 ( .A(n13288), .B(P2_REG0_REG_20__SCAN_IN), .S(n14856), .Z(
        P2_U3487) );
  MUX2_X1 U15315 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13289), .S(n14858), .Z(
        P2_U3486) );
  MUX2_X1 U15316 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13290), .S(n14858), .Z(
        P2_U3484) );
  MUX2_X1 U15317 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13291), .S(n14858), .Z(
        P2_U3481) );
  MUX2_X1 U15318 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13292), .S(n14858), .Z(
        P2_U3478) );
  MUX2_X1 U15319 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13293), .S(n14858), .Z(
        P2_U3475) );
  MUX2_X1 U15320 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n13294), .S(n14858), .Z(
        P2_U3466) );
  INV_X1 U15321 ( .A(n13295), .ZN(n14084) );
  NOR4_X1 U15322 ( .A1(n13297), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13296), .A4(
        P2_U3088), .ZN(n13298) );
  AOI21_X1 U15323 ( .B1(n13299), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13298), 
        .ZN(n13300) );
  OAI21_X1 U15324 ( .B1(n14084), .B2(n6452), .A(n13300), .ZN(P2_U3296) );
  OAI222_X1 U15325 ( .A1(n6452), .A2(n13303), .B1(P2_U3088), .B2(n13302), .C1(
        n13301), .C2(n13314), .ZN(P2_U3297) );
  INV_X1 U15326 ( .A(n9470), .ZN(n14087) );
  OAI222_X1 U15327 ( .A1(n6452), .A2(n14087), .B1(P2_U3088), .B2(n13305), .C1(
        n13304), .C2(n13314), .ZN(P2_U3298) );
  NAND2_X1 U15328 ( .A1(n13307), .A2(n13306), .ZN(n13309) );
  OAI211_X1 U15329 ( .C1(n13314), .C2(n13310), .A(n13309), .B(n13308), .ZN(
        P2_U3299) );
  OAI222_X1 U15330 ( .A1(n13314), .A2(n13313), .B1(n6452), .B2(n13312), .C1(
        n13311), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U15331 ( .A(n13315), .ZN(n13316) );
  MUX2_X1 U15332 ( .A(n13316), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI22_X1 U15333 ( .A1(n14052), .A2(n10594), .B1(n13755), .B2(n6486), .ZN(
        n13317) );
  XNOR2_X1 U15334 ( .A(n13317), .B(n13463), .ZN(n13321) );
  OR2_X1 U15335 ( .A1(n14052), .A2(n6486), .ZN(n13319) );
  NAND2_X1 U15336 ( .A1(n13790), .A2(n10598), .ZN(n13318) );
  NAND2_X1 U15337 ( .A1(n13319), .A2(n13318), .ZN(n13320) );
  NOR2_X1 U15338 ( .A1(n13321), .A2(n13320), .ZN(n13460) );
  AOI21_X1 U15339 ( .B1(n13321), .B2(n13320), .A(n13460), .ZN(n13423) );
  INV_X1 U15340 ( .A(n13322), .ZN(n13323) );
  NAND2_X1 U15341 ( .A1(n13324), .A2(n13323), .ZN(n13325) );
  NAND2_X1 U15342 ( .A1(n13326), .A2(n13325), .ZN(n14329) );
  INV_X1 U15343 ( .A(n14329), .ZN(n13333) );
  NAND2_X1 U15344 ( .A1(n14336), .A2(n13465), .ZN(n13328) );
  OR2_X1 U15345 ( .A1(n13330), .A2(n6486), .ZN(n13327) );
  NAND2_X1 U15346 ( .A1(n13328), .A2(n13327), .ZN(n13329) );
  XNOR2_X1 U15347 ( .A(n13329), .B(n13404), .ZN(n13335) );
  NOR2_X1 U15348 ( .A1(n13330), .A2(n13360), .ZN(n13331) );
  AOI21_X1 U15349 ( .B1(n14336), .B2(n13462), .A(n13331), .ZN(n13334) );
  XNOR2_X1 U15350 ( .A(n13335), .B(n13334), .ZN(n14328) );
  NAND2_X1 U15351 ( .A1(n13335), .A2(n13334), .ZN(n13336) );
  NAND2_X1 U15352 ( .A1(n14332), .A2(n13336), .ZN(n13340) );
  AOI22_X1 U15353 ( .A1(n14362), .A2(n13465), .B1(n6449), .B2(n13587), .ZN(
        n13337) );
  XOR2_X1 U15354 ( .A(n13463), .B(n13337), .Z(n13338) );
  XNOR2_X1 U15355 ( .A(n13340), .B(n13338), .ZN(n13573) );
  OAI22_X1 U15356 ( .A1(n13581), .A2(n6486), .B1(n14324), .B2(n13360), .ZN(
        n13572) );
  NAND2_X1 U15357 ( .A1(n13573), .A2(n13572), .ZN(n13571) );
  INV_X1 U15358 ( .A(n13338), .ZN(n13339) );
  OR2_X1 U15359 ( .A1(n13340), .A2(n13339), .ZN(n13341) );
  OAI22_X1 U15360 ( .A1(n14355), .A2(n10594), .B1(n13947), .B2(n6486), .ZN(
        n13342) );
  XNOR2_X1 U15361 ( .A(n13342), .B(n13463), .ZN(n13343) );
  OAI22_X1 U15362 ( .A1(n14355), .A2(n6486), .B1(n13947), .B2(n13360), .ZN(
        n13344) );
  XNOR2_X1 U15363 ( .A(n13343), .B(n13344), .ZN(n13506) );
  INV_X1 U15364 ( .A(n13343), .ZN(n13346) );
  INV_X1 U15365 ( .A(n13344), .ZN(n13345) );
  AOI22_X1 U15366 ( .A1(n14034), .A2(n13465), .B1(n13462), .B2(n13928), .ZN(
        n13347) );
  XOR2_X1 U15367 ( .A(n13463), .B(n13347), .Z(n13515) );
  AOI22_X1 U15368 ( .A1(n14034), .A2(n6449), .B1(n10598), .B2(n13928), .ZN(
        n13514) );
  NAND2_X1 U15369 ( .A1(n13348), .A2(n13514), .ZN(n13349) );
  AOI22_X1 U15370 ( .A1(n13936), .A2(n13462), .B1(n10598), .B2(n13912), .ZN(
        n13353) );
  AOI22_X1 U15371 ( .A1(n13936), .A2(n13465), .B1(n13462), .B2(n13912), .ZN(
        n13350) );
  XNOR2_X1 U15372 ( .A(n13350), .B(n13463), .ZN(n13354) );
  XOR2_X1 U15373 ( .A(n13353), .B(n13354), .Z(n13551) );
  NOR2_X1 U15374 ( .A1(n13553), .A2(n13360), .ZN(n13351) );
  AOI21_X1 U15375 ( .B1(n13917), .B2(n6449), .A(n13351), .ZN(n13356) );
  AOI22_X1 U15376 ( .A1(n13917), .A2(n13465), .B1(n6449), .B2(n13930), .ZN(
        n13352) );
  XNOR2_X1 U15377 ( .A(n13352), .B(n13463), .ZN(n13355) );
  XOR2_X1 U15378 ( .A(n13356), .B(n13355), .Z(n13454) );
  NAND2_X1 U15379 ( .A1(n13354), .A2(n13353), .ZN(n13452) );
  NAND2_X1 U15380 ( .A1(n13549), .A2(n7384), .ZN(n13453) );
  INV_X1 U15381 ( .A(n13355), .ZN(n13358) );
  INV_X1 U15382 ( .A(n13356), .ZN(n13357) );
  OAI22_X1 U15383 ( .A1(n14019), .A2(n6486), .B1(n13488), .B2(n13360), .ZN(
        n13362) );
  OAI22_X1 U15384 ( .A1(n14019), .A2(n10594), .B1(n13488), .B2(n6486), .ZN(
        n13361) );
  XNOR2_X1 U15385 ( .A(n13361), .B(n13463), .ZN(n13363) );
  XOR2_X1 U15386 ( .A(n13362), .B(n13363), .Z(n13530) );
  NAND2_X1 U15387 ( .A1(n13879), .A2(n13465), .ZN(n13366) );
  NAND2_X1 U15388 ( .A1(n13585), .A2(n6449), .ZN(n13365) );
  NAND2_X1 U15389 ( .A1(n13366), .A2(n13365), .ZN(n13367) );
  XNOR2_X1 U15390 ( .A(n13367), .B(n13463), .ZN(n13371) );
  NAND2_X1 U15391 ( .A1(n13879), .A2(n6449), .ZN(n13369) );
  NAND2_X1 U15392 ( .A1(n13585), .A2(n10598), .ZN(n13368) );
  NAND2_X1 U15393 ( .A1(n13369), .A2(n13368), .ZN(n13370) );
  NOR2_X1 U15394 ( .A1(n13371), .A2(n13370), .ZN(n13372) );
  AOI21_X1 U15395 ( .B1(n13371), .B2(n13370), .A(n13372), .ZN(n13483) );
  INV_X1 U15396 ( .A(n13372), .ZN(n13540) );
  NAND2_X1 U15397 ( .A1(n13863), .A2(n13465), .ZN(n13374) );
  NAND2_X1 U15398 ( .A1(n13487), .A2(n13462), .ZN(n13373) );
  NAND2_X1 U15399 ( .A1(n13374), .A2(n13373), .ZN(n13375) );
  XNOR2_X1 U15400 ( .A(n13375), .B(n13404), .ZN(n13377) );
  AND2_X1 U15401 ( .A1(n13487), .A2(n10598), .ZN(n13376) );
  AOI21_X1 U15402 ( .B1(n13863), .B2(n13462), .A(n13376), .ZN(n13378) );
  NAND2_X1 U15403 ( .A1(n13377), .A2(n13378), .ZN(n13382) );
  INV_X1 U15404 ( .A(n13377), .ZN(n13380) );
  INV_X1 U15405 ( .A(n13378), .ZN(n13379) );
  NAND2_X1 U15406 ( .A1(n13380), .A2(n13379), .ZN(n13381) );
  NAND2_X1 U15407 ( .A1(n13382), .A2(n13381), .ZN(n13539) );
  INV_X1 U15408 ( .A(n13382), .ZN(n13433) );
  NAND2_X1 U15409 ( .A1(n14001), .A2(n10578), .ZN(n13384) );
  NAND2_X1 U15410 ( .A1(n13856), .A2(n6449), .ZN(n13383) );
  NAND2_X1 U15411 ( .A1(n13384), .A2(n13383), .ZN(n13385) );
  XNOR2_X1 U15412 ( .A(n13385), .B(n13404), .ZN(n13387) );
  AND2_X1 U15413 ( .A1(n13856), .A2(n10598), .ZN(n13386) );
  AOI21_X1 U15414 ( .B1(n14001), .B2(n13462), .A(n13386), .ZN(n13388) );
  NAND2_X1 U15415 ( .A1(n13387), .A2(n13388), .ZN(n13524) );
  INV_X1 U15416 ( .A(n13387), .ZN(n13390) );
  INV_X1 U15417 ( .A(n13388), .ZN(n13389) );
  NAND2_X1 U15418 ( .A1(n13390), .A2(n13389), .ZN(n13391) );
  NAND2_X1 U15419 ( .A1(n13827), .A2(n13465), .ZN(n13393) );
  NAND2_X1 U15420 ( .A1(n13584), .A2(n13462), .ZN(n13392) );
  NAND2_X1 U15421 ( .A1(n13393), .A2(n13392), .ZN(n13394) );
  XNOR2_X1 U15422 ( .A(n13394), .B(n13404), .ZN(n13396) );
  AND2_X1 U15423 ( .A1(n13584), .A2(n10598), .ZN(n13395) );
  AOI21_X1 U15424 ( .B1(n13827), .B2(n6449), .A(n13395), .ZN(n13397) );
  NAND2_X1 U15425 ( .A1(n13396), .A2(n13397), .ZN(n13401) );
  INV_X1 U15426 ( .A(n13396), .ZN(n13399) );
  INV_X1 U15427 ( .A(n13397), .ZN(n13398) );
  NAND2_X1 U15428 ( .A1(n13399), .A2(n13398), .ZN(n13400) );
  NAND2_X1 U15429 ( .A1(n13401), .A2(n13400), .ZN(n13523) );
  INV_X1 U15430 ( .A(n13401), .ZN(n13497) );
  NAND2_X1 U15431 ( .A1(n13807), .A2(n10578), .ZN(n13403) );
  NAND2_X1 U15432 ( .A1(n13819), .A2(n6449), .ZN(n13402) );
  NAND2_X1 U15433 ( .A1(n13403), .A2(n13402), .ZN(n13405) );
  XNOR2_X1 U15434 ( .A(n13405), .B(n13404), .ZN(n13407) );
  AND2_X1 U15435 ( .A1(n13819), .A2(n10598), .ZN(n13406) );
  AOI21_X1 U15436 ( .B1(n13807), .B2(n13462), .A(n13406), .ZN(n13408) );
  NAND2_X1 U15437 ( .A1(n13407), .A2(n13408), .ZN(n13412) );
  INV_X1 U15438 ( .A(n13407), .ZN(n13410) );
  INV_X1 U15439 ( .A(n13408), .ZN(n13409) );
  NAND2_X1 U15440 ( .A1(n13410), .A2(n13409), .ZN(n13411) );
  NAND2_X1 U15441 ( .A1(n13494), .A2(n13412), .ZN(n13559) );
  NAND2_X1 U15442 ( .A1(n13988), .A2(n13465), .ZN(n13414) );
  NAND2_X1 U15443 ( .A1(n13583), .A2(n13462), .ZN(n13413) );
  NAND2_X1 U15444 ( .A1(n13414), .A2(n13413), .ZN(n13415) );
  XNOR2_X1 U15445 ( .A(n13415), .B(n13463), .ZN(n13419) );
  NAND2_X1 U15446 ( .A1(n13988), .A2(n6449), .ZN(n13417) );
  NAND2_X1 U15447 ( .A1(n13583), .A2(n10598), .ZN(n13416) );
  NAND2_X1 U15448 ( .A1(n13417), .A2(n13416), .ZN(n13418) );
  NOR2_X1 U15449 ( .A1(n13419), .A2(n13418), .ZN(n13420) );
  AOI21_X1 U15450 ( .B1(n13419), .B2(n13418), .A(n13420), .ZN(n13560) );
  NAND2_X1 U15451 ( .A1(n13559), .A2(n13560), .ZN(n13558) );
  INV_X1 U15452 ( .A(n13420), .ZN(n13421) );
  OAI21_X1 U15453 ( .B1(n13423), .B2(n13422), .A(n13461), .ZN(n13424) );
  NAND2_X1 U15454 ( .A1(n13424), .A2(n13570), .ZN(n13429) );
  AOI22_X1 U15455 ( .A1(n13425), .A2(n13562), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13426) );
  OAI21_X1 U15456 ( .B1(n13501), .B2(n14326), .A(n13426), .ZN(n13427) );
  AOI21_X1 U15457 ( .B1(n13567), .B2(n13759), .A(n13427), .ZN(n13428) );
  OAI211_X1 U15458 ( .C1(n14052), .C2(n13580), .A(n13429), .B(n13428), .ZN(
        P1_U3214) );
  INV_X1 U15459 ( .A(n13430), .ZN(n13435) );
  NOR3_X1 U15460 ( .A1(n13431), .A2(n13433), .A3(n13432), .ZN(n13434) );
  OAI21_X1 U15461 ( .B1(n13435), .B2(n13434), .A(n13570), .ZN(n13442) );
  NAND2_X1 U15462 ( .A1(n13584), .A2(n14507), .ZN(n13437) );
  NAND2_X1 U15463 ( .A1(n13487), .A2(n13929), .ZN(n13436) );
  NAND2_X1 U15464 ( .A1(n13437), .A2(n13436), .ZN(n13839) );
  INV_X1 U15465 ( .A(n13843), .ZN(n13439) );
  OAI22_X1 U15466 ( .A1(n13439), .A2(n14339), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13438), .ZN(n13440) );
  AOI21_X1 U15467 ( .B1(n13839), .B2(n13534), .A(n13440), .ZN(n13441) );
  OAI211_X1 U15468 ( .C1(n13845), .C2(n13580), .A(n13442), .B(n13441), .ZN(
        P1_U3216) );
  AOI21_X1 U15469 ( .B1(n13444), .B2(n13443), .A(n14330), .ZN(n13445) );
  NAND2_X1 U15470 ( .A1(n13445), .A2(n10617), .ZN(n13451) );
  AOI22_X1 U15471 ( .A1(n13577), .A2(n13599), .B1(n13446), .B2(n14335), .ZN(
        n13450) );
  AOI22_X1 U15472 ( .A1(n13567), .A2(n13597), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13449) );
  NAND2_X1 U15473 ( .A1(n13562), .A2(n13447), .ZN(n13448) );
  NAND4_X1 U15474 ( .A1(n13451), .A2(n13450), .A3(n13449), .A4(n13448), .ZN(
        P1_U3218) );
  INV_X1 U15475 ( .A(n13917), .ZN(n14073) );
  AND2_X1 U15476 ( .A1(n13549), .A2(n13452), .ZN(n13455) );
  OAI211_X1 U15477 ( .C1(n13455), .C2(n13454), .A(n13570), .B(n13453), .ZN(
        n13459) );
  NAND2_X1 U15478 ( .A1(n13577), .A2(n13912), .ZN(n13456) );
  NAND2_X1 U15479 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13728)
         );
  OAI211_X1 U15480 ( .C1(n13488), .C2(n14325), .A(n13456), .B(n13728), .ZN(
        n13457) );
  AOI21_X1 U15481 ( .B1(n13918), .B2(n13562), .A(n13457), .ZN(n13458) );
  OAI211_X1 U15482 ( .C1(n14073), .C2(n13580), .A(n13459), .B(n13458), .ZN(
        P1_U3219) );
  AOI22_X1 U15483 ( .A1(n13980), .A2(n6449), .B1(n10598), .B2(n13759), .ZN(
        n13464) );
  XNOR2_X1 U15484 ( .A(n13464), .B(n13463), .ZN(n13467) );
  AOI22_X1 U15485 ( .A1(n13980), .A2(n13465), .B1(n13462), .B2(n13759), .ZN(
        n13466) );
  XNOR2_X1 U15486 ( .A(n13467), .B(n13466), .ZN(n13468) );
  AOI22_X1 U15487 ( .A1(n13582), .A2(n14507), .B1(n13790), .B2(n13929), .ZN(
        n13771) );
  INV_X1 U15488 ( .A(n13469), .ZN(n13777) );
  AOI22_X1 U15489 ( .A1(n13777), .A2(n13562), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13470) );
  OAI21_X1 U15490 ( .B1(n13771), .B2(n13544), .A(n13470), .ZN(n13471) );
  AOI21_X1 U15491 ( .B1(n13980), .B2(n14335), .A(n13471), .ZN(n13472) );
  OAI21_X1 U15492 ( .B1(n13473), .B2(n14330), .A(n13472), .ZN(P1_U3220) );
  OAI21_X1 U15493 ( .B1(n13476), .B2(n13475), .A(n13474), .ZN(n13477) );
  NAND2_X1 U15494 ( .A1(n13477), .A2(n13570), .ZN(n13482) );
  AOI22_X1 U15495 ( .A1(n14335), .A2(n13479), .B1(n13478), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n13481) );
  AOI22_X1 U15496 ( .A1(n13577), .A2(n14518), .B1(n13567), .B2(n13599), .ZN(
        n13480) );
  NAND3_X1 U15497 ( .A1(n13482), .A2(n13481), .A3(n13480), .ZN(P1_U3222) );
  INV_X1 U15498 ( .A(n13879), .ZN(n14068) );
  OAI21_X1 U15499 ( .B1(n13484), .B2(n13483), .A(n13541), .ZN(n13485) );
  NAND2_X1 U15500 ( .A1(n13485), .A2(n13570), .ZN(n13493) );
  INV_X1 U15501 ( .A(n13486), .ZN(n13880) );
  NAND2_X1 U15502 ( .A1(n13487), .A2(n14507), .ZN(n13490) );
  OR2_X1 U15503 ( .A1(n13488), .A2(n14523), .ZN(n13489) );
  AND2_X1 U15504 ( .A1(n13490), .A2(n13489), .ZN(n13874) );
  OAI22_X1 U15505 ( .A1(n13874), .A2(n13544), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15112), .ZN(n13491) );
  AOI21_X1 U15506 ( .B1(n13880), .B2(n13562), .A(n13491), .ZN(n13492) );
  OAI211_X1 U15507 ( .C1(n14068), .C2(n13580), .A(n13493), .B(n13492), .ZN(
        P1_U3223) );
  INV_X1 U15508 ( .A(n13494), .ZN(n13499) );
  NOR3_X1 U15509 ( .A1(n13495), .A2(n13497), .A3(n13496), .ZN(n13498) );
  OAI21_X1 U15510 ( .B1(n13499), .B2(n13498), .A(n13570), .ZN(n13504) );
  OAI22_X1 U15511 ( .A1(n13501), .A2(n14533), .B1(n13500), .B2(n14523), .ZN(
        n13802) );
  OAI22_X1 U15512 ( .A1(n13810), .A2(n14339), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15171), .ZN(n13502) );
  AOI21_X1 U15513 ( .B1(n13802), .B2(n13534), .A(n13502), .ZN(n13503) );
  OAI211_X1 U15514 ( .C1(n6945), .C2(n13580), .A(n13504), .B(n13503), .ZN(
        P1_U3225) );
  AOI21_X1 U15515 ( .B1(n13506), .B2(n13505), .A(n6512), .ZN(n13513) );
  NAND2_X1 U15516 ( .A1(n13562), .A2(n13507), .ZN(n13508) );
  NAND2_X1 U15517 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14462)
         );
  OAI211_X1 U15518 ( .C1(n13509), .C2(n13544), .A(n13508), .B(n14462), .ZN(
        n13510) );
  AOI21_X1 U15519 ( .B1(n13511), .B2(n14335), .A(n13510), .ZN(n13512) );
  OAI21_X1 U15520 ( .B1(n13513), .B2(n14330), .A(n13512), .ZN(P1_U3226) );
  XNOR2_X1 U15521 ( .A(n13515), .B(n13514), .ZN(n13516) );
  XNOR2_X1 U15522 ( .A(n13517), .B(n13516), .ZN(n13522) );
  NAND2_X1 U15523 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14474)
         );
  OAI21_X1 U15524 ( .B1(n14326), .B2(n13947), .A(n14474), .ZN(n13518) );
  AOI21_X1 U15525 ( .B1(n13567), .B2(n13912), .A(n13518), .ZN(n13519) );
  OAI21_X1 U15526 ( .B1(n14339), .B2(n13953), .A(n13519), .ZN(n13520) );
  AOI21_X1 U15527 ( .B1(n14034), .B2(n14335), .A(n13520), .ZN(n13521) );
  OAI21_X1 U15528 ( .B1(n13522), .B2(n14330), .A(n13521), .ZN(P1_U3228) );
  INV_X1 U15529 ( .A(n13827), .ZN(n14059) );
  AND3_X1 U15530 ( .A1(n13430), .A2(n13524), .A3(n13523), .ZN(n13525) );
  OAI21_X1 U15531 ( .B1(n13495), .B2(n13525), .A(n13570), .ZN(n13529) );
  AOI22_X1 U15532 ( .A1(n13828), .A2(n13562), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13526) );
  OAI21_X1 U15533 ( .B1(n13565), .B2(n14325), .A(n13526), .ZN(n13527) );
  AOI21_X1 U15534 ( .B1(n13577), .B2(n13856), .A(n13527), .ZN(n13528) );
  OAI211_X1 U15535 ( .C1(n14059), .C2(n13580), .A(n13529), .B(n13528), .ZN(
        P1_U3229) );
  XNOR2_X1 U15536 ( .A(n13531), .B(n13530), .ZN(n13538) );
  NAND2_X1 U15537 ( .A1(n13585), .A2(n14507), .ZN(n13533) );
  OR2_X1 U15538 ( .A1(n13553), .A2(n14523), .ZN(n13532) );
  NAND2_X1 U15539 ( .A1(n13533), .A2(n13532), .ZN(n13893) );
  AOI22_X1 U15540 ( .A1(n13893), .A2(n13534), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13535) );
  OAI21_X1 U15541 ( .B1(n14339), .B2(n13896), .A(n13535), .ZN(n13536) );
  AOI21_X1 U15542 ( .B1(n13902), .B2(n14335), .A(n13536), .ZN(n13537) );
  OAI21_X1 U15543 ( .B1(n13538), .B2(n14330), .A(n13537), .ZN(P1_U3233) );
  AND3_X1 U15544 ( .A1(n13541), .A2(n13540), .A3(n13539), .ZN(n13542) );
  OAI21_X1 U15545 ( .B1(n13431), .B2(n13542), .A(n13570), .ZN(n13548) );
  NOR2_X1 U15546 ( .A1(n14339), .A2(n13857), .ZN(n13546) );
  NAND2_X1 U15547 ( .A1(n13585), .A2(n13929), .ZN(n13853) );
  OAI22_X1 U15548 ( .A1(n13853), .A2(n13544), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13543), .ZN(n13545) );
  AOI211_X1 U15549 ( .C1(n13567), .C2(n13856), .A(n13546), .B(n13545), .ZN(
        n13547) );
  OAI211_X1 U15550 ( .C1(n13580), .C2(n14064), .A(n13548), .B(n13547), .ZN(
        P1_U3235) );
  OAI21_X1 U15551 ( .B1(n13551), .B2(n13550), .A(n13549), .ZN(n13552) );
  NAND2_X1 U15552 ( .A1(n13552), .A2(n13570), .ZN(n13557) );
  NAND2_X1 U15553 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14490)
         );
  OAI21_X1 U15554 ( .B1(n14325), .B2(n13553), .A(n14490), .ZN(n13555) );
  NOR2_X1 U15555 ( .A1(n14339), .A2(n13937), .ZN(n13554) );
  AOI211_X1 U15556 ( .C1(n13577), .C2(n13928), .A(n13555), .B(n13554), .ZN(
        n13556) );
  OAI211_X1 U15557 ( .C1(n6943), .C2(n13580), .A(n13557), .B(n13556), .ZN(
        P1_U3238) );
  INV_X1 U15558 ( .A(n13988), .ZN(n13796) );
  OAI21_X1 U15559 ( .B1(n13560), .B2(n13559), .A(n13558), .ZN(n13561) );
  NAND2_X1 U15560 ( .A1(n13561), .A2(n13570), .ZN(n13569) );
  INV_X1 U15561 ( .A(n13792), .ZN(n13563) );
  AOI22_X1 U15562 ( .A1(n13563), .A2(n13562), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13564) );
  OAI21_X1 U15563 ( .B1(n13565), .B2(n14326), .A(n13564), .ZN(n13566) );
  AOI21_X1 U15564 ( .B1(n13790), .B2(n13567), .A(n13566), .ZN(n13568) );
  OAI211_X1 U15565 ( .C1(n13796), .C2(n13580), .A(n13569), .B(n13568), .ZN(
        P1_U3240) );
  OAI211_X1 U15566 ( .C1(n13573), .C2(n13572), .A(n13571), .B(n13570), .ZN(
        n13579) );
  NAND2_X1 U15567 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14444)
         );
  OAI21_X1 U15568 ( .B1(n14325), .B2(n13947), .A(n14444), .ZN(n13576) );
  NOR2_X1 U15569 ( .A1(n14339), .A2(n13574), .ZN(n13575) );
  AOI211_X1 U15570 ( .C1(n13577), .C2(n13588), .A(n13576), .B(n13575), .ZN(
        n13578) );
  OAI211_X1 U15571 ( .C1(n13581), .C2(n13580), .A(n13579), .B(n13578), .ZN(
        P1_U3241) );
  MUX2_X1 U15572 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13734), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15573 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13745), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15574 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13582), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15575 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13759), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15576 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13790), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15577 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13583), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15578 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13819), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15579 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13584), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15580 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13856), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15581 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13585), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15582 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13913), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15583 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13930), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15584 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13912), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15585 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13928), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15586 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13586), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15587 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13587), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15588 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13588), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15589 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13589), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15590 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13590), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15591 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14506), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15592 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13591), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15593 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13592), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15594 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13593), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U15595 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13594), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15596 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13595), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15597 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13596), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15598 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13597), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15599 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13598), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15600 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13599), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15601 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n8100), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15602 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14518), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI22_X1 U15603 ( .A1(n14492), .A2(n6876), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13600), .ZN(n13601) );
  AOI21_X1 U15604 ( .B1(n13602), .B2(n14489), .A(n13601), .ZN(n13610) );
  OAI211_X1 U15605 ( .C1(n13605), .C2(n13604), .A(n14442), .B(n13603), .ZN(
        n13609) );
  OAI211_X1 U15606 ( .C1(n13607), .C2(n13612), .A(n14440), .B(n13606), .ZN(
        n13608) );
  NAND3_X1 U15607 ( .A1(n13610), .A2(n13609), .A3(n13608), .ZN(P1_U3244) );
  MUX2_X1 U15608 ( .A(n13612), .B(n13611), .S(n8684), .Z(n13614) );
  NAND2_X1 U15609 ( .A1(n13614), .A2(n13613), .ZN(n13615) );
  OAI211_X1 U15610 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n13616), .A(n13615), .B(
        P1_U4016), .ZN(n13657) );
  OAI22_X1 U15611 ( .A1(n14492), .A2(n6879), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13617), .ZN(n13618) );
  AOI21_X1 U15612 ( .B1(n13619), .B2(n14489), .A(n13618), .ZN(n13628) );
  OAI211_X1 U15613 ( .C1(n13622), .C2(n13621), .A(n14440), .B(n13620), .ZN(
        n13627) );
  OAI211_X1 U15614 ( .C1(n13625), .C2(n13624), .A(n14442), .B(n13623), .ZN(
        n13626) );
  NAND4_X1 U15615 ( .A1(n13657), .A2(n13628), .A3(n13627), .A4(n13626), .ZN(
        P1_U3245) );
  INV_X1 U15616 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14140) );
  NAND2_X1 U15617 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n13629) );
  OAI21_X1 U15618 ( .B1(n14492), .B2(n14140), .A(n13629), .ZN(n13630) );
  AOI21_X1 U15619 ( .B1(n13631), .B2(n14489), .A(n13630), .ZN(n13640) );
  OAI211_X1 U15620 ( .C1(n13634), .C2(n13633), .A(n14440), .B(n13632), .ZN(
        n13639) );
  OAI211_X1 U15621 ( .C1(n13637), .C2(n13636), .A(n14442), .B(n13635), .ZN(
        n13638) );
  NAND3_X1 U15622 ( .A1(n13640), .A2(n13639), .A3(n13638), .ZN(P1_U3246) );
  AOI21_X1 U15623 ( .B1(n13642), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n13641), .ZN(
        n13656) );
  INV_X1 U15624 ( .A(n13643), .ZN(n13644) );
  NAND2_X1 U15625 ( .A1(n14489), .A2(n13644), .ZN(n13650) );
  OAI21_X1 U15626 ( .B1(n13647), .B2(n13646), .A(n13645), .ZN(n13648) );
  OR2_X1 U15627 ( .A1(n14482), .A2(n13648), .ZN(n13649) );
  AND2_X1 U15628 ( .A1(n13650), .A2(n13649), .ZN(n13655) );
  OAI211_X1 U15629 ( .C1(n13653), .C2(n13652), .A(n14440), .B(n13651), .ZN(
        n13654) );
  NAND4_X1 U15630 ( .A1(n13657), .A2(n13656), .A3(n13655), .A4(n13654), .ZN(
        P1_U3247) );
  INV_X1 U15631 ( .A(n13658), .ZN(n13661) );
  INV_X1 U15632 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14150) );
  NAND2_X1 U15633 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n13659) );
  OAI21_X1 U15634 ( .B1(n14492), .B2(n14150), .A(n13659), .ZN(n13660) );
  AOI21_X1 U15635 ( .B1(n13661), .B2(n14489), .A(n13660), .ZN(n13670) );
  OAI211_X1 U15636 ( .C1(n13664), .C2(n13663), .A(n14442), .B(n13662), .ZN(
        n13669) );
  OAI211_X1 U15637 ( .C1(n13667), .C2(n13666), .A(n14440), .B(n13665), .ZN(
        n13668) );
  NAND3_X1 U15638 ( .A1(n13670), .A2(n13669), .A3(n13668), .ZN(P1_U3249) );
  INV_X1 U15639 ( .A(n13671), .ZN(n13675) );
  INV_X1 U15640 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n13673) );
  NAND2_X1 U15641 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n13672) );
  OAI21_X1 U15642 ( .B1(n14492), .B2(n13673), .A(n13672), .ZN(n13674) );
  AOI21_X1 U15643 ( .B1(n13675), .B2(n14489), .A(n13674), .ZN(n13684) );
  OAI211_X1 U15644 ( .C1(n13678), .C2(n13677), .A(n14440), .B(n13676), .ZN(
        n13683) );
  OAI211_X1 U15645 ( .C1(n13681), .C2(n13680), .A(n14442), .B(n13679), .ZN(
        n13682) );
  NAND3_X1 U15646 ( .A1(n13684), .A2(n13683), .A3(n13682), .ZN(P1_U3250) );
  OAI211_X1 U15647 ( .C1(n13687), .C2(n13686), .A(n13685), .B(n14442), .ZN(
        n13697) );
  INV_X1 U15648 ( .A(n13688), .ZN(n13691) );
  INV_X1 U15649 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14110) );
  OAI21_X1 U15650 ( .B1(n14492), .B2(n14110), .A(n13689), .ZN(n13690) );
  AOI21_X1 U15651 ( .B1(n13691), .B2(n14489), .A(n13690), .ZN(n13696) );
  OAI211_X1 U15652 ( .C1(n13694), .C2(n13693), .A(n13692), .B(n14440), .ZN(
        n13695) );
  NAND3_X1 U15653 ( .A1(n13697), .A2(n13696), .A3(n13695), .ZN(P1_U3253) );
  INV_X1 U15654 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14484) );
  NAND2_X1 U15655 ( .A1(n14459), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n13699) );
  NAND2_X1 U15656 ( .A1(n13717), .A2(n8350), .ZN(n13698) );
  AND2_X1 U15657 ( .A1(n13699), .A2(n13698), .ZN(n14452) );
  MUX2_X1 U15658 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n13700), .S(n13714), .Z(
        n14423) );
  INV_X1 U15659 ( .A(n14417), .ZN(n13712) );
  AOI21_X1 U15660 ( .B1(n13702), .B2(n13710), .A(n13701), .ZN(n14409) );
  INV_X1 U15661 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n14372) );
  MUX2_X1 U15662 ( .A(n14372), .B(P1_REG1_REG_13__SCAN_IN), .S(n14417), .Z(
        n14410) );
  NAND2_X1 U15663 ( .A1(n14423), .A2(n14424), .ZN(n14422) );
  NAND2_X1 U15664 ( .A1(n14437), .A2(n13703), .ZN(n13704) );
  INV_X1 U15665 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14435) );
  NAND2_X1 U15666 ( .A1(n13704), .A2(n14434), .ZN(n14453) );
  NOR2_X1 U15667 ( .A1(n14452), .A2(n14453), .ZN(n14454) );
  XNOR2_X1 U15668 ( .A(n14473), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n14469) );
  NOR2_X1 U15669 ( .A1(n14470), .A2(n14469), .ZN(n14468) );
  XNOR2_X1 U15670 ( .A(n14477), .B(n13705), .ZN(n14485) );
  NOR2_X1 U15671 ( .A1(n14484), .A2(n14485), .ZN(n14483) );
  NOR2_X1 U15672 ( .A1(n13705), .A2(n14477), .ZN(n13706) );
  NOR2_X1 U15673 ( .A1(n14483), .A2(n13706), .ZN(n13707) );
  XOR2_X1 U15674 ( .A(n13707), .B(P1_REG1_REG_19__SCAN_IN), .Z(n13724) );
  AOI21_X1 U15675 ( .B1(n13724), .B2(n14442), .A(n14489), .ZN(n13723) );
  NAND2_X1 U15676 ( .A1(n13717), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n13708) );
  OAI21_X1 U15677 ( .B1(n13717), .B2(P1_REG2_REG_16__SCAN_IN), .A(n13708), 
        .ZN(n14447) );
  AOI21_X1 U15678 ( .B1(n13711), .B2(n13710), .A(n13709), .ZN(n14413) );
  MUX2_X1 U15679 ( .A(n8298), .B(P1_REG2_REG_13__SCAN_IN), .S(n14417), .Z(
        n14414) );
  AOI21_X1 U15680 ( .B1(n13712), .B2(P1_REG2_REG_13__SCAN_IN), .A(n14411), 
        .ZN(n14428) );
  MUX2_X1 U15681 ( .A(n13713), .B(P1_REG2_REG_14__SCAN_IN), .S(n13714), .Z(
        n14427) );
  NOR2_X1 U15682 ( .A1(n14428), .A2(n14427), .ZN(n14426) );
  AOI21_X1 U15683 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n13714), .A(n14426), 
        .ZN(n13715) );
  NAND2_X1 U15684 ( .A1(n13715), .A2(n14437), .ZN(n13716) );
  XOR2_X1 U15685 ( .A(n13715), .B(n14437), .Z(n14439) );
  NAND2_X1 U15686 ( .A1(n14439), .A2(n11770), .ZN(n14438) );
  NAND2_X1 U15687 ( .A1(n13716), .A2(n14438), .ZN(n14448) );
  NOR2_X1 U15688 ( .A1(n14447), .A2(n14448), .ZN(n14449) );
  AOI21_X1 U15689 ( .B1(n13717), .B2(P1_REG2_REG_16__SCAN_IN), .A(n14449), 
        .ZN(n14467) );
  NAND2_X1 U15690 ( .A1(n14473), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n13718) );
  OAI21_X1 U15691 ( .B1(n14473), .B2(P1_REG2_REG_17__SCAN_IN), .A(n13718), 
        .ZN(n14466) );
  NOR2_X1 U15692 ( .A1(n14467), .A2(n14466), .ZN(n14465) );
  AOI21_X1 U15693 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n14473), .A(n14465), 
        .ZN(n13719) );
  NOR2_X1 U15694 ( .A1(n13719), .A2(n14477), .ZN(n13720) );
  XNOR2_X1 U15695 ( .A(n14477), .B(n13719), .ZN(n14481) );
  NOR2_X1 U15696 ( .A1(n14480), .A2(n14481), .ZN(n14479) );
  NOR2_X1 U15697 ( .A1(n13720), .A2(n14479), .ZN(n13721) );
  XOR2_X1 U15698 ( .A(n13721), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13725) );
  NAND2_X1 U15699 ( .A1(n13725), .A2(n14440), .ZN(n13722) );
  NAND2_X1 U15700 ( .A1(n13723), .A2(n13722), .ZN(n13727) );
  OAI22_X1 U15701 ( .A1(n13725), .A2(n14478), .B1(n13724), .B2(n14482), .ZN(
        n13726) );
  OAI21_X1 U15702 ( .B1(n14492), .B2(n7410), .A(n13728), .ZN(n13729) );
  NOR2_X1 U15703 ( .A1(n14543), .A2(n13731), .ZN(n13735) );
  INV_X1 U15704 ( .A(P1_B_REG_SCAN_IN), .ZN(n13732) );
  NOR2_X1 U15705 ( .A1(n8684), .A2(n13732), .ZN(n13733) );
  NOR2_X1 U15706 ( .A1(n14533), .A2(n13733), .ZN(n13746) );
  NAND2_X1 U15707 ( .A1(n13746), .A2(n13734), .ZN(n13965) );
  NOR2_X1 U15708 ( .A1(n14545), .A2(n13965), .ZN(n13741) );
  AOI211_X1 U15709 ( .C1(n13736), .C2(n14501), .A(n13735), .B(n13741), .ZN(
        n13737) );
  OAI21_X1 U15710 ( .B1(n13964), .B2(n13899), .A(n13737), .ZN(P1_U3263) );
  INV_X1 U15711 ( .A(n13740), .ZN(n14045) );
  INV_X1 U15712 ( .A(n13738), .ZN(n13739) );
  AOI211_X1 U15713 ( .C1(n13740), .C2(n13744), .A(n14526), .B(n13739), .ZN(
        n13967) );
  NAND2_X1 U15714 ( .A1(n13967), .A2(n14511), .ZN(n13743) );
  AOI21_X1 U15715 ( .B1(n14545), .B2(P1_REG2_REG_30__SCAN_IN), .A(n13741), 
        .ZN(n13742) );
  OAI211_X1 U15716 ( .C1(n14045), .C2(n13958), .A(n13743), .B(n13742), .ZN(
        P1_U3264) );
  OAI211_X1 U15717 ( .C1(n13970), .C2(n13776), .A(n14508), .B(n13744), .ZN(
        n13974) );
  NAND2_X1 U15718 ( .A1(n13746), .A2(n13745), .ZN(n13971) );
  OAI21_X1 U15719 ( .B1(n13974), .B2(n13747), .A(n13971), .ZN(n13748) );
  INV_X1 U15720 ( .A(n13748), .ZN(n13768) );
  INV_X1 U15721 ( .A(n13759), .ZN(n13751) );
  AND2_X1 U15722 ( .A1(n13980), .A2(n13751), .ZN(n13752) );
  XNOR2_X1 U15723 ( .A(n13753), .B(n13757), .ZN(n13754) );
  NAND2_X1 U15724 ( .A1(n13754), .A2(n14519), .ZN(n13758) );
  NAND2_X1 U15725 ( .A1(n13759), .A2(n13929), .ZN(n13972) );
  INV_X1 U15726 ( .A(n13972), .ZN(n13760) );
  INV_X1 U15727 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n13761) );
  OAI22_X1 U15728 ( .A1(n13762), .A2(n13952), .B1(n13761), .B2(n14543), .ZN(
        n13763) );
  AOI21_X1 U15729 ( .B1(n13764), .B2(n14501), .A(n13763), .ZN(n13765) );
  OAI211_X1 U15730 ( .C1(n13768), .C2(n13767), .A(n13766), .B(n13765), .ZN(
        P1_U3356) );
  XNOR2_X1 U15731 ( .A(n13769), .B(n13770), .ZN(n13773) );
  INV_X1 U15732 ( .A(n13771), .ZN(n13772) );
  AND2_X1 U15733 ( .A1(n13980), .A2(n13774), .ZN(n13775) );
  NOR3_X1 U15734 ( .A1(n13776), .A2(n13775), .A3(n14526), .ZN(n13979) );
  NAND2_X1 U15735 ( .A1(n13980), .A2(n14501), .ZN(n13779) );
  AOI22_X1 U15736 ( .A1(n13777), .A2(n14542), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n14545), .ZN(n13778) );
  NAND2_X1 U15737 ( .A1(n13779), .A2(n13778), .ZN(n13784) );
  NOR2_X1 U15738 ( .A1(n13983), .A2(n13963), .ZN(n13783) );
  AOI211_X1 U15739 ( .C1(n13979), .C2(n14511), .A(n13784), .B(n13783), .ZN(
        n13785) );
  OAI21_X1 U15740 ( .B1(n14545), .B2(n13982), .A(n13785), .ZN(P1_U3265) );
  OAI21_X1 U15741 ( .B1(n13787), .B2(n6706), .A(n13786), .ZN(n13991) );
  XNOR2_X1 U15742 ( .A(n13788), .B(n13789), .ZN(n13791) );
  AOI222_X1 U15743 ( .A1(n14519), .A2(n13791), .B1(n13790), .B2(n14507), .C1(
        n13819), .C2(n13929), .ZN(n13990) );
  OAI21_X1 U15744 ( .B1(n13792), .B2(n13952), .A(n13990), .ZN(n13793) );
  NAND2_X1 U15745 ( .A1(n13793), .A2(n14543), .ZN(n13799) );
  AOI211_X1 U15746 ( .C1(n13988), .C2(n13808), .A(n14526), .B(n13794), .ZN(
        n13987) );
  INV_X1 U15747 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n13795) );
  OAI22_X1 U15748 ( .A1(n13796), .A2(n13958), .B1(n14543), .B2(n13795), .ZN(
        n13797) );
  AOI21_X1 U15749 ( .B1(n13987), .B2(n14511), .A(n13797), .ZN(n13798) );
  OAI211_X1 U15750 ( .C1(n13991), .C2(n13963), .A(n13799), .B(n13798), .ZN(
        P1_U3267) );
  OAI21_X1 U15751 ( .B1(n13800), .B2(n7223), .A(n13801), .ZN(n13803) );
  NAND2_X1 U15752 ( .A1(n13804), .A2(n7223), .ZN(n13805) );
  AOI21_X1 U15753 ( .B1(n13826), .B2(n13807), .A(n14526), .ZN(n13809) );
  NAND2_X1 U15754 ( .A1(n13994), .A2(n14511), .ZN(n13813) );
  INV_X1 U15755 ( .A(n13810), .ZN(n13811) );
  AOI22_X1 U15756 ( .A1(n13811), .A2(n14542), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n14545), .ZN(n13812) );
  OAI211_X1 U15757 ( .C1(n6945), .C2(n13958), .A(n13813), .B(n13812), .ZN(
        n13814) );
  AOI21_X1 U15758 ( .B1(n13995), .B2(n14512), .A(n13814), .ZN(n13815) );
  OAI21_X1 U15759 ( .B1(n13992), .B2(n14545), .A(n13815), .ZN(P1_U3268) );
  INV_X1 U15760 ( .A(n13816), .ZN(n13817) );
  AOI21_X1 U15761 ( .B1(n13821), .B2(n13818), .A(n13817), .ZN(n13825) );
  AOI22_X1 U15762 ( .A1(n13819), .A2(n14507), .B1(n13929), .B2(n13856), .ZN(
        n13824) );
  OAI211_X1 U15763 ( .C1(n13822), .C2(n13821), .A(n14519), .B(n13820), .ZN(
        n13823) );
  OAI211_X1 U15764 ( .C1(n13825), .C2(n14549), .A(n13824), .B(n13823), .ZN(
        n13999) );
  INV_X1 U15765 ( .A(n13999), .ZN(n13832) );
  AOI211_X1 U15766 ( .C1(n13827), .C2(n13842), .A(n14526), .B(n6946), .ZN(
        n13998) );
  AOI22_X1 U15767 ( .A1(n13828), .A2(n14542), .B1(n14545), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n13829) );
  OAI21_X1 U15768 ( .B1(n14059), .B2(n13958), .A(n13829), .ZN(n13830) );
  AOI21_X1 U15769 ( .B1(n13998), .B2(n14511), .A(n13830), .ZN(n13831) );
  OAI21_X1 U15770 ( .B1(n13832), .B2(n14545), .A(n13831), .ZN(P1_U3269) );
  NAND2_X1 U15771 ( .A1(n13833), .A2(n13837), .ZN(n13834) );
  NAND2_X1 U15772 ( .A1(n13835), .A2(n13834), .ZN(n14004) );
  XNOR2_X1 U15773 ( .A(n13836), .B(n13837), .ZN(n13838) );
  NAND2_X1 U15774 ( .A1(n13838), .A2(n14519), .ZN(n13841) );
  INV_X1 U15775 ( .A(n13839), .ZN(n13840) );
  NAND2_X1 U15776 ( .A1(n13841), .A2(n13840), .ZN(n14006) );
  NAND2_X1 U15777 ( .A1(n14006), .A2(n14543), .ZN(n13849) );
  OAI211_X1 U15778 ( .C1(n13845), .C2(n13860), .A(n14508), .B(n13842), .ZN(
        n14002) );
  INV_X1 U15779 ( .A(n14002), .ZN(n13847) );
  AOI22_X1 U15780 ( .A1(n14545), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n13843), 
        .B2(n14542), .ZN(n13844) );
  OAI21_X1 U15781 ( .B1(n13845), .B2(n13958), .A(n13844), .ZN(n13846) );
  AOI21_X1 U15782 ( .B1(n13847), .B2(n14511), .A(n13846), .ZN(n13848) );
  OAI211_X1 U15783 ( .C1(n14004), .C2(n13963), .A(n13849), .B(n13848), .ZN(
        P1_U3270) );
  NAND2_X1 U15784 ( .A1(n13850), .A2(n13861), .ZN(n13851) );
  NAND2_X1 U15785 ( .A1(n13852), .A2(n13851), .ZN(n13855) );
  INV_X1 U15786 ( .A(n13853), .ZN(n13854) );
  AOI21_X1 U15787 ( .B1(n13855), .B2(n14519), .A(n13854), .ZN(n14011) );
  NAND2_X1 U15788 ( .A1(n13856), .A2(n14507), .ZN(n14009) );
  OAI211_X1 U15789 ( .C1(n13952), .C2(n13857), .A(n14011), .B(n14009), .ZN(
        n13867) );
  NAND2_X1 U15790 ( .A1(n13863), .A2(n13878), .ZN(n13858) );
  NAND2_X1 U15791 ( .A1(n13858), .A2(n14508), .ZN(n13859) );
  OR2_X1 U15792 ( .A1(n13860), .A2(n13859), .ZN(n14008) );
  XNOR2_X1 U15793 ( .A(n13862), .B(n13861), .ZN(n14007) );
  NAND2_X1 U15794 ( .A1(n14007), .A2(n14512), .ZN(n13865) );
  AOI22_X1 U15795 ( .A1(n13863), .A2(n14501), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n14545), .ZN(n13864) );
  OAI211_X1 U15796 ( .C1(n14008), .C2(n13899), .A(n13865), .B(n13864), .ZN(
        n13866) );
  AOI21_X1 U15797 ( .B1(n13867), .B2(n14543), .A(n13866), .ZN(n13868) );
  INV_X1 U15798 ( .A(n13868), .ZN(P1_U3271) );
  NAND3_X1 U15799 ( .A1(n13869), .A2(n6450), .A3(n13871), .ZN(n13872) );
  NAND3_X1 U15800 ( .A1(n13873), .A2(n14519), .A3(n13872), .ZN(n13875) );
  NAND2_X1 U15801 ( .A1(n13875), .A2(n13874), .ZN(n14014) );
  INV_X1 U15802 ( .A(n14014), .ZN(n13885) );
  OAI21_X1 U15803 ( .B1(n13877), .B2(n6450), .A(n13876), .ZN(n14016) );
  AOI211_X1 U15804 ( .C1(n13879), .C2(n13898), .A(n14526), .B(n6617), .ZN(
        n14015) );
  NAND2_X1 U15805 ( .A1(n14015), .A2(n14511), .ZN(n13882) );
  AOI22_X1 U15806 ( .A1(n14545), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n13880), 
        .B2(n14542), .ZN(n13881) );
  OAI211_X1 U15807 ( .C1(n14068), .C2(n13958), .A(n13882), .B(n13881), .ZN(
        n13883) );
  AOI21_X1 U15808 ( .B1(n14016), .B2(n14512), .A(n13883), .ZN(n13884) );
  OAI21_X1 U15809 ( .B1(n13885), .B2(n14545), .A(n13884), .ZN(P1_U3272) );
  NAND2_X1 U15810 ( .A1(n13887), .A2(n13888), .ZN(n13889) );
  NAND2_X1 U15811 ( .A1(n13886), .A2(n13889), .ZN(n14022) );
  NAND2_X1 U15812 ( .A1(n13891), .A2(n13890), .ZN(n13892) );
  NAND3_X1 U15813 ( .A1(n13869), .A2(n14519), .A3(n13892), .ZN(n13895) );
  INV_X1 U15814 ( .A(n13893), .ZN(n13894) );
  NAND2_X1 U15815 ( .A1(n13895), .A2(n13894), .ZN(n14024) );
  NAND2_X1 U15816 ( .A1(n14024), .A2(n14543), .ZN(n13904) );
  INV_X1 U15817 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n13897) );
  OAI22_X1 U15818 ( .A1(n14543), .A2(n13897), .B1(n13896), .B2(n13952), .ZN(
        n13901) );
  OAI211_X1 U15819 ( .C1(n13916), .C2(n14019), .A(n14508), .B(n13898), .ZN(
        n14020) );
  NOR2_X1 U15820 ( .A1(n14020), .A2(n13899), .ZN(n13900) );
  AOI211_X1 U15821 ( .C1(n14501), .C2(n13902), .A(n13901), .B(n13900), .ZN(
        n13903) );
  OAI211_X1 U15822 ( .C1(n14022), .C2(n13963), .A(n13904), .B(n13903), .ZN(
        P1_U3273) );
  INV_X1 U15823 ( .A(n13907), .ZN(n13906) );
  NAND2_X1 U15824 ( .A1(n13906), .A2(n14588), .ZN(n13911) );
  AOI22_X1 U15825 ( .A1(n13908), .A2(n14519), .B1(n14588), .B2(n13907), .ZN(
        n13910) );
  MUX2_X1 U15826 ( .A(n13911), .B(n13910), .S(n13909), .Z(n13915) );
  AOI22_X1 U15827 ( .A1(n13913), .A2(n14507), .B1(n13929), .B2(n13912), .ZN(
        n13914) );
  OAI211_X1 U15828 ( .C1(n14548), .C2(n13905), .A(n13915), .B(n13914), .ZN(
        n14026) );
  INV_X1 U15829 ( .A(n14026), .ZN(n13922) );
  AOI211_X1 U15830 ( .C1(n13917), .C2(n13934), .A(n14526), .B(n13916), .ZN(
        n14025) );
  AOI22_X1 U15831 ( .A1(n14545), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n13918), 
        .B2(n14542), .ZN(n13919) );
  OAI21_X1 U15832 ( .B1(n14073), .B2(n13958), .A(n13919), .ZN(n13920) );
  AOI21_X1 U15833 ( .B1(n14025), .B2(n14511), .A(n13920), .ZN(n13921) );
  OAI21_X1 U15834 ( .B1(n13922), .B2(n14545), .A(n13921), .ZN(P1_U3274) );
  XNOR2_X1 U15835 ( .A(n13923), .B(n13924), .ZN(n13933) );
  OAI211_X1 U15836 ( .C1(n13927), .C2(n13926), .A(n13925), .B(n14519), .ZN(
        n13932) );
  AOI22_X1 U15837 ( .A1(n13930), .A2(n14507), .B1(n13929), .B2(n13928), .ZN(
        n13931) );
  OAI211_X1 U15838 ( .C1(n13933), .C2(n14549), .A(n13932), .B(n13931), .ZN(
        n14030) );
  INV_X1 U15839 ( .A(n14030), .ZN(n13942) );
  INV_X1 U15840 ( .A(n13934), .ZN(n13935) );
  AOI211_X1 U15841 ( .C1(n13936), .C2(n13955), .A(n14526), .B(n13935), .ZN(
        n14029) );
  INV_X1 U15842 ( .A(n13937), .ZN(n13938) );
  AOI22_X1 U15843 ( .A1(n14545), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n13938), 
        .B2(n14542), .ZN(n13939) );
  OAI21_X1 U15844 ( .B1(n6943), .B2(n13958), .A(n13939), .ZN(n13940) );
  AOI21_X1 U15845 ( .B1(n14029), .B2(n14511), .A(n13940), .ZN(n13941) );
  OAI21_X1 U15846 ( .B1(n13942), .B2(n14545), .A(n13941), .ZN(P1_U3275) );
  XNOR2_X1 U15847 ( .A(n13944), .B(n13943), .ZN(n14037) );
  AOI21_X1 U15848 ( .B1(n13946), .B2(n13945), .A(n14548), .ZN(n13951) );
  OAI22_X1 U15849 ( .A1(n13948), .A2(n14533), .B1(n13947), .B2(n14523), .ZN(
        n13949) );
  AOI21_X1 U15850 ( .B1(n13951), .B2(n13950), .A(n13949), .ZN(n14036) );
  OAI21_X1 U15851 ( .B1(n13953), .B2(n13952), .A(n14036), .ZN(n13954) );
  NAND2_X1 U15852 ( .A1(n13954), .A2(n14543), .ZN(n13962) );
  AOI211_X1 U15853 ( .C1(n14034), .C2(n13956), .A(n14526), .B(n6944), .ZN(
        n14033) );
  INV_X1 U15854 ( .A(n14034), .ZN(n13959) );
  OAI22_X1 U15855 ( .A1(n13959), .A2(n13958), .B1(n14543), .B2(n13957), .ZN(
        n13960) );
  AOI21_X1 U15856 ( .B1(n14033), .B2(n14511), .A(n13960), .ZN(n13961) );
  OAI211_X1 U15857 ( .C1(n14037), .C2(n13963), .A(n13962), .B(n13961), .ZN(
        P1_U3276) );
  INV_X1 U15858 ( .A(n13965), .ZN(n13966) );
  NOR2_X1 U15859 ( .A1(n13967), .A2(n13966), .ZN(n14042) );
  MUX2_X1 U15860 ( .A(n13968), .B(n14042), .S(n14597), .Z(n13969) );
  OAI21_X1 U15861 ( .B1(n14045), .B2(n14032), .A(n13969), .ZN(P1_U3558) );
  OR2_X1 U15862 ( .A1(n13970), .A2(n14584), .ZN(n13973) );
  NAND4_X1 U15863 ( .A1(n13974), .A2(n13973), .A3(n13972), .A4(n13971), .ZN(
        n13975) );
  NOR2_X1 U15864 ( .A1(n13976), .A2(n13975), .ZN(n14046) );
  INV_X1 U15865 ( .A(n13978), .ZN(P1_U3557) );
  AOI21_X1 U15866 ( .B1(n13980), .B2(n14574), .A(n13979), .ZN(n13981) );
  OAI211_X1 U15867 ( .C1(n14549), .C2(n13983), .A(n13982), .B(n13981), .ZN(
        n14049) );
  MUX2_X1 U15868 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14049), .S(n14597), .Z(
        P1_U3556) );
  OAI21_X1 U15869 ( .B1(n14052), .B2(n14032), .A(n13986), .ZN(P1_U3555) );
  AOI21_X1 U15870 ( .B1(n13988), .B2(n14574), .A(n13987), .ZN(n13989) );
  OAI211_X1 U15871 ( .C1(n14549), .C2(n13991), .A(n13990), .B(n13989), .ZN(
        n14053) );
  MUX2_X1 U15872 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14053), .S(n14597), .Z(
        P1_U3554) );
  INV_X1 U15873 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n13996) );
  INV_X1 U15874 ( .A(n13992), .ZN(n13993) );
  AOI211_X2 U15875 ( .C1(n14588), .C2(n13995), .A(n13994), .B(n13993), .ZN(
        n14054) );
  MUX2_X1 U15876 ( .A(n13996), .B(n14054), .S(n14597), .Z(n13997) );
  NOR2_X1 U15877 ( .A1(n13999), .A2(n13998), .ZN(n14056) );
  MUX2_X1 U15878 ( .A(n15108), .B(n14056), .S(n14597), .Z(n14000) );
  OAI21_X1 U15879 ( .B1(n14059), .B2(n14032), .A(n14000), .ZN(P1_U3552) );
  NAND2_X1 U15880 ( .A1(n14001), .A2(n14574), .ZN(n14003) );
  OAI211_X1 U15881 ( .C1(n14004), .C2(n14549), .A(n14003), .B(n14002), .ZN(
        n14005) );
  MUX2_X1 U15882 ( .A(n14060), .B(P1_REG1_REG_23__SCAN_IN), .S(n14595), .Z(
        P1_U3551) );
  NAND2_X1 U15883 ( .A1(n14007), .A2(n14588), .ZN(n14010) );
  NAND4_X1 U15884 ( .A1(n14011), .A2(n14010), .A3(n14009), .A4(n14008), .ZN(
        n14061) );
  MUX2_X1 U15885 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14061), .S(n14597), .Z(
        n14012) );
  INV_X1 U15886 ( .A(n14012), .ZN(n14013) );
  OAI21_X1 U15887 ( .B1(n14032), .B2(n14064), .A(n14013), .ZN(P1_U3550) );
  AOI211_X1 U15888 ( .C1(n14588), .C2(n14016), .A(n14015), .B(n14014), .ZN(
        n14065) );
  MUX2_X1 U15889 ( .A(n14017), .B(n14065), .S(n14597), .Z(n14018) );
  OAI21_X1 U15890 ( .B1(n14068), .B2(n14032), .A(n14018), .ZN(P1_U3549) );
  OR2_X1 U15891 ( .A1(n14019), .A2(n14584), .ZN(n14021) );
  OAI211_X1 U15892 ( .C1(n14022), .C2(n14549), .A(n14021), .B(n14020), .ZN(
        n14023) );
  MUX2_X1 U15893 ( .A(n14069), .B(P1_REG1_REG_20__SCAN_IN), .S(n14595), .Z(
        P1_U3548) );
  NOR2_X1 U15894 ( .A1(n14026), .A2(n14025), .ZN(n14070) );
  MUX2_X1 U15895 ( .A(n14027), .B(n14070), .S(n14597), .Z(n14028) );
  OAI21_X1 U15896 ( .B1(n14073), .B2(n14032), .A(n14028), .ZN(P1_U3547) );
  NOR2_X1 U15897 ( .A1(n14030), .A2(n14029), .ZN(n14074) );
  MUX2_X1 U15898 ( .A(n14484), .B(n14074), .S(n14597), .Z(n14031) );
  OAI21_X1 U15899 ( .B1(n6943), .B2(n14032), .A(n14031), .ZN(P1_U3546) );
  AOI21_X1 U15900 ( .B1(n14034), .B2(n14574), .A(n14033), .ZN(n14035) );
  OAI211_X1 U15901 ( .C1(n14549), .C2(n14037), .A(n14036), .B(n14035), .ZN(
        n14078) );
  MUX2_X1 U15902 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14078), .S(n14597), .Z(
        P1_U3545) );
  MUX2_X1 U15903 ( .A(n14039), .B(n14038), .S(n14589), .Z(n14040) );
  OAI21_X1 U15904 ( .B1(n14041), .B2(n14077), .A(n14040), .ZN(P1_U3527) );
  INV_X1 U15905 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14043) );
  MUX2_X1 U15906 ( .A(n14043), .B(n14042), .S(n14589), .Z(n14044) );
  OAI21_X1 U15907 ( .B1(n14045), .B2(n14077), .A(n14044), .ZN(P1_U3526) );
  INV_X1 U15908 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n14047) );
  INV_X1 U15909 ( .A(n14048), .ZN(P1_U3525) );
  MUX2_X1 U15910 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14049), .S(n14589), .Z(
        P1_U3524) );
  OAI21_X1 U15911 ( .B1(n14052), .B2(n14077), .A(n14051), .ZN(P1_U3523) );
  MUX2_X1 U15912 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14053), .S(n14589), .Z(
        P1_U3522) );
  MUX2_X1 U15913 ( .A(n15135), .B(n14054), .S(n14589), .Z(n14055) );
  OAI21_X1 U15914 ( .B1(n6945), .B2(n14077), .A(n14055), .ZN(P1_U3521) );
  INV_X1 U15915 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n14057) );
  MUX2_X1 U15916 ( .A(n14057), .B(n14056), .S(n14589), .Z(n14058) );
  OAI21_X1 U15917 ( .B1(n14059), .B2(n14077), .A(n14058), .ZN(P1_U3520) );
  MUX2_X1 U15918 ( .A(n14060), .B(P1_REG0_REG_23__SCAN_IN), .S(n6712), .Z(
        P1_U3519) );
  MUX2_X1 U15919 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14061), .S(n14589), .Z(
        n14062) );
  INV_X1 U15920 ( .A(n14062), .ZN(n14063) );
  OAI21_X1 U15921 ( .B1(n14077), .B2(n14064), .A(n14063), .ZN(P1_U3518) );
  INV_X1 U15922 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n14066) );
  MUX2_X1 U15923 ( .A(n14066), .B(n14065), .S(n14589), .Z(n14067) );
  OAI21_X1 U15924 ( .B1(n14068), .B2(n14077), .A(n14067), .ZN(P1_U3517) );
  MUX2_X1 U15925 ( .A(n14069), .B(P1_REG0_REG_20__SCAN_IN), .S(n6712), .Z(
        P1_U3516) );
  INV_X1 U15926 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n14071) );
  MUX2_X1 U15927 ( .A(n14071), .B(n14070), .S(n14589), .Z(n14072) );
  OAI21_X1 U15928 ( .B1(n14073), .B2(n14077), .A(n14072), .ZN(P1_U3515) );
  INV_X1 U15929 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n14075) );
  MUX2_X1 U15930 ( .A(n14075), .B(n14074), .S(n14589), .Z(n14076) );
  OAI21_X1 U15931 ( .B1(n6943), .B2(n14077), .A(n14076), .ZN(P1_U3513) );
  MUX2_X1 U15932 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14078), .S(n14589), .Z(
        P1_U3510) );
  NOR4_X1 U15933 ( .A1(n14079), .A2(P1_IR_REG_30__SCAN_IN), .A3(n8325), .A4(
        P1_U3086), .ZN(n14080) );
  AOI21_X1 U15934 ( .B1(n14081), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14080), 
        .ZN(n14082) );
  OAI21_X1 U15935 ( .B1(n14084), .B2(n14083), .A(n14082), .ZN(P1_U3324) );
  OAI222_X1 U15936 ( .A1(n8056), .A2(P1_U3086), .B1(n14088), .B2(n14087), .C1(
        n14086), .C2(n14085), .ZN(P1_U3326) );
  MUX2_X1 U15937 ( .A(n14090), .B(n14089), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U15938 ( .A(n14091), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U15939 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14715) );
  INV_X1 U15940 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14702) );
  INV_X1 U15941 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14464) );
  XOR2_X1 U15942 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n14464), .Z(n14118) );
  INV_X1 U15943 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14446) );
  NOR2_X1 U15944 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14446), .ZN(n14117) );
  INV_X1 U15945 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15149) );
  NOR2_X1 U15946 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n12367), .ZN(n14115) );
  INV_X1 U15947 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14121) );
  XNOR2_X1 U15948 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(n10190), .ZN(n14173) );
  XOR2_X1 U15949 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(n14112), .Z(n14124) );
  XOR2_X1 U15950 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(P3_ADDR_REG_9__SCAN_IN), .Z(
        n14163) );
  XOR2_X1 U15951 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n14107), .Z(n14128) );
  XOR2_X1 U15952 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n15168), .Z(n14131) );
  NAND2_X1 U15953 ( .A1(n14131), .A2(n14132), .ZN(n14092) );
  NAND2_X1 U15954 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14093), .ZN(n14094) );
  NAND2_X1 U15955 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14095), .ZN(n14097) );
  NAND2_X1 U15956 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14098), .ZN(n14100) );
  OR2_X1 U15957 ( .A1(n14150), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n14101) );
  INV_X1 U15958 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n14102) );
  NAND2_X1 U15959 ( .A1(n14103), .A2(n14102), .ZN(n14105) );
  XOR2_X1 U15960 ( .A(n14103), .B(n14102), .Z(n14154) );
  NAND2_X1 U15961 ( .A1(n14154), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14104) );
  NAND2_X1 U15962 ( .A1(n14105), .A2(n14104), .ZN(n14129) );
  NAND2_X1 U15963 ( .A1(n14128), .A2(n14129), .ZN(n14106) );
  XOR2_X1 U15964 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n14110), .Z(n14126) );
  NAND2_X1 U15965 ( .A1(n14127), .A2(n14126), .ZN(n14109) );
  NAND2_X1 U15966 ( .A1(n14124), .A2(n14125), .ZN(n14111) );
  INV_X1 U15967 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14421) );
  NOR2_X1 U15968 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14421), .ZN(n14114) );
  OAI22_X1 U15969 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14121), .B1(n14123), 
        .B2(n14114), .ZN(n14119) );
  OAI22_X1 U15970 ( .A1(P3_ADDR_REG_14__SCAN_IN), .A2(n15149), .B1(n14115), 
        .B2(n14119), .ZN(n14174) );
  INV_X1 U15971 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14116) );
  OAI22_X1 U15972 ( .A1(n14117), .A2(n14174), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n14116), .ZN(n14178) );
  XNOR2_X1 U15973 ( .A(n14118), .B(n14178), .ZN(n14405) );
  INV_X1 U15974 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15142) );
  XOR2_X1 U15975 ( .A(n15149), .B(P3_ADDR_REG_14__SCAN_IN), .Z(n14120) );
  XNOR2_X1 U15976 ( .A(n14120), .B(n14119), .ZN(n14397) );
  XNOR2_X1 U15977 ( .A(n14121), .B(P1_ADDR_REG_13__SCAN_IN), .ZN(n14122) );
  XNOR2_X1 U15978 ( .A(n14123), .B(n14122), .ZN(n14393) );
  XOR2_X1 U15979 ( .A(n14125), .B(n14124), .Z(n14171) );
  XOR2_X1 U15980 ( .A(n14127), .B(n14126), .Z(n14167) );
  XOR2_X1 U15981 ( .A(n14129), .B(n14128), .Z(n14159) );
  XNOR2_X1 U15982 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n14130), .ZN(n14142) );
  NOR2_X1 U15983 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14142), .ZN(n14144) );
  XNOR2_X1 U15984 ( .A(n14132), .B(n14131), .ZN(n14202) );
  NAND2_X1 U15985 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14136), .ZN(n14138) );
  AOI21_X1 U15986 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14135), .A(n14134), .ZN(
        n15199) );
  INV_X1 U15987 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15198) );
  NOR2_X1 U15988 ( .A1(n15199), .A2(n15198), .ZN(n15208) );
  NAND2_X1 U15989 ( .A1(n15208), .A2(n15207), .ZN(n14137) );
  XOR2_X1 U15990 ( .A(n14140), .B(n14139), .Z(n15204) );
  INV_X1 U15991 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15205) );
  NAND2_X1 U15992 ( .A1(n15203), .A2(n15204), .ZN(n15202) );
  OAI21_X1 U15993 ( .B1(n14141), .B2(n15205), .A(n15202), .ZN(n15195) );
  XNOR2_X1 U15994 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n14142), .ZN(n15194) );
  NOR2_X1 U15995 ( .A1(n15195), .A2(n15194), .ZN(n14143) );
  NAND2_X1 U15996 ( .A1(n14149), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14153) );
  INV_X1 U15997 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n14623) );
  XNOR2_X1 U15998 ( .A(n14149), .B(n14623), .ZN(n14212) );
  XOR2_X1 U15999 ( .A(n14150), .B(P3_ADDR_REG_6__SCAN_IN), .Z(n14152) );
  XNOR2_X1 U16000 ( .A(n14152), .B(n14151), .ZN(n14211) );
  NAND2_X1 U16001 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14155), .ZN(n14157) );
  XOR2_X1 U16002 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14154), .Z(n15201) );
  INV_X1 U16003 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14636) );
  NAND2_X1 U16004 ( .A1(n14157), .A2(n14156), .ZN(n14158) );
  NOR2_X1 U16005 ( .A1(n14159), .A2(n14158), .ZN(n14161) );
  XNOR2_X1 U16006 ( .A(n14159), .B(n14158), .ZN(n14226) );
  NOR2_X1 U16007 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n14226), .ZN(n14160) );
  XNOR2_X1 U16008 ( .A(n14163), .B(n14162), .ZN(n14165) );
  NAND2_X1 U16009 ( .A1(n14164), .A2(n14165), .ZN(n14166) );
  NOR2_X1 U16010 ( .A1(n14167), .A2(n14168), .ZN(n14229) );
  NOR2_X1 U16011 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n14228), .ZN(n14169) );
  NOR2_X1 U16012 ( .A1(n14171), .A2(n14170), .ZN(n14385) );
  XNOR2_X1 U16013 ( .A(n14173), .B(n14172), .ZN(n14389) );
  INV_X1 U16014 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14390) );
  INV_X1 U16015 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14667) );
  NAND2_X1 U16016 ( .A1(n14393), .A2(n14394), .ZN(n14392) );
  XOR2_X1 U16017 ( .A(n14446), .B(P3_ADDR_REG_15__SCAN_IN), .Z(n14175) );
  XOR2_X1 U16018 ( .A(n14175), .B(n14174), .Z(n14401) );
  INV_X1 U16019 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14690) );
  NAND2_X1 U16020 ( .A1(n14400), .A2(n14401), .ZN(n14399) );
  NAND2_X1 U16021 ( .A1(n14405), .A2(n14404), .ZN(n14177) );
  NOR2_X1 U16022 ( .A1(n14405), .A2(n14404), .ZN(n14403) );
  INV_X1 U16023 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14476) );
  AND2_X1 U16024 ( .A1(n14464), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n14179) );
  XOR2_X1 U16025 ( .A(n14476), .B(n14180), .Z(n14181) );
  XOR2_X1 U16026 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14181), .Z(n14248) );
  NOR2_X1 U16027 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14180), .ZN(n14184) );
  INV_X1 U16028 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14182) );
  NOR2_X1 U16029 ( .A1(n14182), .A2(n14181), .ZN(n14183) );
  NOR2_X1 U16030 ( .A1(n14184), .A2(n14183), .ZN(n14191) );
  INV_X1 U16031 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14192) );
  XNOR2_X1 U16032 ( .A(n14192), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(n14185) );
  XNOR2_X1 U16033 ( .A(n14191), .B(n14185), .ZN(n14186) );
  NOR2_X1 U16034 ( .A1(n14187), .A2(n14186), .ZN(n14188) );
  INV_X1 U16035 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14493) );
  NOR2_X1 U16036 ( .A1(P3_ADDR_REG_18__SCAN_IN), .A2(n14493), .ZN(n14190) );
  OAI22_X1 U16037 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n14192), .B1(n14191), 
        .B2(n14190), .ZN(n14195) );
  XNOR2_X1 U16038 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n14193) );
  XNOR2_X1 U16039 ( .A(n14193), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n14194) );
  XNOR2_X1 U16040 ( .A(n14195), .B(n14194), .ZN(n14196) );
  XNOR2_X1 U16041 ( .A(n14197), .B(n14196), .ZN(SUB_1596_U4) );
  INV_X1 U16042 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n14732) );
  XOR2_X1 U16043 ( .A(n14732), .B(n14198), .Z(SUB_1596_U62) );
  AOI21_X1 U16044 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14199) );
  OAI21_X1 U16045 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14199), 
        .ZN(U28) );
  AOI21_X1 U16046 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14200) );
  OAI21_X1 U16047 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14200), 
        .ZN(U29) );
  AOI21_X1 U16048 ( .B1(n14203), .B2(n14202), .A(n14201), .ZN(n14204) );
  XOR2_X1 U16049 ( .A(n14204), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  AOI22_X1 U16050 ( .A1(n14205), .A2(n14223), .B1(SI_9_), .B2(n14222), .ZN(
        n14206) );
  OAI21_X1 U16051 ( .B1(P3_U3151), .B2(n14207), .A(n14206), .ZN(P3_U3286) );
  INV_X1 U16052 ( .A(n14208), .ZN(n14209) );
  AOI22_X1 U16053 ( .A1(n14209), .A2(n14223), .B1(SI_11_), .B2(n14222), .ZN(
        n14210) );
  OAI21_X1 U16054 ( .B1(P3_U3151), .B2(n14899), .A(n14210), .ZN(P3_U3284) );
  XOR2_X1 U16055 ( .A(n14212), .B(n14211), .Z(SUB_1596_U57) );
  OAI22_X1 U16056 ( .A1(n14216), .A2(n14215), .B1(n14214), .B2(n14213), .ZN(
        n14217) );
  INV_X1 U16057 ( .A(n14217), .ZN(n14218) );
  OAI21_X1 U16058 ( .B1(P3_U3151), .B2(n14219), .A(n14218), .ZN(P3_U3281) );
  AOI22_X1 U16059 ( .A1(n14220), .A2(n14223), .B1(SI_15_), .B2(n14222), .ZN(
        n14221) );
  OAI21_X1 U16060 ( .B1(P3_U3151), .B2(n14266), .A(n14221), .ZN(P3_U3280) );
  AOI22_X1 U16061 ( .A1(n14224), .A2(n14223), .B1(SI_16_), .B2(n14222), .ZN(
        n14225) );
  OAI21_X1 U16062 ( .B1(P3_U3151), .B2(n14288), .A(n14225), .ZN(P3_U3279) );
  INV_X1 U16063 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14649) );
  XOR2_X1 U16064 ( .A(n14649), .B(n14226), .Z(SUB_1596_U55) );
  XOR2_X1 U16065 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14227), .Z(SUB_1596_U54) );
  NOR2_X1 U16066 ( .A1(n14229), .A2(n14228), .ZN(n14230) );
  XNOR2_X1 U16067 ( .A(n14231), .B(n14230), .ZN(SUB_1596_U70) );
  INV_X1 U16068 ( .A(n14233), .ZN(n14234) );
  NOR2_X1 U16069 ( .A1(n14235), .A2(n14234), .ZN(n14236) );
  AOI21_X1 U16070 ( .B1(n11633), .B2(n14236), .A(n14548), .ZN(n14238) );
  AOI21_X1 U16071 ( .B1(n14232), .B2(n14238), .A(n14237), .ZN(n14368) );
  INV_X1 U16072 ( .A(n14239), .ZN(n14240) );
  AOI222_X1 U16073 ( .A1(n14241), .A2(n14501), .B1(P1_REG2_REG_13__SCAN_IN), 
        .B2(n14545), .C1(n14240), .C2(n14542), .ZN(n14247) );
  XNOR2_X1 U16074 ( .A(n14242), .B(n14243), .ZN(n14371) );
  OAI211_X1 U16075 ( .C1(n14244), .C2(n14369), .A(n14508), .B(n6594), .ZN(
        n14367) );
  INV_X1 U16076 ( .A(n14367), .ZN(n14245) );
  AOI22_X1 U16077 ( .A1(n14371), .A2(n14512), .B1(n14511), .B2(n14245), .ZN(
        n14246) );
  OAI211_X1 U16078 ( .C1(n14545), .C2(n14368), .A(n14247), .B(n14246), .ZN(
        P1_U3280) );
  AOI21_X1 U16079 ( .B1(n14249), .B2(n6438), .A(n6577), .ZN(n14250) );
  XOR2_X1 U16080 ( .A(n14250), .B(P2_ADDR_REG_17__SCAN_IN), .Z(SUB_1596_U63)
         );
  XOR2_X1 U16081 ( .A(n14252), .B(n14251), .Z(n14258) );
  NAND2_X1 U16082 ( .A1(n14253), .A2(n14884), .ZN(n14254) );
  OAI211_X1 U16083 ( .C1(n14298), .C2(n14889), .A(n14255), .B(n14254), .ZN(
        n14256) );
  AOI21_X1 U16084 ( .B1(n14258), .B2(n14257), .A(n14256), .ZN(n14259) );
  OAI21_X1 U16085 ( .B1(n14260), .B2(n14893), .A(n14259), .ZN(P3_U3155) );
  AOI21_X1 U16086 ( .B1(n14263), .B2(n14262), .A(n14261), .ZN(n14278) );
  INV_X1 U16087 ( .A(n14264), .ZN(n14265) );
  OAI21_X1 U16088 ( .B1(n14917), .B2(n14266), .A(n14265), .ZN(n14276) );
  AOI21_X1 U16089 ( .B1(n14269), .B2(n14268), .A(n14267), .ZN(n14274) );
  AOI21_X1 U16090 ( .B1(n14272), .B2(n14271), .A(n14270), .ZN(n14273) );
  OAI22_X1 U16091 ( .A1(n14274), .A2(n14927), .B1(n14273), .B2(n14906), .ZN(
        n14275) );
  AOI211_X1 U16092 ( .C1(n14931), .C2(P3_ADDR_REG_15__SCAN_IN), .A(n14276), 
        .B(n14275), .ZN(n14277) );
  OAI21_X1 U16093 ( .B1(n14278), .B2(n14933), .A(n14277), .ZN(P3_U3197) );
  AOI21_X1 U16094 ( .B1(n14280), .B2(n14279), .A(n6529), .ZN(n14296) );
  INV_X1 U16095 ( .A(n14281), .ZN(n14283) );
  NAND2_X1 U16096 ( .A1(n14283), .A2(n14282), .ZN(n14284) );
  XNOR2_X1 U16097 ( .A(n14285), .B(n14284), .ZN(n14294) );
  NAND2_X1 U16098 ( .A1(n14931), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n14286) );
  OAI211_X1 U16099 ( .C1(n14917), .C2(n14288), .A(n14287), .B(n14286), .ZN(
        n14293) );
  AOI21_X1 U16100 ( .B1(n6533), .B2(n14290), .A(n14289), .ZN(n14291) );
  NOR2_X1 U16101 ( .A1(n14291), .A2(n14927), .ZN(n14292) );
  AOI211_X1 U16102 ( .C1(n14924), .C2(n14294), .A(n14293), .B(n14292), .ZN(
        n14295) );
  OAI21_X1 U16103 ( .B1(n14296), .B2(n14933), .A(n14295), .ZN(P3_U3198) );
  INV_X1 U16104 ( .A(n14297), .ZN(n14301) );
  OAI22_X1 U16105 ( .A1(n14299), .A2(n14304), .B1(n14298), .B2(n15001), .ZN(
        n14300) );
  NOR2_X1 U16106 ( .A1(n14301), .A2(n14300), .ZN(n14317) );
  INV_X1 U16107 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n14302) );
  AOI22_X1 U16108 ( .A1(n15034), .A2(n14317), .B1(n14302), .B2(n15039), .ZN(
        P3_U3473) );
  OAI22_X1 U16109 ( .A1(n14305), .A2(n14304), .B1(n14303), .B2(n15001), .ZN(
        n14307) );
  NOR2_X1 U16110 ( .A1(n14307), .A2(n14306), .ZN(n14319) );
  AOI22_X1 U16111 ( .A1(n15034), .A2(n14319), .B1(n14920), .B2(n15039), .ZN(
        P3_U3472) );
  AOI22_X1 U16112 ( .A1(n14309), .A2(n15007), .B1(n15014), .B2(n14308), .ZN(
        n14310) );
  AND2_X1 U16113 ( .A1(n14311), .A2(n14310), .ZN(n14321) );
  AOI22_X1 U16114 ( .A1(n15034), .A2(n14321), .B1(n15132), .B2(n15039), .ZN(
        P3_U3471) );
  AOI22_X1 U16115 ( .A1(n14313), .A2(n15007), .B1(n14312), .B2(n15014), .ZN(
        n14314) );
  AND2_X1 U16116 ( .A1(n14315), .A2(n14314), .ZN(n14323) );
  AOI22_X1 U16117 ( .A1(n15034), .A2(n14323), .B1(n14902), .B2(n15039), .ZN(
        P3_U3470) );
  INV_X1 U16118 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14316) );
  AOI22_X1 U16119 ( .A1(n15025), .A2(n14317), .B1(n14316), .B2(n15023), .ZN(
        P3_U3432) );
  INV_X1 U16120 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14318) );
  AOI22_X1 U16121 ( .A1(n15025), .A2(n14319), .B1(n14318), .B2(n15023), .ZN(
        P3_U3429) );
  INV_X1 U16122 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14320) );
  AOI22_X1 U16123 ( .A1(n15025), .A2(n14321), .B1(n14320), .B2(n15023), .ZN(
        P3_U3426) );
  INV_X1 U16124 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14322) );
  AOI22_X1 U16125 ( .A1(n15025), .A2(n14323), .B1(n14322), .B2(n15023), .ZN(
        P3_U3423) );
  OAI22_X1 U16126 ( .A1(n14327), .A2(n14326), .B1(n14325), .B2(n14324), .ZN(
        n14334) );
  NAND2_X1 U16127 ( .A1(n14329), .A2(n14328), .ZN(n14331) );
  AOI21_X1 U16128 ( .B1(n14332), .B2(n14331), .A(n14330), .ZN(n14333) );
  AOI211_X1 U16129 ( .C1(n14336), .C2(n14335), .A(n14334), .B(n14333), .ZN(
        n14337) );
  NAND2_X1 U16130 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14432)
         );
  OAI211_X1 U16131 ( .C1(n14339), .C2(n14338), .A(n14337), .B(n14432), .ZN(
        P1_U3215) );
  AOI21_X1 U16132 ( .B1(n6595), .B2(n14346), .A(n14548), .ZN(n14342) );
  AOI21_X1 U16133 ( .B1(n14342), .B2(n14341), .A(n14340), .ZN(n14375) );
  INV_X1 U16134 ( .A(n14343), .ZN(n14344) );
  AOI222_X1 U16135 ( .A1(n14373), .A2(n14501), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n14545), .C1(n14542), .C2(n14344), .ZN(n14353) );
  XNOR2_X1 U16136 ( .A(n14345), .B(n14346), .ZN(n14378) );
  NAND2_X1 U16137 ( .A1(n14347), .A2(n14373), .ZN(n14348) );
  NAND2_X1 U16138 ( .A1(n14348), .A2(n14508), .ZN(n14350) );
  OR2_X1 U16139 ( .A1(n14350), .A2(n14349), .ZN(n14374) );
  INV_X1 U16140 ( .A(n14374), .ZN(n14351) );
  AOI22_X1 U16141 ( .A1(n14378), .A2(n14512), .B1(n14511), .B2(n14351), .ZN(
        n14352) );
  OAI211_X1 U16142 ( .C1(n14545), .C2(n14375), .A(n14353), .B(n14352), .ZN(
        P1_U3282) );
  OAI21_X1 U16143 ( .B1(n14355), .B2(n14584), .A(n14354), .ZN(n14358) );
  INV_X1 U16144 ( .A(n14356), .ZN(n14357) );
  AOI211_X1 U16145 ( .C1(n14588), .C2(n14359), .A(n14358), .B(n14357), .ZN(
        n14379) );
  AOI22_X1 U16146 ( .A1(n14597), .A2(n14379), .B1(n8350), .B2(n14595), .ZN(
        P1_U3544) );
  AOI211_X1 U16147 ( .C1(n14362), .C2(n14574), .A(n14361), .B(n14360), .ZN(
        n14364) );
  OAI211_X1 U16148 ( .C1(n14365), .C2(n14549), .A(n14364), .B(n14363), .ZN(
        n14366) );
  INV_X1 U16149 ( .A(n14366), .ZN(n14380) );
  AOI22_X1 U16150 ( .A1(n14597), .A2(n14380), .B1(n14435), .B2(n14595), .ZN(
        P1_U3543) );
  OAI211_X1 U16151 ( .C1(n14369), .C2(n14584), .A(n14368), .B(n14367), .ZN(
        n14370) );
  AOI21_X1 U16152 ( .B1(n14588), .B2(n14371), .A(n14370), .ZN(n14381) );
  AOI22_X1 U16153 ( .A1(n14597), .A2(n14381), .B1(n14372), .B2(n14595), .ZN(
        P1_U3541) );
  INV_X1 U16154 ( .A(n14373), .ZN(n14376) );
  OAI211_X1 U16155 ( .C1(n14376), .C2(n14584), .A(n14375), .B(n14374), .ZN(
        n14377) );
  AOI21_X1 U16156 ( .B1(n14588), .B2(n14378), .A(n14377), .ZN(n14383) );
  AOI22_X1 U16157 ( .A1(n14597), .A2(n14383), .B1(n10187), .B2(n14595), .ZN(
        P1_U3539) );
  AOI22_X1 U16158 ( .A1(n14589), .A2(n14379), .B1(n8351), .B2(n6712), .ZN(
        P1_U3507) );
  AOI22_X1 U16159 ( .A1(n14589), .A2(n14380), .B1(n8331), .B2(n6712), .ZN(
        P1_U3504) );
  AOI22_X1 U16160 ( .A1(n14589), .A2(n14381), .B1(n8295), .B2(n6712), .ZN(
        P1_U3498) );
  INV_X1 U16161 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14382) );
  AOI22_X1 U16162 ( .A1(n14589), .A2(n14383), .B1(n14382), .B2(n6712), .ZN(
        P1_U3492) );
  NOR2_X1 U16163 ( .A1(n14385), .A2(n14384), .ZN(n14386) );
  XOR2_X1 U16164 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n14386), .Z(SUB_1596_U69)
         );
  OAI21_X1 U16165 ( .B1(n14389), .B2(n14388), .A(n14387), .ZN(n14391) );
  XOR2_X1 U16166 ( .A(n14391), .B(n14390), .Z(SUB_1596_U68) );
  OAI21_X1 U16167 ( .B1(n14394), .B2(n14393), .A(n14392), .ZN(n14395) );
  XOR2_X1 U16168 ( .A(n14395), .B(n14667), .Z(SUB_1596_U67) );
  AOI21_X1 U16169 ( .B1(n14397), .B2(n14396), .A(n6589), .ZN(n14398) );
  XOR2_X1 U16170 ( .A(n14398), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  OAI21_X1 U16171 ( .B1(n14401), .B2(n14400), .A(n14399), .ZN(n14402) );
  XOR2_X1 U16172 ( .A(n14402), .B(n14690), .Z(SUB_1596_U65) );
  AOI21_X1 U16173 ( .B1(n14405), .B2(n14404), .A(n14403), .ZN(n14406) );
  XOR2_X1 U16174 ( .A(n14406), .B(P2_ADDR_REG_16__SCAN_IN), .Z(SUB_1596_U64)
         );
  INV_X1 U16175 ( .A(n14489), .ZN(n14460) );
  INV_X1 U16176 ( .A(n14407), .ZN(n14408) );
  OAI211_X1 U16177 ( .C1(n14410), .C2(n14409), .A(n14408), .B(n14442), .ZN(
        n14416) );
  INV_X1 U16178 ( .A(n14411), .ZN(n14412) );
  OAI211_X1 U16179 ( .C1(n14414), .C2(n14413), .A(n14412), .B(n14440), .ZN(
        n14415) );
  OAI211_X1 U16180 ( .C1(n14460), .C2(n14417), .A(n14416), .B(n14415), .ZN(
        n14418) );
  INV_X1 U16181 ( .A(n14418), .ZN(n14420) );
  OAI211_X1 U16182 ( .C1(n14421), .C2(n14492), .A(n14420), .B(n14419), .ZN(
        P1_U3256) );
  OAI21_X1 U16183 ( .B1(n14424), .B2(n14423), .A(n14422), .ZN(n14431) );
  NOR2_X1 U16184 ( .A1(n14460), .A2(n14425), .ZN(n14430) );
  AOI211_X1 U16185 ( .C1(n14428), .C2(n14427), .A(n14426), .B(n14478), .ZN(
        n14429) );
  AOI211_X1 U16186 ( .C1(n14431), .C2(n14442), .A(n14430), .B(n14429), .ZN(
        n14433) );
  OAI211_X1 U16187 ( .C1(n15149), .C2(n14492), .A(n14433), .B(n14432), .ZN(
        P1_U3257) );
  OAI21_X1 U16188 ( .B1(n14436), .B2(n14435), .A(n14434), .ZN(n14443) );
  OAI21_X1 U16189 ( .B1(n14439), .B2(n11770), .A(n14438), .ZN(n14441) );
  AOI222_X1 U16190 ( .A1(n14443), .A2(n14442), .B1(n6621), .B2(n14489), .C1(
        n14441), .C2(n14440), .ZN(n14445) );
  OAI211_X1 U16191 ( .C1(n14446), .C2(n14492), .A(n14445), .B(n14444), .ZN(
        P1_U3258) );
  NAND2_X1 U16192 ( .A1(n14448), .A2(n14447), .ZN(n14451) );
  NOR2_X1 U16193 ( .A1(n14478), .A2(n14449), .ZN(n14450) );
  NAND2_X1 U16194 ( .A1(n14451), .A2(n14450), .ZN(n14458) );
  NAND2_X1 U16195 ( .A1(n14453), .A2(n14452), .ZN(n14456) );
  NOR2_X1 U16196 ( .A1(n14482), .A2(n14454), .ZN(n14455) );
  NAND2_X1 U16197 ( .A1(n14456), .A2(n14455), .ZN(n14457) );
  OAI211_X1 U16198 ( .C1(n14460), .C2(n14459), .A(n14458), .B(n14457), .ZN(
        n14461) );
  INV_X1 U16199 ( .A(n14461), .ZN(n14463) );
  OAI211_X1 U16200 ( .C1(n14464), .C2(n14492), .A(n14463), .B(n14462), .ZN(
        P1_U3259) );
  AOI211_X1 U16201 ( .C1(n14467), .C2(n14466), .A(n14465), .B(n14478), .ZN(
        n14472) );
  AOI211_X1 U16202 ( .C1(n14470), .C2(n14469), .A(n14468), .B(n14482), .ZN(
        n14471) );
  AOI211_X1 U16203 ( .C1(n14489), .C2(n14473), .A(n14472), .B(n14471), .ZN(
        n14475) );
  OAI211_X1 U16204 ( .C1(n14476), .C2(n14492), .A(n14475), .B(n14474), .ZN(
        P1_U3260) );
  INV_X1 U16205 ( .A(n14477), .ZN(n14488) );
  AOI211_X1 U16206 ( .C1(n14481), .C2(n14480), .A(n14479), .B(n14478), .ZN(
        n14487) );
  AOI211_X1 U16207 ( .C1(n14485), .C2(n14484), .A(n14483), .B(n14482), .ZN(
        n14486) );
  AOI211_X1 U16208 ( .C1(n14489), .C2(n14488), .A(n14487), .B(n14486), .ZN(
        n14491) );
  OAI211_X1 U16209 ( .C1(n14493), .C2(n14492), .A(n14491), .B(n14490), .ZN(
        P1_U3261) );
  AOI21_X1 U16210 ( .B1(n14494), .B2(n14504), .A(n14548), .ZN(n14498) );
  INV_X1 U16211 ( .A(n14495), .ZN(n14496) );
  AOI21_X1 U16212 ( .B1(n14498), .B2(n14497), .A(n14496), .ZN(n14583) );
  INV_X1 U16213 ( .A(n14499), .ZN(n14500) );
  AOI222_X1 U16214 ( .A1(n14502), .A2(n14501), .B1(P1_REG2_REG_10__SCAN_IN), 
        .B2(n14545), .C1(n14500), .C2(n14542), .ZN(n14514) );
  XNOR2_X1 U16215 ( .A(n14503), .B(n14504), .ZN(n14587) );
  XNOR2_X1 U16216 ( .A(n14505), .B(n14585), .ZN(n14509) );
  AOI22_X1 U16217 ( .A1(n14509), .A2(n14508), .B1(n14507), .B2(n14506), .ZN(
        n14582) );
  INV_X1 U16218 ( .A(n14582), .ZN(n14510) );
  AOI22_X1 U16219 ( .A1(n14587), .A2(n14512), .B1(n14511), .B2(n14510), .ZN(
        n14513) );
  OAI211_X1 U16220 ( .C1(n14545), .C2(n14583), .A(n14514), .B(n14513), .ZN(
        P1_U3283) );
  XNOR2_X1 U16221 ( .A(n10397), .B(n14515), .ZN(n14525) );
  OAI21_X1 U16222 ( .B1(n10397), .B2(n14516), .A(n14519), .ZN(n14522) );
  OAI21_X1 U16223 ( .B1(n14556), .B2(n14535), .A(n14517), .ZN(n14527) );
  XNOR2_X1 U16224 ( .A(n14527), .B(n8100), .ZN(n14520) );
  AOI21_X1 U16225 ( .B1(n14520), .B2(n14519), .A(n14518), .ZN(n14521) );
  AOI21_X1 U16226 ( .B1(n14523), .B2(n14522), .A(n14521), .ZN(n14524) );
  AOI21_X1 U16227 ( .B1(n14588), .B2(n14525), .A(n14524), .ZN(n14555) );
  NOR2_X1 U16228 ( .A1(n14527), .A2(n14526), .ZN(n14558) );
  NOR2_X1 U16229 ( .A1(n14556), .A2(n14528), .ZN(n14530) );
  NOR2_X1 U16230 ( .A1(n14529), .A2(n14533), .ZN(n14559) );
  AOI211_X1 U16231 ( .C1(n14558), .C2(n14536), .A(n14530), .B(n14559), .ZN(
        n14532) );
  AOI22_X1 U16232 ( .A1(n14542), .A2(P1_REG3_REG_1__SCAN_IN), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(n14545), .ZN(n14531) );
  OAI221_X1 U16233 ( .B1(n14545), .B2(n14555), .C1(n14545), .C2(n14532), .A(
        n14531), .ZN(P1_U3292) );
  NOR2_X1 U16234 ( .A1(n10398), .A2(n14533), .ZN(n14550) );
  INV_X1 U16235 ( .A(n14550), .ZN(n14540) );
  NAND3_X1 U16236 ( .A1(n14553), .A2(n10041), .A3(n14534), .ZN(n14539) );
  NOR2_X1 U16237 ( .A1(n14535), .A2(n10041), .ZN(n14551) );
  OAI21_X1 U16238 ( .B1(n14537), .B2(n14536), .A(n14551), .ZN(n14538) );
  NAND3_X1 U16239 ( .A1(n14540), .A2(n14539), .A3(n14538), .ZN(n14541) );
  AOI21_X1 U16240 ( .B1(n14542), .B2(P1_REG3_REG_0__SCAN_IN), .A(n14541), .ZN(
        n14544) );
  AOI22_X1 U16241 ( .A1(n14545), .A2(n8057), .B1(n14544), .B2(n14543), .ZN(
        P1_U3293) );
  AND2_X1 U16242 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14546), .ZN(P1_U3294) );
  AND2_X1 U16243 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14546), .ZN(P1_U3295) );
  AND2_X1 U16244 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14546), .ZN(P1_U3296) );
  AND2_X1 U16245 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14546), .ZN(P1_U3297) );
  AND2_X1 U16246 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14546), .ZN(P1_U3298) );
  AND2_X1 U16247 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14546), .ZN(P1_U3299) );
  AND2_X1 U16248 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14546), .ZN(P1_U3300) );
  AND2_X1 U16249 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14546), .ZN(P1_U3301) );
  AND2_X1 U16250 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14546), .ZN(P1_U3302) );
  AND2_X1 U16251 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14546), .ZN(P1_U3303) );
  AND2_X1 U16252 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14546), .ZN(P1_U3304) );
  AND2_X1 U16253 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14546), .ZN(P1_U3305) );
  INV_X1 U16254 ( .A(n14546), .ZN(n14547) );
  INV_X1 U16255 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n15099) );
  NOR2_X1 U16256 ( .A1(n14547), .A2(n15099), .ZN(P1_U3306) );
  AND2_X1 U16257 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14546), .ZN(P1_U3307) );
  AND2_X1 U16258 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14546), .ZN(P1_U3308) );
  AND2_X1 U16259 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14546), .ZN(P1_U3309) );
  AND2_X1 U16260 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14546), .ZN(P1_U3310) );
  AND2_X1 U16261 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14546), .ZN(P1_U3311) );
  AND2_X1 U16262 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14546), .ZN(P1_U3312) );
  AND2_X1 U16263 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14546), .ZN(P1_U3313) );
  AND2_X1 U16264 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14546), .ZN(P1_U3314) );
  AND2_X1 U16265 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14546), .ZN(P1_U3315) );
  AND2_X1 U16266 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14546), .ZN(P1_U3316) );
  AND2_X1 U16267 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14546), .ZN(P1_U3317) );
  AND2_X1 U16268 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14546), .ZN(P1_U3318) );
  AND2_X1 U16269 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14546), .ZN(P1_U3319) );
  AND2_X1 U16270 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14546), .ZN(P1_U3320) );
  AND2_X1 U16271 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14546), .ZN(P1_U3321) );
  AND2_X1 U16272 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14546), .ZN(P1_U3322) );
  INV_X1 U16273 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15131) );
  NOR2_X1 U16274 ( .A1(n14547), .A2(n15131), .ZN(P1_U3323) );
  NAND2_X1 U16275 ( .A1(n14549), .A2(n14548), .ZN(n14552) );
  AOI211_X1 U16276 ( .C1(n14553), .C2(n14552), .A(n14551), .B(n14550), .ZN(
        n14590) );
  INV_X1 U16277 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n14554) );
  AOI22_X1 U16278 ( .A1(n14589), .A2(n14590), .B1(n14554), .B2(n6712), .ZN(
        P1_U3459) );
  INV_X1 U16279 ( .A(n14555), .ZN(n14560) );
  NOR2_X1 U16280 ( .A1(n14584), .A2(n14556), .ZN(n14557) );
  NOR4_X1 U16281 ( .A1(n14560), .A2(n14559), .A3(n14558), .A4(n14557), .ZN(
        n14591) );
  INV_X1 U16282 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14561) );
  AOI22_X1 U16283 ( .A1(n14589), .A2(n14591), .B1(n14561), .B2(n6712), .ZN(
        P1_U3462) );
  OAI211_X1 U16284 ( .C1(n14564), .C2(n14584), .A(n14563), .B(n14562), .ZN(
        n14565) );
  AOI21_X1 U16285 ( .B1(n14588), .B2(n14566), .A(n14565), .ZN(n14592) );
  INV_X1 U16286 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14567) );
  AOI22_X1 U16287 ( .A1(n14589), .A2(n14592), .B1(n14567), .B2(n6712), .ZN(
        P1_U3465) );
  OAI21_X1 U16288 ( .B1(n14569), .B2(n14584), .A(n14568), .ZN(n14571) );
  AOI211_X1 U16289 ( .C1(n14588), .C2(n14572), .A(n14571), .B(n14570), .ZN(
        n14593) );
  AOI22_X1 U16290 ( .A1(n14589), .A2(n14593), .B1(n8137), .B2(n6712), .ZN(
        P1_U3471) );
  AOI21_X1 U16291 ( .B1(n14575), .B2(n14574), .A(n14573), .ZN(n14577) );
  NAND3_X1 U16292 ( .A1(n14578), .A2(n14577), .A3(n14576), .ZN(n14579) );
  AOI21_X1 U16293 ( .B1(n14588), .B2(n14580), .A(n14579), .ZN(n14594) );
  INV_X1 U16294 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14581) );
  AOI22_X1 U16295 ( .A1(n14589), .A2(n14594), .B1(n14581), .B2(n6712), .ZN(
        P1_U3483) );
  OAI211_X1 U16296 ( .C1(n14585), .C2(n14584), .A(n14583), .B(n14582), .ZN(
        n14586) );
  AOI21_X1 U16297 ( .B1(n14588), .B2(n14587), .A(n14586), .ZN(n14596) );
  AOI22_X1 U16298 ( .A1(n14589), .A2(n14596), .B1(n8239), .B2(n6712), .ZN(
        P1_U3489) );
  AOI22_X1 U16299 ( .A1(n14597), .A2(n14590), .B1(n8055), .B2(n14595), .ZN(
        P1_U3528) );
  AOI22_X1 U16300 ( .A1(n14597), .A2(n14591), .B1(n8072), .B2(n14595), .ZN(
        P1_U3529) );
  AOI22_X1 U16301 ( .A1(n14597), .A2(n14592), .B1(n8109), .B2(n14595), .ZN(
        P1_U3530) );
  AOI22_X1 U16302 ( .A1(n14597), .A2(n14593), .B1(n9933), .B2(n14595), .ZN(
        P1_U3532) );
  AOI22_X1 U16303 ( .A1(n14597), .A2(n14594), .B1(n9937), .B2(n14595), .ZN(
        P1_U3536) );
  AOI22_X1 U16304 ( .A1(n14597), .A2(n14596), .B1(n9939), .B2(n14595), .ZN(
        P1_U3538) );
  NOR2_X1 U16305 ( .A1(n14598), .A2(P2_U3947), .ZN(P2_U3087) );
  OAI211_X1 U16306 ( .C1(n14601), .C2(n14600), .A(n14724), .B(n14599), .ZN(
        n14606) );
  OAI211_X1 U16307 ( .C1(n14604), .C2(n14603), .A(n14657), .B(n14602), .ZN(
        n14605) );
  NAND2_X1 U16308 ( .A1(n14606), .A2(n14605), .ZN(n14607) );
  AOI21_X1 U16309 ( .B1(n14608), .B2(n14728), .A(n14607), .ZN(n14610) );
  NAND2_X1 U16310 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n14609) );
  OAI211_X1 U16311 ( .C1(n14731), .C2(n15205), .A(n14610), .B(n14609), .ZN(
        P2_U3217) );
  OAI211_X1 U16312 ( .C1(n14613), .C2(n14612), .A(n14657), .B(n14611), .ZN(
        n14618) );
  OAI211_X1 U16313 ( .C1(n14616), .C2(n14615), .A(n14724), .B(n14614), .ZN(
        n14617) );
  OAI211_X1 U16314 ( .C1(n14659), .C2(n14619), .A(n14618), .B(n14617), .ZN(
        n14620) );
  INV_X1 U16315 ( .A(n14620), .ZN(n14622) );
  OAI211_X1 U16316 ( .C1(n14731), .C2(n14623), .A(n14622), .B(n14621), .ZN(
        P2_U3220) );
  OAI211_X1 U16317 ( .C1(n14626), .C2(n14625), .A(n14657), .B(n14624), .ZN(
        n14631) );
  OAI211_X1 U16318 ( .C1(n14629), .C2(n14628), .A(n14724), .B(n14627), .ZN(
        n14630) );
  OAI211_X1 U16319 ( .C1(n14659), .C2(n14632), .A(n14631), .B(n14630), .ZN(
        n14633) );
  INV_X1 U16320 ( .A(n14633), .ZN(n14635) );
  OAI211_X1 U16321 ( .C1(n14636), .C2(n14731), .A(n14635), .B(n14634), .ZN(
        P2_U3221) );
  OAI211_X1 U16322 ( .C1(n14639), .C2(n14638), .A(n14724), .B(n14637), .ZN(
        n14644) );
  OAI211_X1 U16323 ( .C1(n14642), .C2(n14641), .A(n14657), .B(n14640), .ZN(
        n14643) );
  OAI211_X1 U16324 ( .C1(n14659), .C2(n14645), .A(n14644), .B(n14643), .ZN(
        n14646) );
  INV_X1 U16325 ( .A(n14646), .ZN(n14648) );
  NAND2_X1 U16326 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n14647) );
  OAI211_X1 U16327 ( .C1(n14649), .C2(n14731), .A(n14648), .B(n14647), .ZN(
        P2_U3222) );
  NAND2_X1 U16328 ( .A1(n14651), .A2(n14650), .ZN(n14652) );
  NAND2_X1 U16329 ( .A1(n14652), .A2(n14724), .ZN(n14653) );
  NOR2_X1 U16330 ( .A1(n14654), .A2(n14653), .ZN(n14664) );
  NAND2_X1 U16331 ( .A1(n14656), .A2(n14655), .ZN(n14658) );
  NAND2_X1 U16332 ( .A1(n14658), .A2(n14657), .ZN(n14661) );
  OAI22_X1 U16333 ( .A1(n14662), .A2(n14661), .B1(n14660), .B2(n14659), .ZN(
        n14663) );
  NOR2_X1 U16334 ( .A1(n14664), .A2(n14663), .ZN(n14666) );
  NAND2_X1 U16335 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n14665)
         );
  OAI211_X1 U16336 ( .C1(n14667), .C2(n14731), .A(n14666), .B(n14665), .ZN(
        P2_U3227) );
  AOI211_X1 U16337 ( .C1(n14669), .C2(n15134), .A(n14668), .B(n14706), .ZN(
        n14674) );
  AOI211_X1 U16338 ( .C1(n14672), .C2(n14671), .A(n14670), .B(n14716), .ZN(
        n14673) );
  AOI211_X1 U16339 ( .C1(n14728), .C2(n14675), .A(n14674), .B(n14673), .ZN(
        n14677) );
  NAND2_X1 U16340 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14676)
         );
  OAI211_X1 U16341 ( .C1(n15142), .C2(n14731), .A(n14677), .B(n14676), .ZN(
        P2_U3228) );
  INV_X1 U16342 ( .A(n14678), .ZN(n14687) );
  AOI211_X1 U16343 ( .C1(n14681), .C2(n14680), .A(n14679), .B(n14716), .ZN(
        n14686) );
  AOI211_X1 U16344 ( .C1(n14684), .C2(n14683), .A(n14682), .B(n14706), .ZN(
        n14685) );
  AOI211_X1 U16345 ( .C1(n14728), .C2(n14687), .A(n14686), .B(n14685), .ZN(
        n14689) );
  NAND2_X1 U16346 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n14688)
         );
  OAI211_X1 U16347 ( .C1(n14690), .C2(n14731), .A(n14689), .B(n14688), .ZN(
        P2_U3229) );
  AOI211_X1 U16348 ( .C1(n14693), .C2(n14692), .A(n14691), .B(n14716), .ZN(
        n14698) );
  AOI211_X1 U16349 ( .C1(n14696), .C2(n14695), .A(n14694), .B(n14706), .ZN(
        n14697) );
  AOI211_X1 U16350 ( .C1(n14728), .C2(n14699), .A(n14698), .B(n14697), .ZN(
        n14701) );
  NAND2_X1 U16351 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n14700)
         );
  OAI211_X1 U16352 ( .C1(n14702), .C2(n14731), .A(n14701), .B(n14700), .ZN(
        P2_U3230) );
  AOI211_X1 U16353 ( .C1(n14705), .C2(n14704), .A(n14703), .B(n14716), .ZN(
        n14711) );
  AOI211_X1 U16354 ( .C1(n14709), .C2(n14708), .A(n14707), .B(n14706), .ZN(
        n14710) );
  AOI211_X1 U16355 ( .C1(n14728), .C2(n14712), .A(n14711), .B(n14710), .ZN(
        n14714) );
  NAND2_X1 U16356 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3088), .ZN(n14713)
         );
  OAI211_X1 U16357 ( .C1(n14715), .C2(n14731), .A(n14714), .B(n14713), .ZN(
        P2_U3231) );
  AOI211_X1 U16358 ( .C1(n14719), .C2(n14718), .A(n14717), .B(n14716), .ZN(
        n14726) );
  OAI21_X1 U16359 ( .B1(n14722), .B2(n14721), .A(n14720), .ZN(n14723) );
  AND2_X1 U16360 ( .A1(n14724), .A2(n14723), .ZN(n14725) );
  AOI211_X1 U16361 ( .C1(n14728), .C2(n14727), .A(n14726), .B(n14725), .ZN(
        n14730) );
  OAI211_X1 U16362 ( .C1(n14732), .C2(n14731), .A(n14730), .B(n14729), .ZN(
        P2_U3232) );
  CLKBUF_X1 U16363 ( .A(n14757), .Z(n14761) );
  NOR2_X1 U16364 ( .A1(n14761), .A2(n15159), .ZN(P2_U3266) );
  INV_X1 U16365 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n14734) );
  NOR2_X1 U16366 ( .A1(n14761), .A2(n14734), .ZN(P2_U3267) );
  INV_X1 U16367 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n14735) );
  NOR2_X1 U16368 ( .A1(n14761), .A2(n14735), .ZN(P2_U3268) );
  INV_X1 U16369 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n14736) );
  NOR2_X1 U16370 ( .A1(n14757), .A2(n14736), .ZN(P2_U3269) );
  INV_X1 U16371 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n14737) );
  NOR2_X1 U16372 ( .A1(n14757), .A2(n14737), .ZN(P2_U3270) );
  INV_X1 U16373 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n14738) );
  NOR2_X1 U16374 ( .A1(n14757), .A2(n14738), .ZN(P2_U3271) );
  INV_X1 U16375 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n14739) );
  NOR2_X1 U16376 ( .A1(n14757), .A2(n14739), .ZN(P2_U3272) );
  NOR2_X1 U16377 ( .A1(n14757), .A2(n15169), .ZN(P2_U3273) );
  INV_X1 U16378 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n14740) );
  NOR2_X1 U16379 ( .A1(n14757), .A2(n14740), .ZN(P2_U3274) );
  INV_X1 U16380 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n14741) );
  NOR2_X1 U16381 ( .A1(n14757), .A2(n14741), .ZN(P2_U3275) );
  NOR2_X1 U16382 ( .A1(n14757), .A2(n15141), .ZN(P2_U3276) );
  INV_X1 U16383 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n14742) );
  NOR2_X1 U16384 ( .A1(n14757), .A2(n14742), .ZN(P2_U3277) );
  INV_X1 U16385 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n14743) );
  NOR2_X1 U16386 ( .A1(n14761), .A2(n14743), .ZN(P2_U3278) );
  INV_X1 U16387 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n14744) );
  NOR2_X1 U16388 ( .A1(n14761), .A2(n14744), .ZN(P2_U3279) );
  INV_X1 U16389 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n14745) );
  NOR2_X1 U16390 ( .A1(n14761), .A2(n14745), .ZN(P2_U3280) );
  INV_X1 U16391 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n14746) );
  NOR2_X1 U16392 ( .A1(n14761), .A2(n14746), .ZN(P2_U3281) );
  INV_X1 U16393 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n14747) );
  NOR2_X1 U16394 ( .A1(n14761), .A2(n14747), .ZN(P2_U3282) );
  INV_X1 U16395 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n14748) );
  NOR2_X1 U16396 ( .A1(n14761), .A2(n14748), .ZN(P2_U3283) );
  NOR2_X1 U16397 ( .A1(n14761), .A2(n15126), .ZN(P2_U3284) );
  INV_X1 U16398 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n14749) );
  NOR2_X1 U16399 ( .A1(n14761), .A2(n14749), .ZN(P2_U3285) );
  INV_X1 U16400 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n14750) );
  NOR2_X1 U16401 ( .A1(n14761), .A2(n14750), .ZN(P2_U3286) );
  INV_X1 U16402 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n14751) );
  NOR2_X1 U16403 ( .A1(n14761), .A2(n14751), .ZN(P2_U3287) );
  INV_X1 U16404 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n14752) );
  NOR2_X1 U16405 ( .A1(n14761), .A2(n14752), .ZN(P2_U3288) );
  INV_X1 U16406 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n14753) );
  NOR2_X1 U16407 ( .A1(n14761), .A2(n14753), .ZN(P2_U3289) );
  INV_X1 U16408 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n14754) );
  NOR2_X1 U16409 ( .A1(n14757), .A2(n14754), .ZN(P2_U3290) );
  INV_X1 U16410 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n14755) );
  NOR2_X1 U16411 ( .A1(n14761), .A2(n14755), .ZN(P2_U3291) );
  INV_X1 U16412 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n14756) );
  NOR2_X1 U16413 ( .A1(n14757), .A2(n14756), .ZN(P2_U3292) );
  INV_X1 U16414 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n14758) );
  NOR2_X1 U16415 ( .A1(n14761), .A2(n14758), .ZN(P2_U3293) );
  INV_X1 U16416 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n14759) );
  NOR2_X1 U16417 ( .A1(n14761), .A2(n14759), .ZN(P2_U3294) );
  INV_X1 U16418 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n14760) );
  NOR2_X1 U16419 ( .A1(n14761), .A2(n14760), .ZN(P2_U3295) );
  AOI22_X1 U16420 ( .A1(n14767), .A2(n14763), .B1(n14762), .B2(n14764), .ZN(
        P2_U3416) );
  AOI22_X1 U16421 ( .A1(n14767), .A2(n14766), .B1(n14765), .B2(n14764), .ZN(
        P2_U3417) );
  NOR2_X1 U16422 ( .A1(n14768), .A2(n14838), .ZN(n14771) );
  INV_X1 U16423 ( .A(n14769), .ZN(n14770) );
  AOI211_X1 U16424 ( .C1(n14773), .C2(n14772), .A(n14771), .B(n14770), .ZN(
        n14859) );
  INV_X1 U16425 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14774) );
  AOI22_X1 U16426 ( .A1(n14858), .A2(n14859), .B1(n14774), .B2(n14856), .ZN(
        P2_U3430) );
  INV_X1 U16427 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15095) );
  AOI22_X1 U16428 ( .A1(n14858), .A2(n14775), .B1(n15095), .B2(n14856), .ZN(
        P2_U3433) );
  INV_X1 U16429 ( .A(n14776), .ZN(n14782) );
  NOR2_X1 U16430 ( .A1(n14776), .A2(n14838), .ZN(n14781) );
  OAI211_X1 U16431 ( .C1(n14779), .C2(n14852), .A(n14778), .B(n14777), .ZN(
        n14780) );
  AOI211_X1 U16432 ( .C1(n14836), .C2(n14782), .A(n14781), .B(n14780), .ZN(
        n14860) );
  INV_X1 U16433 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14783) );
  AOI22_X1 U16434 ( .A1(n14858), .A2(n14860), .B1(n14783), .B2(n14856), .ZN(
        P2_U3436) );
  AOI21_X1 U16435 ( .B1(n14841), .B2(n14785), .A(n14784), .ZN(n14786) );
  OAI211_X1 U16436 ( .C1(n14798), .C2(n14788), .A(n14787), .B(n14786), .ZN(
        n14789) );
  INV_X1 U16437 ( .A(n14789), .ZN(n14861) );
  INV_X1 U16438 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14790) );
  AOI22_X1 U16439 ( .A1(n14858), .A2(n14861), .B1(n14790), .B2(n14856), .ZN(
        P2_U3439) );
  AOI211_X1 U16440 ( .C1(n14841), .C2(n14793), .A(n14792), .B(n14791), .ZN(
        n14794) );
  OAI21_X1 U16441 ( .B1(n14798), .B2(n14795), .A(n14794), .ZN(n14796) );
  INV_X1 U16442 ( .A(n14796), .ZN(n14862) );
  INV_X1 U16443 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14797) );
  AOI22_X1 U16444 ( .A1(n14858), .A2(n14862), .B1(n14797), .B2(n14856), .ZN(
        P2_U3442) );
  NOR2_X1 U16445 ( .A1(n14799), .A2(n14798), .ZN(n14804) );
  OAI21_X1 U16446 ( .B1(n14801), .B2(n14852), .A(n14800), .ZN(n14802) );
  NOR3_X1 U16447 ( .A1(n14804), .A2(n14803), .A3(n14802), .ZN(n14863) );
  INV_X1 U16448 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14805) );
  AOI22_X1 U16449 ( .A1(n14858), .A2(n14863), .B1(n14805), .B2(n14856), .ZN(
        P2_U3445) );
  AND2_X1 U16450 ( .A1(n14806), .A2(n8001), .ZN(n14810) );
  OAI21_X1 U16451 ( .B1(n14808), .B2(n14852), .A(n14807), .ZN(n14809) );
  NOR3_X1 U16452 ( .A1(n14811), .A2(n14810), .A3(n14809), .ZN(n14865) );
  INV_X1 U16453 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n14812) );
  AOI22_X1 U16454 ( .A1(n14858), .A2(n14865), .B1(n14812), .B2(n14856), .ZN(
        P2_U3448) );
  INV_X1 U16455 ( .A(n14813), .ZN(n14814) );
  OAI21_X1 U16456 ( .B1(n14815), .B2(n14852), .A(n14814), .ZN(n14818) );
  INV_X1 U16457 ( .A(n14816), .ZN(n14817) );
  AOI211_X1 U16458 ( .C1(n14819), .C2(n8001), .A(n14818), .B(n14817), .ZN(
        n14867) );
  INV_X1 U16459 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n14820) );
  AOI22_X1 U16460 ( .A1(n14858), .A2(n14867), .B1(n14820), .B2(n14856), .ZN(
        P2_U3451) );
  OAI21_X1 U16461 ( .B1(n14822), .B2(n14852), .A(n14821), .ZN(n14826) );
  NOR2_X1 U16462 ( .A1(n14823), .A2(n14838), .ZN(n14825) );
  NOR2_X1 U16463 ( .A1(n14823), .A2(n14839), .ZN(n14824) );
  NOR4_X1 U16464 ( .A1(n14827), .A2(n14826), .A3(n14825), .A4(n14824), .ZN(
        n14869) );
  INV_X1 U16465 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14828) );
  AOI22_X1 U16466 ( .A1(n14858), .A2(n14869), .B1(n14828), .B2(n14856), .ZN(
        P2_U3454) );
  NAND2_X1 U16467 ( .A1(n14829), .A2(n14841), .ZN(n14831) );
  OAI211_X1 U16468 ( .C1(n14832), .C2(n14838), .A(n14831), .B(n14830), .ZN(
        n14833) );
  AOI211_X1 U16469 ( .C1(n14836), .C2(n14835), .A(n14834), .B(n14833), .ZN(
        n14871) );
  INV_X1 U16470 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n14837) );
  AOI22_X1 U16471 ( .A1(n14858), .A2(n14871), .B1(n14837), .B2(n14856), .ZN(
        P2_U3457) );
  NOR2_X1 U16472 ( .A1(n14840), .A2(n14838), .ZN(n14848) );
  NOR2_X1 U16473 ( .A1(n14840), .A2(n14839), .ZN(n14847) );
  NAND2_X1 U16474 ( .A1(n14842), .A2(n14841), .ZN(n14843) );
  NAND2_X1 U16475 ( .A1(n14844), .A2(n14843), .ZN(n14845) );
  NOR4_X1 U16476 ( .A1(n14848), .A2(n14847), .A3(n14846), .A4(n14845), .ZN(
        n14872) );
  INV_X1 U16477 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14849) );
  AOI22_X1 U16478 ( .A1(n14858), .A2(n14872), .B1(n14849), .B2(n14856), .ZN(
        P2_U3460) );
  AND2_X1 U16479 ( .A1(n14850), .A2(n8001), .ZN(n14854) );
  OAI21_X1 U16480 ( .B1(n6821), .B2(n14852), .A(n14851), .ZN(n14853) );
  NOR3_X1 U16481 ( .A1(n14855), .A2(n14854), .A3(n14853), .ZN(n14875) );
  INV_X1 U16482 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14857) );
  AOI22_X1 U16483 ( .A1(n14858), .A2(n14875), .B1(n14857), .B2(n14856), .ZN(
        P2_U3463) );
  AOI22_X1 U16484 ( .A1(n14876), .A2(n14859), .B1(n7729), .B2(n14873), .ZN(
        P2_U3499) );
  AOI22_X1 U16485 ( .A1(n14876), .A2(n14860), .B1(n7739), .B2(n14873), .ZN(
        P2_U3501) );
  AOI22_X1 U16486 ( .A1(n14876), .A2(n14861), .B1(n9882), .B2(n14873), .ZN(
        P2_U3502) );
  AOI22_X1 U16487 ( .A1(n14876), .A2(n14862), .B1(n9884), .B2(n14873), .ZN(
        P2_U3503) );
  AOI22_X1 U16488 ( .A1(n14876), .A2(n14863), .B1(n10000), .B2(n14873), .ZN(
        P2_U3504) );
  AOI22_X1 U16489 ( .A1(n14876), .A2(n14865), .B1(n14864), .B2(n14873), .ZN(
        P2_U3505) );
  AOI22_X1 U16490 ( .A1(n14876), .A2(n14867), .B1(n14866), .B2(n14873), .ZN(
        P2_U3506) );
  AOI22_X1 U16491 ( .A1(n14876), .A2(n14869), .B1(n14868), .B2(n14873), .ZN(
        P2_U3507) );
  AOI22_X1 U16492 ( .A1(n14876), .A2(n14871), .B1(n14870), .B2(n14873), .ZN(
        P2_U3508) );
  AOI22_X1 U16493 ( .A1(n14876), .A2(n14872), .B1(n9999), .B2(n14873), .ZN(
        P2_U3509) );
  AOI22_X1 U16494 ( .A1(n14876), .A2(n14875), .B1(n14874), .B2(n14873), .ZN(
        P2_U3510) );
  NOR2_X1 U16495 ( .A1(P3_U3897), .A2(n14931), .ZN(P3_U3150) );
  INV_X1 U16496 ( .A(n14877), .ZN(n14883) );
  AOI21_X1 U16497 ( .B1(n14880), .B2(n14879), .A(n14878), .ZN(n14882) );
  NOR3_X1 U16498 ( .A1(n14883), .A2(n14882), .A3(n14881), .ZN(n14891) );
  NAND2_X1 U16499 ( .A1(n14885), .A2(n14884), .ZN(n14887) );
  OAI211_X1 U16500 ( .C1(n14889), .C2(n14888), .A(n14887), .B(n14886), .ZN(
        n14890) );
  NOR2_X1 U16501 ( .A1(n14891), .A2(n14890), .ZN(n14892) );
  OAI21_X1 U16502 ( .B1(n14894), .B2(n14893), .A(n14892), .ZN(P3_U3157) );
  AOI21_X1 U16503 ( .B1(n14897), .B2(n14896), .A(n14895), .ZN(n14912) );
  OAI21_X1 U16504 ( .B1(n14917), .B2(n14899), .A(n14898), .ZN(n14910) );
  AOI21_X1 U16505 ( .B1(n14902), .B2(n14901), .A(n14900), .ZN(n14908) );
  AOI21_X1 U16506 ( .B1(n14905), .B2(n14904), .A(n14903), .ZN(n14907) );
  OAI22_X1 U16507 ( .A1(n14908), .A2(n14927), .B1(n14907), .B2(n14906), .ZN(
        n14909) );
  AOI211_X1 U16508 ( .C1(n14931), .C2(P3_ADDR_REG_11__SCAN_IN), .A(n14910), 
        .B(n14909), .ZN(n14911) );
  OAI21_X1 U16509 ( .B1(n14912), .B2(n14933), .A(n14911), .ZN(P3_U3193) );
  AOI21_X1 U16510 ( .B1(n11590), .B2(n14914), .A(n14913), .ZN(n14934) );
  OAI21_X1 U16511 ( .B1(n14917), .B2(n14916), .A(n14915), .ZN(n14930) );
  AOI21_X1 U16512 ( .B1(n14920), .B2(n14919), .A(n14918), .ZN(n14928) );
  OAI21_X1 U16513 ( .B1(n14923), .B2(n14922), .A(n14921), .ZN(n14925) );
  NAND2_X1 U16514 ( .A1(n14925), .A2(n14924), .ZN(n14926) );
  OAI21_X1 U16515 ( .B1(n14928), .B2(n14927), .A(n14926), .ZN(n14929) );
  AOI211_X1 U16516 ( .C1(n14931), .C2(P3_ADDR_REG_13__SCAN_IN), .A(n14930), 
        .B(n14929), .ZN(n14932) );
  OAI21_X1 U16517 ( .B1(n14934), .B2(n14933), .A(n14932), .ZN(P3_U3195) );
  XNOR2_X1 U16518 ( .A(n14935), .B(n14938), .ZN(n14974) );
  INV_X1 U16519 ( .A(n14936), .ZN(n15022) );
  XNOR2_X1 U16520 ( .A(n14937), .B(n14938), .ZN(n14940) );
  NOR2_X1 U16521 ( .A1(n14940), .A2(n14939), .ZN(n14941) );
  AOI211_X1 U16522 ( .C1(n14974), .C2(n15022), .A(n14942), .B(n14941), .ZN(
        n14970) );
  NOR2_X1 U16523 ( .A1(n14943), .A2(n15001), .ZN(n14972) );
  AOI22_X1 U16524 ( .A1(n14972), .A2(n14955), .B1(P3_REG3_REG_2__SCAN_IN), 
        .B2(n14959), .ZN(n14946) );
  INV_X1 U16525 ( .A(n14944), .ZN(n14960) );
  AOI22_X1 U16526 ( .A1(n14974), .A2(n14960), .B1(P3_REG2_REG_2__SCAN_IN), 
        .B2(n14965), .ZN(n14945) );
  OAI221_X1 U16527 ( .B1(n14965), .B2(n14970), .C1(n14965), .C2(n14946), .A(
        n14945), .ZN(P3_U3231) );
  XNOR2_X1 U16528 ( .A(n14947), .B(n10236), .ZN(n14949) );
  NAND2_X1 U16529 ( .A1(n14949), .A2(n14948), .ZN(n14952) );
  INV_X1 U16530 ( .A(n14950), .ZN(n14951) );
  NAND2_X1 U16531 ( .A1(n14952), .A2(n14951), .ZN(n14966) );
  INV_X1 U16532 ( .A(n14966), .ZN(n14958) );
  XNOR2_X1 U16533 ( .A(n14953), .B(n10236), .ZN(n14968) );
  NAND2_X1 U16534 ( .A1(n14968), .A2(n15022), .ZN(n14957) );
  AND2_X1 U16535 ( .A1(n14954), .A2(n15014), .ZN(n14967) );
  NAND2_X1 U16536 ( .A1(n14967), .A2(n14955), .ZN(n14956) );
  AND3_X1 U16537 ( .A1(n14958), .A2(n14957), .A3(n14956), .ZN(n14964) );
  AOI22_X1 U16538 ( .A1(n14968), .A2(n14960), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n14959), .ZN(n14961) );
  OAI221_X1 U16539 ( .B1(n14965), .B2(n14964), .C1(n14963), .C2(n14962), .A(
        n14961), .ZN(P3_U3232) );
  AOI211_X1 U16540 ( .C1(n15007), .C2(n14968), .A(n14967), .B(n14966), .ZN(
        n15027) );
  INV_X1 U16541 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n14969) );
  AOI22_X1 U16542 ( .A1(n15025), .A2(n15027), .B1(n14969), .B2(n15023), .ZN(
        P3_U3393) );
  INV_X1 U16543 ( .A(n15018), .ZN(n14973) );
  INV_X1 U16544 ( .A(n14970), .ZN(n14971) );
  AOI211_X1 U16545 ( .C1(n14974), .C2(n14973), .A(n14972), .B(n14971), .ZN(
        n15028) );
  INV_X1 U16546 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n14975) );
  AOI22_X1 U16547 ( .A1(n15025), .A2(n15028), .B1(n14975), .B2(n15023), .ZN(
        P3_U3396) );
  INV_X1 U16548 ( .A(n14979), .ZN(n14981) );
  NAND2_X1 U16549 ( .A1(n14976), .A2(n15014), .ZN(n14977) );
  OAI211_X1 U16550 ( .C1(n15018), .C2(n14979), .A(n14978), .B(n14977), .ZN(
        n14980) );
  AOI21_X1 U16551 ( .B1(n14981), .B2(n15022), .A(n14980), .ZN(n15029) );
  INV_X1 U16552 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n14982) );
  AOI22_X1 U16553 ( .A1(n15025), .A2(n15029), .B1(n14982), .B2(n15023), .ZN(
        P3_U3399) );
  AOI21_X1 U16554 ( .B1(n14984), .B2(n15014), .A(n14983), .ZN(n14985) );
  OAI21_X1 U16555 ( .B1(n15018), .B2(n14986), .A(n14985), .ZN(n14987) );
  AOI21_X1 U16556 ( .B1(n14988), .B2(n15022), .A(n14987), .ZN(n15031) );
  INV_X1 U16557 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n14989) );
  AOI22_X1 U16558 ( .A1(n15025), .A2(n15031), .B1(n14989), .B2(n15023), .ZN(
        P3_U3402) );
  OAI22_X1 U16559 ( .A1(n14991), .A2(n15018), .B1(n14990), .B2(n15001), .ZN(
        n14992) );
  NOR2_X1 U16560 ( .A1(n14993), .A2(n14992), .ZN(n15032) );
  INV_X1 U16561 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n14994) );
  AOI22_X1 U16562 ( .A1(n15025), .A2(n15032), .B1(n14994), .B2(n15023), .ZN(
        P3_U3405) );
  INV_X1 U16563 ( .A(n14999), .ZN(n14996) );
  OAI22_X1 U16564 ( .A1(n14996), .A2(n15018), .B1(n14995), .B2(n15001), .ZN(
        n14998) );
  AOI211_X1 U16565 ( .C1(n15022), .C2(n14999), .A(n14998), .B(n14997), .ZN(
        n15033) );
  INV_X1 U16566 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15000) );
  AOI22_X1 U16567 ( .A1(n15025), .A2(n15033), .B1(n15000), .B2(n15023), .ZN(
        P3_U3408) );
  OAI22_X1 U16568 ( .A1(n15003), .A2(n15018), .B1(n15002), .B2(n15001), .ZN(
        n15004) );
  NOR2_X1 U16569 ( .A1(n15005), .A2(n15004), .ZN(n15036) );
  INV_X1 U16570 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15006) );
  AOI22_X1 U16571 ( .A1(n15025), .A2(n15036), .B1(n15006), .B2(n15023), .ZN(
        P3_U3411) );
  AND2_X1 U16572 ( .A1(n15008), .A2(n15007), .ZN(n15011) );
  AND2_X1 U16573 ( .A1(n15009), .A2(n15014), .ZN(n15010) );
  NOR3_X1 U16574 ( .A1(n15012), .A2(n15011), .A3(n15010), .ZN(n15038) );
  INV_X1 U16575 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15013) );
  AOI22_X1 U16576 ( .A1(n15025), .A2(n15038), .B1(n15013), .B2(n15023), .ZN(
        P3_U3414) );
  NAND2_X1 U16577 ( .A1(n15015), .A2(n15014), .ZN(n15016) );
  OAI211_X1 U16578 ( .C1(n15019), .C2(n15018), .A(n15017), .B(n15016), .ZN(
        n15020) );
  AOI21_X1 U16579 ( .B1(n15022), .B2(n15021), .A(n15020), .ZN(n15041) );
  INV_X1 U16580 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15024) );
  AOI22_X1 U16581 ( .A1(n15025), .A2(n15041), .B1(n15024), .B2(n15023), .ZN(
        P3_U3417) );
  AOI22_X1 U16582 ( .A1(n15034), .A2(n15027), .B1(n15026), .B2(n15039), .ZN(
        P3_U3460) );
  AOI22_X1 U16583 ( .A1(n15034), .A2(n15028), .B1(n10259), .B2(n15039), .ZN(
        P3_U3461) );
  AOI22_X1 U16584 ( .A1(n15034), .A2(n15029), .B1(n10265), .B2(n15039), .ZN(
        P3_U3462) );
  AOI22_X1 U16585 ( .A1(n15034), .A2(n15031), .B1(n15030), .B2(n15039), .ZN(
        P3_U3463) );
  AOI22_X1 U16586 ( .A1(n15034), .A2(n15032), .B1(n10305), .B2(n15039), .ZN(
        P3_U3464) );
  AOI22_X1 U16587 ( .A1(n15034), .A2(n15033), .B1(n10324), .B2(n15039), .ZN(
        P3_U3465) );
  AOI22_X1 U16588 ( .A1(n15034), .A2(n15036), .B1(n15035), .B2(n15039), .ZN(
        P3_U3466) );
  INV_X1 U16589 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15037) );
  AOI22_X1 U16590 ( .A1(n15034), .A2(n15038), .B1(n15037), .B2(n15039), .ZN(
        P3_U3467) );
  AOI22_X1 U16591 ( .A1(n15034), .A2(n15041), .B1(n15040), .B2(n15039), .ZN(
        P3_U3468) );
  NAND2_X1 U16592 ( .A1(keyinput29), .A2(keyinput3), .ZN(n15048) );
  NOR2_X1 U16593 ( .A1(keyinput49), .A2(keyinput33), .ZN(n15046) );
  NAND3_X1 U16594 ( .A1(keyinput19), .A2(keyinput23), .A3(keyinput55), .ZN(
        n15044) );
  INV_X1 U16595 ( .A(keyinput18), .ZN(n15042) );
  NAND3_X1 U16596 ( .A1(keyinput54), .A2(keyinput24), .A3(n15042), .ZN(n15043)
         );
  NOR4_X1 U16597 ( .A1(keyinput2), .A2(keyinput28), .A3(n15044), .A4(n15043), 
        .ZN(n15045) );
  NAND4_X1 U16598 ( .A1(keyinput59), .A2(keyinput25), .A3(n15046), .A4(n15045), 
        .ZN(n15047) );
  NOR4_X1 U16599 ( .A1(keyinput21), .A2(keyinput26), .A3(n15048), .A4(n15047), 
        .ZN(n15189) );
  NOR3_X1 U16600 ( .A1(keyinput10), .A2(keyinput52), .A3(keyinput63), .ZN(
        n15054) );
  INV_X1 U16601 ( .A(keyinput7), .ZN(n15049) );
  NOR4_X1 U16602 ( .A1(keyinput61), .A2(keyinput60), .A3(keyinput8), .A4(
        n15049), .ZN(n15053) );
  NAND4_X1 U16603 ( .A1(keyinput11), .A2(keyinput41), .A3(keyinput39), .A4(
        keyinput1), .ZN(n15051) );
  NAND2_X1 U16604 ( .A1(keyinput0), .A2(keyinput43), .ZN(n15050) );
  NOR4_X1 U16605 ( .A1(keyinput14), .A2(keyinput20), .A3(n15051), .A4(n15050), 
        .ZN(n15052) );
  NAND4_X1 U16606 ( .A1(keyinput12), .A2(n15054), .A3(n15053), .A4(n15052), 
        .ZN(n15068) );
  NOR4_X1 U16607 ( .A1(keyinput51), .A2(keyinput31), .A3(keyinput45), .A4(
        keyinput57), .ZN(n15060) );
  NOR3_X1 U16608 ( .A1(keyinput34), .A2(keyinput22), .A3(keyinput4), .ZN(
        n15059) );
  NAND2_X1 U16609 ( .A1(keyinput16), .A2(keyinput40), .ZN(n15057) );
  INV_X1 U16610 ( .A(keyinput30), .ZN(n15055) );
  NAND4_X1 U16611 ( .A1(keyinput44), .A2(keyinput36), .A3(keyinput50), .A4(
        n15055), .ZN(n15056) );
  NOR4_X1 U16612 ( .A1(keyinput56), .A2(keyinput6), .A3(n15057), .A4(n15056), 
        .ZN(n15058) );
  NAND4_X1 U16613 ( .A1(n15060), .A2(keyinput32), .A3(n15059), .A4(n15058), 
        .ZN(n15067) );
  NOR4_X1 U16614 ( .A1(keyinput47), .A2(keyinput15), .A3(keyinput58), .A4(
        keyinput53), .ZN(n15062) );
  NOR2_X1 U16615 ( .A1(keyinput5), .A2(keyinput38), .ZN(n15061) );
  NAND4_X1 U16616 ( .A1(n15062), .A2(keyinput48), .A3(keyinput27), .A4(n15061), 
        .ZN(n15066) );
  NOR3_X1 U16617 ( .A1(keyinput37), .A2(keyinput9), .A3(keyinput46), .ZN(
        n15064) );
  NOR3_X1 U16618 ( .A1(keyinput13), .A2(keyinput62), .A3(keyinput42), .ZN(
        n15063) );
  NAND4_X1 U16619 ( .A1(keyinput35), .A2(n15064), .A3(keyinput17), .A4(n15063), 
        .ZN(n15065) );
  NOR4_X1 U16620 ( .A1(n15068), .A2(n15067), .A3(n15066), .A4(n15065), .ZN(
        n15188) );
  AOI22_X1 U16621 ( .A1(n15070), .A2(keyinput39), .B1(keyinput1), .B2(n10818), 
        .ZN(n15069) );
  OAI221_X1 U16622 ( .B1(n15070), .B2(keyinput39), .C1(n10818), .C2(keyinput1), 
        .A(n15069), .ZN(n15080) );
  AOI22_X1 U16623 ( .A1(n8137), .A2(keyinput63), .B1(n15072), .B2(keyinput12), 
        .ZN(n15071) );
  OAI221_X1 U16624 ( .B1(n8137), .B2(keyinput63), .C1(n15072), .C2(keyinput12), 
        .A(n15071), .ZN(n15079) );
  AOI22_X1 U16625 ( .A1(n7967), .A2(keyinput11), .B1(keyinput41), .B2(n15074), 
        .ZN(n15073) );
  OAI221_X1 U16626 ( .B1(n7967), .B2(keyinput11), .C1(n15074), .C2(keyinput41), 
        .A(n15073), .ZN(n15078) );
  XOR2_X1 U16627 ( .A(n8331), .B(keyinput52), .Z(n15076) );
  XNOR2_X1 U16628 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput10), .ZN(n15075)
         );
  NAND2_X1 U16629 ( .A1(n15076), .A2(n15075), .ZN(n15077) );
  NOR4_X1 U16630 ( .A1(n15080), .A2(n15079), .A3(n15078), .A4(n15077), .ZN(
        n15123) );
  AOI22_X1 U16631 ( .A1(n10963), .A2(keyinput60), .B1(n15082), .B2(keyinput8), 
        .ZN(n15081) );
  OAI221_X1 U16632 ( .B1(n10963), .B2(keyinput60), .C1(n15082), .C2(keyinput8), 
        .A(n15081), .ZN(n15093) );
  AOI22_X1 U16633 ( .A1(n15085), .A2(keyinput61), .B1(n15084), .B2(keyinput7), 
        .ZN(n15083) );
  OAI221_X1 U16634 ( .B1(n15085), .B2(keyinput61), .C1(n15084), .C2(keyinput7), 
        .A(n15083), .ZN(n15092) );
  AOI22_X1 U16635 ( .A1(n6876), .A2(keyinput0), .B1(n15087), .B2(keyinput43), 
        .ZN(n15086) );
  OAI221_X1 U16636 ( .B1(n6876), .B2(keyinput0), .C1(n15087), .C2(keyinput43), 
        .A(n15086), .ZN(n15091) );
  XNOR2_X1 U16637 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput20), .ZN(n15088) );
  NAND2_X1 U16638 ( .A1(n15089), .A2(n15088), .ZN(n15090) );
  NOR4_X1 U16639 ( .A1(n15093), .A2(n15092), .A3(n15091), .A4(n15090), .ZN(
        n15122) );
  AOI22_X1 U16640 ( .A1(n15096), .A2(keyinput40), .B1(keyinput6), .B2(n15095), 
        .ZN(n15094) );
  OAI221_X1 U16641 ( .B1(n15096), .B2(keyinput40), .C1(n15095), .C2(keyinput6), 
        .A(n15094), .ZN(n15106) );
  AOI22_X1 U16642 ( .A1(n15099), .A2(keyinput16), .B1(n15098), .B2(keyinput56), 
        .ZN(n15097) );
  OAI221_X1 U16643 ( .B1(n15099), .B2(keyinput16), .C1(n15098), .C2(keyinput56), .A(n15097), .ZN(n15105) );
  XNOR2_X1 U16644 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput31), .ZN(n15103) );
  XNOR2_X1 U16645 ( .A(P1_REG3_REG_8__SCAN_IN), .B(keyinput51), .ZN(n15102) );
  XNOR2_X1 U16646 ( .A(P3_IR_REG_6__SCAN_IN), .B(keyinput45), .ZN(n15101) );
  XNOR2_X1 U16647 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(keyinput57), .ZN(n15100)
         );
  NAND4_X1 U16648 ( .A1(n15103), .A2(n15102), .A3(n15101), .A4(n15100), .ZN(
        n15104) );
  NOR3_X1 U16649 ( .A1(n15106), .A2(n15105), .A3(n15104), .ZN(n15121) );
  AOI22_X1 U16650 ( .A1(n15108), .A2(keyinput34), .B1(n9882), .B2(keyinput22), 
        .ZN(n15107) );
  OAI221_X1 U16651 ( .B1(n15108), .B2(keyinput34), .C1(n9882), .C2(keyinput22), 
        .A(n15107), .ZN(n15119) );
  AOI22_X1 U16652 ( .A1(n12535), .A2(keyinput36), .B1(keyinput44), .B2(n15110), 
        .ZN(n15109) );
  OAI221_X1 U16653 ( .B1(n12535), .B2(keyinput36), .C1(n15110), .C2(keyinput44), .A(n15109), .ZN(n15118) );
  AOI22_X1 U16654 ( .A1(n15113), .A2(keyinput32), .B1(n15112), .B2(keyinput4), 
        .ZN(n15111) );
  OAI221_X1 U16655 ( .B1(n15113), .B2(keyinput32), .C1(n15112), .C2(keyinput4), 
        .A(n15111), .ZN(n15117) );
  XNOR2_X1 U16656 ( .A(P3_REG2_REG_31__SCAN_IN), .B(keyinput50), .ZN(n15115)
         );
  XNOR2_X1 U16657 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput30), .ZN(n15114)
         );
  NAND2_X1 U16658 ( .A1(n15115), .A2(n15114), .ZN(n15116) );
  NOR4_X1 U16659 ( .A1(n15119), .A2(n15118), .A3(n15117), .A4(n15116), .ZN(
        n15120) );
  NAND4_X1 U16660 ( .A1(n15123), .A2(n15122), .A3(n15121), .A4(n15120), .ZN(
        n15187) );
  AOI22_X1 U16661 ( .A1(n12367), .A2(keyinput54), .B1(n9935), .B2(keyinput18), 
        .ZN(n15124) );
  OAI221_X1 U16662 ( .B1(n12367), .B2(keyinput54), .C1(n9935), .C2(keyinput18), 
        .A(n15124), .ZN(n15129) );
  XNOR2_X1 U16663 ( .A(n15125), .B(keyinput49), .ZN(n15128) );
  XNOR2_X1 U16664 ( .A(n15126), .B(keyinput59), .ZN(n15127) );
  OR3_X1 U16665 ( .A1(n15129), .A2(n15128), .A3(n15127), .ZN(n15138) );
  AOI22_X1 U16666 ( .A1(n15132), .A2(keyinput24), .B1(keyinput28), .B2(n15131), 
        .ZN(n15130) );
  OAI221_X1 U16667 ( .B1(n15132), .B2(keyinput24), .C1(n15131), .C2(keyinput28), .A(n15130), .ZN(n15137) );
  AOI22_X1 U16668 ( .A1(n15135), .A2(keyinput25), .B1(n15134), .B2(keyinput33), 
        .ZN(n15133) );
  OAI221_X1 U16669 ( .B1(n15135), .B2(keyinput25), .C1(n15134), .C2(keyinput33), .A(n15133), .ZN(n15136) );
  NOR3_X1 U16670 ( .A1(n15138), .A2(n15137), .A3(n15136), .ZN(n15185) );
  AOI22_X1 U16671 ( .A1(n15141), .A2(keyinput21), .B1(keyinput29), .B2(n15140), 
        .ZN(n15139) );
  OAI221_X1 U16672 ( .B1(n15141), .B2(keyinput21), .C1(n15140), .C2(keyinput29), .A(n15139), .ZN(n15145) );
  XNOR2_X1 U16673 ( .A(n15142), .B(keyinput19), .ZN(n15144) );
  XOR2_X1 U16674 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput23), .Z(n15143) );
  OR3_X1 U16675 ( .A1(n15145), .A2(n15144), .A3(n15143), .ZN(n15152) );
  AOI22_X1 U16676 ( .A1(n15147), .A2(keyinput2), .B1(keyinput55), .B2(n9931), 
        .ZN(n15146) );
  OAI221_X1 U16677 ( .B1(n15147), .B2(keyinput2), .C1(n9931), .C2(keyinput55), 
        .A(n15146), .ZN(n15151) );
  AOI22_X1 U16678 ( .A1(n15149), .A2(keyinput3), .B1(n10988), .B2(keyinput26), 
        .ZN(n15148) );
  OAI221_X1 U16679 ( .B1(n15149), .B2(keyinput3), .C1(n10988), .C2(keyinput26), 
        .A(n15148), .ZN(n15150) );
  NOR3_X1 U16680 ( .A1(n15152), .A2(n15151), .A3(n15150), .ZN(n15184) );
  AOI22_X1 U16681 ( .A1(n15155), .A2(keyinput5), .B1(keyinput38), .B2(n15154), 
        .ZN(n15153) );
  OAI221_X1 U16682 ( .B1(n15155), .B2(keyinput5), .C1(n15154), .C2(keyinput38), 
        .A(n15153), .ZN(n15166) );
  AOI22_X1 U16683 ( .A1(n15157), .A2(keyinput48), .B1(keyinput27), .B2(n7901), 
        .ZN(n15156) );
  OAI221_X1 U16684 ( .B1(n15157), .B2(keyinput48), .C1(n7901), .C2(keyinput27), 
        .A(n15156), .ZN(n15165) );
  AOI22_X1 U16685 ( .A1(n10251), .A2(keyinput62), .B1(keyinput42), .B2(n15159), 
        .ZN(n15158) );
  OAI221_X1 U16686 ( .B1(n10251), .B2(keyinput62), .C1(n15159), .C2(keyinput42), .A(n15158), .ZN(n15164) );
  AOI22_X1 U16687 ( .A1(n15162), .A2(keyinput17), .B1(n15161), .B2(keyinput13), 
        .ZN(n15160) );
  OAI221_X1 U16688 ( .B1(n15162), .B2(keyinput17), .C1(n15161), .C2(keyinput13), .A(n15160), .ZN(n15163) );
  NOR4_X1 U16689 ( .A1(n15166), .A2(n15165), .A3(n15164), .A4(n15163), .ZN(
        n15183) );
  AOI22_X1 U16690 ( .A1(n15169), .A2(keyinput35), .B1(keyinput46), .B2(n15168), 
        .ZN(n15167) );
  OAI221_X1 U16691 ( .B1(n15169), .B2(keyinput35), .C1(n15168), .C2(keyinput46), .A(n15167), .ZN(n15181) );
  AOI22_X1 U16692 ( .A1(n15172), .A2(keyinput37), .B1(keyinput9), .B2(n15171), 
        .ZN(n15170) );
  OAI221_X1 U16693 ( .B1(n15172), .B2(keyinput37), .C1(n15171), .C2(keyinput9), 
        .A(n15170), .ZN(n15180) );
  INV_X1 U16694 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n15175) );
  AOI22_X1 U16695 ( .A1(n15175), .A2(keyinput58), .B1(keyinput53), .B2(n15174), 
        .ZN(n15173) );
  OAI221_X1 U16696 ( .B1(n15175), .B2(keyinput58), .C1(n15174), .C2(keyinput53), .A(n15173), .ZN(n15179) );
  INV_X1 U16697 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n15177) );
  AOI22_X1 U16698 ( .A1(n8059), .A2(keyinput47), .B1(n15177), .B2(keyinput15), 
        .ZN(n15176) );
  OAI221_X1 U16699 ( .B1(n8059), .B2(keyinput47), .C1(n15177), .C2(keyinput15), 
        .A(n15176), .ZN(n15178) );
  NOR4_X1 U16700 ( .A1(n15181), .A2(n15180), .A3(n15179), .A4(n15178), .ZN(
        n15182) );
  NAND4_X1 U16701 ( .A1(n15185), .A2(n15184), .A3(n15183), .A4(n15182), .ZN(
        n15186) );
  AOI211_X1 U16702 ( .C1(n15189), .C2(n15188), .A(n15187), .B(n15186), .ZN(
        n15193) );
  MUX2_X1 U16703 ( .A(n15191), .B(n15190), .S(P1_U4016), .Z(n15192) );
  XNOR2_X1 U16704 ( .A(n15193), .B(n15192), .ZN(P1_U3582) );
  XNOR2_X1 U16705 ( .A(n15195), .B(n15194), .ZN(SUB_1596_U59) );
  XOR2_X1 U16706 ( .A(n15197), .B(n15196), .Z(SUB_1596_U58) );
  AOI21_X1 U16707 ( .B1(n15199), .B2(n15198), .A(n15208), .ZN(SUB_1596_U53) );
  XOR2_X1 U16708 ( .A(n15201), .B(n15200), .Z(SUB_1596_U56) );
  OAI21_X1 U16709 ( .B1(n15204), .B2(n15203), .A(n15202), .ZN(n15206) );
  XOR2_X1 U16710 ( .A(n15206), .B(n15205), .Z(SUB_1596_U60) );
  XOR2_X1 U16711 ( .A(n15208), .B(n15207), .Z(SUB_1596_U5) );
  AND2_X1 U7266 ( .A1(n10511), .A2(n10510), .ZN(n10630) );
  CLKBUF_X1 U7205 ( .A(n10279), .Z(n6447) );
  CLKBUF_X1 U7210 ( .A(n7538), .Z(n9862) );
  CLKBUF_X1 U7279 ( .A(n6444), .Z(n12090) );
  INV_X1 U7308 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8973) );
endmodule

