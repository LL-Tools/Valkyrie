

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n5031, n5032, n5033, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028;

  NAND2_X1 U5096 ( .A1(n9287), .A2(n8212), .ZN(n9261) );
  NAND2_X2 U5097 ( .A1(n5135), .A2(n7782), .ZN(n10970) );
  XNOR2_X1 U5098 ( .A(n9850), .B(n10857), .ZN(n9764) );
  BUF_X2 U5099 ( .A(n7104), .Z(n5039) );
  CLKBUF_X2 U5100 ( .A(n5854), .Z(n8430) );
  OR2_X1 U5102 ( .A1(n8581), .A2(n9316), .ZN(n8579) );
  INV_X2 U5103 ( .A(n8535), .ZN(n8562) );
  INV_X1 U5104 ( .A(n8374), .ZN(n8266) );
  NAND2_X2 U5105 ( .A1(n6521), .A2(n6519), .ZN(n8321) );
  INV_X1 U5106 ( .A(n9940), .ZN(n9973) );
  AND3_X1 U5107 ( .A1(n5846), .A2(n5847), .A3(n5845), .ZN(n10870) );
  INV_X1 U5108 ( .A(n8266), .ZN(n8324) );
  NAND4_X1 U5109 ( .A1(n5787), .A2(n5785), .A3(n5786), .A4(n5788), .ZN(n7241)
         );
  NAND4_X2 U5110 ( .A1(n6526), .A2(n6525), .A3(n6524), .A4(n6523), .ZN(n8998)
         );
  INV_X2 U5111 ( .A(n10829), .ZN(n9303) );
  INV_X1 U5112 ( .A(n6519), .ZN(n9423) );
  INV_X1 U5113 ( .A(n10806), .ZN(n6793) );
  NAND4_X2 U5114 ( .A1(n5772), .A2(n5771), .A3(n5770), .A4(n5769), .ZN(n6891)
         );
  INV_X1 U5115 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10261) );
  AND4_X1 U5116 ( .A1(n6449), .A2(n6451), .A3(n6450), .A4(n6453), .ZN(n5031)
         );
  NAND2_X2 U5117 ( .A1(n7461), .A2(n7460), .ZN(n7522) );
  NAND2_X2 U5118 ( .A1(n10108), .A2(n10107), .ZN(n10106) );
  NOR2_X2 U5119 ( .A1(n6113), .A2(n6110), .ZN(n6108) );
  INV_X2 U5120 ( .A(n7288), .ZN(n5913) );
  OAI21_X2 U5121 ( .B1(n6116), .B2(n6115), .A(n6114), .ZN(n6142) );
  OAI21_X2 U5122 ( .B1(n9014), .B2(P2_REG2_REG_14__SCAN_IN), .A(n9013), .ZN(
        n9026) );
  INV_X1 U5123 ( .A(n7400), .ZN(n10851) );
  NOR2_X2 U5124 ( .A1(n5740), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5744) );
  AOI21_X2 U5125 ( .B1(n9573), .B2(n8616), .A(n8615), .ZN(n9098) );
  NAND2_X1 U5126 ( .A1(n6435), .A2(n8463), .ZN(n5032) );
  NAND2_X1 U5127 ( .A1(n6435), .A2(n8463), .ZN(n5033) );
  AOI211_X2 U5128 ( .C1(n10115), .C2(n10169), .A(n9956), .B(n9955), .ZN(n9957)
         );
  NAND2_X1 U5129 ( .A1(n6520), .A2(n6519), .ZN(n8374) );
  NAND2_X2 U5132 ( .A1(n5413), .A2(n5412), .ZN(n9945) );
  NOR2_X2 U5133 ( .A1(n7718), .A2(n7717), .ZN(n7839) );
  XNOR2_X2 U5134 ( .A(n6064), .B(n5649), .ZN(n7991) );
  AOI22_X2 U5135 ( .A1(n10806), .A2(n6522), .B1(P2_REG2_REG_2__SCAN_IN), .B2(
        n6793), .ZN(n10804) );
  AOI21_X2 U5136 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n10806), .A(n10802), .ZN(
        n6829) );
  XNOR2_X2 U5137 ( .A(n6536), .B(P2_IR_REG_2__SCAN_IN), .ZN(n10806) );
  XNOR2_X2 U5138 ( .A(n6543), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6791) );
  OR2_X1 U5139 ( .A1(n8955), .A2(n8954), .ZN(n8956) );
  NOR2_X1 U5140 ( .A1(n7942), .A2(n7944), .ZN(n7946) );
  AND2_X1 U5141 ( .A1(n6010), .A2(n6009), .ZN(n7941) );
  NAND2_X2 U5142 ( .A1(n9698), .A2(n9694), .ZN(n9780) );
  AND2_X1 U5143 ( .A1(n7628), .A2(n7704), .ZN(n7629) );
  OR2_X1 U5144 ( .A1(n7679), .A2(n7564), .ZN(n9660) );
  OR2_X1 U5145 ( .A1(n5966), .A2(n5965), .ZN(n5692) );
  INV_X4 U5146 ( .A(n6208), .ZN(n8422) );
  INV_X2 U5147 ( .A(n8551), .ZN(n8563) );
  INV_X2 U5148 ( .A(n7315), .ZN(n10877) );
  NAND2_X1 U5149 ( .A1(n5795), .A2(n5794), .ZN(n10839) );
  INV_X1 U5150 ( .A(n7296), .ZN(n9594) );
  INV_X2 U5151 ( .A(n8233), .ZN(n8811) );
  CLKBUF_X2 U5152 ( .A(n5806), .Z(n8432) );
  INV_X2 U5153 ( .A(n6473), .ZN(n5814) );
  CLKBUF_X2 U5154 ( .A(n7104), .Z(n5038) );
  NAND2_X1 U5155 ( .A1(n7537), .A2(n6535), .ZN(n6544) );
  OR2_X1 U5156 ( .A1(n5762), .A2(n9798), .ZN(n7248) );
  NAND2_X1 U5157 ( .A1(n7537), .A2(n5668), .ZN(n7104) );
  NAND2_X1 U5158 ( .A1(n6535), .A2(P1_U3084), .ZN(n10267) );
  CLKBUF_X2 U5159 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n10753) );
  OR2_X1 U5160 ( .A1(n8813), .A2(n8812), .ZN(n8815) );
  AND2_X1 U5161 ( .A1(n10154), .A2(n10153), .ZN(n10155) );
  NAND2_X1 U5162 ( .A1(n5197), .A2(n5196), .ZN(n8814) );
  AND2_X1 U5163 ( .A1(n8560), .A2(n8559), .ZN(n8830) );
  AOI211_X1 U5164 ( .C1(n10115), .C2(n10164), .A(n9942), .B(n9941), .ZN(n9943)
         );
  OR2_X1 U5165 ( .A1(n6385), .A2(n6384), .ZN(n8445) );
  AND2_X1 U5166 ( .A1(n5449), .A2(n5199), .ZN(n5198) );
  AOI211_X1 U5167 ( .C1(n10131), .C2(n9940), .A(n9939), .B(n9938), .ZN(n10166)
         );
  OAI21_X1 U5168 ( .B1(n9969), .B2(n5141), .A(n10125), .ZN(n5140) );
  NOR2_X1 U5169 ( .A1(n9969), .A2(n8451), .ZN(n9952) );
  AND2_X1 U5170 ( .A1(n5622), .A2(n9738), .ZN(n9969) );
  NOR2_X1 U5171 ( .A1(n8557), .A2(n5444), .ZN(n5443) );
  NOR2_X1 U5172 ( .A1(n8581), .A2(n5331), .ZN(n9097) );
  XNOR2_X1 U5173 ( .A(n8612), .B(n8611), .ZN(n10260) );
  AND2_X1 U5174 ( .A1(n8609), .A2(n8507), .ZN(n9573) );
  OR2_X1 U5175 ( .A1(n8506), .A2(n8505), .ZN(n8507) );
  NAND2_X1 U5176 ( .A1(n8343), .A2(SI_29_), .ZN(n8501) );
  XNOR2_X1 U5177 ( .A(n8497), .B(n8498), .ZN(n8343) );
  OAI21_X1 U5178 ( .B1(n6368), .B2(n5514), .A(n5512), .ZN(n8497) );
  NAND2_X1 U5179 ( .A1(n8263), .A2(n8262), .ZN(n9347) );
  NAND2_X1 U5180 ( .A1(n8278), .A2(n8277), .ZN(n9162) );
  OAI21_X1 U5181 ( .B1(n6347), .B2(n6346), .A(n6345), .ZN(n6366) );
  NAND2_X1 U5182 ( .A1(n8074), .A2(n8073), .ZN(n8392) );
  OAI21_X1 U5183 ( .B1(n6325), .B2(n6324), .A(n6323), .ZN(n6347) );
  NAND2_X1 U5184 ( .A1(n5421), .A2(n5419), .ZN(n8074) );
  NAND2_X1 U5185 ( .A1(n6303), .A2(n6302), .ZN(n6325) );
  AOI21_X1 U5186 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n9054), .A(n9053), .ZN(
        n9056) );
  INV_X1 U5187 ( .A(n5603), .ZN(n5602) );
  AND2_X1 U5188 ( .A1(n8095), .A2(n8094), .ZN(n8115) );
  AOI21_X1 U5189 ( .B1(n7941), .B2(n5604), .A(n5085), .ZN(n5603) );
  AOI21_X1 U5190 ( .B1(n5620), .B2(n5050), .A(n5617), .ZN(n5616) );
  NAND2_X1 U5191 ( .A1(n6235), .A2(n6234), .ZN(n6237) );
  NAND2_X1 U5192 ( .A1(n7864), .A2(n9775), .ZN(n7961) );
  OR2_X1 U5193 ( .A1(n8020), .A2(n7957), .ZN(n9678) );
  NAND2_X1 U5194 ( .A1(n6053), .A2(n6052), .ZN(n8146) );
  NAND2_X1 U5195 ( .A1(n6025), .A2(n6024), .ZN(n10233) );
  NAND2_X1 U5196 ( .A1(n7751), .A2(n7750), .ZN(n7856) );
  AND2_X1 U5197 ( .A1(n9669), .A2(n9670), .ZN(n9772) );
  XNOR2_X1 U5198 ( .A(n6015), .B(n5066), .ZN(n7781) );
  NAND2_X1 U5199 ( .A1(n5485), .A2(n5486), .ZN(n6015) );
  OR2_X1 U5200 ( .A1(n5692), .A2(n5489), .ZN(n5485) );
  AND3_X1 U5201 ( .A1(n7452), .A2(n7451), .A3(n7450), .ZN(n10931) );
  NAND2_X1 U5202 ( .A1(n5682), .A2(n5681), .ZN(n5946) );
  INV_X2 U5203 ( .A(n10093), .ZN(n10141) );
  AND3_X1 U5204 ( .A1(n7109), .A2(n7108), .A3(n7107), .ZN(n10898) );
  AND2_X1 U5205 ( .A1(n8633), .A2(n8634), .ZN(n8629) );
  OAI211_X1 U5206 ( .C1(n7103), .C2(n8453), .A(n5894), .B(n5893), .ZN(n7500)
         );
  NAND2_X1 U5207 ( .A1(n5675), .A2(n5674), .ZN(n5905) );
  AND2_X2 U5208 ( .A1(n6648), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  CLKBUF_X1 U5209 ( .A(n7199), .Z(n10820) );
  OR2_X2 U5210 ( .A1(n5779), .A2(n7248), .ZN(n6208) );
  NAND4_X1 U5211 ( .A1(n5889), .A2(n5888), .A3(n5887), .A4(n5886), .ZN(n9849)
         );
  NAND2_X1 U5212 ( .A1(n5671), .A2(n5670), .ZN(n5891) );
  CLKBUF_X1 U5214 ( .A(n5755), .Z(n6471) );
  AND4_X1 U5215 ( .A1(n6552), .A2(n6551), .A3(n6550), .A4(n6549), .ZN(n7221)
         );
  NAND2_X2 U5216 ( .A1(n7255), .A2(n7248), .ZN(n7288) );
  OR2_X1 U5217 ( .A1(n8374), .A2(n6790), .ZN(n6524) );
  NAND2_X1 U5218 ( .A1(n5667), .A2(n5666), .ZN(n5863) );
  AND2_X1 U5219 ( .A1(n6520), .A2(n9423), .ZN(n7118) );
  AND2_X2 U5220 ( .A1(n6513), .A2(n6512), .ZN(n8233) );
  NAND2_X1 U5221 ( .A1(n5142), .A2(n5662), .ZN(n5840) );
  NAND2_X1 U5222 ( .A1(n5729), .A2(n5728), .ZN(n8130) );
  INV_X1 U5223 ( .A(n10269), .ZN(n5748) );
  CLKBUF_X2 U5224 ( .A(n6544), .Z(n5037) );
  NAND2_X1 U5225 ( .A1(n5745), .A2(n10262), .ZN(n10269) );
  MUX2_X1 U5226 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5743), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5745) );
  OR2_X1 U5227 ( .A1(n5744), .A2(n10261), .ZN(n5741) );
  NAND2_X1 U5228 ( .A1(n5595), .A2(n5594), .ZN(n8463) );
  XNOR2_X1 U5229 ( .A(n6534), .B(n6533), .ZN(n8375) );
  NOR2_X1 U5230 ( .A1(n10783), .A2(n5068), .ZN(n10803) );
  INV_X2 U5231 ( .A(n9420), .ZN(n8494) );
  INV_X2 U5232 ( .A(n10660), .ZN(n10265) );
  INV_X2 U5233 ( .A(n6701), .ZN(n5036) );
  INV_X1 U5234 ( .A(n6093), .ZN(n5736) );
  OAI21_X1 U5235 ( .B1(n5176), .B2(n10261), .A(n10420), .ZN(n5175) );
  AND2_X1 U5236 ( .A1(n5640), .A2(n10633), .ZN(n5639) );
  AND2_X1 U5237 ( .A1(n5647), .A2(n5704), .ZN(n5176) );
  AND2_X1 U5238 ( .A1(n5527), .A2(n5526), .ZN(n6666) );
  AND3_X1 U5239 ( .A1(n10619), .A2(n5704), .A3(n6070), .ZN(n5056) );
  INV_X1 U5240 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n10630) );
  INV_X4 U5241 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U5242 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5527) );
  NOR2_X1 U5243 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5526) );
  INV_X2 U5244 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n10618) );
  INV_X4 U5245 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U5246 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10619) );
  NOR2_X1 U5247 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n6453) );
  INV_X1 U5248 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6070) );
  INV_X1 U5249 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6021) );
  INV_X1 U5250 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n10593) );
  INV_X1 U5251 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n10592) );
  INV_X1 U5252 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U5253 ( .A1(n8470), .A2(n8469), .ZN(n10124) );
  NOR2_X2 U5254 ( .A1(n9199), .A2(n9347), .ZN(n9180) );
  INV_X2 U5255 ( .A(n5656), .ZN(n5663) );
  OR2_X1 U5256 ( .A1(n5039), .A2(n5137), .ZN(n6566) );
  NOR2_X2 U5257 ( .A1(n9936), .A2(n9937), .ZN(n9935) );
  OAI21_X2 U5258 ( .B1(n9971), .B2(n5626), .A(n5623), .ZN(n9936) );
  NAND4_X4 U5259 ( .A1(n5835), .A2(n5837), .A3(n5836), .A4(n5834), .ZN(n7246)
         );
  NAND2_X1 U5260 ( .A1(n5804), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5772) );
  XNOR2_X2 U5261 ( .A(n7241), .B(n10839), .ZN(n7284) );
  NAND2_X2 U5262 ( .A1(n5951), .A2(n5950), .ZN(n7679) );
  AOI21_X2 U5263 ( .B1(n10124), .B2(n10123), .A(n8471), .ZN(n10105) );
  AND2_X2 U5264 ( .A1(n9673), .A2(n9674), .ZN(n9773) );
  AOI21_X2 U5265 ( .B1(n9061), .B2(P2_REG2_REG_17__SCAN_IN), .A(n9060), .ZN(
        n9082) );
  NAND2_X1 U5266 ( .A1(n5747), .A2(n10269), .ZN(n5854) );
  XNOR2_X1 U5267 ( .A(n5658), .B(n10511), .ZN(n5791) );
  NAND2_X1 U5268 ( .A1(n5657), .A2(n6547), .ZN(n5658) );
  INV_X2 U5269 ( .A(n5842), .ZN(n9574) );
  OAI21_X2 U5270 ( .B1(n9931), .B2(n9788), .A(n5393), .ZN(n9918) );
  BUF_X4 U5271 ( .A(n5804), .Z(n5040) );
  INV_X1 U5272 ( .A(SI_21_), .ZN(n10484) );
  INV_X1 U5273 ( .A(n6042), .ZN(n5202) );
  OR2_X1 U5274 ( .A1(n9316), .A2(n8833), .ZN(n8749) );
  AND2_X1 U5275 ( .A1(n9133), .A2(n8871), .ZN(n8737) );
  NOR2_X1 U5276 ( .A1(n6170), .A2(n5568), .ZN(n5567) );
  INV_X1 U5277 ( .A(n9494), .ZN(n5568) );
  NAND2_X1 U5278 ( .A1(n6216), .A2(n6215), .ZN(n6235) );
  NAND2_X1 U5279 ( .A1(n6144), .A2(n6143), .ZN(n6174) );
  INV_X1 U5280 ( .A(n8253), .ZN(n8370) );
  NAND2_X1 U5281 ( .A1(n6511), .A2(n6510), .ZN(n6512) );
  OR2_X1 U5282 ( .A1(n9311), .A2(n9316), .ZN(n5331) );
  INV_X2 U5283 ( .A(n5855), .ZN(n6429) );
  INV_X1 U5284 ( .A(n5634), .ZN(n5633) );
  AND2_X1 U5285 ( .A1(n9620), .A2(n5631), .ZN(n5630) );
  NAND2_X1 U5286 ( .A1(n7863), .A2(n7862), .ZN(n7864) );
  NAND2_X1 U5287 ( .A1(n10479), .A2(keyinput_132), .ZN(n5336) );
  AOI21_X1 U5288 ( .B1(n8842), .B2(n8841), .A(n8539), .ZN(n8543) );
  INV_X1 U5289 ( .A(n6520), .ZN(n6521) );
  OR3_X1 U5290 ( .A1(n8281), .A2(n8280), .A3(n8279), .ZN(n8294) );
  NAND2_X1 U5291 ( .A1(n5456), .A2(n8692), .ZN(n5454) );
  OR2_X1 U5292 ( .A1(n9389), .A2(n8390), .ZN(n8689) );
  OAI22_X1 U5293 ( .A1(n7178), .A2(n7398), .B1(n7185), .B2(n10851), .ZN(n7207)
         );
  AND2_X1 U5294 ( .A1(n7185), .A2(n10851), .ZN(n7178) );
  NAND2_X1 U5295 ( .A1(n9262), .A2(n8764), .ZN(n8364) );
  AOI21_X1 U5296 ( .B1(n9249), .B2(n5468), .A(n5467), .ZN(n5466) );
  INV_X1 U5297 ( .A(n8706), .ZN(n5467) );
  INV_X1 U5298 ( .A(n8363), .ZN(n5468) );
  NAND2_X1 U5299 ( .A1(n9493), .A2(n6169), .ZN(n5566) );
  OR2_X1 U5300 ( .A1(n10179), .A2(n9974), .ZN(n9656) );
  NAND2_X1 U5301 ( .A1(n10179), .A2(n9974), .ZN(n9655) );
  OR2_X1 U5302 ( .A1(n10223), .A2(n9558), .ZN(n9705) );
  OR2_X1 U5303 ( .A1(n9567), .A2(n9429), .ZN(n9699) );
  INV_X1 U5304 ( .A(n9674), .ZN(n5635) );
  AND2_X1 U5305 ( .A1(n10077), .A2(n8472), .ZN(n5411) );
  NAND2_X1 U5306 ( .A1(n5765), .A2(n10659), .ZN(n9731) );
  NAND2_X1 U5307 ( .A1(n6395), .A2(n5734), .ZN(n5755) );
  NOR2_X1 U5308 ( .A1(n8130), .A2(n7976), .ZN(n5734) );
  INV_X1 U5309 ( .A(n6264), .ZN(n5505) );
  AND2_X1 U5310 ( .A1(n6236), .A2(n6219), .ZN(n6234) );
  AOI21_X1 U5311 ( .B1(n5494), .B2(n5496), .A(n5093), .ZN(n5493) );
  INV_X1 U5312 ( .A(n5643), .ZN(n5433) );
  NOR2_X1 U5313 ( .A1(n7033), .A2(n7032), .ZN(n7031) );
  OR2_X1 U5314 ( .A1(n7374), .A2(n7373), .ZN(n7376) );
  NAND2_X1 U5315 ( .A1(n5216), .A2(n8763), .ZN(n8798) );
  XNOR2_X1 U5316 ( .A(n5509), .B(n8811), .ZN(n5508) );
  NOR2_X1 U5317 ( .A1(n8795), .A2(n8794), .ZN(n5510) );
  AOI21_X1 U5318 ( .B1(n8582), .B2(n8353), .A(n8337), .ZN(n8833) );
  NAND2_X1 U5319 ( .A1(n5436), .A2(n5435), .ZN(n5434) );
  INV_X1 U5320 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U5321 ( .A1(n5534), .A2(n5546), .ZN(n5533) );
  INV_X1 U5322 ( .A(n5539), .ZN(n5534) );
  AOI21_X1 U5323 ( .B1(n5542), .B2(n5541), .A(n5540), .ZN(n5539) );
  INV_X1 U5324 ( .A(n5544), .ZN(n5541) );
  INV_X1 U5325 ( .A(n5546), .ZN(n5537) );
  NOR2_X1 U5326 ( .A1(n9119), .A2(n9136), .ZN(n5544) );
  OR2_X1 U5327 ( .A1(n9162), .A2(n9168), .ZN(n8289) );
  OR2_X1 U5328 ( .A1(n9221), .A2(n9233), .ZN(n5645) );
  NAND2_X1 U5329 ( .A1(n8688), .A2(n8689), .ZN(n8161) );
  NAND2_X1 U5330 ( .A1(n8007), .A2(n5558), .ZN(n8064) );
  AND2_X1 U5331 ( .A1(n8781), .A2(n8006), .ZN(n5558) );
  INV_X1 U5332 ( .A(n5038), .ZN(n8235) );
  INV_X1 U5333 ( .A(n7537), .ZN(n8234) );
  INV_X1 U5334 ( .A(n9272), .ZN(n9254) );
  NAND2_X1 U5335 ( .A1(n7184), .A2(n8812), .ZN(n10822) );
  NAND2_X1 U5336 ( .A1(n8331), .A2(n8330), .ZN(n9316) );
  AND2_X1 U5337 ( .A1(n6480), .A2(n6479), .ZN(n7231) );
  AND2_X2 U5338 ( .A1(n5235), .A2(n6518), .ZN(n6519) );
  NOR2_X1 U5339 ( .A1(n6669), .A2(n5525), .ZN(n5524) );
  INV_X1 U5340 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6448) );
  INV_X1 U5341 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6508) );
  AND2_X1 U5342 ( .A1(n5160), .A2(n5167), .ZN(n5158) );
  INV_X1 U5343 ( .A(n9465), .ZN(n5167) );
  INV_X1 U5344 ( .A(n8432), .ZN(n8458) );
  INV_X1 U5345 ( .A(n5040), .ZN(n8462) );
  NAND2_X1 U5346 ( .A1(n5047), .A2(n5079), .ZN(n5594) );
  NOR2_X1 U5347 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5596) );
  OR2_X1 U5348 ( .A1(n10184), .A2(n10015), .ZN(n8478) );
  OR2_X1 U5349 ( .A1(n10198), .A2(n10068), .ZN(n8475) );
  INV_X1 U5350 ( .A(n5613), .ZN(n5612) );
  OAI21_X1 U5351 ( .B1(n5045), .B2(n5614), .A(n10067), .ZN(n5613) );
  INV_X1 U5352 ( .A(n9713), .ZN(n5614) );
  AND4_X1 U5353 ( .A1(n6061), .A2(n6060), .A3(n6059), .A4(n6058), .ZN(n8106)
         );
  BUF_X1 U5354 ( .A(n5838), .Z(n6176) );
  NAND2_X1 U5355 ( .A1(n7816), .A2(n7815), .ZN(n5410) );
  NAND2_X1 U5356 ( .A1(n5628), .A2(n5081), .ZN(n7808) );
  BUF_X1 U5357 ( .A(n5842), .Z(n6199) );
  AOI21_X1 U5358 ( .B1(n5765), .B2(n7248), .A(n10659), .ZN(n5763) );
  NAND2_X1 U5359 ( .A1(n5033), .A2(n6535), .ZN(n5842) );
  INV_X1 U5360 ( .A(n8453), .ZN(n5838) );
  CLKBUF_X1 U5361 ( .A(n5722), .Z(n5723) );
  NAND2_X1 U5362 ( .A1(n5479), .A2(n5073), .ZN(n6216) );
  INV_X1 U5363 ( .A(n6196), .ZN(n5478) );
  OAI21_X1 U5364 ( .B1(n6174), .B2(n6173), .A(n6172), .ZN(n6190) );
  AND2_X1 U5365 ( .A1(n5422), .A2(n5420), .ZN(n5419) );
  NAND2_X1 U5366 ( .A1(n5044), .A2(n7838), .ZN(n5420) );
  INV_X1 U5367 ( .A(n9998), .ZN(n10184) );
  NAND2_X1 U5368 ( .A1(n9536), .A2(n5563), .ZN(n9449) );
  INV_X1 U5369 ( .A(n9537), .ZN(n5569) );
  NAND2_X1 U5370 ( .A1(keyinput_131), .A2(SI_29_), .ZN(n5335) );
  NAND2_X1 U5371 ( .A1(n5334), .A2(SI_28_), .ZN(n5333) );
  XNOR2_X1 U5372 ( .A(n5338), .B(SI_30_), .ZN(n5337) );
  INV_X1 U5373 ( .A(keyinput_4), .ZN(n5270) );
  INV_X1 U5374 ( .A(keyinput_3), .ZN(n5268) );
  XNOR2_X1 U5375 ( .A(n5272), .B(keyinput_2), .ZN(n5271) );
  NAND2_X1 U5376 ( .A1(n5341), .A2(n5339), .ZN(n10487) );
  INV_X1 U5377 ( .A(n5340), .ZN(n5339) );
  AOI21_X1 U5378 ( .B1(n5289), .B2(n5286), .A(n5283), .ZN(n10331) );
  AND2_X1 U5379 ( .A1(n5288), .A2(n5287), .ZN(n5286) );
  NAND2_X1 U5380 ( .A1(n5285), .A2(n5284), .ZN(n5283) );
  OAI21_X1 U5381 ( .B1(n10321), .B2(n5127), .A(n5290), .ZN(n5289) );
  NAND2_X1 U5382 ( .A1(n5255), .A2(n5254), .ZN(n5253) );
  AOI22_X1 U5383 ( .A1(n10336), .A2(n10498), .B1(keyinput_22), .B2(SI_10_), 
        .ZN(n5254) );
  NAND2_X1 U5384 ( .A1(n5258), .A2(n5256), .ZN(n5255) );
  NAND2_X1 U5385 ( .A1(n5227), .A2(n5472), .ZN(n5226) );
  AOI21_X1 U5386 ( .B1(n5250), .B2(n10342), .A(n5128), .ZN(n10343) );
  NAND2_X1 U5387 ( .A1(n5369), .A2(n5368), .ZN(n5367) );
  AOI22_X1 U5388 ( .A1(n10520), .A2(n10519), .B1(keyinput_164), .B2(
        P2_REG3_REG_27__SCAN_IN), .ZN(n5368) );
  NAND2_X1 U5389 ( .A1(n5371), .A2(n5370), .ZN(n5369) );
  NAND2_X1 U5390 ( .A1(n5363), .A2(n5119), .ZN(n5362) );
  NOR2_X1 U5391 ( .A1(n10528), .A2(n10529), .ZN(n5363) );
  AND2_X1 U5392 ( .A1(n5366), .A2(n5365), .ZN(n5364) );
  NAND2_X1 U5393 ( .A1(n10522), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U5394 ( .A1(n10521), .A2(keyinput_165), .ZN(n5365) );
  NAND2_X1 U5395 ( .A1(n8677), .A2(n8760), .ZN(n5222) );
  NAND2_X1 U5396 ( .A1(n8673), .A2(n5223), .ZN(n8671) );
  AND2_X1 U5397 ( .A1(n8668), .A2(n8667), .ZN(n5223) );
  NAND2_X1 U5398 ( .A1(n5280), .A2(n5279), .ZN(n5278) );
  AOI22_X1 U5399 ( .A1(n10520), .A2(n10350), .B1(keyinput_36), .B2(
        P2_REG3_REG_27__SCAN_IN), .ZN(n5279) );
  NAND2_X1 U5400 ( .A1(n5282), .A2(n5281), .ZN(n5280) );
  NAND2_X1 U5401 ( .A1(n5274), .A2(n5120), .ZN(n5273) );
  NOR2_X1 U5402 ( .A1(n10354), .A2(n10355), .ZN(n5274) );
  AND2_X1 U5403 ( .A1(n5277), .A2(n5276), .ZN(n5275) );
  NAND2_X1 U5404 ( .A1(n10351), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U5405 ( .A1(n10521), .A2(keyinput_37), .ZN(n5276) );
  AND2_X1 U5406 ( .A1(n8784), .A2(n8687), .ZN(n5218) );
  OAI21_X1 U5407 ( .B1(n10553), .B2(n10552), .A(n5349), .ZN(n5348) );
  AND2_X1 U5408 ( .A1(n10551), .A2(n5350), .ZN(n5349) );
  NAND2_X1 U5409 ( .A1(n5247), .A2(n5246), .ZN(n5245) );
  INV_X1 U5410 ( .A(n10380), .ZN(n5246) );
  OAI21_X1 U5411 ( .B1(n10371), .B2(n10372), .A(n5248), .ZN(n5247) );
  OAI21_X1 U5412 ( .B1(n10579), .B2(n10580), .A(n5375), .ZN(n5374) );
  XNOR2_X1 U5413 ( .A(n5992), .B(n5376), .ZN(n5375) );
  NOR4_X1 U5414 ( .A1(n10578), .A2(n10577), .A3(n10576), .A4(n10575), .ZN(
        n10579) );
  NOR2_X1 U5415 ( .A1(n10590), .A2(n10591), .ZN(n5373) );
  AOI21_X1 U5416 ( .B1(n10387), .B2(n10388), .A(n5261), .ZN(n5260) );
  XNOR2_X1 U5417 ( .A(keyinput_86), .B(P2_DATAO_REG_10__SCAN_IN), .ZN(n5261)
         );
  NAND2_X1 U5418 ( .A1(n10389), .A2(n10390), .ZN(n5259) );
  NAND2_X1 U5419 ( .A1(n8743), .A2(n5540), .ZN(n5214) );
  MUX2_X1 U5420 ( .A(n8741), .B(n8740), .S(n8752), .Z(n8743) );
  AND2_X1 U5421 ( .A1(n5706), .A2(n5609), .ZN(n5608) );
  INV_X1 U5422 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5609) );
  INV_X1 U5423 ( .A(SI_23_), .ZN(n10473) );
  AND2_X1 U5424 ( .A1(n5427), .A2(n7841), .ZN(n5426) );
  NAND2_X1 U5425 ( .A1(n5427), .A2(n8023), .ZN(n5425) );
  NAND2_X1 U5426 ( .A1(n5095), .A2(n5450), .ZN(n5449) );
  NAND2_X1 U5427 ( .A1(n8809), .A2(n5452), .ZN(n5450) );
  NAND2_X1 U5428 ( .A1(n8806), .A2(n5200), .ZN(n5199) );
  INV_X1 U5429 ( .A(n8804), .ZN(n5200) );
  NAND2_X1 U5430 ( .A1(n8808), .A2(n5452), .ZN(n5448) );
  INV_X1 U5431 ( .A(n8806), .ZN(n5201) );
  INV_X1 U5432 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6964) );
  NOR2_X1 U5433 ( .A1(n6683), .A2(n6502), .ZN(n6503) );
  INV_X1 U5434 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6501) );
  OR2_X1 U5435 ( .A1(n9321), .A2(n9122), .ZN(n8744) );
  NAND2_X1 U5436 ( .A1(n9106), .A2(n9122), .ZN(n5546) );
  OR2_X1 U5437 ( .A1(n9330), .A2(n9158), .ZN(n9118) );
  OR2_X1 U5438 ( .A1(n9162), .A2(n8890), .ZN(n8734) );
  NOR2_X1 U5439 ( .A1(n5477), .A2(n8714), .ZN(n5185) );
  INV_X1 U5440 ( .A(n5061), .ZN(n5477) );
  NAND2_X1 U5441 ( .A1(n9205), .A2(n9213), .ZN(n5557) );
  NAND2_X1 U5442 ( .A1(n7753), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7790) );
  NOR2_X1 U5443 ( .A1(n8777), .A2(n5144), .ZN(n5548) );
  INV_X1 U5444 ( .A(n7763), .ZN(n5144) );
  NOR2_X1 U5445 ( .A1(n5471), .A2(n7442), .ZN(n5470) );
  INV_X1 U5446 ( .A(n7446), .ZN(n5471) );
  NAND2_X1 U5447 ( .A1(n5472), .A2(n7446), .ZN(n5474) );
  NAND2_X1 U5448 ( .A1(n7444), .A2(n5238), .ZN(n7446) );
  NAND2_X1 U5449 ( .A1(n5239), .A2(n8644), .ZN(n5238) );
  NAND2_X1 U5450 ( .A1(n7445), .A2(n8648), .ZN(n5239) );
  AOI21_X1 U5451 ( .B1(n6496), .B2(n6495), .A(n7051), .ZN(n6467) );
  NAND2_X1 U5452 ( .A1(n6457), .A2(n5562), .ZN(n5561) );
  INV_X1 U5453 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6457) );
  INV_X1 U5454 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5562) );
  INV_X1 U5455 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6445) );
  NAND2_X1 U5456 ( .A1(n7643), .A2(n5987), .ZN(n6010) );
  AND2_X1 U5457 ( .A1(n9545), .A2(n5586), .ZN(n5585) );
  NAND2_X1 U5458 ( .A1(n5587), .A2(n6344), .ZN(n5586) );
  INV_X1 U5459 ( .A(n6343), .ZN(n5587) );
  OR2_X1 U5460 ( .A1(n5878), .A2(n5880), .ZN(n5879) );
  XNOR2_X1 U5461 ( .A(n5611), .B(n5913), .ZN(n5853) );
  OAI21_X1 U5462 ( .B1(n10870), .B2(n6300), .A(n5850), .ZN(n5611) );
  AND2_X1 U5463 ( .A1(n7424), .A2(n5943), .ZN(n5574) );
  OR2_X1 U5464 ( .A1(n7673), .A2(n5964), .ZN(n5575) );
  AND2_X1 U5465 ( .A1(n5575), .A2(n5943), .ZN(n5572) );
  AND2_X1 U5466 ( .A1(n7645), .A2(n5581), .ZN(n5580) );
  NAND2_X1 U5467 ( .A1(n7673), .A2(n5964), .ZN(n5581) );
  INV_X1 U5468 ( .A(n10152), .ZN(n8487) );
  NAND2_X1 U5469 ( .A1(n5400), .A2(n5399), .ZN(n5398) );
  INV_X1 U5470 ( .A(n9919), .ZN(n5399) );
  INV_X1 U5471 ( .A(n5393), .ZN(n5389) );
  NAND2_X1 U5472 ( .A1(n9653), .A2(n9970), .ZN(n5627) );
  NOR2_X1 U5473 ( .A1(n10168), .A2(n10175), .ZN(n5309) );
  OR2_X1 U5474 ( .A1(n10175), .A2(n8450), .ZN(n9654) );
  AND2_X1 U5475 ( .A1(n6292), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6306) );
  OR2_X1 U5476 ( .A1(n10216), .A2(n10082), .ZN(n9708) );
  NAND2_X1 U5477 ( .A1(n7276), .A2(n7259), .ZN(n9600) );
  INV_X1 U5478 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10563) );
  INV_X1 U5479 ( .A(n5513), .ZN(n5512) );
  OAI21_X1 U5480 ( .B1(n5516), .B2(n5514), .A(n8342), .ZN(n5513) );
  INV_X1 U5481 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5724) );
  NOR2_X1 U5482 ( .A1(n6258), .A2(n5504), .ZN(n5503) );
  INV_X1 U5483 ( .A(n6236), .ZN(n5504) );
  INV_X1 U5484 ( .A(SI_22_), .ZN(n6260) );
  INV_X1 U5485 ( .A(n5703), .ZN(n5404) );
  NAND2_X1 U5486 ( .A1(n6237), .A2(n5503), .ZN(n5507) );
  OR2_X1 U5487 ( .A1(n6257), .A2(n10484), .ZN(n5506) );
  AND2_X1 U5488 ( .A1(n6143), .A2(n6120), .ZN(n6141) );
  NAND2_X1 U5489 ( .A1(n5043), .A2(n5965), .ZN(n5204) );
  AOI21_X1 U5490 ( .B1(n5043), .B2(n5489), .A(n5092), .ZN(n5484) );
  AND2_X1 U5491 ( .A1(n5696), .A2(n5695), .ZN(n5648) );
  OR2_X1 U5492 ( .A1(n5947), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5967) );
  INV_X1 U5493 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5523) );
  OR2_X1 U5494 ( .A1(n8319), .A2(n10520), .ZN(n8332) );
  OR2_X1 U5495 ( .A1(n6544), .A2(n6658), .ZN(n5327) );
  OR2_X1 U5496 ( .A1(n7104), .A2(n6659), .ZN(n5328) );
  OR2_X1 U5497 ( .A1(n7185), .A2(n8562), .ZN(n6545) );
  NAND2_X1 U5498 ( .A1(n7493), .A2(n5442), .ZN(n5441) );
  INV_X1 U5499 ( .A(n5653), .ZN(n5442) );
  NOR2_X1 U5500 ( .A1(n6580), .A2(n6494), .ZN(n6591) );
  MUX2_X1 U5501 ( .A(n8800), .B(n8799), .S(n8798), .Z(n5215) );
  AND3_X1 U5502 ( .A1(n8269), .A2(n8268), .A3(n8267), .ZN(n8530) );
  NAND2_X1 U5503 ( .A1(n6503), .A2(n5436), .ZN(n7057) );
  NAND2_X1 U5504 ( .A1(n6507), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6511) );
  INV_X1 U5505 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6506) );
  INV_X1 U5506 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6510) );
  NOR2_X1 U5507 ( .A1(n8314), .A2(n8737), .ZN(n9119) );
  AND2_X1 U5508 ( .A1(n8306), .A2(n8295), .ZN(n9138) );
  NAND2_X1 U5509 ( .A1(n5206), .A2(n5205), .ZN(n9153) );
  AND2_X1 U5510 ( .A1(n9154), .A2(n8622), .ZN(n5205) );
  OR2_X1 U5511 ( .A1(n9347), .A2(n8530), .ZN(n8722) );
  AND2_X1 U5512 ( .A1(n5061), .A2(n8719), .ZN(n9207) );
  NOR2_X1 U5513 ( .A1(n9207), .A2(n5556), .ZN(n5555) );
  INV_X1 U5514 ( .A(n5645), .ZN(n5556) );
  NAND2_X1 U5515 ( .A1(n9216), .A2(n9215), .ZN(n9214) );
  AOI21_X1 U5516 ( .B1(n5466), .B2(n5469), .A(n5465), .ZN(n5464) );
  NAND2_X1 U5517 ( .A1(n5459), .A2(n5190), .ZN(n5189) );
  NOR2_X1 U5518 ( .A1(n7998), .A2(n5192), .ZN(n5190) );
  AND2_X1 U5519 ( .A1(n8698), .A2(n8697), .ZN(n9283) );
  INV_X1 U5520 ( .A(n5454), .ZN(n5195) );
  OR2_X1 U5521 ( .A1(n7790), .A2(n7774), .ZN(n7985) );
  NAND2_X1 U5522 ( .A1(n8064), .A2(n5077), .ZN(n8153) );
  AND4_X1 U5523 ( .A1(n7990), .A2(n7989), .A3(n7988), .A4(n7987), .ZN(n8390)
         );
  NAND2_X1 U5524 ( .A1(n7787), .A2(n7786), .ZN(n8028) );
  OR2_X1 U5525 ( .A1(n7529), .A2(n6721), .ZN(n7530) );
  NAND2_X1 U5526 ( .A1(n7443), .A2(n7442), .ZN(n5476) );
  OR2_X1 U5527 ( .A1(n6582), .A2(n6777), .ZN(n9272) );
  NAND2_X1 U5528 ( .A1(n6582), .A2(n7176), .ZN(n9270) );
  NAND2_X1 U5529 ( .A1(n8347), .A2(n8346), .ZN(n9311) );
  OR2_X1 U5530 ( .A1(n10268), .A2(n5037), .ZN(n8347) );
  INV_X1 U5531 ( .A(n9175), .ZN(n9341) );
  NAND2_X1 U5532 ( .A1(n8205), .A2(n8204), .ZN(n9352) );
  NAND2_X1 U5533 ( .A1(n8248), .A2(n8247), .ZN(n9357) );
  NAND2_X1 U5534 ( .A1(n8801), .A2(n10830), .ZN(n10994) );
  OR2_X1 U5535 ( .A1(n10994), .A2(n8811), .ZN(n7234) );
  AND2_X1 U5536 ( .A1(n7029), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7237) );
  AND2_X1 U5537 ( .A1(n6477), .A2(n6476), .ZN(n10700) );
  AND2_X1 U5538 ( .A1(n6780), .A2(n10772), .ZN(n10702) );
  NAND2_X1 U5539 ( .A1(n9449), .A2(n5161), .ZN(n5159) );
  AOI21_X1 U5540 ( .B1(n5161), .B2(n9447), .A(n5090), .ZN(n5160) );
  XNOR2_X1 U5541 ( .A(n5897), .B(n5913), .ZN(n7063) );
  AOI21_X1 U5542 ( .B1(n8422), .B2(n7296), .A(n5780), .ZN(n5781) );
  INV_X1 U5543 ( .A(n6891), .ZN(n5155) );
  NOR2_X1 U5544 ( .A1(n8013), .A2(n8101), .ZN(n5148) );
  XNOR2_X1 U5545 ( .A(n5825), .B(n5913), .ZN(n5830) );
  NAND2_X1 U5546 ( .A1(n7274), .A2(n8416), .ZN(n5823) );
  NAND2_X1 U5547 ( .A1(n5565), .A2(n5566), .ZN(n6189) );
  NAND2_X1 U5548 ( .A1(n5601), .A2(n5597), .ZN(n5170) );
  AND2_X1 U5549 ( .A1(n5600), .A2(n5599), .ZN(n5597) );
  OR2_X1 U5550 ( .A1(n7063), .A2(n7062), .ZN(n5599) );
  AND2_X1 U5551 ( .A1(n9823), .A2(n10030), .ZN(n6417) );
  NAND2_X1 U5552 ( .A1(n5387), .A2(n5384), .ZN(n5383) );
  AND2_X1 U5553 ( .A1(n5396), .A2(n5385), .ZN(n5384) );
  NAND2_X1 U5554 ( .A1(n5391), .A2(n5389), .ZN(n5387) );
  OAI22_X1 U5555 ( .A1(n9790), .A2(n8481), .B1(n5400), .B2(n5052), .ZN(n5396)
         );
  NOR2_X1 U5556 ( .A1(n5398), .A2(n5389), .ZN(n5388) );
  AND2_X1 U5557 ( .A1(n5395), .A2(n5392), .ZN(n5391) );
  NAND2_X1 U5558 ( .A1(n9788), .A2(n5393), .ZN(n5392) );
  NOR2_X1 U5559 ( .A1(n5400), .A2(n8481), .ZN(n5395) );
  AND2_X1 U5560 ( .A1(n9577), .A2(n9751), .ZN(n9919) );
  AOI21_X1 U5561 ( .B1(n5414), .B2(n9980), .A(n5086), .ZN(n5412) );
  AND2_X1 U5562 ( .A1(n9970), .A2(n5106), .ZN(n5414) );
  AND2_X1 U5563 ( .A1(n9656), .A2(n9655), .ZN(n9980) );
  OR2_X1 U5564 ( .A1(n9978), .A2(n9980), .ZN(n5415) );
  NAND2_X1 U5565 ( .A1(n10188), .A2(n10025), .ZN(n5143) );
  NOR2_X1 U5566 ( .A1(n10023), .A2(n5409), .ZN(n5408) );
  INV_X1 U5567 ( .A(n8475), .ZN(n5409) );
  AND2_X1 U5568 ( .A1(n9615), .A2(n9721), .ZN(n10023) );
  NAND2_X1 U5569 ( .A1(n10106), .A2(n5045), .ZN(n10080) );
  NAND2_X1 U5570 ( .A1(n10105), .A2(n10104), .ZN(n10103) );
  NAND2_X1 U5571 ( .A1(n10126), .A2(n9705), .ZN(n10108) );
  AND2_X1 U5572 ( .A1(n9699), .A2(n9695), .ZN(n9782) );
  INV_X1 U5573 ( .A(n9698), .ZN(n5617) );
  NAND2_X1 U5574 ( .A1(n8097), .A2(n9780), .ZN(n8174) );
  NAND2_X1 U5575 ( .A1(n5621), .A2(n9683), .ZN(n8086) );
  NAND2_X1 U5576 ( .A1(n8116), .A2(n9778), .ZN(n5621) );
  AND4_X1 U5577 ( .A1(n6104), .A2(n6103), .A3(n6102), .A4(n6101), .ZN(n9429)
         );
  AND4_X1 U5578 ( .A1(n6032), .A2(n6031), .A3(n6030), .A4(n6029), .ZN(n8117)
         );
  NAND2_X1 U5579 ( .A1(n7865), .A2(n9773), .ZN(n5636) );
  NAND2_X1 U5580 ( .A1(n5410), .A2(n5078), .ZN(n7863) );
  AND2_X1 U5581 ( .A1(n7562), .A2(n9661), .ZN(n5629) );
  AOI21_X1 U5582 ( .B1(n7597), .B2(n9769), .A(n7576), .ZN(n7659) );
  INV_X1 U5583 ( .A(n7608), .ZN(n10921) );
  INV_X1 U5584 ( .A(n5762), .ZN(n9760) );
  NAND2_X1 U5585 ( .A1(n5032), .A2(n5668), .ZN(n8453) );
  NAND2_X1 U5586 ( .A1(n9600), .A2(n5637), .ZN(n7416) );
  NOR2_X1 U5587 ( .A1(n9762), .A2(n5638), .ZN(n5637) );
  INV_X1 U5588 ( .A(n9598), .ZN(n5638) );
  AND2_X1 U5589 ( .A1(n6893), .A2(n9828), .ZN(n10946) );
  NAND2_X1 U5590 ( .A1(n5733), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U5591 ( .A1(n5726), .A2(n5724), .ZN(n5728) );
  NAND2_X1 U5592 ( .A1(n5172), .A2(n5171), .ZN(n5737) );
  AOI21_X1 U5593 ( .B1(n5174), .B2(n10261), .A(n10261), .ZN(n5171) );
  INV_X1 U5594 ( .A(n5175), .ZN(n5174) );
  NAND2_X1 U5595 ( .A1(n5737), .A2(n10628), .ZN(n5758) );
  XNOR2_X1 U5596 ( .A(n5739), .B(P1_IR_REG_20__SCAN_IN), .ZN(n9798) );
  AND4_X1 U5597 ( .A1(n7457), .A2(n7456), .A3(n7455), .A4(n7454), .ZN(n7711)
         );
  NAND2_X1 U5598 ( .A1(n8045), .A2(n8044), .ZN(n9389) );
  NAND2_X1 U5599 ( .A1(n8043), .A2(n8616), .ZN(n8045) );
  XNOR2_X1 U5600 ( .A(n8538), .B(n8536), .ZN(n8842) );
  NAND2_X1 U5601 ( .A1(n5429), .A2(n5428), .ZN(n8901) );
  OR2_X1 U5602 ( .A1(n5062), .A2(n5432), .ZN(n5428) );
  NOR2_X1 U5603 ( .A1(n8509), .A2(n5433), .ZN(n5432) );
  XNOR2_X1 U5604 ( .A(n6545), .B(n6556), .ZN(n7226) );
  AND4_X1 U5605 ( .A1(n8259), .A2(n8258), .A3(n8257), .A4(n8256), .ZN(n9233)
         );
  NAND2_X1 U5606 ( .A1(n8529), .A2(n8859), .ZN(n8913) );
  AND4_X1 U5607 ( .A1(n8055), .A2(n8054), .A3(n8053), .A4(n8052), .ZN(n8881)
         );
  OAI21_X1 U5608 ( .B1(n7031), .B2(n6574), .A(n6573), .ZN(n7358) );
  OR2_X1 U5609 ( .A1(n7716), .A2(n7715), .ZN(n7717) );
  NOR2_X1 U5610 ( .A1(n8233), .A2(n6590), .ZN(n5446) );
  NAND2_X1 U5611 ( .A1(n8156), .A2(n8155), .ZN(n9383) );
  INV_X1 U5612 ( .A(n8530), .ZN(n9197) );
  AOI21_X1 U5613 ( .B1(n5535), .B2(n5041), .A(n5055), .ZN(n5530) );
  AOI21_X1 U5614 ( .B1(n8377), .B2(n10822), .A(n5242), .ZN(n9314) );
  INV_X1 U5615 ( .A(n5243), .ZN(n5242) );
  AOI22_X1 U5616 ( .A1(n8979), .A2(n9254), .B1(n9093), .B2(n8977), .ZN(n5243)
         );
  NAND2_X1 U5617 ( .A1(n10829), .A2(n10980), .ZN(n9300) );
  NAND2_X1 U5618 ( .A1(n10829), .A2(n7205), .ZN(n10819) );
  AND2_X1 U5619 ( .A1(n5559), .A2(n5233), .ZN(n5232) );
  AND2_X1 U5620 ( .A1(n6530), .A2(n5234), .ZN(n5233) );
  INV_X1 U5621 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5234) );
  AND4_X1 U5622 ( .A1(n5959), .A2(n5958), .A3(n5957), .A4(n5956), .ZN(n7564)
         );
  NAND2_X1 U5623 ( .A1(n6063), .A2(n5150), .ZN(n5149) );
  NAND2_X1 U5624 ( .A1(n8138), .A2(n5152), .ZN(n5151) );
  INV_X1 U5625 ( .A(n8136), .ZN(n5150) );
  AND2_X1 U5626 ( .A1(n6313), .A2(n6312), .ZN(n9974) );
  NAND2_X1 U5627 ( .A1(n5589), .A2(n5592), .ZN(n9503) );
  AOI22_X1 U5628 ( .A1(n5094), .A2(n9438), .B1(n9439), .B2(n5593), .ZN(n5592)
         );
  AND4_X1 U5629 ( .A1(n6003), .A2(n6002), .A3(n6001), .A4(n6000), .ZN(n7866)
         );
  NAND2_X1 U5630 ( .A1(n6221), .A2(n6220), .ZN(n10198) );
  NAND2_X1 U5631 ( .A1(n6181), .A2(n6180), .ZN(n10096) );
  INV_X1 U5632 ( .A(n9934), .ZN(n9840) );
  INV_X1 U5633 ( .A(n9974), .ZN(n10002) );
  INV_X1 U5634 ( .A(n9451), .ZN(n10068) );
  INV_X1 U5635 ( .A(n8140), .ZN(n9841) );
  INV_X1 U5636 ( .A(n7957), .ZN(n9844) );
  NAND2_X1 U5637 ( .A1(n9572), .A2(n9571), .ZN(n10149) );
  XNOR2_X1 U5638 ( .A(n5302), .B(n5301), .ZN(n10150) );
  INV_X1 U5639 ( .A(n10149), .ZN(n5301) );
  NOR2_X1 U5640 ( .A1(n9906), .A2(n9900), .ZN(n5302) );
  OR3_X1 U5641 ( .A1(n10923), .A2(n9760), .A3(n10666), .ZN(n10090) );
  AND2_X1 U5642 ( .A1(n6410), .A2(n6409), .ZN(n10259) );
  NAND2_X1 U5643 ( .A1(n5479), .A2(n5481), .ZN(n6197) );
  XNOR2_X1 U5644 ( .A(n5761), .B(P1_IR_REG_19__SCAN_IN), .ZN(n10659) );
  NAND2_X1 U5645 ( .A1(n5736), .A2(n5647), .ZN(n5760) );
  OAI211_X1 U5646 ( .C1(n10651), .C2(n10650), .A(n10649), .B(n10648), .ZN(
        n10653) );
  OAI21_X1 U5647 ( .B1(n10439), .B2(n10438), .A(n5134), .ZN(n5265) );
  INV_X1 U5648 ( .A(keyinput_130), .ZN(n5338) );
  INV_X1 U5649 ( .A(keyinput_132), .ZN(n5334) );
  INV_X1 U5650 ( .A(SI_24_), .ZN(n10471) );
  NAND2_X1 U5651 ( .A1(n10482), .A2(n10481), .ZN(n5347) );
  AOI21_X1 U5652 ( .B1(SI_25_), .B2(keyinput_135), .A(n10477), .ZN(n10482) );
  XNOR2_X1 U5653 ( .A(n5346), .B(SI_22_), .ZN(n5345) );
  INV_X1 U5654 ( .A(keyinput_138), .ZN(n5346) );
  NAND2_X1 U5655 ( .A1(n5268), .A2(SI_29_), .ZN(n5267) );
  NAND2_X1 U5656 ( .A1(SI_28_), .A2(n5270), .ZN(n5269) );
  NAND2_X1 U5657 ( .A1(n10316), .A2(keyinput_3), .ZN(n5266) );
  OAI22_X1 U5658 ( .A1(n10485), .A2(keyinput_140), .B1(n10486), .B2(SI_20_), 
        .ZN(n5340) );
  NAND2_X1 U5659 ( .A1(n5344), .A2(n5342), .ZN(n5341) );
  INV_X1 U5660 ( .A(n5343), .ZN(n5342) );
  NAND2_X1 U5661 ( .A1(n5347), .A2(n5345), .ZN(n5344) );
  OAI22_X1 U5662 ( .A1(n10483), .A2(n10484), .B1(SI_21_), .B2(keyinput_139), 
        .ZN(n5343) );
  AOI22_X1 U5663 ( .A1(n10322), .A2(n10484), .B1(keyinput_11), .B2(SI_21_), 
        .ZN(n5290) );
  NAND2_X1 U5664 ( .A1(n10489), .A2(n10324), .ZN(n5285) );
  NAND2_X1 U5665 ( .A1(keyinput_13), .A2(SI_19_), .ZN(n5284) );
  NAND2_X1 U5666 ( .A1(n10485), .A2(keyinput_12), .ZN(n5288) );
  NAND2_X1 U5667 ( .A1(n10323), .A2(SI_20_), .ZN(n5287) );
  NAND2_X1 U5668 ( .A1(n5361), .A2(n5360), .ZN(n5359) );
  NOR2_X1 U5669 ( .A1(n10492), .A2(n10493), .ZN(n5360) );
  NAND2_X1 U5670 ( .A1(n10494), .A2(n10495), .ZN(n5361) );
  INV_X1 U5671 ( .A(n10496), .ZN(n5358) );
  INV_X1 U5672 ( .A(keyinput_149), .ZN(n5356) );
  NAND2_X1 U5673 ( .A1(n10498), .A2(keyinput_150), .ZN(n5353) );
  NAND2_X1 U5674 ( .A1(n10499), .A2(SI_10_), .ZN(n5354) );
  NAND2_X1 U5675 ( .A1(n10335), .A2(n10334), .ZN(n5258) );
  NOR2_X1 U5676 ( .A1(n10333), .A2(n5257), .ZN(n5256) );
  AND2_X1 U5677 ( .A1(n10497), .A2(keyinput_21), .ZN(n5257) );
  AOI21_X1 U5678 ( .B1(n5357), .B2(n5355), .A(n5352), .ZN(n10506) );
  NAND2_X1 U5679 ( .A1(n5354), .A2(n5353), .ZN(n5352) );
  XNOR2_X1 U5680 ( .A(n10497), .B(n5356), .ZN(n5355) );
  NAND2_X1 U5681 ( .A1(n5359), .A2(n5358), .ZN(n5357) );
  NAND2_X1 U5682 ( .A1(n5252), .A2(n5251), .ZN(n5250) );
  AND2_X1 U5683 ( .A1(n10341), .A2(n10340), .ZN(n5251) );
  NAND2_X1 U5684 ( .A1(n5253), .A2(n5123), .ZN(n5252) );
  NAND2_X1 U5685 ( .A1(n10517), .A2(n10518), .ZN(n5371) );
  INV_X1 U5686 ( .A(n10516), .ZN(n5370) );
  NAND2_X1 U5687 ( .A1(n5225), .A2(n5224), .ZN(n8673) );
  NOR2_X1 U5688 ( .A1(n8665), .A2(n8666), .ZN(n5224) );
  NAND2_X1 U5689 ( .A1(n10348), .A2(n10349), .ZN(n5282) );
  INV_X1 U5690 ( .A(n10347), .ZN(n5281) );
  AOI21_X1 U5691 ( .B1(n5367), .B2(n5364), .A(n5362), .ZN(n10531) );
  AND2_X1 U5692 ( .A1(n10550), .A2(n5351), .ZN(n5350) );
  XNOR2_X1 U5693 ( .A(n10286), .B(keyinput_195), .ZN(n5351) );
  AOI21_X1 U5694 ( .B1(n5278), .B2(n5275), .A(n5273), .ZN(n10358) );
  NAND2_X1 U5695 ( .A1(n5219), .A2(n5218), .ZN(n5217) );
  NOR3_X1 U5696 ( .A1(n10374), .A2(n10373), .A3(n5249), .ZN(n5248) );
  OAI21_X1 U5697 ( .B1(keyinput_66), .B2(P2_DATAO_REG_30__SCAN_IN), .A(n10370), 
        .ZN(n5249) );
  AOI211_X1 U5698 ( .C1(n5348), .C2(n10560), .A(n10558), .B(n10559), .ZN(
        n10565) );
  INV_X1 U5699 ( .A(keyinput_214), .ZN(n5376) );
  NAND2_X1 U5700 ( .A1(n5244), .A2(n10382), .ZN(n10383) );
  NAND2_X1 U5701 ( .A1(n5245), .A2(n5058), .ZN(n5244) );
  AOI21_X1 U5702 ( .B1(n5374), .B2(n5373), .A(n5372), .ZN(n10595) );
  NAND2_X1 U5703 ( .A1(n5130), .A2(n5059), .ZN(n5372) );
  NAND2_X1 U5704 ( .A1(n5229), .A2(n8723), .ZN(n5228) );
  AOI21_X1 U5705 ( .B1(n5231), .B2(n8722), .A(n8721), .ZN(n5230) );
  OAI21_X1 U5706 ( .B1(n5260), .B2(n5259), .A(n5133), .ZN(n10394) );
  INV_X1 U5707 ( .A(SI_25_), .ZN(n10311) );
  INV_X1 U5708 ( .A(SI_15_), .ZN(n10491) );
  INV_X1 U5709 ( .A(SI_12_), .ZN(n10467) );
  INV_X1 U5710 ( .A(SI_10_), .ZN(n10498) );
  OR2_X1 U5711 ( .A1(n9094), .A2(n8807), .ZN(n5452) );
  NAND2_X1 U5712 ( .A1(n5213), .A2(n5211), .ZN(n5210) );
  NAND2_X1 U5713 ( .A1(n5212), .A2(n8760), .ZN(n5211) );
  INV_X1 U5714 ( .A(n8746), .ZN(n5212) );
  AND2_X1 U5715 ( .A1(n8750), .A2(n8752), .ZN(n5209) );
  NAND2_X1 U5716 ( .A1(n6505), .A2(n5438), .ZN(n5437) );
  INV_X1 U5717 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5438) );
  AND3_X1 U5718 ( .A1(n6960), .A2(n6964), .A3(n6504), .ZN(n6505) );
  INV_X1 U5719 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U5720 ( .A1(n6499), .A2(n6500), .ZN(n6683) );
  INV_X1 U5721 ( .A(n6372), .ZN(n6424) );
  NAND2_X1 U5722 ( .A1(n5515), .A2(n8191), .ZN(n5514) );
  INV_X1 U5723 ( .A(n8338), .ZN(n5515) );
  AND2_X1 U5724 ( .A1(n5646), .A2(n5707), .ZN(n5640) );
  NOR2_X1 U5725 ( .A1(n5703), .A2(n5713), .ZN(n5305) );
  INV_X1 U5726 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n10420) );
  AND2_X1 U5727 ( .A1(n10628), .A2(keyinput_240), .ZN(n5381) );
  AOI22_X1 U5728 ( .A1(n10630), .A2(n10629), .B1(keyinput_241), .B2(
        P1_IR_REG_22__SCAN_IN), .ZN(n5380) );
  XNOR2_X1 U5729 ( .A(n10628), .B(keyinput_112), .ZN(n5295) );
  NOR2_X1 U5730 ( .A1(n10427), .A2(n10426), .ZN(n5292) );
  NOR2_X1 U5731 ( .A1(n5495), .A2(n5492), .ZN(n5491) );
  INV_X1 U5732 ( .A(n6044), .ZN(n5492) );
  INV_X1 U5733 ( .A(n5496), .ZN(n5495) );
  NOR2_X1 U5734 ( .A1(n6086), .A2(n5497), .ZN(n5496) );
  INV_X1 U5735 ( .A(n6065), .ZN(n5497) );
  INV_X1 U5736 ( .A(n5649), .ZN(n5494) );
  INV_X1 U5737 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5520) );
  INV_X1 U5738 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5519) );
  INV_X1 U5739 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5521) );
  AND2_X1 U5740 ( .A1(n8888), .A2(n8399), .ZN(n8400) );
  NOR2_X1 U5741 ( .A1(n5437), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5436) );
  INV_X1 U5742 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7774) );
  NOR2_X1 U5743 ( .A1(n8781), .A2(n5462), .ZN(n5461) );
  AND2_X1 U5744 ( .A1(n6922), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7753) );
  CLKBUF_X1 U5745 ( .A(n7798), .Z(n7887) );
  NOR2_X1 U5746 ( .A1(n5551), .A2(n7548), .ZN(n5550) );
  INV_X1 U5747 ( .A(n7521), .ZN(n5551) );
  NAND2_X1 U5748 ( .A1(n7215), .A2(n5063), .ZN(n5322) );
  NAND2_X1 U5749 ( .A1(n10816), .A2(n7392), .ZN(n7391) );
  NAND2_X1 U5750 ( .A1(n7185), .A2(n7400), .ZN(n7392) );
  NOR2_X1 U5751 ( .A1(n8002), .A2(n8028), .ZN(n8003) );
  NAND2_X1 U5752 ( .A1(n6462), .A2(n6461), .ZN(n6468) );
  INV_X1 U5753 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6461) );
  INV_X1 U5754 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6960) );
  INV_X1 U5755 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6500) );
  INV_X1 U5756 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6692) );
  INV_X1 U5757 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6695) );
  INV_X1 U5758 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6447) );
  INV_X1 U5759 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6446) );
  INV_X1 U5760 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5972) );
  NOR2_X1 U5761 ( .A1(n5607), .A2(n5610), .ZN(n5606) );
  INV_X1 U5762 ( .A(n5608), .ZN(n5607) );
  INV_X1 U5763 ( .A(n5646), .ZN(n5610) );
  AND3_X1 U5764 ( .A1(n5072), .A2(n5304), .A3(n5305), .ZN(n5712) );
  AND2_X1 U5765 ( .A1(n5306), .A2(n5640), .ZN(n5304) );
  INV_X1 U5766 ( .A(n8481), .ZN(n5397) );
  OR2_X1 U5767 ( .A1(n5398), .A2(n5386), .ZN(n5385) );
  NAND2_X1 U5768 ( .A1(n9788), .A2(n5393), .ZN(n5386) );
  AND2_X1 U5769 ( .A1(n10158), .A2(n9840), .ZN(n8481) );
  OR2_X1 U5770 ( .A1(n10163), .A2(n9547), .ZN(n9649) );
  NOR2_X1 U5771 ( .A1(n10163), .A2(n5308), .ZN(n5307) );
  INV_X1 U5772 ( .A(n5309), .ZN(n5308) );
  INV_X1 U5773 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6154) );
  INV_X1 U5774 ( .A(n9780), .ZN(n5620) );
  NAND2_X1 U5775 ( .A1(n5634), .A2(n5632), .ZN(n5631) );
  NAND2_X1 U5776 ( .A1(n7814), .A2(n7810), .ZN(n7870) );
  NOR2_X1 U5777 ( .A1(n7471), .A2(n7500), .ZN(n7514) );
  NAND2_X1 U5778 ( .A1(n9606), .A2(n9608), .ZN(n7484) );
  NOR2_X1 U5779 ( .A1(n8192), .A2(n5517), .ZN(n5516) );
  INV_X1 U5780 ( .A(n6367), .ZN(n5517) );
  INV_X1 U5781 ( .A(SI_27_), .ZN(n10474) );
  AND2_X1 U5782 ( .A1(n6367), .A2(n6350), .ZN(n6365) );
  NAND2_X1 U5783 ( .A1(n5379), .A2(n5377), .ZN(n10641) );
  NOR2_X1 U5784 ( .A1(n10632), .A2(n5378), .ZN(n5377) );
  OAI21_X1 U5785 ( .B1(n10627), .B2(n5381), .A(n5380), .ZN(n5379) );
  XNOR2_X1 U5786 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_243), .ZN(n5378) );
  AOI21_X1 U5787 ( .B1(n5294), .B2(n5293), .A(n5291), .ZN(n10431) );
  AOI22_X1 U5788 ( .A1(n10630), .A2(n10425), .B1(keyinput_113), .B2(
        P1_IR_REG_22__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U5789 ( .A1(n5292), .A2(n5132), .ZN(n5291) );
  NAND2_X1 U5790 ( .A1(n10424), .A2(n5295), .ZN(n5294) );
  AOI21_X1 U5791 ( .B1(n5648), .B2(n5488), .A(n5487), .ZN(n5486) );
  INV_X1 U5792 ( .A(n5696), .ZN(n5487) );
  INV_X1 U5793 ( .A(n5691), .ZN(n5488) );
  INV_X1 U5794 ( .A(n5648), .ZN(n5489) );
  OAI21_X1 U5795 ( .B1(n5668), .B2(n5137), .A(n5136), .ZN(n5665) );
  NAND2_X1 U5796 ( .A1(n5668), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5136) );
  INV_X1 U5797 ( .A(n8549), .ZN(n5444) );
  OAI21_X1 U5798 ( .B1(n8529), .B2(n5418), .A(n5416), .ZN(n8538) );
  AOI21_X1 U5799 ( .B1(n8532), .B2(n5417), .A(n5053), .ZN(n5416) );
  INV_X1 U5800 ( .A(n8532), .ZN(n5418) );
  NAND2_X1 U5801 ( .A1(n6927), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8281) );
  INV_X1 U5802 ( .A(n8264), .ZN(n6927) );
  INV_X1 U5803 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10524) );
  NOR2_X1 U5804 ( .A1(n5062), .A2(n5431), .ZN(n5430) );
  INV_X1 U5805 ( .A(n8400), .ZN(n5431) );
  AOI21_X1 U5806 ( .B1(n5423), .B2(n5044), .A(n5121), .ZN(n5422) );
  INV_X1 U5807 ( .A(n5426), .ZN(n5423) );
  INV_X1 U5808 ( .A(n8870), .ZN(n5445) );
  OR2_X1 U5809 ( .A1(n8403), .A2(n8402), .ZN(n5643) );
  NAND2_X1 U5810 ( .A1(n8877), .A2(n8400), .ZN(n8884) );
  INV_X1 U5811 ( .A(n10959), .ZN(n7762) );
  NAND2_X1 U5812 ( .A1(n7842), .A2(n5426), .ZN(n5424) );
  AOI21_X1 U5813 ( .B1(n5198), .B2(n5201), .A(n5447), .ZN(n5196) );
  AND2_X1 U5814 ( .A1(n8313), .A2(n8312), .ZN(n8871) );
  AND4_X1 U5815 ( .A1(n6727), .A2(n6726), .A3(n6725), .A4(n6724), .ZN(n8929)
         );
  AOI21_X1 U5816 ( .B1(n8266), .B2(P2_REG1_REG_1__SCAN_IN), .A(n5046), .ZN(
        n5236) );
  AOI21_X1 U5817 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7749), .A(n7620), .ZN(
        n9001) );
  AOI21_X1 U5818 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7785), .A(n7693), .ZN(
        n7696) );
  NOR2_X1 U5819 ( .A1(n6903), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6957) );
  AND2_X1 U5820 ( .A1(n8820), .A2(n8796), .ZN(n7176) );
  NAND2_X1 U5821 ( .A1(n8585), .A2(n8793), .ZN(n8590) );
  AND2_X1 U5822 ( .A1(n8328), .A2(n8327), .ZN(n9122) );
  NAND2_X1 U5823 ( .A1(n9153), .A2(n8734), .ZN(n9141) );
  NAND2_X1 U5824 ( .A1(n9141), .A2(n9136), .ZN(n9145) );
  AND2_X1 U5825 ( .A1(n8734), .A2(n8730), .ZN(n9154) );
  AOI21_X1 U5826 ( .B1(n9138), .B2(n8353), .A(n8299), .ZN(n9158) );
  NOR2_X1 U5827 ( .A1(n8791), .A2(n5208), .ZN(n5207) );
  INV_X1 U5828 ( .A(n8722), .ZN(n5208) );
  AOI21_X1 U5829 ( .B1(n5185), .B2(n9215), .A(n5183), .ZN(n5182) );
  INV_X1 U5830 ( .A(n5185), .ZN(n5184) );
  INV_X1 U5831 ( .A(n8719), .ZN(n5183) );
  NAND2_X1 U5832 ( .A1(n5554), .A2(n5557), .ZN(n5553) );
  INV_X1 U5833 ( .A(n5555), .ZN(n5554) );
  NOR2_X1 U5834 ( .A1(n5042), .A2(n5318), .ZN(n5317) );
  NAND2_X1 U5835 ( .A1(n9236), .A2(n9221), .ZN(n5318) );
  OR2_X1 U5836 ( .A1(n8238), .A2(n10524), .ZN(n8250) );
  NAND2_X1 U5837 ( .A1(n6926), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8252) );
  INV_X1 U5838 ( .A(n8250), .ZN(n6926) );
  NOR2_X1 U5839 ( .A1(n5316), .A2(n9296), .ZN(n9237) );
  OR2_X1 U5840 ( .A1(n5042), .A2(n9361), .ZN(n5316) );
  NAND2_X1 U5841 ( .A1(n6925), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8238) );
  INV_X1 U5842 ( .A(n8225), .ZN(n6925) );
  NAND2_X1 U5843 ( .A1(n8364), .A2(n8363), .ZN(n9246) );
  AND4_X1 U5844 ( .A1(n8168), .A2(n8167), .A3(n8166), .A4(n8165), .ZN(n9273)
         );
  AOI21_X1 U5845 ( .B1(n5459), .B2(n5458), .A(n5457), .ZN(n5456) );
  INV_X1 U5846 ( .A(n8689), .ZN(n5457) );
  INV_X1 U5847 ( .A(n5461), .ZN(n5458) );
  AND2_X1 U5848 ( .A1(n8692), .A2(n8691), .ZN(n8785) );
  INV_X1 U5849 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10521) );
  NAND2_X1 U5850 ( .A1(n8003), .A2(n10993), .ZN(n8058) );
  AND4_X1 U5851 ( .A1(n7759), .A2(n7758), .A3(n7757), .A4(n7756), .ZN(n8033)
         );
  NAND2_X1 U5852 ( .A1(n7780), .A2(n8669), .ZN(n7881) );
  NAND2_X1 U5853 ( .A1(n5324), .A2(n5323), .ZN(n8002) );
  INV_X1 U5854 ( .A(n10970), .ZN(n5323) );
  AND2_X1 U5855 ( .A1(n8668), .A2(n8669), .ZN(n8777) );
  NAND2_X1 U5856 ( .A1(n7747), .A2(n8667), .ZN(n7780) );
  AND2_X1 U5857 ( .A1(n7631), .A2(n8661), .ZN(n7549) );
  AND2_X1 U5858 ( .A1(n8672), .A2(n8667), .ZN(n8772) );
  NAND2_X1 U5859 ( .A1(n7549), .A2(n8772), .ZN(n7747) );
  NAND2_X1 U5860 ( .A1(n7522), .A2(n7521), .ZN(n7634) );
  AND2_X1 U5861 ( .A1(n5473), .A2(n5237), .ZN(n7632) );
  AOI21_X1 U5862 ( .B1(n5470), .B2(n5472), .A(n5069), .ZN(n5473) );
  OR2_X1 U5863 ( .A1(n7443), .A2(n5474), .ZN(n5237) );
  NOR2_X1 U5864 ( .A1(n5322), .A2(n7365), .ZN(n7434) );
  INV_X1 U5865 ( .A(n8995), .ZN(n7384) );
  NAND2_X1 U5866 ( .A1(n7215), .A2(n10864), .ZN(n7311) );
  AND2_X1 U5867 ( .A1(n8627), .A2(n8624), .ZN(n8623) );
  NAND2_X1 U5868 ( .A1(n8293), .A2(n8292), .ZN(n9330) );
  CLKBUF_X1 U5869 ( .A(n9170), .Z(n9346) );
  OAI21_X1 U5870 ( .B1(n8364), .B2(n5469), .A(n5466), .ZN(n9232) );
  AND2_X1 U5871 ( .A1(n8007), .A2(n8006), .ZN(n8008) );
  AND3_X1 U5872 ( .A1(n7330), .A2(n7329), .A3(n7328), .ZN(n10912) );
  NAND2_X1 U5873 ( .A1(n10851), .A2(n10817), .ZN(n10848) );
  INV_X1 U5874 ( .A(n10971), .ZN(n10992) );
  AND2_X1 U5875 ( .A1(n8620), .A2(n8807), .ZN(n10830) );
  INV_X1 U5876 ( .A(n10990), .ZN(n10980) );
  INV_X1 U5877 ( .A(n8133), .ZN(n6477) );
  AND2_X1 U5878 ( .A1(n6455), .A2(n5560), .ZN(n5559) );
  NOR2_X1 U5879 ( .A1(n5561), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5560) );
  INV_X1 U5880 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6530) );
  NOR2_X1 U5881 ( .A1(n5561), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U5882 ( .A1(n6460), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6496) );
  INV_X1 U5883 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6495) );
  OR2_X1 U5884 ( .A1(n6499), .A2(n7051), .ZN(n6677) );
  AND2_X1 U5885 ( .A1(n6662), .A2(n6663), .ZN(n6809) );
  NAND2_X1 U5886 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6543) );
  NAND2_X1 U5887 ( .A1(n5656), .A2(n5655), .ZN(n6547) );
  NOR2_X1 U5888 ( .A1(n5089), .A2(n5169), .ZN(n5168) );
  INV_X1 U5889 ( .A(n5598), .ZN(n5169) );
  INV_X1 U5890 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U5891 ( .A1(n5153), .A2(n8136), .ZN(n5152) );
  XNOR2_X1 U5892 ( .A(n5187), .B(n6066), .ZN(n8043) );
  NAND2_X1 U5893 ( .A1(n5188), .A2(n6065), .ZN(n5187) );
  NAND2_X1 U5894 ( .A1(n6064), .A2(n5649), .ZN(n5188) );
  AOI21_X1 U5895 ( .B1(n5585), .B2(n5588), .A(n5116), .ZN(n5584) );
  NAND2_X1 U5896 ( .A1(n5577), .A2(n5943), .ZN(n5582) );
  NAND2_X1 U5897 ( .A1(n5579), .A2(n5578), .ZN(n5577) );
  OR2_X1 U5898 ( .A1(n5882), .A2(n8382), .ZN(n5600) );
  NOR2_X1 U5899 ( .A1(n5076), .A2(n5591), .ZN(n5590) );
  INV_X1 U5900 ( .A(n9524), .ZN(n5591) );
  AND2_X1 U5901 ( .A1(n5580), .A2(n5573), .ZN(n5576) );
  NAND2_X1 U5902 ( .A1(n5574), .A2(n5575), .ZN(n5573) );
  OR2_X1 U5903 ( .A1(n6222), .A2(n9516), .ZN(n6241) );
  INV_X1 U5904 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9516) );
  INV_X1 U5905 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6055) );
  AOI21_X1 U5906 ( .B1(n5158), .B2(n5162), .A(n5115), .ZN(n5156) );
  INV_X1 U5907 ( .A(n5158), .ZN(n5157) );
  NAND2_X1 U5908 ( .A1(n9523), .A2(n9524), .ZN(n9522) );
  INV_X1 U5909 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5749) );
  NOR2_X1 U5910 ( .A1(n5998), .A2(n5749), .ZN(n6027) );
  OR2_X1 U5911 ( .A1(n5996), .A2(n6885), .ZN(n5998) );
  OR2_X1 U5912 ( .A1(n7946), .A2(n7941), .ZN(n5605) );
  INV_X1 U5913 ( .A(n6935), .ZN(n5777) );
  XNOR2_X1 U5914 ( .A(n5798), .B(n7288), .ZN(n5801) );
  INV_X1 U5915 ( .A(n6188), .ZN(n5564) );
  NAND2_X1 U5916 ( .A1(n7063), .A2(n7062), .ZN(n5598) );
  INV_X1 U5917 ( .A(n5778), .ZN(n8420) );
  AND2_X1 U5918 ( .A1(n9646), .A2(n9819), .ZN(n9827) );
  AND4_X1 U5919 ( .A1(n6337), .A2(n6336), .A3(n6335), .A4(n6334), .ZN(n8450)
         );
  NAND2_X1 U5920 ( .A1(n5394), .A2(n9547), .ZN(n5393) );
  AND2_X1 U5921 ( .A1(n9649), .A2(n9650), .ZN(n9788) );
  AOI21_X1 U5922 ( .B1(n5625), .B2(n8451), .A(n5624), .ZN(n5623) );
  INV_X1 U5923 ( .A(n6332), .ZN(n6333) );
  NAND2_X1 U5924 ( .A1(n9986), .A2(n9964), .ZN(n9961) );
  AND2_X1 U5925 ( .A1(n9733), .A2(n9732), .ZN(n10001) );
  INV_X1 U5926 ( .A(n9527), .ZN(n10010) );
  AND2_X1 U5927 ( .A1(n5049), .A2(n5314), .ZN(n5313) );
  NAND2_X1 U5928 ( .A1(n5406), .A2(n5060), .ZN(n5405) );
  INV_X1 U5929 ( .A(n5408), .ZN(n5406) );
  NAND2_X1 U5930 ( .A1(n10114), .A2(n5049), .ZN(n10048) );
  AND2_X1 U5931 ( .A1(n10114), .A2(n5065), .ZN(n10061) );
  AND2_X1 U5932 ( .A1(n10114), .A2(n10208), .ZN(n10089) );
  NAND2_X1 U5933 ( .A1(n10106), .A2(n9708), .ZN(n10078) );
  AND3_X1 U5934 ( .A1(n6207), .A2(n6206), .A3(n6205), .ZN(n10084) );
  NAND2_X1 U5935 ( .A1(n6124), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6155) );
  INV_X1 U5936 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7143) );
  NOR2_X1 U5937 ( .A1(n6075), .A2(n7143), .ZN(n6098) );
  OR2_X1 U5938 ( .A1(n6056), .A2(n6055), .ZN(n6075) );
  AND2_X1 U5939 ( .A1(n8122), .A2(n10983), .ZN(n8124) );
  AND4_X1 U5940 ( .A1(n6081), .A2(n6080), .A3(n6079), .A4(n6078), .ZN(n8140)
         );
  OR2_X1 U5941 ( .A1(n7870), .A2(n8020), .ZN(n7965) );
  AND4_X1 U5942 ( .A1(n5754), .A2(n5753), .A3(n5752), .A4(n5751), .ZN(n7957)
         );
  NAND2_X1 U5943 ( .A1(n5636), .A2(n5634), .ZN(n8084) );
  NOR2_X1 U5944 ( .A1(n7667), .A2(n10945), .ZN(n7810) );
  NAND2_X1 U5945 ( .A1(n9802), .A2(n9661), .ZN(n7662) );
  NAND2_X1 U5946 ( .A1(n5312), .A2(n5311), .ZN(n7667) );
  CLKBUF_X1 U5947 ( .A(n7559), .Z(n7509) );
  INV_X1 U5948 ( .A(n7484), .ZN(n9766) );
  NAND2_X1 U5949 ( .A1(n7412), .A2(n7411), .ZN(n7471) );
  NAND2_X1 U5950 ( .A1(n9600), .A2(n9598), .ZN(n7260) );
  NOR2_X1 U5951 ( .A1(n7274), .A2(n7294), .ZN(n7273) );
  AND2_X1 U5952 ( .A1(n7273), .A2(n10870), .ZN(n7412) );
  NAND2_X1 U5953 ( .A1(n6202), .A2(n6201), .ZN(n10203) );
  NAND2_X1 U5954 ( .A1(n10103), .A2(n8472), .ZN(n10074) );
  NAND2_X1 U5955 ( .A1(n6151), .A2(n6150), .ZN(n10216) );
  NAND2_X1 U5956 ( .A1(n6123), .A2(n6122), .ZN(n10223) );
  AND2_X1 U5957 ( .A1(n7255), .A2(n10923), .ZN(n10232) );
  INV_X1 U5958 ( .A(n11009), .ZN(n11021) );
  INV_X1 U5959 ( .A(n10946), .ZN(n11018) );
  INV_X1 U5960 ( .A(SI_29_), .ZN(n10316) );
  CLKBUF_X1 U5961 ( .A(n6435), .Z(n6979) );
  XNOR2_X1 U5962 ( .A(n8339), .B(n8338), .ZN(n8413) );
  NAND2_X1 U5963 ( .A1(n5511), .A2(n8191), .ZN(n8339) );
  NAND2_X1 U5964 ( .A1(n6368), .A2(n5516), .ZN(n5511) );
  OAI21_X1 U5965 ( .B1(n6237), .B2(n5502), .A(n5498), .ZN(n6288) );
  AOI21_X1 U5966 ( .B1(n5500), .B2(n5501), .A(n5499), .ZN(n5498) );
  INV_X1 U5967 ( .A(n6281), .ZN(n5499) );
  INV_X1 U5968 ( .A(n5503), .ZN(n5500) );
  AND2_X1 U5969 ( .A1(n6302), .A2(n6286), .ZN(n6287) );
  NAND2_X1 U5970 ( .A1(n5507), .A2(n5501), .ZN(n6282) );
  NAND2_X1 U5971 ( .A1(n5507), .A2(n5506), .ZN(n6265) );
  NAND2_X1 U5972 ( .A1(n6237), .A2(n6236), .ZN(n6259) );
  AOI21_X1 U5973 ( .B1(n5483), .B2(n5482), .A(n5117), .ZN(n5481) );
  INV_X1 U5974 ( .A(n6172), .ZN(n5482) );
  NAND2_X1 U5975 ( .A1(n5480), .A2(n5483), .ZN(n5479) );
  INV_X1 U5976 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n10415) );
  NAND2_X1 U5977 ( .A1(n5203), .A2(n5064), .ZN(n6043) );
  OR2_X1 U5978 ( .A1(n5967), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U5979 ( .A1(n5692), .A2(n5691), .ZN(n5988) );
  CLKBUF_X1 U5980 ( .A(n5713), .Z(n5714) );
  AND2_X1 U5981 ( .A1(n5698), .A2(n5697), .ZN(n5865) );
  NOR2_X1 U5982 ( .A1(n7491), .A2(n5653), .ZN(n7494) );
  AND2_X1 U5983 ( .A1(n8288), .A2(n8287), .ZN(n8890) );
  NOR2_X1 U5984 ( .A1(n7839), .A2(n7838), .ZN(n7842) );
  NAND2_X1 U5985 ( .A1(n7842), .A2(n7841), .ZN(n8925) );
  AND2_X1 U5986 ( .A1(n8348), .A2(n8333), .ZN(n8582) );
  INV_X1 U5987 ( .A(n7640), .ZN(n7704) );
  AND4_X1 U5988 ( .A1(n7535), .A2(n7534), .A3(n7533), .A4(n7532), .ZN(n7761)
         );
  NAND2_X1 U5989 ( .A1(n7226), .A2(n6555), .ZN(n7219) );
  AND2_X1 U5990 ( .A1(n7220), .A2(n6554), .ZN(n6555) );
  INV_X1 U5991 ( .A(n7398), .ZN(n6553) );
  AND4_X1 U5992 ( .A1(n7779), .A2(n7778), .A3(n7777), .A4(n7776), .ZN(n8596)
         );
  NAND2_X1 U5993 ( .A1(n8892), .A2(n8544), .ZN(n8869) );
  NAND2_X1 U5994 ( .A1(n8884), .A2(n5643), .ZN(n8943) );
  NAND2_X1 U5995 ( .A1(n7358), .A2(n7100), .ZN(n7357) );
  AOI21_X1 U5996 ( .B1(n7376), .B2(n5074), .A(n5439), .ZN(n7718) );
  INV_X1 U5997 ( .A(n5440), .ZN(n5439) );
  AOI21_X1 U5998 ( .B1(n5441), .B2(n7587), .A(n7586), .ZN(n5440) );
  AND4_X1 U5999 ( .A1(n7795), .A2(n7794), .A3(n7793), .A4(n7792), .ZN(n8928)
         );
  NAND2_X1 U6000 ( .A1(n8913), .A2(n8532), .ZN(n8912) );
  INV_X1 U6001 ( .A(n8953), .ZN(n8915) );
  AND2_X1 U6002 ( .A1(n6581), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8935) );
  AND4_X1 U6003 ( .A1(n6563), .A2(n6562), .A3(n6561), .A4(n6560), .ZN(n7192)
         );
  AND2_X1 U6004 ( .A1(n7376), .A2(n7375), .ZN(n7491) );
  AND2_X1 U6005 ( .A1(n10823), .A2(n6592), .ZN(n8963) );
  OAI21_X1 U6006 ( .B1(n8397), .B2(n8396), .A(n8607), .ZN(n8972) );
  INV_X1 U6007 ( .A(n8935), .ZN(n8968) );
  INV_X1 U6008 ( .A(n8963), .ZN(n8975) );
  NAND2_X1 U6009 ( .A1(n8797), .A2(n8807), .ZN(n8803) );
  AOI21_X1 U6010 ( .B1(n8798), .B2(n8801), .A(n5508), .ZN(n8797) );
  NAND2_X1 U6011 ( .A1(n8801), .A2(n8811), .ZN(n8819) );
  INV_X1 U6012 ( .A(n8620), .ZN(n8820) );
  OR2_X1 U6013 ( .A1(n6780), .A2(n6470), .ZN(n8999) );
  AOI21_X1 U6014 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n6788), .A(n6828), .ZN(
        n6785) );
  AOI21_X1 U6015 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n6809), .A(n6818), .ZN(
        n6807) );
  AOI21_X1 U6016 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n6946), .A(n6945), .ZN(
        n6947) );
  AND2_X1 U6017 ( .A1(n6966), .A2(n7045), .ZN(n9014) );
  OR2_X1 U6018 ( .A1(n6511), .A2(n6510), .ZN(n6513) );
  AND2_X1 U6019 ( .A1(n9098), .A2(n5330), .ZN(n5329) );
  NOR2_X1 U6020 ( .A1(n5331), .A2(n9321), .ZN(n5330) );
  NAND2_X1 U6021 ( .A1(n5531), .A2(n5533), .ZN(n8578) );
  NAND2_X1 U6022 ( .A1(n5532), .A2(n5536), .ZN(n5531) );
  INV_X1 U6023 ( .A(n9135), .ZN(n5532) );
  NAND2_X1 U6024 ( .A1(n5538), .A2(n5542), .ZN(n9102) );
  NAND2_X1 U6025 ( .A1(n8303), .A2(n8302), .ZN(n9133) );
  AND2_X1 U6026 ( .A1(n8273), .A2(n8272), .ZN(n9175) );
  NAND2_X1 U6027 ( .A1(n9214), .A2(n5645), .ZN(n9206) );
  NAND2_X1 U6028 ( .A1(n5186), .A2(n8713), .ZN(n9195) );
  NAND2_X1 U6029 ( .A1(n9211), .A2(n8788), .ZN(n5186) );
  INV_X1 U6030 ( .A(n9357), .ZN(n9221) );
  NAND2_X1 U6031 ( .A1(n8224), .A2(n8223), .ZN(n9369) );
  NAND2_X1 U6032 ( .A1(n8210), .A2(n8209), .ZN(n9379) );
  NAND2_X1 U6033 ( .A1(n5194), .A2(n8691), .ZN(n9284) );
  AND2_X1 U6034 ( .A1(n10998), .A2(n8063), .ZN(n8065) );
  NAND2_X1 U6035 ( .A1(n5476), .A2(n5475), .ZN(n7547) );
  INV_X1 U6036 ( .A(n10912), .ZN(n8648) );
  CLKBUF_X1 U6037 ( .A(n7461), .Z(n10916) );
  INV_X1 U6038 ( .A(n10819), .ZN(n9292) );
  NAND2_X1 U6039 ( .A1(n6589), .A2(n10702), .ZN(n10823) );
  AND2_X2 U6040 ( .A1(n7237), .A2(n7195), .ZN(n11002) );
  AND2_X2 U6041 ( .A1(n7237), .A2(n7236), .ZN(n11006) );
  AND2_X1 U6042 ( .A1(n6679), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10772) );
  NAND2_X1 U6043 ( .A1(n5235), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6515) );
  INV_X1 U6044 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8261) );
  XNOR2_X1 U6045 ( .A(n6496), .B(n6495), .ZN(n8620) );
  INV_X1 U6046 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8246) );
  CLKBUF_X1 U6047 ( .A(n6579), .Z(n8801) );
  INV_X1 U6048 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8495) );
  INV_X1 U6049 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7054) );
  INV_X1 U6050 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6958) );
  INV_X1 U6051 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6906) );
  INV_X1 U6052 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6698) );
  NOR2_X1 U6053 ( .A1(n6471), .A2(n6444), .ZN(n6648) );
  NAND2_X1 U6054 ( .A1(n5159), .A2(n5158), .ZN(n9467) );
  NAND2_X1 U6055 ( .A1(n5159), .A2(n5160), .ZN(n9464) );
  NOR2_X1 U6056 ( .A1(n5602), .A2(n5122), .ZN(n8104) );
  AND4_X1 U6057 ( .A1(n5903), .A2(n5902), .A3(n5901), .A4(n5900), .ZN(n7572)
         );
  AOI21_X1 U6058 ( .B1(n9483), .B2(n9494), .A(n9493), .ZN(n9496) );
  AND2_X1 U6059 ( .A1(n6299), .A2(n6298), .ZN(n9508) );
  OR2_X1 U6060 ( .A1(n6436), .A2(n9830), .ZN(n9559) );
  NAND2_X1 U6061 ( .A1(n5164), .A2(n9446), .ZN(n9515) );
  NAND2_X1 U6062 ( .A1(n5166), .A2(n5165), .ZN(n5164) );
  INV_X1 U6063 ( .A(n9449), .ZN(n5166) );
  AOI21_X1 U6064 ( .B1(n7946), .B2(n5148), .A(n5147), .ZN(n5145) );
  NAND2_X1 U6065 ( .A1(n5602), .A2(n5154), .ZN(n5146) );
  NOR2_X1 U6066 ( .A1(n8101), .A2(n8100), .ZN(n5147) );
  AND2_X1 U6067 ( .A1(n6248), .A2(n6247), .ZN(n10038) );
  INV_X1 U6068 ( .A(n5605), .ZN(n8014) );
  AOI21_X1 U6069 ( .B1(n5178), .B2(n6343), .A(n5588), .ZN(n5177) );
  NAND2_X1 U6070 ( .A1(n6343), .A2(n5181), .ZN(n5179) );
  NOR2_X1 U6071 ( .A1(n9504), .A2(n5180), .ZN(n5178) );
  NAND2_X1 U6072 ( .A1(n6352), .A2(n6351), .ZN(n10168) );
  INV_X1 U6073 ( .A(n9535), .ZN(n9566) );
  INV_X1 U6074 ( .A(n9508), .ZN(n10015) );
  INV_X1 U6075 ( .A(n10038), .ZN(n10016) );
  OR2_X1 U6076 ( .A1(n6159), .A2(n6158), .ZN(n10129) );
  INV_X1 U6077 ( .A(n7564), .ZN(n7648) );
  INV_X1 U6078 ( .A(n7572), .ZN(n9848) );
  AND3_X1 U6079 ( .A1(n5091), .A2(n5859), .A3(n5858), .ZN(n5861) );
  OR2_X1 U6080 ( .A1(n5806), .A2(n5833), .ZN(n5836) );
  CLKBUF_X1 U6081 ( .A(n7241), .Z(n9851) );
  NAND2_X1 U6082 ( .A1(n5855), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5770) );
  OR2_X1 U6083 ( .A1(n5806), .A2(n5767), .ZN(n5771) );
  INV_X1 U6084 ( .A(n10659), .ZN(n10030) );
  AND2_X1 U6085 ( .A1(n9576), .A2(n9575), .ZN(n11019) );
  NAND2_X1 U6086 ( .A1(n8455), .A2(n8454), .ZN(n10152) );
  INV_X1 U6087 ( .A(n5391), .ZN(n5390) );
  NAND2_X1 U6088 ( .A1(n8466), .A2(n8465), .ZN(n8467) );
  AOI21_X1 U6089 ( .B1(n9916), .B2(n10125), .A(n9915), .ZN(n10161) );
  NAND2_X1 U6090 ( .A1(n9914), .A2(n9913), .ZN(n9915) );
  NAND2_X1 U6091 ( .A1(n5140), .A2(n5138), .ZN(n10173) );
  AOI21_X1 U6092 ( .B1(n9940), .B2(n10130), .A(n5139), .ZN(n5138) );
  NOR2_X1 U6093 ( .A1(n9974), .A2(n10081), .ZN(n5139) );
  NAND2_X1 U6094 ( .A1(n5415), .A2(n5414), .ZN(n9958) );
  AND2_X1 U6095 ( .A1(n5415), .A2(n5106), .ZN(n9959) );
  NAND2_X1 U6096 ( .A1(n6305), .A2(n6304), .ZN(n10179) );
  AND2_X1 U6097 ( .A1(n6291), .A2(n6290), .ZN(n9998) );
  NAND2_X1 U6098 ( .A1(n10041), .A2(n8475), .ZN(n10021) );
  INV_X1 U6099 ( .A(n10198), .ZN(n10054) );
  NAND2_X1 U6100 ( .A1(n10080), .A2(n9713), .ZN(n10066) );
  NAND2_X1 U6101 ( .A1(n8174), .A2(n8173), .ZN(n8176) );
  NAND2_X1 U6102 ( .A1(n6097), .A2(n6096), .ZN(n9567) );
  NAND2_X1 U6103 ( .A1(n5619), .A2(n5621), .ZN(n8178) );
  NAND2_X1 U6104 ( .A1(n7961), .A2(n7960), .ZN(n7963) );
  NAND2_X1 U6105 ( .A1(n5636), .A2(n9674), .ZN(n7955) );
  NAND2_X1 U6106 ( .A1(n5410), .A2(n7817), .ZN(n7819) );
  AND2_X1 U6107 ( .A1(n5628), .A2(n9660), .ZN(n7563) );
  AND2_X1 U6108 ( .A1(n5926), .A2(n5925), .ZN(n7608) );
  INV_X1 U6109 ( .A(n10903), .ZN(n7571) );
  NAND2_X1 U6110 ( .A1(n5838), .A2(n5813), .ZN(n5822) );
  OR2_X1 U6111 ( .A1(n5842), .A2(n5819), .ZN(n5820) );
  INV_X1 U6112 ( .A(n10095), .ZN(n10144) );
  OAI21_X1 U6113 ( .B1(n6473), .B2(n5775), .A(n5774), .ZN(n7296) );
  NAND2_X1 U6114 ( .A1(n6473), .A2(n10664), .ZN(n5774) );
  AND2_X1 U6115 ( .A1(n10093), .A2(n7078), .ZN(n10115) );
  INV_X1 U6116 ( .A(n11024), .ZN(n11023) );
  OAI21_X1 U6117 ( .B1(n10150), .B2(n11009), .A(n5299), .ZN(n10240) );
  NOR2_X1 U6118 ( .A1(n5070), .A2(n5300), .ZN(n5299) );
  INV_X1 U6119 ( .A(n11017), .ZN(n5300) );
  AND2_X1 U6120 ( .A1(n6471), .A2(n6392), .ZN(n10257) );
  NAND2_X1 U6121 ( .A1(n8609), .A2(n8608), .ZN(n8612) );
  XNOR2_X1 U6122 ( .A(n8193), .B(n8189), .ZN(n8315) );
  NAND2_X1 U6123 ( .A1(n6368), .A2(n6367), .ZN(n8193) );
  INV_X1 U6124 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10445) );
  INV_X1 U6125 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10443) );
  INV_X1 U6126 ( .A(n5726), .ZN(n5727) );
  INV_X1 U6127 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10555) );
  NAND2_X1 U6128 ( .A1(n5733), .A2(n5732), .ZN(n7976) );
  INV_X1 U6129 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7709) );
  NAND2_X1 U6130 ( .A1(n5758), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5759) );
  OR2_X1 U6131 ( .A1(n5737), .A2(n10628), .ZN(n5738) );
  INV_X1 U6132 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10562) );
  INV_X1 U6133 ( .A(n9798), .ZN(n9823) );
  XNOR2_X1 U6134 ( .A(n10668), .B(n5264), .ZN(n5263) );
  INV_X1 U6135 ( .A(keyinput_126), .ZN(n5264) );
  INV_X1 U6136 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10569) );
  INV_X1 U6137 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10574) );
  INV_X1 U6138 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10442) );
  INV_X1 U6139 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10272) );
  INV_X1 U6140 ( .A(n8999), .ZN(P2_U3966) );
  OAI21_X1 U6141 ( .B1(n9314), .B2(n9303), .A(n5087), .ZN(P2_U3267) );
  OR2_X1 U6142 ( .A1(n9315), .A2(n9300), .ZN(n5240) );
  AOI21_X1 U6143 ( .B1(n9312), .B2(n9226), .A(n8378), .ZN(n5241) );
  INV_X1 U6144 ( .A(n5296), .ZN(P1_U3554) );
  AOI21_X1 U6145 ( .B1(n10240), .B2(n11024), .A(n5297), .ZN(n5296) );
  NOR2_X1 U6146 ( .A1(n11024), .A2(n5298), .ZN(n5297) );
  INV_X1 U6147 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n5298) );
  AOI21_X1 U6148 ( .B1(n5265), .B2(n5262), .A(n10656), .ZN(n10663) );
  AND2_X1 U6149 ( .A1(n10657), .A2(n5263), .ZN(n5262) );
  AND2_X1 U6150 ( .A1(n5533), .A2(n8586), .ZN(n5041) );
  NAND2_X1 U6151 ( .A1(n5320), .A2(n5319), .ZN(n5042) );
  INV_X1 U6152 ( .A(n8791), .ZN(n5229) );
  AND2_X1 U6153 ( .A1(n5486), .A2(n5066), .ZN(n5043) );
  INV_X4 U6154 ( .A(n5656), .ZN(n5668) );
  AND2_X1 U6155 ( .A1(n5425), .A2(n8035), .ZN(n5044) );
  INV_X1 U6156 ( .A(n9229), .ZN(n5465) );
  AND3_X1 U6157 ( .A1(n5870), .A2(n5869), .A3(n5868), .ZN(n7411) );
  NOR2_X1 U6158 ( .A1(n5543), .A2(n5537), .ZN(n5536) );
  AND2_X1 U6159 ( .A1(n10073), .A2(n9708), .ZN(n5045) );
  AND2_X1 U6160 ( .A1(n7118), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5046) );
  NAND2_X1 U6161 ( .A1(n6388), .A2(n5606), .ZN(n5047) );
  AND2_X1 U6162 ( .A1(n9986), .A2(n5307), .ZN(n5048) );
  AND2_X1 U6163 ( .A1(n5065), .A2(n10054), .ZN(n5049) );
  INV_X1 U6164 ( .A(n9652), .ZN(n5624) );
  INV_X1 U6165 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7051) );
  INV_X1 U6166 ( .A(n9447), .ZN(n5165) );
  AND2_X1 U6167 ( .A1(n5618), .A2(n9683), .ZN(n5050) );
  AND2_X1 U6168 ( .A1(n9189), .A2(n8722), .ZN(n5051) );
  AOI21_X1 U6169 ( .B1(n6173), .B2(n6172), .A(n5113), .ZN(n5483) );
  AND2_X1 U6170 ( .A1(n9919), .A2(n5397), .ZN(n5052) );
  NOR2_X1 U6171 ( .A1(n8534), .A2(n8533), .ZN(n5053) );
  AND3_X1 U6172 ( .A1(n6021), .A2(n10608), .A3(n6070), .ZN(n5054) );
  NOR2_X1 U6173 ( .A1(n9316), .A2(n8979), .ZN(n5055) );
  INV_X1 U6174 ( .A(n6280), .ZN(n5593) );
  AND2_X1 U6175 ( .A1(n7962), .A2(n7960), .ZN(n5057) );
  INV_X1 U6176 ( .A(n10163), .ZN(n5394) );
  AND2_X1 U6177 ( .A1(n9609), .A2(n7598), .ZN(n7558) );
  INV_X1 U6178 ( .A(n6344), .ZN(n5588) );
  NAND2_X1 U6179 ( .A1(n7998), .A2(n5461), .ZN(n5460) );
  INV_X1 U6180 ( .A(n9369), .ZN(n5320) );
  INV_X1 U6181 ( .A(n6063), .ZN(n5153) );
  AND3_X1 U6182 ( .A1(n10379), .A2(n10378), .A3(n5131), .ZN(n5058) );
  XOR2_X1 U6183 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_222), .Z(n5059) );
  NAND2_X1 U6184 ( .A1(n10194), .A2(n10016), .ZN(n5060) );
  NAND2_X1 U6185 ( .A1(n5861), .A2(n5860), .ZN(n5875) );
  XNOR2_X1 U6186 ( .A(n5759), .B(n10630), .ZN(n5765) );
  XNOR2_X1 U6187 ( .A(n6515), .B(n9416), .ZN(n6520) );
  OR2_X1 U6188 ( .A1(n9352), .A2(n9213), .ZN(n5061) );
  AND2_X1 U6189 ( .A1(n8706), .A2(n8705), .ZN(n9249) );
  INV_X1 U6190 ( .A(n9249), .ZN(n5469) );
  INV_X1 U6191 ( .A(n5162), .ZN(n5161) );
  OR2_X1 U6192 ( .A1(n6233), .A2(n5163), .ZN(n5162) );
  OAI211_X1 U6193 ( .C1(n7537), .C2(n6837), .A(n6567), .B(n6566), .ZN(n7315)
         );
  INV_X1 U6194 ( .A(n9470), .ZN(n10025) );
  NOR2_X1 U6195 ( .A1(n8516), .A2(n8850), .ZN(n5062) );
  AND2_X1 U6196 ( .A1(n10877), .A2(n10864), .ZN(n5063) );
  AND2_X1 U6197 ( .A1(n5484), .A2(n5204), .ZN(n5064) );
  NAND2_X1 U6198 ( .A1(n8237), .A2(n8236), .ZN(n9361) );
  NAND2_X1 U6199 ( .A1(n8496), .A2(n10269), .ZN(n5806) );
  NAND2_X1 U6200 ( .A1(n9522), .A2(n6280), .ZN(n9437) );
  AND2_X1 U6201 ( .A1(n10064), .A2(n10208), .ZN(n5065) );
  XOR2_X1 U6202 ( .A(n6014), .B(SI_11_), .Z(n5066) );
  AND3_X1 U6203 ( .A1(n5705), .A2(n6021), .A3(n10630), .ZN(n5067) );
  NOR2_X1 U6204 ( .A1(n8160), .A2(n8161), .ZN(n5459) );
  AND2_X1 U6205 ( .A1(n6791), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5068) );
  NAND2_X1 U6206 ( .A1(n5173), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5739) );
  AND2_X1 U6207 ( .A1(n8993), .A2(n10931), .ZN(n5069) );
  AND2_X1 U6208 ( .A1(n10149), .A2(n10946), .ZN(n5070) );
  INV_X1 U6209 ( .A(n8416), .ZN(n6300) );
  INV_X1 U6210 ( .A(n8013), .ZN(n5604) );
  OR2_X1 U6211 ( .A1(n8729), .A2(n8760), .ZN(n5071) );
  NAND2_X1 U6212 ( .A1(n8474), .A2(n5641), .ZN(n10041) );
  AND3_X1 U6213 ( .A1(n5067), .A2(n5608), .A3(n5056), .ZN(n5072) );
  NAND2_X2 U6214 ( .A1(n6579), .A2(n5446), .ZN(n8535) );
  AND2_X1 U6215 ( .A1(n5481), .A2(n5478), .ZN(n5073) );
  AND2_X1 U6216 ( .A1(n8713), .A2(n8712), .ZN(n8788) );
  INV_X1 U6217 ( .A(n8788), .ZN(n9215) );
  NAND2_X1 U6218 ( .A1(n5528), .A2(n8232), .ZN(n9228) );
  NAND2_X1 U6219 ( .A1(n6454), .A2(n6499), .ZN(n6497) );
  AND2_X1 U6220 ( .A1(n7587), .A2(n7375), .ZN(n5074) );
  NAND2_X1 U6221 ( .A1(n6370), .A2(n6369), .ZN(n10163) );
  INV_X1 U6222 ( .A(n8742), .ZN(n5540) );
  INV_X1 U6223 ( .A(n5543), .ZN(n5542) );
  OAI22_X1 U6224 ( .A1(n9119), .A2(n5547), .B1(n8981), .B2(n9133), .ZN(n5543)
         );
  AND2_X1 U6225 ( .A1(n8749), .A2(n8746), .ZN(n8793) );
  NAND2_X1 U6226 ( .A1(n6330), .A2(n6329), .ZN(n10175) );
  NOR2_X1 U6227 ( .A1(n9383), .A2(n8986), .ZN(n5075) );
  NOR2_X1 U6228 ( .A1(n9439), .A2(n9438), .ZN(n5076) );
  INV_X1 U6229 ( .A(n9547), .ZN(n9953) );
  AND4_X1 U6230 ( .A1(n6377), .A2(n6376), .A3(n6375), .A4(n6374), .ZN(n9547)
         );
  AND2_X1 U6231 ( .A1(n8161), .A2(n8063), .ZN(n5077) );
  NAND2_X1 U6232 ( .A1(n9986), .A2(n5309), .ZN(n5310) );
  AND2_X1 U6233 ( .A1(n5632), .A2(n7817), .ZN(n5078) );
  XNOR2_X1 U6234 ( .A(n8998), .B(n10864), .ZN(n7209) );
  AND2_X1 U6235 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5079) );
  INV_X1 U6236 ( .A(n9321), .ZN(n9106) );
  NAND2_X1 U6237 ( .A1(n8318), .A2(n8317), .ZN(n9321) );
  AND2_X1 U6238 ( .A1(n5566), .A2(n5564), .ZN(n5080) );
  AND2_X1 U6239 ( .A1(n9660), .A2(n9772), .ZN(n5081) );
  AND2_X1 U6240 ( .A1(n9214), .A2(n5555), .ZN(n5082) );
  AND2_X1 U6241 ( .A1(n10041), .A2(n5408), .ZN(n5083) );
  OR2_X1 U6242 ( .A1(n6208), .A2(n5155), .ZN(n5084) );
  AND2_X1 U6243 ( .A1(n6013), .A2(n6012), .ZN(n5085) );
  INV_X1 U6244 ( .A(n8101), .ZN(n5154) );
  NAND2_X1 U6245 ( .A1(n8415), .A2(n8414), .ZN(n10158) );
  NOR2_X1 U6246 ( .A1(n10175), .A2(n9982), .ZN(n5086) );
  AND2_X1 U6247 ( .A1(n5241), .A2(n5240), .ZN(n5087) );
  AND4_X1 U6248 ( .A1(n6452), .A2(n6500), .A3(n6692), .A4(n6960), .ZN(n5088)
         );
  INV_X1 U6249 ( .A(n9136), .ZN(n9142) );
  AND2_X1 U6250 ( .A1(n9118), .A2(n8732), .ZN(n9136) );
  AND2_X1 U6251 ( .A1(n7167), .A2(n7166), .ZN(n5089) );
  INV_X1 U6252 ( .A(n5547), .ZN(n5545) );
  NAND2_X1 U6253 ( .A1(n9140), .A2(n9158), .ZN(n5547) );
  INV_X1 U6254 ( .A(n9773), .ZN(n5632) );
  NOR2_X1 U6255 ( .A1(n9513), .A2(n9512), .ZN(n5090) );
  OR2_X1 U6256 ( .A1(n5854), .A2(n6605), .ZN(n5091) );
  AND2_X1 U6257 ( .A1(n6014), .A2(SI_11_), .ZN(n5092) );
  AND2_X1 U6258 ( .A1(n6085), .A2(SI_14_), .ZN(n5093) );
  INV_X1 U6259 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5326) );
  AND2_X1 U6260 ( .A1(n9685), .A2(n9683), .ZN(n9778) );
  INV_X1 U6261 ( .A(n9778), .ZN(n5618) );
  NAND2_X1 U6262 ( .A1(n5565), .A2(n5080), .ZN(n5570) );
  INV_X1 U6263 ( .A(n5615), .ZN(n5619) );
  NAND2_X1 U6264 ( .A1(n5620), .A2(n9683), .ZN(n5615) );
  INV_X1 U6265 ( .A(n5626), .ZN(n5625) );
  NAND2_X1 U6266 ( .A1(n9944), .A2(n5627), .ZN(n5626) );
  OAI21_X1 U6267 ( .B1(n5451), .B2(n5448), .A(n8810), .ZN(n5447) );
  AND2_X1 U6268 ( .A1(n9712), .A2(n9713), .ZN(n10073) );
  OR2_X1 U6269 ( .A1(n9439), .A2(n5593), .ZN(n5094) );
  INV_X1 U6270 ( .A(n5536), .ZN(n5535) );
  INV_X1 U6271 ( .A(n9361), .ZN(n9236) );
  INV_X1 U6272 ( .A(n8809), .ZN(n5451) );
  AND2_X1 U6273 ( .A1(n8618), .A2(n8755), .ZN(n8809) );
  OR2_X1 U6274 ( .A1(n5451), .A2(n9307), .ZN(n5095) );
  NAND2_X1 U6275 ( .A1(n9654), .A2(n9653), .ZN(n9970) );
  NAND2_X1 U6276 ( .A1(n9754), .A2(n9756), .ZN(n9790) );
  INV_X1 U6277 ( .A(n9790), .ZN(n5400) );
  OR2_X1 U6278 ( .A1(n9357), .A2(n9233), .ZN(n8713) );
  INV_X1 U6279 ( .A(n7424), .ZN(n5578) );
  AND2_X1 U6280 ( .A1(n8810), .A2(n8756), .ZN(n5096) );
  AND2_X1 U6281 ( .A1(n5307), .A2(n9920), .ZN(n5097) );
  NOR2_X1 U6282 ( .A1(n10480), .A2(n5332), .ZN(n5098) );
  AND2_X1 U6283 ( .A1(n5465), .A2(n8232), .ZN(n5099) );
  AND2_X1 U6284 ( .A1(n8544), .A2(n5445), .ZN(n5100) );
  AND2_X1 U6285 ( .A1(n8660), .A2(n7548), .ZN(n5101) );
  OR2_X1 U6286 ( .A1(n7537), .A2(n10791), .ZN(n5102) );
  AND2_X1 U6287 ( .A1(n9215), .A2(n5557), .ZN(n5103) );
  AND2_X1 U6288 ( .A1(n5060), .A2(n5641), .ZN(n5104) );
  AND2_X1 U6289 ( .A1(n5206), .A2(n8622), .ZN(n5105) );
  NAND2_X1 U6290 ( .A1(n10179), .A2(n10002), .ZN(n5106) );
  AND2_X1 U6291 ( .A1(n5064), .A2(n5202), .ZN(n5107) );
  AND2_X1 U6292 ( .A1(n8175), .A2(n8173), .ZN(n5108) );
  INV_X1 U6293 ( .A(n5193), .ZN(n5192) );
  NOR2_X1 U6294 ( .A1(n8361), .A2(n8693), .ZN(n5193) );
  AND2_X1 U6295 ( .A1(n8690), .A2(n8785), .ZN(n5109) );
  AND2_X1 U6296 ( .A1(n8728), .A2(n5071), .ZN(n5110) );
  INV_X1 U6297 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n10633) );
  INV_X2 U6298 ( .A(n5854), .ZN(n5768) );
  AND2_X1 U6299 ( .A1(n5424), .A2(n5425), .ZN(n5111) );
  INV_X1 U6300 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5137) );
  OR2_X1 U6301 ( .A1(n9296), .A2(n9375), .ZN(n5112) );
  XOR2_X1 U6302 ( .A(n6191), .B(SI_18_), .Z(n5113) );
  NAND2_X1 U6303 ( .A1(n5151), .A2(n5149), .ZN(n9425) );
  AND2_X1 U6304 ( .A1(n5455), .A2(n5456), .ZN(n5114) );
  AND3_X1 U6305 ( .A1(n5403), .A2(n5306), .A3(n5054), .ZN(n6090) );
  AND2_X1 U6306 ( .A1(n6254), .A2(n6253), .ZN(n5115) );
  INV_X1 U6307 ( .A(n8859), .ZN(n5417) );
  AND2_X1 U6308 ( .A1(n6364), .A2(n6363), .ZN(n5116) );
  NAND2_X1 U6309 ( .A1(n5403), .A2(n5306), .ZN(n6019) );
  INV_X1 U6310 ( .A(n5181), .ZN(n5180) );
  AND2_X1 U6311 ( .A1(n6268), .A2(n6267), .ZN(n10012) );
  INV_X1 U6312 ( .A(n10012), .ZN(n10188) );
  INV_X1 U6313 ( .A(n5502), .ZN(n5501) );
  NAND2_X1 U6314 ( .A1(n5505), .A2(n5506), .ZN(n5502) );
  AND2_X1 U6315 ( .A1(n6192), .A2(SI_18_), .ZN(n5117) );
  NOR2_X1 U6316 ( .A1(n9296), .A2(n5042), .ZN(n5118) );
  NAND2_X1 U6317 ( .A1(n7332), .A2(n8640), .ZN(n7443) );
  XNOR2_X1 U6318 ( .A(n5725), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6395) );
  NAND2_X1 U6319 ( .A1(n7674), .A2(n7673), .ZN(n7644) );
  OR2_X1 U6320 ( .A1(n7491), .A2(n5441), .ZN(n7588) );
  XNOR2_X1 U6321 ( .A(n6509), .B(n6508), .ZN(n6579) );
  NAND2_X1 U6322 ( .A1(n7262), .A2(n9760), .ZN(n6387) );
  NAND2_X1 U6323 ( .A1(n8215), .A2(n8214), .ZN(n9375) );
  INV_X1 U6324 ( .A(n9375), .ZN(n5319) );
  NAND2_X1 U6325 ( .A1(n5170), .A2(n5598), .ZN(n7165) );
  AND2_X1 U6326 ( .A1(n5601), .A2(n5600), .ZN(n7061) );
  AND2_X1 U6327 ( .A1(n9684), .A2(n9686), .ZN(n9777) );
  INV_X1 U6328 ( .A(n9446), .ZN(n5163) );
  OAI21_X1 U6329 ( .B1(n7206), .B2(n7209), .A(n7188), .ZN(n8632) );
  NAND2_X1 U6330 ( .A1(n6239), .A2(n6238), .ZN(n10194) );
  INV_X1 U6331 ( .A(n10194), .ZN(n5314) );
  XNOR2_X1 U6332 ( .A(n8573), .B(keyinput_170), .ZN(n5119) );
  XNOR2_X1 U6333 ( .A(n10527), .B(keyinput_39), .ZN(n5120) );
  NAND2_X1 U6334 ( .A1(n8072), .A2(n8032), .ZN(n5121) );
  AND2_X1 U6335 ( .A1(n7946), .A2(n5604), .ZN(n5122) );
  XOR2_X1 U6336 ( .A(SI_9_), .B(keyinput_23), .Z(n5123) );
  NAND2_X1 U6337 ( .A1(n7764), .A2(n7763), .ZN(n5124) );
  INV_X1 U6338 ( .A(n5312), .ZN(n7669) );
  NOR2_X1 U6339 ( .A1(n7604), .A2(n10921), .ZN(n5312) );
  NAND2_X1 U6340 ( .A1(n5571), .A2(n5576), .ZN(n7643) );
  INV_X1 U6341 ( .A(n5324), .ZN(n7880) );
  NOR2_X1 U6342 ( .A1(n7771), .A2(n7856), .ZN(n5324) );
  AND2_X1 U6343 ( .A1(n5605), .A2(n5604), .ZN(n5125) );
  AND2_X1 U6344 ( .A1(n5476), .A2(n7446), .ZN(n5126) );
  AND2_X1 U6345 ( .A1(SI_22_), .A2(keyinput_10), .ZN(n5127) );
  AND2_X1 U6346 ( .A1(SI_2_), .A2(keyinput_30), .ZN(n5128) );
  OR2_X1 U6347 ( .A1(n6464), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n5129) );
  INV_X1 U6348 ( .A(n5474), .ZN(n5475) );
  NAND2_X1 U6349 ( .A1(n5763), .A2(n6387), .ZN(n7255) );
  INV_X1 U6350 ( .A(n7679), .ZN(n5311) );
  NAND2_X2 U6351 ( .A1(n8233), .A2(n8621), .ZN(n8752) );
  INV_X1 U6352 ( .A(n10125), .ZN(n9972) );
  OR2_X1 U6353 ( .A1(n9830), .A2(n6387), .ZN(n10083) );
  INV_X1 U6354 ( .A(n10083), .ZN(n10130) );
  INV_X1 U6355 ( .A(n7411), .ZN(n5871) );
  NAND2_X1 U6356 ( .A1(n5776), .A2(n5084), .ZN(n6935) );
  INV_X1 U6357 ( .A(SI_28_), .ZN(n10479) );
  INV_X1 U6358 ( .A(SI_30_), .ZN(n5272) );
  XOR2_X1 U6359 ( .A(n10592), .B(keyinput_223), .Z(n5130) );
  XOR2_X1 U6360 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .Z(n5131) );
  XNOR2_X1 U6361 ( .A(n6498), .B(n5326), .ZN(n8807) );
  XNOR2_X1 U6362 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_115), .ZN(n5132) );
  AND2_X1 U6363 ( .A1(n10392), .A2(n10391), .ZN(n5133) );
  INV_X1 U6364 ( .A(n5747), .ZN(n8496) );
  INV_X2 U6365 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n10628) );
  AND2_X1 U6366 ( .A1(n10436), .A2(n10437), .ZN(n5134) );
  INV_X1 U6367 ( .A(n10257), .ZN(n10666) );
  NAND2_X1 U6368 ( .A1(n7781), .A2(n8616), .ZN(n5135) );
  NAND2_X1 U6369 ( .A1(n7632), .A2(n7548), .ZN(n7631) );
  NAND2_X1 U6370 ( .A1(n6529), .A2(n6530), .ZN(n6516) );
  INV_X1 U6371 ( .A(n8924), .ZN(n5427) );
  INV_X1 U6372 ( .A(n9186), .ZN(n8367) );
  INV_X1 U6373 ( .A(n6174), .ZN(n5480) );
  NAND2_X1 U6374 ( .A1(n6288), .A2(n6287), .ZN(n6303) );
  NAND2_X1 U6375 ( .A1(n8501), .A2(n8345), .ZN(n10268) );
  NAND2_X1 U6376 ( .A1(n5203), .A2(n5107), .ZN(n6045) );
  NAND2_X1 U6377 ( .A1(n8479), .A2(n8478), .ZN(n9978) );
  OAI22_X2 U6378 ( .A1(n9945), .A2(n8480), .B1(n9973), .B2(n9950), .ZN(n9931)
         );
  NAND2_X1 U6379 ( .A1(n5407), .A2(n5405), .ZN(n10008) );
  NAND2_X1 U6380 ( .A1(n10008), .A2(n5143), .ZN(n8477) );
  NAND2_X1 U6381 ( .A1(n5214), .A2(n8793), .ZN(n5213) );
  NAND2_X1 U6382 ( .A1(n5226), .A2(n5101), .ZN(n5225) );
  NAND2_X1 U6383 ( .A1(n5217), .A2(n5109), .ZN(n8696) );
  AOI21_X1 U6384 ( .B1(n5210), .B2(n8751), .A(n5209), .ZN(n8754) );
  NAND2_X1 U6385 ( .A1(n8676), .A2(n8752), .ZN(n5221) );
  OAI21_X1 U6386 ( .B1(n5230), .B2(n5228), .A(n5110), .ZN(n8735) );
  NAND3_X1 U6387 ( .A1(n5328), .A2(n5102), .A3(n5327), .ZN(n7400) );
  OR2_X2 U6388 ( .A1(n6529), .A2(n7051), .ZN(n6531) );
  AND2_X2 U6389 ( .A1(n6459), .A2(n5559), .ZN(n6529) );
  NAND2_X1 U6390 ( .A1(n8655), .A2(n8654), .ZN(n5227) );
  OAI22_X1 U6391 ( .A1(n8720), .A2(n9194), .B1(n8760), .B2(n8719), .ZN(n5231)
         );
  NAND2_X2 U6392 ( .A1(n5686), .A2(n5685), .ZN(n5966) );
  OAI21_X2 U6393 ( .B1(n8116), .B2(n5615), .A(n5616), .ZN(n8179) );
  AND2_X1 U6394 ( .A1(n9971), .A2(n9970), .ZN(n5141) );
  NAND2_X1 U6395 ( .A1(n5812), .A2(n5811), .ZN(n5142) );
  NAND2_X1 U6396 ( .A1(n7502), .A2(n7501), .ZN(n7506) );
  NAND2_X1 U6397 ( .A1(n10076), .A2(n5642), .ZN(n10039) );
  NOR2_X1 U6398 ( .A1(n9918), .A2(n9919), .ZN(n9917) );
  NOR2_X1 U6399 ( .A1(n9171), .A2(n5229), .ZN(n9170) );
  NAND2_X2 U6400 ( .A1(n9151), .A2(n8289), .ZN(n9135) );
  XNOR2_X2 U6401 ( .A(n5988), .B(n5648), .ZN(n7748) );
  AOI211_X2 U6402 ( .C1(n9125), .C2(n10980), .A(n9124), .B(n9123), .ZN(n9327)
         );
  OAI22_X2 U6403 ( .A1(n9261), .A2(n8764), .B1(n9253), .B2(n9375), .ZN(n9247)
         );
  NOR2_X1 U6404 ( .A1(n10803), .A2(n10804), .ZN(n10802) );
  NAND2_X1 U6405 ( .A1(n5146), .A2(n5145), .ZN(n8138) );
  OAI21_X2 U6406 ( .B1(n9449), .B2(n5157), .A(n5156), .ZN(n9523) );
  NAND2_X1 U6407 ( .A1(n5170), .A2(n5168), .ZN(n5919) );
  NAND2_X1 U6408 ( .A1(n5736), .A2(n5174), .ZN(n5172) );
  NAND2_X1 U6409 ( .A1(n5736), .A2(n5176), .ZN(n5173) );
  NAND4_X1 U6410 ( .A1(n5403), .A2(n5306), .A3(n5054), .A4(n5735), .ZN(n6093)
         );
  AOI21_X1 U6411 ( .B1(n9503), .B2(n9504), .A(n5180), .ZN(n9477) );
  OAI21_X1 U6412 ( .B1(n9503), .B2(n5179), .A(n5177), .ZN(n9544) );
  NAND2_X1 U6413 ( .A1(n6319), .A2(n6318), .ZN(n5181) );
  OAI21_X1 U6414 ( .B1(n9211), .B2(n5184), .A(n5182), .ZN(n9186) );
  NAND2_X1 U6415 ( .A1(n5454), .A2(n5193), .ZN(n5191) );
  NAND3_X1 U6416 ( .A1(n5191), .A2(n5189), .A3(n8698), .ZN(n9262) );
  NAND2_X1 U6417 ( .A1(n5459), .A2(n5453), .ZN(n5455) );
  NAND2_X1 U6418 ( .A1(n5195), .A2(n5455), .ZN(n5194) );
  NAND2_X1 U6419 ( .A1(n8805), .A2(n5198), .ZN(n5197) );
  NAND2_X1 U6420 ( .A1(n5966), .A2(n5043), .ZN(n5203) );
  NAND2_X1 U6421 ( .A1(n9189), .A2(n5207), .ZN(n5206) );
  NAND2_X1 U6422 ( .A1(n5215), .A2(n8801), .ZN(n8802) );
  NAND2_X1 U6423 ( .A1(n8758), .A2(n8759), .ZN(n5216) );
  NAND3_X1 U6424 ( .A1(n5220), .A2(n8683), .A3(n8682), .ZN(n5219) );
  NAND3_X1 U6425 ( .A1(n5222), .A2(n5221), .A3(n7800), .ZN(n5220) );
  NAND2_X1 U6426 ( .A1(n6459), .A2(n5232), .ZN(n5235) );
  INV_X1 U6427 ( .A(n7199), .ZN(n7185) );
  NAND3_X1 U6428 ( .A1(n6542), .A2(n5236), .A3(n6541), .ZN(n7199) );
  AND3_X2 U6429 ( .A1(n6499), .A2(n5326), .A3(n6454), .ZN(n6459) );
  AND2_X2 U6430 ( .A1(n5031), .A2(n5088), .ZN(n6454) );
  NAND4_X1 U6431 ( .A1(n5271), .A2(n5269), .A3(n5267), .A4(n5266), .ZN(n10317)
         );
  AND2_X1 U6432 ( .A1(n5305), .A2(n5306), .ZN(n5303) );
  AND2_X2 U6433 ( .A1(n5072), .A2(n5303), .ZN(n5722) );
  INV_X1 U6434 ( .A(n5702), .ZN(n5306) );
  INV_X1 U6435 ( .A(n5713), .ZN(n5403) );
  NAND2_X1 U6436 ( .A1(n9986), .A2(n5097), .ZN(n9921) );
  INV_X1 U6437 ( .A(n5310), .ZN(n9946) );
  NAND2_X1 U6438 ( .A1(n10114), .A2(n5313), .ZN(n10027) );
  INV_X1 U6439 ( .A(n9296), .ZN(n5315) );
  NAND2_X1 U6440 ( .A1(n5317), .A2(n5315), .ZN(n9201) );
  NAND2_X1 U6441 ( .A1(n5321), .A2(n8638), .ZN(n7463) );
  AND3_X1 U6442 ( .A1(n7215), .A2(n5063), .A3(n10898), .ZN(n5321) );
  INV_X1 U6443 ( .A(n5322), .ZN(n7310) );
  NAND4_X1 U6444 ( .A1(n6454), .A2(n6499), .A3(n6455), .A4(n5326), .ZN(n6464)
         );
  NAND4_X1 U6445 ( .A1(n6454), .A2(n6499), .A3(n6455), .A4(n5325), .ZN(n6532)
         );
  NAND2_X1 U6446 ( .A1(n9129), .A2(n5329), .ZN(n9092) );
  NAND2_X1 U6447 ( .A1(n9129), .A2(n9106), .ZN(n8581) );
  NAND4_X1 U6448 ( .A1(n5337), .A2(n5336), .A3(n5335), .A4(n5333), .ZN(n5332)
         );
  AOI21_X1 U6449 ( .B1(n9931), .B2(n5388), .A(n5383), .ZN(n5382) );
  OAI21_X1 U6450 ( .B1(n9931), .B2(n5390), .A(n5382), .ZN(n8482) );
  NOR2_X2 U6451 ( .A1(n5402), .A2(n5401), .ZN(n6388) );
  NAND2_X1 U6452 ( .A1(n5403), .A2(n5404), .ZN(n5401) );
  NAND3_X1 U6453 ( .A1(n5306), .A2(n5056), .A3(n5067), .ZN(n5402) );
  NAND2_X1 U6454 ( .A1(n8474), .A2(n5104), .ZN(n5407) );
  NAND2_X1 U6455 ( .A1(n8174), .A2(n5108), .ZN(n8470) );
  NAND2_X1 U6456 ( .A1(n7961), .A2(n5057), .ZN(n8095) );
  NAND2_X1 U6457 ( .A1(n10103), .A2(n5411), .ZN(n10076) );
  NAND2_X1 U6458 ( .A1(n9978), .A2(n5414), .ZN(n5413) );
  INV_X1 U6459 ( .A(n5415), .ZN(n9977) );
  NAND3_X1 U6460 ( .A1(n7483), .A2(n7484), .A3(n7482), .ZN(n7502) );
  NAND2_X1 U6461 ( .A1(n7483), .A2(n7482), .ZN(n7486) );
  NOR2_X1 U6462 ( .A1(n5712), .A2(n5596), .ZN(n5595) );
  OAI21_X1 U6463 ( .B1(n10616), .B2(n10615), .A(n10614), .ZN(n10622) );
  NAND2_X1 U6464 ( .A1(n5742), .A2(n5711), .ZN(n6435) );
  NAND2_X1 U6465 ( .A1(n7839), .A2(n5044), .ZN(n5421) );
  NAND2_X1 U6466 ( .A1(n8877), .A2(n5430), .ZN(n5429) );
  OAI21_X1 U6467 ( .B1(n6903), .B2(n5434), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n7406) );
  NOR2_X1 U6468 ( .A1(n6903), .A2(n5437), .ZN(n7049) );
  NAND2_X1 U6469 ( .A1(n8892), .A2(n5100), .ZN(n8867) );
  NAND2_X1 U6470 ( .A1(n8867), .A2(n8549), .ZN(n8955) );
  NAND2_X1 U6471 ( .A1(n8867), .A2(n5443), .ZN(n8560) );
  INV_X1 U6472 ( .A(n7998), .ZN(n5453) );
  NAND2_X1 U6473 ( .A1(n7998), .A2(n8680), .ZN(n7999) );
  INV_X1 U6474 ( .A(n5460), .ZN(n8162) );
  INV_X1 U6475 ( .A(n8680), .ZN(n5462) );
  NAND2_X1 U6476 ( .A1(n8364), .A2(n5466), .ZN(n5463) );
  NAND2_X1 U6477 ( .A1(n5463), .A2(n5464), .ZN(n8366) );
  INV_X1 U6478 ( .A(n8775), .ZN(n5472) );
  NAND2_X1 U6479 ( .A1(n10820), .A2(n10851), .ZN(n8624) );
  NAND2_X1 U6480 ( .A1(n6045), .A2(n5491), .ZN(n5490) );
  NAND2_X1 U6481 ( .A1(n6045), .A2(n6044), .ZN(n6064) );
  NAND2_X1 U6482 ( .A1(n5490), .A2(n5493), .ZN(n6116) );
  NAND3_X1 U6483 ( .A1(n8809), .A2(n5096), .A3(n5510), .ZN(n5509) );
  AND2_X2 U6484 ( .A1(n5522), .A2(n5518), .ZN(n5656) );
  NAND3_X1 U6485 ( .A1(n5521), .A2(n5520), .A3(n5519), .ZN(n5518) );
  NAND3_X1 U6486 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .A3(n5523), .ZN(n5522) );
  NAND2_X1 U6487 ( .A1(n6448), .A2(n6445), .ZN(n5525) );
  NAND3_X1 U6488 ( .A1(n5527), .A2(n5526), .A3(n6445), .ZN(n6660) );
  AND2_X2 U6489 ( .A1(n6666), .A2(n5524), .ZN(n6499) );
  NAND2_X1 U6490 ( .A1(n6447), .A2(n6446), .ZN(n6669) );
  NAND2_X1 U6491 ( .A1(n9247), .A2(n5469), .ZN(n5528) );
  NAND2_X1 U6492 ( .A1(n5528), .A2(n5099), .ZN(n9231) );
  NAND2_X1 U6493 ( .A1(n9135), .A2(n5544), .ZN(n5538) );
  NAND2_X1 U6494 ( .A1(n5530), .A2(n5529), .ZN(n8355) );
  NAND2_X1 U6495 ( .A1(n5041), .A2(n9135), .ZN(n5529) );
  AOI21_X1 U6496 ( .B1(n9135), .B2(n9142), .A(n5545), .ZN(n9117) );
  NAND2_X1 U6497 ( .A1(n7764), .A2(n5548), .ZN(n7798) );
  NAND2_X1 U6498 ( .A1(n7798), .A2(n7885), .ZN(n5549) );
  NAND2_X1 U6499 ( .A1(n5549), .A2(n7884), .ZN(n7883) );
  NAND2_X1 U6500 ( .A1(n7522), .A2(n5550), .ZN(n7543) );
  NAND2_X1 U6501 ( .A1(n9216), .A2(n5103), .ZN(n5552) );
  NAND2_X1 U6502 ( .A1(n5552), .A2(n5553), .ZN(n9179) );
  NAND2_X1 U6503 ( .A1(n9483), .A2(n5567), .ZN(n5565) );
  NAND2_X1 U6504 ( .A1(n5570), .A2(n5569), .ZN(n5563) );
  INV_X1 U6505 ( .A(n7425), .ZN(n5579) );
  NAND2_X1 U6506 ( .A1(n7425), .A2(n5572), .ZN(n5571) );
  OR2_X1 U6507 ( .A1(n5582), .A2(n5963), .ZN(n7676) );
  NAND2_X1 U6508 ( .A1(n5582), .A2(n5963), .ZN(n7674) );
  NAND2_X1 U6509 ( .A1(n5583), .A2(n5584), .ZN(n6385) );
  NAND2_X1 U6510 ( .A1(n9477), .A2(n5585), .ZN(n5583) );
  NAND2_X1 U6511 ( .A1(n9523), .A2(n5590), .ZN(n5589) );
  NAND2_X4 U6512 ( .A1(n6435), .A2(n8463), .ZN(n6473) );
  NAND2_X1 U6513 ( .A1(n8380), .A2(n5883), .ZN(n5601) );
  NAND2_X1 U6514 ( .A1(n7038), .A2(n7039), .ZN(n8380) );
  NAND2_X1 U6515 ( .A1(n6388), .A2(n5706), .ZN(n5730) );
  OAI21_X2 U6516 ( .B1(n10106), .B2(n5614), .A(n5612), .ZN(n10065) );
  INV_X1 U6517 ( .A(n9971), .ZN(n5622) );
  NAND2_X1 U6518 ( .A1(n9802), .A2(n5629), .ZN(n5628) );
  OAI21_X1 U6519 ( .B1(n7865), .B2(n5633), .A(n5630), .ZN(n8085) );
  NOR2_X2 U6520 ( .A1(n7954), .A2(n5635), .ZN(n5634) );
  NAND2_X1 U6521 ( .A1(n7416), .A2(n9602), .ZN(n7473) );
  XNOR2_X2 U6522 ( .A(n7246), .B(n10870), .ZN(n9762) );
  NAND2_X1 U6523 ( .A1(n5722), .A2(n5639), .ZN(n5740) );
  NAND3_X1 U6524 ( .A1(n5697), .A2(n5698), .A3(n10592), .ZN(n5713) );
  NOR2_X2 U6525 ( .A1(n10135), .A2(n10216), .ZN(n10114) );
  NAND2_X1 U6526 ( .A1(n6512), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U6527 ( .A1(n8541), .A2(n8540), .ZN(n8892) );
  AOI21_X1 U6528 ( .B1(n8819), .B2(n7176), .A(n6578), .ZN(n7029) );
  AND2_X1 U6529 ( .A1(n8819), .A2(n10830), .ZN(n10971) );
  NAND2_X1 U6530 ( .A1(n8266), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6550) );
  OR2_X1 U6531 ( .A1(n8253), .A2(n10775), .ZN(n6549) );
  NAND2_X1 U6532 ( .A1(n8445), .A2(n8428), .ZN(n8444) );
  CLKBUF_X1 U6533 ( .A(n9261), .Z(n9266) );
  NOR2_X2 U6534 ( .A1(n10179), .A2(n9993), .ZN(n9986) );
  NAND2_X2 U6535 ( .A1(n7801), .A2(n8684), .ZN(n8007) );
  AND2_X2 U6536 ( .A1(n8496), .A2(n5748), .ZN(n5804) );
  XNOR2_X1 U6537 ( .A(n5874), .B(n5913), .ZN(n5881) );
  CLKBUF_X1 U6538 ( .A(n8064), .Z(n10998) );
  BUF_X1 U6539 ( .A(n5740), .Z(n5742) );
  AND2_X1 U6540 ( .A1(n9231), .A2(n9230), .ZN(n9366) );
  OR2_X1 U6541 ( .A1(n9103), .A2(n8321), .ZN(n8328) );
  OR2_X1 U6542 ( .A1(n9127), .A2(n8321), .ZN(n8313) );
  OR2_X1 U6543 ( .A1(n8321), .A2(n10824), .ZN(n6551) );
  OR2_X1 U6544 ( .A1(n8321), .A2(n10785), .ZN(n6542) );
  OR2_X1 U6545 ( .A1(n8321), .A2(n10451), .ZN(n6525) );
  OAI21_X1 U6546 ( .B1(n7284), .B2(n7243), .A(n7242), .ZN(n7272) );
  AND2_X1 U6547 ( .A1(n10042), .A2(n8473), .ZN(n5641) );
  INV_X1 U6548 ( .A(n9283), .ZN(n8211) );
  OR2_X1 U6549 ( .A1(n10208), .A2(n9499), .ZN(n5642) );
  OR2_X1 U6550 ( .A1(n9236), .A2(n9212), .ZN(n5644) );
  AND2_X1 U6551 ( .A1(n5724), .A2(n10634), .ZN(n5646) );
  AND3_X1 U6552 ( .A1(n10619), .A2(n10415), .A3(n10618), .ZN(n5647) );
  INV_X1 U6553 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8276) );
  INV_X1 U6554 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6533) );
  AND2_X1 U6555 ( .A1(n6411), .A2(n6413), .ZN(n9525) );
  AND2_X1 U6556 ( .A1(n6065), .A2(n6048), .ZN(n5649) );
  AND2_X1 U6557 ( .A1(n5998), .A2(n5749), .ZN(n5650) );
  NAND2_X2 U6558 ( .A1(n7605), .A2(n10090), .ZN(n10093) );
  INV_X1 U6559 ( .A(n5668), .ZN(n6535) );
  INV_X1 U6560 ( .A(n7284), .ZN(n7285) );
  NAND2_X1 U6561 ( .A1(n7284), .A2(n7291), .ZN(n7290) );
  NAND2_X1 U6562 ( .A1(n5783), .A2(n6936), .ZN(n5800) );
  OR3_X1 U6563 ( .A1(n8814), .A2(n8233), .A3(n10994), .ZN(n5651) );
  INV_X1 U6564 ( .A(n10753), .ZN(n5775) );
  OR2_X1 U6565 ( .A1(n9998), .A2(n9508), .ZN(n5652) );
  OR2_X1 U6566 ( .A1(n6514), .A2(n10971), .ZN(n8953) );
  NAND2_X2 U6567 ( .A1(n7214), .A2(n10823), .ZN(n10829) );
  AND2_X1 U6568 ( .A1(n7490), .A2(n7489), .ZN(n5653) );
  INV_X1 U6569 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5704) );
  INV_X1 U6570 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n10634) );
  NOR3_X1 U6571 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n6455) );
  NAND2_X1 U6572 ( .A1(n10203), .A2(n10040), .ZN(n8473) );
  INV_X1 U6573 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5707) );
  OR2_X1 U6574 ( .A1(n9474), .A2(n9475), .ZN(n6343) );
  INV_X1 U6575 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5706) );
  INV_X1 U6576 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U6577 ( .A1(n6553), .A2(n8535), .ZN(n6554) );
  INV_X1 U6578 ( .A(n8049), .ZN(n6923) );
  AND2_X1 U6579 ( .A1(n9341), .A2(n9155), .ZN(n8274) );
  INV_X1 U6580 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10361) );
  INV_X1 U6581 ( .A(n8773), .ZN(n7548) );
  INV_X1 U6582 ( .A(P2_B_REG_SCAN_IN), .ZN(n10547) );
  INV_X1 U6583 ( .A(n8807), .ZN(n8796) );
  INV_X1 U6584 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U6585 ( .A1(n5871), .A2(n8416), .ZN(n5872) );
  AND2_X1 U6586 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n6424), .ZN(n6425) );
  INV_X1 U6587 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U6588 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n10633), .ZN(n5709) );
  INV_X1 U6589 ( .A(n10096), .ZN(n10208) );
  INV_X1 U6590 ( .A(SI_26_), .ZN(n10309) );
  INV_X1 U6591 ( .A(SI_20_), .ZN(n10485) );
  INV_X1 U6592 ( .A(SI_16_), .ZN(n6117) );
  INV_X1 U6593 ( .A(SI_13_), .ZN(n10466) );
  INV_X1 U6594 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10357) );
  NAND2_X1 U6595 ( .A1(n6924), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8216) );
  AND2_X1 U6596 ( .A1(n8082), .A2(n8072), .ZN(n8073) );
  AND2_X1 U6597 ( .A1(n8914), .A2(n8531), .ZN(n8532) );
  AND2_X1 U6598 ( .A1(n7383), .A2(n7372), .ZN(n7373) );
  NAND2_X1 U6599 ( .A1(n6923), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8163) );
  OR2_X1 U6600 ( .A1(n8294), .A2(n10461), .ZN(n8306) );
  INV_X1 U6601 ( .A(n7118), .ZN(n6730) );
  OR2_X1 U6602 ( .A1(n8216), .A2(n10361), .ZN(n8225) );
  OR2_X1 U6603 ( .A1(n7985), .A2(n10521), .ZN(n8049) );
  NAND2_X1 U6604 ( .A1(n6279), .A2(n6278), .ZN(n6280) );
  OR2_X1 U6605 ( .A1(n6155), .A2(n6154), .ZN(n6183) );
  NAND2_X1 U6606 ( .A1(n5873), .A2(n5872), .ZN(n5874) );
  NOR2_X1 U6607 ( .A1(n6269), .A2(n9528), .ZN(n6292) );
  NAND2_X1 U6608 ( .A1(n9425), .A2(n9426), .ZN(n6111) );
  NOR2_X1 U6609 ( .A1(n6183), .A2(n6182), .ZN(n6203) );
  OR2_X1 U6610 ( .A1(n5973), .A2(n5972), .ZN(n5996) );
  NAND2_X1 U6611 ( .A1(n5710), .A2(n5709), .ZN(n5711) );
  AND2_X1 U6612 ( .A1(n6098), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6124) );
  INV_X1 U6613 ( .A(n5765), .ZN(n7262) );
  INV_X1 U6614 ( .A(n7558), .ZN(n7503) );
  AOI21_X1 U6615 ( .B1(n7473), .B2(n9605), .A(n9601), .ZN(n7507) );
  OR2_X1 U6616 ( .A1(n8332), .A2(n8573), .ZN(n8348) );
  OR2_X1 U6617 ( .A1(n8252), .A2(n10357), .ZN(n8264) );
  AND2_X1 U6618 ( .A1(n7360), .A2(n7099), .ZN(n7100) );
  OR2_X1 U6619 ( .A1(n8953), .A2(n8562), .ZN(n8922) );
  OR2_X1 U6620 ( .A1(n7845), .A2(n9270), .ZN(n8964) );
  INV_X1 U6621 ( .A(n8321), .ZN(n8353) );
  INV_X2 U6622 ( .A(n5037), .ZN(n8616) );
  INV_X1 U6623 ( .A(n9154), .ZN(n9152) );
  INV_X1 U6624 ( .A(n7234), .ZN(n6589) );
  AOI21_X1 U6625 ( .B1(n8207), .B2(n8206), .A(n5075), .ZN(n9288) );
  INV_X1 U6626 ( .A(n10822), .ZN(n9264) );
  INV_X1 U6627 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9416) );
  INV_X1 U6628 ( .A(n6459), .ZN(n6460) );
  NOR2_X1 U6629 ( .A1(n5928), .A2(n5927), .ZN(n5953) );
  NAND2_X1 U6630 ( .A1(n6385), .A2(n6384), .ZN(n6386) );
  NOR2_X1 U6631 ( .A1(n8426), .A2(n9569), .ZN(n8427) );
  OR2_X1 U6632 ( .A1(n6241), .A2(n6240), .ZN(n6269) );
  INV_X1 U6633 ( .A(n10129), .ZN(n10082) );
  AND3_X1 U6634 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5898) );
  INV_X1 U6635 ( .A(n6413), .ZN(n6938) );
  OR2_X1 U6636 ( .A1(n6429), .A2(n9923), .ZN(n6432) );
  INV_X1 U6637 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6885) );
  NAND2_X1 U6638 ( .A1(n9953), .A2(n10131), .ZN(n9914) );
  INV_X1 U6639 ( .A(n8146), .ZN(n10983) );
  INV_X1 U6640 ( .A(n10131), .ZN(n10081) );
  INV_X1 U6641 ( .A(n8964), .ZN(n8960) );
  NAND2_X1 U6642 ( .A1(n8803), .A2(n8802), .ZN(n8817) );
  AND4_X1 U6643 ( .A1(n8231), .A2(n8230), .A3(n8229), .A4(n8228), .ZN(n9271)
         );
  INV_X1 U6644 ( .A(n10773), .ZN(n10809) );
  INV_X1 U6645 ( .A(n10801), .ZN(n10776) );
  INV_X1 U6646 ( .A(n10792), .ZN(n10807) );
  INV_X1 U6647 ( .A(n10818), .ZN(n9226) );
  INV_X1 U6648 ( .A(n9270), .ZN(n10821) );
  INV_X1 U6649 ( .A(n9300), .ZN(n10827) );
  AND4_X1 U6650 ( .A1(n7235), .A2(n7231), .A3(n7234), .A4(n7232), .ZN(n7195)
         );
  NAND2_X1 U6651 ( .A1(n8551), .A2(n7177), .ZN(n10990) );
  INV_X1 U6652 ( .A(n10994), .ZN(n10881) );
  INV_X1 U6653 ( .A(n10700), .ZN(n10701) );
  XNOR2_X1 U6654 ( .A(n6463), .B(P2_IR_REG_24__SCAN_IN), .ZN(n6478) );
  AND2_X1 U6655 ( .A1(n6699), .A2(n6697), .ZN(n7749) );
  INV_X1 U6656 ( .A(n9559), .ZN(n9532) );
  NAND2_X1 U6657 ( .A1(n6423), .A2(n6939), .ZN(n9505) );
  INV_X1 U6658 ( .A(n6417), .ZN(n9828) );
  AND4_X1 U6659 ( .A1(n6434), .A2(n6433), .A3(n6432), .A4(n6431), .ZN(n9934)
         );
  AND2_X1 U6660 ( .A1(n6229), .A2(n6228), .ZN(n9451) );
  INV_X1 U6661 ( .A(n9899), .ZN(n10760) );
  INV_X1 U6662 ( .A(n9788), .ZN(n9937) );
  AND2_X1 U6663 ( .A1(n7265), .A2(n9830), .ZN(n10131) );
  AND2_X1 U6664 ( .A1(n10093), .A2(n7077), .ZN(n10095) );
  OR2_X1 U6665 ( .A1(n7293), .A2(n9798), .ZN(n11009) );
  OR2_X1 U6666 ( .A1(n9731), .A2(n9798), .ZN(n10923) );
  INV_X1 U6667 ( .A(n10259), .ZN(n6899) );
  INV_X1 U6668 ( .A(n6406), .ZN(n10665) );
  AND2_X1 U6669 ( .A1(n6177), .A2(n6149), .ZN(n9875) );
  AND2_X1 U6670 ( .A1(n6022), .A2(n6049), .ZN(n6643) );
  AND2_X1 U6671 ( .A1(n5949), .A2(n5967), .ZN(n6675) );
  INV_X1 U6672 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7896) );
  NOR2_X1 U6673 ( .A1(n10716), .A2(n7905), .ZN(n7906) );
  NOR2_X1 U6674 ( .A1(n10727), .A2(n10726), .ZN(n7923) );
  INV_X1 U6675 ( .A(n10787), .ZN(n10800) );
  INV_X1 U6676 ( .A(n9162), .ZN(n9334) );
  AND3_X1 U6677 ( .A1(n8202), .A2(n8201), .A3(n8200), .ZN(n9213) );
  INV_X1 U6678 ( .A(n8871), .ZN(n8981) );
  NAND2_X1 U6679 ( .A1(n6787), .A2(n6784), .ZN(n10801) );
  XNOR2_X1 U6680 ( .A(n8355), .B(n8354), .ZN(n9315) );
  OR2_X1 U6681 ( .A1(n7214), .A2(n8535), .ZN(n10818) );
  INV_X1 U6682 ( .A(n11002), .ZN(n11000) );
  INV_X1 U6683 ( .A(n11006), .ZN(n11003) );
  NAND2_X1 U6684 ( .A1(n10702), .A2(n10701), .ZN(n10769) );
  INV_X1 U6685 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8271) );
  INV_X1 U6686 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7048) );
  INV_X1 U6687 ( .A(n9505), .ZN(n9564) );
  AND2_X1 U6688 ( .A1(n6414), .A2(n10090), .ZN(n9535) );
  INV_X1 U6689 ( .A(n9525), .ZN(n9569) );
  INV_X1 U6690 ( .A(n8450), .ZN(n9982) );
  INV_X1 U6691 ( .A(n8117), .ZN(n9843) );
  OR2_X1 U6692 ( .A1(n6908), .A2(n6979), .ZN(n9869) );
  OR2_X1 U6693 ( .A1(n6908), .A2(n9830), .ZN(n9899) );
  NAND2_X1 U6694 ( .A1(n10093), .A2(n7289), .ZN(n10148) );
  AND2_X2 U6695 ( .A1(n6900), .A2(n10259), .ZN(n11024) );
  AND3_X1 U6696 ( .A1(n10952), .A2(n10951), .A3(n10950), .ZN(n10954) );
  AND2_X2 U6697 ( .A1(n6900), .A2(n6899), .ZN(n11028) );
  CLKBUF_X1 U6698 ( .A(n10698), .Z(n10686) );
  INV_X1 U6699 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10571) );
  INV_X1 U6700 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10568) );
  NOR2_X1 U6701 ( .A1(n7924), .A2(n7923), .ZN(n10729) );
  MUX2_X1 U6702 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5663), .Z(n5661) );
  INV_X1 U6703 ( .A(SI_2_), .ZN(n5654) );
  XNOR2_X1 U6704 ( .A(n5661), .B(n5654), .ZN(n5811) );
  NAND3_X1 U6705 ( .A1(n5663), .A2(SI_0_), .A3(P2_DATAO_REG_0__SCAN_IN), .ZN(
        n5657) );
  AND2_X1 U6706 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5655) );
  MUX2_X1 U6707 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5663), .Z(n5790) );
  NAND2_X1 U6708 ( .A1(n5791), .A2(n5790), .ZN(n5660) );
  NAND2_X1 U6709 ( .A1(n5658), .A2(SI_1_), .ZN(n5659) );
  NAND2_X1 U6710 ( .A1(n5660), .A2(n5659), .ZN(n5812) );
  NAND2_X1 U6711 ( .A1(n5661), .A2(SI_2_), .ZN(n5662) );
  INV_X1 U6712 ( .A(SI_3_), .ZN(n5664) );
  XNOR2_X1 U6713 ( .A(n5665), .B(n5664), .ZN(n5839) );
  NAND2_X1 U6714 ( .A1(n5840), .A2(n5839), .ZN(n5667) );
  NAND2_X1 U6715 ( .A1(n5665), .A2(SI_3_), .ZN(n5666) );
  MUX2_X1 U6716 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5668), .Z(n5669) );
  INV_X1 U6717 ( .A(SI_4_), .ZN(n10307) );
  XNOR2_X1 U6718 ( .A(n5669), .B(n10307), .ZN(n5862) );
  NAND2_X1 U6719 ( .A1(n5863), .A2(n5862), .ZN(n5671) );
  NAND2_X1 U6720 ( .A1(n5669), .A2(SI_4_), .ZN(n5670) );
  MUX2_X1 U6721 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5668), .Z(n5673) );
  INV_X1 U6722 ( .A(SI_5_), .ZN(n5672) );
  XNOR2_X1 U6723 ( .A(n5673), .B(n5672), .ZN(n5890) );
  NAND2_X1 U6724 ( .A1(n5891), .A2(n5890), .ZN(n5675) );
  NAND2_X1 U6725 ( .A1(n5673), .A2(SI_5_), .ZN(n5674) );
  MUX2_X1 U6726 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5668), .Z(n5676) );
  INV_X1 U6727 ( .A(SI_6_), .ZN(n10338) );
  XNOR2_X1 U6728 ( .A(n5676), .B(n10338), .ZN(n5904) );
  NAND2_X1 U6729 ( .A1(n5905), .A2(n5904), .ZN(n5678) );
  NAND2_X1 U6730 ( .A1(n5676), .A2(SI_6_), .ZN(n5677) );
  NAND2_X1 U6731 ( .A1(n5678), .A2(n5677), .ZN(n5921) );
  MUX2_X1 U6732 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5668), .Z(n5680) );
  INV_X1 U6733 ( .A(SI_7_), .ZN(n5679) );
  XNOR2_X1 U6734 ( .A(n5680), .B(n5679), .ZN(n5920) );
  NAND2_X1 U6735 ( .A1(n5921), .A2(n5920), .ZN(n5682) );
  NAND2_X1 U6736 ( .A1(n5680), .A2(SI_7_), .ZN(n5681) );
  INV_X1 U6737 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7524) );
  INV_X1 U6738 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6676) );
  MUX2_X1 U6739 ( .A(n7524), .B(n6676), .S(n5668), .Z(n5683) );
  XNOR2_X1 U6740 ( .A(n5683), .B(SI_8_), .ZN(n5944) );
  NAND2_X1 U6741 ( .A1(n5946), .A2(n5944), .ZN(n5686) );
  INV_X1 U6742 ( .A(n5683), .ZN(n5684) );
  NAND2_X1 U6743 ( .A1(n5684), .A2(SI_8_), .ZN(n5685) );
  INV_X1 U6744 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6685) );
  MUX2_X1 U6745 ( .A(n6685), .B(n10272), .S(n5668), .Z(n5688) );
  INV_X1 U6746 ( .A(SI_9_), .ZN(n5687) );
  NAND2_X1 U6747 ( .A1(n5688), .A2(n5687), .ZN(n5691) );
  INV_X1 U6748 ( .A(n5688), .ZN(n5689) );
  NAND2_X1 U6749 ( .A1(n5689), .A2(SI_9_), .ZN(n5690) );
  NAND2_X1 U6750 ( .A1(n5691), .A2(n5690), .ZN(n5965) );
  MUX2_X1 U6751 ( .A(n6698), .B(n5992), .S(n5668), .Z(n5693) );
  NAND2_X1 U6752 ( .A1(n5693), .A2(n10498), .ZN(n5696) );
  INV_X1 U6753 ( .A(n5693), .ZN(n5694) );
  NAND2_X1 U6754 ( .A1(n5694), .A2(SI_10_), .ZN(n5695) );
  MUX2_X1 U6755 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n5668), .Z(n6014) );
  NOR2_X2 U6756 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5698) );
  NOR2_X2 U6757 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5697) );
  NOR2_X1 U6758 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5701) );
  NOR2_X1 U6759 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5700) );
  NOR2_X1 U6760 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5699) );
  NAND4_X1 U6761 ( .A1(n5701), .A2(n5700), .A3(n5699), .A4(n10593), .ZN(n5702)
         );
  INV_X2 U6762 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10608) );
  NAND4_X1 U6763 ( .A1(n10608), .A2(n10628), .A3(n10618), .A4(n5735), .ZN(
        n5703) );
  NOR2_X1 U6764 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5705) );
  OR2_X1 U6765 ( .A1(n5712), .A2(n10261), .ZN(n5708) );
  NAND2_X1 U6766 ( .A1(n5708), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U6767 ( .A1(n7781), .A2(n6176), .ZN(n5721) );
  INV_X1 U6768 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10279) );
  NOR2_X1 U6769 ( .A1(n5714), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5906) );
  NOR2_X1 U6770 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5715) );
  NAND2_X1 U6771 ( .A1(n5906), .A2(n5715), .ZN(n5947) );
  NAND2_X1 U6772 ( .A1(n5716), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5991) );
  INV_X1 U6773 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U6774 ( .A1(n5991), .A2(n5990), .ZN(n5989) );
  NAND2_X1 U6775 ( .A1(n5989), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5718) );
  INV_X1 U6776 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5717) );
  XNOR2_X1 U6777 ( .A(n5718), .B(n5717), .ZN(n6920) );
  OAI22_X1 U6778 ( .A1(n6199), .A2(n10279), .B1(n6473), .B2(n6920), .ZN(n5719)
         );
  INV_X1 U6779 ( .A(n5719), .ZN(n5720) );
  NAND2_X2 U6780 ( .A1(n5721), .A2(n5720), .ZN(n8020) );
  INV_X1 U6781 ( .A(n5723), .ZN(n5733) );
  NAND2_X1 U6782 ( .A1(n5728), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U6783 ( .A1(n5727), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U6784 ( .A1(n5730), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5731) );
  MUX2_X1 U6785 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5731), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5732) );
  NAND2_X1 U6786 ( .A1(n5738), .A2(n5758), .ZN(n5762) );
  AND2_X4 U6787 ( .A1(n6471), .A2(n7248), .ZN(n8416) );
  NAND2_X1 U6788 ( .A1(n8020), .A2(n8416), .ZN(n5757) );
  XNOR2_X2 U6789 ( .A(n5741), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5747) );
  NAND2_X1 U6790 ( .A1(n5742), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5743) );
  INV_X1 U6791 ( .A(n5744), .ZN(n10262) );
  NAND2_X1 U6792 ( .A1(n5040), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5754) );
  INV_X1 U6793 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5746) );
  OR2_X1 U6794 ( .A1(n8430), .A2(n5746), .ZN(n5753) );
  AND2_X4 U6795 ( .A1(n5747), .A2(n5748), .ZN(n5855) );
  NAND2_X1 U6796 ( .A1(n5898), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U6797 ( .A1(n5953), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5973) );
  OR2_X1 U6798 ( .A1(n5650), .A2(n6027), .ZN(n8018) );
  OR2_X1 U6799 ( .A1(n6429), .A2(n8018), .ZN(n5752) );
  INV_X1 U6800 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5750) );
  OR2_X1 U6801 ( .A1(n8432), .A2(n5750), .ZN(n5751) );
  INV_X1 U6802 ( .A(n5755), .ZN(n5779) );
  NAND2_X1 U6803 ( .A1(n9844), .A2(n8422), .ZN(n5756) );
  NAND2_X1 U6804 ( .A1(n5757), .A2(n5756), .ZN(n5764) );
  NAND2_X1 U6805 ( .A1(n5760), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5761) );
  XNOR2_X1 U6806 ( .A(n5764), .B(n7288), .ZN(n6011) );
  INV_X1 U6807 ( .A(n6011), .ZN(n6013) );
  NAND2_X1 U6808 ( .A1(n5765), .A2(n6417), .ZN(n5766) );
  AND2_X2 U6809 ( .A1(n5766), .A2(n8416), .ZN(n5778) );
  AOI22_X1 U6810 ( .A1(n8020), .A2(n8422), .B1(n5778), .B2(n9844), .ZN(n6012)
         );
  INV_X1 U6811 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5767) );
  NAND2_X1 U6812 ( .A1(n5768), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U6813 ( .A1(n5668), .A2(SI_0_), .ZN(n5773) );
  XNOR2_X1 U6814 ( .A(n5773), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10664) );
  AOI22_X1 U6815 ( .A1(n7296), .A2(n8416), .B1(n5779), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n5776) );
  NAND2_X1 U6816 ( .A1(n5777), .A2(n7288), .ZN(n5783) );
  NAND2_X1 U6817 ( .A1(n6891), .A2(n5778), .ZN(n5782) );
  AND2_X1 U6818 ( .A1(n5779), .A2(n10753), .ZN(n5780) );
  AND2_X1 U6819 ( .A1(n5782), .A2(n5781), .ZN(n6937) );
  NAND2_X1 U6820 ( .A1(n6937), .A2(n6935), .ZN(n6936) );
  NAND2_X1 U6821 ( .A1(n5768), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U6822 ( .A1(n5855), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5787) );
  INV_X1 U6823 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5784) );
  OR2_X1 U6824 ( .A1(n5806), .A2(n5784), .ZN(n5786) );
  NAND2_X1 U6825 ( .A1(n5804), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U6826 ( .A1(n7241), .A2(n8422), .ZN(n5797) );
  NAND2_X1 U6827 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n10753), .ZN(n5789) );
  XNOR2_X1 U6828 ( .A(n5789), .B(P1_IR_REG_1__SCAN_IN), .ZN(n10759) );
  NAND2_X1 U6829 ( .A1(n5814), .A2(n10759), .ZN(n5795) );
  XNOR2_X1 U6830 ( .A(n5791), .B(n5790), .ZN(n6658) );
  NAND2_X1 U6831 ( .A1(n6658), .A2(n5668), .ZN(n5793) );
  INV_X1 U6832 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6654) );
  NAND2_X1 U6833 ( .A1(n6535), .A2(n6654), .ZN(n5792) );
  NAND3_X1 U6834 ( .A1(n6473), .A2(n5793), .A3(n5792), .ZN(n5794) );
  NAND2_X1 U6835 ( .A1(n10839), .A2(n8416), .ZN(n5796) );
  NAND2_X1 U6836 ( .A1(n5797), .A2(n5796), .ZN(n5798) );
  XNOR2_X1 U6837 ( .A(n5800), .B(n5801), .ZN(n9457) );
  INV_X2 U6838 ( .A(n10839), .ZN(n9593) );
  NOR2_X1 U6839 ( .A1(n9593), .A2(n6208), .ZN(n5799) );
  AOI21_X1 U6840 ( .B1(n9851), .B2(n5778), .A(n5799), .ZN(n9458) );
  NAND2_X1 U6841 ( .A1(n9457), .A2(n9458), .ZN(n9456) );
  INV_X1 U6842 ( .A(n5801), .ZN(n5802) );
  NAND2_X1 U6843 ( .A1(n5800), .A2(n5802), .ZN(n5803) );
  NAND2_X1 U6844 ( .A1(n9456), .A2(n5803), .ZN(n6971) );
  NAND2_X1 U6845 ( .A1(n5855), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5810) );
  INV_X1 U6846 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6599) );
  OR2_X1 U6847 ( .A1(n5854), .A2(n6599), .ZN(n5809) );
  NAND2_X1 U6848 ( .A1(n5804), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5808) );
  INV_X1 U6849 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5805) );
  OR2_X1 U6850 ( .A1(n5806), .A2(n5805), .ZN(n5807) );
  NAND4_X2 U6851 ( .A1(n5810), .A2(n5809), .A3(n5808), .A4(n5807), .ZN(n9850)
         );
  NAND2_X1 U6852 ( .A1(n9850), .A2(n8422), .ZN(n5824) );
  XNOR2_X1 U6853 ( .A(n5812), .B(n5811), .ZN(n6673) );
  INV_X1 U6854 ( .A(n6673), .ZN(n5813) );
  NOR2_X1 U6855 ( .A1(n10753), .A2(P1_IR_REG_1__SCAN_IN), .ZN(n5817) );
  INV_X1 U6856 ( .A(n5817), .ZN(n5815) );
  NAND2_X1 U6857 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5815), .ZN(n5816) );
  INV_X1 U6858 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n10583) );
  MUX2_X1 U6859 ( .A(n5816), .B(P1_IR_REG_31__SCAN_IN), .S(n10583), .Z(n5818)
         );
  NAND2_X1 U6860 ( .A1(n10583), .A2(n5817), .ZN(n5843) );
  AND2_X1 U6861 ( .A1(n5818), .A2(n5843), .ZN(n6672) );
  NAND2_X1 U6862 ( .A1(n5814), .A2(n6672), .ZN(n5821) );
  INV_X1 U6863 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U6864 ( .A1(n5824), .A2(n5823), .ZN(n5825) );
  NAND2_X1 U6865 ( .A1(n9850), .A2(n5778), .ZN(n5827) );
  OR2_X1 U6866 ( .A1(n10857), .A2(n6208), .ZN(n5826) );
  NAND2_X1 U6867 ( .A1(n5827), .A2(n5826), .ZN(n5828) );
  XNOR2_X1 U6868 ( .A(n5830), .B(n5828), .ZN(n6970) );
  NAND2_X1 U6869 ( .A1(n6971), .A2(n6970), .ZN(n5832) );
  INV_X1 U6870 ( .A(n5828), .ZN(n5829) );
  NAND2_X1 U6871 ( .A1(n5830), .A2(n5829), .ZN(n5831) );
  NAND2_X1 U6872 ( .A1(n5832), .A2(n5831), .ZN(n7038) );
  OR2_X1 U6873 ( .A1(n6429), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5837) );
  INV_X1 U6874 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U6875 ( .A1(n5040), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5835) );
  OR2_X1 U6876 ( .A1(n8430), .A2(n6597), .ZN(n5834) );
  NAND2_X1 U6877 ( .A1(n7246), .A2(n5778), .ZN(n5849) );
  XNOR2_X1 U6878 ( .A(n5840), .B(n5839), .ZN(n6665) );
  INV_X1 U6879 ( .A(n6665), .ZN(n5841) );
  NAND2_X1 U6880 ( .A1(n5838), .A2(n5841), .ZN(n5847) );
  NAND2_X1 U6881 ( .A1(n9574), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5846) );
  NAND2_X1 U6882 ( .A1(n5843), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5844) );
  XNOR2_X1 U6883 ( .A(n5844), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6858) );
  NAND2_X1 U6884 ( .A1(n5814), .A2(n6858), .ZN(n5845) );
  OR2_X1 U6885 ( .A1(n10870), .A2(n6208), .ZN(n5848) );
  NAND2_X1 U6886 ( .A1(n5849), .A2(n5848), .ZN(n5851) );
  NAND2_X1 U6887 ( .A1(n7246), .A2(n8422), .ZN(n5850) );
  XNOR2_X1 U6888 ( .A(n5851), .B(n5853), .ZN(n7039) );
  INV_X1 U6889 ( .A(n5851), .ZN(n5852) );
  NAND2_X1 U6890 ( .A1(n5853), .A2(n5852), .ZN(n8379) );
  INV_X1 U6891 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6605) );
  INV_X1 U6892 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5856) );
  XNOR2_X1 U6893 ( .A(n5856), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n8386) );
  NAND2_X1 U6894 ( .A1(n5855), .A2(n8386), .ZN(n5859) );
  INV_X1 U6895 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5857) );
  OR2_X1 U6896 ( .A1(n5806), .A2(n5857), .ZN(n5858) );
  NAND2_X1 U6897 ( .A1(n5040), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U6898 ( .A1(n5875), .A2(n8422), .ZN(n5873) );
  XNOR2_X1 U6899 ( .A(n5863), .B(n5862), .ZN(n7095) );
  INV_X1 U6900 ( .A(n7095), .ZN(n5864) );
  NAND2_X1 U6901 ( .A1(n5838), .A2(n5864), .ZN(n5870) );
  NAND2_X1 U6902 ( .A1(n9574), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5869) );
  NOR2_X1 U6903 ( .A1(n5865), .A2(n10261), .ZN(n5866) );
  MUX2_X1 U6904 ( .A(n10261), .B(n5866), .S(P1_IR_REG_4__SCAN_IN), .Z(n5867)
         );
  NOR2_X1 U6905 ( .A1(n5867), .A2(n5403), .ZN(n6626) );
  NAND2_X1 U6906 ( .A1(n5814), .A2(n6626), .ZN(n5868) );
  INV_X1 U6907 ( .A(n5881), .ZN(n5878) );
  NAND2_X1 U6908 ( .A1(n5875), .A2(n5778), .ZN(n5877) );
  OR2_X1 U6909 ( .A1(n7411), .A2(n6208), .ZN(n5876) );
  NAND2_X1 U6910 ( .A1(n5877), .A2(n5876), .ZN(n5880) );
  AND2_X1 U6911 ( .A1(n8379), .A2(n5879), .ZN(n5883) );
  INV_X1 U6912 ( .A(n5879), .ZN(n5882) );
  XNOR2_X1 U6913 ( .A(n5881), .B(n5880), .ZN(n8382) );
  NAND2_X1 U6914 ( .A1(n5040), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5889) );
  AOI21_X1 U6915 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5884) );
  NOR2_X1 U6916 ( .A1(n5884), .A2(n5898), .ZN(n7476) );
  NAND2_X1 U6917 ( .A1(n5855), .A2(n7476), .ZN(n5888) );
  INV_X1 U6918 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7478) );
  OR2_X1 U6919 ( .A1(n8430), .A2(n7478), .ZN(n5887) );
  INV_X1 U6920 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5885) );
  OR2_X1 U6921 ( .A1(n8432), .A2(n5885), .ZN(n5886) );
  NAND2_X1 U6922 ( .A1(n9849), .A2(n8422), .ZN(n5896) );
  XNOR2_X1 U6923 ( .A(n5891), .B(n5890), .ZN(n7103) );
  NAND2_X1 U6924 ( .A1(n9574), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U6925 ( .A1(n5714), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5892) );
  XNOR2_X1 U6926 ( .A(n5892), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6711) );
  NAND2_X1 U6927 ( .A1(n5814), .A2(n6711), .ZN(n5893) );
  NAND2_X1 U6928 ( .A1(n7500), .A2(n8416), .ZN(n5895) );
  NAND2_X1 U6929 ( .A1(n5896), .A2(n5895), .ZN(n5897) );
  AOI22_X1 U6930 ( .A1(n9849), .A2(n5778), .B1(n8422), .B2(n7500), .ZN(n7062)
         );
  NAND2_X1 U6931 ( .A1(n5040), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5903) );
  INV_X1 U6932 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7513) );
  OR2_X1 U6933 ( .A1(n8430), .A2(n7513), .ZN(n5902) );
  OAI21_X1 U6934 ( .B1(n5898), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5928), .ZN(
        n7517) );
  OR2_X1 U6935 ( .A1(n6429), .A2(n7517), .ZN(n5901) );
  INV_X1 U6936 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5899) );
  OR2_X1 U6937 ( .A1(n8432), .A2(n5899), .ZN(n5900) );
  XNOR2_X1 U6938 ( .A(n5905), .B(n5904), .ZN(n7325) );
  OR2_X1 U6939 ( .A1(n8453), .A2(n7325), .ZN(n5912) );
  INV_X1 U6940 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10584) );
  OR2_X1 U6941 ( .A1(n5906), .A2(n10261), .ZN(n5908) );
  INV_X1 U6942 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U6943 ( .A1(n5908), .A2(n5907), .ZN(n5922) );
  OR2_X1 U6944 ( .A1(n5908), .A2(n5907), .ZN(n5909) );
  NAND2_X1 U6945 ( .A1(n5922), .A2(n5909), .ZN(n6872) );
  OAI22_X1 U6946 ( .A1(n6199), .A2(n10584), .B1(n6473), .B2(n6872), .ZN(n5910)
         );
  INV_X1 U6947 ( .A(n5910), .ZN(n5911) );
  NAND2_X1 U6948 ( .A1(n5912), .A2(n5911), .ZN(n10903) );
  OAI22_X1 U6949 ( .A1(n7572), .A2(n6208), .B1(n7571), .B2(n6300), .ZN(n5914)
         );
  XNOR2_X1 U6950 ( .A(n5914), .B(n5913), .ZN(n7167) );
  AND2_X1 U6951 ( .A1(n10903), .A2(n8422), .ZN(n5915) );
  AOI21_X1 U6952 ( .B1(n9848), .B2(n5778), .A(n5915), .ZN(n7166) );
  INV_X1 U6953 ( .A(n7167), .ZN(n5917) );
  INV_X1 U6954 ( .A(n7166), .ZN(n5916) );
  NAND2_X1 U6955 ( .A1(n5917), .A2(n5916), .ZN(n5918) );
  NAND2_X1 U6956 ( .A1(n5919), .A2(n5918), .ZN(n7425) );
  XNOR2_X1 U6957 ( .A(n5921), .B(n5920), .ZN(n7447) );
  OR2_X1 U6958 ( .A1(n7447), .A2(n8453), .ZN(n5926) );
  INV_X1 U6959 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10586) );
  NAND2_X1 U6960 ( .A1(n5922), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5923) );
  INV_X1 U6961 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n10396) );
  XNOR2_X1 U6962 ( .A(n5923), .B(n10396), .ZN(n6740) );
  OAI22_X1 U6963 ( .A1(n6199), .A2(n10586), .B1(n6473), .B2(n6740), .ZN(n5924)
         );
  INV_X1 U6964 ( .A(n5924), .ZN(n5925) );
  NAND2_X1 U6965 ( .A1(n5040), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5934) );
  AND2_X1 U6966 ( .A1(n5928), .A2(n5927), .ZN(n5929) );
  NOR2_X1 U6967 ( .A1(n5953), .A2(n5929), .ZN(n7606) );
  NAND2_X1 U6968 ( .A1(n5855), .A2(n7606), .ZN(n5933) );
  INV_X1 U6969 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7603) );
  OR2_X1 U6970 ( .A1(n8430), .A2(n7603), .ZN(n5932) );
  INV_X1 U6971 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5930) );
  OR2_X1 U6972 ( .A1(n8432), .A2(n5930), .ZN(n5931) );
  NAND4_X1 U6973 ( .A1(n5934), .A2(n5933), .A3(n5932), .A4(n5931), .ZN(n9847)
         );
  NAND2_X1 U6974 ( .A1(n9847), .A2(n8422), .ZN(n5935) );
  OAI21_X1 U6975 ( .B1(n7608), .B2(n6300), .A(n5935), .ZN(n5936) );
  XNOR2_X1 U6976 ( .A(n5936), .B(n7288), .ZN(n5939) );
  OR2_X1 U6977 ( .A1(n7608), .A2(n6208), .ZN(n5938) );
  NAND2_X1 U6978 ( .A1(n9847), .A2(n5778), .ZN(n5937) );
  NAND2_X1 U6979 ( .A1(n5938), .A2(n5937), .ZN(n5940) );
  XNOR2_X1 U6980 ( .A(n5939), .B(n5940), .ZN(n7424) );
  INV_X1 U6981 ( .A(n5939), .ZN(n5942) );
  INV_X1 U6982 ( .A(n5940), .ZN(n5941) );
  NAND2_X1 U6983 ( .A1(n5942), .A2(n5941), .ZN(n5943) );
  INV_X1 U6984 ( .A(n5944), .ZN(n5945) );
  XNOR2_X1 U6985 ( .A(n5946), .B(n5945), .ZN(n7523) );
  NAND2_X1 U6986 ( .A1(n7523), .A2(n6176), .ZN(n5951) );
  NAND2_X1 U6987 ( .A1(n5947), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5948) );
  MUX2_X1 U6988 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5948), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5949) );
  AOI22_X1 U6989 ( .A1(n9574), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5814), .B2(
        n6675), .ZN(n5950) );
  NAND2_X1 U6990 ( .A1(n5040), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5959) );
  INV_X1 U6991 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5952) );
  OR2_X1 U6992 ( .A1(n8430), .A2(n5952), .ZN(n5958) );
  OR2_X1 U6993 ( .A1(n5953), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U6994 ( .A1(n5973), .A2(n5954), .ZN(n7680) );
  OR2_X1 U6995 ( .A1(n6429), .A2(n7680), .ZN(n5957) );
  INV_X1 U6996 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5955) );
  OR2_X1 U6997 ( .A1(n8432), .A2(n5955), .ZN(n5956) );
  AOI22_X1 U6998 ( .A1(n7679), .A2(n8422), .B1(n7648), .B2(n5778), .ZN(n5963)
         );
  NAND2_X1 U6999 ( .A1(n7679), .A2(n8416), .ZN(n5961) );
  NAND2_X1 U7000 ( .A1(n7648), .A2(n8422), .ZN(n5960) );
  NAND2_X1 U7001 ( .A1(n5961), .A2(n5960), .ZN(n5962) );
  XNOR2_X1 U7002 ( .A(n5962), .B(n7288), .ZN(n7673) );
  INV_X1 U7003 ( .A(n5963), .ZN(n5964) );
  XNOR2_X1 U7004 ( .A(n5966), .B(n5965), .ZN(n7536) );
  NAND2_X1 U7005 ( .A1(n7536), .A2(n6176), .ZN(n5971) );
  NAND2_X1 U7006 ( .A1(n5967), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5968) );
  XNOR2_X1 U7007 ( .A(n5968), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6771) );
  INV_X1 U7008 ( .A(n6771), .ZN(n6682) );
  OAI22_X1 U7009 ( .A1(n6199), .A2(n10272), .B1(n5033), .B2(n6682), .ZN(n5969)
         );
  INV_X1 U7010 ( .A(n5969), .ZN(n5970) );
  NAND2_X2 U7011 ( .A1(n5971), .A2(n5970), .ZN(n10945) );
  NAND2_X1 U7012 ( .A1(n10945), .A2(n8416), .ZN(n5981) );
  NAND2_X1 U7013 ( .A1(n5973), .A2(n5972), .ZN(n5974) );
  NAND2_X1 U7014 ( .A1(n5996), .A2(n5974), .ZN(n7568) );
  OR2_X1 U7015 ( .A1(n6429), .A2(n7568), .ZN(n5979) );
  NAND2_X1 U7016 ( .A1(n5040), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5978) );
  NAND2_X1 U7017 ( .A1(n8458), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5977) );
  INV_X1 U7018 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n5975) );
  OR2_X1 U7019 ( .A1(n8430), .A2(n5975), .ZN(n5976) );
  NAND4_X1 U7020 ( .A1(n5979), .A2(n5978), .A3(n5977), .A4(n5976), .ZN(n9846)
         );
  NAND2_X1 U7021 ( .A1(n9846), .A2(n8422), .ZN(n5980) );
  NAND2_X1 U7022 ( .A1(n5981), .A2(n5980), .ZN(n5982) );
  XNOR2_X1 U7023 ( .A(n5982), .B(n7288), .ZN(n5984) );
  AND2_X1 U7024 ( .A1(n9846), .A2(n5778), .ZN(n5983) );
  AOI21_X1 U7025 ( .B1(n10945), .B2(n8422), .A(n5983), .ZN(n5985) );
  XNOR2_X1 U7026 ( .A(n5984), .B(n5985), .ZN(n7645) );
  INV_X1 U7027 ( .A(n5984), .ZN(n5986) );
  NAND2_X1 U7028 ( .A1(n5986), .A2(n5985), .ZN(n5987) );
  NAND2_X1 U7029 ( .A1(n7748), .A2(n6176), .ZN(n5995) );
  OAI21_X1 U7030 ( .B1(n5991), .B2(n5990), .A(n5989), .ZN(n6886) );
  OAI22_X1 U7031 ( .A1(n6199), .A2(n5992), .B1(n6473), .B2(n6886), .ZN(n5993)
         );
  INV_X1 U7032 ( .A(n5993), .ZN(n5994) );
  NAND2_X2 U7033 ( .A1(n5995), .A2(n5994), .ZN(n7978) );
  NAND2_X1 U7034 ( .A1(n7978), .A2(n8416), .ZN(n6005) );
  NAND2_X1 U7035 ( .A1(n5040), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6003) );
  INV_X1 U7036 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6611) );
  OR2_X1 U7037 ( .A1(n8430), .A2(n6611), .ZN(n6002) );
  NAND2_X1 U7038 ( .A1(n5996), .A2(n6885), .ZN(n5997) );
  NAND2_X1 U7039 ( .A1(n5998), .A2(n5997), .ZN(n7950) );
  OR2_X1 U7040 ( .A1(n6429), .A2(n7950), .ZN(n6001) );
  INV_X1 U7041 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5999) );
  OR2_X1 U7042 ( .A1(n8432), .A2(n5999), .ZN(n6000) );
  INV_X1 U7043 ( .A(n7866), .ZN(n9845) );
  NAND2_X1 U7044 ( .A1(n9845), .A2(n8422), .ZN(n6004) );
  NAND2_X1 U7045 ( .A1(n6005), .A2(n6004), .ZN(n6006) );
  XNOR2_X1 U7046 ( .A(n6006), .B(n5913), .ZN(n6009) );
  NOR2_X1 U7047 ( .A1(n6010), .A2(n6009), .ZN(n7942) );
  NAND2_X1 U7048 ( .A1(n7978), .A2(n8422), .ZN(n6008) );
  NAND2_X1 U7049 ( .A1(n9845), .A2(n5778), .ZN(n6007) );
  NAND2_X1 U7050 ( .A1(n6008), .A2(n6007), .ZN(n7944) );
  XOR2_X1 U7051 ( .A(n6012), .B(n6011), .Z(n8013) );
  MUX2_X1 U7052 ( .A(n6906), .B(n10442), .S(n5668), .Z(n6016) );
  NAND2_X1 U7053 ( .A1(n6016), .A2(n10467), .ZN(n6044) );
  INV_X1 U7054 ( .A(n6016), .ZN(n6017) );
  NAND2_X1 U7055 ( .A1(n6017), .A2(SI_12_), .ZN(n6018) );
  NAND2_X1 U7056 ( .A1(n6044), .A2(n6018), .ZN(n6042) );
  XNOR2_X1 U7057 ( .A(n6043), .B(n6042), .ZN(n7784) );
  NAND2_X1 U7058 ( .A1(n7784), .A2(n6176), .ZN(n6025) );
  NAND2_X1 U7059 ( .A1(n6019), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6069) );
  INV_X1 U7060 ( .A(n6069), .ZN(n6020) );
  NAND2_X1 U7061 ( .A1(n6020), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U7062 ( .A1(n6069), .A2(n6021), .ZN(n6049) );
  INV_X1 U7063 ( .A(n6643), .ZN(n7022) );
  OAI22_X1 U7064 ( .A1(n6199), .A2(n10442), .B1(n6473), .B2(n7022), .ZN(n6023)
         );
  INV_X1 U7065 ( .A(n6023), .ZN(n6024) );
  NAND2_X1 U7066 ( .A1(n10233), .A2(n8416), .ZN(n6034) );
  NAND2_X1 U7067 ( .A1(n5040), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6032) );
  INV_X1 U7068 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7968) );
  OR2_X1 U7069 ( .A1(n8430), .A2(n7968), .ZN(n6031) );
  INV_X1 U7070 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n6026) );
  OR2_X1 U7071 ( .A1(n8432), .A2(n6026), .ZN(n6030) );
  NAND2_X1 U7072 ( .A1(n6027), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6056) );
  OR2_X1 U7073 ( .A1(n6027), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U7074 ( .A1(n6056), .A2(n6028), .ZN(n8110) );
  OR2_X1 U7075 ( .A1(n6429), .A2(n8110), .ZN(n6029) );
  NAND2_X1 U7076 ( .A1(n9843), .A2(n8422), .ZN(n6033) );
  NAND2_X1 U7077 ( .A1(n6034), .A2(n6033), .ZN(n6035) );
  XNOR2_X1 U7078 ( .A(n6035), .B(n7288), .ZN(n6041) );
  INV_X1 U7079 ( .A(n6041), .ZN(n6039) );
  NAND2_X1 U7080 ( .A1(n10233), .A2(n8422), .ZN(n6037) );
  NAND2_X1 U7081 ( .A1(n9843), .A2(n5778), .ZN(n6036) );
  NAND2_X1 U7082 ( .A1(n6037), .A2(n6036), .ZN(n6040) );
  INV_X1 U7083 ( .A(n6040), .ZN(n6038) );
  NAND2_X1 U7084 ( .A1(n6039), .A2(n6038), .ZN(n8100) );
  AND2_X1 U7085 ( .A1(n6041), .A2(n6040), .ZN(n8101) );
  MUX2_X1 U7086 ( .A(n6958), .B(n10568), .S(n5668), .Z(n6046) );
  NAND2_X1 U7087 ( .A1(n6046), .A2(n10466), .ZN(n6065) );
  INV_X1 U7088 ( .A(n6046), .ZN(n6047) );
  NAND2_X1 U7089 ( .A1(n6047), .A2(SI_13_), .ZN(n6048) );
  NAND2_X1 U7090 ( .A1(n7991), .A2(n6176), .ZN(n6053) );
  NAND2_X1 U7091 ( .A1(n6049), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6050) );
  XNOR2_X1 U7092 ( .A(n6050), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6644) );
  INV_X1 U7093 ( .A(n6644), .ZN(n7085) );
  OAI22_X1 U7094 ( .A1(n6199), .A2(n10568), .B1(n5033), .B2(n7085), .ZN(n6051)
         );
  INV_X1 U7095 ( .A(n6051), .ZN(n6052) );
  NAND2_X1 U7096 ( .A1(n5040), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6061) );
  INV_X1 U7097 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n8121) );
  OR2_X1 U7098 ( .A1(n8430), .A2(n8121), .ZN(n6060) );
  INV_X1 U7099 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n6054) );
  OR2_X1 U7100 ( .A1(n8432), .A2(n6054), .ZN(n6059) );
  NAND2_X1 U7101 ( .A1(n6056), .A2(n6055), .ZN(n6057) );
  NAND2_X1 U7102 ( .A1(n6075), .A2(n6057), .ZN(n8144) );
  OR2_X1 U7103 ( .A1(n6429), .A2(n8144), .ZN(n6058) );
  OAI22_X1 U7104 ( .A1(n10983), .A2(n6300), .B1(n8106), .B2(n6208), .ZN(n6062)
         );
  XOR2_X1 U7105 ( .A(n7288), .B(n6062), .Z(n6063) );
  OAI22_X1 U7106 ( .A1(n10983), .A2(n6208), .B1(n8106), .B2(n8420), .ZN(n8136)
         );
  MUX2_X1 U7107 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n5668), .Z(n6085) );
  XNOR2_X1 U7108 ( .A(n6085), .B(SI_14_), .ZN(n6086) );
  INV_X1 U7109 ( .A(n6086), .ZN(n6066) );
  NAND2_X1 U7110 ( .A1(n8043), .A2(n6176), .ZN(n6074) );
  INV_X1 U7111 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10573) );
  OR2_X1 U7112 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n6067) );
  NAND2_X1 U7113 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n6067), .ZN(n6068) );
  NAND2_X1 U7114 ( .A1(n6069), .A2(n6068), .ZN(n6071) );
  XNOR2_X1 U7115 ( .A(n6071), .B(n6070), .ZN(n7144) );
  INV_X1 U7116 ( .A(n7144), .ZN(n6969) );
  OAI22_X1 U7117 ( .A1(n6199), .A2(n10573), .B1(n6969), .B2(n5033), .ZN(n6072)
         );
  INV_X1 U7118 ( .A(n6072), .ZN(n6073) );
  NAND2_X2 U7119 ( .A1(n6074), .A2(n6073), .ZN(n10228) );
  NAND2_X1 U7120 ( .A1(n5040), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6081) );
  INV_X1 U7121 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8091) );
  OR2_X1 U7122 ( .A1(n8430), .A2(n8091), .ZN(n6080) );
  AND2_X1 U7123 ( .A1(n6075), .A2(n7143), .ZN(n6076) );
  OR2_X1 U7124 ( .A1(n6076), .A2(n6098), .ZN(n9433) );
  OR2_X1 U7125 ( .A1(n6429), .A2(n9433), .ZN(n6079) );
  INV_X1 U7126 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n6077) );
  OR2_X1 U7127 ( .A1(n8432), .A2(n6077), .ZN(n6078) );
  AOI22_X1 U7128 ( .A1(n10228), .A2(n8422), .B1(n5778), .B2(n9841), .ZN(n9426)
         );
  INV_X1 U7129 ( .A(n6111), .ZN(n6109) );
  NAND2_X1 U7130 ( .A1(n10228), .A2(n8416), .ZN(n6083) );
  NAND2_X1 U7131 ( .A1(n9841), .A2(n8422), .ZN(n6082) );
  NAND2_X1 U7132 ( .A1(n6083), .A2(n6082), .ZN(n6084) );
  XNOR2_X1 U7133 ( .A(n6084), .B(n7288), .ZN(n6112) );
  INV_X1 U7134 ( .A(n6112), .ZN(n9427) );
  NOR2_X1 U7135 ( .A1(n9425), .A2(n9426), .ZN(n6113) );
  MUX2_X1 U7136 ( .A(n7048), .B(n10574), .S(n5668), .Z(n6087) );
  NAND2_X1 U7137 ( .A1(n6087), .A2(n10491), .ZN(n6114) );
  INV_X1 U7138 ( .A(n6087), .ZN(n6088) );
  NAND2_X1 U7139 ( .A1(n6088), .A2(SI_15_), .ZN(n6089) );
  NAND2_X1 U7140 ( .A1(n6114), .A2(n6089), .ZN(n6115) );
  XNOR2_X1 U7141 ( .A(n6116), .B(n6115), .ZN(n8154) );
  NAND2_X1 U7142 ( .A1(n8154), .A2(n6176), .ZN(n6097) );
  NOR2_X1 U7143 ( .A1(n6090), .A2(n10261), .ZN(n6091) );
  MUX2_X1 U7144 ( .A(n10261), .B(n6091), .S(P1_IR_REG_15__SCAN_IN), .Z(n6092)
         );
  INV_X1 U7145 ( .A(n6092), .ZN(n6094) );
  NAND2_X1 U7146 ( .A1(n6094), .A2(n6093), .ZN(n7730) );
  OAI22_X1 U7147 ( .A1(n6199), .A2(n10574), .B1(n6473), .B2(n7730), .ZN(n6095)
         );
  INV_X1 U7148 ( .A(n6095), .ZN(n6096) );
  NAND2_X1 U7149 ( .A1(n9567), .A2(n8416), .ZN(n6106) );
  NAND2_X1 U7150 ( .A1(n5040), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6104) );
  INV_X1 U7151 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8182) );
  OR2_X1 U7152 ( .A1(n8430), .A2(n8182), .ZN(n6103) );
  NOR2_X1 U7153 ( .A1(n6098), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6099) );
  OR2_X1 U7154 ( .A1(n6124), .A2(n6099), .ZN(n9563) );
  OR2_X1 U7155 ( .A1(n6429), .A2(n9563), .ZN(n6102) );
  INV_X1 U7156 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n6100) );
  OR2_X1 U7157 ( .A1(n8432), .A2(n6100), .ZN(n6101) );
  INV_X1 U7158 ( .A(n9429), .ZN(n10132) );
  NAND2_X1 U7159 ( .A1(n10132), .A2(n8422), .ZN(n6105) );
  NAND2_X1 U7160 ( .A1(n6106), .A2(n6105), .ZN(n6107) );
  XNOR2_X1 U7161 ( .A(n6107), .B(n7288), .ZN(n6110) );
  OAI21_X1 U7162 ( .B1(n6109), .B2(n9427), .A(n6108), .ZN(n9553) );
  INV_X1 U7163 ( .A(n9567), .ZN(n11008) );
  OAI22_X1 U7164 ( .A1(n11008), .A2(n6208), .B1(n9429), .B2(n8420), .ZN(n9556)
         );
  NAND2_X1 U7165 ( .A1(n9553), .A2(n9556), .ZN(n9485) );
  OAI211_X1 U7166 ( .C1(n6113), .C2(n6112), .A(n6111), .B(n6110), .ZN(n9554)
         );
  MUX2_X1 U7167 ( .A(n7054), .B(n10569), .S(n5668), .Z(n6118) );
  NAND2_X1 U7168 ( .A1(n6118), .A2(n6117), .ZN(n6143) );
  INV_X1 U7169 ( .A(n6118), .ZN(n6119) );
  NAND2_X1 U7170 ( .A1(n6119), .A2(SI_16_), .ZN(n6120) );
  XNOR2_X1 U7171 ( .A(n6142), .B(n6141), .ZN(n8208) );
  NAND2_X1 U7172 ( .A1(n8208), .A2(n6176), .ZN(n6123) );
  NAND2_X1 U7173 ( .A1(n6093), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6146) );
  XNOR2_X1 U7174 ( .A(n6146), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9860) );
  INV_X1 U7175 ( .A(n9860), .ZN(n7743) );
  OAI22_X1 U7176 ( .A1(n6199), .A2(n10569), .B1(n6473), .B2(n7743), .ZN(n6121)
         );
  INV_X1 U7177 ( .A(n6121), .ZN(n6122) );
  NAND2_X1 U7178 ( .A1(n10223), .A2(n8416), .ZN(n6133) );
  NAND2_X1 U7179 ( .A1(n5040), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6131) );
  OR2_X1 U7180 ( .A1(n6124), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6125) );
  AND2_X1 U7181 ( .A1(n6155), .A2(n6125), .ZN(n10140) );
  NAND2_X1 U7182 ( .A1(n5855), .A2(n10140), .ZN(n6130) );
  INV_X1 U7183 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n6126) );
  OR2_X1 U7184 ( .A1(n8430), .A2(n6126), .ZN(n6129) );
  INV_X1 U7185 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n6127) );
  OR2_X1 U7186 ( .A1(n8432), .A2(n6127), .ZN(n6128) );
  NAND4_X1 U7187 ( .A1(n6131), .A2(n6130), .A3(n6129), .A4(n6128), .ZN(n10109)
         );
  NAND2_X1 U7188 ( .A1(n10109), .A2(n8422), .ZN(n6132) );
  NAND2_X1 U7189 ( .A1(n6133), .A2(n6132), .ZN(n6134) );
  XNOR2_X1 U7190 ( .A(n6134), .B(n5913), .ZN(n6136) );
  AND2_X1 U7191 ( .A1(n10109), .A2(n5778), .ZN(n6135) );
  AOI21_X1 U7192 ( .B1(n10223), .B2(n8422), .A(n6135), .ZN(n6137) );
  NAND2_X1 U7193 ( .A1(n6136), .A2(n6137), .ZN(n9494) );
  INV_X1 U7194 ( .A(n6136), .ZN(n6139) );
  INV_X1 U7195 ( .A(n6137), .ZN(n6138) );
  NAND2_X1 U7196 ( .A1(n6139), .A2(n6138), .ZN(n6140) );
  AND2_X1 U7197 ( .A1(n9494), .A2(n6140), .ZN(n9484) );
  NAND3_X1 U7198 ( .A1(n9485), .A2(n9554), .A3(n9484), .ZN(n9483) );
  NAND2_X1 U7199 ( .A1(n6142), .A2(n6141), .ZN(n6144) );
  MUX2_X1 U7200 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n5668), .Z(n6171) );
  XNOR2_X1 U7201 ( .A(n6171), .B(SI_17_), .ZN(n6173) );
  INV_X1 U7202 ( .A(n6173), .ZN(n6145) );
  XNOR2_X1 U7203 ( .A(n6174), .B(n6145), .ZN(n8213) );
  NAND2_X1 U7204 ( .A1(n8213), .A2(n6176), .ZN(n6151) );
  NAND2_X1 U7205 ( .A1(n6146), .A2(n10619), .ZN(n6147) );
  NAND2_X1 U7206 ( .A1(n6147), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7207 ( .A1(n6148), .A2(n10415), .ZN(n6177) );
  OR2_X1 U7208 ( .A1(n6148), .A2(n10415), .ZN(n6149) );
  AOI22_X1 U7209 ( .A1(n9574), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5814), .B2(
        n9875), .ZN(n6150) );
  NAND2_X1 U7210 ( .A1(n10216), .A2(n8416), .ZN(n6161) );
  INV_X1 U7211 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7212 ( .A1(n5768), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6152) );
  OAI21_X1 U7213 ( .B1(n6153), .B2(n8462), .A(n6152), .ZN(n6159) );
  NAND2_X1 U7214 ( .A1(n6155), .A2(n6154), .ZN(n6156) );
  NAND2_X1 U7215 ( .A1(n6183), .A2(n6156), .ZN(n9497) );
  NAND2_X1 U7216 ( .A1(n8458), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6157) );
  OAI21_X1 U7217 ( .B1(n9497), .B2(n6429), .A(n6157), .ZN(n6158) );
  NAND2_X1 U7218 ( .A1(n10129), .A2(n8422), .ZN(n6160) );
  NAND2_X1 U7219 ( .A1(n6161), .A2(n6160), .ZN(n6162) );
  XNOR2_X1 U7220 ( .A(n6162), .B(n5913), .ZN(n6164) );
  AND2_X1 U7221 ( .A1(n10129), .A2(n5778), .ZN(n6163) );
  AOI21_X1 U7222 ( .B1(n10216), .B2(n8422), .A(n6163), .ZN(n6165) );
  NAND2_X1 U7223 ( .A1(n6164), .A2(n6165), .ZN(n6169) );
  INV_X1 U7224 ( .A(n6164), .ZN(n6167) );
  INV_X1 U7225 ( .A(n6165), .ZN(n6166) );
  NAND2_X1 U7226 ( .A1(n6167), .A2(n6166), .ZN(n6168) );
  NAND2_X1 U7227 ( .A1(n6169), .A2(n6168), .ZN(n9493) );
  INV_X1 U7228 ( .A(n6169), .ZN(n6170) );
  NAND2_X1 U7229 ( .A1(n6171), .A2(SI_17_), .ZN(n6172) );
  MUX2_X1 U7230 ( .A(n6175), .B(n10571), .S(n5668), .Z(n6191) );
  XNOR2_X1 U7231 ( .A(n6190), .B(n5113), .ZN(n8222) );
  NAND2_X1 U7232 ( .A1(n8222), .A2(n6176), .ZN(n6181) );
  NAND2_X1 U7233 ( .A1(n6177), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6178) );
  XNOR2_X1 U7234 ( .A(n6178), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9891) );
  INV_X1 U7235 ( .A(n9891), .ZN(n9873) );
  OAI22_X1 U7236 ( .A1(n6199), .A2(n10571), .B1(n6473), .B2(n9873), .ZN(n6179)
         );
  INV_X1 U7237 ( .A(n6179), .ZN(n6180) );
  AND2_X1 U7238 ( .A1(n6183), .A2(n6182), .ZN(n6184) );
  OR2_X1 U7239 ( .A1(n6184), .A2(n6203), .ZN(n10091) );
  AOI22_X1 U7240 ( .A1(n5040), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n5768), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n6186) );
  NAND2_X1 U7241 ( .A1(n8458), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6185) );
  OAI211_X1 U7242 ( .C1(n10091), .C2(n6429), .A(n6186), .B(n6185), .ZN(n10110)
         );
  INV_X1 U7243 ( .A(n10110), .ZN(n9499) );
  OAI22_X1 U7244 ( .A1(n10208), .A2(n6300), .B1(n9499), .B2(n6208), .ZN(n6187)
         );
  XNOR2_X1 U7245 ( .A(n6187), .B(n7288), .ZN(n6188) );
  AOI22_X1 U7246 ( .A1(n10096), .A2(n8422), .B1(n5778), .B2(n10110), .ZN(n9537) );
  NAND2_X1 U7247 ( .A1(n6189), .A2(n6188), .ZN(n9536) );
  INV_X1 U7248 ( .A(n6191), .ZN(n6192) );
  MUX2_X1 U7249 ( .A(n8495), .B(n10563), .S(n5668), .Z(n6193) );
  INV_X1 U7250 ( .A(SI_19_), .ZN(n10489) );
  NAND2_X1 U7251 ( .A1(n6193), .A2(n10489), .ZN(n6215) );
  INV_X1 U7252 ( .A(n6193), .ZN(n6194) );
  NAND2_X1 U7253 ( .A1(n6194), .A2(SI_19_), .ZN(n6195) );
  NAND2_X1 U7254 ( .A1(n6215), .A2(n6195), .ZN(n6196) );
  NAND2_X1 U7255 ( .A1(n6197), .A2(n6196), .ZN(n6198) );
  NAND2_X1 U7256 ( .A1(n6216), .A2(n6198), .ZN(n10661) );
  NAND2_X1 U7257 ( .A1(n10661), .A2(n6176), .ZN(n6202) );
  OAI22_X1 U7258 ( .A1(n6199), .A2(n10563), .B1(n10030), .B2(n5033), .ZN(n6200) );
  INV_X1 U7259 ( .A(n6200), .ZN(n6201) );
  NAND2_X1 U7260 ( .A1(n10203), .A2(n8416), .ZN(n6210) );
  NAND2_X1 U7261 ( .A1(n6203), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6222) );
  OR2_X1 U7262 ( .A1(n6203), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6204) );
  AND2_X1 U7263 ( .A1(n6222), .A2(n6204), .ZN(n10062) );
  NAND2_X1 U7264 ( .A1(n10062), .A2(n5855), .ZN(n6207) );
  AOI22_X1 U7265 ( .A1(n5040), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n5768), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7266 ( .A1(n8458), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6205) );
  OR2_X1 U7267 ( .A1(n10084), .A2(n6208), .ZN(n6209) );
  NAND2_X1 U7268 ( .A1(n6210), .A2(n6209), .ZN(n6211) );
  XNOR2_X1 U7269 ( .A(n6211), .B(n5913), .ZN(n6214) );
  NOR2_X1 U7270 ( .A1(n10084), .A2(n8420), .ZN(n6212) );
  AOI21_X1 U7271 ( .B1(n10203), .B2(n8422), .A(n6212), .ZN(n6213) );
  NOR2_X1 U7272 ( .A1(n6214), .A2(n6213), .ZN(n9447) );
  NAND2_X1 U7273 ( .A1(n6214), .A2(n6213), .ZN(n9446) );
  MUX2_X1 U7274 ( .A(n8246), .B(n10562), .S(n5668), .Z(n6217) );
  NAND2_X1 U7275 ( .A1(n6217), .A2(n10485), .ZN(n6236) );
  INV_X1 U7276 ( .A(n6217), .ZN(n6218) );
  NAND2_X1 U7277 ( .A1(n6218), .A2(SI_20_), .ZN(n6219) );
  XNOR2_X1 U7278 ( .A(n6235), .B(n6234), .ZN(n8245) );
  NAND2_X1 U7279 ( .A1(n8245), .A2(n6176), .ZN(n6221) );
  NAND2_X1 U7280 ( .A1(n9574), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7281 ( .A1(n6222), .A2(n9516), .ZN(n6223) );
  NAND2_X1 U7282 ( .A1(n6241), .A2(n6223), .ZN(n10051) );
  OR2_X1 U7283 ( .A1(n10051), .A2(n6429), .ZN(n6229) );
  INV_X1 U7284 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U7285 ( .A1(n5768), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U7286 ( .A1(n8458), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6224) );
  OAI211_X1 U7287 ( .C1(n6226), .C2(n8462), .A(n6225), .B(n6224), .ZN(n6227)
         );
  INV_X1 U7288 ( .A(n6227), .ZN(n6228) );
  OAI22_X1 U7289 ( .A1(n10054), .A2(n6300), .B1(n9451), .B2(n6208), .ZN(n6230)
         );
  XOR2_X1 U7290 ( .A(n7288), .B(n6230), .Z(n9513) );
  INV_X1 U7291 ( .A(n9513), .ZN(n6231) );
  OAI22_X1 U7292 ( .A1(n10054), .A2(n6208), .B1(n9451), .B2(n8420), .ZN(n6232)
         );
  NOR2_X1 U7293 ( .A1(n6231), .A2(n6232), .ZN(n6233) );
  INV_X1 U7294 ( .A(n6232), .ZN(n9512) );
  MUX2_X1 U7295 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n5668), .Z(n6256) );
  XNOR2_X1 U7296 ( .A(n6256), .B(n10484), .ZN(n6255) );
  XNOR2_X1 U7297 ( .A(n6259), .B(n6255), .ZN(n8203) );
  NAND2_X1 U7298 ( .A1(n8203), .A2(n6176), .ZN(n6239) );
  NAND2_X1 U7299 ( .A1(n9574), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U7300 ( .A1(n10194), .A2(n8416), .ZN(n6250) );
  INV_X1 U7301 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U7302 ( .A1(n6241), .A2(n6240), .ZN(n6242) );
  AND2_X1 U7303 ( .A1(n6269), .A2(n6242), .ZN(n10029) );
  NAND2_X1 U7304 ( .A1(n10029), .A2(n5855), .ZN(n6248) );
  INV_X1 U7305 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7306 ( .A1(n5768), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U7307 ( .A1(n8458), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6243) );
  OAI211_X1 U7308 ( .C1(n8462), .C2(n6245), .A(n6244), .B(n6243), .ZN(n6246)
         );
  INV_X1 U7309 ( .A(n6246), .ZN(n6247) );
  NAND2_X1 U7310 ( .A1(n10016), .A2(n8422), .ZN(n6249) );
  NAND2_X1 U7311 ( .A1(n6250), .A2(n6249), .ZN(n6251) );
  XNOR2_X1 U7312 ( .A(n6251), .B(n5913), .ZN(n6254) );
  NOR2_X1 U7313 ( .A1(n10038), .A2(n8420), .ZN(n6252) );
  AOI21_X1 U7314 ( .B1(n10194), .B2(n8422), .A(n6252), .ZN(n6253) );
  NOR2_X1 U7315 ( .A1(n6254), .A2(n6253), .ZN(n9465) );
  INV_X1 U7316 ( .A(n6255), .ZN(n6258) );
  INV_X1 U7317 ( .A(n6256), .ZN(n6257) );
  MUX2_X1 U7318 ( .A(n8261), .B(n7709), .S(n5668), .Z(n6261) );
  NAND2_X1 U7319 ( .A1(n6261), .A2(n6260), .ZN(n6281) );
  INV_X1 U7320 ( .A(n6261), .ZN(n6262) );
  NAND2_X1 U7321 ( .A1(n6262), .A2(SI_22_), .ZN(n6263) );
  NAND2_X1 U7322 ( .A1(n6281), .A2(n6263), .ZN(n6264) );
  NAND2_X1 U7323 ( .A1(n6265), .A2(n6264), .ZN(n6266) );
  NAND2_X1 U7324 ( .A1(n6282), .A2(n6266), .ZN(n8260) );
  NAND2_X1 U7325 ( .A1(n8260), .A2(n6176), .ZN(n6268) );
  NAND2_X1 U7326 ( .A1(n9574), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6267) );
  INV_X1 U7327 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9528) );
  AND2_X1 U7328 ( .A1(n6269), .A2(n9528), .ZN(n6270) );
  OR2_X1 U7329 ( .A1(n6270), .A2(n6292), .ZN(n9527) );
  INV_X1 U7330 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U7331 ( .A1(n5768), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U7332 ( .A1(n8458), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6271) );
  OAI211_X1 U7333 ( .C1(n6273), .C2(n8462), .A(n6272), .B(n6271), .ZN(n6274)
         );
  AOI21_X1 U7334 ( .B1(n10010), .B2(n5855), .A(n6274), .ZN(n9470) );
  OAI22_X1 U7335 ( .A1(n10012), .A2(n6208), .B1(n9470), .B2(n8420), .ZN(n6277)
         );
  OAI22_X1 U7336 ( .A1(n10012), .A2(n6300), .B1(n9470), .B2(n6208), .ZN(n6275)
         );
  XNOR2_X1 U7337 ( .A(n6275), .B(n7288), .ZN(n6276) );
  XOR2_X1 U7338 ( .A(n6277), .B(n6276), .Z(n9524) );
  INV_X1 U7339 ( .A(n6276), .ZN(n6279) );
  INV_X1 U7340 ( .A(n6277), .ZN(n6278) );
  INV_X1 U7341 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n6283) );
  MUX2_X1 U7342 ( .A(n8271), .B(n6283), .S(n5668), .Z(n6284) );
  NAND2_X1 U7343 ( .A1(n6284), .A2(n10473), .ZN(n6302) );
  INV_X1 U7344 ( .A(n6284), .ZN(n6285) );
  NAND2_X1 U7345 ( .A1(n6285), .A2(SI_23_), .ZN(n6286) );
  OR2_X1 U7346 ( .A1(n6288), .A2(n6287), .ZN(n6289) );
  NAND2_X1 U7347 ( .A1(n6303), .A2(n6289), .ZN(n8270) );
  NAND2_X1 U7348 ( .A1(n8270), .A2(n6176), .ZN(n6291) );
  NAND2_X1 U7349 ( .A1(n9574), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6290) );
  NOR2_X1 U7350 ( .A1(n6292), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6293) );
  NOR2_X1 U7351 ( .A1(n6306), .A2(n6293), .ZN(n9996) );
  NAND2_X1 U7352 ( .A1(n9996), .A2(n5855), .ZN(n6299) );
  INV_X1 U7353 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U7354 ( .A1(n5768), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U7355 ( .A1(n8458), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6294) );
  OAI211_X1 U7356 ( .C1(n8462), .C2(n6296), .A(n6295), .B(n6294), .ZN(n6297)
         );
  INV_X1 U7357 ( .A(n6297), .ZN(n6298) );
  OAI22_X1 U7358 ( .A1(n9998), .A2(n6300), .B1(n9508), .B2(n6208), .ZN(n6301)
         );
  XOR2_X1 U7359 ( .A(n7288), .B(n6301), .Z(n9439) );
  AOI22_X1 U7360 ( .A1(n10184), .A2(n8422), .B1(n5778), .B2(n10015), .ZN(n9438) );
  MUX2_X1 U7361 ( .A(n8276), .B(n10555), .S(n5668), .Z(n6321) );
  XNOR2_X1 U7362 ( .A(n6321), .B(SI_24_), .ZN(n6320) );
  XNOR2_X1 U7363 ( .A(n6325), .B(n6320), .ZN(n8275) );
  NAND2_X1 U7364 ( .A1(n8275), .A2(n6176), .ZN(n6305) );
  NAND2_X1 U7365 ( .A1(n9574), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6304) );
  NAND2_X1 U7366 ( .A1(n10179), .A2(n8416), .ZN(n6315) );
  OR2_X1 U7367 ( .A1(n6306), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6307) );
  NAND2_X1 U7368 ( .A1(n6306), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6332) );
  AND2_X1 U7369 ( .A1(n6307), .A2(n6332), .ZN(n9987) );
  NAND2_X1 U7370 ( .A1(n9987), .A2(n5855), .ZN(n6313) );
  INV_X1 U7371 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U7372 ( .A1(n5768), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6309) );
  NAND2_X1 U7373 ( .A1(n8458), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6308) );
  OAI211_X1 U7374 ( .C1(n6310), .C2(n8462), .A(n6309), .B(n6308), .ZN(n6311)
         );
  INV_X1 U7375 ( .A(n6311), .ZN(n6312) );
  NAND2_X1 U7376 ( .A1(n10002), .A2(n8422), .ZN(n6314) );
  NAND2_X1 U7377 ( .A1(n6315), .A2(n6314), .ZN(n6316) );
  XNOR2_X1 U7378 ( .A(n6316), .B(n7288), .ZN(n6317) );
  AOI22_X1 U7379 ( .A1(n10179), .A2(n8422), .B1(n5778), .B2(n10002), .ZN(n6318) );
  XNOR2_X1 U7380 ( .A(n6317), .B(n6318), .ZN(n9504) );
  INV_X1 U7381 ( .A(n6317), .ZN(n6319) );
  INV_X1 U7382 ( .A(n6320), .ZN(n6324) );
  INV_X1 U7383 ( .A(n6321), .ZN(n6322) );
  NAND2_X1 U7384 ( .A1(n6322), .A2(SI_24_), .ZN(n6323) );
  INV_X1 U7385 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8291) );
  MUX2_X1 U7386 ( .A(n8291), .B(n10443), .S(n5668), .Z(n6326) );
  NAND2_X1 U7387 ( .A1(n6326), .A2(n10311), .ZN(n6345) );
  INV_X1 U7388 ( .A(n6326), .ZN(n6327) );
  NAND2_X1 U7389 ( .A1(n6327), .A2(SI_25_), .ZN(n6328) );
  NAND2_X1 U7390 ( .A1(n6345), .A2(n6328), .ZN(n6346) );
  XNOR2_X1 U7391 ( .A(n6347), .B(n6346), .ZN(n8290) );
  NAND2_X1 U7392 ( .A1(n8290), .A2(n6176), .ZN(n6330) );
  NAND2_X1 U7393 ( .A1(n9574), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6329) );
  NAND2_X1 U7394 ( .A1(n10175), .A2(n8416), .ZN(n6339) );
  NAND2_X1 U7395 ( .A1(n5040), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6337) );
  INV_X1 U7396 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9966) );
  OR2_X1 U7397 ( .A1(n8430), .A2(n9966), .ZN(n6336) );
  INV_X1 U7398 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n6331) );
  OR2_X1 U7399 ( .A1(n8432), .A2(n6331), .ZN(n6335) );
  NAND2_X1 U7400 ( .A1(n6333), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6353) );
  OAI21_X1 U7401 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n6333), .A(n6353), .ZN(
        n9965) );
  OR2_X1 U7402 ( .A1(n6429), .A2(n9965), .ZN(n6334) );
  NAND2_X1 U7403 ( .A1(n9982), .A2(n8422), .ZN(n6338) );
  NAND2_X1 U7404 ( .A1(n6339), .A2(n6338), .ZN(n6340) );
  XNOR2_X1 U7405 ( .A(n6340), .B(n7288), .ZN(n9474) );
  NAND2_X1 U7406 ( .A1(n10175), .A2(n8422), .ZN(n6342) );
  NAND2_X1 U7407 ( .A1(n9982), .A2(n5778), .ZN(n6341) );
  NAND2_X1 U7408 ( .A1(n6342), .A2(n6341), .ZN(n9475) );
  NAND2_X1 U7409 ( .A1(n9474), .A2(n9475), .ZN(n6344) );
  INV_X1 U7410 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8301) );
  MUX2_X1 U7411 ( .A(n8301), .B(n10445), .S(n5668), .Z(n6348) );
  NAND2_X1 U7412 ( .A1(n6348), .A2(n10309), .ZN(n6367) );
  INV_X1 U7413 ( .A(n6348), .ZN(n6349) );
  NAND2_X1 U7414 ( .A1(n6349), .A2(SI_26_), .ZN(n6350) );
  XNOR2_X1 U7415 ( .A(n6366), .B(n6365), .ZN(n8300) );
  NAND2_X1 U7416 ( .A1(n8300), .A2(n6176), .ZN(n6352) );
  NAND2_X1 U7417 ( .A1(n9574), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6351) );
  INV_X1 U7418 ( .A(n10168), .ZN(n9950) );
  INV_X1 U7419 ( .A(n6353), .ZN(n6354) );
  NAND2_X1 U7420 ( .A1(n6354), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6372) );
  OAI21_X1 U7421 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n6354), .A(n6372), .ZN(
        n9947) );
  OR2_X1 U7422 ( .A1(n6429), .A2(n9947), .ZN(n6359) );
  NAND2_X1 U7423 ( .A1(n5768), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U7424 ( .A1(n5040), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6357) );
  INV_X1 U7425 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n6355) );
  OR2_X1 U7426 ( .A1(n8432), .A2(n6355), .ZN(n6356) );
  NAND4_X1 U7427 ( .A1(n6359), .A2(n6358), .A3(n6357), .A4(n6356), .ZN(n9940)
         );
  OAI22_X1 U7428 ( .A1(n9950), .A2(n6208), .B1(n9973), .B2(n8420), .ZN(n6363)
         );
  NAND2_X1 U7429 ( .A1(n10168), .A2(n8416), .ZN(n6361) );
  NAND2_X1 U7430 ( .A1(n9940), .A2(n8422), .ZN(n6360) );
  NAND2_X1 U7431 ( .A1(n6361), .A2(n6360), .ZN(n6362) );
  XNOR2_X1 U7432 ( .A(n6362), .B(n7288), .ZN(n6364) );
  XOR2_X1 U7433 ( .A(n6363), .B(n6364), .Z(n9545) );
  NAND2_X1 U7434 ( .A1(n6366), .A2(n6365), .ZN(n6368) );
  MUX2_X1 U7435 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n5668), .Z(n8190) );
  XNOR2_X1 U7436 ( .A(n8190), .B(n10474), .ZN(n8189) );
  NAND2_X1 U7437 ( .A1(n8315), .A2(n6176), .ZN(n6370) );
  NAND2_X1 U7438 ( .A1(n9574), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6369) );
  NAND2_X1 U7439 ( .A1(n10163), .A2(n8416), .ZN(n6379) );
  NAND2_X1 U7440 ( .A1(n5040), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6377) );
  INV_X1 U7441 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6371) );
  OR2_X1 U7442 ( .A1(n8430), .A2(n6371), .ZN(n6376) );
  XNOR2_X1 U7443 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n6424), .ZN(n6415) );
  OR2_X1 U7444 ( .A1(n6429), .A2(n6415), .ZN(n6375) );
  INV_X1 U7445 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n6373) );
  OR2_X1 U7446 ( .A1(n8432), .A2(n6373), .ZN(n6374) );
  NAND2_X1 U7447 ( .A1(n9953), .A2(n8422), .ZN(n6378) );
  NAND2_X1 U7448 ( .A1(n6379), .A2(n6378), .ZN(n6380) );
  XNOR2_X1 U7449 ( .A(n6380), .B(n5913), .ZN(n6383) );
  NOR2_X1 U7450 ( .A1(n9547), .A2(n8420), .ZN(n6381) );
  AOI21_X1 U7451 ( .B1(n10163), .B2(n8422), .A(n6381), .ZN(n6382) );
  NAND2_X1 U7452 ( .A1(n6383), .A2(n6382), .ZN(n8439) );
  OAI21_X1 U7453 ( .B1(n6383), .B2(n6382), .A(n8439), .ZN(n6384) );
  NAND2_X1 U7454 ( .A1(n8445), .A2(n6386), .ZN(n6412) );
  NAND2_X1 U7455 ( .A1(n5765), .A2(n5762), .ZN(n7293) );
  INV_X1 U7456 ( .A(n7293), .ZN(n6893) );
  INV_X1 U7457 ( .A(n6387), .ZN(n7265) );
  OR2_X1 U7458 ( .A1(n10946), .A2(n7265), .ZN(n6416) );
  INV_X1 U7459 ( .A(n6388), .ZN(n6389) );
  NAND2_X1 U7460 ( .A1(n6389), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6390) );
  MUX2_X1 U7461 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6390), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n6391) );
  NAND2_X1 U7462 ( .A1(n6391), .A2(n5730), .ZN(n7852) );
  AND2_X1 U7463 ( .A1(n7852), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6392) );
  NOR2_X1 U7464 ( .A1(n6416), .A2(n10666), .ZN(n6411) );
  NAND2_X1 U7465 ( .A1(n8130), .A2(P1_B_REG_SCAN_IN), .ZN(n6394) );
  INV_X1 U7466 ( .A(n7976), .ZN(n6393) );
  MUX2_X1 U7467 ( .A(n6394), .B(P1_B_REG_SCAN_IN), .S(n6393), .Z(n6396) );
  NAND2_X1 U7468 ( .A1(n6396), .A2(n6395), .ZN(n6406) );
  INV_X1 U7469 ( .A(n6395), .ZN(n8135) );
  NAND2_X1 U7470 ( .A1(n8135), .A2(n8130), .ZN(n6397) );
  OAI21_X1 U7471 ( .B1(n6406), .B2(P1_D_REG_1__SCAN_IN), .A(n6397), .ZN(n6895)
         );
  INV_X1 U7472 ( .A(n6895), .ZN(n10258) );
  NOR4_X1 U7473 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n6401) );
  NOR4_X1 U7474 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6400) );
  NOR4_X1 U7475 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6399) );
  NOR4_X1 U7476 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6398) );
  NAND4_X1 U7477 ( .A1(n6401), .A2(n6400), .A3(n6399), .A4(n6398), .ZN(n6408)
         );
  NOR2_X1 U7478 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n6405) );
  NOR4_X1 U7479 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_31__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n6404) );
  NOR4_X1 U7480 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n6403) );
  NOR4_X1 U7481 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n6402) );
  NAND4_X1 U7482 ( .A1(n6405), .A2(n6404), .A3(n6403), .A4(n6402), .ZN(n6407)
         );
  OAI21_X1 U7483 ( .B1(n6408), .B2(n6407), .A(n10665), .ZN(n6894) );
  AND2_X1 U7484 ( .A1(n10258), .A2(n6894), .ZN(n7075) );
  INV_X1 U7485 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10646) );
  NAND2_X1 U7486 ( .A1(n10665), .A2(n10646), .ZN(n6410) );
  NAND2_X1 U7487 ( .A1(n8135), .A2(n7976), .ZN(n6409) );
  AND2_X1 U7488 ( .A1(n7075), .A2(n10259), .ZN(n6413) );
  NAND2_X1 U7489 ( .A1(n6412), .A2(n9525), .ZN(n6443) );
  OR3_X1 U7490 ( .A1(n10666), .A2(n7293), .A3(n9823), .ZN(n6421) );
  OR2_X1 U7491 ( .A1(n6938), .A2(n6421), .ZN(n6414) );
  INV_X1 U7492 ( .A(n6415), .ZN(n9932) );
  INV_X1 U7493 ( .A(n6416), .ZN(n6419) );
  OR2_X1 U7494 ( .A1(n6387), .A2(n6417), .ZN(n7073) );
  NAND3_X1 U7495 ( .A1(n7073), .A2(n6471), .A3(n7852), .ZN(n6418) );
  AOI21_X1 U7496 ( .B1(n6419), .B2(n6938), .A(n6418), .ZN(n6420) );
  OR2_X1 U7497 ( .A1(n6420), .A2(P1_U3084), .ZN(n6423) );
  OR2_X1 U7498 ( .A1(n6387), .A2(n9828), .ZN(n7287) );
  OR2_X1 U7499 ( .A1(n7287), .A2(n10666), .ZN(n9835) );
  NAND2_X1 U7500 ( .A1(n9835), .A2(n6421), .ZN(n6422) );
  NAND2_X1 U7501 ( .A1(n6938), .A2(n6422), .ZN(n6939) );
  NAND2_X1 U7502 ( .A1(n5040), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6434) );
  INV_X1 U7503 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9924) );
  OR2_X1 U7504 ( .A1(n8430), .A2(n9924), .ZN(n6433) );
  NAND2_X1 U7505 ( .A1(n6425), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8483) );
  INV_X1 U7506 ( .A(n6425), .ZN(n6427) );
  INV_X1 U7507 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6426) );
  NAND2_X1 U7508 ( .A1(n6427), .A2(n6426), .ZN(n6428) );
  NAND2_X1 U7509 ( .A1(n8483), .A2(n6428), .ZN(n9923) );
  INV_X1 U7510 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6430) );
  OR2_X1 U7511 ( .A1(n8432), .A2(n6430), .ZN(n6431) );
  NOR2_X1 U7512 ( .A1(n6938), .A2(n9835), .ZN(n6437) );
  INV_X1 U7513 ( .A(n6437), .ZN(n6436) );
  INV_X1 U7514 ( .A(n6979), .ZN(n9830) );
  AND2_X2 U7515 ( .A1(n6437), .A2(n9830), .ZN(n9561) );
  AOI22_X1 U7516 ( .A1(n9561), .A2(n9940), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n6438) );
  OAI21_X1 U7517 ( .B1(n9934), .B2(n9559), .A(n6438), .ZN(n6439) );
  AOI21_X1 U7518 ( .B1(n9932), .B2(n9505), .A(n6439), .ZN(n6440) );
  OAI21_X1 U7519 ( .B1(n5394), .B2(n9535), .A(n6440), .ZN(n6441) );
  INV_X1 U7520 ( .A(n6441), .ZN(n6442) );
  NAND2_X1 U7521 ( .A1(n6443), .A2(n6442), .ZN(P1_U3212) );
  INV_X1 U7522 ( .A(n7852), .ZN(n6444) );
  NOR2_X1 U7523 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n6452) );
  NOR2_X1 U7524 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6451) );
  NOR2_X1 U7525 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n6450) );
  NOR2_X1 U7526 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6449) );
  NAND2_X1 U7527 ( .A1(n5129), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6456) );
  MUX2_X1 U7528 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6456), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6458) );
  NAND2_X1 U7529 ( .A1(n6458), .A2(n6532), .ZN(n8133) );
  INV_X1 U7530 ( .A(n6467), .ZN(n6462) );
  NAND2_X1 U7531 ( .A1(n6468), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U7532 ( .A1(n6464), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6465) );
  MUX2_X1 U7533 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6465), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6466) );
  AND2_X1 U7534 ( .A1(n6466), .A2(n5129), .ZN(n6481) );
  NAND3_X1 U7535 ( .A1(n6477), .A2(n6478), .A3(n6481), .ZN(n6780) );
  NAND2_X1 U7536 ( .A1(n6467), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n6469) );
  NAND2_X1 U7537 ( .A1(n6469), .A2(n6468), .ZN(n6679) );
  INV_X1 U7538 ( .A(n10772), .ZN(n6470) );
  NAND2_X1 U7539 ( .A1(n6387), .A2(n6471), .ZN(n6472) );
  NAND2_X1 U7540 ( .A1(n6472), .A2(n7852), .ZN(n10742) );
  NAND2_X1 U7541 ( .A1(n10742), .A2(n5033), .ZN(n6474) );
  NAND2_X1 U7542 ( .A1(n6474), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U7543 ( .A(n6478), .ZN(n7974) );
  AOI22_X1 U7544 ( .A1(P2_B_REG_SCAN_IN), .A2(n7974), .B1(n6478), .B2(n10547), 
        .ZN(n6475) );
  OR2_X1 U7545 ( .A1(n6481), .A2(n6475), .ZN(n6476) );
  INV_X1 U7546 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10770) );
  NAND2_X1 U7547 ( .A1(n10700), .A2(n10770), .ZN(n6480) );
  NOR2_X1 U7548 ( .A1(n6478), .A2(n6477), .ZN(n10771) );
  INV_X1 U7549 ( .A(n10771), .ZN(n6479) );
  INV_X1 U7550 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10703) );
  NAND2_X1 U7551 ( .A1(n10700), .A2(n10703), .ZN(n6482) );
  INV_X1 U7552 ( .A(n6481), .ZN(n8131) );
  NAND2_X1 U7553 ( .A1(n8131), .A2(n8133), .ZN(n10699) );
  AND2_X1 U7554 ( .A1(n6482), .A2(n10699), .ZN(n7194) );
  NOR4_X1 U7555 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6486) );
  NOR4_X1 U7556 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6485) );
  NOR4_X1 U7557 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6484) );
  NOR4_X1 U7558 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6483) );
  NAND4_X1 U7559 ( .A1(n6486), .A2(n6485), .A3(n6484), .A4(n6483), .ZN(n6492)
         );
  NOR2_X1 U7560 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6490) );
  NOR4_X1 U7561 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6489) );
  NOR4_X1 U7562 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6488) );
  NOR4_X1 U7563 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6487) );
  NAND4_X1 U7564 ( .A1(n6490), .A2(n6489), .A3(n6488), .A4(n6487), .ZN(n6491)
         );
  OAI21_X1 U7565 ( .B1(n6492), .B2(n6491), .A(n10700), .ZN(n7235) );
  NAND2_X1 U7566 ( .A1(n7194), .A2(n7235), .ZN(n7203) );
  INV_X1 U7567 ( .A(n7203), .ZN(n6493) );
  NAND2_X1 U7568 ( .A1(n7231), .A2(n6493), .ZN(n6580) );
  INV_X1 U7569 ( .A(n10702), .ZN(n6494) );
  NAND2_X1 U7570 ( .A1(n6497), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6498) );
  INV_X1 U7571 ( .A(n7176), .ZN(n6777) );
  NAND2_X1 U7572 ( .A1(n6591), .A2(n6777), .ZN(n6514) );
  NAND3_X1 U7573 ( .A1(n6692), .A2(n6695), .A3(n6501), .ZN(n6502) );
  INV_X1 U7574 ( .A(n6503), .ZN(n6903) );
  NAND2_X1 U7575 ( .A1(n7406), .A2(n6506), .ZN(n6507) );
  INV_X1 U7576 ( .A(n10830), .ZN(n6590) );
  INV_X1 U7577 ( .A(n8922), .ZN(n8840) );
  NAND2_X1 U7578 ( .A1(n6516), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6517) );
  MUX2_X1 U7579 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6517), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n6518) );
  NAND2_X1 U7580 ( .A1(n7118), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6526) );
  INV_X1 U7581 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10451) );
  INV_X1 U7582 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6790) );
  INV_X1 U7583 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6522) );
  OR2_X1 U7584 ( .A1(n8253), .A2(n6522), .ZN(n6523) );
  NAND2_X1 U7585 ( .A1(n6579), .A2(n8796), .ZN(n6528) );
  NAND2_X1 U7586 ( .A1(n8811), .A2(n8820), .ZN(n6527) );
  NAND2_X4 U7587 ( .A1(n6528), .A2(n6527), .ZN(n8551) );
  XNOR2_X2 U7588 ( .A(n6531), .B(n6530), .ZN(n6582) );
  NAND2_X1 U7589 ( .A1(n6532), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6534) );
  NAND2_X4 U7590 ( .A1(n6582), .A2(n8375), .ZN(n7537) );
  INV_X1 U7591 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6668) );
  OR2_X1 U7592 ( .A1(n5038), .A2(n6668), .ZN(n6539) );
  OR2_X1 U7593 ( .A1(n5037), .A2(n6673), .ZN(n6538) );
  OR2_X1 U7594 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6564) );
  NAND2_X1 U7595 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n6564), .ZN(n6536) );
  OR2_X1 U7596 ( .A1(n7537), .A2(n6793), .ZN(n6537) );
  AND3_X2 U7597 ( .A1(n6539), .A2(n6538), .A3(n6537), .ZN(n10864) );
  XNOR2_X1 U7598 ( .A(n8563), .B(n10864), .ZN(n6559) );
  NAND3_X1 U7599 ( .A1(n8840), .A2(n8998), .A3(n6559), .ZN(n6577) );
  INV_X1 U7600 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10785) );
  INV_X1 U7601 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6792) );
  INV_X1 U7602 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6540) );
  OR2_X1 U7603 ( .A1(n8253), .A2(n6540), .ZN(n6541) );
  INV_X1 U7604 ( .A(n6545), .ZN(n6557) );
  INV_X1 U7605 ( .A(n6791), .ZN(n10791) );
  INV_X1 U7606 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6659) );
  XNOR2_X1 U7607 ( .A(n8551), .B(n7400), .ZN(n6556) );
  INV_X1 U7608 ( .A(SI_0_), .ZN(n10305) );
  INV_X1 U7609 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6546) );
  OAI21_X1 U7610 ( .B1(n5668), .B2(n10305), .A(n6546), .ZN(n6548) );
  AND2_X1 U7611 ( .A1(n6548), .A2(n6547), .ZN(n9424) );
  MUX2_X1 U7612 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9424), .S(n7537), .Z(n10831)
         );
  OR2_X1 U7613 ( .A1(n10831), .A2(n8551), .ZN(n7220) );
  NAND2_X1 U7614 ( .A1(n7118), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6552) );
  INV_X1 U7615 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10824) );
  INV_X1 U7616 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10775) );
  INV_X1 U7617 ( .A(n10831), .ZN(n10817) );
  OR2_X2 U7618 ( .A1(n7221), .A2(n10817), .ZN(n7398) );
  OAI21_X1 U7619 ( .B1(n6557), .B2(n6556), .A(n7219), .ZN(n7033) );
  AND2_X1 U7620 ( .A1(n8998), .A2(n8535), .ZN(n6558) );
  NAND2_X1 U7621 ( .A1(n6559), .A2(n6558), .ZN(n6572) );
  OAI21_X1 U7622 ( .B1(n6559), .B2(n6558), .A(n6572), .ZN(n7032) );
  NAND2_X1 U7623 ( .A1(n7118), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6563) );
  OR2_X1 U7624 ( .A1(n8321), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6562) );
  INV_X1 U7625 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6789) );
  OR2_X1 U7626 ( .A1(n8374), .A2(n6789), .ZN(n6561) );
  INV_X1 U7627 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7313) );
  OR2_X1 U7628 ( .A1(n8253), .A2(n7313), .ZN(n6560) );
  NOR2_X1 U7629 ( .A1(n7192), .A2(n8562), .ZN(n6568) );
  OAI21_X1 U7630 ( .B1(P2_IR_REG_2__SCAN_IN), .B2(n6564), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6565) );
  XNOR2_X1 U7631 ( .A(n6565), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6788) );
  INV_X1 U7632 ( .A(n6788), .ZN(n6837) );
  OR2_X1 U7633 ( .A1(n5037), .A2(n6665), .ZN(n6567) );
  XNOR2_X1 U7634 ( .A(n8551), .B(n7315), .ZN(n6569) );
  NAND2_X1 U7635 ( .A1(n6568), .A2(n6569), .ZN(n7099) );
  INV_X1 U7636 ( .A(n6568), .ZN(n6570) );
  INV_X1 U7637 ( .A(n6569), .ZN(n7359) );
  NAND2_X1 U7638 ( .A1(n6570), .A2(n7359), .ZN(n6571) );
  AND2_X1 U7639 ( .A1(n7099), .A2(n6571), .ZN(n6573) );
  OAI21_X1 U7640 ( .B1(n7031), .B2(n6573), .A(n8915), .ZN(n6576) );
  INV_X1 U7641 ( .A(n6572), .ZN(n6574) );
  INV_X1 U7642 ( .A(n7358), .ZN(n6575) );
  AOI21_X1 U7643 ( .B1(n6577), .B2(n6576), .A(n6575), .ZN(n6595) );
  NAND2_X1 U7644 ( .A1(n6780), .A2(n6679), .ZN(n6578) );
  NAND2_X1 U7645 ( .A1(n7234), .A2(n6580), .ZN(n7030) );
  NAND2_X1 U7646 ( .A1(n7029), .A2(n7030), .ZN(n6581) );
  MUX2_X1 U7647 ( .A(n8935), .B(P2_U3152), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n6594) );
  NAND2_X1 U7648 ( .A1(n7118), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6587) );
  NAND2_X1 U7649 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n7110) );
  OAI21_X1 U7650 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n7110), .ZN(n7368) );
  OR2_X1 U7651 ( .A1(n8321), .A2(n7368), .ZN(n6586) );
  INV_X1 U7652 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6794) );
  OR2_X1 U7653 ( .A1(n8374), .A2(n6794), .ZN(n6585) );
  INV_X1 U7654 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6583) );
  OR2_X1 U7655 ( .A1(n8253), .A2(n6583), .ZN(n6584) );
  NAND4_X1 U7656 ( .A1(n6587), .A2(n6586), .A3(n6585), .A4(n6584), .ZN(n8996)
         );
  AOI22_X1 U7657 ( .A1(n10821), .A2(n8996), .B1(n8998), .B2(n9254), .ZN(n7307)
         );
  INV_X1 U7658 ( .A(n8819), .ZN(n6588) );
  NAND2_X1 U7659 ( .A1(n6591), .A2(n6588), .ZN(n7845) );
  NOR2_X1 U7660 ( .A1(n8801), .A2(n6590), .ZN(n7205) );
  NAND2_X1 U7661 ( .A1(n6591), .A2(n7205), .ZN(n6592) );
  OAI22_X1 U7662 ( .A1(n7307), .A2(n7845), .B1(n8963), .B2(n10877), .ZN(n6593)
         );
  OR3_X1 U7663 ( .A1(n6595), .A2(n6594), .A3(n6593), .ZN(P2_U3220) );
  AOI22_X1 U7664 ( .A1(n6969), .A2(n8091), .B1(P1_REG2_REG_14__SCAN_IN), .B2(
        n7144), .ZN(n7138) );
  NAND2_X1 U7665 ( .A1(n6771), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6610) );
  MUX2_X1 U7666 ( .A(n5975), .B(P1_REG2_REG_9__SCAN_IN), .S(n6771), .Z(n6596)
         );
  INV_X1 U7667 ( .A(n6596), .ZN(n6766) );
  NOR2_X1 U7668 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n6675), .ZN(n6609) );
  INV_X1 U7669 ( .A(n6872), .ZN(n6631) );
  NOR2_X1 U7670 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6711), .ZN(n6607) );
  INV_X1 U7671 ( .A(n6626), .ZN(n6985) );
  NAND2_X1 U7672 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(n6858), .ZN(n6603) );
  INV_X1 U7673 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6597) );
  MUX2_X1 U7674 ( .A(n6597), .B(P1_REG2_REG_3__SCAN_IN), .S(n6858), .Z(n6598)
         );
  INV_X1 U7675 ( .A(n6598), .ZN(n6860) );
  NAND2_X1 U7676 ( .A1(n6672), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6602) );
  MUX2_X1 U7677 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6599), .S(n6672), .Z(n6999)
         );
  NAND2_X1 U7678 ( .A1(P1_REG2_REG_1__SCAN_IN), .A2(n10759), .ZN(n6601) );
  INV_X1 U7679 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6600) );
  MUX2_X1 U7680 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6600), .S(n10759), .Z(n10764) );
  NAND3_X1 U7681 ( .A1(n10753), .A2(P1_REG2_REG_0__SCAN_IN), .A3(n10764), .ZN(
        n10762) );
  NAND2_X1 U7682 ( .A1(n6601), .A2(n10762), .ZN(n7000) );
  NAND2_X1 U7683 ( .A1(n6999), .A2(n7000), .ZN(n6998) );
  NAND2_X1 U7684 ( .A1(n6602), .A2(n6998), .ZN(n6861) );
  NAND2_X1 U7685 ( .A1(n6860), .A2(n6861), .ZN(n6859) );
  NAND2_X1 U7686 ( .A1(n6603), .A2(n6859), .ZN(n6988) );
  MUX2_X1 U7687 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6605), .S(n6626), .Z(n6604)
         );
  INV_X1 U7688 ( .A(n6604), .ZN(n6987) );
  NOR2_X1 U7689 ( .A1(n6988), .A2(n6987), .ZN(n6986) );
  AOI21_X1 U7690 ( .B1(n6985), .B2(n6605), .A(n6986), .ZN(n6704) );
  MUX2_X1 U7691 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7478), .S(n6711), .Z(n6606)
         );
  INV_X1 U7692 ( .A(n6606), .ZN(n6705) );
  NOR2_X1 U7693 ( .A1(n6704), .A2(n6705), .ZN(n6703) );
  OR2_X1 U7694 ( .A1(n6607), .A2(n6703), .ZN(n6875) );
  MUX2_X1 U7695 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7513), .S(n6872), .Z(n6874)
         );
  NOR2_X1 U7696 ( .A1(n6875), .A2(n6874), .ZN(n6873) );
  AOI21_X1 U7697 ( .B1(n6631), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6873), .ZN(
        n6737) );
  MUX2_X1 U7698 ( .A(n7603), .B(P1_REG2_REG_7__SCAN_IN), .S(n6740), .Z(n6736)
         );
  AND2_X1 U7699 ( .A1(n6737), .A2(n6736), .ZN(n6738) );
  AOI21_X1 U7700 ( .B1(n7603), .B2(n6740), .A(n6738), .ZN(n6760) );
  MUX2_X1 U7701 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n5952), .S(n6675), .Z(n6608)
         );
  INV_X1 U7702 ( .A(n6608), .ZN(n6759) );
  NOR2_X1 U7703 ( .A1(n6760), .A2(n6759), .ZN(n6758) );
  NOR2_X1 U7704 ( .A1(n6609), .A2(n6758), .ZN(n6767) );
  NAND2_X1 U7705 ( .A1(n6766), .A2(n6767), .ZN(n6765) );
  NAND2_X1 U7706 ( .A1(n6610), .A2(n6765), .ZN(n6881) );
  MUX2_X1 U7707 ( .A(n6611), .B(P1_REG2_REG_10__SCAN_IN), .S(n6886), .Z(n6880)
         );
  NAND2_X1 U7708 ( .A1(n6881), .A2(n6880), .ZN(n6879) );
  OR2_X1 U7709 ( .A1(n6886), .A2(n6611), .ZN(n6612) );
  NAND2_X1 U7710 ( .A1(n6879), .A2(n6612), .ZN(n6911) );
  NOR2_X1 U7711 ( .A1(n6920), .A2(n5746), .ZN(n6614) );
  INV_X1 U7712 ( .A(n6920), .ZN(n6613) );
  OAI22_X1 U7713 ( .A1(n6911), .A2(n6614), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n6613), .ZN(n7025) );
  NAND2_X1 U7714 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6643), .ZN(n6615) );
  OAI21_X1 U7715 ( .B1(n6643), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6615), .ZN(
        n7024) );
  NOR2_X1 U7716 ( .A1(n7025), .A2(n7024), .ZN(n7023) );
  AOI21_X1 U7717 ( .B1(n6643), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7023), .ZN(
        n7090) );
  NAND2_X1 U7718 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n6644), .ZN(n6616) );
  OAI21_X1 U7719 ( .B1(n6644), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6616), .ZN(
        n7089) );
  NOR2_X1 U7720 ( .A1(n7090), .A2(n7089), .ZN(n7088) );
  AOI21_X1 U7721 ( .B1(n6644), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7088), .ZN(
        n7137) );
  NAND2_X1 U7722 ( .A1(n7138), .A2(n7137), .ZN(n7136) );
  OR2_X1 U7723 ( .A1(n7144), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6617) );
  NAND2_X1 U7724 ( .A1(n7136), .A2(n6617), .ZN(n7729) );
  XNOR2_X1 U7725 ( .A(n7729), .B(n7730), .ZN(n6619) );
  INV_X1 U7726 ( .A(n8463), .ZN(n10746) );
  NAND2_X1 U7727 ( .A1(n10746), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8149) );
  INV_X1 U7728 ( .A(n8149), .ZN(n6618) );
  NAND2_X1 U7729 ( .A1(n10742), .A2(n6618), .ZN(n6908) );
  NOR2_X1 U7730 ( .A1(n6619), .A2(n8182), .ZN(n7731) );
  AOI211_X1 U7731 ( .C1(n8182), .C2(n6619), .A(n9869), .B(n7731), .ZN(n6653)
         );
  INV_X1 U7732 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11015) );
  INV_X1 U7733 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6620) );
  AOI22_X1 U7734 ( .A1(n6969), .A2(n6620), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n7144), .ZN(n7142) );
  INV_X1 U7735 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10988) );
  NOR2_X1 U7736 ( .A1(n7085), .A2(n10988), .ZN(n6621) );
  AOI21_X1 U7737 ( .B1(n10988), .B2(n7085), .A(n6621), .ZN(n7083) );
  INV_X1 U7738 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6637) );
  MUX2_X1 U7739 ( .A(n6637), .B(P1_REG1_REG_10__SCAN_IN), .S(n6886), .Z(n6884)
         );
  OR2_X1 U7740 ( .A1(n6771), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6636) );
  INV_X1 U7741 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6622) );
  MUX2_X1 U7742 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n6622), .S(n6771), .Z(n6769)
         );
  INV_X1 U7743 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6623) );
  XNOR2_X1 U7744 ( .A(n6626), .B(n6623), .ZN(n6982) );
  INV_X1 U7745 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10744) );
  NAND2_X1 U7746 ( .A1(P1_REG1_REG_1__SCAN_IN), .A2(n10759), .ZN(n6624) );
  OAI21_X1 U7747 ( .B1(n10759), .B2(P1_REG1_REG_1__SCAN_IN), .A(n6624), .ZN(
        n10756) );
  NOR3_X1 U7748 ( .A1(n5775), .A2(n10744), .A3(n10756), .ZN(n10755) );
  AOI21_X1 U7749 ( .B1(n10759), .B2(P1_REG1_REG_1__SCAN_IN), .A(n10755), .ZN(
        n6994) );
  XNOR2_X1 U7750 ( .A(n6672), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n6993) );
  NOR2_X1 U7751 ( .A1(n6994), .A2(n6993), .ZN(n6992) );
  AOI21_X1 U7752 ( .B1(n6672), .B2(P1_REG1_REG_2__SCAN_IN), .A(n6992), .ZN(
        n6856) );
  NAND2_X1 U7753 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(n6858), .ZN(n6625) );
  OAI21_X1 U7754 ( .B1(n6858), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6625), .ZN(
        n6855) );
  NOR2_X1 U7755 ( .A1(n6856), .A2(n6855), .ZN(n6854) );
  AOI21_X1 U7756 ( .B1(n6858), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6854), .ZN(
        n6981) );
  NAND2_X1 U7757 ( .A1(n6982), .A2(n6981), .ZN(n6628) );
  OR2_X1 U7758 ( .A1(n6626), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6627) );
  NAND2_X1 U7759 ( .A1(n6628), .A2(n6627), .ZN(n6709) );
  OR2_X1 U7760 ( .A1(n6711), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6629) );
  NAND2_X1 U7761 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6711), .ZN(n6630) );
  NAND2_X1 U7762 ( .A1(n6629), .A2(n6630), .ZN(n6708) );
  OR2_X1 U7763 ( .A1(n6709), .A2(n6708), .ZN(n6706) );
  NAND2_X1 U7764 ( .A1(n6706), .A2(n6630), .ZN(n6868) );
  XNOR2_X1 U7765 ( .A(n6872), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n6869) );
  NAND2_X1 U7766 ( .A1(n6868), .A2(n6869), .ZN(n6867) );
  NAND2_X1 U7767 ( .A1(n6631), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U7768 ( .A1(n6867), .A2(n6632), .ZN(n6742) );
  INV_X1 U7769 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6633) );
  XNOR2_X1 U7770 ( .A(n6740), .B(n6633), .ZN(n6741) );
  OR2_X1 U7771 ( .A1(n6742), .A2(n6741), .ZN(n6744) );
  NAND2_X1 U7772 ( .A1(n6740), .A2(n6633), .ZN(n6634) );
  NAND2_X1 U7773 ( .A1(n6744), .A2(n6634), .ZN(n6752) );
  INV_X1 U7774 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6635) );
  MUX2_X1 U7775 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6635), .S(n6675), .Z(n6753)
         );
  NAND2_X1 U7776 ( .A1(n6752), .A2(n6753), .ZN(n6751) );
  OAI21_X1 U7777 ( .B1(n6675), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6751), .ZN(
        n6770) );
  NAND2_X1 U7778 ( .A1(n6769), .A2(n6770), .ZN(n6768) );
  NAND2_X1 U7779 ( .A1(n6636), .A2(n6768), .ZN(n6883) );
  NAND2_X1 U7780 ( .A1(n6884), .A2(n6883), .ZN(n6882) );
  NAND2_X1 U7781 ( .A1(n6886), .A2(n6637), .ZN(n6638) );
  NAND2_X1 U7782 ( .A1(n6882), .A2(n6638), .ZN(n6913) );
  INV_X1 U7783 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6639) );
  MUX2_X1 U7784 ( .A(n6639), .B(P1_REG1_REG_11__SCAN_IN), .S(n6920), .Z(n6914)
         );
  NAND2_X1 U7785 ( .A1(n6913), .A2(n6914), .ZN(n6912) );
  NAND2_X1 U7786 ( .A1(n6920), .A2(n6639), .ZN(n6640) );
  NAND2_X1 U7787 ( .A1(n6912), .A2(n6640), .ZN(n7018) );
  OR2_X1 U7788 ( .A1(n6643), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6642) );
  NAND2_X1 U7789 ( .A1(n6643), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6641) );
  AND2_X1 U7790 ( .A1(n6642), .A2(n6641), .ZN(n7019) );
  NAND2_X1 U7791 ( .A1(n7018), .A2(n7019), .ZN(n7017) );
  OAI21_X1 U7792 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n6643), .A(n7017), .ZN(
        n7084) );
  NAND2_X1 U7793 ( .A1(n7083), .A2(n7084), .ZN(n7082) );
  OAI21_X1 U7794 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n6644), .A(n7082), .ZN(
        n7141) );
  NAND2_X1 U7795 ( .A1(n7142), .A2(n7141), .ZN(n7140) );
  OR2_X1 U7796 ( .A1(n7144), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6645) );
  NAND2_X1 U7797 ( .A1(n7140), .A2(n6645), .ZN(n7736) );
  XNOR2_X1 U7798 ( .A(n7736), .B(n7730), .ZN(n6647) );
  NOR2_X1 U7799 ( .A1(n6979), .A2(P1_U3084), .ZN(n8194) );
  AND2_X1 U7800 ( .A1(n8194), .A2(n8463), .ZN(n6646) );
  NAND2_X1 U7801 ( .A1(n10742), .A2(n6646), .ZN(n10754) );
  NOR2_X1 U7802 ( .A1(n6647), .A2(n11015), .ZN(n7737) );
  AOI211_X1 U7803 ( .C1(n11015), .C2(n6647), .A(n10754), .B(n7737), .ZN(n6652)
         );
  OR2_X1 U7804 ( .A1(P1_U3083), .A2(n6648), .ZN(n9884) );
  INV_X1 U7805 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n6649) );
  NOR2_X1 U7806 ( .A1(n9884), .A2(n6649), .ZN(n6651) );
  NAND2_X1 U7807 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9557) );
  OAI21_X1 U7808 ( .B1(n9899), .B2(n7730), .A(n9557), .ZN(n6650) );
  OR4_X1 U7809 ( .A1(n6653), .A2(n6652), .A3(n6651), .A4(n6650), .ZN(P1_U3256)
         );
  INV_X1 U7810 ( .A(n10759), .ZN(n6655) );
  AND2_X1 U7811 ( .A1(n5668), .A2(P1_U3084), .ZN(n10660) );
  OAI222_X1 U7812 ( .A1(P1_U3084), .A2(n6655), .B1(n10265), .B2(n6658), .C1(
        n6654), .C2(n10267), .ZN(P1_U3352) );
  OAI222_X1 U7813 ( .A1(n6872), .A2(P1_U3084), .B1(n10265), .B2(n7325), .C1(
        n10584), .C2(n10267), .ZN(P1_U3347) );
  INV_X1 U7814 ( .A(n10267), .ZN(n10658) );
  AOI22_X1 U7815 ( .A1(n10658), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n6858), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6656) );
  OAI21_X1 U7816 ( .B1(n6665), .B2(n10265), .A(n6656), .ZN(P1_U3350) );
  AOI22_X1 U7817 ( .A1(n6711), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n10658), .ZN(n6657) );
  OAI21_X1 U7818 ( .B1(n7103), .B2(n10265), .A(n6657), .ZN(P1_U3348) );
  AND2_X1 U7819 ( .A1(n5668), .A2(P2_U3152), .ZN(n6701) );
  NOR2_X1 U7820 ( .A1(n5668), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9420) );
  OAI222_X1 U7821 ( .A1(n5036), .A2(n6659), .B1(n8494), .B2(n6658), .C1(
        P2_U3152), .C2(n10791), .ZN(P2_U3357) );
  INV_X1 U7822 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7105) );
  NAND2_X1 U7823 ( .A1(n6660), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6661) );
  MUX2_X1 U7824 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6661), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n6662) );
  OR2_X1 U7825 ( .A1(n6660), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n6663) );
  INV_X1 U7826 ( .A(n6809), .ZN(n7106) );
  OAI222_X1 U7827 ( .A1(n5036), .A2(n7105), .B1(n8494), .B2(n7103), .C1(
        P2_U3152), .C2(n7106), .ZN(P2_U3353) );
  INV_X1 U7828 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7326) );
  NAND2_X1 U7829 ( .A1(n6663), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6664) );
  XNOR2_X1 U7830 ( .A(n6664), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6844) );
  INV_X1 U7831 ( .A(n6844), .ZN(n7327) );
  OAI222_X1 U7832 ( .A1(n5036), .A2(n7326), .B1(n8494), .B2(n7325), .C1(
        P2_U3152), .C2(n7327), .ZN(P2_U3352) );
  OAI222_X1 U7833 ( .A1(n5036), .A2(n5137), .B1(n8494), .B2(n6665), .C1(
        P2_U3152), .C2(n6837), .ZN(P2_U3355) );
  OR2_X1 U7834 ( .A1(n6666), .A2(n7051), .ZN(n6667) );
  XNOR2_X1 U7835 ( .A(n6667), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6805) );
  INV_X1 U7836 ( .A(n6805), .ZN(n7098) );
  INV_X1 U7837 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6866) );
  OAI222_X1 U7838 ( .A1(n7098), .A2(P2_U3152), .B1(n8494), .B2(n7095), .C1(
        n5036), .C2(n6866), .ZN(P2_U3354) );
  OAI222_X1 U7839 ( .A1(n5036), .A2(n6668), .B1(n8494), .B2(n6673), .C1(
        P2_U3152), .C2(n6793), .ZN(P2_U3356) );
  INV_X1 U7840 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7448) );
  NOR2_X1 U7841 ( .A1(n6660), .A2(n6669), .ZN(n6670) );
  OR2_X1 U7842 ( .A1(n6670), .A2(n7051), .ZN(n6671) );
  XNOR2_X1 U7843 ( .A(n6671), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6946) );
  INV_X1 U7844 ( .A(n6946), .ZN(n7449) );
  OAI222_X1 U7845 ( .A1(n5036), .A2(n7448), .B1(n8494), .B2(n7447), .C1(
        P2_U3152), .C2(n7449), .ZN(P2_U3351) );
  OAI222_X1 U7846 ( .A1(n6740), .A2(P1_U3084), .B1(n10265), .B2(n7447), .C1(
        n10586), .C2(n10267), .ZN(P1_U3346) );
  INV_X1 U7847 ( .A(n6672), .ZN(n6997) );
  OAI222_X1 U7848 ( .A1(n6997), .A2(P1_U3084), .B1(n10265), .B2(n6673), .C1(
        n5819), .C2(n10267), .ZN(P1_U3351) );
  INV_X1 U7849 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6674) );
  OAI222_X1 U7850 ( .A1(n6985), .A2(P1_U3084), .B1(n10265), .B2(n7095), .C1(
        n6674), .C2(n10267), .ZN(P1_U3349) );
  INV_X1 U7851 ( .A(n6675), .ZN(n6757) );
  INV_X1 U7852 ( .A(n7523), .ZN(n6678) );
  OAI222_X1 U7853 ( .A1(n6757), .A2(P1_U3084), .B1(n10265), .B2(n6678), .C1(
        n6676), .C2(n10267), .ZN(P1_U3345) );
  XNOR2_X1 U7854 ( .A(n6677), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7007) );
  INV_X1 U7855 ( .A(n7007), .ZN(n7527) );
  OAI222_X1 U7856 ( .A1(n7527), .A2(P2_U3152), .B1(n8494), .B2(n6678), .C1(
        n5036), .C2(n7524), .ZN(P2_U3350) );
  NOR2_X1 U7857 ( .A1(n6679), .A2(P2_U3152), .ZN(n6778) );
  NAND2_X1 U7858 ( .A1(n10702), .A2(n7176), .ZN(n6680) );
  NAND2_X1 U7859 ( .A1(n6680), .A2(n7537), .ZN(n6681) );
  OAI21_X1 U7860 ( .B1(n10702), .B2(n6778), .A(n6681), .ZN(n10787) );
  NOR2_X1 U7861 ( .A1(n10800), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7862 ( .A(n7536), .ZN(n6684) );
  OAI222_X1 U7863 ( .A1(n6682), .A2(P1_U3084), .B1(n10265), .B2(n6684), .C1(
        n10272), .C2(n10267), .ZN(P1_U3344) );
  NAND2_X1 U7864 ( .A1(n6683), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6693) );
  XNOR2_X1 U7865 ( .A(n6693), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7538) );
  INV_X1 U7866 ( .A(n7538), .ZN(n7156) );
  OAI222_X1 U7867 ( .A1(n5036), .A2(n6685), .B1(n8494), .B2(n6684), .C1(
        P2_U3152), .C2(n7156), .ZN(P2_U3349) );
  INV_X1 U7868 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9903) );
  NAND2_X1 U7869 ( .A1(n5040), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6688) );
  INV_X1 U7870 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6686) );
  OR2_X1 U7871 ( .A1(n8432), .A2(n6686), .ZN(n6687) );
  OAI211_X1 U7872 ( .C1(n8430), .C2(n9903), .A(n6688), .B(n6687), .ZN(n9902)
         );
  NAND2_X1 U7873 ( .A1(n9902), .A2(P1_U4006), .ZN(n6689) );
  OAI21_X1 U7874 ( .B1(P1_U4006), .B2(n9417), .A(n6689), .ZN(P1_U3586) );
  INV_X1 U7875 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6691) );
  INV_X1 U7876 ( .A(n7221), .ZN(n7198) );
  NAND2_X1 U7877 ( .A1(n7198), .A2(P2_U3966), .ZN(n6690) );
  OAI21_X1 U7878 ( .B1(P2_U3966), .B2(n6691), .A(n6690), .ZN(P2_U3552) );
  INV_X1 U7879 ( .A(n7748), .ZN(n6716) );
  NAND2_X1 U7880 ( .A1(n6693), .A2(n6692), .ZN(n6694) );
  NAND2_X1 U7881 ( .A1(n6694), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6696) );
  NAND2_X1 U7882 ( .A1(n6696), .A2(n6695), .ZN(n6699) );
  OR2_X1 U7883 ( .A1(n6696), .A2(n6695), .ZN(n6697) );
  INV_X1 U7884 ( .A(n7749), .ZN(n7613) );
  OAI222_X1 U7885 ( .A1(n8494), .A2(n6716), .B1(n7613), .B2(P2_U3152), .C1(
        n6698), .C2(n5036), .ZN(P2_U3348) );
  INV_X1 U7886 ( .A(n7781), .ZN(n6729) );
  NAND2_X1 U7887 ( .A1(n6699), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6700) );
  XNOR2_X1 U7888 ( .A(n6700), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9004) );
  AOI22_X1 U7889 ( .A1(n9004), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n6701), .ZN(n6702) );
  OAI21_X1 U7890 ( .B1(n6729), .B2(n8494), .A(n6702), .ZN(P2_U3347) );
  AOI21_X1 U7891 ( .B1(n6705), .B2(n6704), .A(n6703), .ZN(n6714) );
  AND2_X1 U7892 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7065) );
  INV_X1 U7893 ( .A(n6706), .ZN(n6707) );
  AOI211_X1 U7894 ( .C1(n6709), .C2(n6708), .A(n6707), .B(n10754), .ZN(n6710)
         );
  AOI211_X1 U7895 ( .C1(n10760), .C2(n6711), .A(n7065), .B(n6710), .ZN(n6713)
         );
  INV_X1 U7896 ( .A(n9884), .ZN(n10761) );
  NAND2_X1 U7897 ( .A1(n10761), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n6712) );
  OAI211_X1 U7898 ( .C1(n6714), .C2(n9869), .A(n6713), .B(n6712), .ZN(P1_U3246) );
  NAND2_X1 U7899 ( .A1(n10110), .A2(P1_U4006), .ZN(n6715) );
  OAI21_X1 U7900 ( .B1(n6175), .B2(P1_U4006), .A(n6715), .ZN(P1_U3573) );
  OAI222_X1 U7901 ( .A1(n6886), .A2(P1_U3084), .B1(n10267), .B2(n5992), .C1(
        n6716), .C2(n10265), .ZN(P1_U3343) );
  NAND2_X1 U7902 ( .A1(n7648), .A2(P1_U4006), .ZN(n6717) );
  OAI21_X1 U7903 ( .B1(P1_U4006), .B2(n7524), .A(n6717), .ZN(P1_U3563) );
  INV_X2 U7904 ( .A(n6730), .ZN(n8047) );
  NAND2_X1 U7905 ( .A1(n8047), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6727) );
  INV_X1 U7906 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7769) );
  OR2_X1 U7907 ( .A1(n8253), .A2(n7769), .ZN(n6726) );
  INV_X1 U7908 ( .A(n7110), .ZN(n6718) );
  NAND2_X1 U7909 ( .A1(n6718), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7119) );
  INV_X1 U7910 ( .A(n7119), .ZN(n6719) );
  NAND2_X1 U7911 ( .A1(n6719), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7318) );
  INV_X1 U7912 ( .A(n7318), .ZN(n6720) );
  NAND2_X1 U7913 ( .A1(n6720), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7529) );
  NAND2_X1 U7914 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n6721) );
  INV_X1 U7915 ( .A(n7530), .ZN(n6722) );
  NAND2_X1 U7916 ( .A1(n6722), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7754) );
  INV_X1 U7917 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10527) );
  NAND2_X1 U7918 ( .A1(n7530), .A2(n10527), .ZN(n6723) );
  NAND2_X1 U7919 ( .A1(n7754), .A2(n6723), .ZN(n7843) );
  OR2_X1 U7920 ( .A1(n8321), .A2(n7843), .ZN(n6725) );
  INV_X1 U7921 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7157) );
  OR2_X1 U7922 ( .A1(n8324), .A2(n7157), .ZN(n6724) );
  INV_X1 U7923 ( .A(n8929), .ZN(n7882) );
  NAND2_X1 U7924 ( .A1(n7882), .A2(P2_U3966), .ZN(n6728) );
  OAI21_X1 U7925 ( .B1(P2_U3966), .B2(n5992), .A(n6728), .ZN(P2_U3562) );
  OAI222_X1 U7926 ( .A1(P1_U3084), .A2(n6920), .B1(n10265), .B2(n6729), .C1(
        n10279), .C2(n10267), .ZN(P1_U3342) );
  INV_X1 U7927 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10287) );
  INV_X1 U7928 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6733) );
  NAND2_X1 U7929 ( .A1(n8370), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6732) );
  NAND2_X1 U7930 ( .A1(n8047), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6731) );
  OAI211_X1 U7931 ( .C1(n8324), .C2(n6733), .A(n6732), .B(n6731), .ZN(n9094)
         );
  NAND2_X1 U7932 ( .A1(n9094), .A2(P2_U3966), .ZN(n6734) );
  OAI21_X1 U7933 ( .B1(P2_U3966), .B2(n10287), .A(n6734), .ZN(P2_U3583) );
  INV_X1 U7934 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7059) );
  NAND2_X1 U7935 ( .A1(n10129), .A2(P1_U4006), .ZN(n6735) );
  OAI21_X1 U7936 ( .B1(n7059), .B2(P1_U4006), .A(n6735), .ZN(P1_U3572) );
  INV_X1 U7937 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6750) );
  NOR2_X1 U7938 ( .A1(n6737), .A2(n6736), .ZN(n6739) );
  INV_X1 U7939 ( .A(n9869), .ZN(n10763) );
  OAI21_X1 U7940 ( .B1(n6739), .B2(n6738), .A(n10763), .ZN(n6749) );
  INV_X1 U7941 ( .A(n6740), .ZN(n6747) );
  NAND2_X1 U7942 ( .A1(n6742), .A2(n6741), .ZN(n6743) );
  AND2_X1 U7943 ( .A1(n6744), .A2(n6743), .ZN(n6745) );
  NAND2_X1 U7944 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7426) );
  OAI21_X1 U7945 ( .B1(n10754), .B2(n6745), .A(n7426), .ZN(n6746) );
  AOI21_X1 U7946 ( .B1(n10760), .B2(n6747), .A(n6746), .ZN(n6748) );
  OAI211_X1 U7947 ( .C1(n9884), .C2(n6750), .A(n6749), .B(n6748), .ZN(P1_U3248) );
  INV_X1 U7948 ( .A(n10754), .ZN(n10745) );
  OAI21_X1 U7949 ( .B1(n6753), .B2(n6752), .A(n6751), .ZN(n6755) );
  INV_X1 U7950 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6754) );
  NOR2_X1 U7951 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6754), .ZN(n7678) );
  AOI21_X1 U7952 ( .B1(n10745), .B2(n6755), .A(n7678), .ZN(n6756) );
  OAI21_X1 U7953 ( .B1(n6757), .B2(n9899), .A(n6756), .ZN(n6763) );
  AOI21_X1 U7954 ( .B1(n6760), .B2(n6759), .A(n6758), .ZN(n6761) );
  NOR2_X1 U7955 ( .A1(n6761), .A2(n9869), .ZN(n6762) );
  AOI211_X1 U7956 ( .C1(n10761), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n6763), .B(
        n6762), .ZN(n6764) );
  INV_X1 U7957 ( .A(n6764), .ZN(P1_U3249) );
  OAI211_X1 U7958 ( .C1(n6767), .C2(n6766), .A(n10763), .B(n6765), .ZN(n6776)
         );
  OAI21_X1 U7959 ( .B1(n6770), .B2(n6769), .A(n6768), .ZN(n6774) );
  INV_X1 U7960 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7916) );
  AND2_X1 U7961 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7649) );
  AOI21_X1 U7962 ( .B1(n10760), .B2(n6771), .A(n7649), .ZN(n6772) );
  OAI21_X1 U7963 ( .B1(n7916), .B2(n9884), .A(n6772), .ZN(n6773) );
  AOI21_X1 U7964 ( .B1(n10745), .B2(n6774), .A(n6773), .ZN(n6775) );
  NAND2_X1 U7965 ( .A1(n6776), .A2(n6775), .ZN(P1_U3250) );
  AOI22_X1 U7966 ( .A1(n6805), .A2(n6583), .B1(P2_REG2_REG_4__SCAN_IN), .B2(
        n7098), .ZN(n6786) );
  INV_X1 U7967 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10794) );
  AOI22_X1 U7968 ( .A1(n6791), .A2(n6540), .B1(P2_REG2_REG_1__SCAN_IN), .B2(
        n10791), .ZN(n10781) );
  NOR3_X1 U7969 ( .A1(n10794), .A2(n10775), .A3(n10781), .ZN(n10783) );
  AOI22_X1 U7970 ( .A1(n6788), .A2(n7313), .B1(P2_REG2_REG_3__SCAN_IN), .B2(
        n6837), .ZN(n6830) );
  NOR2_X1 U7971 ( .A1(n6829), .A2(n6830), .ZN(n6828) );
  NOR2_X1 U7972 ( .A1(n6785), .A2(n6786), .ZN(n6804) );
  NAND2_X1 U7973 ( .A1(n10702), .A2(n6777), .ZN(n6779) );
  INV_X1 U7974 ( .A(n6778), .ZN(n8823) );
  OAI211_X1 U7975 ( .C1(n6780), .C2(P2_U3152), .A(n6779), .B(n8823), .ZN(n6781) );
  NAND2_X1 U7976 ( .A1(n6781), .A2(n7537), .ZN(n6795) );
  NAND2_X1 U7977 ( .A1(n6795), .A2(n8999), .ZN(n6787) );
  INV_X1 U7978 ( .A(n6582), .ZN(n6783) );
  INV_X1 U7979 ( .A(n8375), .ZN(n6782) );
  NAND2_X1 U7980 ( .A1(n6783), .A2(n6782), .ZN(n8818) );
  INV_X1 U7981 ( .A(n8818), .ZN(n6784) );
  AOI211_X1 U7982 ( .C1(n6786), .C2(n6785), .A(n6804), .B(n10801), .ZN(n6802)
         );
  NAND2_X1 U7983 ( .A1(n6787), .A2(n6582), .ZN(n10792) );
  MUX2_X1 U7984 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6789), .S(n6788), .Z(n6832)
         );
  MUX2_X1 U7985 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6790), .S(n10806), .Z(n10810) );
  MUX2_X1 U7986 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6792), .S(n6791), .Z(n10796)
         );
  NAND3_X1 U7987 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n10796), .ZN(n10795) );
  OAI21_X1 U7988 ( .B1(n10791), .B2(n6792), .A(n10795), .ZN(n10811) );
  NAND2_X1 U7989 ( .A1(n10810), .A2(n10811), .ZN(n10808) );
  OAI21_X1 U7990 ( .B1(n6793), .B2(n6790), .A(n10808), .ZN(n6833) );
  NAND2_X1 U7991 ( .A1(n6832), .A2(n6833), .ZN(n6831) );
  OAI21_X1 U7992 ( .B1(n6837), .B2(n6789), .A(n6831), .ZN(n6798) );
  MUX2_X1 U7993 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6794), .S(n6805), .Z(n6797)
         );
  INV_X1 U7994 ( .A(n6795), .ZN(n6796) );
  NAND2_X1 U7995 ( .A1(n6796), .A2(n8375), .ZN(n10773) );
  NAND2_X1 U7996 ( .A1(n6797), .A2(n6798), .ZN(n6810) );
  OAI211_X1 U7997 ( .C1(n6798), .C2(n6797), .A(n10809), .B(n6810), .ZN(n6800)
         );
  INV_X1 U7998 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10292) );
  NOR2_X1 U7999 ( .A1(n10292), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7362) );
  AOI21_X1 U8000 ( .B1(n10800), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n7362), .ZN(
        n6799) );
  OAI211_X1 U8001 ( .C1(n10792), .C2(n7098), .A(n6800), .B(n6799), .ZN(n6801)
         );
  OR2_X1 U8002 ( .A1(n6802), .A2(n6801), .ZN(P2_U3249) );
  NAND2_X1 U8003 ( .A1(n6844), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6803) );
  OAI21_X1 U8004 ( .B1(n6844), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6803), .ZN(
        n6808) );
  AOI21_X1 U8005 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n6805), .A(n6804), .ZN(
        n6819) );
  NAND2_X1 U8006 ( .A1(n6809), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6806) );
  OAI21_X1 U8007 ( .B1(n6809), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6806), .ZN(
        n6820) );
  NOR2_X1 U8008 ( .A1(n6819), .A2(n6820), .ZN(n6818) );
  NOR2_X1 U8009 ( .A1(n6807), .A2(n6808), .ZN(n6841) );
  AOI211_X1 U8010 ( .C1(n6808), .C2(n6807), .A(n6841), .B(n10801), .ZN(n6817)
         );
  NAND2_X1 U8011 ( .A1(n6809), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6811) );
  INV_X1 U8012 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7112) );
  MUX2_X1 U8013 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n7112), .S(n6809), .Z(n6822)
         );
  OAI21_X1 U8014 ( .B1(n7098), .B2(n6794), .A(n6810), .ZN(n6823) );
  NAND2_X1 U8015 ( .A1(n6822), .A2(n6823), .ZN(n6821) );
  NAND2_X1 U8016 ( .A1(n6811), .A2(n6821), .ZN(n6813) );
  INV_X1 U8017 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7121) );
  MUX2_X1 U8018 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n7121), .S(n6844), .Z(n6812)
         );
  NAND2_X1 U8019 ( .A1(n6812), .A2(n6813), .ZN(n6845) );
  OAI211_X1 U8020 ( .C1(n6813), .C2(n6812), .A(n10809), .B(n6845), .ZN(n6815)
         );
  INV_X1 U8021 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10539) );
  NOR2_X1 U8022 ( .A1(n10539), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7377) );
  AOI21_X1 U8023 ( .B1(n10800), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7377), .ZN(
        n6814) );
  OAI211_X1 U8024 ( .C1(n10792), .C2(n7327), .A(n6815), .B(n6814), .ZN(n6816)
         );
  OR2_X1 U8025 ( .A1(n6817), .A2(n6816), .ZN(P2_U3251) );
  AOI211_X1 U8026 ( .C1(n6820), .C2(n6819), .A(n6818), .B(n10801), .ZN(n6827)
         );
  OAI211_X1 U8027 ( .C1(n6823), .C2(n6822), .A(n10809), .B(n6821), .ZN(n6825)
         );
  INV_X1 U8028 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10459) );
  NOR2_X1 U8029 ( .A1(n10459), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7126) );
  AOI21_X1 U8030 ( .B1(n10800), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7126), .ZN(
        n6824) );
  OAI211_X1 U8031 ( .C1(n10792), .C2(n7106), .A(n6825), .B(n6824), .ZN(n6826)
         );
  OR2_X1 U8032 ( .A1(n6827), .A2(n6826), .ZN(P2_U3250) );
  AOI211_X1 U8033 ( .C1(n6830), .C2(n6829), .A(n6828), .B(n10801), .ZN(n6839)
         );
  OAI211_X1 U8034 ( .C1(n6833), .C2(n6832), .A(n10809), .B(n6831), .ZN(n6836)
         );
  INV_X1 U8035 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10525) );
  NOR2_X1 U8036 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10525), .ZN(n6834) );
  AOI21_X1 U8037 ( .B1(n10800), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6834), .ZN(
        n6835) );
  OAI211_X1 U8038 ( .C1(n10792), .C2(n6837), .A(n6836), .B(n6835), .ZN(n6838)
         );
  OR2_X1 U8039 ( .A1(n6839), .A2(n6838), .ZN(P2_U3248) );
  INV_X1 U8040 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6840) );
  AOI22_X1 U8041 ( .A1(n6946), .A2(n6840), .B1(P2_REG2_REG_7__SCAN_IN), .B2(
        n7449), .ZN(n6843) );
  AOI21_X1 U8042 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n6844), .A(n6841), .ZN(
        n6842) );
  NOR2_X1 U8043 ( .A1(n6842), .A2(n6843), .ZN(n6945) );
  AOI211_X1 U8044 ( .C1(n6843), .C2(n6842), .A(n6945), .B(n10801), .ZN(n6853)
         );
  NAND2_X1 U8045 ( .A1(n6844), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6846) );
  NAND2_X1 U8046 ( .A1(n6846), .A2(n6845), .ZN(n6848) );
  INV_X1 U8047 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7320) );
  MUX2_X1 U8048 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7320), .S(n6946), .Z(n6847)
         );
  NAND2_X1 U8049 ( .A1(n6847), .A2(n6848), .ZN(n6949) );
  OAI211_X1 U8050 ( .C1(n6848), .C2(n6847), .A(n10809), .B(n6949), .ZN(n6851)
         );
  INV_X1 U8051 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10514) );
  NOR2_X1 U8052 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10514), .ZN(n6849) );
  AOI21_X1 U8053 ( .B1(n10800), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6849), .ZN(
        n6850) );
  OAI211_X1 U8054 ( .C1(n10792), .C2(n7449), .A(n6851), .B(n6850), .ZN(n6852)
         );
  OR2_X1 U8055 ( .A1(n6853), .A2(n6852), .ZN(P2_U3252) );
  INV_X1 U8056 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6864) );
  INV_X1 U8057 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7253) );
  NOR2_X1 U8058 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7253), .ZN(n7042) );
  AOI211_X1 U8059 ( .C1(n6856), .C2(n6855), .A(n6854), .B(n10754), .ZN(n6857)
         );
  AOI211_X1 U8060 ( .C1(n10760), .C2(n6858), .A(n7042), .B(n6857), .ZN(n6863)
         );
  OAI211_X1 U8061 ( .C1(n6861), .C2(n6860), .A(n10763), .B(n6859), .ZN(n6862)
         );
  OAI211_X1 U8062 ( .C1(n9884), .C2(n6864), .A(n6863), .B(n6862), .ZN(P1_U3244) );
  NAND2_X1 U8063 ( .A1(n5875), .A2(P1_U4006), .ZN(n6865) );
  OAI21_X1 U8064 ( .B1(P1_U4006), .B2(n6866), .A(n6865), .ZN(P1_U3559) );
  OAI211_X1 U8065 ( .C1(n6869), .C2(n6868), .A(n10745), .B(n6867), .ZN(n6871)
         );
  INV_X1 U8066 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6870) );
  OR2_X1 U8067 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6870), .ZN(n7169) );
  OAI211_X1 U8068 ( .C1(n9899), .C2(n6872), .A(n6871), .B(n7169), .ZN(n6877)
         );
  AOI211_X1 U8069 ( .C1(n6875), .C2(n6874), .A(n9869), .B(n6873), .ZN(n6876)
         );
  AOI211_X1 U8070 ( .C1(n10761), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n6877), .B(
        n6876), .ZN(n6878) );
  INV_X1 U8071 ( .A(n6878), .ZN(P1_U3247) );
  INV_X1 U8072 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7895) );
  OAI211_X1 U8073 ( .C1(n6881), .C2(n6880), .A(n6879), .B(n10763), .ZN(n6890)
         );
  OAI21_X1 U8074 ( .B1(n6884), .B2(n6883), .A(n6882), .ZN(n6888) );
  NOR2_X1 U8075 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6885), .ZN(n7948) );
  NOR2_X1 U8076 ( .A1(n9899), .A2(n6886), .ZN(n6887) );
  AOI211_X1 U8077 ( .C1(n10745), .C2(n6888), .A(n7948), .B(n6887), .ZN(n6889)
         );
  OAI211_X1 U8078 ( .C1(n7895), .C2(n9884), .A(n6890), .B(n6889), .ZN(P1_U3251) );
  INV_X1 U8079 ( .A(n7241), .ZN(n7256) );
  XNOR2_X1 U8080 ( .A(n6891), .B(n9594), .ZN(n9763) );
  NAND3_X1 U8081 ( .A1(n9763), .A2(n7287), .A3(n7293), .ZN(n6892) );
  OAI21_X1 U8082 ( .B1(n7256), .B2(n10083), .A(n6892), .ZN(n7072) );
  AOI21_X1 U8083 ( .B1(n7296), .B2(n6893), .A(n7072), .ZN(n6902) );
  OR2_X1 U8084 ( .A1(n10923), .A2(n9760), .ZN(n6897) );
  AND3_X1 U8085 ( .A1(n6895), .A2(n6894), .A3(n10257), .ZN(n6896) );
  AND3_X1 U8086 ( .A1(n6897), .A2(n6896), .A3(n7073), .ZN(n6900) );
  NAND2_X1 U8087 ( .A1(n11023), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6898) );
  OAI21_X1 U8088 ( .B1(n6902), .B2(n11023), .A(n6898), .ZN(P1_U3523) );
  INV_X1 U8089 ( .A(n11028), .ZN(n11025) );
  OR2_X1 U8090 ( .A1(n11028), .A2(n5767), .ZN(n6901) );
  OAI21_X1 U8091 ( .B1(n6902), .B2(n11025), .A(n6901), .ZN(P1_U3454) );
  INV_X1 U8092 ( .A(n7784), .ZN(n6905) );
  OAI222_X1 U8093 ( .A1(n7022), .A2(P1_U3084), .B1(n10265), .B2(n6905), .C1(
        n10442), .C2(n10267), .ZN(P1_U3341) );
  NAND2_X1 U8094 ( .A1(n6903), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6904) );
  XNOR2_X1 U8095 ( .A(n6904), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7785) );
  INV_X1 U8096 ( .A(n7785), .ZN(n7690) );
  OAI222_X1 U8097 ( .A1(n5036), .A2(n6906), .B1(n8494), .B2(n6905), .C1(
        P2_U3152), .C2(n7690), .ZN(P2_U3346) );
  INV_X1 U8098 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7658) );
  NAND2_X1 U8099 ( .A1(n10016), .A2(P1_U4006), .ZN(n6907) );
  OAI21_X1 U8100 ( .B1(n7658), .B2(P1_U4006), .A(n6907), .ZN(P1_U3576) );
  NOR2_X1 U8101 ( .A1(n6908), .A2(n5746), .ZN(n6909) );
  AOI21_X1 U8102 ( .B1(n6911), .B2(n6909), .A(n10760), .ZN(n6921) );
  NAND2_X1 U8103 ( .A1(n6920), .A2(n5746), .ZN(n6910) );
  OAI211_X1 U8104 ( .C1(n6911), .C2(n6910), .A(n7025), .B(n10763), .ZN(n6919)
         );
  OAI21_X1 U8105 ( .B1(n6914), .B2(n6913), .A(n6912), .ZN(n6917) );
  AND2_X1 U8106 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8016) );
  INV_X1 U8107 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6915) );
  NOR2_X1 U8108 ( .A1(n9884), .A2(n6915), .ZN(n6916) );
  AOI211_X1 U8109 ( .C1(n10745), .C2(n6917), .A(n8016), .B(n6916), .ZN(n6918)
         );
  OAI211_X1 U8110 ( .C1(n6921), .C2(n6920), .A(n6919), .B(n6918), .ZN(P1_U3252) );
  INV_X1 U8111 ( .A(n7754), .ZN(n6922) );
  INV_X1 U8112 ( .A(n8163), .ZN(n6924) );
  XNOR2_X1 U8113 ( .A(n8281), .B(P2_REG3_REG_23__SCAN_IN), .ZN(n9173) );
  NAND2_X1 U8114 ( .A1(n9173), .A2(n8353), .ZN(n6933) );
  INV_X1 U8115 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n6930) );
  NAND2_X1 U8116 ( .A1(n8370), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6929) );
  NAND2_X1 U8117 ( .A1(n8047), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6928) );
  OAI211_X1 U8118 ( .C1(n6930), .C2(n8324), .A(n6929), .B(n6928), .ZN(n6931)
         );
  INV_X1 U8119 ( .A(n6931), .ZN(n6932) );
  NAND2_X1 U8120 ( .A1(n6933), .A2(n6932), .ZN(n9155) );
  NAND2_X1 U8121 ( .A1(n9155), .A2(P2_U3966), .ZN(n6934) );
  OAI21_X1 U8122 ( .B1(P2_U3966), .B2(n6283), .A(n6934), .ZN(P2_U3575) );
  OAI21_X1 U8123 ( .B1(n6937), .B2(n6935), .A(n6936), .ZN(n6976) );
  INV_X1 U8124 ( .A(n6976), .ZN(n6943) );
  NAND2_X1 U8125 ( .A1(n6938), .A2(n11018), .ZN(n6940) );
  NAND4_X1 U8126 ( .A1(n6940), .A2(n10257), .A3(n6939), .A4(n7073), .ZN(n9460)
         );
  OAI22_X1 U8127 ( .A1(n7256), .A2(n9559), .B1(n9535), .B2(n9594), .ZN(n6941)
         );
  AOI21_X1 U8128 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n9460), .A(n6941), .ZN(
        n6942) );
  OAI21_X1 U8129 ( .B1(n6943), .B2(n9569), .A(n6942), .ZN(P1_U3230) );
  INV_X1 U8130 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6944) );
  AOI22_X1 U8131 ( .A1(n7007), .A2(n6944), .B1(P2_REG2_REG_8__SCAN_IN), .B2(
        n7527), .ZN(n6948) );
  NOR2_X1 U8132 ( .A1(n6947), .A2(n6948), .ZN(n7006) );
  AOI211_X1 U8133 ( .C1(n6948), .C2(n6947), .A(n7006), .B(n10801), .ZN(n6956)
         );
  OAI21_X1 U8134 ( .B1(n7449), .B2(n7320), .A(n6949), .ZN(n6951) );
  INV_X1 U8135 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7453) );
  MUX2_X1 U8136 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7453), .S(n7007), .Z(n6950)
         );
  NAND2_X1 U8137 ( .A1(n6950), .A2(n6951), .ZN(n7010) );
  OAI211_X1 U8138 ( .C1(n6951), .C2(n6950), .A(n10809), .B(n7010), .ZN(n6954)
         );
  NOR2_X1 U8139 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7592), .ZN(n6952) );
  AOI21_X1 U8140 ( .B1(n10800), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6952), .ZN(
        n6953) );
  OAI211_X1 U8141 ( .C1(n10792), .C2(n7527), .A(n6954), .B(n6953), .ZN(n6955)
         );
  OR2_X1 U8142 ( .A1(n6956), .A2(n6955), .ZN(P2_U3253) );
  INV_X1 U8143 ( .A(n7991), .ZN(n6959) );
  OR2_X1 U8144 ( .A1(n6957), .A2(n7051), .ZN(n6961) );
  XNOR2_X1 U8145 ( .A(n6961), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7992) );
  INV_X1 U8146 ( .A(n7992), .ZN(n7824) );
  OAI222_X1 U8147 ( .A1(n8494), .A2(n6959), .B1(n7824), .B2(P2_U3152), .C1(
        n6958), .C2(n5036), .ZN(P2_U3345) );
  OAI222_X1 U8148 ( .A1(P1_U3084), .A2(n7085), .B1(n10265), .B2(n6959), .C1(
        n10568), .C2(n10267), .ZN(P1_U3340) );
  INV_X1 U8149 ( .A(n8043), .ZN(n6968) );
  NAND2_X1 U8150 ( .A1(n6961), .A2(n6960), .ZN(n6962) );
  NAND2_X1 U8151 ( .A1(n6962), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6965) );
  INV_X1 U8152 ( .A(n6965), .ZN(n6963) );
  NAND2_X1 U8153 ( .A1(n6963), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n6966) );
  NAND2_X1 U8154 ( .A1(n6965), .A2(n6964), .ZN(n7045) );
  INV_X1 U8155 ( .A(n9014), .ZN(n9021) );
  INV_X1 U8156 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6967) );
  OAI222_X1 U8157 ( .A1(n8494), .A2(n6968), .B1(n9021), .B2(P2_U3152), .C1(
        n6967), .C2(n5036), .ZN(P2_U3344) );
  OAI222_X1 U8158 ( .A1(n10267), .A2(n10573), .B1(P1_U3084), .B2(n6969), .C1(
        n6968), .C2(n10265), .ZN(P1_U3339) );
  XOR2_X1 U8159 ( .A(n6971), .B(n6970), .Z(n6974) );
  INV_X1 U8160 ( .A(n10857), .ZN(n7274) );
  AOI22_X1 U8161 ( .A1(n9561), .A2(n9851), .B1(n9566), .B2(n7274), .ZN(n6973)
         );
  AOI22_X1 U8162 ( .A1(P1_REG3_REG_2__SCAN_IN), .A2(n9460), .B1(n9532), .B2(
        n7246), .ZN(n6972) );
  OAI211_X1 U8163 ( .C1(n6974), .C2(n9569), .A(n6973), .B(n6972), .ZN(P1_U3235) );
  NAND2_X1 U8164 ( .A1(n10002), .A2(P1_U4006), .ZN(n6975) );
  OAI21_X1 U8165 ( .B1(n8276), .B2(P1_U4006), .A(n6975), .ZN(P1_U3579) );
  INV_X1 U8166 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7076) );
  NOR2_X1 U8167 ( .A1(n5775), .A2(n7076), .ZN(n10765) );
  INV_X1 U8168 ( .A(n10765), .ZN(n6977) );
  MUX2_X1 U8169 ( .A(n6977), .B(n6976), .S(n8463), .Z(n6978) );
  NOR2_X1 U8170 ( .A1(n6978), .A2(n6979), .ZN(n6980) );
  AOI21_X1 U8171 ( .B1(n10746), .B2(n7076), .A(n6979), .ZN(n10741) );
  NOR2_X1 U8172 ( .A1(n10741), .A2(n10753), .ZN(n10752) );
  INV_X1 U8173 ( .A(P1_U4006), .ZN(n9852) );
  NOR3_X1 U8174 ( .A1(n6980), .A2(n10752), .A3(n9852), .ZN(n7004) );
  XNOR2_X1 U8175 ( .A(n6982), .B(n6981), .ZN(n6983) );
  AND2_X1 U8176 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n8385) );
  AOI21_X1 U8177 ( .B1(n10745), .B2(n6983), .A(n8385), .ZN(n6984) );
  OAI21_X1 U8178 ( .B1(n6985), .B2(n9899), .A(n6984), .ZN(n6991) );
  AOI21_X1 U8179 ( .B1(n6988), .B2(n6987), .A(n6986), .ZN(n6989) );
  OAI22_X1 U8180 ( .A1(n9884), .A2(n7896), .B1(n9869), .B2(n6989), .ZN(n6990)
         );
  OR3_X1 U8181 ( .A1(n7004), .A2(n6991), .A3(n6990), .ZN(P1_U3245) );
  AOI211_X1 U8182 ( .C1(n6994), .C2(n6993), .A(n6992), .B(n10754), .ZN(n6995)
         );
  AOI21_X1 U8183 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(P1_U3084), .A(n6995), .ZN(
        n6996) );
  OAI21_X1 U8184 ( .B1(n6997), .B2(n9899), .A(n6996), .ZN(n7003) );
  INV_X1 U8185 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7897) );
  OAI21_X1 U8186 ( .B1(n7000), .B2(n6999), .A(n6998), .ZN(n7001) );
  OAI22_X1 U8187 ( .A1(n9884), .A2(n7897), .B1(n9869), .B2(n7001), .ZN(n7002)
         );
  OR3_X1 U8188 ( .A1(n7004), .A2(n7003), .A3(n7002), .ZN(P1_U3243) );
  INV_X1 U8189 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7005) );
  AOI22_X1 U8190 ( .A1(n7538), .A2(n7005), .B1(P2_REG2_REG_9__SCAN_IN), .B2(
        n7156), .ZN(n7009) );
  AOI21_X1 U8191 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7007), .A(n7006), .ZN(
        n7008) );
  NOR2_X1 U8192 ( .A1(n7008), .A2(n7009), .ZN(n7151) );
  AOI211_X1 U8193 ( .C1(n7009), .C2(n7008), .A(n7151), .B(n10801), .ZN(n7016)
         );
  OAI21_X1 U8194 ( .B1(n7527), .B2(n7453), .A(n7010), .ZN(n7012) );
  INV_X1 U8195 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7528) );
  MUX2_X1 U8196 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7528), .S(n7538), .Z(n7011)
         );
  NAND2_X1 U8197 ( .A1(n7011), .A2(n7012), .ZN(n7155) );
  OAI211_X1 U8198 ( .C1(n7012), .C2(n7011), .A(n10809), .B(n7155), .ZN(n7014)
         );
  INV_X1 U8199 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10450) );
  NOR2_X1 U8200 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10450), .ZN(n7720) );
  AOI21_X1 U8201 ( .B1(n10800), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7720), .ZN(
        n7013) );
  OAI211_X1 U8202 ( .C1(n10792), .C2(n7156), .A(n7014), .B(n7013), .ZN(n7015)
         );
  OR2_X1 U8203 ( .A1(n7016), .A2(n7015), .ZN(P2_U3254) );
  NAND2_X1 U8204 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8105) );
  OAI21_X1 U8205 ( .B1(n7019), .B2(n7018), .A(n7017), .ZN(n7020) );
  NAND2_X1 U8206 ( .A1(n10745), .A2(n7020), .ZN(n7021) );
  OAI211_X1 U8207 ( .C1(n9899), .C2(n7022), .A(n8105), .B(n7021), .ZN(n7027)
         );
  AOI211_X1 U8208 ( .C1(n7025), .C2(n7024), .A(n9869), .B(n7023), .ZN(n7026)
         );
  AOI211_X1 U8209 ( .C1(n10761), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n7027), .B(
        n7026), .ZN(n7028) );
  INV_X1 U8210 ( .A(n7028), .ZN(P1_U3253) );
  AND2_X1 U8211 ( .A1(n7237), .A2(n7030), .ZN(n7225) );
  AOI211_X1 U8212 ( .C1(n7033), .C2(n7032), .A(n8953), .B(n7031), .ZN(n7034)
         );
  INV_X1 U8213 ( .A(n7034), .ZN(n7037) );
  INV_X1 U8214 ( .A(n10864), .ZN(n7186) );
  OR2_X1 U8215 ( .A1(n7845), .A2(n9272), .ZN(n8930) );
  OAI22_X1 U8216 ( .A1(n7192), .A2(n8964), .B1(n8930), .B2(n7185), .ZN(n7035)
         );
  AOI21_X1 U8217 ( .B1(n7186), .B2(n8975), .A(n7035), .ZN(n7036) );
  OAI211_X1 U8218 ( .C1(n7225), .C2(n10451), .A(n7037), .B(n7036), .ZN(
        P2_U3239) );
  XNOR2_X1 U8219 ( .A(n7039), .B(n7038), .ZN(n7040) );
  NAND2_X1 U8220 ( .A1(n7040), .A2(n9525), .ZN(n7044) );
  INV_X1 U8221 ( .A(n10870), .ZN(n7414) );
  INV_X1 U8222 ( .A(n9561), .ZN(n9529) );
  INV_X1 U8223 ( .A(n9850), .ZN(n7258) );
  INV_X1 U8224 ( .A(n5875), .ZN(n7481) );
  OAI22_X1 U8225 ( .A1(n9529), .A2(n7258), .B1(n7481), .B2(n9559), .ZN(n7041)
         );
  AOI211_X1 U8226 ( .C1(n7414), .C2(n9566), .A(n7042), .B(n7041), .ZN(n7043)
         );
  OAI211_X1 U8227 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9564), .A(n7044), .B(
        n7043), .ZN(P1_U3216) );
  INV_X1 U8228 ( .A(n8154), .ZN(n7047) );
  OAI222_X1 U8229 ( .A1(n7730), .A2(P1_U3084), .B1(n10265), .B2(n7047), .C1(
        n10574), .C2(n10267), .ZN(P1_U3338) );
  NAND2_X1 U8230 ( .A1(n7045), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7046) );
  XNOR2_X1 U8231 ( .A(n7046), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9034) );
  INV_X1 U8232 ( .A(n9034), .ZN(n9027) );
  OAI222_X1 U8233 ( .A1(n5036), .A2(n7048), .B1(n8494), .B2(n7047), .C1(
        P2_U3152), .C2(n9027), .ZN(P2_U3343) );
  INV_X1 U8234 ( .A(n8208), .ZN(n7055) );
  NOR2_X1 U8235 ( .A1(n7049), .A2(n7051), .ZN(n7050) );
  MUX2_X1 U8236 ( .A(n7051), .B(n7050), .S(P2_IR_REG_16__SCAN_IN), .Z(n7052)
         );
  INV_X1 U8237 ( .A(n7052), .ZN(n7053) );
  AND2_X1 U8238 ( .A1(n7053), .A2(n7057), .ZN(n9054) );
  INV_X1 U8239 ( .A(n9054), .ZN(n9047) );
  OAI222_X1 U8240 ( .A1(n8494), .A2(n7055), .B1(n9047), .B2(P2_U3152), .C1(
        n7054), .C2(n5036), .ZN(P2_U3342) );
  OAI222_X1 U8241 ( .A1(P1_U3084), .A2(n7743), .B1(n10265), .B2(n7055), .C1(
        n10569), .C2(n10267), .ZN(P1_U3337) );
  INV_X1 U8242 ( .A(n8213), .ZN(n7060) );
  AOI22_X1 U8243 ( .A1(n9875), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10658), .ZN(n7056) );
  OAI21_X1 U8244 ( .B1(n7060), .B2(n10265), .A(n7056), .ZN(P1_U3336) );
  NAND2_X1 U8245 ( .A1(n7057), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7058) );
  XNOR2_X1 U8246 ( .A(n7058), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9061) );
  INV_X1 U8247 ( .A(n9061), .ZN(n9066) );
  OAI222_X1 U8248 ( .A1(n8494), .A2(n7060), .B1(n5036), .B2(n7059), .C1(
        P2_U3152), .C2(n9066), .ZN(P2_U3341) );
  XNOR2_X1 U8249 ( .A(n7063), .B(n7062), .ZN(n7064) );
  XNOR2_X1 U8250 ( .A(n7061), .B(n7064), .ZN(n7071) );
  INV_X1 U8251 ( .A(n7500), .ZN(n10890) );
  NOR2_X1 U8252 ( .A1(n9535), .A2(n10890), .ZN(n7069) );
  NAND2_X1 U8253 ( .A1(n9561), .A2(n5875), .ZN(n7067) );
  INV_X1 U8254 ( .A(n7065), .ZN(n7066) );
  OAI211_X1 U8255 ( .C1(n7572), .C2(n9559), .A(n7067), .B(n7066), .ZN(n7068)
         );
  AOI211_X1 U8256 ( .C1(n7476), .C2(n9505), .A(n7069), .B(n7068), .ZN(n7070)
         );
  OAI21_X1 U8257 ( .B1(n7071), .B2(n9569), .A(n7070), .ZN(P1_U3225) );
  INV_X1 U8258 ( .A(n7072), .ZN(n7081) );
  NOR2_X1 U8259 ( .A1(n10259), .A2(n10666), .ZN(n7074) );
  NAND3_X1 U8260 ( .A1(n7075), .A2(n7074), .A3(n7073), .ZN(n7605) );
  INV_X1 U8261 ( .A(n10090), .ZN(n10139) );
  AOI22_X1 U8262 ( .A1(n10141), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n10139), .ZN(n7080) );
  NOR2_X1 U8263 ( .A1(n7293), .A2(n9823), .ZN(n7077) );
  NOR2_X1 U8264 ( .A1(n7293), .A2(n9828), .ZN(n7078) );
  OAI21_X1 U8265 ( .B1(n10095), .B2(n10115), .A(n7296), .ZN(n7079) );
  OAI211_X1 U8266 ( .C1(n7081), .C2(n10141), .A(n7080), .B(n7079), .ZN(
        P1_U3291) );
  OAI21_X1 U8267 ( .B1(n7084), .B2(n7083), .A(n7082), .ZN(n7093) );
  INV_X1 U8268 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7087) );
  NAND2_X1 U8269 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8139) );
  OR2_X1 U8270 ( .A1(n9899), .A2(n7085), .ZN(n7086) );
  OAI211_X1 U8271 ( .C1(n9884), .C2(n7087), .A(n8139), .B(n7086), .ZN(n7092)
         );
  AOI211_X1 U8272 ( .C1(n7090), .C2(n7089), .A(n7088), .B(n9869), .ZN(n7091)
         );
  AOI211_X1 U8273 ( .C1(n10745), .C2(n7093), .A(n7092), .B(n7091), .ZN(n7094)
         );
  INV_X1 U8274 ( .A(n7094), .ZN(P1_U3254) );
  NAND2_X1 U8275 ( .A1(n8996), .A2(n8535), .ZN(n7102) );
  OR2_X1 U8276 ( .A1(n5039), .A2(n6866), .ZN(n7097) );
  OR2_X1 U8277 ( .A1(n5037), .A2(n7095), .ZN(n7096) );
  OAI211_X1 U8278 ( .C1(n7537), .C2(n7098), .A(n7097), .B(n7096), .ZN(n7365)
         );
  XNOR2_X1 U8279 ( .A(n8551), .B(n7365), .ZN(n7101) );
  XNOR2_X1 U8280 ( .A(n7102), .B(n7101), .ZN(n7360) );
  INV_X1 U8281 ( .A(n7101), .ZN(n7131) );
  NAND2_X1 U8282 ( .A1(n7131), .A2(n7102), .ZN(n7117) );
  OR2_X1 U8283 ( .A1(n5037), .A2(n7103), .ZN(n7109) );
  OR2_X1 U8284 ( .A1(n5039), .A2(n7105), .ZN(n7108) );
  OR2_X1 U8285 ( .A1(n7537), .A2(n7106), .ZN(n7107) );
  XNOR2_X1 U8286 ( .A(n10898), .B(n8551), .ZN(n7383) );
  NAND2_X1 U8287 ( .A1(n8047), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7116) );
  NAND2_X1 U8288 ( .A1(n7110), .A2(n10459), .ZN(n7111) );
  NAND2_X1 U8289 ( .A1(n7119), .A2(n7111), .ZN(n7435) );
  OR2_X1 U8290 ( .A1(n8321), .A2(n7435), .ZN(n7115) );
  OR2_X1 U8291 ( .A1(n8324), .A2(n7112), .ZN(n7114) );
  INV_X1 U8292 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7436) );
  OR2_X1 U8293 ( .A1(n8253), .A2(n7436), .ZN(n7113) );
  NAND4_X1 U8294 ( .A1(n7116), .A2(n7115), .A3(n7114), .A4(n7113), .ZN(n8995)
         );
  NAND2_X1 U8295 ( .A1(n8995), .A2(n8535), .ZN(n7372) );
  XNOR2_X1 U8296 ( .A(n7383), .B(n7372), .ZN(n7133) );
  AOI21_X1 U8297 ( .B1(n7357), .B2(n7117), .A(n7133), .ZN(n7374) );
  INV_X1 U8298 ( .A(n7374), .ZN(n7387) );
  INV_X1 U8299 ( .A(n10898), .ZN(n7438) );
  NAND2_X1 U8300 ( .A1(n7118), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7125) );
  NAND2_X1 U8301 ( .A1(n7119), .A2(n10539), .ZN(n7120) );
  NAND2_X1 U8302 ( .A1(n7318), .A2(n7120), .ZN(n7381) );
  OR2_X1 U8303 ( .A1(n8321), .A2(n7381), .ZN(n7124) );
  OR2_X1 U8304 ( .A1(n8324), .A2(n7121), .ZN(n7123) );
  INV_X1 U8305 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7336) );
  OR2_X1 U8306 ( .A1(n8253), .A2(n7336), .ZN(n7122) );
  NAND4_X1 U8307 ( .A1(n7125), .A2(n7124), .A3(n7123), .A4(n7122), .ZN(n8994)
         );
  INV_X1 U8308 ( .A(n8994), .ZN(n7445) );
  INV_X1 U8309 ( .A(n8930), .ZN(n8966) );
  NAND2_X1 U8310 ( .A1(n8966), .A2(n8996), .ZN(n7128) );
  INV_X1 U8311 ( .A(n7126), .ZN(n7127) );
  OAI211_X1 U8312 ( .C1(n7445), .C2(n8964), .A(n7128), .B(n7127), .ZN(n7130)
         );
  NOR2_X1 U8313 ( .A1(n8968), .A2(n7435), .ZN(n7129) );
  AOI211_X1 U8314 ( .C1(n7438), .C2(n8975), .A(n7130), .B(n7129), .ZN(n7135)
         );
  INV_X1 U8315 ( .A(n8996), .ZN(n7339) );
  OAI22_X1 U8316 ( .A1(n7339), .A2(n8922), .B1(n7131), .B2(n8953), .ZN(n7132)
         );
  NAND3_X1 U8317 ( .A1(n7357), .A2(n7133), .A3(n7132), .ZN(n7134) );
  OAI211_X1 U8318 ( .C1(n7387), .C2(n8953), .A(n7135), .B(n7134), .ZN(P2_U3229) );
  OAI21_X1 U8319 ( .B1(n7138), .B2(n7137), .A(n7136), .ZN(n7139) );
  INV_X1 U8320 ( .A(n7139), .ZN(n7150) );
  OAI21_X1 U8321 ( .B1(n7142), .B2(n7141), .A(n7140), .ZN(n7148) );
  INV_X1 U8322 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7146) );
  NOR2_X1 U8323 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7143), .ZN(n9431) );
  AOI21_X1 U8324 ( .B1(n10760), .B2(n7144), .A(n9431), .ZN(n7145) );
  OAI21_X1 U8325 ( .B1(n7146), .B2(n9884), .A(n7145), .ZN(n7147) );
  AOI21_X1 U8326 ( .B1(n7148), .B2(n10745), .A(n7147), .ZN(n7149) );
  OAI21_X1 U8327 ( .B1(n7150), .B2(n9869), .A(n7149), .ZN(P1_U3255) );
  AOI21_X1 U8328 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n7538), .A(n7151), .ZN(
        n7154) );
  NAND2_X1 U8329 ( .A1(n7749), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7152) );
  OAI21_X1 U8330 ( .B1(n7749), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7152), .ZN(
        n7153) );
  NOR2_X1 U8331 ( .A1(n7154), .A2(n7153), .ZN(n7620) );
  AOI211_X1 U8332 ( .C1(n7154), .C2(n7153), .A(n7620), .B(n10801), .ZN(n7164)
         );
  OAI21_X1 U8333 ( .B1(n7156), .B2(n7528), .A(n7155), .ZN(n7159) );
  MUX2_X1 U8334 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7157), .S(n7749), .Z(n7158)
         );
  NAND2_X1 U8335 ( .A1(n7158), .A2(n7159), .ZN(n7612) );
  OAI211_X1 U8336 ( .C1(n7159), .C2(n7158), .A(n10809), .B(n7612), .ZN(n7162)
         );
  NOR2_X1 U8337 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10527), .ZN(n7160) );
  AOI21_X1 U8338 ( .B1(n10800), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7160), .ZN(
        n7161) );
  OAI211_X1 U8339 ( .C1(n10792), .C2(n7613), .A(n7162), .B(n7161), .ZN(n7163)
         );
  OR2_X1 U8340 ( .A1(n7164), .A2(n7163), .ZN(P2_U3255) );
  XNOR2_X1 U8341 ( .A(n7167), .B(n7166), .ZN(n7168) );
  XNOR2_X1 U8342 ( .A(n7165), .B(n7168), .ZN(n7175) );
  INV_X1 U8343 ( .A(n7517), .ZN(n7173) );
  NOR2_X1 U8344 ( .A1(n9535), .A2(n7571), .ZN(n7172) );
  INV_X1 U8345 ( .A(n9847), .ZN(n7561) );
  NAND2_X1 U8346 ( .A1(n9561), .A2(n9849), .ZN(n7170) );
  OAI211_X1 U8347 ( .C1(n7561), .C2(n9559), .A(n7170), .B(n7169), .ZN(n7171)
         );
  AOI211_X1 U8348 ( .C1(n7173), .C2(n9505), .A(n7172), .B(n7171), .ZN(n7174)
         );
  OAI21_X1 U8349 ( .B1(n7175), .B2(n9569), .A(n7174), .ZN(P1_U3237) );
  NAND2_X1 U8350 ( .A1(n8801), .A2(n7176), .ZN(n7177) );
  INV_X1 U8351 ( .A(n7207), .ZN(n7179) );
  NAND2_X1 U8352 ( .A1(n7179), .A2(n7209), .ZN(n7303) );
  INV_X1 U8353 ( .A(n8998), .ZN(n7187) );
  NAND2_X1 U8354 ( .A1(n7187), .A2(n10864), .ZN(n7302) );
  NAND2_X1 U8355 ( .A1(n7303), .A2(n7302), .ZN(n7180) );
  NAND2_X1 U8356 ( .A1(n7192), .A2(n7315), .ZN(n8633) );
  INV_X1 U8357 ( .A(n7192), .ZN(n8997) );
  NAND2_X1 U8358 ( .A1(n8997), .A2(n10877), .ZN(n8634) );
  INV_X1 U8359 ( .A(n8629), .ZN(n8765) );
  NAND2_X1 U8360 ( .A1(n7180), .A2(n8765), .ZN(n7309) );
  NAND2_X1 U8361 ( .A1(n7192), .A2(n10877), .ZN(n7181) );
  NAND2_X1 U8362 ( .A1(n7309), .A2(n7181), .ZN(n7182) );
  XNOR2_X1 U8363 ( .A(n8996), .B(n7365), .ZN(n8768) );
  INV_X1 U8364 ( .A(n8768), .ZN(n7190) );
  NAND2_X1 U8365 ( .A1(n7182), .A2(n7190), .ZN(n7341) );
  OAI21_X1 U8366 ( .B1(n7182), .B2(n7190), .A(n7341), .ZN(n7349) );
  INV_X1 U8367 ( .A(n10848), .ZN(n7215) );
  INV_X1 U8368 ( .A(n7365), .ZN(n8638) );
  NOR2_X1 U8369 ( .A1(n7310), .A2(n8638), .ZN(n7183) );
  OR2_X1 U8370 ( .A1(n7434), .A2(n7183), .ZN(n7351) );
  OAI22_X1 U8371 ( .A1(n7351), .A2(n10994), .B1(n8638), .B2(n10992), .ZN(n7193) );
  NOR2_X1 U8372 ( .A1(n8811), .A2(n8620), .ZN(n8800) );
  INV_X1 U8373 ( .A(n8800), .ZN(n7184) );
  OR2_X1 U8374 ( .A1(n8801), .A2(n8807), .ZN(n8812) );
  NAND2_X1 U8375 ( .A1(n7221), .A2(n10831), .ZN(n10816) );
  NAND2_X1 U8376 ( .A1(n7391), .A2(n8624), .ZN(n7206) );
  NAND2_X1 U8377 ( .A1(n7187), .A2(n7186), .ZN(n7188) );
  NAND2_X1 U8378 ( .A1(n8632), .A2(n8629), .ZN(n7189) );
  NAND2_X1 U8379 ( .A1(n7189), .A2(n8633), .ZN(n7331) );
  XNOR2_X1 U8380 ( .A(n7331), .B(n7190), .ZN(n7191) );
  OAI222_X1 U8381 ( .A1(n9270), .A2(n7384), .B1(n9272), .B2(n7192), .C1(n9264), 
        .C2(n7191), .ZN(n7350) );
  AOI211_X1 U8382 ( .C1(n10980), .C2(n7349), .A(n7193), .B(n7350), .ZN(n7238)
         );
  INV_X1 U8383 ( .A(n7194), .ZN(n7232) );
  NAND2_X1 U8384 ( .A1(n11000), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7196) );
  OAI21_X1 U8385 ( .B1(n7238), .B2(n11000), .A(n7196), .ZN(P2_U3524) );
  AOI21_X1 U8386 ( .B1(n7198), .B2(n8535), .A(n8953), .ZN(n7197) );
  OAI21_X1 U8387 ( .B1(n7197), .B2(n8975), .A(n10831), .ZN(n7202) );
  NAND2_X1 U8388 ( .A1(n7198), .A2(n10817), .ZN(n10815) );
  INV_X1 U8389 ( .A(n10815), .ZN(n7200) );
  AOI22_X1 U8390 ( .A1(n8840), .A2(n7200), .B1(n8960), .B2(n10820), .ZN(n7201)
         );
  OAI211_X1 U8391 ( .C1(n7225), .C2(n10824), .A(n7202), .B(n7201), .ZN(
        P2_U3234) );
  NOR2_X1 U8392 ( .A1(n7231), .A2(n7203), .ZN(n7204) );
  NAND2_X1 U8393 ( .A1(n7237), .A2(n7204), .ZN(n7214) );
  NAND2_X1 U8394 ( .A1(n7206), .A2(n10822), .ZN(n7211) );
  INV_X1 U8395 ( .A(n7206), .ZN(n7208) );
  AOI22_X1 U8396 ( .A1(n7208), .A2(n10822), .B1(n7207), .B2(n10980), .ZN(n7210) );
  INV_X1 U8397 ( .A(n7209), .ZN(n8769) );
  MUX2_X1 U8398 ( .A(n7211), .B(n7210), .S(n8769), .Z(n7213) );
  AOI22_X1 U8399 ( .A1(n10821), .A2(n8997), .B1(n10820), .B2(n9254), .ZN(n7212) );
  OAI211_X1 U8400 ( .C1(n10990), .C2(n7303), .A(n7213), .B(n7212), .ZN(n10867)
         );
  NAND2_X1 U8401 ( .A1(n10867), .A2(n10829), .ZN(n7218) );
  OAI21_X1 U8402 ( .B1(n7215), .B2(n10864), .A(n7311), .ZN(n10865) );
  OAI22_X1 U8403 ( .A1(n10818), .A2(n10865), .B1(n10451), .B2(n10823), .ZN(
        n7216) );
  AOI21_X1 U8404 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n9303), .A(n7216), .ZN(
        n7217) );
  OAI211_X1 U8405 ( .C1(n10864), .C2(n10819), .A(n7218), .B(n7217), .ZN(
        P2_U3294) );
  OAI21_X1 U8406 ( .B1(n7220), .B2(n7226), .A(n7219), .ZN(n7229) );
  OR2_X1 U8407 ( .A1(n7221), .A2(n9272), .ZN(n7223) );
  NAND2_X1 U8408 ( .A1(n8998), .A2(n10821), .ZN(n7222) );
  NAND2_X1 U8409 ( .A1(n7223), .A2(n7222), .ZN(n7394) );
  INV_X1 U8410 ( .A(n7845), .ZN(n8882) );
  AOI22_X1 U8411 ( .A1(n8975), .A2(n7400), .B1(n7394), .B2(n8882), .ZN(n7224)
         );
  OAI21_X1 U8412 ( .B1(n7225), .B2(n10785), .A(n7224), .ZN(n7228) );
  NOR3_X1 U8413 ( .A1(n7226), .A2(n7398), .A3(n8922), .ZN(n7227) );
  AOI211_X1 U8414 ( .C1(n8915), .C2(n7229), .A(n7228), .B(n7227), .ZN(n7230)
         );
  INV_X1 U8415 ( .A(n7230), .ZN(P2_U3224) );
  INV_X1 U8416 ( .A(n7231), .ZN(n7233) );
  AND4_X1 U8417 ( .A1(n7235), .A2(n7234), .A3(n7233), .A4(n7232), .ZN(n7236)
         );
  INV_X1 U8418 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7240) );
  OR2_X1 U8419 ( .A1(n7238), .A2(n11003), .ZN(n7239) );
  OAI21_X1 U8420 ( .B1(n11006), .B2(n7240), .A(n7239), .ZN(P2_U3463) );
  NAND2_X1 U8421 ( .A1(n6891), .A2(n7296), .ZN(n7286) );
  INV_X1 U8422 ( .A(n7286), .ZN(n7243) );
  NAND2_X1 U8423 ( .A1(n7256), .A2(n9593), .ZN(n7242) );
  NAND2_X1 U8424 ( .A1(n7272), .A2(n9764), .ZN(n7245) );
  NAND2_X1 U8425 ( .A1(n7258), .A2(n10857), .ZN(n7244) );
  NAND2_X1 U8426 ( .A1(n7245), .A2(n7244), .ZN(n7408) );
  INV_X1 U8427 ( .A(n9762), .ZN(n7247) );
  XNOR2_X1 U8428 ( .A(n7408), .B(n7247), .ZN(n7268) );
  INV_X1 U8429 ( .A(n7268), .ZN(n10874) );
  NOR2_X1 U8430 ( .A1(n7248), .A2(n10030), .ZN(n7249) );
  NAND2_X1 U8431 ( .A1(n10093), .A2(n7249), .ZN(n10055) );
  INV_X1 U8432 ( .A(n10055), .ZN(n10121) );
  NAND2_X1 U8433 ( .A1(n9594), .A2(n9593), .ZN(n7294) );
  INV_X1 U8434 ( .A(n7412), .ZN(n7252) );
  INV_X1 U8435 ( .A(n7273), .ZN(n7250) );
  NAND2_X1 U8436 ( .A1(n7250), .A2(n7414), .ZN(n7251) );
  NAND2_X1 U8437 ( .A1(n7252), .A2(n7251), .ZN(n10871) );
  INV_X1 U8438 ( .A(n10115), .ZN(n10098) );
  AOI22_X1 U8439 ( .A1(n10095), .A2(n7414), .B1(n7253), .B2(n10139), .ZN(n7254) );
  OAI21_X1 U8440 ( .B1(n10871), .B2(n10098), .A(n7254), .ZN(n7270) );
  NOR2_X1 U8441 ( .A1(n6891), .A2(n9594), .ZN(n7291) );
  NAND2_X1 U8442 ( .A1(n7256), .A2(n10839), .ZN(n7257) );
  AND2_X2 U8443 ( .A1(n7290), .A2(n7257), .ZN(n7276) );
  NAND2_X1 U8444 ( .A1(n7258), .A2(n7274), .ZN(n7259) );
  NAND2_X1 U8445 ( .A1(n9850), .A2(n10857), .ZN(n9598) );
  NAND2_X1 U8446 ( .A1(n7260), .A2(n9762), .ZN(n7261) );
  NAND2_X1 U8447 ( .A1(n7416), .A2(n7261), .ZN(n7264) );
  NAND2_X1 U8448 ( .A1(n7262), .A2(n10659), .ZN(n7263) );
  OR2_X1 U8449 ( .A1(n5762), .A2(n9823), .ZN(n9818) );
  NAND2_X2 U8450 ( .A1(n7263), .A2(n9818), .ZN(n10125) );
  NAND2_X1 U8451 ( .A1(n7264), .A2(n10125), .ZN(n7267) );
  AOI22_X1 U8452 ( .A1(n10131), .A2(n9850), .B1(n5875), .B2(n10130), .ZN(n7266) );
  OAI211_X1 U8453 ( .C1(n7268), .C2(n7255), .A(n7267), .B(n7266), .ZN(n10872)
         );
  MUX2_X1 U8454 ( .A(n10872), .B(P1_REG2_REG_3__SCAN_IN), .S(n10141), .Z(n7269) );
  AOI211_X1 U8455 ( .C1(n10874), .C2(n10121), .A(n7270), .B(n7269), .ZN(n7271)
         );
  INV_X1 U8456 ( .A(n7271), .ZN(P1_U3288) );
  XNOR2_X1 U8457 ( .A(n7272), .B(n9764), .ZN(n10861) );
  AOI21_X1 U8458 ( .B1(n7274), .B2(n7294), .A(n7273), .ZN(n10856) );
  AOI22_X1 U8459 ( .A1(n10856), .A2(n10115), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n10139), .ZN(n7275) );
  OAI21_X1 U8460 ( .B1(n10857), .B2(n10144), .A(n7275), .ZN(n7282) );
  XNOR2_X1 U8461 ( .A(n7276), .B(n9764), .ZN(n7277) );
  NAND2_X1 U8462 ( .A1(n7277), .A2(n10125), .ZN(n7280) );
  INV_X1 U8463 ( .A(n7255), .ZN(n10929) );
  NAND2_X1 U8464 ( .A1(n10861), .A2(n10929), .ZN(n7279) );
  AOI22_X1 U8465 ( .A1(n10130), .A2(n7246), .B1(n9851), .B2(n10131), .ZN(n7278) );
  NAND3_X1 U8466 ( .A1(n7280), .A2(n7279), .A3(n7278), .ZN(n10859) );
  MUX2_X1 U8467 ( .A(n10859), .B(P1_REG2_REG_2__SCAN_IN), .S(n10141), .Z(n7281) );
  AOI211_X1 U8468 ( .C1(n10861), .C2(n10121), .A(n7282), .B(n7281), .ZN(n7283)
         );
  INV_X1 U8469 ( .A(n7283), .ZN(P1_U3289) );
  XNOR2_X1 U8470 ( .A(n7285), .B(n7286), .ZN(n10844) );
  AND2_X1 U8471 ( .A1(n7288), .A2(n7287), .ZN(n7289) );
  INV_X1 U8472 ( .A(n10148), .ZN(n9929) );
  OAI22_X1 U8473 ( .A1(n10144), .A2(n9593), .B1(n6600), .B2(n10093), .ZN(n7299) );
  OAI21_X1 U8474 ( .B1(n7284), .B2(n7291), .A(n7290), .ZN(n7292) );
  AOI222_X1 U8475 ( .A1(n10125), .A2(n7292), .B1(n9850), .B2(n10130), .C1(
        n6891), .C2(n10131), .ZN(n10841) );
  INV_X1 U8476 ( .A(n7294), .ZN(n7295) );
  AOI211_X1 U8477 ( .C1(n7296), .C2(n10839), .A(n11009), .B(n7295), .ZN(n10838) );
  AOI22_X1 U8478 ( .A1(n10838), .A2(n10030), .B1(n10139), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7297) );
  AOI21_X1 U8479 ( .B1(n10841), .B2(n7297), .A(n10141), .ZN(n7298) );
  AOI211_X1 U8480 ( .C1(n10844), .C2(n9929), .A(n7299), .B(n7298), .ZN(n7300)
         );
  INV_X1 U8481 ( .A(n7300), .ZN(P1_U3290) );
  INV_X1 U8482 ( .A(n8632), .ZN(n7301) );
  NAND2_X1 U8483 ( .A1(n7301), .A2(n10822), .ZN(n7306) );
  AND3_X1 U8484 ( .A1(n7303), .A2(n10980), .A3(n7302), .ZN(n7304) );
  AOI21_X1 U8485 ( .B1(n8632), .B2(n10822), .A(n7304), .ZN(n7305) );
  MUX2_X1 U8486 ( .A(n7306), .B(n7305), .S(n8629), .Z(n7308) );
  OAI211_X1 U8487 ( .C1(n10990), .C2(n7309), .A(n7308), .B(n7307), .ZN(n10878)
         );
  INV_X1 U8488 ( .A(n10878), .ZN(n7317) );
  AOI21_X1 U8489 ( .B1(n7315), .B2(n7311), .A(n7310), .ZN(n10880) );
  INV_X1 U8490 ( .A(n10823), .ZN(n9202) );
  AOI22_X1 U8491 ( .A1(n10880), .A2(n9226), .B1(n9202), .B2(n10525), .ZN(n7312) );
  OAI21_X1 U8492 ( .B1(n7313), .B2(n10829), .A(n7312), .ZN(n7314) );
  AOI21_X1 U8493 ( .B1(n9292), .B2(n7315), .A(n7314), .ZN(n7316) );
  OAI21_X1 U8494 ( .B1(n7317), .B2(n9303), .A(n7316), .ZN(P2_U3293) );
  NAND2_X1 U8495 ( .A1(n8047), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7324) );
  NAND2_X1 U8496 ( .A1(n7318), .A2(n10514), .ZN(n7319) );
  NAND2_X1 U8497 ( .A1(n7529), .A2(n7319), .ZN(n7495) );
  OR2_X1 U8498 ( .A1(n8321), .A2(n7495), .ZN(n7323) );
  OR2_X1 U8499 ( .A1(n8324), .A2(n7320), .ZN(n7322) );
  OR2_X1 U8500 ( .A1(n8253), .A2(n6840), .ZN(n7321) );
  NAND4_X1 U8501 ( .A1(n7324), .A2(n7323), .A3(n7322), .A4(n7321), .ZN(n8993)
         );
  INV_X1 U8502 ( .A(n8993), .ZN(n8656) );
  OR2_X1 U8503 ( .A1(n5037), .A2(n7325), .ZN(n7330) );
  OR2_X1 U8504 ( .A1(n5039), .A2(n7326), .ZN(n7329) );
  OR2_X1 U8505 ( .A1(n7537), .A2(n7327), .ZN(n7328) );
  NAND2_X1 U8506 ( .A1(n7445), .A2(n10912), .ZN(n8651) );
  NAND2_X1 U8507 ( .A1(n8994), .A2(n8648), .ZN(n8650) );
  NAND2_X1 U8508 ( .A1(n8651), .A2(n8650), .ZN(n8770) );
  NAND2_X1 U8509 ( .A1(n7331), .A2(n8768), .ZN(n7332) );
  NAND2_X1 U8510 ( .A1(n7339), .A2(n7365), .ZN(n8640) );
  NAND2_X1 U8511 ( .A1(n8995), .A2(n10898), .ZN(n8645) );
  NAND2_X1 U8512 ( .A1(n7443), .A2(n8645), .ZN(n7333) );
  NAND2_X1 U8513 ( .A1(n7384), .A2(n7438), .ZN(n8644) );
  NAND2_X1 U8514 ( .A1(n7333), .A2(n8644), .ZN(n7334) );
  XOR2_X1 U8515 ( .A(n8770), .B(n7334), .Z(n7335) );
  OAI222_X1 U8516 ( .A1(n9270), .A2(n8656), .B1(n9272), .B2(n7384), .C1(n9264), 
        .C2(n7335), .ZN(n10914) );
  INV_X1 U8517 ( .A(n10914), .ZN(n7348) );
  OAI22_X1 U8518 ( .A1(n10829), .A2(n7336), .B1(n7381), .B2(n10823), .ZN(n7338) );
  XNOR2_X1 U8519 ( .A(n7463), .B(n8648), .ZN(n10913) );
  NOR2_X1 U8520 ( .A1(n10913), .A2(n10818), .ZN(n7337) );
  AOI211_X1 U8521 ( .C1(n9292), .C2(n8648), .A(n7338), .B(n7337), .ZN(n7347)
         );
  NAND2_X1 U8522 ( .A1(n7339), .A2(n8638), .ZN(n7340) );
  NAND2_X1 U8523 ( .A1(n7341), .A2(n7340), .ZN(n7433) );
  NAND2_X1 U8524 ( .A1(n8644), .A2(n8645), .ZN(n8766) );
  NAND2_X1 U8525 ( .A1(n7433), .A2(n8766), .ZN(n7343) );
  NAND2_X1 U8526 ( .A1(n7384), .A2(n10898), .ZN(n7342) );
  NAND2_X1 U8527 ( .A1(n7343), .A2(n7342), .ZN(n7344) );
  AND2_X1 U8528 ( .A1(n7344), .A2(n8770), .ZN(n10911) );
  INV_X1 U8529 ( .A(n10911), .ZN(n7345) );
  OR2_X2 U8530 ( .A1(n7344), .A2(n8770), .ZN(n7461) );
  NAND3_X1 U8531 ( .A1(n7345), .A2(n10827), .A3(n10916), .ZN(n7346) );
  OAI211_X1 U8532 ( .C1(n7348), .C2(n9303), .A(n7347), .B(n7346), .ZN(P2_U3290) );
  INV_X1 U8533 ( .A(n7349), .ZN(n7356) );
  NAND2_X1 U8534 ( .A1(n7350), .A2(n10829), .ZN(n7355) );
  OAI22_X1 U8535 ( .A1(n10829), .A2(n6583), .B1(n7368), .B2(n10823), .ZN(n7353) );
  NOR2_X1 U8536 ( .A1(n7351), .A2(n10818), .ZN(n7352) );
  AOI211_X1 U8537 ( .C1(n9292), .C2(n7365), .A(n7353), .B(n7352), .ZN(n7354)
         );
  OAI211_X1 U8538 ( .C1(n7356), .C2(n9300), .A(n7355), .B(n7354), .ZN(P2_U3292) );
  OAI21_X1 U8539 ( .B1(n7360), .B2(n7358), .A(n7357), .ZN(n7370) );
  NOR3_X1 U8540 ( .A1(n7360), .A2(n7359), .A3(n8922), .ZN(n7361) );
  OAI21_X1 U8541 ( .B1(n7361), .B2(n8966), .A(n8997), .ZN(n7367) );
  INV_X1 U8542 ( .A(n7362), .ZN(n7363) );
  OAI21_X1 U8543 ( .B1(n8964), .B2(n7384), .A(n7363), .ZN(n7364) );
  AOI21_X1 U8544 ( .B1(n8975), .B2(n7365), .A(n7364), .ZN(n7366) );
  OAI211_X1 U8545 ( .C1(n8968), .C2(n7368), .A(n7367), .B(n7366), .ZN(n7369)
         );
  AOI21_X1 U8546 ( .B1(n7370), .B2(n8915), .A(n7369), .ZN(n7371) );
  INV_X1 U8547 ( .A(n7371), .ZN(P2_U3232) );
  XNOR2_X1 U8548 ( .A(n10912), .B(n8551), .ZN(n7489) );
  NAND2_X1 U8549 ( .A1(n8994), .A2(n8535), .ZN(n7490) );
  XNOR2_X1 U8550 ( .A(n7489), .B(n7490), .ZN(n7386) );
  INV_X1 U8551 ( .A(n7386), .ZN(n7375) );
  INV_X1 U8552 ( .A(n7491), .ZN(n7390) );
  INV_X1 U8553 ( .A(n7377), .ZN(n7378) );
  OAI21_X1 U8554 ( .B1(n8930), .B2(n7384), .A(n7378), .ZN(n7379) );
  AOI21_X1 U8555 ( .B1(n8960), .B2(n8993), .A(n7379), .ZN(n7380) );
  OAI21_X1 U8556 ( .B1(n7381), .B2(n8968), .A(n7380), .ZN(n7382) );
  AOI21_X1 U8557 ( .B1(n8648), .B2(n8975), .A(n7382), .ZN(n7389) );
  OAI22_X1 U8558 ( .A1(n8922), .A2(n7384), .B1(n7383), .B2(n8953), .ZN(n7385)
         );
  NAND3_X1 U8559 ( .A1(n7387), .A2(n7386), .A3(n7385), .ZN(n7388) );
  OAI211_X1 U8560 ( .C1(n7390), .C2(n8953), .A(n7389), .B(n7388), .ZN(P2_U3241) );
  INV_X1 U8561 ( .A(n7391), .ZN(n8627) );
  INV_X1 U8562 ( .A(n8623), .ZN(n7396) );
  NAND2_X1 U8563 ( .A1(n7392), .A2(n8624), .ZN(n7399) );
  INV_X1 U8564 ( .A(n10816), .ZN(n7393) );
  AOI21_X1 U8565 ( .B1(n7399), .B2(n7393), .A(n9264), .ZN(n7395) );
  AOI21_X1 U8566 ( .B1(n7396), .B2(n7395), .A(n7394), .ZN(n10850) );
  INV_X1 U8567 ( .A(n10850), .ZN(n7397) );
  AOI21_X1 U8568 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n9202), .A(n7397), .ZN(
        n7405) );
  XNOR2_X1 U8569 ( .A(n7399), .B(n7398), .ZN(n10853) );
  NAND2_X1 U8570 ( .A1(n7400), .A2(n10831), .ZN(n10847) );
  NAND3_X1 U8571 ( .A1(n9226), .A2(n10848), .A3(n10847), .ZN(n7402) );
  NAND2_X1 U8572 ( .A1(n9303), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7401) );
  OAI211_X1 U8573 ( .C1(n10819), .C2(n10851), .A(n7402), .B(n7401), .ZN(n7403)
         );
  AOI21_X1 U8574 ( .B1(n10827), .B2(n10853), .A(n7403), .ZN(n7404) );
  OAI21_X1 U8575 ( .B1(n7405), .B2(n9303), .A(n7404), .ZN(P2_U3295) );
  INV_X1 U8576 ( .A(n8222), .ZN(n7407) );
  OAI222_X1 U8577 ( .A1(n9873), .A2(P1_U3084), .B1(n10265), .B2(n7407), .C1(
        n10571), .C2(n10267), .ZN(P1_U3335) );
  XNOR2_X1 U8578 ( .A(n7406), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9073) );
  INV_X1 U8579 ( .A(n9073), .ZN(n9081) );
  OAI222_X1 U8580 ( .A1(n9081), .A2(P2_U3152), .B1(n8494), .B2(n7407), .C1(
        n5036), .C2(n6175), .ZN(P2_U3340) );
  NAND2_X1 U8581 ( .A1(n7408), .A2(n9762), .ZN(n7410) );
  INV_X1 U8582 ( .A(n7246), .ZN(n7415) );
  NAND2_X1 U8583 ( .A1(n7415), .A2(n10870), .ZN(n7409) );
  NAND2_X1 U8584 ( .A1(n7410), .A2(n7409), .ZN(n7480) );
  XNOR2_X1 U8585 ( .A(n5875), .B(n7411), .ZN(n7479) );
  INV_X1 U8586 ( .A(n7479), .ZN(n9765) );
  XNOR2_X1 U8587 ( .A(n7480), .B(n9765), .ZN(n7420) );
  INV_X1 U8588 ( .A(n7420), .ZN(n10887) );
  OAI21_X1 U8589 ( .B1(n7412), .B2(n7411), .A(n7471), .ZN(n10884) );
  AOI22_X1 U8590 ( .A1(n10095), .A2(n5871), .B1(n10139), .B2(n8386), .ZN(n7413) );
  OAI21_X1 U8591 ( .B1(n10884), .B2(n10098), .A(n7413), .ZN(n7422) );
  NAND2_X1 U8592 ( .A1(n7415), .A2(n7414), .ZN(n9602) );
  XNOR2_X1 U8593 ( .A(n7473), .B(n9765), .ZN(n7417) );
  NAND2_X1 U8594 ( .A1(n7417), .A2(n10125), .ZN(n7419) );
  AOI22_X1 U8595 ( .A1(n10131), .A2(n7246), .B1(n9849), .B2(n10130), .ZN(n7418) );
  OAI211_X1 U8596 ( .C1(n7420), .C2(n7255), .A(n7419), .B(n7418), .ZN(n10885)
         );
  MUX2_X1 U8597 ( .A(n10885), .B(P1_REG2_REG_4__SCAN_IN), .S(n10141), .Z(n7421) );
  AOI211_X1 U8598 ( .C1(n10887), .C2(n10121), .A(n7422), .B(n7421), .ZN(n7423)
         );
  INV_X1 U8599 ( .A(n7423), .ZN(P1_U3287) );
  XOR2_X1 U8600 ( .A(n7425), .B(n7424), .Z(n7431) );
  NOR2_X1 U8601 ( .A1(n9535), .A2(n7608), .ZN(n7429) );
  NAND2_X1 U8602 ( .A1(n9561), .A2(n9848), .ZN(n7427) );
  OAI211_X1 U8603 ( .C1(n7564), .C2(n9559), .A(n7427), .B(n7426), .ZN(n7428)
         );
  AOI211_X1 U8604 ( .C1(n7606), .C2(n9505), .A(n7429), .B(n7428), .ZN(n7430)
         );
  OAI21_X1 U8605 ( .B1(n7431), .B2(n9569), .A(n7430), .ZN(P1_U3211) );
  INV_X1 U8606 ( .A(n8766), .ZN(n8642) );
  XNOR2_X1 U8607 ( .A(n7443), .B(n8642), .ZN(n7432) );
  AOI222_X1 U8608 ( .A1(n10822), .A2(n7432), .B1(n8994), .B2(n10821), .C1(
        n8996), .C2(n9254), .ZN(n10897) );
  XNOR2_X1 U8609 ( .A(n7433), .B(n8766), .ZN(n10900) );
  OAI211_X1 U8610 ( .C1(n7434), .C2(n10898), .A(n10881), .B(n7463), .ZN(n10896) );
  NAND2_X1 U8611 ( .A1(n10829), .A2(n8811), .ZN(n9280) );
  OAI22_X1 U8612 ( .A1(n10829), .A2(n7436), .B1(n7435), .B2(n10823), .ZN(n7437) );
  AOI21_X1 U8613 ( .B1(n9292), .B2(n7438), .A(n7437), .ZN(n7439) );
  OAI21_X1 U8614 ( .B1(n10896), .B2(n9280), .A(n7439), .ZN(n7440) );
  AOI21_X1 U8615 ( .B1(n10900), .B2(n10827), .A(n7440), .ZN(n7441) );
  OAI21_X1 U8616 ( .B1(n10897), .B2(n9303), .A(n7441), .ZN(P2_U3291) );
  NAND2_X1 U8617 ( .A1(n8994), .A2(n10912), .ZN(n7444) );
  AND2_X1 U8618 ( .A1(n8645), .A2(n7444), .ZN(n7442) );
  OR2_X1 U8619 ( .A1(n5037), .A2(n7447), .ZN(n7452) );
  OR2_X1 U8620 ( .A1(n5039), .A2(n7448), .ZN(n7451) );
  OR2_X1 U8621 ( .A1(n7537), .A2(n7449), .ZN(n7450) );
  XNOR2_X1 U8622 ( .A(n8993), .B(n10931), .ZN(n8775) );
  OAI211_X1 U8623 ( .C1(n5126), .C2(n5472), .A(n7547), .B(n10822), .ZN(n7459)
         );
  NAND2_X1 U8624 ( .A1(n8047), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7457) );
  OR2_X1 U8625 ( .A1(n8253), .A2(n6944), .ZN(n7456) );
  INV_X1 U8626 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7592) );
  XNOR2_X1 U8627 ( .A(n7529), .B(n7592), .ZN(n7638) );
  OR2_X1 U8628 ( .A1(n8321), .A2(n7638), .ZN(n7455) );
  OR2_X1 U8629 ( .A1(n8324), .A2(n7453), .ZN(n7454) );
  INV_X1 U8630 ( .A(n7711), .ZN(n8992) );
  AOI22_X1 U8631 ( .A1(n8992), .A2(n10821), .B1(n9254), .B2(n8994), .ZN(n7458)
         );
  NAND2_X1 U8632 ( .A1(n7459), .A2(n7458), .ZN(n10933) );
  INV_X1 U8633 ( .A(n10933), .ZN(n7470) );
  AND2_X1 U8634 ( .A1(n10916), .A2(n8650), .ZN(n7462) );
  AND2_X1 U8635 ( .A1(n8775), .A2(n8650), .ZN(n7460) );
  OAI21_X1 U8636 ( .B1(n7462), .B2(n8775), .A(n7522), .ZN(n10935) );
  OR2_X1 U8637 ( .A1(n7463), .A2(n8648), .ZN(n7464) );
  INV_X1 U8638 ( .A(n10931), .ZN(n8657) );
  AND2_X1 U8639 ( .A1(n7464), .A2(n8657), .ZN(n7465) );
  NOR2_X1 U8640 ( .A1(n7464), .A2(n8657), .ZN(n7628) );
  OR2_X1 U8641 ( .A1(n7465), .A2(n7628), .ZN(n10932) );
  OAI22_X1 U8642 ( .A1(n10829), .A2(n6840), .B1(n7495), .B2(n10823), .ZN(n7466) );
  AOI21_X1 U8643 ( .B1(n9292), .B2(n8657), .A(n7466), .ZN(n7467) );
  OAI21_X1 U8644 ( .B1(n10932), .B2(n10818), .A(n7467), .ZN(n7468) );
  AOI21_X1 U8645 ( .B1(n10935), .B2(n10827), .A(n7468), .ZN(n7469) );
  OAI21_X1 U8646 ( .B1(n9303), .B2(n7470), .A(n7469), .ZN(P2_U3289) );
  INV_X1 U8647 ( .A(n7471), .ZN(n7472) );
  INV_X1 U8648 ( .A(n7514), .ZN(n7516) );
  OAI211_X1 U8649 ( .C1(n10890), .C2(n7472), .A(n7516), .B(n11021), .ZN(n10889) );
  NOR2_X1 U8650 ( .A1(n10889), .A2(n10659), .ZN(n7475) );
  NAND2_X1 U8651 ( .A1(n5875), .A2(n7411), .ZN(n9605) );
  NOR2_X1 U8652 ( .A1(n5875), .A2(n7411), .ZN(n9601) );
  INV_X1 U8653 ( .A(n9849), .ZN(n8383) );
  NAND2_X1 U8654 ( .A1(n8383), .A2(n7500), .ZN(n9608) );
  NAND2_X1 U8655 ( .A1(n9849), .A2(n10890), .ZN(n9606) );
  XNOR2_X1 U8656 ( .A(n7507), .B(n9766), .ZN(n7474) );
  OAI222_X1 U8657 ( .A1(n10083), .A2(n7572), .B1(n10081), .B2(n7481), .C1(
        n7474), .C2(n9972), .ZN(n10891) );
  AOI211_X1 U8658 ( .C1(n10139), .C2(n7476), .A(n7475), .B(n10891), .ZN(n7477)
         );
  MUX2_X1 U8659 ( .A(n7478), .B(n7477), .S(n10093), .Z(n7488) );
  NAND2_X1 U8660 ( .A1(n7480), .A2(n7479), .ZN(n7483) );
  NAND2_X1 U8661 ( .A1(n7481), .A2(n7411), .ZN(n7482) );
  INV_X1 U8662 ( .A(n7502), .ZN(n7485) );
  AOI21_X1 U8663 ( .B1(n9766), .B2(n7486), .A(n7485), .ZN(n10893) );
  AOI22_X1 U8664 ( .A1(n10893), .A2(n9929), .B1(n10095), .B2(n7500), .ZN(n7487) );
  NAND2_X1 U8665 ( .A1(n7488), .A2(n7487), .ZN(P1_U3286) );
  XNOR2_X1 U8666 ( .A(n10931), .B(n8551), .ZN(n7580) );
  NAND2_X1 U8667 ( .A1(n8993), .A2(n8535), .ZN(n7492) );
  NOR2_X1 U8668 ( .A1(n7580), .A2(n7492), .ZN(n7585) );
  AOI21_X1 U8669 ( .B1(n7580), .B2(n7492), .A(n7585), .ZN(n7493) );
  OAI211_X1 U8670 ( .C1(n7494), .C2(n7493), .A(n7588), .B(n8915), .ZN(n7499)
         );
  OAI22_X1 U8671 ( .A1(n8964), .A2(n7711), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10514), .ZN(n7497) );
  NOR2_X1 U8672 ( .A1(n8968), .A2(n7495), .ZN(n7496) );
  AOI211_X1 U8673 ( .C1(n8966), .C2(n8994), .A(n7497), .B(n7496), .ZN(n7498)
         );
  OAI211_X1 U8674 ( .C1(n10931), .C2(n8963), .A(n7499), .B(n7498), .ZN(
        P2_U3215) );
  NAND2_X1 U8675 ( .A1(n7572), .A2(n10903), .ZN(n9609) );
  NAND2_X1 U8676 ( .A1(n9848), .A2(n7571), .ZN(n7598) );
  NAND2_X1 U8677 ( .A1(n9849), .A2(n7500), .ZN(n7501) );
  INV_X1 U8678 ( .A(n7506), .ZN(n7504) );
  NAND2_X1 U8679 ( .A1(n7504), .A2(n7503), .ZN(n7574) );
  INV_X1 U8680 ( .A(n7574), .ZN(n7505) );
  AOI21_X1 U8681 ( .B1(n7558), .B2(n7506), .A(n7505), .ZN(n10907) );
  NAND2_X1 U8682 ( .A1(n7507), .A2(n9766), .ZN(n7508) );
  NAND2_X1 U8683 ( .A1(n7508), .A2(n9606), .ZN(n7559) );
  XNOR2_X1 U8684 ( .A(n7509), .B(n7503), .ZN(n7512) );
  AOI22_X1 U8685 ( .A1(n10131), .A2(n9849), .B1(n9847), .B2(n10130), .ZN(n7510) );
  OAI21_X1 U8686 ( .B1(n10907), .B2(n7255), .A(n7510), .ZN(n7511) );
  AOI21_X1 U8687 ( .B1(n10125), .B2(n7512), .A(n7511), .ZN(n10906) );
  MUX2_X1 U8688 ( .A(n7513), .B(n10906), .S(n10093), .Z(n7520) );
  NAND2_X1 U8689 ( .A1(n7514), .A2(n7571), .ZN(n7604) );
  INV_X1 U8690 ( .A(n7604), .ZN(n7515) );
  AOI21_X1 U8691 ( .B1(n10903), .B2(n7516), .A(n7515), .ZN(n10904) );
  OAI22_X1 U8692 ( .A1(n10144), .A2(n7571), .B1(n7517), .B2(n10090), .ZN(n7518) );
  AOI21_X1 U8693 ( .B1(n10904), .B2(n10115), .A(n7518), .ZN(n7519) );
  OAI211_X1 U8694 ( .C1(n10907), .C2(n10055), .A(n7520), .B(n7519), .ZN(
        P1_U3285) );
  NAND2_X1 U8695 ( .A1(n8656), .A2(n10931), .ZN(n7521) );
  NAND2_X1 U8696 ( .A1(n7523), .A2(n8616), .ZN(n7526) );
  OR2_X1 U8697 ( .A1(n5039), .A2(n7524), .ZN(n7525) );
  OAI211_X1 U8698 ( .C1(n7537), .C2(n7527), .A(n7526), .B(n7525), .ZN(n7640)
         );
  NAND2_X1 U8699 ( .A1(n7711), .A2(n7640), .ZN(n8661) );
  NAND2_X1 U8700 ( .A1(n8992), .A2(n7704), .ZN(n8662) );
  NAND2_X1 U8701 ( .A1(n8661), .A2(n8662), .ZN(n8773) );
  INV_X1 U8702 ( .A(n7543), .ZN(n7633) );
  NOR2_X1 U8703 ( .A1(n7711), .A2(n7704), .ZN(n7541) );
  NAND2_X1 U8704 ( .A1(n8047), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7535) );
  OR2_X1 U8705 ( .A1(n8324), .A2(n7528), .ZN(n7534) );
  OAI21_X1 U8706 ( .B1(n7529), .B2(n7592), .A(n10450), .ZN(n7531) );
  NAND2_X1 U8707 ( .A1(n7531), .A2(n7530), .ZN(n7723) );
  OR2_X1 U8708 ( .A1(n8321), .A2(n7723), .ZN(n7533) );
  OR2_X1 U8709 ( .A1(n8253), .A2(n7005), .ZN(n7532) );
  NAND2_X1 U8710 ( .A1(n7536), .A2(n8616), .ZN(n7540) );
  AOI22_X1 U8711 ( .A1(n8235), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8234), .B2(
        n7538), .ZN(n7539) );
  NAND2_X1 U8712 ( .A1(n7540), .A2(n7539), .ZN(n10959) );
  NAND2_X1 U8713 ( .A1(n7761), .A2(n10959), .ZN(n8672) );
  INV_X1 U8714 ( .A(n7761), .ZN(n8991) );
  NAND2_X1 U8715 ( .A1(n7762), .A2(n8991), .ZN(n8667) );
  OAI21_X1 U8716 ( .B1(n7633), .B2(n7541), .A(n8772), .ZN(n7544) );
  NOR2_X1 U8717 ( .A1(n8772), .A2(n7541), .ZN(n7542) );
  NAND2_X1 U8718 ( .A1(n7543), .A2(n7542), .ZN(n7764) );
  AOI21_X1 U8719 ( .B1(n7544), .B2(n7764), .A(n10990), .ZN(n7546) );
  OR2_X1 U8720 ( .A1(n7711), .A2(n9272), .ZN(n7545) );
  OAI21_X1 U8721 ( .B1(n8929), .B2(n9270), .A(n7545), .ZN(n7719) );
  NOR2_X1 U8722 ( .A1(n7546), .A2(n7719), .ZN(n7551) );
  OAI211_X1 U8723 ( .C1(n7549), .C2(n8772), .A(n7747), .B(n10822), .ZN(n7550)
         );
  NAND2_X1 U8724 ( .A1(n7551), .A2(n7550), .ZN(n10957) );
  INV_X1 U8725 ( .A(n10957), .ZN(n7555) );
  OAI22_X1 U8726 ( .A1(n10829), .A2(n7005), .B1(n7723), .B2(n10823), .ZN(n7553) );
  NOR2_X1 U8727 ( .A1(n7629), .A2(n7762), .ZN(n10956) );
  NAND2_X1 U8728 ( .A1(n7629), .A2(n7762), .ZN(n7771) );
  INV_X1 U8729 ( .A(n7771), .ZN(n10955) );
  NOR3_X1 U8730 ( .A1(n10956), .A2(n10955), .A3(n10818), .ZN(n7552) );
  AOI211_X1 U8731 ( .C1(n9292), .C2(n10959), .A(n7553), .B(n7552), .ZN(n7554)
         );
  OAI21_X1 U8732 ( .B1(n7555), .B2(n9303), .A(n7554), .ZN(P2_U3287) );
  INV_X1 U8733 ( .A(n8245), .ZN(n7556) );
  OAI222_X1 U8734 ( .A1(n8494), .A2(n7556), .B1(n8801), .B2(P2_U3152), .C1(
        n8246), .C2(n5036), .ZN(P2_U3338) );
  OAI222_X1 U8735 ( .A1(P1_U3084), .A2(n9823), .B1(n10265), .B2(n7556), .C1(
        n10562), .C2(n10267), .ZN(P1_U3333) );
  INV_X1 U8736 ( .A(n9846), .ZN(n7557) );
  OR2_X1 U8737 ( .A1(n10945), .A2(n7557), .ZN(n9669) );
  NAND2_X1 U8738 ( .A1(n10945), .A2(n7557), .ZN(n9670) );
  NAND2_X1 U8739 ( .A1(n7559), .A2(n7558), .ZN(n7560) );
  NAND2_X1 U8740 ( .A1(n7608), .A2(n9847), .ZN(n7575) );
  AND2_X1 U8741 ( .A1(n7575), .A2(n7598), .ZN(n9611) );
  NAND2_X2 U8742 ( .A1(n7560), .A2(n9611), .ZN(n9802) );
  NAND2_X1 U8743 ( .A1(n7561), .A2(n10921), .ZN(n9661) );
  NAND2_X1 U8744 ( .A1(n7679), .A2(n7564), .ZN(n9659) );
  NAND2_X1 U8745 ( .A1(n9660), .A2(n9659), .ZN(n9658) );
  INV_X1 U8746 ( .A(n9658), .ZN(n7562) );
  OAI21_X1 U8747 ( .B1(n9772), .B2(n7563), .A(n7808), .ZN(n7566) );
  OAI22_X1 U8748 ( .A1(n7564), .A2(n10081), .B1(n7866), .B2(n10083), .ZN(n7565) );
  AOI21_X1 U8749 ( .B1(n7566), .B2(n10125), .A(n7565), .ZN(n10952) );
  AND2_X1 U8750 ( .A1(n7667), .A2(n10945), .ZN(n7567) );
  NOR2_X1 U8751 ( .A1(n7810), .A2(n7567), .ZN(n10947) );
  INV_X1 U8752 ( .A(n10945), .ZN(n7652) );
  INV_X1 U8753 ( .A(n7568), .ZN(n7655) );
  AOI22_X1 U8754 ( .A1(n10141), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7655), .B2(
        n10139), .ZN(n7569) );
  OAI21_X1 U8755 ( .B1(n7652), .B2(n10144), .A(n7569), .ZN(n7570) );
  AOI21_X1 U8756 ( .B1(n10947), .B2(n10115), .A(n7570), .ZN(n7579) );
  NAND2_X1 U8757 ( .A1(n7572), .A2(n7571), .ZN(n7573) );
  NAND2_X1 U8758 ( .A1(n7574), .A2(n7573), .ZN(n7597) );
  NAND2_X1 U8759 ( .A1(n7575), .A2(n9661), .ZN(n9769) );
  NOR2_X1 U8760 ( .A1(n10921), .A2(n9847), .ZN(n7576) );
  NAND2_X1 U8761 ( .A1(n7659), .A2(n9658), .ZN(n7661) );
  NAND2_X1 U8762 ( .A1(n7679), .A2(n7648), .ZN(n7577) );
  NAND2_X1 U8763 ( .A1(n7661), .A2(n7577), .ZN(n7816) );
  XNOR2_X1 U8764 ( .A(n7816), .B(n9772), .ZN(n10949) );
  NAND2_X1 U8765 ( .A1(n10949), .A2(n9929), .ZN(n7578) );
  OAI211_X1 U8766 ( .C1(n10952), .C2(n10141), .A(n7579), .B(n7578), .ZN(
        P1_U3282) );
  NOR3_X1 U8767 ( .A1(n8922), .A2(n7580), .A3(n8656), .ZN(n7591) );
  NOR2_X1 U8768 ( .A1(n7711), .A2(n8562), .ZN(n7581) );
  XNOR2_X1 U8769 ( .A(n7640), .B(n8551), .ZN(n7582) );
  NAND2_X1 U8770 ( .A1(n7581), .A2(n7582), .ZN(n7714) );
  INV_X1 U8771 ( .A(n7581), .ZN(n7583) );
  INV_X1 U8772 ( .A(n7582), .ZN(n7712) );
  NAND2_X1 U8773 ( .A1(n7583), .A2(n7712), .ZN(n7584) );
  NAND2_X1 U8774 ( .A1(n7714), .A2(n7584), .ZN(n7586) );
  AOI21_X1 U8775 ( .B1(n7588), .B2(n7586), .A(n8953), .ZN(n7590) );
  INV_X1 U8776 ( .A(n7585), .ZN(n7587) );
  INV_X1 U8777 ( .A(n7718), .ZN(n7589) );
  OAI21_X1 U8778 ( .B1(n7591), .B2(n7590), .A(n7589), .ZN(n7596) );
  OAI22_X1 U8779 ( .A1(n8964), .A2(n7761), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7592), .ZN(n7594) );
  NOR2_X1 U8780 ( .A1(n8968), .A2(n7638), .ZN(n7593) );
  AOI211_X1 U8781 ( .C1(n8966), .C2(n8993), .A(n7594), .B(n7593), .ZN(n7595)
         );
  OAI211_X1 U8782 ( .C1(n7704), .C2(n8963), .A(n7596), .B(n7595), .ZN(P2_U3223) );
  XOR2_X1 U8783 ( .A(n9769), .B(n7597), .Z(n10924) );
  INV_X1 U8784 ( .A(n7598), .ZN(n7599) );
  OR2_X1 U8785 ( .A1(n7509), .A2(n7599), .ZN(n7600) );
  NAND2_X1 U8786 ( .A1(n7600), .A2(n9609), .ZN(n7601) );
  XOR2_X1 U8787 ( .A(n9769), .B(n7601), .Z(n7602) );
  AOI222_X1 U8788 ( .A1(n10125), .A2(n7602), .B1(n9848), .B2(n10131), .C1(
        n7648), .C2(n10130), .ZN(n10925) );
  MUX2_X1 U8789 ( .A(n7603), .B(n10925), .S(n10093), .Z(n7611) );
  AOI211_X1 U8790 ( .C1(n10921), .C2(n7604), .A(n11009), .B(n5312), .ZN(n10920) );
  NOR2_X1 U8791 ( .A1(n7605), .A2(n10659), .ZN(n10138) );
  INV_X1 U8792 ( .A(n7606), .ZN(n7607) );
  OAI22_X1 U8793 ( .A1(n10144), .A2(n7608), .B1(n7607), .B2(n10090), .ZN(n7609) );
  AOI21_X1 U8794 ( .B1(n10920), .B2(n10138), .A(n7609), .ZN(n7610) );
  OAI211_X1 U8795 ( .C1(n10148), .C2(n10924), .A(n7611), .B(n7610), .ZN(
        P1_U3284) );
  INV_X1 U8796 ( .A(n9004), .ZN(n7614) );
  INV_X1 U8797 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10972) );
  MUX2_X1 U8798 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10972), .S(n9004), .Z(n9007) );
  OAI21_X1 U8799 ( .B1(n7613), .B2(n7157), .A(n7612), .ZN(n9008) );
  NAND2_X1 U8800 ( .A1(n9007), .A2(n9008), .ZN(n9006) );
  OAI21_X1 U8801 ( .B1(n7614), .B2(n10972), .A(n9006), .ZN(n7616) );
  INV_X1 U8802 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7791) );
  MUX2_X1 U8803 ( .A(n7791), .B(P2_REG1_REG_12__SCAN_IN), .S(n7785), .Z(n7615)
         );
  NOR2_X1 U8804 ( .A1(n7615), .A2(n7616), .ZN(n7689) );
  AOI21_X1 U8805 ( .B1(n7616), .B2(n7615), .A(n7689), .ZN(n7619) );
  INV_X1 U8806 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10302) );
  NOR2_X1 U8807 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10302), .ZN(n7617) );
  AOI21_X1 U8808 ( .B1(n10800), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7617), .ZN(
        n7618) );
  OAI21_X1 U8809 ( .B1(n7619), .B2(n10773), .A(n7618), .ZN(n7626) );
  NOR2_X1 U8810 ( .A1(n9004), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7621) );
  AOI21_X1 U8811 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n9004), .A(n7621), .ZN(
        n9002) );
  NAND2_X1 U8812 ( .A1(n9001), .A2(n9002), .ZN(n9000) );
  OAI21_X1 U8813 ( .B1(n9004), .B2(P2_REG2_REG_11__SCAN_IN), .A(n9000), .ZN(
        n7624) );
  NAND2_X1 U8814 ( .A1(n7785), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7622) );
  OAI21_X1 U8815 ( .B1(n7785), .B2(P2_REG2_REG_12__SCAN_IN), .A(n7622), .ZN(
        n7623) );
  NOR2_X1 U8816 ( .A1(n7623), .A2(n7624), .ZN(n7693) );
  AOI211_X1 U8817 ( .C1(n7624), .C2(n7623), .A(n7693), .B(n10801), .ZN(n7625)
         );
  AOI211_X1 U8818 ( .C1(n10807), .C2(n7785), .A(n7626), .B(n7625), .ZN(n7627)
         );
  INV_X1 U8819 ( .A(n7627), .ZN(P2_U3257) );
  OAI21_X1 U8820 ( .B1(n7628), .B2(n7704), .A(n10881), .ZN(n7630) );
  OR2_X1 U8821 ( .A1(n7630), .A2(n7629), .ZN(n7702) );
  OAI21_X1 U8822 ( .B1(n7632), .B2(n7548), .A(n7631), .ZN(n7637) );
  OAI22_X1 U8823 ( .A1(n8656), .A2(n9272), .B1(n7761), .B2(n9270), .ZN(n7636)
         );
  AOI211_X1 U8824 ( .C1(n7548), .C2(n7634), .A(n10990), .B(n7633), .ZN(n7635)
         );
  AOI211_X1 U8825 ( .C1(n10822), .C2(n7637), .A(n7636), .B(n7635), .ZN(n7703)
         );
  OR2_X1 U8826 ( .A1(n7703), .A2(n9303), .ZN(n7642) );
  OAI22_X1 U8827 ( .A1(n10829), .A2(n6944), .B1(n7638), .B2(n10823), .ZN(n7639) );
  AOI21_X1 U8828 ( .B1(n9292), .B2(n7640), .A(n7639), .ZN(n7641) );
  OAI211_X1 U8829 ( .C1(n7702), .C2(n9280), .A(n7642), .B(n7641), .ZN(P2_U3288) );
  INV_X1 U8830 ( .A(n7643), .ZN(n7647) );
  AOI21_X1 U8831 ( .B1(n7644), .B2(n7676), .A(n7645), .ZN(n7646) );
  OAI21_X1 U8832 ( .B1(n7647), .B2(n7646), .A(n9525), .ZN(n7657) );
  NAND2_X1 U8833 ( .A1(n9561), .A2(n7648), .ZN(n7651) );
  INV_X1 U8834 ( .A(n7649), .ZN(n7650) );
  OAI211_X1 U8835 ( .C1(n7866), .C2(n9559), .A(n7651), .B(n7650), .ZN(n7654)
         );
  NOR2_X1 U8836 ( .A1(n7652), .A2(n9535), .ZN(n7653) );
  AOI211_X1 U8837 ( .C1(n7655), .C2(n9505), .A(n7654), .B(n7653), .ZN(n7656)
         );
  NAND2_X1 U8838 ( .A1(n7657), .A2(n7656), .ZN(P1_U3229) );
  INV_X1 U8839 ( .A(n8203), .ZN(n7688) );
  OAI222_X1 U8840 ( .A1(n8494), .A2(n7688), .B1(n5036), .B2(n7658), .C1(n8807), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  OR2_X1 U8841 ( .A1(n7659), .A2(n9658), .ZN(n7660) );
  NAND2_X1 U8842 ( .A1(n7661), .A2(n7660), .ZN(n10938) );
  XNOR2_X1 U8843 ( .A(n7662), .B(n7562), .ZN(n7663) );
  NAND2_X1 U8844 ( .A1(n7663), .A2(n10125), .ZN(n7665) );
  AOI22_X1 U8845 ( .A1(n10130), .A2(n9846), .B1(n9847), .B2(n10131), .ZN(n7664) );
  OAI211_X1 U8846 ( .C1(n7255), .C2(n10938), .A(n7665), .B(n7664), .ZN(n10941)
         );
  MUX2_X1 U8847 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10941), .S(n10093), .Z(n7666) );
  INV_X1 U8848 ( .A(n7666), .ZN(n7672) );
  INV_X1 U8849 ( .A(n7667), .ZN(n7668) );
  AOI21_X1 U8850 ( .B1(n7679), .B2(n7669), .A(n7668), .ZN(n10939) );
  OAI22_X1 U8851 ( .A1(n10144), .A2(n5311), .B1(n10090), .B2(n7680), .ZN(n7670) );
  AOI21_X1 U8852 ( .B1(n10939), .B2(n10115), .A(n7670), .ZN(n7671) );
  OAI211_X1 U8853 ( .C1(n10938), .C2(n10055), .A(n7672), .B(n7671), .ZN(
        P1_U3283) );
  INV_X1 U8854 ( .A(n7644), .ZN(n7677) );
  AOI21_X1 U8855 ( .B1(n7676), .B2(n7674), .A(n7673), .ZN(n7675) );
  AOI211_X1 U8856 ( .C1(n7677), .C2(n7676), .A(n9569), .B(n7675), .ZN(n7687)
         );
  AOI21_X1 U8857 ( .B1(n9561), .B2(n9847), .A(n7678), .ZN(n7685) );
  NAND2_X1 U8858 ( .A1(n9566), .A2(n7679), .ZN(n7684) );
  INV_X1 U8859 ( .A(n7680), .ZN(n7681) );
  NAND2_X1 U8860 ( .A1(n9505), .A2(n7681), .ZN(n7683) );
  NAND2_X1 U8861 ( .A1(n9532), .A2(n9846), .ZN(n7682) );
  NAND4_X1 U8862 ( .A1(n7685), .A2(n7684), .A3(n7683), .A4(n7682), .ZN(n7686)
         );
  OR2_X1 U8863 ( .A1(n7687), .A2(n7686), .ZN(P1_U3219) );
  INV_X1 U8864 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10557) );
  OAI222_X1 U8865 ( .A1(P1_U3084), .A2(n5762), .B1(n10265), .B2(n7688), .C1(
        n10557), .C2(n10267), .ZN(P1_U3332) );
  AOI21_X1 U8866 ( .B1(n7690), .B2(n7791), .A(n7689), .ZN(n7692) );
  INV_X1 U8867 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11001) );
  AOI22_X1 U8868 ( .A1(n7992), .A2(n11001), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7824), .ZN(n7691) );
  NOR2_X1 U8869 ( .A1(n7692), .A2(n7691), .ZN(n7823) );
  AOI21_X1 U8870 ( .B1(n7692), .B2(n7691), .A(n7823), .ZN(n7701) );
  NOR2_X1 U8871 ( .A1(n7992), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7694) );
  AOI21_X1 U8872 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n7992), .A(n7694), .ZN(
        n7695) );
  NAND2_X1 U8873 ( .A1(n7696), .A2(n7695), .ZN(n7828) );
  OAI21_X1 U8874 ( .B1(n7696), .B2(n7695), .A(n7828), .ZN(n7697) );
  NAND2_X1 U8875 ( .A1(n7697), .A2(n10776), .ZN(n7700) );
  INV_X1 U8876 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7925) );
  NAND2_X1 U8877 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3152), .ZN(n8075) );
  OAI21_X1 U8878 ( .B1(n10787), .B2(n7925), .A(n8075), .ZN(n7698) );
  AOI21_X1 U8879 ( .B1(n10807), .B2(n7992), .A(n7698), .ZN(n7699) );
  OAI211_X1 U8880 ( .C1(n7701), .C2(n10773), .A(n7700), .B(n7699), .ZN(
        P2_U3258) );
  INV_X1 U8881 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7706) );
  OAI211_X1 U8882 ( .C1(n7704), .C2(n10992), .A(n7703), .B(n7702), .ZN(n7707)
         );
  NAND2_X1 U8883 ( .A1(n7707), .A2(n11006), .ZN(n7705) );
  OAI21_X1 U8884 ( .B1(n11006), .B2(n7706), .A(n7705), .ZN(P2_U3475) );
  NAND2_X1 U8885 ( .A1(n7707), .A2(n11002), .ZN(n7708) );
  OAI21_X1 U8886 ( .B1(n11002), .B2(n7453), .A(n7708), .ZN(P2_U3528) );
  INV_X1 U8887 ( .A(n8260), .ZN(n7710) );
  OAI222_X1 U8888 ( .A1(n5765), .A2(P1_U3084), .B1(n10265), .B2(n7710), .C1(
        n7709), .C2(n10267), .ZN(P1_U3331) );
  OAI222_X1 U8889 ( .A1(n5036), .A2(n8261), .B1(n8494), .B2(n7710), .C1(n8620), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  NOR3_X1 U8890 ( .A1(n7712), .A2(n8922), .A3(n7711), .ZN(n7713) );
  AOI21_X1 U8891 ( .B1(n7718), .B2(n8915), .A(n7713), .ZN(n7728) );
  XNOR2_X1 U8892 ( .A(n10959), .B(n8563), .ZN(n7837) );
  OR2_X1 U8893 ( .A1(n7761), .A2(n8562), .ZN(n7836) );
  XNOR2_X1 U8894 ( .A(n7837), .B(n7836), .ZN(n7716) );
  INV_X1 U8895 ( .A(n7716), .ZN(n7727) );
  INV_X1 U8896 ( .A(n7714), .ZN(n7715) );
  NOR2_X1 U8897 ( .A1(n8963), .A2(n7762), .ZN(n7725) );
  NAND2_X1 U8898 ( .A1(n7719), .A2(n8882), .ZN(n7722) );
  INV_X1 U8899 ( .A(n7720), .ZN(n7721) );
  OAI211_X1 U8900 ( .C1(n8968), .C2(n7723), .A(n7722), .B(n7721), .ZN(n7724)
         );
  AOI211_X1 U8901 ( .C1(n7839), .C2(n8915), .A(n7725), .B(n7724), .ZN(n7726)
         );
  OAI21_X1 U8902 ( .B1(n7728), .B2(n7727), .A(n7726), .ZN(P2_U3233) );
  INV_X1 U8903 ( .A(n7729), .ZN(n7732) );
  INV_X1 U8904 ( .A(n7730), .ZN(n7738) );
  AOI21_X1 U8905 ( .B1(n7732), .B2(n7738), .A(n7731), .ZN(n7735) );
  NAND2_X1 U8906 ( .A1(n9860), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7733) );
  OAI21_X1 U8907 ( .B1(n9860), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7733), .ZN(
        n7734) );
  NOR2_X1 U8908 ( .A1(n7735), .A2(n7734), .ZN(n9859) );
  AOI211_X1 U8909 ( .C1(n7735), .C2(n7734), .A(n9859), .B(n9869), .ZN(n7746)
         );
  INV_X1 U8910 ( .A(n7736), .ZN(n7739) );
  AOI21_X1 U8911 ( .B1(n7739), .B2(n7738), .A(n7737), .ZN(n7741) );
  XNOR2_X1 U8912 ( .A(n9860), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7740) );
  NOR2_X1 U8913 ( .A1(n7741), .A2(n7740), .ZN(n9854) );
  AOI211_X1 U8914 ( .C1(n7741), .C2(n7740), .A(n9854), .B(n10754), .ZN(n7745)
         );
  NAND2_X1 U8915 ( .A1(n10761), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7742) );
  NAND2_X1 U8916 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9488) );
  OAI211_X1 U8917 ( .C1(n7743), .C2(n9899), .A(n7742), .B(n9488), .ZN(n7744)
         );
  OR3_X1 U8918 ( .A1(n7746), .A2(n7745), .A3(n7744), .ZN(P1_U3257) );
  NAND2_X1 U8919 ( .A1(n7748), .A2(n8616), .ZN(n7751) );
  AOI22_X1 U8920 ( .A1(n8235), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8234), .B2(
        n7749), .ZN(n7750) );
  OR2_X1 U8921 ( .A1(n7856), .A2(n8929), .ZN(n8668) );
  NAND2_X1 U8922 ( .A1(n7856), .A2(n8929), .ZN(n8669) );
  INV_X1 U8923 ( .A(n8777), .ZN(n7765) );
  XNOR2_X1 U8924 ( .A(n7780), .B(n7765), .ZN(n7768) );
  NAND2_X1 U8925 ( .A1(n8047), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7759) );
  INV_X1 U8926 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7752) );
  OR2_X1 U8927 ( .A1(n8253), .A2(n7752), .ZN(n7758) );
  INV_X1 U8928 ( .A(n7753), .ZN(n7788) );
  NAND2_X1 U8929 ( .A1(n7754), .A2(n10448), .ZN(n7755) );
  NAND2_X1 U8930 ( .A1(n7788), .A2(n7755), .ZN(n8933) );
  OR2_X1 U8931 ( .A1(n8321), .A2(n8933), .ZN(n7757) );
  OR2_X1 U8932 ( .A1(n8324), .A2(n10972), .ZN(n7756) );
  OR2_X1 U8933 ( .A1(n7761), .A2(n9272), .ZN(n7760) );
  OAI21_X1 U8934 ( .B1(n8033), .B2(n9270), .A(n7760), .ZN(n7844) );
  NAND2_X1 U8935 ( .A1(n7762), .A2(n7761), .ZN(n7763) );
  INV_X1 U8936 ( .A(n7887), .ZN(n7766) );
  AOI211_X1 U8937 ( .C1(n8777), .C2(n5124), .A(n10990), .B(n7766), .ZN(n7767)
         );
  AOI211_X1 U8938 ( .C1(n10822), .C2(n7768), .A(n7844), .B(n7767), .ZN(n7859)
         );
  OAI22_X1 U8939 ( .A1(n10829), .A2(n7769), .B1(n7843), .B2(n10823), .ZN(n7770) );
  AOI21_X1 U8940 ( .B1(n9292), .B2(n7856), .A(n7770), .ZN(n7773) );
  AOI21_X1 U8941 ( .B1(n7856), .B2(n7771), .A(n5324), .ZN(n7857) );
  NAND2_X1 U8942 ( .A1(n7857), .A2(n9226), .ZN(n7772) );
  OAI211_X1 U8943 ( .C1(n7859), .C2(n9303), .A(n7773), .B(n7772), .ZN(P2_U3286) );
  NAND2_X1 U8944 ( .A1(n8047), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7779) );
  INV_X1 U8945 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8001) );
  OR2_X1 U8946 ( .A1(n8253), .A2(n8001), .ZN(n7778) );
  NAND2_X1 U8947 ( .A1(n7790), .A2(n7774), .ZN(n7775) );
  NAND2_X1 U8948 ( .A1(n7985), .A2(n7775), .ZN(n8076) );
  OR2_X1 U8949 ( .A1(n8321), .A2(n8076), .ZN(n7777) );
  OR2_X1 U8950 ( .A1(n8324), .A2(n11001), .ZN(n7776) );
  AOI22_X1 U8951 ( .A1(n8235), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8234), .B2(
        n9004), .ZN(n7782) );
  OR2_X1 U8952 ( .A1(n10970), .A2(n8033), .ZN(n7996) );
  AND2_X1 U8953 ( .A1(n7996), .A2(n8668), .ZN(n8674) );
  NAND2_X1 U8954 ( .A1(n10970), .A2(n8033), .ZN(n8670) );
  INV_X1 U8955 ( .A(n8670), .ZN(n7783) );
  AOI21_X1 U8956 ( .B1(n7881), .B2(n8674), .A(n7783), .ZN(n7796) );
  NAND2_X1 U8957 ( .A1(n7784), .A2(n8616), .ZN(n7787) );
  AOI22_X1 U8958 ( .A1(n8235), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8234), .B2(
        n7785), .ZN(n7786) );
  NAND2_X1 U8959 ( .A1(n8047), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7795) );
  INV_X1 U8960 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7802) );
  OR2_X1 U8961 ( .A1(n8253), .A2(n7802), .ZN(n7794) );
  NAND2_X1 U8962 ( .A1(n7788), .A2(n10302), .ZN(n7789) );
  NAND2_X1 U8963 ( .A1(n7790), .A2(n7789), .ZN(n8038) );
  OR2_X1 U8964 ( .A1(n8321), .A2(n8038), .ZN(n7793) );
  OR2_X1 U8965 ( .A1(n8324), .A2(n7791), .ZN(n7792) );
  OR2_X1 U8966 ( .A1(n8028), .A2(n8928), .ZN(n8679) );
  NAND2_X1 U8967 ( .A1(n8028), .A2(n8928), .ZN(n7997) );
  NAND2_X1 U8968 ( .A1(n8679), .A2(n7997), .ZN(n8684) );
  INV_X1 U8969 ( .A(n8684), .ZN(n7800) );
  XNOR2_X1 U8970 ( .A(n7796), .B(n7800), .ZN(n7797) );
  OAI222_X1 U8971 ( .A1(n9270), .A2(n8596), .B1(n9272), .B2(n8033), .C1(n7797), 
        .C2(n9264), .ZN(n10977) );
  INV_X1 U8972 ( .A(n10977), .ZN(n7807) );
  NAND2_X1 U8973 ( .A1(n7856), .A2(n7882), .ZN(n7885) );
  NAND2_X1 U8974 ( .A1(n7996), .A2(n8670), .ZN(n7884) );
  INV_X1 U8975 ( .A(n8033), .ZN(n8990) );
  NAND2_X1 U8976 ( .A1(n10970), .A2(n8990), .ZN(n7799) );
  AND2_X2 U8977 ( .A1(n7883), .A2(n7799), .ZN(n7801) );
  OAI21_X1 U8978 ( .B1(n7801), .B2(n8684), .A(n8007), .ZN(n10979) );
  XNOR2_X1 U8979 ( .A(n8002), .B(n8028), .ZN(n10976) );
  OAI22_X1 U8980 ( .A1(n10829), .A2(n7802), .B1(n8038), .B2(n10823), .ZN(n7803) );
  AOI21_X1 U8981 ( .B1(n9292), .B2(n8028), .A(n7803), .ZN(n7804) );
  OAI21_X1 U8982 ( .B1(n10976), .B2(n10818), .A(n7804), .ZN(n7805) );
  AOI21_X1 U8983 ( .B1(n10979), .B2(n10827), .A(n7805), .ZN(n7806) );
  OAI21_X1 U8984 ( .B1(n7807), .B2(n9303), .A(n7806), .ZN(P2_U3284) );
  NAND2_X1 U8985 ( .A1(n7808), .A2(n9670), .ZN(n7865) );
  OR2_X1 U8986 ( .A1(n7978), .A2(n7866), .ZN(n9673) );
  NAND2_X1 U8987 ( .A1(n7978), .A2(n7866), .ZN(n9674) );
  XNOR2_X1 U8988 ( .A(n7865), .B(n9773), .ZN(n7809) );
  AOI222_X1 U8989 ( .A1(n10125), .A2(n7809), .B1(n9844), .B2(n10130), .C1(
        n9846), .C2(n10131), .ZN(n7980) );
  INV_X1 U8990 ( .A(n7810), .ZN(n7811) );
  INV_X1 U8991 ( .A(n7978), .ZN(n7814) );
  INV_X1 U8992 ( .A(n7870), .ZN(n7871) );
  AOI211_X1 U8993 ( .C1(n7978), .C2(n7811), .A(n11009), .B(n7871), .ZN(n7977)
         );
  INV_X1 U8994 ( .A(n7950), .ZN(n7812) );
  AOI22_X1 U8995 ( .A1(n10141), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7812), .B2(
        n10139), .ZN(n7813) );
  OAI21_X1 U8996 ( .B1(n7814), .B2(n10144), .A(n7813), .ZN(n7821) );
  OR2_X1 U8997 ( .A1(n10945), .A2(n9846), .ZN(n7815) );
  NAND2_X1 U8998 ( .A1(n10945), .A2(n9846), .ZN(n7817) );
  INV_X1 U8999 ( .A(n7863), .ZN(n7818) );
  AOI21_X1 U9000 ( .B1(n9773), .B2(n7819), .A(n7818), .ZN(n7981) );
  NOR2_X1 U9001 ( .A1(n7981), .A2(n10148), .ZN(n7820) );
  AOI211_X1 U9002 ( .C1(n7977), .C2(n10138), .A(n7821), .B(n7820), .ZN(n7822)
         );
  OAI21_X1 U9003 ( .B1(n10141), .B2(n7980), .A(n7822), .ZN(P1_U3281) );
  AOI21_X1 U9004 ( .B1(n7824), .B2(n11001), .A(n7823), .ZN(n7826) );
  INV_X1 U9005 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9020) );
  AOI22_X1 U9006 ( .A1(n9014), .A2(n9020), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n9021), .ZN(n7825) );
  NOR2_X1 U9007 ( .A1(n7826), .A2(n7825), .ZN(n9019) );
  AOI21_X1 U9008 ( .B1(n7826), .B2(n7825), .A(n9019), .ZN(n7835) );
  NOR2_X1 U9009 ( .A1(n9014), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7827) );
  AOI21_X1 U9010 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n9014), .A(n7827), .ZN(
        n7830) );
  OAI21_X1 U9011 ( .B1(n7992), .B2(P2_REG2_REG_13__SCAN_IN), .A(n7828), .ZN(
        n7829) );
  NAND2_X1 U9012 ( .A1(n7830), .A2(n7829), .ZN(n9013) );
  OAI21_X1 U9013 ( .B1(n7830), .B2(n7829), .A(n9013), .ZN(n7831) );
  NAND2_X1 U9014 ( .A1(n7831), .A2(n10776), .ZN(n7834) );
  INV_X1 U9015 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7928) );
  NAND2_X1 U9016 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n8595) );
  OAI21_X1 U9017 ( .B1(n10787), .B2(n7928), .A(n8595), .ZN(n7832) );
  AOI21_X1 U9018 ( .B1(n10807), .B2(n9014), .A(n7832), .ZN(n7833) );
  OAI211_X1 U9019 ( .C1(n7835), .C2(n10773), .A(n7834), .B(n7833), .ZN(
        P2_U3259) );
  INV_X1 U9020 ( .A(n7856), .ZN(n7851) );
  AND2_X1 U9021 ( .A1(n7837), .A2(n7836), .ZN(n7838) );
  XNOR2_X1 U9022 ( .A(n7856), .B(n8563), .ZN(n8923) );
  OR2_X1 U9023 ( .A1(n8929), .A2(n8562), .ZN(n7840) );
  NOR2_X1 U9024 ( .A1(n8923), .A2(n7840), .ZN(n8023) );
  AOI21_X1 U9025 ( .B1(n8923), .B2(n7840), .A(n8023), .ZN(n7841) );
  OAI211_X1 U9026 ( .C1(n7842), .C2(n7841), .A(n8925), .B(n8915), .ZN(n7850)
         );
  INV_X1 U9027 ( .A(n7843), .ZN(n7848) );
  INV_X1 U9028 ( .A(n7844), .ZN(n7846) );
  OAI22_X1 U9029 ( .A1(n7846), .A2(n7845), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10527), .ZN(n7847) );
  AOI21_X1 U9030 ( .B1(n7848), .B2(n8935), .A(n7847), .ZN(n7849) );
  OAI211_X1 U9031 ( .C1(n7851), .C2(n8963), .A(n7850), .B(n7849), .ZN(P2_U3219) );
  INV_X1 U9032 ( .A(n8270), .ZN(n7854) );
  NOR2_X1 U9033 ( .A1(n7852), .A2(P1_U3084), .ZN(n9832) );
  AOI21_X1 U9034 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n10658), .A(n9832), .ZN(
        n7853) );
  OAI21_X1 U9035 ( .B1(n7854), .B2(n10265), .A(n7853), .ZN(P1_U3330) );
  NAND2_X1 U9036 ( .A1(n8270), .A2(n9420), .ZN(n7855) );
  OAI211_X1 U9037 ( .C1(n8271), .C2(n5036), .A(n7855), .B(n8823), .ZN(P2_U3335) );
  INV_X1 U9038 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7861) );
  AOI22_X1 U9039 ( .A1(n7857), .A2(n10881), .B1(n10971), .B2(n7856), .ZN(n7858) );
  NAND2_X1 U9040 ( .A1(n7859), .A2(n7858), .ZN(n7877) );
  NAND2_X1 U9041 ( .A1(n7877), .A2(n11006), .ZN(n7860) );
  OAI21_X1 U9042 ( .B1(n11006), .B2(n7861), .A(n7860), .ZN(P2_U3481) );
  OR2_X1 U9043 ( .A1(n7978), .A2(n9845), .ZN(n7862) );
  NAND2_X1 U9044 ( .A1(n8020), .A2(n7957), .ZN(n9679) );
  NAND2_X1 U9045 ( .A1(n9678), .A2(n9679), .ZN(n9775) );
  OAI21_X1 U9046 ( .B1(n7864), .B2(n9775), .A(n7961), .ZN(n10966) );
  INV_X1 U9047 ( .A(n10966), .ZN(n7876) );
  XNOR2_X1 U9048 ( .A(n7955), .B(n9775), .ZN(n7869) );
  OAI22_X1 U9049 ( .A1(n7866), .A2(n10081), .B1(n8117), .B2(n10083), .ZN(n7867) );
  AOI21_X1 U9050 ( .B1(n10966), .B2(n10929), .A(n7867), .ZN(n7868) );
  OAI21_X1 U9051 ( .B1(n7869), .B2(n9972), .A(n7868), .ZN(n10964) );
  NAND2_X1 U9052 ( .A1(n10964), .A2(n10093), .ZN(n7875) );
  OAI22_X1 U9053 ( .A1(n10093), .A2(n5746), .B1(n8018), .B2(n10090), .ZN(n7873) );
  INV_X1 U9054 ( .A(n8020), .ZN(n10963) );
  OAI211_X1 U9055 ( .C1(n7871), .C2(n10963), .A(n11021), .B(n7965), .ZN(n10962) );
  INV_X1 U9056 ( .A(n10138), .ZN(n7971) );
  NOR2_X1 U9057 ( .A1(n10962), .A2(n7971), .ZN(n7872) );
  AOI211_X1 U9058 ( .C1(n10095), .C2(n8020), .A(n7873), .B(n7872), .ZN(n7874)
         );
  OAI211_X1 U9059 ( .C1(n7876), .C2(n10055), .A(n7875), .B(n7874), .ZN(
        P1_U3280) );
  NAND2_X1 U9060 ( .A1(n7877), .A2(n11002), .ZN(n7878) );
  OAI21_X1 U9061 ( .B1(n11002), .B2(n7157), .A(n7878), .ZN(P2_U3530) );
  INV_X1 U9062 ( .A(n8002), .ZN(n7879) );
  AOI211_X1 U9063 ( .C1(n10970), .C2(n7880), .A(n10994), .B(n7879), .ZN(n10969) );
  NOR2_X1 U9064 ( .A1(n10823), .A2(n8933), .ZN(n7892) );
  NAND2_X1 U9065 ( .A1(n7881), .A2(n8668), .ZN(n7995) );
  XOR2_X1 U9066 ( .A(n7995), .B(n7884), .Z(n7891) );
  INV_X1 U9067 ( .A(n8928), .ZN(n8989) );
  AOI22_X1 U9068 ( .A1(n9254), .A2(n7882), .B1(n8989), .B2(n10821), .ZN(n7890)
         );
  INV_X1 U9069 ( .A(n7884), .ZN(n7886) );
  NAND3_X1 U9070 ( .A1(n7887), .A2(n7886), .A3(n7885), .ZN(n7888) );
  NAND3_X1 U9071 ( .A1(n7883), .A2(n10980), .A3(n7888), .ZN(n7889) );
  OAI211_X1 U9072 ( .C1(n7891), .C2(n9264), .A(n7890), .B(n7889), .ZN(n10968)
         );
  AOI211_X1 U9073 ( .C1(n10969), .C2(n8811), .A(n7892), .B(n10968), .ZN(n7894)
         );
  AOI22_X1 U9074 ( .A1(n9292), .A2(n10970), .B1(P2_REG2_REG_11__SCAN_IN), .B2(
        n9303), .ZN(n7893) );
  OAI21_X1 U9075 ( .B1(n7894), .B2(n9303), .A(n7893), .ZN(P2_U3285) );
  NOR2_X1 U9076 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7936) );
  NOR2_X1 U9077 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7934) );
  NOR2_X1 U9078 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7932) );
  NOR2_X1 U9079 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7930) );
  NOR2_X1 U9080 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7927) );
  NOR2_X1 U9081 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7924) );
  NAND2_X1 U9082 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7922) );
  XOR2_X1 U9083 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10725) );
  NAND2_X1 U9084 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7920) );
  XNOR2_X1 U9085 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n7895), .ZN(n10723) );
  NOR2_X1 U9086 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7903) );
  XOR2_X1 U9087 ( .A(n7896), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10714) );
  NAND2_X1 U9088 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7901) );
  XOR2_X1 U9089 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10712) );
  NAND2_X1 U9090 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7899) );
  XNOR2_X1 U9091 ( .A(n7897), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(n10710) );
  AOI21_X1 U9092 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10705) );
  INV_X1 U9093 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10786) );
  NAND3_X1 U9094 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10707) );
  OAI21_X1 U9095 ( .B1(n10705), .B2(n10786), .A(n10707), .ZN(n10709) );
  NAND2_X1 U9096 ( .A1(n10710), .A2(n10709), .ZN(n7898) );
  NAND2_X1 U9097 ( .A1(n7899), .A2(n7898), .ZN(n10711) );
  NAND2_X1 U9098 ( .A1(n10712), .A2(n10711), .ZN(n7900) );
  NAND2_X1 U9099 ( .A1(n7901), .A2(n7900), .ZN(n10713) );
  NOR2_X1 U9100 ( .A1(n10714), .A2(n10713), .ZN(n7902) );
  NOR2_X1 U9101 ( .A1(n7903), .A2(n7902), .ZN(n7904) );
  NOR2_X1 U9102 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7904), .ZN(n10716) );
  AND2_X1 U9103 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7904), .ZN(n10715) );
  NOR2_X1 U9104 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10715), .ZN(n7905) );
  NAND2_X1 U9105 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n7906), .ZN(n7908) );
  XOR2_X1 U9106 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n7906), .Z(n10718) );
  NAND2_X1 U9107 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10718), .ZN(n7907) );
  NAND2_X1 U9108 ( .A1(n7908), .A2(n7907), .ZN(n7909) );
  NAND2_X1 U9109 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7909), .ZN(n7911) );
  XOR2_X1 U9110 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7909), .Z(n10719) );
  NAND2_X1 U9111 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10719), .ZN(n7910) );
  NAND2_X1 U9112 ( .A1(n7911), .A2(n7910), .ZN(n7912) );
  NAND2_X1 U9113 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7912), .ZN(n7914) );
  XOR2_X1 U9114 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7912), .Z(n10720) );
  NAND2_X1 U9115 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10720), .ZN(n7913) );
  NAND2_X1 U9116 ( .A1(n7914), .A2(n7913), .ZN(n7915) );
  NAND2_X1 U9117 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n7915), .ZN(n7918) );
  XNOR2_X1 U9118 ( .A(n7916), .B(n7915), .ZN(n10721) );
  NAND2_X1 U9119 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10721), .ZN(n7917) );
  NAND2_X1 U9120 ( .A1(n7918), .A2(n7917), .ZN(n10722) );
  NAND2_X1 U9121 ( .A1(n10723), .A2(n10722), .ZN(n7919) );
  NAND2_X1 U9122 ( .A1(n7920), .A2(n7919), .ZN(n10724) );
  NAND2_X1 U9123 ( .A1(n10725), .A2(n10724), .ZN(n7921) );
  NAND2_X1 U9124 ( .A1(n7922), .A2(n7921), .ZN(n10727) );
  XNOR2_X1 U9125 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10726) );
  XOR2_X1 U9126 ( .A(n7925), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n10728) );
  NOR2_X1 U9127 ( .A1(n10729), .A2(n10728), .ZN(n7926) );
  NOR2_X1 U9128 ( .A1(n7927), .A2(n7926), .ZN(n10731) );
  XOR2_X1 U9129 ( .A(n7928), .B(P1_ADDR_REG_14__SCAN_IN), .Z(n10730) );
  NOR2_X1 U9130 ( .A1(n10731), .A2(n10730), .ZN(n7929) );
  NOR2_X1 U9131 ( .A1(n7930), .A2(n7929), .ZN(n10733) );
  XNOR2_X1 U9132 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10732) );
  NOR2_X1 U9133 ( .A1(n10733), .A2(n10732), .ZN(n7931) );
  NOR2_X1 U9134 ( .A1(n7932), .A2(n7931), .ZN(n10735) );
  XNOR2_X1 U9135 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10734) );
  NOR2_X1 U9136 ( .A1(n10735), .A2(n10734), .ZN(n7933) );
  NOR2_X1 U9137 ( .A1(n7934), .A2(n7933), .ZN(n10737) );
  XNOR2_X1 U9138 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10736) );
  NOR2_X1 U9139 ( .A1(n10737), .A2(n10736), .ZN(n7935) );
  NOR2_X1 U9140 ( .A1(n7936), .A2(n7935), .ZN(n7937) );
  AND2_X1 U9141 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n7937), .ZN(n10738) );
  NOR2_X1 U9142 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10738), .ZN(n7938) );
  NOR2_X1 U9143 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n7937), .ZN(n10739) );
  NOR2_X1 U9144 ( .A1(n7938), .A2(n10739), .ZN(n7940) );
  XNOR2_X1 U9145 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7939) );
  XNOR2_X1 U9146 ( .A(n7940), .B(n7939), .ZN(ADD_1071_U4) );
  INV_X1 U9147 ( .A(n7941), .ZN(n7945) );
  OR2_X1 U9148 ( .A1(n7942), .A2(n7941), .ZN(n7943) );
  AOI22_X1 U9149 ( .A1(n7946), .A2(n7945), .B1(n7944), .B2(n7943), .ZN(n7953)
         );
  NOR2_X1 U9150 ( .A1(n9559), .A2(n7957), .ZN(n7947) );
  AOI211_X1 U9151 ( .C1(n9561), .C2(n9846), .A(n7948), .B(n7947), .ZN(n7949)
         );
  OAI21_X1 U9152 ( .B1(n9564), .B2(n7950), .A(n7949), .ZN(n7951) );
  AOI21_X1 U9153 ( .B1(n7978), .B2(n9566), .A(n7951), .ZN(n7952) );
  OAI21_X1 U9154 ( .B1(n7953), .B2(n9569), .A(n7952), .ZN(P1_U3215) );
  INV_X1 U9155 ( .A(n9679), .ZN(n7954) );
  NAND2_X1 U9156 ( .A1(n8084), .A2(n9678), .ZN(n7956) );
  OR2_X1 U9157 ( .A1(n10233), .A2(n8117), .ZN(n9684) );
  NAND2_X1 U9158 ( .A1(n10233), .A2(n8117), .ZN(n9686) );
  XNOR2_X1 U9159 ( .A(n7956), .B(n7962), .ZN(n7959) );
  OAI22_X1 U9160 ( .A1(n7957), .A2(n10081), .B1(n8106), .B2(n10083), .ZN(n7958) );
  AOI21_X1 U9161 ( .B1(n7959), .B2(n10125), .A(n7958), .ZN(n10239) );
  OR2_X1 U9162 ( .A1(n8020), .A2(n9844), .ZN(n7960) );
  INV_X1 U9163 ( .A(n9777), .ZN(n7962) );
  NAND2_X1 U9164 ( .A1(n7963), .A2(n9777), .ZN(n7964) );
  AND2_X1 U9165 ( .A1(n8095), .A2(n7964), .ZN(n10237) );
  NOR2_X1 U9166 ( .A1(n7965), .A2(n10233), .ZN(n8122) );
  NAND2_X1 U9167 ( .A1(n7965), .A2(n10233), .ZN(n7966) );
  NAND2_X1 U9168 ( .A1(n7966), .A2(n11021), .ZN(n7967) );
  OR2_X1 U9169 ( .A1(n8122), .A2(n7967), .ZN(n10235) );
  OAI22_X1 U9170 ( .A1(n10093), .A2(n7968), .B1(n8110), .B2(n10090), .ZN(n7969) );
  AOI21_X1 U9171 ( .B1(n10233), .B2(n10095), .A(n7969), .ZN(n7970) );
  OAI21_X1 U9172 ( .B1(n10235), .B2(n7971), .A(n7970), .ZN(n7972) );
  AOI21_X1 U9173 ( .B1(n10237), .B2(n9929), .A(n7972), .ZN(n7973) );
  OAI21_X1 U9174 ( .B1(n10239), .B2(n10141), .A(n7973), .ZN(P1_U3279) );
  INV_X1 U9175 ( .A(n8275), .ZN(n7975) );
  OAI222_X1 U9176 ( .A1(n8494), .A2(n7975), .B1(n5036), .B2(n8276), .C1(
        P2_U3152), .C2(n7974), .ZN(P2_U3334) );
  OAI222_X1 U9177 ( .A1(n7976), .A2(P1_U3084), .B1(n10265), .B2(n7975), .C1(
        n10555), .C2(n10267), .ZN(P1_U3329) );
  AOI21_X1 U9178 ( .B1(n10946), .B2(n7978), .A(n7977), .ZN(n7979) );
  OAI211_X1 U9179 ( .C1(n10232), .C2(n7981), .A(n7980), .B(n7979), .ZN(n7983)
         );
  NAND2_X1 U9180 ( .A1(n7983), .A2(n11028), .ZN(n7982) );
  OAI21_X1 U9181 ( .B1(n11028), .B2(n5999), .A(n7982), .ZN(P1_U3484) );
  NAND2_X1 U9182 ( .A1(n7983), .A2(n11024), .ZN(n7984) );
  OAI21_X1 U9183 ( .B1(n11024), .B2(n6637), .A(n7984), .ZN(P1_U3533) );
  NAND2_X1 U9184 ( .A1(n8047), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7990) );
  INV_X1 U9185 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8060) );
  OR2_X1 U9186 ( .A1(n8253), .A2(n8060), .ZN(n7989) );
  NAND2_X1 U9187 ( .A1(n7985), .A2(n10521), .ZN(n7986) );
  NAND2_X1 U9188 ( .A1(n8049), .A2(n7986), .ZN(n8599) );
  OR2_X1 U9189 ( .A1(n8321), .A2(n8599), .ZN(n7988) );
  OR2_X1 U9190 ( .A1(n8324), .A2(n9020), .ZN(n7987) );
  NAND2_X1 U9191 ( .A1(n7991), .A2(n8616), .ZN(n7994) );
  AOI22_X1 U9192 ( .A1(n8235), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8234), .B2(
        n7992), .ZN(n7993) );
  NAND2_X1 U9193 ( .A1(n7994), .A2(n7993), .ZN(n8071) );
  OR2_X1 U9194 ( .A1(n8071), .A2(n8596), .ZN(n8686) );
  NAND2_X1 U9195 ( .A1(n8071), .A2(n8596), .ZN(n8685) );
  NAND2_X1 U9196 ( .A1(n8686), .A2(n8685), .ZN(n8781) );
  AND2_X1 U9197 ( .A1(n7997), .A2(n8670), .ZN(n8678) );
  NAND2_X1 U9198 ( .A1(n7995), .A2(n8678), .ZN(n7998) );
  NAND2_X1 U9199 ( .A1(n8679), .A2(n7996), .ZN(n8779) );
  NAND2_X1 U9200 ( .A1(n8779), .A2(n7997), .ZN(n8680) );
  AOI21_X1 U9201 ( .B1(n8781), .B2(n7999), .A(n8162), .ZN(n8000) );
  OAI222_X1 U9202 ( .A1(n9270), .A2(n8390), .B1(n9272), .B2(n8928), .C1(n9264), 
        .C2(n8000), .ZN(n10996) );
  INV_X1 U9203 ( .A(n10996), .ZN(n8012) );
  OAI22_X1 U9204 ( .A1(n10829), .A2(n8001), .B1(n8076), .B2(n10823), .ZN(n8005) );
  INV_X1 U9205 ( .A(n8071), .ZN(n10993) );
  OAI21_X1 U9206 ( .B1(n8003), .B2(n10993), .A(n8058), .ZN(n10995) );
  NOR2_X1 U9207 ( .A1(n10995), .A2(n10818), .ZN(n8004) );
  AOI211_X1 U9208 ( .C1(n9292), .C2(n8071), .A(n8005), .B(n8004), .ZN(n8011)
         );
  OR2_X1 U9209 ( .A1(n8028), .A2(n8989), .ZN(n8006) );
  NOR2_X1 U9210 ( .A1(n8008), .A2(n8781), .ZN(n10991) );
  INV_X1 U9211 ( .A(n10991), .ZN(n8009) );
  NAND3_X1 U9212 ( .A1(n8009), .A2(n10827), .A3(n10998), .ZN(n8010) );
  OAI211_X1 U9213 ( .C1(n8012), .C2(n9303), .A(n8011), .B(n8010), .ZN(P2_U3283) );
  AOI21_X1 U9214 ( .B1(n8014), .B2(n8013), .A(n5125), .ZN(n8022) );
  NOR2_X1 U9215 ( .A1(n9559), .A2(n8117), .ZN(n8015) );
  AOI211_X1 U9216 ( .C1(n9561), .C2(n9845), .A(n8016), .B(n8015), .ZN(n8017)
         );
  OAI21_X1 U9217 ( .B1(n9564), .B2(n8018), .A(n8017), .ZN(n8019) );
  AOI21_X1 U9218 ( .B1(n8020), .B2(n9566), .A(n8019), .ZN(n8021) );
  OAI21_X1 U9219 ( .B1(n8022), .B2(n9569), .A(n8021), .ZN(P1_U3234) );
  INV_X1 U9220 ( .A(n8028), .ZN(n10975) );
  XNOR2_X1 U9221 ( .A(n10970), .B(n8551), .ZN(n8024) );
  NOR2_X1 U9222 ( .A1(n8033), .A2(n8562), .ZN(n8025) );
  NAND2_X1 U9223 ( .A1(n8024), .A2(n8025), .ZN(n8035) );
  INV_X1 U9224 ( .A(n8024), .ZN(n8034) );
  INV_X1 U9225 ( .A(n8025), .ZN(n8026) );
  NAND2_X1 U9226 ( .A1(n8034), .A2(n8026), .ZN(n8027) );
  NAND2_X1 U9227 ( .A1(n8035), .A2(n8027), .ZN(n8924) );
  XNOR2_X1 U9228 ( .A(n8028), .B(n8551), .ZN(n8029) );
  NOR2_X1 U9229 ( .A1(n8928), .A2(n8562), .ZN(n8030) );
  NAND2_X1 U9230 ( .A1(n8029), .A2(n8030), .ZN(n8072) );
  INV_X1 U9231 ( .A(n8029), .ZN(n8068) );
  INV_X1 U9232 ( .A(n8030), .ZN(n8031) );
  NAND2_X1 U9233 ( .A1(n8068), .A2(n8031), .ZN(n8032) );
  AOI21_X1 U9234 ( .B1(n5111), .B2(n5121), .A(n8953), .ZN(n8037) );
  NOR3_X1 U9235 ( .A1(n8034), .A2(n8033), .A3(n8922), .ZN(n8036) );
  OAI21_X1 U9236 ( .B1(n8037), .B2(n8036), .A(n8074), .ZN(n8042) );
  OAI22_X1 U9237 ( .A1(n8964), .A2(n8596), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10302), .ZN(n8040) );
  NOR2_X1 U9238 ( .A1(n8968), .A2(n8038), .ZN(n8039) );
  AOI211_X1 U9239 ( .C1(n8966), .C2(n8990), .A(n8040), .B(n8039), .ZN(n8041)
         );
  OAI211_X1 U9240 ( .C1(n10975), .C2(n8963), .A(n8042), .B(n8041), .ZN(
        P2_U3226) );
  NAND2_X1 U9241 ( .A1(n5460), .A2(n8685), .ZN(n8046) );
  AOI22_X1 U9242 ( .A1(n8235), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8234), .B2(
        n9014), .ZN(n8044) );
  NAND2_X1 U9243 ( .A1(n9389), .A2(n8390), .ZN(n8688) );
  INV_X1 U9244 ( .A(n8161), .ZN(n8784) );
  XNOR2_X1 U9245 ( .A(n8046), .B(n8784), .ZN(n8056) );
  NAND2_X1 U9246 ( .A1(n8047), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8055) );
  INV_X1 U9247 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8048) );
  OR2_X1 U9248 ( .A1(n8253), .A2(n8048), .ZN(n8054) );
  INV_X1 U9249 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10545) );
  NAND2_X1 U9250 ( .A1(n8049), .A2(n10545), .ZN(n8050) );
  NAND2_X1 U9251 ( .A1(n8163), .A2(n8050), .ZN(n8969) );
  OR2_X1 U9252 ( .A1(n8321), .A2(n8969), .ZN(n8053) );
  INV_X1 U9253 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8051) );
  OR2_X1 U9254 ( .A1(n8324), .A2(n8051), .ZN(n8052) );
  INV_X1 U9255 ( .A(n8881), .ZN(n8986) );
  INV_X1 U9256 ( .A(n8596), .ZN(n8988) );
  AOI222_X1 U9257 ( .A1(n10822), .A2(n8056), .B1(n8986), .B2(n10821), .C1(
        n8988), .C2(n9254), .ZN(n9392) );
  OR2_X2 U9258 ( .A1(n8058), .A2(n9389), .ZN(n8356) );
  INV_X1 U9259 ( .A(n8356), .ZN(n8057) );
  AOI21_X1 U9260 ( .B1(n9389), .B2(n8058), .A(n8057), .ZN(n9390) );
  INV_X1 U9261 ( .A(n9389), .ZN(n8059) );
  NOR2_X1 U9262 ( .A1(n8059), .A2(n10819), .ZN(n8062) );
  OAI22_X1 U9263 ( .A1(n10829), .A2(n8060), .B1(n8599), .B2(n10823), .ZN(n8061) );
  AOI211_X1 U9264 ( .C1(n9390), .C2(n9226), .A(n8062), .B(n8061), .ZN(n8067)
         );
  NAND2_X1 U9265 ( .A1(n8071), .A2(n8988), .ZN(n8063) );
  OAI21_X1 U9266 ( .B1(n8065), .B2(n8161), .A(n8153), .ZN(n9388) );
  NAND2_X1 U9267 ( .A1(n9388), .A2(n10827), .ZN(n8066) );
  OAI211_X1 U9268 ( .C1(n9392), .C2(n9303), .A(n8067), .B(n8066), .ZN(P2_U3282) );
  INV_X1 U9269 ( .A(n8074), .ZN(n8070) );
  NOR3_X1 U9270 ( .A1(n8068), .A2(n8928), .A3(n8922), .ZN(n8069) );
  AOI21_X1 U9271 ( .B1(n8070), .B2(n8915), .A(n8069), .ZN(n8083) );
  XNOR2_X1 U9272 ( .A(n8071), .B(n8563), .ZN(n8391) );
  NOR2_X1 U9273 ( .A1(n8596), .A2(n8562), .ZN(n8393) );
  XNOR2_X1 U9274 ( .A(n8391), .B(n8393), .ZN(n8082) );
  INV_X1 U9275 ( .A(n8392), .ZN(n8603) );
  INV_X1 U9276 ( .A(n8390), .ZN(n8987) );
  OAI21_X1 U9277 ( .B1(n8930), .B2(n8928), .A(n8075), .ZN(n8078) );
  NOR2_X1 U9278 ( .A1(n8968), .A2(n8076), .ZN(n8077) );
  AOI211_X1 U9279 ( .C1(n8960), .C2(n8987), .A(n8078), .B(n8077), .ZN(n8079)
         );
  OAI21_X1 U9280 ( .B1(n10993), .B2(n8963), .A(n8079), .ZN(n8080) );
  AOI21_X1 U9281 ( .B1(n8603), .B2(n8915), .A(n8080), .ZN(n8081) );
  OAI21_X1 U9282 ( .B1(n8083), .B2(n8082), .A(n8081), .ZN(P2_U3236) );
  AND2_X1 U9283 ( .A1(n9684), .A2(n9678), .ZN(n9620) );
  NAND2_X1 U9284 ( .A1(n8085), .A2(n9686), .ZN(n8116) );
  OR2_X1 U9285 ( .A1(n8146), .A2(n8106), .ZN(n9685) );
  NAND2_X1 U9286 ( .A1(n8146), .A2(n8106), .ZN(n9683) );
  OR2_X2 U9287 ( .A1(n10228), .A2(n8140), .ZN(n9698) );
  NAND2_X1 U9288 ( .A1(n10228), .A2(n8140), .ZN(n9694) );
  AOI21_X1 U9289 ( .B1(n8086), .B2(n9780), .A(n9972), .ZN(n8088) );
  OAI22_X1 U9290 ( .A1(n8106), .A2(n10081), .B1(n9429), .B2(n10083), .ZN(n8087) );
  AOI21_X1 U9291 ( .B1(n8088), .B2(n8178), .A(n8087), .ZN(n10230) );
  INV_X1 U9292 ( .A(n8124), .ZN(n8089) );
  INV_X1 U9293 ( .A(n10228), .ZN(n8090) );
  NAND2_X1 U9294 ( .A1(n8124), .A2(n8090), .ZN(n8183) );
  INV_X1 U9295 ( .A(n8183), .ZN(n8184) );
  AOI211_X1 U9296 ( .C1(n10228), .C2(n8089), .A(n11009), .B(n8184), .ZN(n10227) );
  NOR2_X1 U9297 ( .A1(n8090), .A2(n10144), .ZN(n8093) );
  OAI22_X1 U9298 ( .A1(n10093), .A2(n8091), .B1(n9433), .B2(n10090), .ZN(n8092) );
  AOI211_X1 U9299 ( .C1(n10227), .C2(n10138), .A(n8093), .B(n8092), .ZN(n8099)
         );
  NAND2_X1 U9300 ( .A1(n10233), .A2(n9843), .ZN(n8094) );
  NAND2_X1 U9301 ( .A1(n8115), .A2(n5618), .ZN(n8114) );
  INV_X1 U9302 ( .A(n8106), .ZN(n9842) );
  OR2_X1 U9303 ( .A1(n8146), .A2(n9842), .ZN(n8096) );
  NAND2_X1 U9304 ( .A1(n8114), .A2(n8096), .ZN(n8097) );
  OAI21_X1 U9305 ( .B1(n8097), .B2(n9780), .A(n8174), .ZN(n10226) );
  NAND2_X1 U9306 ( .A1(n10226), .A2(n9929), .ZN(n8098) );
  OAI211_X1 U9307 ( .C1(n10230), .C2(n10141), .A(n8099), .B(n8098), .ZN(
        P1_U3277) );
  INV_X1 U9308 ( .A(n8100), .ZN(n8102) );
  NOR2_X1 U9309 ( .A1(n8102), .A2(n8101), .ZN(n8103) );
  XNOR2_X1 U9310 ( .A(n8104), .B(n8103), .ZN(n8113) );
  INV_X1 U9311 ( .A(n8105), .ZN(n8108) );
  NOR2_X1 U9312 ( .A1(n9559), .A2(n8106), .ZN(n8107) );
  AOI211_X1 U9313 ( .C1(n9561), .C2(n9844), .A(n8108), .B(n8107), .ZN(n8109)
         );
  OAI21_X1 U9314 ( .B1(n9564), .B2(n8110), .A(n8109), .ZN(n8111) );
  AOI21_X1 U9315 ( .B1(n10233), .B2(n9566), .A(n8111), .ZN(n8112) );
  OAI21_X1 U9316 ( .B1(n8113), .B2(n9569), .A(n8112), .ZN(P1_U3222) );
  OAI21_X1 U9317 ( .B1(n8115), .B2(n5618), .A(n8114), .ZN(n10987) );
  INV_X1 U9318 ( .A(n10987), .ZN(n8129) );
  XOR2_X1 U9319 ( .A(n8116), .B(n9778), .Z(n8120) );
  OAI22_X1 U9320 ( .A1(n8117), .A2(n10081), .B1(n8140), .B2(n10083), .ZN(n8118) );
  AOI21_X1 U9321 ( .B1(n10987), .B2(n10929), .A(n8118), .ZN(n8119) );
  OAI21_X1 U9322 ( .B1(n9972), .B2(n8120), .A(n8119), .ZN(n10985) );
  NAND2_X1 U9323 ( .A1(n10985), .A2(n10093), .ZN(n8128) );
  OAI22_X1 U9324 ( .A1(n10093), .A2(n8121), .B1(n8144), .B2(n10090), .ZN(n8126) );
  NOR2_X1 U9325 ( .A1(n8122), .A2(n10983), .ZN(n8123) );
  OR2_X1 U9326 ( .A1(n8124), .A2(n8123), .ZN(n10984) );
  NOR2_X1 U9327 ( .A1(n10984), .A2(n10098), .ZN(n8125) );
  AOI211_X1 U9328 ( .C1(n10095), .C2(n8146), .A(n8126), .B(n8125), .ZN(n8127)
         );
  OAI211_X1 U9329 ( .C1(n8129), .C2(n10055), .A(n8128), .B(n8127), .ZN(
        P1_U3278) );
  INV_X1 U9330 ( .A(n8290), .ZN(n8132) );
  OAI222_X1 U9331 ( .A1(P1_U3084), .A2(n8130), .B1(n10265), .B2(n8132), .C1(
        n10443), .C2(n10267), .ZN(P1_U3328) );
  OAI222_X1 U9332 ( .A1(n5036), .A2(n8291), .B1(n8494), .B2(n8132), .C1(
        P2_U3152), .C2(n8131), .ZN(P2_U3333) );
  INV_X1 U9333 ( .A(n8300), .ZN(n8134) );
  OAI222_X1 U9334 ( .A1(n8494), .A2(n8134), .B1(n8133), .B2(P2_U3152), .C1(
        n8301), .C2(n5036), .ZN(P2_U3332) );
  OAI222_X1 U9335 ( .A1(n8135), .A2(P1_U3084), .B1(n10265), .B2(n8134), .C1(
        n10445), .C2(n10267), .ZN(P1_U3327) );
  XNOR2_X1 U9336 ( .A(n5153), .B(n8136), .ZN(n8137) );
  XNOR2_X1 U9337 ( .A(n8138), .B(n8137), .ZN(n8148) );
  INV_X1 U9338 ( .A(n8139), .ZN(n8142) );
  NOR2_X1 U9339 ( .A1(n9559), .A2(n8140), .ZN(n8141) );
  AOI211_X1 U9340 ( .C1(n9561), .C2(n9843), .A(n8142), .B(n8141), .ZN(n8143)
         );
  OAI21_X1 U9341 ( .B1(n9564), .B2(n8144), .A(n8143), .ZN(n8145) );
  AOI21_X1 U9342 ( .B1(n8146), .B2(n9566), .A(n8145), .ZN(n8147) );
  OAI21_X1 U9343 ( .B1(n8148), .B2(n9569), .A(n8147), .ZN(P1_U3232) );
  INV_X1 U9344 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10446) );
  NAND2_X1 U9345 ( .A1(n8315), .A2(n10660), .ZN(n8150) );
  OAI211_X1 U9346 ( .C1(n10267), .C2(n10446), .A(n8150), .B(n8149), .ZN(
        P1_U3326) );
  INV_X1 U9347 ( .A(n8315), .ZN(n8151) );
  INV_X1 U9348 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8316) );
  OAI222_X1 U9349 ( .A1(n8494), .A2(n8151), .B1(P2_U3152), .B2(n8375), .C1(
        n8316), .C2(n5036), .ZN(P2_U3331) );
  OR2_X1 U9350 ( .A1(n9389), .A2(n8987), .ZN(n8152) );
  NAND2_X1 U9351 ( .A1(n8153), .A2(n8152), .ZN(n8207) );
  NAND2_X1 U9352 ( .A1(n8154), .A2(n8616), .ZN(n8156) );
  AOI22_X1 U9353 ( .A1(n8235), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8234), .B2(
        n9034), .ZN(n8155) );
  OR2_X1 U9354 ( .A1(n9383), .A2(n8881), .ZN(n8692) );
  NAND2_X1 U9355 ( .A1(n9383), .A2(n8881), .ZN(n8691) );
  XNOR2_X1 U9356 ( .A(n8207), .B(n8785), .ZN(n9387) );
  XOR2_X1 U9357 ( .A(n9383), .B(n8356), .Z(n9384) );
  INV_X1 U9358 ( .A(n9383), .ZN(n8159) );
  INV_X1 U9359 ( .A(n8969), .ZN(n8157) );
  AOI22_X1 U9360 ( .A1(n9303), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8157), .B2(
        n9202), .ZN(n8158) );
  OAI21_X1 U9361 ( .B1(n8159), .B2(n10819), .A(n8158), .ZN(n8171) );
  INV_X1 U9362 ( .A(n8685), .ZN(n8160) );
  XNOR2_X1 U9363 ( .A(n5114), .B(n8785), .ZN(n8169) );
  NAND2_X1 U9364 ( .A1(n8047), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8168) );
  INV_X1 U9365 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9290) );
  OR2_X1 U9366 ( .A1(n8253), .A2(n9290), .ZN(n8167) );
  INV_X1 U9367 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10300) );
  NAND2_X1 U9368 ( .A1(n8163), .A2(n10300), .ZN(n8164) );
  NAND2_X1 U9369 ( .A1(n8216), .A2(n8164), .ZN(n9289) );
  OR2_X1 U9370 ( .A1(n8321), .A2(n9289), .ZN(n8166) );
  INV_X1 U9371 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9046) );
  OR2_X1 U9372 ( .A1(n8324), .A2(n9046), .ZN(n8165) );
  INV_X1 U9373 ( .A(n9273), .ZN(n8985) );
  AOI222_X1 U9374 ( .A1(n10822), .A2(n8169), .B1(n8985), .B2(n10821), .C1(
        n8987), .C2(n9254), .ZN(n9386) );
  NOR2_X1 U9375 ( .A1(n9386), .A2(n9303), .ZN(n8170) );
  AOI211_X1 U9376 ( .C1(n9384), .C2(n9226), .A(n8171), .B(n8170), .ZN(n8172)
         );
  OAI21_X1 U9377 ( .B1(n9387), .B2(n9300), .A(n8172), .ZN(P2_U3281) );
  OR2_X1 U9378 ( .A1(n10228), .A2(n9841), .ZN(n8173) );
  NAND2_X1 U9379 ( .A1(n9567), .A2(n9429), .ZN(n9695) );
  INV_X1 U9380 ( .A(n9782), .ZN(n8175) );
  NAND2_X1 U9381 ( .A1(n8176), .A2(n9782), .ZN(n8177) );
  NAND2_X1 U9382 ( .A1(n8470), .A2(n8177), .ZN(n11007) );
  AOI22_X1 U9383 ( .A1(n9841), .A2(n10131), .B1(n10130), .B2(n10109), .ZN(
        n8181) );
  NAND2_X1 U9384 ( .A1(n8179), .A2(n9782), .ZN(n8447) );
  OAI211_X1 U9385 ( .C1(n9782), .C2(n8179), .A(n8447), .B(n10125), .ZN(n8180)
         );
  OAI211_X1 U9386 ( .C1(n11007), .C2(n7255), .A(n8181), .B(n8180), .ZN(n11011)
         );
  NAND2_X1 U9387 ( .A1(n11011), .A2(n10093), .ZN(n8188) );
  OAI22_X1 U9388 ( .A1(n10093), .A2(n8182), .B1(n9563), .B2(n10090), .ZN(n8186) );
  OR2_X2 U9389 ( .A1(n8183), .A2(n9567), .ZN(n10137) );
  OAI21_X1 U9390 ( .B1(n8184), .B2(n11008), .A(n10137), .ZN(n11010) );
  NOR2_X1 U9391 ( .A1(n11010), .A2(n10098), .ZN(n8185) );
  AOI211_X1 U9392 ( .C1(n10095), .C2(n9567), .A(n8186), .B(n8185), .ZN(n8187)
         );
  OAI211_X1 U9393 ( .C1(n11007), .C2(n10055), .A(n8188), .B(n8187), .ZN(
        P1_U3276) );
  INV_X1 U9394 ( .A(n8189), .ZN(n8192) );
  NAND2_X1 U9395 ( .A1(n8190), .A2(SI_27_), .ZN(n8191) );
  MUX2_X1 U9396 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n5663), .Z(n8340) );
  XNOR2_X1 U9397 ( .A(n8340), .B(SI_28_), .ZN(n8338) );
  INV_X1 U9398 ( .A(n8413), .ZN(n8196) );
  AOI21_X1 U9399 ( .B1(n10658), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n8194), .ZN(
        n8195) );
  OAI21_X1 U9400 ( .B1(n8196), .B2(n10265), .A(n8195), .ZN(P1_U3325) );
  INV_X1 U9401 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8329) );
  OAI222_X1 U9402 ( .A1(n5036), .A2(n8329), .B1(n8494), .B2(n8196), .C1(n6582), 
        .C2(P2_U3152), .ZN(P2_U3330) );
  NAND2_X1 U9403 ( .A1(n8252), .A2(n10357), .ZN(n8197) );
  AND2_X1 U9404 ( .A1(n8264), .A2(n8197), .ZN(n9203) );
  NAND2_X1 U9405 ( .A1(n9203), .A2(n8353), .ZN(n8202) );
  NAND2_X1 U9406 ( .A1(n8370), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8199) );
  NAND2_X1 U9407 ( .A1(n8047), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8198) );
  AND2_X1 U9408 ( .A1(n8199), .A2(n8198), .ZN(n8201) );
  NAND2_X1 U9409 ( .A1(n8266), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U9410 ( .A1(n8203), .A2(n8616), .ZN(n8205) );
  OR2_X1 U9411 ( .A1(n5039), .A2(n7658), .ZN(n8204) );
  INV_X1 U9412 ( .A(n9352), .ZN(n9205) );
  INV_X1 U9413 ( .A(n8785), .ZN(n8206) );
  NAND2_X1 U9414 ( .A1(n8208), .A2(n8616), .ZN(n8210) );
  AOI22_X1 U9415 ( .A1(n8235), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8234), .B2(
        n9054), .ZN(n8209) );
  OR2_X1 U9416 ( .A1(n9379), .A2(n9273), .ZN(n8698) );
  AND2_X1 U9417 ( .A1(n9379), .A2(n9273), .ZN(n8361) );
  INV_X1 U9418 ( .A(n8361), .ZN(n8697) );
  NAND2_X1 U9419 ( .A1(n9288), .A2(n8211), .ZN(n9287) );
  NAND2_X1 U9420 ( .A1(n9379), .A2(n8985), .ZN(n8212) );
  NAND2_X1 U9421 ( .A1(n8213), .A2(n8616), .ZN(n8215) );
  AOI22_X1 U9422 ( .A1(n8235), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8234), .B2(
        n9061), .ZN(n8214) );
  NAND2_X1 U9423 ( .A1(n8047), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8221) );
  NAND2_X1 U9424 ( .A1(n8216), .A2(n10361), .ZN(n8217) );
  NAND2_X1 U9425 ( .A1(n8225), .A2(n8217), .ZN(n9276) );
  OR2_X1 U9426 ( .A1(n8321), .A2(n9276), .ZN(n8220) );
  INV_X1 U9427 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9067) );
  OR2_X1 U9428 ( .A1(n8324), .A2(n9067), .ZN(n8219) );
  INV_X1 U9429 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9277) );
  OR2_X1 U9430 ( .A1(n8253), .A2(n9277), .ZN(n8218) );
  NAND4_X1 U9431 ( .A1(n8221), .A2(n8220), .A3(n8219), .A4(n8218), .ZN(n9253)
         );
  XNOR2_X1 U9432 ( .A(n9375), .B(n9253), .ZN(n8764) );
  NAND2_X1 U9433 ( .A1(n8222), .A2(n8616), .ZN(n8224) );
  AOI22_X1 U9434 ( .A1(n8235), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8234), .B2(
        n9073), .ZN(n8223) );
  NAND2_X1 U9435 ( .A1(n8047), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8231) );
  INV_X1 U9436 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9373) );
  OR2_X1 U9437 ( .A1(n8324), .A2(n9373), .ZN(n8230) );
  INV_X1 U9438 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10540) );
  NAND2_X1 U9439 ( .A1(n8225), .A2(n10540), .ZN(n8226) );
  NAND2_X1 U9440 ( .A1(n8238), .A2(n8226), .ZN(n9257) );
  OR2_X1 U9441 ( .A1(n8321), .A2(n9257), .ZN(n8229) );
  INV_X1 U9442 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8227) );
  OR2_X1 U9443 ( .A1(n8253), .A2(n8227), .ZN(n8228) );
  OR2_X1 U9444 ( .A1(n9369), .A2(n9271), .ZN(n8706) );
  NAND2_X1 U9445 ( .A1(n9369), .A2(n9271), .ZN(n8705) );
  INV_X1 U9446 ( .A(n9271), .ZN(n8984) );
  OR2_X1 U9447 ( .A1(n9369), .A2(n8984), .ZN(n8232) );
  NAND2_X1 U9448 ( .A1(n10661), .A2(n8616), .ZN(n8237) );
  AOI22_X1 U9449 ( .A1(n8235), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8234), .B2(
        n8233), .ZN(n8236) );
  NAND2_X1 U9450 ( .A1(n8238), .A2(n10524), .ZN(n8239) );
  NAND2_X1 U9451 ( .A1(n8250), .A2(n8239), .ZN(n9239) );
  OR2_X1 U9452 ( .A1(n8321), .A2(n9239), .ZN(n8244) );
  INV_X1 U9453 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8240) );
  OR2_X1 U9454 ( .A1(n8253), .A2(n8240), .ZN(n8243) );
  INV_X1 U9455 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9367) );
  OR2_X1 U9456 ( .A1(n8324), .A2(n9367), .ZN(n8242) );
  INV_X1 U9457 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9407) );
  OR2_X1 U9458 ( .A1(n6730), .A2(n9407), .ZN(n8241) );
  NAND4_X1 U9459 ( .A1(n8244), .A2(n8243), .A3(n8242), .A4(n8241), .ZN(n9252)
         );
  XNOR2_X1 U9460 ( .A(n9361), .B(n9252), .ZN(n9229) );
  INV_X1 U9461 ( .A(n9252), .ZN(n9212) );
  NAND2_X1 U9462 ( .A1(n9231), .A2(n5644), .ZN(n9216) );
  NAND2_X1 U9463 ( .A1(n8245), .A2(n8616), .ZN(n8248) );
  OR2_X1 U9464 ( .A1(n5038), .A2(n8246), .ZN(n8247) );
  INV_X1 U9465 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8249) );
  NAND2_X1 U9466 ( .A1(n8250), .A2(n8249), .ZN(n8251) );
  NAND2_X1 U9467 ( .A1(n8252), .A2(n8251), .ZN(n9222) );
  OR2_X1 U9468 ( .A1(n9222), .A2(n8321), .ZN(n8259) );
  INV_X1 U9469 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9223) );
  OR2_X1 U9470 ( .A1(n8253), .A2(n9223), .ZN(n8258) );
  INV_X1 U9471 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8254) );
  OR2_X1 U9472 ( .A1(n6730), .A2(n8254), .ZN(n8257) );
  INV_X1 U9473 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8255) );
  OR2_X1 U9474 ( .A1(n8324), .A2(n8255), .ZN(n8256) );
  NAND2_X1 U9475 ( .A1(n9357), .A2(n9233), .ZN(n8712) );
  NAND2_X1 U9476 ( .A1(n9352), .A2(n9213), .ZN(n8719) );
  NAND2_X1 U9477 ( .A1(n8260), .A2(n8616), .ZN(n8263) );
  OR2_X1 U9478 ( .A1(n5038), .A2(n8261), .ZN(n8262) );
  INV_X1 U9479 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10291) );
  NAND2_X1 U9480 ( .A1(n8264), .A2(n10291), .ZN(n8265) );
  NAND2_X1 U9481 ( .A1(n8281), .A2(n8265), .ZN(n9181) );
  OR2_X1 U9482 ( .A1(n9181), .A2(n8321), .ZN(n8269) );
  AOI22_X1 U9483 ( .A1(n8370), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8047), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n8268) );
  NAND2_X1 U9484 ( .A1(n8266), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8267) );
  NAND2_X1 U9485 ( .A1(n9347), .A2(n8530), .ZN(n8723) );
  NAND2_X1 U9486 ( .A1(n8722), .A2(n8723), .ZN(n9185) );
  INV_X1 U9487 ( .A(n9185), .ZN(n8789) );
  OAI22_X1 U9488 ( .A1(n9179), .A2(n8789), .B1(n9197), .B2(n9347), .ZN(n9171)
         );
  NAND2_X1 U9489 ( .A1(n8270), .A2(n8616), .ZN(n8273) );
  OR2_X1 U9490 ( .A1(n5039), .A2(n8271), .ZN(n8272) );
  NAND2_X1 U9491 ( .A1(n9175), .A2(n9155), .ZN(n8725) );
  INV_X1 U9492 ( .A(n9155), .ZN(n9187) );
  NAND2_X1 U9493 ( .A1(n9341), .A2(n9187), .ZN(n8622) );
  NAND2_X1 U9494 ( .A1(n8725), .A2(n8622), .ZN(n8791) );
  NOR2_X1 U9495 ( .A1(n9170), .A2(n8274), .ZN(n9150) );
  NAND2_X1 U9496 ( .A1(n8275), .A2(n8616), .ZN(n8278) );
  OR2_X1 U9497 ( .A1(n5038), .A2(n8276), .ZN(n8277) );
  INV_X1 U9498 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8280) );
  INV_X1 U9499 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8279) );
  OAI21_X1 U9500 ( .B1(n8281), .B2(n8280), .A(n8279), .ZN(n8282) );
  NAND2_X1 U9501 ( .A1(n8282), .A2(n8294), .ZN(n8894) );
  OR2_X1 U9502 ( .A1(n8894), .A2(n8321), .ZN(n8288) );
  INV_X1 U9503 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8285) );
  NAND2_X1 U9504 ( .A1(n8047), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8284) );
  NAND2_X1 U9505 ( .A1(n8370), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8283) );
  OAI211_X1 U9506 ( .C1(n8324), .C2(n8285), .A(n8284), .B(n8283), .ZN(n8286)
         );
  INV_X1 U9507 ( .A(n8286), .ZN(n8287) );
  NAND2_X1 U9508 ( .A1(n9162), .A2(n8890), .ZN(n8730) );
  NAND2_X1 U9509 ( .A1(n9150), .A2(n9152), .ZN(n9151) );
  INV_X1 U9510 ( .A(n8890), .ZN(n9168) );
  NAND2_X1 U9511 ( .A1(n8290), .A2(n8616), .ZN(n8293) );
  OR2_X1 U9512 ( .A1(n5038), .A2(n8291), .ZN(n8292) );
  INV_X1 U9513 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10461) );
  NAND2_X1 U9514 ( .A1(n8294), .A2(n10461), .ZN(n8295) );
  INV_X1 U9515 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8298) );
  NAND2_X1 U9516 ( .A1(n8047), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8297) );
  NAND2_X1 U9517 ( .A1(n8370), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8296) );
  OAI211_X1 U9518 ( .C1(n8298), .C2(n8324), .A(n8297), .B(n8296), .ZN(n8299)
         );
  NAND2_X1 U9519 ( .A1(n9330), .A2(n9158), .ZN(n8732) );
  INV_X1 U9520 ( .A(n9330), .ZN(n9140) );
  NAND2_X1 U9521 ( .A1(n8300), .A2(n8616), .ZN(n8303) );
  OR2_X1 U9522 ( .A1(n5039), .A2(n8301), .ZN(n8302) );
  INV_X1 U9523 ( .A(n8306), .ZN(n8304) );
  NAND2_X1 U9524 ( .A1(n8304), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8319) );
  INV_X1 U9525 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8305) );
  NAND2_X1 U9526 ( .A1(n8306), .A2(n8305), .ZN(n8307) );
  NAND2_X1 U9527 ( .A1(n8319), .A2(n8307), .ZN(n9127) );
  INV_X1 U9528 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8310) );
  NAND2_X1 U9529 ( .A1(n8047), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8309) );
  NAND2_X1 U9530 ( .A1(n8370), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8308) );
  OAI211_X1 U9531 ( .C1(n8324), .C2(n8310), .A(n8309), .B(n8308), .ZN(n8311)
         );
  INV_X1 U9532 ( .A(n8311), .ZN(n8312) );
  OR2_X1 U9533 ( .A1(n9133), .A2(n8871), .ZN(n8368) );
  INV_X1 U9534 ( .A(n8368), .ZN(n8314) );
  NAND2_X1 U9535 ( .A1(n8315), .A2(n8616), .ZN(n8318) );
  OR2_X1 U9536 ( .A1(n5039), .A2(n8316), .ZN(n8317) );
  INV_X1 U9537 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10520) );
  NAND2_X1 U9538 ( .A1(n8319), .A2(n10520), .ZN(n8320) );
  NAND2_X1 U9539 ( .A1(n8332), .A2(n8320), .ZN(n9103) );
  INV_X1 U9540 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8325) );
  NAND2_X1 U9541 ( .A1(n8370), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8323) );
  NAND2_X1 U9542 ( .A1(n8047), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8322) );
  OAI211_X1 U9543 ( .C1(n8325), .C2(n8324), .A(n8323), .B(n8322), .ZN(n8326)
         );
  INV_X1 U9544 ( .A(n8326), .ZN(n8327) );
  NAND2_X1 U9545 ( .A1(n9321), .A2(n9122), .ZN(n8748) );
  NAND2_X1 U9546 ( .A1(n8744), .A2(n8748), .ZN(n8742) );
  NAND2_X1 U9547 ( .A1(n8413), .A2(n8616), .ZN(n8331) );
  OR2_X1 U9548 ( .A1(n5039), .A2(n8329), .ZN(n8330) );
  INV_X1 U9549 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U9550 ( .A1(n8332), .A2(n8573), .ZN(n8333) );
  INV_X1 U9551 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8336) );
  NAND2_X1 U9552 ( .A1(n8047), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8335) );
  NAND2_X1 U9553 ( .A1(n8370), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8334) );
  OAI211_X1 U9554 ( .C1(n8324), .C2(n8336), .A(n8335), .B(n8334), .ZN(n8337)
         );
  NAND2_X1 U9555 ( .A1(n9316), .A2(n8833), .ZN(n8746) );
  INV_X1 U9556 ( .A(n8833), .ZN(n8979) );
  INV_X1 U9557 ( .A(n8340), .ZN(n8341) );
  NAND2_X1 U9558 ( .A1(n8341), .A2(n10479), .ZN(n8342) );
  MUX2_X1 U9559 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n5668), .Z(n8498) );
  INV_X1 U9560 ( .A(n8343), .ZN(n8344) );
  NAND2_X1 U9561 ( .A1(n8344), .A2(n10316), .ZN(n8345) );
  INV_X1 U9562 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9422) );
  OR2_X1 U9563 ( .A1(n5038), .A2(n9422), .ZN(n8346) );
  INV_X1 U9564 ( .A(n9311), .ZN(n8359) );
  INV_X1 U9565 ( .A(n8348), .ZN(n8357) );
  INV_X1 U9566 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8351) );
  NAND2_X1 U9567 ( .A1(n8370), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8350) );
  NAND2_X1 U9568 ( .A1(n8047), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8349) );
  OAI211_X1 U9569 ( .C1(n8351), .C2(n8324), .A(n8350), .B(n8349), .ZN(n8352)
         );
  AOI21_X1 U9570 ( .B1(n8357), .B2(n8353), .A(n8352), .ZN(n8588) );
  INV_X1 U9571 ( .A(n8588), .ZN(n8978) );
  NAND2_X1 U9572 ( .A1(n8359), .A2(n8978), .ZN(n8806) );
  NAND2_X1 U9573 ( .A1(n9311), .A2(n8588), .ZN(n8804) );
  NAND2_X1 U9574 ( .A1(n8806), .A2(n8804), .ZN(n8795) );
  INV_X1 U9575 ( .A(n8795), .ZN(n8354) );
  NOR2_X1 U9576 ( .A1(n8356), .A2(n9383), .ZN(n9294) );
  INV_X1 U9577 ( .A(n9379), .ZN(n9293) );
  NAND2_X1 U9578 ( .A1(n9294), .A2(n9293), .ZN(n9296) );
  OR2_X2 U9579 ( .A1(n9201), .A2(n9352), .ZN(n9199) );
  AND2_X1 U9580 ( .A1(n9180), .A2(n9175), .ZN(n9160) );
  NAND2_X1 U9581 ( .A1(n9160), .A2(n9334), .ZN(n9159) );
  OR2_X2 U9582 ( .A1(n9159), .A2(n9330), .ZN(n9128) );
  NOR2_X2 U9583 ( .A1(n9128), .A2(n9133), .ZN(n9129) );
  AOI21_X1 U9584 ( .B1(n9311), .B2(n8579), .A(n9097), .ZN(n9312) );
  AOI22_X1 U9585 ( .A1(n8357), .A2(n9202), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n9303), .ZN(n8358) );
  OAI21_X1 U9586 ( .B1(n8359), .B2(n10819), .A(n8358), .ZN(n8378) );
  INV_X1 U9587 ( .A(n8692), .ZN(n8360) );
  INV_X1 U9588 ( .A(n9253), .ZN(n8362) );
  OR2_X1 U9589 ( .A1(n9375), .A2(n8362), .ZN(n8363) );
  NAND2_X1 U9590 ( .A1(n9236), .A2(n9252), .ZN(n8365) );
  NAND2_X1 U9591 ( .A1(n8366), .A2(n8365), .ZN(n9211) );
  NAND2_X1 U9592 ( .A1(n8367), .A2(n8789), .ZN(n9189) );
  AND2_X1 U9593 ( .A1(n8368), .A2(n9118), .ZN(n8736) );
  NAND2_X1 U9594 ( .A1(n9145), .A2(n8736), .ZN(n9109) );
  NOR2_X1 U9595 ( .A1(n8742), .A2(n8737), .ZN(n8369) );
  NAND2_X1 U9596 ( .A1(n9109), .A2(n8369), .ZN(n9107) );
  NAND2_X1 U9597 ( .A1(n9107), .A2(n8744), .ZN(n8585) );
  NAND2_X1 U9598 ( .A1(n8590), .A2(n8749), .ZN(n8805) );
  XNOR2_X1 U9599 ( .A(n8805), .B(n8795), .ZN(n8377) );
  INV_X1 U9600 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8373) );
  NAND2_X1 U9601 ( .A1(n8370), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8372) );
  NAND2_X1 U9602 ( .A1(n8047), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8371) );
  OAI211_X1 U9603 ( .C1(n8324), .C2(n8373), .A(n8372), .B(n8371), .ZN(n8977)
         );
  NOR2_X1 U9604 ( .A1(n8375), .A2(n10547), .ZN(n8376) );
  NOR2_X1 U9605 ( .A1(n9270), .A2(n8376), .ZN(n9093) );
  NAND2_X1 U9606 ( .A1(n8380), .A2(n8379), .ZN(n8381) );
  XOR2_X1 U9607 ( .A(n8382), .B(n8381), .Z(n8389) );
  OAI22_X1 U9608 ( .A1(n8383), .A2(n9559), .B1(n9535), .B2(n7411), .ZN(n8384)
         );
  AOI211_X1 U9609 ( .C1(n9561), .C2(n7246), .A(n8385), .B(n8384), .ZN(n8388)
         );
  NAND2_X1 U9610 ( .A1(n9505), .A2(n8386), .ZN(n8387) );
  OAI211_X1 U9611 ( .C1(n8389), .C2(n9569), .A(n8388), .B(n8387), .ZN(P1_U3228) );
  NOR2_X1 U9612 ( .A1(n8390), .A2(n8562), .ZN(n8397) );
  XNOR2_X1 U9613 ( .A(n9389), .B(n8563), .ZN(n8394) );
  INV_X1 U9614 ( .A(n8394), .ZN(n8396) );
  INV_X1 U9615 ( .A(n8391), .ZN(n8600) );
  OAI21_X1 U9616 ( .B1(n8393), .B2(n8600), .A(n8392), .ZN(n8395) );
  XNOR2_X1 U9617 ( .A(n8394), .B(n8397), .ZN(n8601) );
  NAND2_X1 U9618 ( .A1(n8395), .A2(n8601), .ZN(n8607) );
  XNOR2_X1 U9619 ( .A(n9383), .B(n8551), .ZN(n8878) );
  NOR2_X1 U9620 ( .A1(n8881), .A2(n8562), .ZN(n8398) );
  NAND2_X1 U9621 ( .A1(n8878), .A2(n8398), .ZN(n8399) );
  OAI21_X1 U9622 ( .B1(n8878), .B2(n8398), .A(n8399), .ZN(n8971) );
  OR2_X2 U9623 ( .A1(n8972), .A2(n8971), .ZN(n8877) );
  XNOR2_X1 U9624 ( .A(n9379), .B(n8563), .ZN(n8401) );
  NOR2_X1 U9625 ( .A1(n9273), .A2(n8562), .ZN(n8402) );
  XNOR2_X1 U9626 ( .A(n8401), .B(n8402), .ZN(n8888) );
  INV_X1 U9627 ( .A(n8401), .ZN(n8403) );
  XNOR2_X1 U9628 ( .A(n9375), .B(n8551), .ZN(n8405) );
  AND2_X1 U9629 ( .A1(n9253), .A2(n8535), .ZN(n8404) );
  NOR2_X1 U9630 ( .A1(n8405), .A2(n8404), .ZN(n8942) );
  INV_X1 U9631 ( .A(n8942), .ZN(n8406) );
  NAND2_X1 U9632 ( .A1(n8405), .A2(n8404), .ZN(n8944) );
  NAND2_X1 U9633 ( .A1(n8406), .A2(n8944), .ZN(n8407) );
  XNOR2_X1 U9634 ( .A(n8943), .B(n8407), .ZN(n8412) );
  NAND2_X1 U9635 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9050) );
  OAI21_X1 U9636 ( .B1(n8964), .B2(n9271), .A(n9050), .ZN(n8408) );
  AOI21_X1 U9637 ( .B1(n8966), .B2(n8985), .A(n8408), .ZN(n8409) );
  OAI21_X1 U9638 ( .B1(n9276), .B2(n8968), .A(n8409), .ZN(n8410) );
  AOI21_X1 U9639 ( .B1(n9375), .B2(n8975), .A(n8410), .ZN(n8411) );
  OAI21_X1 U9640 ( .B1(n8412), .B2(n8953), .A(n8411), .ZN(P2_U3230) );
  NAND2_X1 U9641 ( .A1(n8413), .A2(n6176), .ZN(n8415) );
  NAND2_X1 U9642 ( .A1(n9574), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8414) );
  NAND2_X1 U9643 ( .A1(n10158), .A2(n8416), .ZN(n8418) );
  NAND2_X1 U9644 ( .A1(n9840), .A2(n8422), .ZN(n8417) );
  NAND2_X1 U9645 ( .A1(n8418), .A2(n8417), .ZN(n8419) );
  XNOR2_X1 U9646 ( .A(n8419), .B(n5913), .ZN(n8424) );
  NOR2_X1 U9647 ( .A1(n9934), .A2(n8420), .ZN(n8421) );
  AOI21_X1 U9648 ( .B1(n10158), .B2(n8422), .A(n8421), .ZN(n8423) );
  XNOR2_X1 U9649 ( .A(n8424), .B(n8423), .ZN(n8440) );
  INV_X1 U9650 ( .A(n8440), .ZN(n8425) );
  NAND2_X1 U9651 ( .A1(n8425), .A2(n9525), .ZN(n8446) );
  INV_X1 U9652 ( .A(n8439), .ZN(n8426) );
  AND2_X1 U9653 ( .A1(n8440), .A2(n8427), .ZN(n8428) );
  NAND2_X1 U9654 ( .A1(n5040), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8436) );
  INV_X1 U9655 ( .A(n8483), .ZN(n8429) );
  NAND2_X1 U9656 ( .A1(n5855), .A2(n8429), .ZN(n8435) );
  INV_X1 U9657 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8484) );
  OR2_X1 U9658 ( .A1(n8430), .A2(n8484), .ZN(n8434) );
  INV_X1 U9659 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8431) );
  OR2_X1 U9660 ( .A1(n8432), .A2(n8431), .ZN(n8433) );
  NAND4_X1 U9661 ( .A1(n8436), .A2(n8435), .A3(n8434), .A4(n8433), .ZN(n9912)
         );
  AOI22_X1 U9662 ( .A1(n9532), .A2(n9912), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8438) );
  NAND2_X1 U9663 ( .A1(n9561), .A2(n9953), .ZN(n8437) );
  OAI211_X1 U9664 ( .C1(n9564), .C2(n9923), .A(n8438), .B(n8437), .ZN(n8442)
         );
  NOR3_X1 U9665 ( .A1(n8440), .A2(n9569), .A3(n8439), .ZN(n8441) );
  AOI211_X1 U9666 ( .C1(n10158), .C2(n9566), .A(n8442), .B(n8441), .ZN(n8443)
         );
  OAI211_X1 U9667 ( .C1(n8446), .C2(n8445), .A(n8444), .B(n8443), .ZN(P1_U3218) );
  NAND2_X1 U9668 ( .A1(n8447), .A2(n9699), .ZN(n10128) );
  INV_X1 U9669 ( .A(n10109), .ZN(n9558) );
  NAND2_X1 U9670 ( .A1(n10223), .A2(n9558), .ZN(n9704) );
  NAND2_X1 U9671 ( .A1(n9705), .A2(n9704), .ZN(n10123) );
  INV_X1 U9672 ( .A(n10123), .ZN(n10127) );
  NAND2_X1 U9673 ( .A1(n10128), .A2(n10127), .ZN(n10126) );
  NAND2_X1 U9674 ( .A1(n10216), .A2(n10082), .ZN(n9709) );
  NAND2_X1 U9675 ( .A1(n9708), .A2(n9709), .ZN(n10104) );
  INV_X1 U9676 ( .A(n10104), .ZN(n10107) );
  OR2_X1 U9677 ( .A1(n10096), .A2(n9499), .ZN(n9712) );
  NAND2_X1 U9678 ( .A1(n10096), .A2(n9499), .ZN(n9713) );
  INV_X1 U9679 ( .A(n10073), .ZN(n10077) );
  OR2_X1 U9680 ( .A1(n10203), .A2(n10084), .ZN(n9716) );
  NAND2_X1 U9681 ( .A1(n10203), .A2(n10084), .ZN(n9715) );
  NAND2_X1 U9682 ( .A1(n9716), .A2(n9715), .ZN(n10059) );
  INV_X1 U9683 ( .A(n10059), .ZN(n10067) );
  NAND2_X1 U9684 ( .A1(n10065), .A2(n9715), .ZN(n10036) );
  OR2_X1 U9685 ( .A1(n10198), .A2(n9451), .ZN(n9614) );
  NAND2_X1 U9686 ( .A1(n10198), .A2(n9451), .ZN(n9583) );
  NAND2_X1 U9687 ( .A1(n9614), .A2(n9583), .ZN(n10042) );
  INV_X1 U9688 ( .A(n10042), .ZN(n10037) );
  NAND2_X1 U9689 ( .A1(n10036), .A2(n10037), .ZN(n10035) );
  NAND2_X1 U9690 ( .A1(n10035), .A2(n9583), .ZN(n10024) );
  OR2_X1 U9691 ( .A1(n10194), .A2(n10038), .ZN(n9615) );
  NAND2_X1 U9692 ( .A1(n10194), .A2(n10038), .ZN(n9721) );
  INV_X1 U9693 ( .A(n9721), .ZN(n8448) );
  AOI21_X2 U9694 ( .B1(n10024), .B2(n10023), .A(n8448), .ZN(n10014) );
  XNOR2_X1 U9695 ( .A(n10188), .B(n9470), .ZN(n10013) );
  NAND2_X1 U9696 ( .A1(n10188), .A2(n9470), .ZN(n9728) );
  OAI21_X1 U9697 ( .B1(n10014), .B2(n10013), .A(n9728), .ZN(n10000) );
  NAND2_X1 U9698 ( .A1(n9998), .A2(n10015), .ZN(n9733) );
  NAND2_X1 U9699 ( .A1(n10184), .A2(n9508), .ZN(n9732) );
  NAND2_X1 U9700 ( .A1(n10000), .A2(n10001), .ZN(n9999) );
  NAND2_X1 U9701 ( .A1(n9999), .A2(n9732), .ZN(n9981) );
  INV_X1 U9702 ( .A(n9655), .ZN(n8449) );
  AOI21_X2 U9703 ( .B1(n9981), .B2(n9980), .A(n8449), .ZN(n9971) );
  NAND2_X1 U9704 ( .A1(n10175), .A2(n8450), .ZN(n9653) );
  INV_X1 U9705 ( .A(n9653), .ZN(n8451) );
  OR2_X1 U9706 ( .A1(n10168), .A2(n9973), .ZN(n9651) );
  NAND2_X1 U9707 ( .A1(n10168), .A2(n9973), .ZN(n9652) );
  NAND2_X1 U9708 ( .A1(n9651), .A2(n9652), .ZN(n9951) );
  NAND2_X1 U9709 ( .A1(n10163), .A2(n9547), .ZN(n9650) );
  INV_X1 U9710 ( .A(n9649), .ZN(n8452) );
  NOR2_X1 U9711 ( .A1(n9935), .A2(n8452), .ZN(n9911) );
  OR2_X1 U9712 ( .A1(n10158), .A2(n9934), .ZN(n9577) );
  NAND2_X1 U9713 ( .A1(n10158), .A2(n9934), .ZN(n9751) );
  NAND2_X1 U9714 ( .A1(n9911), .A2(n9919), .ZN(n9910) );
  NAND2_X1 U9715 ( .A1(n9910), .A2(n9751), .ZN(n8457) );
  OR2_X1 U9716 ( .A1(n10268), .A2(n8453), .ZN(n8455) );
  NAND2_X1 U9717 ( .A1(n9574), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8454) );
  NAND2_X1 U9718 ( .A1(n8487), .A2(n9912), .ZN(n9754) );
  INV_X1 U9719 ( .A(n9912), .ZN(n8456) );
  NAND2_X1 U9720 ( .A1(n10152), .A2(n8456), .ZN(n9756) );
  XNOR2_X1 U9721 ( .A(n8457), .B(n5400), .ZN(n8468) );
  NAND2_X1 U9722 ( .A1(n9840), .A2(n10131), .ZN(n8466) );
  INV_X1 U9723 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8461) );
  NAND2_X1 U9724 ( .A1(n5768), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8460) );
  NAND2_X1 U9725 ( .A1(n8458), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8459) );
  OAI211_X1 U9726 ( .C1(n8462), .C2(n8461), .A(n8460), .B(n8459), .ZN(n9839)
         );
  INV_X1 U9727 ( .A(P1_B_REG_SCAN_IN), .ZN(n9831) );
  NOR2_X1 U9728 ( .A1(n8463), .A2(n9831), .ZN(n8464) );
  NOR2_X1 U9729 ( .A1(n10083), .A2(n8464), .ZN(n9901) );
  NAND2_X1 U9730 ( .A1(n9839), .A2(n9901), .ZN(n8465) );
  AOI21_X2 U9731 ( .B1(n8468), .B2(n10125), .A(n8467), .ZN(n10154) );
  NAND2_X1 U9732 ( .A1(n9567), .A2(n10132), .ZN(n8469) );
  AND2_X1 U9733 ( .A1(n10223), .A2(n10109), .ZN(n8471) );
  OR2_X1 U9734 ( .A1(n10216), .A2(n10129), .ZN(n8472) );
  NAND2_X1 U9735 ( .A1(n10039), .A2(n10059), .ZN(n8474) );
  INV_X1 U9736 ( .A(n10084), .ZN(n10040) );
  NAND2_X1 U9737 ( .A1(n10012), .A2(n9470), .ZN(n8476) );
  NAND2_X1 U9738 ( .A1(n8477), .A2(n8476), .ZN(n9992) );
  NAND2_X1 U9739 ( .A1(n9992), .A2(n5652), .ZN(n8479) );
  NOR2_X1 U9740 ( .A1(n10168), .A2(n9940), .ZN(n8480) );
  INV_X1 U9741 ( .A(n8482), .ZN(n10156) );
  OAI22_X1 U9742 ( .A1(n10093), .A2(n8484), .B1(n8483), .B2(n10090), .ZN(n8485) );
  AOI21_X1 U9743 ( .B1(n10152), .B2(n10095), .A(n8485), .ZN(n8490) );
  INV_X1 U9744 ( .A(n10158), .ZN(n9920) );
  INV_X1 U9745 ( .A(n10175), .ZN(n9964) );
  OR2_X2 U9746 ( .A1(n10137), .A2(n10223), .ZN(n10135) );
  INV_X1 U9747 ( .A(n10203), .ZN(n10064) );
  NOR2_X1 U9748 ( .A1(n10188), .A2(n10027), .ZN(n10009) );
  NAND2_X1 U9749 ( .A1(n9998), .A2(n10009), .ZN(n9993) );
  INV_X1 U9750 ( .A(n9921), .ZN(n8486) );
  NAND2_X1 U9751 ( .A1(n8487), .A2(n8486), .ZN(n9906) );
  AOI21_X1 U9752 ( .B1(n10152), .B2(n9921), .A(n11009), .ZN(n8488) );
  AND2_X1 U9753 ( .A1(n9906), .A2(n8488), .ZN(n10151) );
  NAND2_X1 U9754 ( .A1(n10151), .A2(n10138), .ZN(n8489) );
  OAI211_X1 U9755 ( .C1(n10156), .C2(n10148), .A(n8490), .B(n8489), .ZN(n8491)
         );
  INV_X1 U9756 ( .A(n8491), .ZN(n8492) );
  OAI21_X1 U9757 ( .B1(n10154), .B2(n10141), .A(n8492), .ZN(P1_U3355) );
  INV_X1 U9758 ( .A(n10661), .ZN(n8493) );
  OAI222_X1 U9759 ( .A1(n5036), .A2(n8495), .B1(n8494), .B2(n8493), .C1(
        P2_U3152), .C2(n8811), .ZN(P2_U3339) );
  INV_X1 U9760 ( .A(n8497), .ZN(n8499) );
  NAND2_X1 U9761 ( .A1(n8499), .A2(n8498), .ZN(n8500) );
  NAND2_X1 U9762 ( .A1(n8501), .A2(n8500), .ZN(n8506) );
  MUX2_X1 U9763 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n5668), .Z(n8502) );
  NAND2_X1 U9764 ( .A1(n8502), .A2(SI_30_), .ZN(n8608) );
  INV_X1 U9765 ( .A(n8502), .ZN(n8503) );
  NAND2_X1 U9766 ( .A1(n8503), .A2(n5272), .ZN(n8504) );
  AND2_X1 U9767 ( .A1(n8608), .A2(n8504), .ZN(n8505) );
  NAND2_X1 U9768 ( .A1(n8506), .A2(n8505), .ZN(n8609) );
  INV_X1 U9769 ( .A(n9573), .ZN(n8826) );
  INV_X1 U9770 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10549) );
  OAI222_X1 U9771 ( .A1(P1_U3084), .A2(n8496), .B1(n10265), .B2(n8826), .C1(
        n10549), .C2(n10267), .ZN(P1_U3323) );
  XNOR2_X1 U9772 ( .A(n9369), .B(n8563), .ZN(n8511) );
  OR2_X1 U9773 ( .A1(n9271), .A2(n8562), .ZN(n8512) );
  NAND2_X1 U9774 ( .A1(n8511), .A2(n8512), .ZN(n8940) );
  INV_X1 U9775 ( .A(n8940), .ZN(n8510) );
  OR2_X1 U9776 ( .A1(n8942), .A2(n8510), .ZN(n8849) );
  XNOR2_X1 U9777 ( .A(n9361), .B(n8563), .ZN(n8902) );
  NAND2_X1 U9778 ( .A1(n9252), .A2(n8535), .ZN(n8508) );
  NOR2_X1 U9779 ( .A1(n8902), .A2(n8508), .ZN(n8517) );
  AOI21_X1 U9780 ( .B1(n8902), .B2(n8508), .A(n8517), .ZN(n8853) );
  INV_X1 U9781 ( .A(n8853), .ZN(n8516) );
  OR2_X1 U9782 ( .A1(n8849), .A2(n8516), .ZN(n8509) );
  OR2_X1 U9783 ( .A1(n8510), .A2(n8944), .ZN(n8515) );
  INV_X1 U9784 ( .A(n8511), .ZN(n8514) );
  INV_X1 U9785 ( .A(n8512), .ZN(n8513) );
  NAND2_X1 U9786 ( .A1(n8514), .A2(n8513), .ZN(n8941) );
  AND2_X1 U9787 ( .A1(n8515), .A2(n8941), .ZN(n8850) );
  INV_X1 U9788 ( .A(n8517), .ZN(n8518) );
  NAND2_X1 U9789 ( .A1(n8901), .A2(n8518), .ZN(n8523) );
  XNOR2_X1 U9790 ( .A(n9357), .B(n8551), .ZN(n8519) );
  NOR2_X1 U9791 ( .A1(n9233), .A2(n8562), .ZN(n8520) );
  NAND2_X1 U9792 ( .A1(n8519), .A2(n8520), .ZN(n8524) );
  INV_X1 U9793 ( .A(n8519), .ZN(n8860) );
  INV_X1 U9794 ( .A(n8520), .ZN(n8521) );
  NAND2_X1 U9795 ( .A1(n8860), .A2(n8521), .ZN(n8522) );
  AND2_X1 U9796 ( .A1(n8524), .A2(n8522), .ZN(n8899) );
  NAND2_X1 U9797 ( .A1(n8523), .A2(n8899), .ZN(n8858) );
  NAND2_X1 U9798 ( .A1(n8858), .A2(n8524), .ZN(n8529) );
  XNOR2_X1 U9799 ( .A(n9352), .B(n8551), .ZN(n8525) );
  NOR2_X1 U9800 ( .A1(n9213), .A2(n8562), .ZN(n8526) );
  NAND2_X1 U9801 ( .A1(n8525), .A2(n8526), .ZN(n8531) );
  INV_X1 U9802 ( .A(n8525), .ZN(n8910) );
  INV_X1 U9803 ( .A(n8526), .ZN(n8527) );
  NAND2_X1 U9804 ( .A1(n8910), .A2(n8527), .ZN(n8528) );
  AND2_X1 U9805 ( .A1(n8531), .A2(n8528), .ZN(n8859) );
  NOR2_X1 U9806 ( .A1(n8530), .A2(n8562), .ZN(n8533) );
  XNOR2_X1 U9807 ( .A(n9347), .B(n8551), .ZN(n8534) );
  XOR2_X1 U9808 ( .A(n8533), .B(n8534), .Z(n8914) );
  XNOR2_X1 U9809 ( .A(n9175), .B(n8563), .ZN(n8536) );
  NAND2_X1 U9810 ( .A1(n9155), .A2(n8535), .ZN(n8841) );
  INV_X1 U9811 ( .A(n8536), .ZN(n8537) );
  AND2_X1 U9812 ( .A1(n8538), .A2(n8537), .ZN(n8539) );
  XNOR2_X1 U9813 ( .A(n9162), .B(n8551), .ZN(n8542) );
  XNOR2_X1 U9814 ( .A(n8543), .B(n8542), .ZN(n8891) );
  INV_X1 U9815 ( .A(n8891), .ZN(n8541) );
  NOR2_X1 U9816 ( .A1(n8890), .A2(n8562), .ZN(n8540) );
  NAND2_X1 U9817 ( .A1(n8543), .A2(n8542), .ZN(n8544) );
  XNOR2_X1 U9818 ( .A(n9330), .B(n8551), .ZN(n8545) );
  NOR2_X1 U9819 ( .A1(n9158), .A2(n8562), .ZN(n8546) );
  XNOR2_X1 U9820 ( .A(n8545), .B(n8546), .ZN(n8870) );
  INV_X1 U9821 ( .A(n8545), .ZN(n8548) );
  INV_X1 U9822 ( .A(n8546), .ZN(n8547) );
  NAND2_X1 U9823 ( .A1(n8548), .A2(n8547), .ZN(n8549) );
  XNOR2_X1 U9824 ( .A(n9133), .B(n8551), .ZN(n8828) );
  NOR2_X1 U9825 ( .A1(n8871), .A2(n8562), .ZN(n8550) );
  NAND2_X1 U9826 ( .A1(n8828), .A2(n8550), .ZN(n8558) );
  OAI21_X1 U9827 ( .B1(n8828), .B2(n8550), .A(n8558), .ZN(n8954) );
  XNOR2_X1 U9828 ( .A(n9321), .B(n8551), .ZN(n8552) );
  NOR2_X1 U9829 ( .A1(n9122), .A2(n8562), .ZN(n8553) );
  NAND2_X1 U9830 ( .A1(n8552), .A2(n8553), .ZN(n8561) );
  INV_X1 U9831 ( .A(n8552), .ZN(n8555) );
  INV_X1 U9832 ( .A(n8553), .ZN(n8554) );
  NAND2_X1 U9833 ( .A1(n8555), .A2(n8554), .ZN(n8556) );
  NAND2_X1 U9834 ( .A1(n8561), .A2(n8556), .ZN(n8827) );
  OR2_X1 U9835 ( .A1(n8954), .A2(n8827), .ZN(n8557) );
  OR2_X1 U9836 ( .A1(n8827), .A2(n8558), .ZN(n8559) );
  NAND2_X1 U9837 ( .A1(n8830), .A2(n8561), .ZN(n8572) );
  NOR2_X1 U9838 ( .A1(n8833), .A2(n8562), .ZN(n8564) );
  MUX2_X1 U9839 ( .A(n8833), .B(n8564), .S(n8563), .Z(n8567) );
  INV_X1 U9840 ( .A(n9316), .ZN(n8584) );
  NOR3_X1 U9841 ( .A1(n8584), .A2(n8567), .A3(n8975), .ZN(n8565) );
  AOI21_X1 U9842 ( .B1(n8567), .B2(n8584), .A(n8565), .ZN(n8571) );
  NAND3_X1 U9843 ( .A1(n9316), .A2(n8567), .A3(n8963), .ZN(n8566) );
  OAI21_X1 U9844 ( .B1(n9316), .B2(n8567), .A(n8566), .ZN(n8568) );
  NAND2_X1 U9845 ( .A1(n8572), .A2(n8568), .ZN(n8570) );
  OAI21_X1 U9846 ( .B1(n8584), .B2(n8963), .A(n8953), .ZN(n8569) );
  OAI211_X1 U9847 ( .C1(n8572), .C2(n8571), .A(n8570), .B(n8569), .ZN(n8577)
         );
  NOR2_X1 U9848 ( .A1(n8573), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8575) );
  OAI22_X1 U9849 ( .A1(n8588), .A2(n8964), .B1(n9122), .B2(n8930), .ZN(n8574)
         );
  AOI211_X1 U9850 ( .C1(n8582), .C2(n8935), .A(n8575), .B(n8574), .ZN(n8576)
         );
  NAND2_X1 U9851 ( .A1(n8577), .A2(n8576), .ZN(P2_U3222) );
  XOR2_X1 U9852 ( .A(n8793), .B(n8578), .Z(n9320) );
  INV_X1 U9853 ( .A(n8579), .ZN(n8580) );
  AOI21_X1 U9854 ( .B1(n9316), .B2(n8581), .A(n8580), .ZN(n9317) );
  AOI22_X1 U9855 ( .A1(n8582), .A2(n9202), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9303), .ZN(n8583) );
  OAI21_X1 U9856 ( .B1(n8584), .B2(n10819), .A(n8583), .ZN(n8593) );
  INV_X1 U9857 ( .A(n8585), .ZN(n8587) );
  INV_X1 U9858 ( .A(n8793), .ZN(n8586) );
  AOI21_X1 U9859 ( .B1(n8587), .B2(n8586), .A(n9264), .ZN(n8591) );
  OAI22_X1 U9860 ( .A1(n8588), .A2(n9270), .B1(n9122), .B2(n9272), .ZN(n8589)
         );
  AOI21_X1 U9861 ( .B1(n8591), .B2(n8590), .A(n8589), .ZN(n9319) );
  NOR2_X1 U9862 ( .A1(n9319), .A2(n9303), .ZN(n8592) );
  AOI211_X1 U9863 ( .C1(n9226), .C2(n9317), .A(n8593), .B(n8592), .ZN(n8594)
         );
  OAI21_X1 U9864 ( .B1(n9320), .B2(n9300), .A(n8594), .ZN(P2_U3268) );
  OAI21_X1 U9865 ( .B1(n8930), .B2(n8596), .A(n8595), .ZN(n8597) );
  AOI21_X1 U9866 ( .B1(n8960), .B2(n8986), .A(n8597), .ZN(n8598) );
  OAI21_X1 U9867 ( .B1(n8599), .B2(n8968), .A(n8598), .ZN(n8605) );
  AOI22_X1 U9868 ( .A1(n8600), .A2(n8915), .B1(n8840), .B2(n8988), .ZN(n8602)
         );
  NOR3_X1 U9869 ( .A1(n8603), .A2(n8602), .A3(n8601), .ZN(n8604) );
  AOI211_X1 U9870 ( .C1(n9389), .C2(n8975), .A(n8605), .B(n8604), .ZN(n8606)
         );
  OAI21_X1 U9871 ( .B1(n8607), .B2(n8953), .A(n8606), .ZN(P2_U3217) );
  MUX2_X1 U9872 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n5663), .Z(n8610) );
  XNOR2_X1 U9873 ( .A(n8610), .B(SI_31_), .ZN(n8611) );
  NAND2_X1 U9874 ( .A1(n10260), .A2(n8616), .ZN(n8614) );
  INV_X1 U9875 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9417) );
  OR2_X1 U9876 ( .A1(n5039), .A2(n9417), .ZN(n8613) );
  NAND2_X2 U9877 ( .A1(n8614), .A2(n8613), .ZN(n9304) );
  INV_X1 U9878 ( .A(n9094), .ZN(n8619) );
  OR2_X1 U9879 ( .A1(n9304), .A2(n8619), .ZN(n8618) );
  INV_X1 U9880 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8825) );
  NOR2_X1 U9881 ( .A1(n5038), .A2(n8825), .ZN(n8615) );
  INV_X1 U9882 ( .A(n9098), .ZN(n9307) );
  INV_X1 U9883 ( .A(n8977), .ZN(n8617) );
  NAND2_X1 U9884 ( .A1(n9307), .A2(n8617), .ZN(n8755) );
  NAND2_X1 U9885 ( .A1(n9304), .A2(n8619), .ZN(n8810) );
  AND2_X1 U9886 ( .A1(n9098), .A2(n8977), .ZN(n8808) );
  INV_X1 U9887 ( .A(n8808), .ZN(n8756) );
  AND2_X1 U9888 ( .A1(n8620), .A2(n8796), .ZN(n8621) );
  MUX2_X1 U9889 ( .A(n8809), .B(n5096), .S(n8752), .Z(n8759) );
  INV_X1 U9890 ( .A(n8752), .ZN(n8760) );
  AND2_X1 U9891 ( .A1(n8730), .A2(n8622), .ZN(n8729) );
  NAND2_X1 U9892 ( .A1(n8623), .A2(n10815), .ZN(n8767) );
  NAND2_X1 U9893 ( .A1(n10815), .A2(n8796), .ZN(n8626) );
  INV_X1 U9894 ( .A(n8624), .ZN(n8625) );
  AOI21_X1 U9895 ( .B1(n8627), .B2(n8626), .A(n8625), .ZN(n8628) );
  MUX2_X1 U9896 ( .A(n8767), .B(n8628), .S(n8752), .Z(n8630) );
  OAI21_X1 U9897 ( .B1(n8630), .B2(n7209), .A(n8629), .ZN(n8637) );
  AND2_X1 U9898 ( .A1(n8998), .A2(n10864), .ZN(n8631) );
  MUX2_X1 U9899 ( .A(n8632), .B(n8631), .S(n8752), .Z(n8636) );
  MUX2_X1 U9900 ( .A(n8634), .B(n8633), .S(n8752), .Z(n8635) );
  OAI211_X1 U9901 ( .C1(n8637), .C2(n8636), .A(n8768), .B(n8635), .ZN(n8643)
         );
  NAND2_X1 U9902 ( .A1(n8996), .A2(n8638), .ZN(n8639) );
  MUX2_X1 U9903 ( .A(n8640), .B(n8639), .S(n8752), .Z(n8641) );
  NAND3_X1 U9904 ( .A1(n8643), .A2(n8642), .A3(n8641), .ZN(n8647) );
  MUX2_X1 U9905 ( .A(n8645), .B(n8644), .S(n8752), .Z(n8646) );
  NAND2_X1 U9906 ( .A1(n8647), .A2(n8646), .ZN(n8653) );
  MUX2_X1 U9907 ( .A(n8994), .B(n8648), .S(n8752), .Z(n8649) );
  OAI21_X1 U9908 ( .B1(n8653), .B2(n8650), .A(n8649), .ZN(n8655) );
  INV_X1 U9909 ( .A(n8651), .ZN(n8652) );
  NAND2_X1 U9910 ( .A1(n8653), .A2(n8652), .ZN(n8654) );
  NAND2_X1 U9911 ( .A1(n8993), .A2(n8760), .ZN(n8659) );
  NAND2_X1 U9912 ( .A1(n8656), .A2(n8752), .ZN(n8658) );
  MUX2_X1 U9913 ( .A(n8659), .B(n8658), .S(n8657), .Z(n8660) );
  INV_X1 U9914 ( .A(n8667), .ZN(n8666) );
  NAND2_X1 U9915 ( .A1(n8672), .A2(n8661), .ZN(n8664) );
  INV_X1 U9916 ( .A(n8662), .ZN(n8663) );
  MUX2_X1 U9917 ( .A(n8664), .B(n8663), .S(n8752), .Z(n8665) );
  NAND3_X1 U9918 ( .A1(n8671), .A2(n8670), .A3(n8669), .ZN(n8677) );
  NAND3_X1 U9919 ( .A1(n8673), .A2(n8777), .A3(n8672), .ZN(n8675) );
  NAND2_X1 U9920 ( .A1(n8675), .A2(n8674), .ZN(n8676) );
  INV_X1 U9921 ( .A(n8781), .ZN(n8683) );
  INV_X1 U9922 ( .A(n8678), .ZN(n8780) );
  NAND2_X1 U9923 ( .A1(n8780), .A2(n8679), .ZN(n8681) );
  MUX2_X1 U9924 ( .A(n8681), .B(n8680), .S(n8760), .Z(n8682) );
  MUX2_X1 U9925 ( .A(n8686), .B(n8685), .S(n8760), .Z(n8687) );
  MUX2_X1 U9926 ( .A(n8689), .B(n8688), .S(n8752), .Z(n8690) );
  INV_X1 U9927 ( .A(n8691), .ZN(n8693) );
  MUX2_X1 U9928 ( .A(n8693), .B(n8360), .S(n8752), .Z(n8694) );
  NOR2_X1 U9929 ( .A1(n8211), .A2(n8694), .ZN(n8695) );
  NAND2_X1 U9930 ( .A1(n8696), .A2(n8695), .ZN(n8700) );
  MUX2_X1 U9931 ( .A(n8698), .B(n8697), .S(n8752), .Z(n8699) );
  NAND3_X1 U9932 ( .A1(n8700), .A2(n8764), .A3(n8699), .ZN(n8704) );
  NAND2_X1 U9933 ( .A1(n9375), .A2(n8760), .ZN(n8702) );
  OR2_X1 U9934 ( .A1(n9375), .A2(n8760), .ZN(n8701) );
  MUX2_X1 U9935 ( .A(n8702), .B(n8701), .S(n9253), .Z(n8703) );
  NAND3_X1 U9936 ( .A1(n8704), .A2(n9249), .A3(n8703), .ZN(n8708) );
  MUX2_X1 U9937 ( .A(n8706), .B(n8705), .S(n8752), .Z(n8707) );
  NAND3_X1 U9938 ( .A1(n8708), .A2(n9229), .A3(n8707), .ZN(n8718) );
  AND2_X1 U9939 ( .A1(n9252), .A2(n8752), .ZN(n8710) );
  NOR2_X1 U9940 ( .A1(n9252), .A2(n8752), .ZN(n8709) );
  MUX2_X1 U9941 ( .A(n8710), .B(n8709), .S(n9361), .Z(n8711) );
  NOR2_X1 U9942 ( .A1(n9215), .A2(n8711), .ZN(n8717) );
  INV_X1 U9943 ( .A(n8712), .ZN(n8715) );
  INV_X1 U9944 ( .A(n8713), .ZN(n8714) );
  MUX2_X1 U9945 ( .A(n8715), .B(n8714), .S(n8760), .Z(n8716) );
  AOI21_X1 U9946 ( .B1(n8718), .B2(n8717), .A(n8716), .ZN(n8720) );
  INV_X1 U9947 ( .A(n9207), .ZN(n9194) );
  AOI21_X1 U9948 ( .B1(n8722), .B2(n5061), .A(n8752), .ZN(n8721) );
  INV_X1 U9949 ( .A(n8723), .ZN(n8724) );
  AND2_X1 U9950 ( .A1(n8734), .A2(n8725), .ZN(n8727) );
  NAND2_X1 U9951 ( .A1(n8725), .A2(n8724), .ZN(n8726) );
  MUX2_X1 U9952 ( .A(n8727), .B(n8726), .S(n8752), .Z(n8728) );
  NAND3_X1 U9953 ( .A1(n8735), .A2(n8732), .A3(n8730), .ZN(n8731) );
  AOI21_X1 U9954 ( .B1(n8731), .B2(n8736), .A(n8737), .ZN(n8741) );
  INV_X1 U9955 ( .A(n8732), .ZN(n8733) );
  AOI21_X1 U9956 ( .B1(n8735), .B2(n8734), .A(n8733), .ZN(n8739) );
  INV_X1 U9957 ( .A(n8736), .ZN(n8738) );
  INV_X1 U9958 ( .A(n8737), .ZN(n9108) );
  OAI21_X1 U9959 ( .B1(n8739), .B2(n8738), .A(n9108), .ZN(n8740) );
  INV_X1 U9960 ( .A(n8744), .ZN(n8745) );
  NAND2_X1 U9961 ( .A1(n8746), .A2(n8745), .ZN(n8747) );
  MUX2_X1 U9962 ( .A(n8748), .B(n8747), .S(n8760), .Z(n8751) );
  INV_X1 U9963 ( .A(n8749), .ZN(n8750) );
  MUX2_X1 U9964 ( .A(n8804), .B(n8806), .S(n8752), .Z(n8753) );
  OAI21_X1 U9965 ( .B1(n8754), .B2(n8795), .A(n8753), .ZN(n8757) );
  NAND3_X1 U9966 ( .A1(n8757), .A2(n8756), .A3(n8755), .ZN(n8758) );
  MUX2_X1 U9967 ( .A(n9094), .B(n9304), .S(n8760), .Z(n8762) );
  NAND2_X1 U9968 ( .A1(n9304), .A2(n9094), .ZN(n8761) );
  NAND2_X1 U9969 ( .A1(n8762), .A2(n8761), .ZN(n8763) );
  INV_X1 U9970 ( .A(n8764), .ZN(n9267) );
  NOR4_X1 U9971 ( .A1(n8767), .A2(n8801), .A3(n8766), .A4(n8765), .ZN(n8771)
         );
  NAND4_X1 U9972 ( .A1(n8771), .A2(n8770), .A3(n8769), .A4(n8768), .ZN(n8776)
         );
  INV_X1 U9973 ( .A(n8772), .ZN(n8774) );
  NOR4_X1 U9974 ( .A1(n8776), .A2(n8775), .A3(n8774), .A4(n8773), .ZN(n8778)
         );
  NAND2_X1 U9975 ( .A1(n8778), .A2(n8777), .ZN(n8782) );
  NOR4_X1 U9976 ( .A1(n8782), .A2(n8781), .A3(n8780), .A4(n8779), .ZN(n8783)
         );
  NAND4_X1 U9977 ( .A1(n9283), .A2(n8785), .A3(n8784), .A4(n8783), .ZN(n8786)
         );
  NOR4_X1 U9978 ( .A1(n5465), .A2(n5469), .A3(n9267), .A4(n8786), .ZN(n8787)
         );
  NAND4_X1 U9979 ( .A1(n8789), .A2(n9207), .A3(n8788), .A4(n8787), .ZN(n8790)
         );
  NOR4_X1 U9980 ( .A1(n9142), .A2(n9152), .A3(n8791), .A4(n8790), .ZN(n8792)
         );
  NAND4_X1 U9981 ( .A1(n8793), .A2(n5540), .A3(n9119), .A4(n8792), .ZN(n8794)
         );
  NOR2_X1 U9982 ( .A1(n8800), .A2(n10830), .ZN(n8799) );
  XNOR2_X1 U9983 ( .A(n8814), .B(n8811), .ZN(n8813) );
  NAND2_X1 U9984 ( .A1(n8815), .A2(n5651), .ZN(n8816) );
  NOR2_X1 U9985 ( .A1(n8817), .A2(n8816), .ZN(n8824) );
  NOR3_X1 U9986 ( .A1(n10787), .A2(n8819), .A3(n8818), .ZN(n8822) );
  OAI21_X1 U9987 ( .B1(n8823), .B2(n8820), .A(P2_B_REG_SCAN_IN), .ZN(n8821) );
  OAI22_X1 U9988 ( .A1(n8824), .A2(n8823), .B1(n8822), .B2(n8821), .ZN(
        P2_U3244) );
  OAI222_X1 U9989 ( .A1(n8494), .A2(n8826), .B1(n6520), .B2(P2_U3152), .C1(
        n8825), .C2(n5036), .ZN(P2_U3328) );
  AOI21_X1 U9990 ( .B1(n8956), .B2(n8827), .A(n8953), .ZN(n8832) );
  INV_X1 U9991 ( .A(n8828), .ZN(n8829) );
  NOR3_X1 U9992 ( .A1(n8829), .A2(n8871), .A3(n8922), .ZN(n8831) );
  OAI21_X1 U9993 ( .B1(n8832), .B2(n8831), .A(n8830), .ZN(n8839) );
  OR2_X1 U9994 ( .A1(n8833), .A2(n9270), .ZN(n8835) );
  NAND2_X1 U9995 ( .A1(n8981), .A2(n9254), .ZN(n8834) );
  NAND2_X1 U9996 ( .A1(n8835), .A2(n8834), .ZN(n9112) );
  OAI22_X1 U9997 ( .A1(n9103), .A2(n8968), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10520), .ZN(n8837) );
  NOR2_X1 U9998 ( .A1(n9106), .A2(n8963), .ZN(n8836) );
  AOI211_X1 U9999 ( .C1(n8882), .C2(n9112), .A(n8837), .B(n8836), .ZN(n8838)
         );
  NAND2_X1 U10000 ( .A1(n8839), .A2(n8838), .ZN(P2_U3216) );
  NAND2_X1 U10001 ( .A1(n8840), .A2(n9155), .ZN(n8844) );
  NAND2_X1 U10002 ( .A1(n8841), .A2(n8915), .ZN(n8843) );
  MUX2_X1 U10003 ( .A(n8844), .B(n8843), .S(n8842), .Z(n8848) );
  AOI22_X1 U10004 ( .A1(n9197), .A2(n8966), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8845) );
  OAI21_X1 U10005 ( .B1(n8890), .B2(n8964), .A(n8845), .ZN(n8846) );
  AOI21_X1 U10006 ( .B1(n9173), .B2(n8935), .A(n8846), .ZN(n8847) );
  OAI211_X1 U10007 ( .C1(n9175), .C2(n8963), .A(n8848), .B(n8847), .ZN(
        P2_U3218) );
  OR2_X1 U10008 ( .A1(n8943), .A2(n8849), .ZN(n8851) );
  NAND2_X1 U10009 ( .A1(n8851), .A2(n8850), .ZN(n8852) );
  OAI211_X1 U10010 ( .C1(n8853), .C2(n8852), .A(n8901), .B(n8915), .ZN(n8857)
         );
  NAND2_X1 U10011 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9087) );
  OAI21_X1 U10012 ( .B1(n8964), .B2(n9233), .A(n9087), .ZN(n8855) );
  NOR2_X1 U10013 ( .A1(n8968), .A2(n9239), .ZN(n8854) );
  AOI211_X1 U10014 ( .C1(n8966), .C2(n8984), .A(n8855), .B(n8854), .ZN(n8856)
         );
  OAI211_X1 U10015 ( .C1(n9236), .C2(n8963), .A(n8857), .B(n8856), .ZN(
        P2_U3221) );
  AOI21_X1 U10016 ( .B1(n8858), .B2(n5417), .A(n8953), .ZN(n8862) );
  NOR3_X1 U10017 ( .A1(n8860), .A2(n9233), .A3(n8922), .ZN(n8861) );
  OAI21_X1 U10018 ( .B1(n8862), .B2(n8861), .A(n8913), .ZN(n8866) );
  AOI22_X1 U10019 ( .A1(n9197), .A2(n8960), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8863) );
  OAI21_X1 U10020 ( .B1(n9233), .B2(n8930), .A(n8863), .ZN(n8864) );
  AOI21_X1 U10021 ( .B1(n9203), .B2(n8935), .A(n8864), .ZN(n8865) );
  OAI211_X1 U10022 ( .C1(n9205), .C2(n8963), .A(n8866), .B(n8865), .ZN(
        P2_U3225) );
  INV_X1 U10023 ( .A(n8867), .ZN(n8868) );
  AOI21_X1 U10024 ( .B1(n8870), .B2(n8869), .A(n8868), .ZN(n8876) );
  OAI22_X1 U10025 ( .A1(n8871), .A2(n9270), .B1(n8890), .B2(n9272), .ZN(n9144)
         );
  INV_X1 U10026 ( .A(n9138), .ZN(n8872) );
  OAI22_X1 U10027 ( .A1(n8872), .A2(n8968), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10461), .ZN(n8874) );
  NOR2_X1 U10028 ( .A1(n9140), .A2(n8963), .ZN(n8873) );
  AOI211_X1 U10029 ( .C1(n8882), .C2(n9144), .A(n8874), .B(n8873), .ZN(n8875)
         );
  OAI21_X1 U10030 ( .B1(n8876), .B2(n8953), .A(n8875), .ZN(P2_U3227) );
  INV_X1 U10031 ( .A(n8877), .ZN(n8970) );
  NOR2_X1 U10032 ( .A1(n8922), .A2(n8881), .ZN(n8879) );
  AOI22_X1 U10033 ( .A1(n8970), .A2(n8915), .B1(n8879), .B2(n8878), .ZN(n8889)
         );
  NAND2_X1 U10034 ( .A1(n9253), .A2(n10821), .ZN(n8880) );
  OAI21_X1 U10035 ( .B1(n8881), .B2(n9272), .A(n8880), .ZN(n9285) );
  AOI22_X1 U10036 ( .A1(n9285), .A2(n8882), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3152), .ZN(n8883) );
  OAI21_X1 U10037 ( .B1(n9289), .B2(n8968), .A(n8883), .ZN(n8886) );
  NOR2_X1 U10038 ( .A1(n8884), .A2(n8953), .ZN(n8885) );
  AOI211_X1 U10039 ( .C1(n9379), .C2(n8975), .A(n8886), .B(n8885), .ZN(n8887)
         );
  OAI21_X1 U10040 ( .B1(n8889), .B2(n8888), .A(n8887), .ZN(P2_U3228) );
  OAI22_X1 U10041 ( .A1(n8891), .A2(n8953), .B1(n8890), .B2(n8922), .ZN(n8893)
         );
  NAND2_X1 U10042 ( .A1(n8893), .A2(n8892), .ZN(n8898) );
  INV_X1 U10043 ( .A(n8894), .ZN(n9161) );
  INV_X1 U10044 ( .A(n9158), .ZN(n8982) );
  AOI22_X1 U10045 ( .A1(n8982), .A2(n8960), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n8895) );
  OAI21_X1 U10046 ( .B1(n9187), .B2(n8930), .A(n8895), .ZN(n8896) );
  AOI21_X1 U10047 ( .B1(n9161), .B2(n8935), .A(n8896), .ZN(n8897) );
  OAI211_X1 U10048 ( .C1(n9334), .C2(n8963), .A(n8898), .B(n8897), .ZN(
        P2_U3231) );
  INV_X1 U10049 ( .A(n8899), .ZN(n8900) );
  AOI21_X1 U10050 ( .B1(n8901), .B2(n8900), .A(n8953), .ZN(n8904) );
  NOR3_X1 U10051 ( .A1(n8902), .A2(n9212), .A3(n8922), .ZN(n8903) );
  OAI21_X1 U10052 ( .B1(n8904), .B2(n8903), .A(n8858), .ZN(n8909) );
  INV_X1 U10053 ( .A(n9222), .ZN(n8907) );
  INV_X1 U10054 ( .A(n9213), .ZN(n8983) );
  AOI22_X1 U10055 ( .A1(n8983), .A2(n8960), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8905) );
  OAI21_X1 U10056 ( .B1(n9212), .B2(n8930), .A(n8905), .ZN(n8906) );
  AOI21_X1 U10057 ( .B1(n8907), .B2(n8935), .A(n8906), .ZN(n8908) );
  OAI211_X1 U10058 ( .C1(n9221), .C2(n8963), .A(n8909), .B(n8908), .ZN(
        P2_U3235) );
  NOR3_X1 U10059 ( .A1(n8914), .A2(n8910), .A3(n8922), .ZN(n8911) );
  NOR2_X1 U10060 ( .A1(n8911), .A2(n8966), .ZN(n8921) );
  OAI21_X1 U10061 ( .B1(n8914), .B2(n8913), .A(n8912), .ZN(n8916) );
  NAND2_X1 U10062 ( .A1(n8916), .A2(n8915), .ZN(n8920) );
  AOI22_X1 U10063 ( .A1(n9155), .A2(n8960), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8917) );
  OAI21_X1 U10064 ( .B1(n9181), .B2(n8968), .A(n8917), .ZN(n8918) );
  AOI21_X1 U10065 ( .B1(n9347), .B2(n8975), .A(n8918), .ZN(n8919) );
  OAI211_X1 U10066 ( .C1(n9213), .C2(n8921), .A(n8920), .B(n8919), .ZN(
        P2_U3237) );
  NOR3_X1 U10067 ( .A1(n8923), .A2(n8929), .A3(n8922), .ZN(n8927) );
  AOI21_X1 U10068 ( .B1(n8925), .B2(n8924), .A(n8953), .ZN(n8926) );
  OAI21_X1 U10069 ( .B1(n8927), .B2(n8926), .A(n5111), .ZN(n8939) );
  INV_X1 U10070 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10448) );
  OAI22_X1 U10071 ( .A1(n8964), .A2(n8928), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10448), .ZN(n8932) );
  NOR2_X1 U10072 ( .A1(n8930), .A2(n8929), .ZN(n8931) );
  NOR2_X1 U10073 ( .A1(n8932), .A2(n8931), .ZN(n8938) );
  NAND2_X1 U10074 ( .A1(n10970), .A2(n8975), .ZN(n8937) );
  INV_X1 U10075 ( .A(n8933), .ZN(n8934) );
  NAND2_X1 U10076 ( .A1(n8935), .A2(n8934), .ZN(n8936) );
  NAND4_X1 U10077 ( .A1(n8939), .A2(n8938), .A3(n8937), .A4(n8936), .ZN(
        P2_U3238) );
  NAND2_X1 U10078 ( .A1(n8941), .A2(n8940), .ZN(n8947) );
  OR2_X1 U10079 ( .A1(n8943), .A2(n8942), .ZN(n8945) );
  NAND2_X1 U10080 ( .A1(n8945), .A2(n8944), .ZN(n8946) );
  XOR2_X1 U10081 ( .A(n8947), .B(n8946), .Z(n8952) );
  NAND2_X1 U10082 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9063) );
  OAI21_X1 U10083 ( .B1(n8964), .B2(n9212), .A(n9063), .ZN(n8948) );
  AOI21_X1 U10084 ( .B1(n8966), .B2(n9253), .A(n8948), .ZN(n8949) );
  OAI21_X1 U10085 ( .B1(n9257), .B2(n8968), .A(n8949), .ZN(n8950) );
  AOI21_X1 U10086 ( .B1(n9369), .B2(n8975), .A(n8950), .ZN(n8951) );
  OAI21_X1 U10087 ( .B1(n8952), .B2(n8953), .A(n8951), .ZN(P2_U3240) );
  INV_X1 U10088 ( .A(n9133), .ZN(n9328) );
  AOI21_X1 U10089 ( .B1(n8955), .B2(n8954), .A(n8953), .ZN(n8957) );
  NAND2_X1 U10090 ( .A1(n8957), .A2(n8956), .ZN(n8962) );
  INV_X1 U10091 ( .A(n9122), .ZN(n8980) );
  AOI22_X1 U10092 ( .A1(n8982), .A2(n8966), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8958) );
  OAI21_X1 U10093 ( .B1(n9127), .B2(n8968), .A(n8958), .ZN(n8959) );
  AOI21_X1 U10094 ( .B1(n8960), .B2(n8980), .A(n8959), .ZN(n8961) );
  OAI211_X1 U10095 ( .C1(n9328), .C2(n8963), .A(n8962), .B(n8961), .ZN(
        P2_U3242) );
  OAI22_X1 U10096 ( .A1(n8964), .A2(n9273), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10545), .ZN(n8965) );
  AOI21_X1 U10097 ( .B1(n8966), .B2(n8987), .A(n8965), .ZN(n8967) );
  OAI21_X1 U10098 ( .B1(n8969), .B2(n8968), .A(n8967), .ZN(n8974) );
  AOI211_X1 U10099 ( .C1(n8972), .C2(n8971), .A(n8953), .B(n8970), .ZN(n8973)
         );
  AOI211_X1 U10100 ( .C1(n9383), .C2(n8975), .A(n8974), .B(n8973), .ZN(n8976)
         );
  INV_X1 U10101 ( .A(n8976), .ZN(P2_U3243) );
  MUX2_X1 U10102 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8977), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U10103 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8978), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U10104 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8979), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U10105 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8980), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10106 ( .A(n8981), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8999), .Z(
        P2_U3578) );
  MUX2_X1 U10107 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8982), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U10108 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9168), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U10109 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9197), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10110 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8983), .S(P2_U3966), .Z(
        P2_U3573) );
  INV_X1 U10111 ( .A(n9233), .ZN(n9196) );
  MUX2_X1 U10112 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9196), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10113 ( .A(n9252), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8999), .Z(
        P2_U3571) );
  MUX2_X1 U10114 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8984), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U10115 ( .A(n9253), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8999), .Z(
        P2_U3569) );
  MUX2_X1 U10116 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8985), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10117 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8986), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10118 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8987), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10119 ( .A(n8988), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8999), .Z(
        P2_U3565) );
  MUX2_X1 U10120 ( .A(n8989), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8999), .Z(
        P2_U3564) );
  MUX2_X1 U10121 ( .A(n8990), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8999), .Z(
        P2_U3563) );
  MUX2_X1 U10122 ( .A(n8991), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8999), .Z(
        P2_U3561) );
  MUX2_X1 U10123 ( .A(n8992), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8999), .Z(
        P2_U3560) );
  MUX2_X1 U10124 ( .A(n8993), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8999), .Z(
        P2_U3559) );
  MUX2_X1 U10125 ( .A(n8994), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8999), .Z(
        P2_U3558) );
  MUX2_X1 U10126 ( .A(n8995), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8999), .Z(
        P2_U3557) );
  MUX2_X1 U10127 ( .A(n8996), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8999), .Z(
        P2_U3556) );
  MUX2_X1 U10128 ( .A(n8997), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8999), .Z(
        P2_U3555) );
  MUX2_X1 U10129 ( .A(n8998), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8999), .Z(
        P2_U3554) );
  MUX2_X1 U10130 ( .A(n10820), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8999), .Z(
        P2_U3553) );
  OAI21_X1 U10131 ( .B1(n9002), .B2(n9001), .A(n9000), .ZN(n9003) );
  NAND2_X1 U10132 ( .A1(n10776), .A2(n9003), .ZN(n9012) );
  NAND2_X1 U10133 ( .A1(n10807), .A2(n9004), .ZN(n9011) );
  NOR2_X1 U10134 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10448), .ZN(n9005) );
  AOI21_X1 U10135 ( .B1(n10800), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n9005), .ZN(
        n9010) );
  OAI211_X1 U10136 ( .C1(n9008), .C2(n9007), .A(n10809), .B(n9006), .ZN(n9009)
         );
  NAND4_X1 U10137 ( .A1(n9012), .A2(n9011), .A3(n9010), .A4(n9009), .ZN(
        P2_U3256) );
  XNOR2_X1 U10138 ( .A(n9034), .B(n9026), .ZN(n9015) );
  NAND2_X1 U10139 ( .A1(n9015), .A2(n8048), .ZN(n9028) );
  OAI21_X1 U10140 ( .B1(n9015), .B2(n8048), .A(n9028), .ZN(n9016) );
  INV_X1 U10141 ( .A(n9016), .ZN(n9025) );
  NOR2_X1 U10142 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10545), .ZN(n9018) );
  NOR2_X1 U10143 ( .A1(n10792), .A2(n9027), .ZN(n9017) );
  AOI211_X1 U10144 ( .C1(n10800), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n9018), .B(
        n9017), .ZN(n9024) );
  AOI21_X1 U10145 ( .B1(n9021), .B2(n9020), .A(n9019), .ZN(n9033) );
  XNOR2_X1 U10146 ( .A(n9033), .B(n9027), .ZN(n9022) );
  NAND2_X1 U10147 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n9022), .ZN(n9035) );
  OAI211_X1 U10148 ( .C1(n9022), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10809), .B(
        n9035), .ZN(n9023) );
  OAI211_X1 U10149 ( .C1(n9025), .C2(n10801), .A(n9024), .B(n9023), .ZN(
        P2_U3260) );
  NAND2_X1 U10150 ( .A1(n9027), .A2(n9026), .ZN(n9029) );
  NAND2_X1 U10151 ( .A1(n9029), .A2(n9028), .ZN(n9032) );
  NAND2_X1 U10152 ( .A1(n9054), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9030) );
  OAI21_X1 U10153 ( .B1(n9054), .B2(P2_REG2_REG_16__SCAN_IN), .A(n9030), .ZN(
        n9031) );
  NOR2_X1 U10154 ( .A1(n9032), .A2(n9031), .ZN(n9053) );
  AOI211_X1 U10155 ( .C1(n9032), .C2(n9031), .A(n9053), .B(n10801), .ZN(n9044)
         );
  NAND2_X1 U10156 ( .A1(n9034), .A2(n9033), .ZN(n9036) );
  NAND2_X1 U10157 ( .A1(n9036), .A2(n9035), .ZN(n9038) );
  XNOR2_X1 U10158 ( .A(n9054), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n9037) );
  NOR2_X1 U10159 ( .A1(n9038), .A2(n9037), .ZN(n9045) );
  AOI21_X1 U10160 ( .B1(n9038), .B2(n9037), .A(n9045), .ZN(n9039) );
  NOR2_X1 U10161 ( .A1(n9039), .A2(n10773), .ZN(n9043) );
  NOR2_X1 U10162 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10300), .ZN(n9040) );
  AOI21_X1 U10163 ( .B1(n10800), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n9040), .ZN(
        n9041) );
  OAI21_X1 U10164 ( .B1(n10792), .B2(n9047), .A(n9041), .ZN(n9042) );
  OR3_X1 U10165 ( .A1(n9044), .A2(n9043), .A3(n9042), .ZN(P2_U3261) );
  INV_X1 U10166 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9052) );
  XNOR2_X1 U10167 ( .A(n9066), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n9049) );
  AOI21_X1 U10168 ( .B1(n9047), .B2(n9046), .A(n9045), .ZN(n9048) );
  NAND2_X1 U10169 ( .A1(n9049), .A2(n9048), .ZN(n9065) );
  OAI211_X1 U10170 ( .C1(n9049), .C2(n9048), .A(n10809), .B(n9065), .ZN(n9051)
         );
  OAI211_X1 U10171 ( .C1(n10787), .C2(n9052), .A(n9051), .B(n9050), .ZN(n9058)
         );
  AOI22_X1 U10172 ( .A1(n9061), .A2(n9277), .B1(P2_REG2_REG_17__SCAN_IN), .B2(
        n9066), .ZN(n9055) );
  NOR2_X1 U10173 ( .A1(n9056), .A2(n9055), .ZN(n9060) );
  AOI211_X1 U10174 ( .C1(n9056), .C2(n9055), .A(n9060), .B(n10801), .ZN(n9057)
         );
  AOI211_X1 U10175 ( .C1(n10807), .C2(n9061), .A(n9058), .B(n9057), .ZN(n9059)
         );
  INV_X1 U10176 ( .A(n9059), .ZN(P2_U3262) );
  NOR2_X1 U10177 ( .A1(n9073), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9083) );
  AOI21_X1 U10178 ( .B1(n9073), .B2(P2_REG2_REG_18__SCAN_IN), .A(n9083), .ZN(
        n9062) );
  XOR2_X1 U10179 ( .A(n9082), .B(n9062), .Z(n9075) );
  INV_X1 U10180 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9064) );
  OAI21_X1 U10181 ( .B1(n10787), .B2(n9064), .A(n9063), .ZN(n9072) );
  OAI21_X1 U10182 ( .B1(n9067), .B2(n9066), .A(n9065), .ZN(n9069) );
  OR2_X1 U10183 ( .A1(n9073), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9076) );
  OAI21_X1 U10184 ( .B1(n9081), .B2(n9373), .A(n9076), .ZN(n9068) );
  NOR2_X1 U10185 ( .A1(n9068), .A2(n9069), .ZN(n9078) );
  AOI21_X1 U10186 ( .B1(n9069), .B2(n9068), .A(n9078), .ZN(n9070) );
  NOR2_X1 U10187 ( .A1(n9070), .A2(n10773), .ZN(n9071) );
  AOI211_X1 U10188 ( .C1(n10807), .C2(n9073), .A(n9072), .B(n9071), .ZN(n9074)
         );
  OAI21_X1 U10189 ( .B1(n9075), .B2(n10801), .A(n9074), .ZN(P2_U3263) );
  INV_X1 U10190 ( .A(n9076), .ZN(n9077) );
  NOR2_X1 U10191 ( .A1(n9078), .A2(n9077), .ZN(n9080) );
  XNOR2_X1 U10192 ( .A(n8233), .B(n9367), .ZN(n9079) );
  XNOR2_X1 U10193 ( .A(n9080), .B(n9079), .ZN(n9091) );
  OAI22_X1 U10194 ( .A1(n9083), .A2(n9082), .B1(n8227), .B2(n9081), .ZN(n9085)
         );
  XNOR2_X1 U10195 ( .A(n8233), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n9084) );
  XNOR2_X1 U10196 ( .A(n9085), .B(n9084), .ZN(n9086) );
  AOI22_X1 U10197 ( .A1(n8233), .A2(n10807), .B1(n10776), .B2(n9086), .ZN(
        n9090) );
  INV_X1 U10198 ( .A(n9087), .ZN(n9088) );
  AOI21_X1 U10199 ( .B1(n10800), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n9088), .ZN(
        n9089) );
  OAI211_X1 U10200 ( .C1(n10773), .C2(n9091), .A(n9090), .B(n9089), .ZN(
        P2_U3264) );
  XNOR2_X1 U10201 ( .A(n9304), .B(n9092), .ZN(n9306) );
  NAND2_X1 U10202 ( .A1(n9094), .A2(n9093), .ZN(n9309) );
  NOR2_X1 U10203 ( .A1(n9303), .A2(n9309), .ZN(n9100) );
  AOI21_X1 U10204 ( .B1(n9303), .B2(P2_REG2_REG_31__SCAN_IN), .A(n9100), .ZN(
        n9096) );
  NAND2_X1 U10205 ( .A1(n9304), .A2(n9292), .ZN(n9095) );
  OAI211_X1 U10206 ( .C1(n9306), .C2(n10818), .A(n9096), .B(n9095), .ZN(
        P2_U3265) );
  XNOR2_X1 U10207 ( .A(n9098), .B(n9097), .ZN(n9310) );
  NOR2_X1 U10208 ( .A1(n9098), .A2(n10819), .ZN(n9099) );
  AOI211_X1 U10209 ( .C1(n9303), .C2(P2_REG2_REG_30__SCAN_IN), .A(n9100), .B(
        n9099), .ZN(n9101) );
  OAI21_X1 U10210 ( .B1(n10818), .B2(n9310), .A(n9101), .ZN(P2_U3266) );
  XNOR2_X1 U10211 ( .A(n9102), .B(n5540), .ZN(n9325) );
  XNOR2_X1 U10212 ( .A(n9129), .B(n9321), .ZN(n9322) );
  INV_X1 U10213 ( .A(n9103), .ZN(n9104) );
  AOI22_X1 U10214 ( .A1(n9104), .A2(n9202), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9303), .ZN(n9105) );
  OAI21_X1 U10215 ( .B1(n9106), .B2(n10819), .A(n9105), .ZN(n9115) );
  INV_X1 U10216 ( .A(n9107), .ZN(n9111) );
  AOI21_X1 U10217 ( .B1(n9109), .B2(n9108), .A(n5540), .ZN(n9110) );
  NOR3_X1 U10218 ( .A1(n9111), .A2(n9110), .A3(n9264), .ZN(n9113) );
  NOR2_X1 U10219 ( .A1(n9113), .A2(n9112), .ZN(n9324) );
  NOR2_X1 U10220 ( .A1(n9324), .A2(n9303), .ZN(n9114) );
  AOI211_X1 U10221 ( .C1(n9226), .C2(n9322), .A(n9115), .B(n9114), .ZN(n9116)
         );
  OAI21_X1 U10222 ( .B1(n9325), .B2(n9300), .A(n9116), .ZN(P2_U3269) );
  XNOR2_X1 U10223 ( .A(n9117), .B(n9119), .ZN(n9125) );
  NAND2_X1 U10224 ( .A1(n9145), .A2(n9118), .ZN(n9120) );
  XNOR2_X1 U10225 ( .A(n9120), .B(n9119), .ZN(n9121) );
  NOR2_X1 U10226 ( .A1(n9121), .A2(n9264), .ZN(n9124) );
  OAI22_X1 U10227 ( .A1(n9122), .A2(n9270), .B1(n9158), .B2(n9272), .ZN(n9123)
         );
  INV_X1 U10228 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9126) );
  OAI22_X1 U10229 ( .A1(n9127), .A2(n10823), .B1(n9126), .B2(n10829), .ZN(
        n9132) );
  INV_X1 U10230 ( .A(n9128), .ZN(n9137) );
  INV_X1 U10231 ( .A(n9129), .ZN(n9130) );
  OAI211_X1 U10232 ( .C1(n9328), .C2(n9137), .A(n9130), .B(n10881), .ZN(n9326)
         );
  NOR2_X1 U10233 ( .A1(n9326), .A2(n9280), .ZN(n9131) );
  AOI211_X1 U10234 ( .C1(n9292), .C2(n9133), .A(n9132), .B(n9131), .ZN(n9134)
         );
  OAI21_X1 U10235 ( .B1(n9327), .B2(n9303), .A(n9134), .ZN(P2_U3270) );
  XNOR2_X1 U10236 ( .A(n9135), .B(n9136), .ZN(n9333) );
  INV_X1 U10237 ( .A(n9280), .ZN(n9297) );
  AOI211_X1 U10238 ( .C1(n9330), .C2(n9159), .A(n10994), .B(n9137), .ZN(n9329)
         );
  AOI22_X1 U10239 ( .A1(n9303), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n9138), .B2(
        n9202), .ZN(n9139) );
  OAI21_X1 U10240 ( .B1(n9140), .B2(n10819), .A(n9139), .ZN(n9148) );
  INV_X1 U10241 ( .A(n9141), .ZN(n9143) );
  AOI21_X1 U10242 ( .B1(n9143), .B2(n9142), .A(n9264), .ZN(n9146) );
  AOI21_X1 U10243 ( .B1(n9146), .B2(n9145), .A(n9144), .ZN(n9332) );
  NOR2_X1 U10244 ( .A1(n9332), .A2(n9303), .ZN(n9147) );
  AOI211_X1 U10245 ( .C1(n9297), .C2(n9329), .A(n9148), .B(n9147), .ZN(n9149)
         );
  OAI21_X1 U10246 ( .B1(n9333), .B2(n9300), .A(n9149), .ZN(P2_U3271) );
  OAI21_X1 U10247 ( .B1(n9150), .B2(n9152), .A(n9151), .ZN(n9338) );
  INV_X1 U10248 ( .A(n9338), .ZN(n9167) );
  OAI211_X1 U10249 ( .C1(n5105), .C2(n9154), .A(n9153), .B(n10822), .ZN(n9157)
         );
  NAND2_X1 U10250 ( .A1(n9155), .A2(n9254), .ZN(n9156) );
  OAI211_X1 U10251 ( .C1(n9158), .C2(n9270), .A(n9157), .B(n9156), .ZN(n9337)
         );
  OAI21_X1 U10252 ( .B1(n9160), .B2(n9334), .A(n9159), .ZN(n9335) );
  AOI22_X1 U10253 ( .A1(n9303), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9161), .B2(
        n9202), .ZN(n9164) );
  NAND2_X1 U10254 ( .A1(n9162), .A2(n9292), .ZN(n9163) );
  OAI211_X1 U10255 ( .C1(n9335), .C2(n10818), .A(n9164), .B(n9163), .ZN(n9165)
         );
  AOI21_X1 U10256 ( .B1(n9337), .B2(n10829), .A(n9165), .ZN(n9166) );
  OAI21_X1 U10257 ( .B1(n9167), .B2(n9300), .A(n9166), .ZN(P2_U3272) );
  OAI21_X1 U10258 ( .B1(n5051), .B2(n5229), .A(n5206), .ZN(n9169) );
  AOI222_X1 U10259 ( .A1(n10822), .A2(n9169), .B1(n9168), .B2(n10821), .C1(
        n9197), .C2(n9254), .ZN(n9344) );
  INV_X1 U10260 ( .A(n9346), .ZN(n9172) );
  NAND2_X1 U10261 ( .A1(n9171), .A2(n5229), .ZN(n9340) );
  NAND3_X1 U10262 ( .A1(n9172), .A2(n10827), .A3(n9340), .ZN(n9178) );
  XNOR2_X1 U10263 ( .A(n9180), .B(n9341), .ZN(n9342) );
  AOI22_X1 U10264 ( .A1(n9303), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9173), .B2(
        n9202), .ZN(n9174) );
  OAI21_X1 U10265 ( .B1(n9175), .B2(n10819), .A(n9174), .ZN(n9176) );
  AOI21_X1 U10266 ( .B1(n9342), .B2(n9226), .A(n9176), .ZN(n9177) );
  OAI211_X1 U10267 ( .C1(n9303), .C2(n9344), .A(n9178), .B(n9177), .ZN(
        P2_U3273) );
  XNOR2_X1 U10268 ( .A(n9179), .B(n9185), .ZN(n9351) );
  AOI21_X1 U10269 ( .B1(n9347), .B2(n9199), .A(n9180), .ZN(n9348) );
  INV_X1 U10270 ( .A(n9347), .ZN(n9184) );
  INV_X1 U10271 ( .A(n9181), .ZN(n9182) );
  AOI22_X1 U10272 ( .A1(n9303), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9182), .B2(
        n9202), .ZN(n9183) );
  OAI21_X1 U10273 ( .B1(n9184), .B2(n10819), .A(n9183), .ZN(n9192) );
  AOI21_X1 U10274 ( .B1(n9186), .B2(n9185), .A(n9264), .ZN(n9190) );
  OAI22_X1 U10275 ( .A1(n9187), .A2(n9270), .B1(n9213), .B2(n9272), .ZN(n9188)
         );
  AOI21_X1 U10276 ( .B1(n9190), .B2(n9189), .A(n9188), .ZN(n9350) );
  NOR2_X1 U10277 ( .A1(n9350), .A2(n9303), .ZN(n9191) );
  AOI211_X1 U10278 ( .C1(n9348), .C2(n9226), .A(n9192), .B(n9191), .ZN(n9193)
         );
  OAI21_X1 U10279 ( .B1(n9351), .B2(n9300), .A(n9193), .ZN(P2_U3274) );
  XNOR2_X1 U10280 ( .A(n9195), .B(n9194), .ZN(n9198) );
  AOI222_X1 U10281 ( .A1(n10822), .A2(n9198), .B1(n9197), .B2(n10821), .C1(
        n9196), .C2(n9254), .ZN(n9355) );
  INV_X1 U10282 ( .A(n9199), .ZN(n9200) );
  AOI21_X1 U10283 ( .B1(n9352), .B2(n9201), .A(n9200), .ZN(n9353) );
  AOI22_X1 U10284 ( .A1(n9303), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9203), .B2(
        n9202), .ZN(n9204) );
  OAI21_X1 U10285 ( .B1(n9205), .B2(n10819), .A(n9204), .ZN(n9209) );
  AOI21_X1 U10286 ( .B1(n9207), .B2(n9206), .A(n5082), .ZN(n9356) );
  NOR2_X1 U10287 ( .A1(n9356), .A2(n9300), .ZN(n9208) );
  AOI211_X1 U10288 ( .C1(n9353), .C2(n9226), .A(n9209), .B(n9208), .ZN(n9210)
         );
  OAI21_X1 U10289 ( .B1(n9303), .B2(n9355), .A(n9210), .ZN(P2_U3275) );
  XNOR2_X1 U10290 ( .A(n9211), .B(n9215), .ZN(n9220) );
  OAI22_X1 U10291 ( .A1(n9213), .A2(n9270), .B1(n9212), .B2(n9272), .ZN(n9219)
         );
  OAI211_X1 U10292 ( .C1(n9216), .C2(n9215), .A(n9214), .B(n10980), .ZN(n9217)
         );
  INV_X1 U10293 ( .A(n9217), .ZN(n9218) );
  AOI211_X1 U10294 ( .C1(n10822), .C2(n9220), .A(n9219), .B(n9218), .ZN(n9360)
         );
  XNOR2_X1 U10295 ( .A(n9237), .B(n9357), .ZN(n9358) );
  NOR2_X1 U10296 ( .A1(n9221), .A2(n10819), .ZN(n9225) );
  OAI22_X1 U10297 ( .A1(n10829), .A2(n9223), .B1(n9222), .B2(n10823), .ZN(
        n9224) );
  AOI211_X1 U10298 ( .C1(n9358), .C2(n9226), .A(n9225), .B(n9224), .ZN(n9227)
         );
  OAI21_X1 U10299 ( .B1(n9360), .B2(n9303), .A(n9227), .ZN(P2_U3276) );
  NAND2_X1 U10300 ( .A1(n9228), .A2(n9229), .ZN(n9230) );
  INV_X1 U10301 ( .A(n9366), .ZN(n9244) );
  AOI22_X1 U10302 ( .A1(n9361), .A2(n9292), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n9303), .ZN(n9243) );
  XNOR2_X1 U10303 ( .A(n9232), .B(n5465), .ZN(n9235) );
  OAI22_X1 U10304 ( .A1(n9271), .A2(n9272), .B1(n9233), .B2(n9270), .ZN(n9234)
         );
  AOI21_X1 U10305 ( .B1(n9235), .B2(n10822), .A(n9234), .ZN(n9364) );
  INV_X1 U10306 ( .A(n9364), .ZN(n9241) );
  OAI21_X1 U10307 ( .B1(n5118), .B2(n9236), .A(n10881), .ZN(n9238) );
  OR2_X1 U10308 ( .A1(n9238), .A2(n9237), .ZN(n9362) );
  OAI22_X1 U10309 ( .A1(n9362), .A2(n8233), .B1(n10823), .B2(n9239), .ZN(n9240) );
  OAI21_X1 U10310 ( .B1(n9241), .B2(n9240), .A(n10829), .ZN(n9242) );
  OAI211_X1 U10311 ( .C1(n9244), .C2(n9300), .A(n9243), .B(n9242), .ZN(
        P2_U3277) );
  AND2_X1 U10312 ( .A1(n5112), .A2(n9369), .ZN(n9245) );
  OR2_X1 U10313 ( .A1(n9245), .A2(n5118), .ZN(n9370) );
  AOI22_X1 U10314 ( .A1(n9247), .A2(n10980), .B1(n9246), .B2(n10822), .ZN(
        n9251) );
  OAI22_X1 U10315 ( .A1(n9247), .A2(n10990), .B1(n9264), .B2(n9246), .ZN(n9248) );
  INV_X1 U10316 ( .A(n9248), .ZN(n9250) );
  MUX2_X1 U10317 ( .A(n9251), .B(n9250), .S(n9249), .Z(n9256) );
  AOI22_X1 U10318 ( .A1(n9254), .A2(n9253), .B1(n9252), .B2(n10821), .ZN(n9255) );
  NAND2_X1 U10319 ( .A1(n9256), .A2(n9255), .ZN(n9372) );
  NOR2_X1 U10320 ( .A1(n10823), .A2(n9257), .ZN(n9258) );
  OAI21_X1 U10321 ( .B1(n9372), .B2(n9258), .A(n10829), .ZN(n9260) );
  AOI22_X1 U10322 ( .A1(n9369), .A2(n9292), .B1(P2_REG2_REG_18__SCAN_IN), .B2(
        n9303), .ZN(n9259) );
  OAI211_X1 U10323 ( .C1(n9370), .C2(n10818), .A(n9260), .B(n9259), .ZN(
        P2_U3278) );
  INV_X1 U10324 ( .A(n9266), .ZN(n9263) );
  OAI22_X1 U10325 ( .A1(n9263), .A2(n10990), .B1(n9264), .B2(n9262), .ZN(n9269) );
  INV_X1 U10326 ( .A(n9262), .ZN(n9265) );
  OAI22_X1 U10327 ( .A1(n9266), .A2(n10990), .B1(n9265), .B2(n9264), .ZN(n9268) );
  MUX2_X1 U10328 ( .A(n9269), .B(n9268), .S(n9267), .Z(n9275) );
  OAI22_X1 U10329 ( .A1(n9273), .A2(n9272), .B1(n9271), .B2(n9270), .ZN(n9274)
         );
  NOR2_X1 U10330 ( .A1(n9275), .A2(n9274), .ZN(n9377) );
  OAI22_X1 U10331 ( .A1(n10829), .A2(n9277), .B1(n9276), .B2(n10823), .ZN(
        n9278) );
  AOI21_X1 U10332 ( .B1(n9375), .B2(n9292), .A(n9278), .ZN(n9282) );
  AOI21_X1 U10333 ( .B1(n9296), .B2(n9375), .A(n10994), .ZN(n9279) );
  NAND2_X1 U10334 ( .A1(n9279), .A2(n5112), .ZN(n9376) );
  OR2_X1 U10335 ( .A1(n9376), .A2(n9280), .ZN(n9281) );
  OAI211_X1 U10336 ( .C1(n9377), .C2(n9303), .A(n9282), .B(n9281), .ZN(
        P2_U3279) );
  XNOR2_X1 U10337 ( .A(n9284), .B(n9283), .ZN(n9286) );
  AOI21_X1 U10338 ( .B1(n9286), .B2(n10822), .A(n9285), .ZN(n9381) );
  OAI21_X1 U10339 ( .B1(n9288), .B2(n8211), .A(n9287), .ZN(n9382) );
  OAI22_X1 U10340 ( .A1(n10829), .A2(n9290), .B1(n9289), .B2(n10823), .ZN(
        n9291) );
  AOI21_X1 U10341 ( .B1(n9379), .B2(n9292), .A(n9291), .ZN(n9299) );
  OR2_X1 U10342 ( .A1(n9294), .A2(n9293), .ZN(n9295) );
  AND3_X1 U10343 ( .A1(n9296), .A2(n10881), .A3(n9295), .ZN(n9378) );
  NAND2_X1 U10344 ( .A1(n9378), .A2(n9297), .ZN(n9298) );
  OAI211_X1 U10345 ( .C1(n9382), .C2(n9300), .A(n9299), .B(n9298), .ZN(n9301)
         );
  INV_X1 U10346 ( .A(n9301), .ZN(n9302) );
  OAI21_X1 U10347 ( .B1(n9303), .B2(n9381), .A(n9302), .ZN(P2_U3280) );
  NAND2_X1 U10348 ( .A1(n9304), .A2(n10971), .ZN(n9305) );
  OAI211_X1 U10349 ( .C1(n9306), .C2(n10994), .A(n9305), .B(n9309), .ZN(n9394)
         );
  MUX2_X1 U10350 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9394), .S(n11002), .Z(
        P2_U3551) );
  NAND2_X1 U10351 ( .A1(n9307), .A2(n10971), .ZN(n9308) );
  OAI211_X1 U10352 ( .C1(n9310), .C2(n10994), .A(n9309), .B(n9308), .ZN(n9395)
         );
  MUX2_X1 U10353 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9395), .S(n11002), .Z(
        P2_U3550) );
  AOI22_X1 U10354 ( .A1(n9312), .A2(n10881), .B1(n10971), .B2(n9311), .ZN(
        n9313) );
  OAI211_X1 U10355 ( .C1(n9315), .C2(n10990), .A(n9314), .B(n9313), .ZN(n9396)
         );
  MUX2_X1 U10356 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9396), .S(n11002), .Z(
        P2_U3549) );
  AOI22_X1 U10357 ( .A1(n9317), .A2(n10881), .B1(n10971), .B2(n9316), .ZN(
        n9318) );
  OAI211_X1 U10358 ( .C1(n9320), .C2(n10990), .A(n9319), .B(n9318), .ZN(n9397)
         );
  MUX2_X1 U10359 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9397), .S(n11002), .Z(
        P2_U3548) );
  AOI22_X1 U10360 ( .A1(n9322), .A2(n10881), .B1(n10971), .B2(n9321), .ZN(
        n9323) );
  OAI211_X1 U10361 ( .C1(n9325), .C2(n10990), .A(n9324), .B(n9323), .ZN(n9398)
         );
  MUX2_X1 U10362 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9398), .S(n11002), .Z(
        P2_U3547) );
  OAI211_X1 U10363 ( .C1(n9328), .C2(n10992), .A(n9327), .B(n9326), .ZN(n9399)
         );
  MUX2_X1 U10364 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9399), .S(n11002), .Z(
        P2_U3546) );
  AOI21_X1 U10365 ( .B1(n10971), .B2(n9330), .A(n9329), .ZN(n9331) );
  OAI211_X1 U10366 ( .C1(n9333), .C2(n10990), .A(n9332), .B(n9331), .ZN(n9400)
         );
  MUX2_X1 U10367 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9400), .S(n11002), .Z(
        P2_U3545) );
  OAI22_X1 U10368 ( .A1(n9335), .A2(n10994), .B1(n9334), .B2(n10992), .ZN(
        n9336) );
  AOI211_X1 U10369 ( .C1(n9338), .C2(n10980), .A(n9337), .B(n9336), .ZN(n9339)
         );
  INV_X1 U10370 ( .A(n9339), .ZN(n9401) );
  MUX2_X1 U10371 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9401), .S(n11002), .Z(
        P2_U3544) );
  NAND2_X1 U10372 ( .A1(n9340), .A2(n10980), .ZN(n9345) );
  AOI22_X1 U10373 ( .A1(n9342), .A2(n10881), .B1(n10971), .B2(n9341), .ZN(
        n9343) );
  OAI211_X1 U10374 ( .C1(n9346), .C2(n9345), .A(n9344), .B(n9343), .ZN(n9402)
         );
  MUX2_X1 U10375 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9402), .S(n11002), .Z(
        P2_U3543) );
  AOI22_X1 U10376 ( .A1(n9348), .A2(n10881), .B1(n10971), .B2(n9347), .ZN(
        n9349) );
  OAI211_X1 U10377 ( .C1(n9351), .C2(n10990), .A(n9350), .B(n9349), .ZN(n9403)
         );
  MUX2_X1 U10378 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9403), .S(n11002), .Z(
        P2_U3542) );
  AOI22_X1 U10379 ( .A1(n9353), .A2(n10881), .B1(n10971), .B2(n9352), .ZN(
        n9354) );
  OAI211_X1 U10380 ( .C1(n9356), .C2(n10990), .A(n9355), .B(n9354), .ZN(n9404)
         );
  MUX2_X1 U10381 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9404), .S(n11002), .Z(
        P2_U3541) );
  AOI22_X1 U10382 ( .A1(n9358), .A2(n10881), .B1(n10971), .B2(n9357), .ZN(
        n9359) );
  NAND2_X1 U10383 ( .A1(n9360), .A2(n9359), .ZN(n9405) );
  MUX2_X1 U10384 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9405), .S(n11002), .Z(
        P2_U3540) );
  NAND2_X1 U10385 ( .A1(n9361), .A2(n10971), .ZN(n9363) );
  NAND3_X1 U10386 ( .A1(n9364), .A2(n9363), .A3(n9362), .ZN(n9365) );
  AOI21_X1 U10387 ( .B1(n9366), .B2(n10980), .A(n9365), .ZN(n9406) );
  MUX2_X1 U10388 ( .A(n9367), .B(n9406), .S(n11002), .Z(n9368) );
  INV_X1 U10389 ( .A(n9368), .ZN(P2_U3539) );
  OAI22_X1 U10390 ( .A1(n9370), .A2(n10994), .B1(n5320), .B2(n10992), .ZN(
        n9371) );
  NOR2_X1 U10391 ( .A1(n9372), .A2(n9371), .ZN(n9409) );
  MUX2_X1 U10392 ( .A(n9373), .B(n9409), .S(n11002), .Z(n9374) );
  INV_X1 U10393 ( .A(n9374), .ZN(P2_U3538) );
  OAI211_X1 U10394 ( .C1(n5319), .C2(n10992), .A(n9377), .B(n9376), .ZN(n9412)
         );
  MUX2_X1 U10395 ( .A(n9412), .B(P2_REG1_REG_17__SCAN_IN), .S(n11000), .Z(
        P2_U3537) );
  AOI21_X1 U10396 ( .B1(n10971), .B2(n9379), .A(n9378), .ZN(n9380) );
  OAI211_X1 U10397 ( .C1(n9382), .C2(n10990), .A(n9381), .B(n9380), .ZN(n9413)
         );
  MUX2_X1 U10398 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9413), .S(n11002), .Z(
        P2_U3536) );
  AOI22_X1 U10399 ( .A1(n9384), .A2(n10881), .B1(n10971), .B2(n9383), .ZN(
        n9385) );
  OAI211_X1 U10400 ( .C1(n9387), .C2(n10990), .A(n9386), .B(n9385), .ZN(n9414)
         );
  MUX2_X1 U10401 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9414), .S(n11002), .Z(
        P2_U3535) );
  INV_X1 U10402 ( .A(n9388), .ZN(n9393) );
  AOI22_X1 U10403 ( .A1(n9390), .A2(n10881), .B1(n10971), .B2(n9389), .ZN(
        n9391) );
  OAI211_X1 U10404 ( .C1(n9393), .C2(n10990), .A(n9392), .B(n9391), .ZN(n9415)
         );
  MUX2_X1 U10405 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9415), .S(n11002), .Z(
        P2_U3534) );
  MUX2_X1 U10406 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9394), .S(n11006), .Z(
        P2_U3519) );
  MUX2_X1 U10407 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9395), .S(n11006), .Z(
        P2_U3518) );
  MUX2_X1 U10408 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9396), .S(n11006), .Z(
        P2_U3517) );
  MUX2_X1 U10409 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9397), .S(n11006), .Z(
        P2_U3516) );
  MUX2_X1 U10410 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9398), .S(n11006), .Z(
        P2_U3515) );
  MUX2_X1 U10411 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9399), .S(n11006), .Z(
        P2_U3514) );
  MUX2_X1 U10412 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9400), .S(n11006), .Z(
        P2_U3513) );
  MUX2_X1 U10413 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9401), .S(n11006), .Z(
        P2_U3512) );
  MUX2_X1 U10414 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9402), .S(n11006), .Z(
        P2_U3511) );
  MUX2_X1 U10415 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9403), .S(n11006), .Z(
        P2_U3510) );
  MUX2_X1 U10416 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9404), .S(n11006), .Z(
        P2_U3509) );
  MUX2_X1 U10417 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9405), .S(n11006), .Z(
        P2_U3508) );
  MUX2_X1 U10418 ( .A(n9407), .B(n9406), .S(n11006), .Z(n9408) );
  INV_X1 U10419 ( .A(n9408), .ZN(P2_U3507) );
  INV_X1 U10420 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9410) );
  MUX2_X1 U10421 ( .A(n9410), .B(n9409), .S(n11006), .Z(n9411) );
  INV_X1 U10422 ( .A(n9411), .ZN(P2_U3505) );
  MUX2_X1 U10423 ( .A(n9412), .B(P2_REG0_REG_17__SCAN_IN), .S(n11003), .Z(
        P2_U3502) );
  MUX2_X1 U10424 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9413), .S(n11006), .Z(
        P2_U3499) );
  MUX2_X1 U10425 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9414), .S(n11006), .Z(
        P2_U3496) );
  MUX2_X1 U10426 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9415), .S(n11006), .Z(
        P2_U3493) );
  NAND3_X1 U10427 ( .A1(n9416), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n9418) );
  OAI22_X1 U10428 ( .A1(n5235), .A2(n9418), .B1(n9417), .B2(n5036), .ZN(n9419)
         );
  AOI21_X1 U10429 ( .B1(n10260), .B2(n9420), .A(n9419), .ZN(n9421) );
  INV_X1 U10430 ( .A(n9421), .ZN(P2_U3327) );
  OAI222_X1 U10431 ( .A1(n8494), .A2(n10268), .B1(n9423), .B2(P2_U3152), .C1(
        n9422), .C2(n5036), .ZN(P2_U3329) );
  MUX2_X1 U10432 ( .A(n9424), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10433 ( .A(n9427), .B(n9426), .ZN(n9428) );
  XNOR2_X1 U10434 ( .A(n9425), .B(n9428), .ZN(n9436) );
  NOR2_X1 U10435 ( .A1(n9559), .A2(n9429), .ZN(n9430) );
  AOI211_X1 U10436 ( .C1(n9561), .C2(n9842), .A(n9431), .B(n9430), .ZN(n9432)
         );
  OAI21_X1 U10437 ( .B1(n9564), .B2(n9433), .A(n9432), .ZN(n9434) );
  AOI21_X1 U10438 ( .B1(n10228), .B2(n9566), .A(n9434), .ZN(n9435) );
  OAI21_X1 U10439 ( .B1(n9436), .B2(n9569), .A(n9435), .ZN(P1_U3213) );
  XNOR2_X1 U10440 ( .A(n9439), .B(n9438), .ZN(n9440) );
  XNOR2_X1 U10441 ( .A(n9437), .B(n9440), .ZN(n9445) );
  AOI22_X1 U10442 ( .A1(n10025), .A2(n9561), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9442) );
  NAND2_X1 U10443 ( .A1(n9996), .A2(n9505), .ZN(n9441) );
  OAI211_X1 U10444 ( .C1(n9974), .C2(n9559), .A(n9442), .B(n9441), .ZN(n9443)
         );
  AOI21_X1 U10445 ( .B1(n10184), .B2(n9566), .A(n9443), .ZN(n9444) );
  OAI21_X1 U10446 ( .B1(n9445), .B2(n9569), .A(n9444), .ZN(P1_U3214) );
  NOR2_X1 U10447 ( .A1(n9447), .A2(n5163), .ZN(n9448) );
  XNOR2_X1 U10448 ( .A(n9449), .B(n9448), .ZN(n9455) );
  NAND2_X1 U10449 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9894) );
  NAND2_X1 U10450 ( .A1(n9561), .A2(n10110), .ZN(n9450) );
  OAI211_X1 U10451 ( .C1(n9451), .C2(n9559), .A(n9894), .B(n9450), .ZN(n9453)
         );
  NOR2_X1 U10452 ( .A1(n10064), .A2(n9535), .ZN(n9452) );
  AOI211_X1 U10453 ( .C1(n10062), .C2(n9505), .A(n9453), .B(n9452), .ZN(n9454)
         );
  OAI21_X1 U10454 ( .B1(n9455), .B2(n9569), .A(n9454), .ZN(P1_U3217) );
  OAI21_X1 U10455 ( .B1(n9458), .B2(n9457), .A(n9456), .ZN(n9459) );
  NAND2_X1 U10456 ( .A1(n9459), .A2(n9525), .ZN(n9463) );
  AOI22_X1 U10457 ( .A1(n9561), .A2(n6891), .B1(n9566), .B2(n10839), .ZN(n9462) );
  AOI22_X1 U10458 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(n9460), .B1(n9532), .B2(
        n9850), .ZN(n9461) );
  NAND3_X1 U10459 ( .A1(n9463), .A2(n9462), .A3(n9461), .ZN(P1_U3220) );
  OAI21_X1 U10460 ( .B1(n9465), .B2(n5115), .A(n9464), .ZN(n9466) );
  OAI21_X1 U10461 ( .B1(n9467), .B2(n5115), .A(n9466), .ZN(n9468) );
  NAND2_X1 U10462 ( .A1(n9468), .A2(n9525), .ZN(n9473) );
  AOI22_X1 U10463 ( .A1(n10068), .A2(n9561), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9469) );
  OAI21_X1 U10464 ( .B1(n9470), .B2(n9559), .A(n9469), .ZN(n9471) );
  AOI21_X1 U10465 ( .B1(n10029), .B2(n9505), .A(n9471), .ZN(n9472) );
  OAI211_X1 U10466 ( .C1(n5314), .C2(n9535), .A(n9473), .B(n9472), .ZN(
        P1_U3221) );
  XOR2_X1 U10467 ( .A(n9475), .B(n9474), .Z(n9476) );
  XNOR2_X1 U10468 ( .A(n9477), .B(n9476), .ZN(n9482) );
  NAND2_X1 U10469 ( .A1(n10002), .A2(n9561), .ZN(n9479) );
  AOI22_X1 U10470 ( .A1(n9532), .A2(n9940), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9478) );
  OAI211_X1 U10471 ( .C1(n9564), .C2(n9965), .A(n9479), .B(n9478), .ZN(n9480)
         );
  AOI21_X1 U10472 ( .B1(n10175), .B2(n9566), .A(n9480), .ZN(n9481) );
  OAI21_X1 U10473 ( .B1(n9482), .B2(n9569), .A(n9481), .ZN(P1_U3223) );
  INV_X1 U10474 ( .A(n10223), .ZN(n10145) );
  INV_X1 U10475 ( .A(n9483), .ZN(n9487) );
  AOI21_X1 U10476 ( .B1(n9554), .B2(n9485), .A(n9484), .ZN(n9486) );
  OAI21_X1 U10477 ( .B1(n9487), .B2(n9486), .A(n9525), .ZN(n9492) );
  NAND2_X1 U10478 ( .A1(n9561), .A2(n10132), .ZN(n9489) );
  OAI211_X1 U10479 ( .C1(n10082), .C2(n9559), .A(n9489), .B(n9488), .ZN(n9490)
         );
  AOI21_X1 U10480 ( .B1(n10140), .B2(n9505), .A(n9490), .ZN(n9491) );
  OAI211_X1 U10481 ( .C1(n10145), .C2(n9535), .A(n9492), .B(n9491), .ZN(
        P1_U3224) );
  INV_X1 U10482 ( .A(n10216), .ZN(n10119) );
  AND3_X1 U10483 ( .A1(n9483), .A2(n9494), .A3(n9493), .ZN(n9495) );
  OAI21_X1 U10484 ( .B1(n9496), .B2(n9495), .A(n9525), .ZN(n9502) );
  INV_X1 U10485 ( .A(n9497), .ZN(n10116) );
  NAND2_X1 U10486 ( .A1(n9561), .A2(n10109), .ZN(n9498) );
  NAND2_X1 U10487 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9853) );
  OAI211_X1 U10488 ( .C1(n9499), .C2(n9559), .A(n9498), .B(n9853), .ZN(n9500)
         );
  AOI21_X1 U10489 ( .B1(n10116), .B2(n9505), .A(n9500), .ZN(n9501) );
  OAI211_X1 U10490 ( .C1(n10119), .C2(n9535), .A(n9502), .B(n9501), .ZN(
        P1_U3226) );
  XOR2_X1 U10491 ( .A(n9504), .B(n9503), .Z(n9511) );
  AOI22_X1 U10492 ( .A1(n9532), .A2(n9982), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9507) );
  NAND2_X1 U10493 ( .A1(n9987), .A2(n9505), .ZN(n9506) );
  OAI211_X1 U10494 ( .C1(n9508), .C2(n9529), .A(n9507), .B(n9506), .ZN(n9509)
         );
  AOI21_X1 U10495 ( .B1(n10179), .B2(n9566), .A(n9509), .ZN(n9510) );
  OAI21_X1 U10496 ( .B1(n9511), .B2(n9569), .A(n9510), .ZN(P1_U3227) );
  XNOR2_X1 U10497 ( .A(n9513), .B(n9512), .ZN(n9514) );
  XNOR2_X1 U10498 ( .A(n9515), .B(n9514), .ZN(n9521) );
  OAI22_X1 U10499 ( .A1(n10038), .A2(n9559), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9516), .ZN(n9517) );
  AOI21_X1 U10500 ( .B1(n9561), .B2(n10040), .A(n9517), .ZN(n9518) );
  OAI21_X1 U10501 ( .B1(n9564), .B2(n10051), .A(n9518), .ZN(n9519) );
  AOI21_X1 U10502 ( .B1(n10198), .B2(n9566), .A(n9519), .ZN(n9520) );
  OAI21_X1 U10503 ( .B1(n9521), .B2(n9569), .A(n9520), .ZN(P1_U3231) );
  OAI21_X1 U10504 ( .B1(n9524), .B2(n9523), .A(n9522), .ZN(n9526) );
  NAND2_X1 U10505 ( .A1(n9526), .A2(n9525), .ZN(n9534) );
  NOR2_X1 U10506 ( .A1(n9527), .A2(n9564), .ZN(n9531) );
  OAI22_X1 U10507 ( .A1(n10038), .A2(n9529), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9528), .ZN(n9530) );
  AOI211_X1 U10508 ( .C1(n10015), .C2(n9532), .A(n9531), .B(n9530), .ZN(n9533)
         );
  OAI211_X1 U10509 ( .C1(n10012), .C2(n9535), .A(n9534), .B(n9533), .ZN(
        P1_U3233) );
  NAND2_X1 U10510 ( .A1(n5570), .A2(n9536), .ZN(n9538) );
  XNOR2_X1 U10511 ( .A(n9538), .B(n9537), .ZN(n9543) );
  NAND2_X1 U10512 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9878) );
  OAI21_X1 U10513 ( .B1(n10084), .B2(n9559), .A(n9878), .ZN(n9539) );
  AOI21_X1 U10514 ( .B1(n9561), .B2(n10129), .A(n9539), .ZN(n9540) );
  OAI21_X1 U10515 ( .B1(n9564), .B2(n10091), .A(n9540), .ZN(n9541) );
  AOI21_X1 U10516 ( .B1(n10096), .B2(n9566), .A(n9541), .ZN(n9542) );
  OAI21_X1 U10517 ( .B1(n9543), .B2(n9569), .A(n9542), .ZN(P1_U3236) );
  XNOR2_X1 U10518 ( .A(n9544), .B(n9545), .ZN(n9552) );
  INV_X1 U10519 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9546) );
  OAI22_X1 U10520 ( .A1(n9559), .A2(n9547), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9546), .ZN(n9548) );
  AOI21_X1 U10521 ( .B1(n9561), .B2(n9982), .A(n9548), .ZN(n9549) );
  OAI21_X1 U10522 ( .B1(n9564), .B2(n9947), .A(n9549), .ZN(n9550) );
  AOI21_X1 U10523 ( .B1(n10168), .B2(n9566), .A(n9550), .ZN(n9551) );
  OAI21_X1 U10524 ( .B1(n9552), .B2(n9569), .A(n9551), .ZN(P1_U3238) );
  NAND2_X1 U10525 ( .A1(n9554), .A2(n9553), .ZN(n9555) );
  XOR2_X1 U10526 ( .A(n9556), .B(n9555), .Z(n9570) );
  OAI21_X1 U10527 ( .B1(n9559), .B2(n9558), .A(n9557), .ZN(n9560) );
  AOI21_X1 U10528 ( .B1(n9561), .B2(n9841), .A(n9560), .ZN(n9562) );
  OAI21_X1 U10529 ( .B1(n9564), .B2(n9563), .A(n9562), .ZN(n9565) );
  AOI21_X1 U10530 ( .B1(n9567), .B2(n9566), .A(n9565), .ZN(n9568) );
  OAI21_X1 U10531 ( .B1(n9570), .B2(n9569), .A(n9568), .ZN(P1_U3239) );
  NAND2_X1 U10532 ( .A1(n10260), .A2(n6176), .ZN(n9572) );
  NAND2_X1 U10533 ( .A1(n9574), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n9571) );
  INV_X1 U10534 ( .A(n9902), .ZN(n9645) );
  NAND2_X1 U10535 ( .A1(n10149), .A2(n9645), .ZN(n9747) );
  NAND2_X1 U10536 ( .A1(n9573), .A2(n6176), .ZN(n9576) );
  NAND2_X1 U10537 ( .A1(n9574), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9575) );
  NAND2_X1 U10538 ( .A1(n11019), .A2(n9839), .ZN(n9647) );
  NAND2_X1 U10539 ( .A1(n9747), .A2(n9647), .ZN(n9793) );
  NAND2_X1 U10540 ( .A1(n9754), .A2(n9577), .ZN(n9810) );
  NAND2_X1 U10541 ( .A1(n9649), .A2(n5624), .ZN(n9578) );
  NAND3_X1 U10542 ( .A1(n9751), .A2(n9650), .A3(n9578), .ZN(n9812) );
  NAND2_X1 U10543 ( .A1(n9653), .A2(n9655), .ZN(n9582) );
  OAI211_X1 U10544 ( .C1(n9656), .C2(n9582), .A(n9651), .B(n9654), .ZN(n9579)
         );
  INV_X1 U10545 ( .A(n9579), .ZN(n9580) );
  NAND2_X1 U10546 ( .A1(n9580), .A2(n9649), .ZN(n9809) );
  INV_X1 U10547 ( .A(n9732), .ZN(n9581) );
  OR2_X1 U10548 ( .A1(n9582), .A2(n9581), .ZN(n9807) );
  NAND2_X1 U10549 ( .A1(n9721), .A2(n9583), .ZN(n9584) );
  NAND2_X1 U10550 ( .A1(n9584), .A2(n9615), .ZN(n9723) );
  NAND2_X1 U10551 ( .A1(n9728), .A2(n9723), .ZN(n9635) );
  INV_X1 U10552 ( .A(n9715), .ZN(n9585) );
  OR2_X1 U10553 ( .A1(n9635), .A2(n9585), .ZN(n9616) );
  AND2_X1 U10554 ( .A1(n9709), .A2(n9704), .ZN(n9586) );
  NAND2_X1 U10555 ( .A1(n9713), .A2(n9586), .ZN(n9617) );
  INV_X1 U10556 ( .A(n9695), .ZN(n9591) );
  NAND2_X1 U10557 ( .A1(n9674), .A2(n9670), .ZN(n9587) );
  NAND2_X1 U10558 ( .A1(n9587), .A2(n9673), .ZN(n9588) );
  AND3_X1 U10559 ( .A1(n9686), .A2(n9679), .A3(n9588), .ZN(n9589) );
  AND2_X1 U10560 ( .A1(n9683), .A2(n9589), .ZN(n9619) );
  NAND4_X1 U10561 ( .A1(n9694), .A2(n9619), .A3(n9659), .A4(n9661), .ZN(n9590)
         );
  OR3_X1 U10562 ( .A1(n9617), .A2(n9591), .A3(n9590), .ZN(n9592) );
  NOR2_X1 U10563 ( .A1(n9616), .A2(n9592), .ZN(n9803) );
  NAND2_X1 U10564 ( .A1(n9851), .A2(n9593), .ZN(n9596) );
  NAND2_X1 U10565 ( .A1(n6891), .A2(n9594), .ZN(n9595) );
  AND3_X1 U10566 ( .A1(n9596), .A2(n9595), .A3(n9760), .ZN(n9599) );
  NAND2_X1 U10567 ( .A1(n7246), .A2(n10870), .ZN(n9597) );
  OAI211_X1 U10568 ( .C1(n9600), .C2(n9599), .A(n9598), .B(n9597), .ZN(n9604)
         );
  INV_X1 U10569 ( .A(n9601), .ZN(n9603) );
  NAND3_X1 U10570 ( .A1(n9604), .A2(n9603), .A3(n9602), .ZN(n9607) );
  NAND3_X1 U10571 ( .A1(n9607), .A2(n9606), .A3(n9605), .ZN(n9610) );
  NAND3_X1 U10572 ( .A1(n9610), .A2(n9609), .A3(n9608), .ZN(n9612) );
  NAND2_X1 U10573 ( .A1(n9612), .A2(n9611), .ZN(n9613) );
  AND2_X1 U10574 ( .A1(n9803), .A2(n9613), .ZN(n9637) );
  NAND2_X1 U10575 ( .A1(n9615), .A2(n9614), .ZN(n9722) );
  INV_X1 U10576 ( .A(n9722), .ZN(n9636) );
  NAND2_X1 U10577 ( .A1(n10012), .A2(n10025), .ZN(n9727) );
  AND2_X1 U10578 ( .A1(n9733), .A2(n9727), .ZN(n9634) );
  INV_X1 U10579 ( .A(n9616), .ZN(n9632) );
  INV_X1 U10580 ( .A(n9617), .ZN(n9627) );
  NAND3_X1 U10581 ( .A1(n9673), .A2(n9660), .A3(n9669), .ZN(n9618) );
  NAND2_X1 U10582 ( .A1(n9619), .A2(n9618), .ZN(n9623) );
  INV_X1 U10583 ( .A(n9620), .ZN(n9621) );
  NAND3_X1 U10584 ( .A1(n9621), .A2(n9683), .A3(n9686), .ZN(n9622) );
  NAND4_X1 U10585 ( .A1(n9623), .A2(n9698), .A3(n9685), .A4(n9622), .ZN(n9624)
         );
  NAND3_X1 U10586 ( .A1(n9695), .A2(n9694), .A3(n9624), .ZN(n9625) );
  NAND3_X1 U10587 ( .A1(n9705), .A2(n9699), .A3(n9625), .ZN(n9626) );
  NAND2_X1 U10588 ( .A1(n9627), .A2(n9626), .ZN(n9630) );
  INV_X1 U10589 ( .A(n9708), .ZN(n9628) );
  NAND2_X1 U10590 ( .A1(n9713), .A2(n9628), .ZN(n9629) );
  NAND4_X1 U10591 ( .A1(n9630), .A2(n9629), .A3(n9716), .A4(n9712), .ZN(n9631)
         );
  NAND2_X1 U10592 ( .A1(n9632), .A2(n9631), .ZN(n9633) );
  OAI211_X1 U10593 ( .C1(n9636), .C2(n9635), .A(n9634), .B(n9633), .ZN(n9804)
         );
  NOR2_X1 U10594 ( .A1(n9637), .A2(n9804), .ZN(n9638) );
  NOR2_X1 U10595 ( .A1(n9807), .A2(n9638), .ZN(n9639) );
  NOR2_X1 U10596 ( .A1(n9809), .A2(n9639), .ZN(n9640) );
  NOR2_X1 U10597 ( .A1(n9812), .A2(n9640), .ZN(n9642) );
  INV_X1 U10598 ( .A(n11019), .ZN(n9900) );
  INV_X1 U10599 ( .A(n9839), .ZN(n9641) );
  NAND2_X1 U10600 ( .A1(n9900), .A2(n9641), .ZN(n9791) );
  OAI211_X1 U10601 ( .C1(n9810), .C2(n9642), .A(n9791), .B(n9756), .ZN(n9643)
         );
  INV_X1 U10602 ( .A(n9643), .ZN(n9644) );
  OR2_X1 U10603 ( .A1(n9793), .A2(n9644), .ZN(n9646) );
  OR2_X1 U10604 ( .A1(n10149), .A2(n9645), .ZN(n9819) );
  NAND2_X1 U10605 ( .A1(n9647), .A2(n9902), .ZN(n9648) );
  NAND2_X1 U10606 ( .A1(n9648), .A2(n10149), .ZN(n9817) );
  INV_X1 U10607 ( .A(n9731), .ZN(n9758) );
  MUX2_X1 U10608 ( .A(n9650), .B(n9649), .S(n9758), .Z(n9744) );
  MUX2_X1 U10609 ( .A(n9652), .B(n9651), .S(n9731), .Z(n9742) );
  INV_X1 U10610 ( .A(n9951), .ZN(n9944) );
  MUX2_X1 U10611 ( .A(n9654), .B(n9653), .S(n9731), .Z(n9740) );
  INV_X1 U10612 ( .A(n9970), .ZN(n9738) );
  MUX2_X1 U10613 ( .A(n9656), .B(n9655), .S(n9758), .Z(n9737) );
  NAND2_X1 U10614 ( .A1(n7562), .A2(n9731), .ZN(n9668) );
  NAND2_X1 U10615 ( .A1(n9661), .A2(n9758), .ZN(n9657) );
  NOR2_X1 U10616 ( .A1(n9658), .A2(n9657), .ZN(n9666) );
  MUX2_X1 U10617 ( .A(n9660), .B(n9659), .S(n9731), .Z(n9664) );
  INV_X1 U10618 ( .A(n9661), .ZN(n9662) );
  NAND3_X1 U10619 ( .A1(n7562), .A2(n9662), .A3(n9731), .ZN(n9663) );
  NAND3_X1 U10620 ( .A1(n9772), .A2(n9664), .A3(n9663), .ZN(n9665) );
  AOI21_X1 U10621 ( .B1(n9802), .B2(n9666), .A(n9665), .ZN(n9667) );
  OAI21_X1 U10622 ( .B1(n9802), .B2(n9668), .A(n9667), .ZN(n9672) );
  MUX2_X1 U10623 ( .A(n9670), .B(n9669), .S(n9731), .Z(n9671) );
  NAND3_X1 U10624 ( .A1(n9672), .A2(n9773), .A3(n9671), .ZN(n9677) );
  INV_X1 U10625 ( .A(n9775), .ZN(n9676) );
  MUX2_X1 U10626 ( .A(n9674), .B(n9673), .S(n9758), .Z(n9675) );
  NAND3_X1 U10627 ( .A1(n9677), .A2(n9676), .A3(n9675), .ZN(n9682) );
  MUX2_X1 U10628 ( .A(n9679), .B(n9678), .S(n9731), .Z(n9680) );
  AND2_X1 U10629 ( .A1(n9777), .A2(n9680), .ZN(n9681) );
  NAND2_X1 U10630 ( .A1(n9682), .A2(n9681), .ZN(n9687) );
  INV_X1 U10631 ( .A(n9683), .ZN(n9697) );
  AOI21_X1 U10632 ( .B1(n9687), .B2(n9684), .A(n9697), .ZN(n9689) );
  INV_X1 U10633 ( .A(n9685), .ZN(n9693) );
  AOI21_X1 U10634 ( .B1(n9687), .B2(n9686), .A(n9693), .ZN(n9688) );
  MUX2_X1 U10635 ( .A(n9689), .B(n9688), .S(n9731), .Z(n9691) );
  MUX2_X1 U10636 ( .A(n9698), .B(n9694), .S(n9758), .Z(n9690) );
  OAI21_X1 U10637 ( .B1(n9691), .B2(n9780), .A(n9690), .ZN(n9692) );
  NAND2_X1 U10638 ( .A1(n9692), .A2(n9782), .ZN(n9701) );
  AND2_X1 U10639 ( .A1(n9694), .A2(n9693), .ZN(n9696) );
  OAI21_X1 U10640 ( .B1(n9701), .B2(n9696), .A(n9695), .ZN(n9703) );
  AND2_X1 U10641 ( .A1(n9698), .A2(n9697), .ZN(n9700) );
  OAI21_X1 U10642 ( .B1(n9701), .B2(n9700), .A(n9699), .ZN(n9702) );
  MUX2_X1 U10643 ( .A(n9703), .B(n9702), .S(n9731), .Z(n9707) );
  MUX2_X1 U10644 ( .A(n9705), .B(n9704), .S(n9731), .Z(n9706) );
  OAI211_X1 U10645 ( .C1(n9707), .C2(n10123), .A(n10107), .B(n9706), .ZN(n9711) );
  MUX2_X1 U10646 ( .A(n9709), .B(n9708), .S(n9731), .Z(n9710) );
  AOI21_X1 U10647 ( .B1(n9711), .B2(n9710), .A(n10077), .ZN(n9719) );
  MUX2_X1 U10648 ( .A(n9713), .B(n9712), .S(n9731), .Z(n9714) );
  NAND2_X1 U10649 ( .A1(n10067), .A2(n9714), .ZN(n9718) );
  MUX2_X1 U10650 ( .A(n9716), .B(n9715), .S(n9731), .Z(n9717) );
  OAI21_X1 U10651 ( .B1(n9719), .B2(n9718), .A(n9717), .ZN(n9720) );
  NAND3_X1 U10652 ( .A1(n9720), .A2(n10037), .A3(n10023), .ZN(n9726) );
  INV_X1 U10653 ( .A(n10013), .ZN(n10007) );
  NAND2_X1 U10654 ( .A1(n9722), .A2(n9721), .ZN(n9724) );
  MUX2_X1 U10655 ( .A(n9724), .B(n9723), .S(n9731), .Z(n9725) );
  NAND3_X1 U10656 ( .A1(n9726), .A2(n10007), .A3(n9725), .ZN(n9730) );
  MUX2_X1 U10657 ( .A(n9728), .B(n9727), .S(n9731), .Z(n9729) );
  NAND3_X1 U10658 ( .A1(n9730), .A2(n10001), .A3(n9729), .ZN(n9735) );
  MUX2_X1 U10659 ( .A(n9733), .B(n9732), .S(n9731), .Z(n9734) );
  NAND3_X1 U10660 ( .A1(n9735), .A2(n9980), .A3(n9734), .ZN(n9736) );
  NAND3_X1 U10661 ( .A1(n9738), .A2(n9737), .A3(n9736), .ZN(n9739) );
  NAND3_X1 U10662 ( .A1(n9944), .A2(n9740), .A3(n9739), .ZN(n9741) );
  NAND3_X1 U10663 ( .A1(n9788), .A2(n9742), .A3(n9741), .ZN(n9743) );
  AND3_X1 U10664 ( .A1(n9919), .A2(n9744), .A3(n9743), .ZN(n9750) );
  OAI21_X1 U10665 ( .B1(n9810), .B2(n9750), .A(n9756), .ZN(n9745) );
  NAND2_X1 U10666 ( .A1(n9817), .A2(n9745), .ZN(n9749) );
  NAND2_X1 U10667 ( .A1(n9902), .A2(n9839), .ZN(n9746) );
  AND2_X1 U10668 ( .A1(n9900), .A2(n9746), .ZN(n9755) );
  NAND2_X1 U10669 ( .A1(n9747), .A2(n9755), .ZN(n9748) );
  AOI21_X1 U10670 ( .B1(n9749), .B2(n9748), .A(n5765), .ZN(n9797) );
  INV_X1 U10671 ( .A(n9750), .ZN(n9752) );
  NAND2_X1 U10672 ( .A1(n9752), .A2(n9751), .ZN(n9753) );
  AND2_X1 U10673 ( .A1(n9754), .A2(n9753), .ZN(n9759) );
  INV_X1 U10674 ( .A(n9755), .ZN(n9757) );
  NAND2_X1 U10675 ( .A1(n9757), .A2(n9756), .ZN(n9801) );
  OAI211_X1 U10676 ( .C1(n9759), .C2(n9801), .A(n9817), .B(n9758), .ZN(n9761)
         );
  NAND3_X1 U10677 ( .A1(n9761), .A2(n9760), .A3(n9819), .ZN(n9796) );
  NOR2_X1 U10678 ( .A1(n9762), .A2(n7285), .ZN(n9768) );
  NOR2_X1 U10679 ( .A1(n9764), .A2(n9763), .ZN(n9767) );
  NAND4_X1 U10680 ( .A1(n9768), .A2(n9767), .A3(n9766), .A4(n9765), .ZN(n9770)
         );
  NOR3_X1 U10681 ( .A1(n9770), .A2(n7503), .A3(n9769), .ZN(n9771) );
  NAND4_X1 U10682 ( .A1(n9773), .A2(n9772), .A3(n7562), .A4(n9771), .ZN(n9774)
         );
  NOR2_X1 U10683 ( .A1(n9775), .A2(n9774), .ZN(n9776) );
  NAND3_X1 U10684 ( .A1(n9778), .A2(n9777), .A3(n9776), .ZN(n9779) );
  NOR2_X1 U10685 ( .A1(n9780), .A2(n9779), .ZN(n9781) );
  NAND4_X1 U10686 ( .A1(n10107), .A2(n10127), .A3(n9782), .A4(n9781), .ZN(
        n9783) );
  NOR2_X1 U10687 ( .A1(n10059), .A2(n9783), .ZN(n9784) );
  AND4_X1 U10688 ( .A1(n10023), .A2(n10037), .A3(n10073), .A4(n9784), .ZN(
        n9785) );
  NAND4_X1 U10689 ( .A1(n9980), .A2(n10001), .A3(n9785), .A4(n10007), .ZN(
        n9786) );
  NOR2_X1 U10690 ( .A1(n9970), .A2(n9786), .ZN(n9787) );
  NAND4_X1 U10691 ( .A1(n9919), .A2(n9788), .A3(n9944), .A4(n9787), .ZN(n9789)
         );
  NOR2_X1 U10692 ( .A1(n9790), .A2(n9789), .ZN(n9792) );
  NAND3_X1 U10693 ( .A1(n9819), .A2(n9792), .A3(n9791), .ZN(n9794) );
  OR2_X1 U10694 ( .A1(n9794), .A2(n9793), .ZN(n9795) );
  NAND2_X1 U10695 ( .A1(n9795), .A2(n5762), .ZN(n9824) );
  OAI21_X1 U10696 ( .B1(n9797), .B2(n9796), .A(n9824), .ZN(n9799) );
  MUX2_X1 U10697 ( .A(n9827), .B(n9799), .S(n9798), .Z(n9800) );
  INV_X1 U10698 ( .A(n9800), .ZN(n9826) );
  INV_X1 U10699 ( .A(n9801), .ZN(n9815) );
  AND2_X1 U10700 ( .A1(n9803), .A2(n9802), .ZN(n9805) );
  NOR2_X1 U10701 ( .A1(n9805), .A2(n9804), .ZN(n9806) );
  NOR2_X1 U10702 ( .A1(n9807), .A2(n9806), .ZN(n9808) );
  NOR2_X1 U10703 ( .A1(n9809), .A2(n9808), .ZN(n9813) );
  INV_X1 U10704 ( .A(n9810), .ZN(n9811) );
  OAI21_X1 U10705 ( .B1(n9813), .B2(n9812), .A(n9811), .ZN(n9814) );
  NAND2_X1 U10706 ( .A1(n9815), .A2(n9814), .ZN(n9816) );
  NAND2_X1 U10707 ( .A1(n9817), .A2(n9816), .ZN(n9821) );
  INV_X1 U10708 ( .A(n9818), .ZN(n9820) );
  NAND3_X1 U10709 ( .A1(n9821), .A2(n9820), .A3(n9819), .ZN(n9822) );
  OAI21_X1 U10710 ( .B1(n9824), .B2(n9823), .A(n9822), .ZN(n9825) );
  MUX2_X1 U10711 ( .A(n9826), .B(n9825), .S(n10030), .Z(n9838) );
  INV_X1 U10712 ( .A(n9827), .ZN(n9829) );
  OAI21_X1 U10713 ( .B1(n9829), .B2(n9828), .A(n9832), .ZN(n9837) );
  NAND2_X1 U10714 ( .A1(n9830), .A2(n10746), .ZN(n9834) );
  AOI21_X1 U10715 ( .B1(n5765), .B2(n9832), .A(n9831), .ZN(n9833) );
  OAI21_X1 U10716 ( .B1(n9835), .B2(n9834), .A(n9833), .ZN(n9836) );
  OAI21_X1 U10717 ( .B1(n9838), .B2(n9837), .A(n9836), .ZN(P1_U3240) );
  MUX2_X1 U10718 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9839), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10719 ( .A(n9912), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9852), .Z(
        P1_U3584) );
  MUX2_X1 U10720 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9840), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10721 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9953), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10722 ( .A(n9940), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9852), .Z(
        P1_U3581) );
  MUX2_X1 U10723 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9982), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10724 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n10015), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10725 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n10025), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10726 ( .A(n10068), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9852), .Z(
        P1_U3575) );
  MUX2_X1 U10727 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10040), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10728 ( .A(n10109), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9852), .Z(
        P1_U3571) );
  MUX2_X1 U10729 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n10132), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10730 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9841), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10731 ( .A(n9842), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9852), .Z(
        P1_U3568) );
  MUX2_X1 U10732 ( .A(n9843), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9852), .Z(
        P1_U3567) );
  MUX2_X1 U10733 ( .A(n9844), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9852), .Z(
        P1_U3566) );
  MUX2_X1 U10734 ( .A(n9845), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9852), .Z(
        P1_U3565) );
  MUX2_X1 U10735 ( .A(n9846), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9852), .Z(
        P1_U3564) );
  MUX2_X1 U10736 ( .A(n9847), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9852), .Z(
        P1_U3562) );
  MUX2_X1 U10737 ( .A(n9848), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9852), .Z(
        P1_U3561) );
  MUX2_X1 U10738 ( .A(n9849), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9852), .Z(
        P1_U3560) );
  MUX2_X1 U10739 ( .A(n7246), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9852), .Z(
        P1_U3558) );
  MUX2_X1 U10740 ( .A(n9850), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9852), .Z(
        P1_U3557) );
  MUX2_X1 U10741 ( .A(n9851), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9852), .Z(
        P1_U3556) );
  MUX2_X1 U10742 ( .A(n6891), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9852), .Z(
        P1_U3555) );
  INV_X1 U10743 ( .A(n9853), .ZN(n9858) );
  AOI21_X1 U10744 ( .B1(n9860), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9854), .ZN(
        n9856) );
  XNOR2_X1 U10745 ( .A(n9875), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9855) );
  NOR2_X1 U10746 ( .A1(n9856), .A2(n9855), .ZN(n9874) );
  AOI211_X1 U10747 ( .C1(n9856), .C2(n9855), .A(n9874), .B(n10754), .ZN(n9857)
         );
  AOI211_X1 U10748 ( .C1(n9875), .C2(n10760), .A(n9858), .B(n9857), .ZN(n9866)
         );
  AOI21_X1 U10749 ( .B1(n9860), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9859), .ZN(
        n9863) );
  NAND2_X1 U10750 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9875), .ZN(n9861) );
  OAI21_X1 U10751 ( .B1(n9875), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9861), .ZN(
        n9862) );
  NOR2_X1 U10752 ( .A1(n9863), .A2(n9862), .ZN(n9867) );
  AOI211_X1 U10753 ( .C1(n9863), .C2(n9862), .A(n9867), .B(n9869), .ZN(n9864)
         );
  AOI21_X1 U10754 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(n10761), .A(n9864), .ZN(
        n9865) );
  NAND2_X1 U10755 ( .A1(n9866), .A2(n9865), .ZN(P1_U3258) );
  INV_X1 U10756 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9883) );
  AOI21_X1 U10757 ( .B1(n9875), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9867), .ZN(
        n9871) );
  NAND2_X1 U10758 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n9891), .ZN(n9868) );
  OAI21_X1 U10759 ( .B1(n9891), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9868), .ZN(
        n9870) );
  NOR2_X1 U10760 ( .A1(n9871), .A2(n9870), .ZN(n9886) );
  AOI211_X1 U10761 ( .C1(n9871), .C2(n9870), .A(n9886), .B(n9869), .ZN(n9872)
         );
  AOI21_X1 U10762 ( .B1(n10760), .B2(n9891), .A(n9872), .ZN(n9882) );
  XNOR2_X1 U10763 ( .A(n9873), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9877) );
  AOI21_X1 U10764 ( .B1(n9875), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9874), .ZN(
        n9876) );
  NAND2_X1 U10765 ( .A1(n9876), .A2(n9877), .ZN(n9890) );
  OAI21_X1 U10766 ( .B1(n9877), .B2(n9876), .A(n9890), .ZN(n9880) );
  INV_X1 U10767 ( .A(n9878), .ZN(n9879) );
  AOI21_X1 U10768 ( .B1(n10745), .B2(n9880), .A(n9879), .ZN(n9881) );
  OAI211_X1 U10769 ( .C1(n9884), .C2(n9883), .A(n9882), .B(n9881), .ZN(
        P1_U3259) );
  INV_X1 U10770 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9885) );
  MUX2_X1 U10771 ( .A(n9885), .B(P1_REG2_REG_19__SCAN_IN), .S(n10659), .Z(
        n9888) );
  AOI21_X1 U10772 ( .B1(n9891), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9886), .ZN(
        n9887) );
  XOR2_X1 U10773 ( .A(n9888), .B(n9887), .Z(n9889) );
  AOI22_X1 U10774 ( .A1(n10761), .A2(P1_ADDR_REG_19__SCAN_IN), .B1(n10763), 
        .B2(n9889), .ZN(n9898) );
  OAI21_X1 U10775 ( .B1(n9891), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9890), .ZN(
        n9893) );
  XNOR2_X1 U10776 ( .A(n10030), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9892) );
  XNOR2_X1 U10777 ( .A(n9893), .B(n9892), .ZN(n9896) );
  INV_X1 U10778 ( .A(n9894), .ZN(n9895) );
  AOI21_X1 U10779 ( .B1(n10745), .B2(n9896), .A(n9895), .ZN(n9897) );
  OAI211_X1 U10780 ( .C1(n10030), .C2(n9899), .A(n9898), .B(n9897), .ZN(
        P1_U3260) );
  NAND2_X1 U10781 ( .A1(n9902), .A2(n9901), .ZN(n11017) );
  NOR2_X1 U10782 ( .A1(n10141), .A2(n11017), .ZN(n9907) );
  NOR2_X1 U10783 ( .A1(n10093), .A2(n9903), .ZN(n9904) );
  AOI211_X1 U10784 ( .C1(n10149), .C2(n10095), .A(n9907), .B(n9904), .ZN(n9905) );
  OAI21_X1 U10785 ( .B1(n10150), .B2(n10098), .A(n9905), .ZN(P1_U3261) );
  XNOR2_X1 U10786 ( .A(n11019), .B(n9906), .ZN(n11022) );
  NAND2_X1 U10787 ( .A1(n11022), .A2(n10115), .ZN(n9909) );
  AOI21_X1 U10788 ( .B1(n10141), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9907), .ZN(
        n9908) );
  OAI211_X1 U10789 ( .C1(n11019), .C2(n10144), .A(n9909), .B(n9908), .ZN(
        P1_U3262) );
  OAI21_X1 U10790 ( .B1(n9919), .B2(n9911), .A(n9910), .ZN(n9916) );
  NAND2_X1 U10791 ( .A1(n9912), .A2(n10130), .ZN(n9913) );
  AOI21_X1 U10792 ( .B1(n9919), .B2(n9918), .A(n9917), .ZN(n10157) );
  OR2_X1 U10793 ( .A1(n9920), .A2(n5048), .ZN(n9922) );
  AND2_X1 U10794 ( .A1(n9922), .A2(n9921), .ZN(n10159) );
  NAND2_X1 U10795 ( .A1(n10159), .A2(n10115), .ZN(n9927) );
  OAI22_X1 U10796 ( .A1(n10093), .A2(n9924), .B1(n9923), .B2(n10090), .ZN(
        n9925) );
  AOI21_X1 U10797 ( .B1(n10158), .B2(n10095), .A(n9925), .ZN(n9926) );
  NAND2_X1 U10798 ( .A1(n9927), .A2(n9926), .ZN(n9928) );
  AOI21_X1 U10799 ( .B1(n10157), .B2(n9929), .A(n9928), .ZN(n9930) );
  OAI21_X1 U10800 ( .B1(n10141), .B2(n10161), .A(n9930), .ZN(P1_U3263) );
  XNOR2_X1 U10801 ( .A(n9931), .B(n9937), .ZN(n10167) );
  AOI21_X1 U10802 ( .B1(n10163), .B2(n5310), .A(n5048), .ZN(n10164) );
  AOI22_X1 U10803 ( .A1(n10141), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n10139), 
        .B2(n9932), .ZN(n9933) );
  OAI21_X1 U10804 ( .B1(n5394), .B2(n10144), .A(n9933), .ZN(n9942) );
  NOR2_X1 U10805 ( .A1(n9934), .A2(n10083), .ZN(n9939) );
  AOI211_X1 U10806 ( .C1(n9937), .C2(n9936), .A(n9972), .B(n9935), .ZN(n9938)
         );
  NOR2_X1 U10807 ( .A1(n10166), .A2(n10141), .ZN(n9941) );
  OAI21_X1 U10808 ( .B1(n10148), .B2(n10167), .A(n9943), .ZN(P1_U3264) );
  XNOR2_X1 U10809 ( .A(n9945), .B(n9944), .ZN(n10172) );
  AOI21_X1 U10810 ( .B1(n10168), .B2(n9961), .A(n9946), .ZN(n10169) );
  INV_X1 U10811 ( .A(n9947), .ZN(n9948) );
  AOI22_X1 U10812 ( .A1(n10141), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9948), 
        .B2(n10139), .ZN(n9949) );
  OAI21_X1 U10813 ( .B1(n9950), .B2(n10144), .A(n9949), .ZN(n9956) );
  XNOR2_X1 U10814 ( .A(n9952), .B(n9951), .ZN(n9954) );
  AOI222_X1 U10815 ( .A1(n10125), .A2(n9954), .B1(n9982), .B2(n10131), .C1(
        n9953), .C2(n10130), .ZN(n10171) );
  NOR2_X1 U10816 ( .A1(n10171), .A2(n10141), .ZN(n9955) );
  OAI21_X1 U10817 ( .B1(n10172), .B2(n10148), .A(n9957), .ZN(P1_U3265) );
  OAI21_X1 U10818 ( .B1(n9959), .B2(n9970), .A(n9958), .ZN(n9960) );
  INV_X1 U10819 ( .A(n9960), .ZN(n10177) );
  INV_X1 U10820 ( .A(n9986), .ZN(n9963) );
  INV_X1 U10821 ( .A(n9961), .ZN(n9962) );
  AOI211_X1 U10822 ( .C1(n10175), .C2(n9963), .A(n11009), .B(n9962), .ZN(
        n10174) );
  NOR2_X1 U10823 ( .A1(n9964), .A2(n10144), .ZN(n9968) );
  OAI22_X1 U10824 ( .A1(n10093), .A2(n9966), .B1(n9965), .B2(n10090), .ZN(
        n9967) );
  AOI211_X1 U10825 ( .C1(n10174), .C2(n10138), .A(n9968), .B(n9967), .ZN(n9976) );
  NAND2_X1 U10826 ( .A1(n10173), .A2(n10093), .ZN(n9975) );
  OAI211_X1 U10827 ( .C1(n10177), .C2(n10148), .A(n9976), .B(n9975), .ZN(
        P1_U3266) );
  AOI21_X1 U10828 ( .B1(n9980), .B2(n9978), .A(n9977), .ZN(n9979) );
  INV_X1 U10829 ( .A(n9979), .ZN(n10182) );
  AOI22_X1 U10830 ( .A1(n10179), .A2(n10095), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10141), .ZN(n9991) );
  XNOR2_X1 U10831 ( .A(n9981), .B(n9980), .ZN(n9983) );
  AOI222_X1 U10832 ( .A1(n10125), .A2(n9983), .B1(n10015), .B2(n10131), .C1(
        n9982), .C2(n10130), .ZN(n10181) );
  NAND2_X1 U10833 ( .A1(n10179), .A2(n9993), .ZN(n9984) );
  NAND2_X1 U10834 ( .A1(n9984), .A2(n11021), .ZN(n9985) );
  NOR2_X1 U10835 ( .A1(n9986), .A2(n9985), .ZN(n10178) );
  AOI22_X1 U10836 ( .A1(n10178), .A2(n10030), .B1(n10139), .B2(n9987), .ZN(
        n9988) );
  AOI21_X1 U10837 ( .B1(n10181), .B2(n9988), .A(n10141), .ZN(n9989) );
  INV_X1 U10838 ( .A(n9989), .ZN(n9990) );
  OAI211_X1 U10839 ( .C1(n10182), .C2(n10148), .A(n9991), .B(n9990), .ZN(
        P1_U3267) );
  XNOR2_X1 U10840 ( .A(n9992), .B(n10001), .ZN(n10187) );
  INV_X1 U10841 ( .A(n10009), .ZN(n9995) );
  INV_X1 U10842 ( .A(n9993), .ZN(n9994) );
  AOI211_X1 U10843 ( .C1(n10184), .C2(n9995), .A(n11009), .B(n9994), .ZN(
        n10183) );
  AOI22_X1 U10844 ( .A1(n9996), .A2(n10139), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10141), .ZN(n9997) );
  OAI21_X1 U10845 ( .B1(n9998), .B2(n10144), .A(n9997), .ZN(n10005) );
  OAI21_X1 U10846 ( .B1(n10001), .B2(n10000), .A(n9999), .ZN(n10003) );
  AOI222_X1 U10847 ( .A1(n10125), .A2(n10003), .B1(n10025), .B2(n10131), .C1(
        n10002), .C2(n10130), .ZN(n10186) );
  NOR2_X1 U10848 ( .A1(n10186), .A2(n10141), .ZN(n10004) );
  AOI211_X1 U10849 ( .C1(n10183), .C2(n10138), .A(n10005), .B(n10004), .ZN(
        n10006) );
  OAI21_X1 U10850 ( .B1(n10187), .B2(n10148), .A(n10006), .ZN(P1_U3268) );
  XNOR2_X1 U10851 ( .A(n10008), .B(n10007), .ZN(n10192) );
  AOI21_X1 U10852 ( .B1(n10188), .B2(n10027), .A(n10009), .ZN(n10189) );
  AOI22_X1 U10853 ( .A1(n10010), .A2(n10139), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10141), .ZN(n10011) );
  OAI21_X1 U10854 ( .B1(n10012), .B2(n10144), .A(n10011), .ZN(n10019) );
  XNOR2_X1 U10855 ( .A(n10014), .B(n10013), .ZN(n10017) );
  AOI222_X1 U10856 ( .A1(n10125), .A2(n10017), .B1(n10016), .B2(n10131), .C1(
        n10015), .C2(n10130), .ZN(n10191) );
  NOR2_X1 U10857 ( .A1(n10191), .A2(n10141), .ZN(n10018) );
  AOI211_X1 U10858 ( .C1(n10189), .C2(n10115), .A(n10019), .B(n10018), .ZN(
        n10020) );
  OAI21_X1 U10859 ( .B1(n10192), .B2(n10148), .A(n10020), .ZN(P1_U3269) );
  AOI21_X1 U10860 ( .B1(n10023), .B2(n10021), .A(n5083), .ZN(n10022) );
  INV_X1 U10861 ( .A(n10022), .ZN(n10197) );
  XNOR2_X1 U10862 ( .A(n10024), .B(n10023), .ZN(n10026) );
  AOI222_X1 U10863 ( .A1(n10125), .A2(n10026), .B1(n10025), .B2(n10130), .C1(
        n10068), .C2(n10131), .ZN(n10196) );
  AOI21_X1 U10864 ( .B1(n10048), .B2(n10194), .A(n11009), .ZN(n10028) );
  AND2_X1 U10865 ( .A1(n10028), .A2(n10027), .ZN(n10193) );
  AOI22_X1 U10866 ( .A1(n10193), .A2(n10030), .B1(n10139), .B2(n10029), .ZN(
        n10031) );
  AOI21_X1 U10867 ( .B1(n10196), .B2(n10031), .A(n10141), .ZN(n10032) );
  INV_X1 U10868 ( .A(n10032), .ZN(n10034) );
  AOI22_X1 U10869 ( .A1(n10194), .A2(n10095), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n10141), .ZN(n10033) );
  OAI211_X1 U10870 ( .C1(n10197), .C2(n10148), .A(n10034), .B(n10033), .ZN(
        P1_U3270) );
  OAI21_X1 U10871 ( .B1(n10037), .B2(n10036), .A(n10035), .ZN(n10047) );
  OAI22_X1 U10872 ( .A1(n10038), .A2(n10083), .B1(n10084), .B2(n10081), .ZN(
        n10046) );
  AOI22_X1 U10873 ( .A1(n10039), .A2(n10059), .B1(n10040), .B2(n10203), .ZN(
        n10043) );
  OAI21_X1 U10874 ( .B1(n10043), .B2(n10042), .A(n10041), .ZN(n10044) );
  INV_X1 U10875 ( .A(n10044), .ZN(n10202) );
  NOR2_X1 U10876 ( .A1(n10202), .A2(n7255), .ZN(n10045) );
  AOI211_X1 U10877 ( .C1(n10125), .C2(n10047), .A(n10046), .B(n10045), .ZN(
        n10201) );
  INV_X1 U10878 ( .A(n10061), .ZN(n10050) );
  INV_X1 U10879 ( .A(n10048), .ZN(n10049) );
  AOI21_X1 U10880 ( .B1(n10198), .B2(n10050), .A(n10049), .ZN(n10199) );
  INV_X1 U10881 ( .A(n10051), .ZN(n10052) );
  AOI22_X1 U10882 ( .A1(n10052), .A2(n10139), .B1(n10141), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n10053) );
  OAI21_X1 U10883 ( .B1(n10054), .B2(n10144), .A(n10053), .ZN(n10057) );
  NOR2_X1 U10884 ( .A1(n10202), .A2(n10055), .ZN(n10056) );
  AOI211_X1 U10885 ( .C1(n10199), .C2(n10115), .A(n10057), .B(n10056), .ZN(
        n10058) );
  OAI21_X1 U10886 ( .B1(n10201), .B2(n10141), .A(n10058), .ZN(P1_U3271) );
  XNOR2_X1 U10887 ( .A(n10039), .B(n10059), .ZN(n10207) );
  NOR2_X1 U10888 ( .A1(n10089), .A2(n10064), .ZN(n10060) );
  NOR2_X1 U10889 ( .A1(n10061), .A2(n10060), .ZN(n10204) );
  AOI22_X1 U10890 ( .A1(n10141), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n10062), 
        .B2(n10139), .ZN(n10063) );
  OAI21_X1 U10891 ( .B1(n10064), .B2(n10144), .A(n10063), .ZN(n10071) );
  OAI21_X1 U10892 ( .B1(n10067), .B2(n10066), .A(n10065), .ZN(n10069) );
  AOI222_X1 U10893 ( .A1(n10125), .A2(n10069), .B1(n10068), .B2(n10130), .C1(
        n10110), .C2(n10131), .ZN(n10206) );
  NOR2_X1 U10894 ( .A1(n10206), .A2(n10141), .ZN(n10070) );
  AOI211_X1 U10895 ( .C1(n10204), .C2(n10115), .A(n10071), .B(n10070), .ZN(
        n10072) );
  OAI21_X1 U10896 ( .B1(n10148), .B2(n10207), .A(n10072), .ZN(P1_U3272) );
  NAND2_X1 U10897 ( .A1(n10074), .A2(n10073), .ZN(n10075) );
  NAND2_X1 U10898 ( .A1(n10076), .A2(n10075), .ZN(n10212) );
  NAND2_X1 U10899 ( .A1(n10078), .A2(n10077), .ZN(n10079) );
  NAND2_X1 U10900 ( .A1(n10080), .A2(n10079), .ZN(n10086) );
  OAI22_X1 U10901 ( .A1(n10084), .A2(n10083), .B1(n10082), .B2(n10081), .ZN(
        n10085) );
  AOI21_X1 U10902 ( .B1(n10086), .B2(n10125), .A(n10085), .ZN(n10087) );
  OAI21_X1 U10903 ( .B1(n10212), .B2(n7255), .A(n10087), .ZN(n10214) );
  INV_X1 U10904 ( .A(n10214), .ZN(n10102) );
  INV_X1 U10905 ( .A(n10212), .ZN(n10100) );
  NOR2_X1 U10906 ( .A1(n10114), .A2(n10208), .ZN(n10088) );
  OR2_X1 U10907 ( .A1(n10089), .A2(n10088), .ZN(n10209) );
  INV_X1 U10908 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10092) );
  OAI22_X1 U10909 ( .A1(n10093), .A2(n10092), .B1(n10091), .B2(n10090), .ZN(
        n10094) );
  AOI21_X1 U10910 ( .B1(n10096), .B2(n10095), .A(n10094), .ZN(n10097) );
  OAI21_X1 U10911 ( .B1(n10209), .B2(n10098), .A(n10097), .ZN(n10099) );
  AOI21_X1 U10912 ( .B1(n10100), .B2(n10121), .A(n10099), .ZN(n10101) );
  OAI21_X1 U10913 ( .B1(n10102), .B2(n10141), .A(n10101), .ZN(P1_U3273) );
  OAI21_X1 U10914 ( .B1(n10105), .B2(n10104), .A(n10103), .ZN(n10215) );
  OAI211_X1 U10915 ( .C1(n10108), .C2(n10107), .A(n10106), .B(n10125), .ZN(
        n10112) );
  AOI22_X1 U10916 ( .A1(n10110), .A2(n10130), .B1(n10131), .B2(n10109), .ZN(
        n10111) );
  NAND2_X1 U10917 ( .A1(n10112), .A2(n10111), .ZN(n10113) );
  AOI21_X1 U10918 ( .B1(n10929), .B2(n10215), .A(n10113), .ZN(n10219) );
  AOI21_X1 U10919 ( .B1(n10216), .B2(n10135), .A(n10114), .ZN(n10217) );
  NAND2_X1 U10920 ( .A1(n10217), .A2(n10115), .ZN(n10118) );
  AOI22_X1 U10921 ( .A1(n10141), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10116), 
        .B2(n10139), .ZN(n10117) );
  OAI211_X1 U10922 ( .C1(n10119), .C2(n10144), .A(n10118), .B(n10117), .ZN(
        n10120) );
  AOI21_X1 U10923 ( .B1(n10215), .B2(n10121), .A(n10120), .ZN(n10122) );
  OAI21_X1 U10924 ( .B1(n10219), .B2(n10141), .A(n10122), .ZN(P1_U3274) );
  XNOR2_X1 U10925 ( .A(n10124), .B(n10123), .ZN(n10225) );
  OAI211_X1 U10926 ( .C1(n10128), .C2(n10127), .A(n10126), .B(n10125), .ZN(
        n10134) );
  AOI22_X1 U10927 ( .A1(n10132), .A2(n10131), .B1(n10130), .B2(n10129), .ZN(
        n10133) );
  NAND2_X1 U10928 ( .A1(n10134), .A2(n10133), .ZN(n10221) );
  INV_X1 U10929 ( .A(n10135), .ZN(n10136) );
  AOI211_X1 U10930 ( .C1(n10223), .C2(n10137), .A(n11009), .B(n10136), .ZN(
        n10222) );
  NAND2_X1 U10931 ( .A1(n10222), .A2(n10138), .ZN(n10143) );
  AOI22_X1 U10932 ( .A1(n10141), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n10140), 
        .B2(n10139), .ZN(n10142) );
  OAI211_X1 U10933 ( .C1(n10145), .C2(n10144), .A(n10143), .B(n10142), .ZN(
        n10146) );
  AOI21_X1 U10934 ( .B1(n10221), .B2(n10093), .A(n10146), .ZN(n10147) );
  OAI21_X1 U10935 ( .B1(n10148), .B2(n10225), .A(n10147), .ZN(P1_U3275) );
  AOI21_X1 U10936 ( .B1(n10946), .B2(n10152), .A(n10151), .ZN(n10153) );
  OAI21_X1 U10937 ( .B1(n10156), .B2(n10232), .A(n10155), .ZN(n10241) );
  MUX2_X1 U10938 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10241), .S(n11024), .Z(
        P1_U3552) );
  INV_X1 U10939 ( .A(n10157), .ZN(n10162) );
  AOI22_X1 U10940 ( .A1(n10159), .A2(n11021), .B1(n10946), .B2(n10158), .ZN(
        n10160) );
  OAI211_X1 U10941 ( .C1(n10162), .C2(n10232), .A(n10161), .B(n10160), .ZN(
        n10242) );
  MUX2_X1 U10942 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10242), .S(n11024), .Z(
        P1_U3551) );
  AOI22_X1 U10943 ( .A1(n10164), .A2(n11021), .B1(n10946), .B2(n10163), .ZN(
        n10165) );
  OAI211_X1 U10944 ( .C1(n10232), .C2(n10167), .A(n10166), .B(n10165), .ZN(
        n10243) );
  MUX2_X1 U10945 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10243), .S(n11024), .Z(
        P1_U3550) );
  AOI22_X1 U10946 ( .A1(n10169), .A2(n11021), .B1(n10946), .B2(n10168), .ZN(
        n10170) );
  OAI211_X1 U10947 ( .C1(n10172), .C2(n10232), .A(n10171), .B(n10170), .ZN(
        n10244) );
  MUX2_X1 U10948 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10244), .S(n11024), .Z(
        P1_U3549) );
  AOI211_X1 U10949 ( .C1(n10946), .C2(n10175), .A(n10174), .B(n10173), .ZN(
        n10176) );
  OAI21_X1 U10950 ( .B1(n10232), .B2(n10177), .A(n10176), .ZN(n10245) );
  MUX2_X1 U10951 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10245), .S(n11024), .Z(
        P1_U3548) );
  AOI21_X1 U10952 ( .B1(n10946), .B2(n10179), .A(n10178), .ZN(n10180) );
  OAI211_X1 U10953 ( .C1(n10182), .C2(n10232), .A(n10181), .B(n10180), .ZN(
        n10246) );
  MUX2_X1 U10954 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10246), .S(n11024), .Z(
        P1_U3547) );
  AOI21_X1 U10955 ( .B1(n10946), .B2(n10184), .A(n10183), .ZN(n10185) );
  OAI211_X1 U10956 ( .C1(n10187), .C2(n10232), .A(n10186), .B(n10185), .ZN(
        n10247) );
  MUX2_X1 U10957 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10247), .S(n11024), .Z(
        P1_U3546) );
  AOI22_X1 U10958 ( .A1(n10189), .A2(n11021), .B1(n10946), .B2(n10188), .ZN(
        n10190) );
  OAI211_X1 U10959 ( .C1(n10192), .C2(n10232), .A(n10191), .B(n10190), .ZN(
        n10248) );
  MUX2_X1 U10960 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10248), .S(n11024), .Z(
        P1_U3545) );
  AOI21_X1 U10961 ( .B1(n10946), .B2(n10194), .A(n10193), .ZN(n10195) );
  OAI211_X1 U10962 ( .C1(n10197), .C2(n10232), .A(n10196), .B(n10195), .ZN(
        n10249) );
  MUX2_X1 U10963 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10249), .S(n11024), .Z(
        P1_U3544) );
  AOI22_X1 U10964 ( .A1(n10199), .A2(n11021), .B1(n10946), .B2(n10198), .ZN(
        n10200) );
  OAI211_X1 U10965 ( .C1(n10202), .C2(n10923), .A(n10201), .B(n10200), .ZN(
        n10250) );
  MUX2_X1 U10966 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10250), .S(n11024), .Z(
        P1_U3543) );
  AOI22_X1 U10967 ( .A1(n10204), .A2(n11021), .B1(n10946), .B2(n10203), .ZN(
        n10205) );
  OAI211_X1 U10968 ( .C1(n10232), .C2(n10207), .A(n10206), .B(n10205), .ZN(
        n10251) );
  MUX2_X1 U10969 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10251), .S(n11024), .Z(
        P1_U3542) );
  OAI22_X1 U10970 ( .A1(n10209), .A2(n11009), .B1(n10208), .B2(n11018), .ZN(
        n10210) );
  INV_X1 U10971 ( .A(n10210), .ZN(n10211) );
  OAI21_X1 U10972 ( .B1(n10212), .B2(n10923), .A(n10211), .ZN(n10213) );
  OR2_X1 U10973 ( .A1(n10214), .A2(n10213), .ZN(n10252) );
  MUX2_X1 U10974 ( .A(n10252), .B(P1_REG1_REG_18__SCAN_IN), .S(n11023), .Z(
        P1_U3541) );
  INV_X1 U10975 ( .A(n10215), .ZN(n10220) );
  AOI22_X1 U10976 ( .A1(n10217), .A2(n11021), .B1(n10946), .B2(n10216), .ZN(
        n10218) );
  OAI211_X1 U10977 ( .C1(n10220), .C2(n10923), .A(n10219), .B(n10218), .ZN(
        n10253) );
  MUX2_X1 U10978 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10253), .S(n11024), .Z(
        P1_U3540) );
  AOI211_X1 U10979 ( .C1(n10946), .C2(n10223), .A(n10222), .B(n10221), .ZN(
        n10224) );
  OAI21_X1 U10980 ( .B1(n10232), .B2(n10225), .A(n10224), .ZN(n10254) );
  MUX2_X1 U10981 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10254), .S(n11024), .Z(
        P1_U3539) );
  INV_X1 U10982 ( .A(n10226), .ZN(n10231) );
  AOI21_X1 U10983 ( .B1(n10946), .B2(n10228), .A(n10227), .ZN(n10229) );
  OAI211_X1 U10984 ( .C1(n10231), .C2(n10232), .A(n10230), .B(n10229), .ZN(
        n10255) );
  MUX2_X1 U10985 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10255), .S(n11024), .Z(
        P1_U3537) );
  INV_X1 U10986 ( .A(n10232), .ZN(n10948) );
  NAND2_X1 U10987 ( .A1(n10233), .A2(n10946), .ZN(n10234) );
  NAND2_X1 U10988 ( .A1(n10235), .A2(n10234), .ZN(n10236) );
  AOI21_X1 U10989 ( .B1(n10237), .B2(n10948), .A(n10236), .ZN(n10238) );
  NAND2_X1 U10990 ( .A1(n10239), .A2(n10238), .ZN(n10256) );
  MUX2_X1 U10991 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10256), .S(n11024), .Z(
        P1_U3535) );
  MUX2_X1 U10992 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10240), .S(n11028), .Z(
        P1_U3522) );
  MUX2_X1 U10993 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10241), .S(n11028), .Z(
        P1_U3520) );
  MUX2_X1 U10994 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10242), .S(n11028), .Z(
        P1_U3519) );
  MUX2_X1 U10995 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10243), .S(n11028), .Z(
        P1_U3518) );
  MUX2_X1 U10996 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10244), .S(n11028), .Z(
        P1_U3517) );
  MUX2_X1 U10997 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10245), .S(n11028), .Z(
        P1_U3516) );
  MUX2_X1 U10998 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10246), .S(n11028), .Z(
        P1_U3515) );
  MUX2_X1 U10999 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10247), .S(n11028), .Z(
        P1_U3514) );
  MUX2_X1 U11000 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10248), .S(n11028), .Z(
        P1_U3513) );
  MUX2_X1 U11001 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10249), .S(n11028), .Z(
        P1_U3512) );
  MUX2_X1 U11002 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10250), .S(n11028), .Z(
        P1_U3511) );
  MUX2_X1 U11003 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10251), .S(n11028), .Z(
        P1_U3510) );
  MUX2_X1 U11004 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10252), .S(n11028), .Z(
        P1_U3508) );
  MUX2_X1 U11005 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10253), .S(n11028), .Z(
        P1_U3505) );
  MUX2_X1 U11006 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10254), .S(n11028), .Z(
        P1_U3502) );
  MUX2_X1 U11007 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10255), .S(n11028), .Z(
        P1_U3496) );
  MUX2_X1 U11008 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n10256), .S(n11028), .Z(
        P1_U3490) );
  MUX2_X1 U11009 ( .A(P1_D_REG_1__SCAN_IN), .B(n10258), .S(n10257), .Z(
        P1_U3441) );
  MUX2_X1 U11010 ( .A(n10259), .B(P1_D_REG_0__SCAN_IN), .S(n10666), .Z(
        P1_U3440) );
  INV_X1 U11011 ( .A(n10260), .ZN(n10266) );
  NOR4_X1 U11012 ( .A1(n10262), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), 
        .A4(n10261), .ZN(n10263) );
  AOI21_X1 U11013 ( .B1(n10658), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10263), 
        .ZN(n10264) );
  OAI21_X1 U11014 ( .B1(n10266), .B2(n10265), .A(n10264), .ZN(P1_U3322) );
  INV_X1 U11015 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10286) );
  OAI222_X1 U11016 ( .A1(P1_U3084), .A2(n10269), .B1(n10265), .B2(n10268), 
        .C1(n10286), .C2(n10267), .ZN(P1_U3324) );
  INV_X1 U11017 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10668) );
  INV_X1 U11018 ( .A(keyinput_113), .ZN(n10425) );
  OAI22_X1 U11019 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput_93), .B1(
        keyinput_88), .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n10270) );
  AOI221_X1 U11020 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput_93), .C1(
        P2_DATAO_REG_8__SCAN_IN), .C2(keyinput_88), .A(n10270), .ZN(n10390) );
  OAI22_X1 U11021 ( .A1(n10272), .A2(keyinput_87), .B1(keyinput_89), .B2(
        P2_DATAO_REG_7__SCAN_IN), .ZN(n10271) );
  AOI221_X1 U11022 ( .B1(n10272), .B2(keyinput_87), .C1(
        P2_DATAO_REG_7__SCAN_IN), .C2(keyinput_89), .A(n10271), .ZN(n10276) );
  INV_X1 U11023 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n10274) );
  OAI22_X1 U11024 ( .A1(n10274), .A2(keyinput_92), .B1(n10584), .B2(
        keyinput_90), .ZN(n10273) );
  AOI221_X1 U11025 ( .B1(n10274), .B2(keyinput_92), .C1(keyinput_90), .C2(
        n10584), .A(n10273), .ZN(n10275) );
  OAI211_X1 U11026 ( .C1(n10753), .C2(keyinput_91), .A(n10276), .B(n10275), 
        .ZN(n10277) );
  AOI21_X1 U11027 ( .B1(n10753), .B2(keyinput_91), .A(n10277), .ZN(n10389) );
  OAI22_X1 U11028 ( .A1(n10279), .A2(keyinput_85), .B1(keyinput_84), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n10278) );
  AOI221_X1 U11029 ( .B1(n10279), .B2(keyinput_85), .C1(
        P2_DATAO_REG_12__SCAN_IN), .C2(keyinput_84), .A(n10278), .ZN(n10388)
         );
  OAI22_X1 U11030 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(keyinput_78), .B1(
        keyinput_80), .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n10280) );
  AOI221_X1 U11031 ( .B1(P2_DATAO_REG_18__SCAN_IN), .B2(keyinput_78), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput_80), .A(n10280), .ZN(n10386)
         );
  OAI22_X1 U11032 ( .A1(n10573), .A2(keyinput_82), .B1(keyinput_81), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n10281) );
  AOI221_X1 U11033 ( .B1(n10573), .B2(keyinput_82), .C1(
        P2_DATAO_REG_15__SCAN_IN), .C2(keyinput_81), .A(n10281), .ZN(n10385)
         );
  OAI22_X1 U11034 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(keyinput_79), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_83), .ZN(n10282) );
  AOI221_X1 U11035 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_79), .C1(
        keyinput_83), .C2(P2_DATAO_REG_13__SCAN_IN), .A(n10282), .ZN(n10384)
         );
  INV_X1 U11036 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U11037 ( .A1(n10547), .A2(keyinput_64), .B1(n10284), .B2(
        keyinput_68), .ZN(n10283) );
  OAI221_X1 U11038 ( .B1(n10547), .B2(keyinput_64), .C1(n10284), .C2(
        keyinput_68), .A(n10283), .ZN(n10374) );
  AOI22_X1 U11039 ( .A1(n10287), .A2(keyinput_65), .B1(n10286), .B2(
        keyinput_67), .ZN(n10285) );
  OAI221_X1 U11040 ( .B1(n10287), .B2(keyinput_65), .C1(n10286), .C2(
        keyinput_67), .A(n10285), .ZN(n10373) );
  AOI22_X1 U11041 ( .A1(n8305), .A2(keyinput_62), .B1(n10545), .B2(keyinput_63), .ZN(n10288) );
  OAI221_X1 U11042 ( .B1(n8305), .B2(keyinput_62), .C1(n10545), .C2(
        keyinput_63), .A(n10288), .ZN(n10372) );
  AOI22_X1 U11043 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_56), .B1(n10450), .B2(keyinput_53), .ZN(n10289) );
  OAI221_X1 U11044 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_56), .C1(
        n10450), .C2(keyinput_53), .A(n10289), .ZN(n10298) );
  AOI22_X1 U11045 ( .A1(n10292), .A2(keyinput_52), .B1(keyinput_57), .B2(
        n10291), .ZN(n10290) );
  OAI221_X1 U11046 ( .B1(n10292), .B2(keyinput_52), .C1(n10291), .C2(
        keyinput_57), .A(n10290), .ZN(n10297) );
  AOI22_X1 U11047 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_54), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(keyinput_59), .ZN(n10293) );
  OAI221_X1 U11048 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_54), .C1(
        P2_REG3_REG_2__SCAN_IN), .C2(keyinput_59), .A(n10293), .ZN(n10296) );
  AOI22_X1 U11049 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_55), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_58), .ZN(n10294) );
  OAI221_X1 U11050 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_55), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_58), .A(n10294), .ZN(n10295) );
  NOR4_X1 U11051 ( .A1(n10298), .A2(n10297), .A3(n10296), .A4(n10295), .ZN(
        n10369) );
  AOI22_X1 U11052 ( .A1(n10459), .A2(keyinput_49), .B1(keyinput_48), .B2(
        n10300), .ZN(n10299) );
  OAI221_X1 U11053 ( .B1(n10459), .B2(keyinput_49), .C1(n10300), .C2(
        keyinput_48), .A(n10299), .ZN(n10365) );
  OAI22_X1 U11054 ( .A1(n10302), .A2(keyinput_46), .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_47), .ZN(n10301) );
  AOI221_X1 U11055 ( .B1(n10302), .B2(keyinput_46), .C1(keyinput_47), .C2(
        P2_REG3_REG_25__SCAN_IN), .A(n10301), .ZN(n10364) );
  AOI22_X1 U11056 ( .A1(n10785), .A2(keyinput_44), .B1(n7592), .B2(keyinput_43), .ZN(n10303) );
  OAI221_X1 U11057 ( .B1(n10785), .B2(keyinput_44), .C1(n7592), .C2(
        keyinput_43), .A(n10303), .ZN(n10359) );
  INV_X1 U11058 ( .A(keyinput_37), .ZN(n10351) );
  INV_X1 U11059 ( .A(keyinput_36), .ZN(n10350) );
  OAI22_X1 U11060 ( .A1(n10305), .A2(keyinput_32), .B1(P2_RD_REG_SCAN_IN), 
        .B2(keyinput_33), .ZN(n10304) );
  AOI221_X1 U11061 ( .B1(n10305), .B2(keyinput_32), .C1(keyinput_33), .C2(
        P2_RD_REG_SCAN_IN), .A(n10304), .ZN(n10349) );
  INV_X1 U11062 ( .A(SI_1_), .ZN(n10511) );
  INV_X1 U11063 ( .A(keyinput_31), .ZN(n10345) );
  OAI22_X1 U11064 ( .A1(n10307), .A2(keyinput_28), .B1(keyinput_29), .B2(SI_3_), .ZN(n10306) );
  AOI221_X1 U11065 ( .B1(n10307), .B2(keyinput_28), .C1(SI_3_), .C2(
        keyinput_29), .A(n10306), .ZN(n10342) );
  INV_X1 U11066 ( .A(keyinput_22), .ZN(n10336) );
  INV_X1 U11067 ( .A(keyinput_13), .ZN(n10324) );
  INV_X1 U11068 ( .A(keyinput_12), .ZN(n10323) );
  INV_X1 U11069 ( .A(keyinput_11), .ZN(n10322) );
  AOI22_X1 U11070 ( .A1(n10471), .A2(keyinput_8), .B1(n10309), .B2(keyinput_6), 
        .ZN(n10308) );
  OAI221_X1 U11071 ( .B1(n10471), .B2(keyinput_8), .C1(n10309), .C2(keyinput_6), .A(n10308), .ZN(n10313) );
  AOI22_X1 U11072 ( .A1(SI_23_), .A2(keyinput_9), .B1(n10311), .B2(keyinput_7), 
        .ZN(n10310) );
  OAI221_X1 U11073 ( .B1(SI_23_), .B2(keyinput_9), .C1(n10311), .C2(keyinput_7), .A(n10310), .ZN(n10312) );
  AOI211_X1 U11074 ( .C1(keyinput_5), .C2(SI_27_), .A(n10313), .B(n10312), 
        .ZN(n10314) );
  OAI21_X1 U11075 ( .B1(keyinput_5), .B2(SI_27_), .A(n10314), .ZN(n10320) );
  OAI22_X1 U11076 ( .A1(SI_31_), .A2(keyinput_1), .B1(keyinput_0), .B2(
        P2_WR_REG_SCAN_IN), .ZN(n10315) );
  AOI221_X1 U11077 ( .B1(SI_31_), .B2(keyinput_1), .C1(P2_WR_REG_SCAN_IN), 
        .C2(keyinput_0), .A(n10315), .ZN(n10318) );
  AOI211_X1 U11078 ( .C1(n10479), .C2(keyinput_4), .A(n10318), .B(n10317), 
        .ZN(n10319) );
  OAI22_X1 U11079 ( .A1(n10320), .A2(n10319), .B1(keyinput_10), .B2(SI_22_), 
        .ZN(n10321) );
  INV_X1 U11080 ( .A(SI_17_), .ZN(n10326) );
  INV_X1 U11081 ( .A(SI_18_), .ZN(n10469) );
  AOI22_X1 U11082 ( .A1(n10326), .A2(keyinput_15), .B1(n10469), .B2(
        keyinput_14), .ZN(n10325) );
  OAI221_X1 U11083 ( .B1(n10326), .B2(keyinput_15), .C1(n10469), .C2(
        keyinput_14), .A(n10325), .ZN(n10330) );
  XOR2_X1 U11084 ( .A(SI_16_), .B(keyinput_16), .Z(n10329) );
  OAI22_X1 U11085 ( .A1(SI_15_), .A2(keyinput_17), .B1(keyinput_18), .B2(
        SI_14_), .ZN(n10327) );
  AOI221_X1 U11086 ( .B1(SI_15_), .B2(keyinput_17), .C1(SI_14_), .C2(
        keyinput_18), .A(n10327), .ZN(n10328) );
  OAI211_X1 U11087 ( .C1(n10331), .C2(n10330), .A(n10329), .B(n10328), .ZN(
        n10335) );
  OAI22_X1 U11088 ( .A1(SI_13_), .A2(keyinput_19), .B1(keyinput_20), .B2(
        SI_12_), .ZN(n10332) );
  AOI221_X1 U11089 ( .B1(SI_13_), .B2(keyinput_19), .C1(SI_12_), .C2(
        keyinput_20), .A(n10332), .ZN(n10334) );
  INV_X1 U11090 ( .A(SI_11_), .ZN(n10497) );
  NOR2_X1 U11091 ( .A1(n10497), .A2(keyinput_21), .ZN(n10333) );
  INV_X1 U11092 ( .A(SI_8_), .ZN(n10501) );
  OAI22_X1 U11093 ( .A1(n10501), .A2(keyinput_24), .B1(n10338), .B2(
        keyinput_26), .ZN(n10337) );
  AOI221_X1 U11094 ( .B1(n10501), .B2(keyinput_24), .C1(keyinput_26), .C2(
        n10338), .A(n10337), .ZN(n10341) );
  OAI22_X1 U11095 ( .A1(SI_7_), .A2(keyinput_25), .B1(SI_5_), .B2(keyinput_27), 
        .ZN(n10339) );
  AOI221_X1 U11096 ( .B1(SI_7_), .B2(keyinput_25), .C1(keyinput_27), .C2(SI_5_), .A(n10339), .ZN(n10340) );
  OAI21_X1 U11097 ( .B1(keyinput_30), .B2(SI_2_), .A(n10343), .ZN(n10344) );
  OAI221_X1 U11098 ( .B1(SI_1_), .B2(keyinput_31), .C1(n10511), .C2(n10345), 
        .A(n10344), .ZN(n10348) );
  AOI22_X1 U11099 ( .A1(n10514), .A2(keyinput_35), .B1(keyinput_34), .B2(
        P2_U3152), .ZN(n10346) );
  OAI221_X1 U11100 ( .B1(n10514), .B2(keyinput_35), .C1(P2_U3152), .C2(
        keyinput_34), .A(n10346), .ZN(n10347) );
  AOI22_X1 U11101 ( .A1(n10524), .A2(keyinput_41), .B1(keyinput_42), .B2(n8573), .ZN(n10352) );
  OAI221_X1 U11102 ( .B1(n10524), .B2(keyinput_41), .C1(n8573), .C2(
        keyinput_42), .A(n10352), .ZN(n10355) );
  AOI22_X1 U11103 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_40), .B1(n8280), 
        .B2(keyinput_38), .ZN(n10353) );
  OAI221_X1 U11104 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_40), .C1(n8280), 
        .C2(keyinput_38), .A(n10353), .ZN(n10354) );
  NAND2_X1 U11105 ( .A1(n10357), .A2(keyinput_45), .ZN(n10356) );
  OAI221_X1 U11106 ( .B1(n10359), .B2(n10358), .C1(n10357), .C2(keyinput_45), 
        .A(n10356), .ZN(n10363) );
  OAI22_X1 U11107 ( .A1(n10361), .A2(keyinput_50), .B1(keyinput_51), .B2(
        P2_REG3_REG_24__SCAN_IN), .ZN(n10360) );
  AOI221_X1 U11108 ( .B1(n10361), .B2(keyinput_50), .C1(
        P2_REG3_REG_24__SCAN_IN), .C2(keyinput_51), .A(n10360), .ZN(n10362) );
  OAI221_X1 U11109 ( .B1(n10365), .B2(n10364), .C1(n10365), .C2(n10363), .A(
        n10362), .ZN(n10368) );
  AOI22_X1 U11110 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_60), .B1(
        P2_REG3_REG_6__SCAN_IN), .B2(keyinput_61), .ZN(n10366) );
  OAI221_X1 U11111 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_60), .C1(
        P2_REG3_REG_6__SCAN_IN), .C2(keyinput_61), .A(n10366), .ZN(n10367) );
  AOI21_X1 U11112 ( .B1(n10369), .B2(n10368), .A(n10367), .ZN(n10371) );
  NAND2_X1 U11113 ( .A1(keyinput_66), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(
        n10370) );
  AOI22_X1 U11114 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(keyinput_69), .B1(
        n10445), .B2(keyinput_70), .ZN(n10375) );
  OAI221_X1 U11115 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_69), .C1(
        n10445), .C2(keyinput_70), .A(n10375), .ZN(n10380) );
  OAI22_X1 U11116 ( .A1(n10557), .A2(keyinput_75), .B1(keyinput_72), .B2(
        P2_DATAO_REG_24__SCAN_IN), .ZN(n10376) );
  AOI221_X1 U11117 ( .B1(n10557), .B2(keyinput_75), .C1(
        P2_DATAO_REG_24__SCAN_IN), .C2(keyinput_72), .A(n10376), .ZN(n10379)
         );
  OAI22_X1 U11118 ( .A1(n6283), .A2(keyinput_73), .B1(P2_DATAO_REG_22__SCAN_IN), .B2(keyinput_74), .ZN(n10377) );
  AOI221_X1 U11119 ( .B1(n6283), .B2(keyinput_73), .C1(keyinput_74), .C2(
        P2_DATAO_REG_22__SCAN_IN), .A(n10377), .ZN(n10378) );
  OAI22_X1 U11120 ( .A1(n10562), .A2(keyinput_76), .B1(keyinput_77), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n10381) );
  AOI221_X1 U11121 ( .B1(n10562), .B2(keyinput_76), .C1(
        P2_DATAO_REG_19__SCAN_IN), .C2(keyinput_77), .A(n10381), .ZN(n10382)
         );
  NAND4_X1 U11122 ( .A1(n10386), .A2(n10385), .A3(n10384), .A4(n10383), .ZN(
        n10387) );
  XOR2_X1 U11123 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_94), .Z(n10392) );
  XNOR2_X1 U11124 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_95), .ZN(n10391) );
  XNOR2_X1 U11125 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_96), .ZN(n10393) );
  NAND2_X1 U11126 ( .A1(n10394), .A2(n10393), .ZN(n10400) );
  INV_X1 U11127 ( .A(keyinput_97), .ZN(n10395) );
  MUX2_X1 U11128 ( .A(keyinput_97), .B(n10395), .S(P1_IR_REG_6__SCAN_IN), .Z(
        n10399) );
  XNOR2_X1 U11129 ( .A(n10396), .B(keyinput_98), .ZN(n10398) );
  XNOR2_X1 U11130 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_99), .ZN(n10397) );
  AOI211_X1 U11131 ( .C1(n10400), .C2(n10399), .A(n10398), .B(n10397), .ZN(
        n10404) );
  XNOR2_X1 U11132 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_100), .ZN(n10403) );
  INV_X1 U11133 ( .A(keyinput_101), .ZN(n10401) );
  MUX2_X1 U11134 ( .A(n10401), .B(keyinput_101), .S(P1_IR_REG_10__SCAN_IN), 
        .Z(n10402) );
  OAI21_X1 U11135 ( .B1(n10404), .B2(n10403), .A(n10402), .ZN(n10410) );
  INV_X1 U11136 ( .A(keyinput_102), .ZN(n10405) );
  MUX2_X1 U11137 ( .A(keyinput_102), .B(n10405), .S(P1_IR_REG_11__SCAN_IN), 
        .Z(n10409) );
  OAI22_X1 U11138 ( .A1(n10608), .A2(keyinput_104), .B1(keyinput_103), .B2(
        P1_IR_REG_12__SCAN_IN), .ZN(n10406) );
  AOI221_X1 U11139 ( .B1(n10608), .B2(keyinput_104), .C1(P1_IR_REG_12__SCAN_IN), .C2(keyinput_103), .A(n10406), .ZN(n10407) );
  INV_X1 U11140 ( .A(n10407), .ZN(n10408) );
  AOI21_X1 U11141 ( .B1(n10410), .B2(n10409), .A(n10408), .ZN(n10414) );
  XNOR2_X1 U11142 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_105), .ZN(n10413)
         );
  INV_X1 U11143 ( .A(keyinput_106), .ZN(n10411) );
  MUX2_X1 U11144 ( .A(keyinput_106), .B(n10411), .S(P1_IR_REG_15__SCAN_IN), 
        .Z(n10412) );
  OAI21_X1 U11145 ( .B1(n10414), .B2(n10413), .A(n10412), .ZN(n10419) );
  XNOR2_X1 U11146 ( .A(n10415), .B(keyinput_108), .ZN(n10418) );
  OAI22_X1 U11147 ( .A1(n10618), .A2(keyinput_109), .B1(keyinput_107), .B2(
        P1_IR_REG_16__SCAN_IN), .ZN(n10416) );
  AOI221_X1 U11148 ( .B1(n10618), .B2(keyinput_109), .C1(P1_IR_REG_16__SCAN_IN), .C2(keyinput_107), .A(n10416), .ZN(n10417) );
  NAND3_X1 U11149 ( .A1(n10419), .A2(n10418), .A3(n10417), .ZN(n10423) );
  XNOR2_X1 U11150 ( .A(n10420), .B(keyinput_111), .ZN(n10422) );
  XNOR2_X1 U11151 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_110), .ZN(n10421)
         );
  NAND3_X1 U11152 ( .A1(n10423), .A2(n10422), .A3(n10421), .ZN(n10424) );
  XNOR2_X1 U11153 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_114), .ZN(n10427)
         );
  XNOR2_X1 U11154 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_116), .ZN(n10426)
         );
  XNOR2_X1 U11155 ( .A(n10633), .B(keyinput_119), .ZN(n10430) );
  XNOR2_X1 U11156 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_117), .ZN(n10429)
         );
  XNOR2_X1 U11157 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_118), .ZN(n10428)
         );
  NOR4_X1 U11158 ( .A1(n10431), .A2(n10430), .A3(n10429), .A4(n10428), .ZN(
        n10434) );
  INV_X1 U11159 ( .A(keyinput_120), .ZN(n10432) );
  MUX2_X1 U11160 ( .A(keyinput_120), .B(n10432), .S(P1_IR_REG_29__SCAN_IN), 
        .Z(n10433) );
  NOR2_X1 U11161 ( .A1(n10434), .A2(n10433), .ZN(n10439) );
  INV_X1 U11162 ( .A(keyinput_121), .ZN(n10435) );
  MUX2_X1 U11163 ( .A(keyinput_121), .B(n10435), .S(P1_IR_REG_30__SCAN_IN), 
        .Z(n10438) );
  XNOR2_X1 U11164 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_123), .ZN(n10437) );
  XNOR2_X1 U11165 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_122), .ZN(n10436)
         );
  OAI22_X1 U11166 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput_125), .B1(
        keyinput_124), .B2(P1_D_REG_1__SCAN_IN), .ZN(n10440) );
  AOI221_X1 U11167 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput_125), .C1(
        P1_D_REG_1__SCAN_IN), .C2(keyinput_124), .A(n10440), .ZN(n10657) );
  INV_X1 U11168 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10669) );
  INV_X1 U11169 ( .A(keyinput_241), .ZN(n10629) );
  AOI22_X1 U11170 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput_213), .B1(
        n10442), .B2(keyinput_212), .ZN(n10441) );
  OAI221_X1 U11171 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_213), .C1(
        n10442), .C2(keyinput_212), .A(n10441), .ZN(n10580) );
  XNOR2_X1 U11172 ( .A(n10443), .B(keyinput_199), .ZN(n10566) );
  OAI22_X1 U11173 ( .A1(n10446), .A2(keyinput_197), .B1(n10445), .B2(
        keyinput_198), .ZN(n10444) );
  AOI221_X1 U11174 ( .B1(n10446), .B2(keyinput_197), .C1(keyinput_198), .C2(
        n10445), .A(n10444), .ZN(n10560) );
  AOI22_X1 U11175 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_184), .B1(
        n10448), .B2(keyinput_186), .ZN(n10447) );
  OAI221_X1 U11176 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_184), .C1(
        n10448), .C2(keyinput_186), .A(n10447), .ZN(n10457) );
  AOI22_X1 U11177 ( .A1(n10451), .A2(keyinput_187), .B1(n10450), .B2(
        keyinput_181), .ZN(n10449) );
  OAI221_X1 U11178 ( .B1(n10451), .B2(keyinput_187), .C1(n10450), .C2(
        keyinput_181), .A(n10449), .ZN(n10456) );
  AOI22_X1 U11179 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_185), .B1(
        P2_REG3_REG_4__SCAN_IN), .B2(keyinput_180), .ZN(n10452) );
  OAI221_X1 U11180 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_185), .C1(
        P2_REG3_REG_4__SCAN_IN), .C2(keyinput_180), .A(n10452), .ZN(n10455) );
  AOI22_X1 U11181 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_182), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput_183), .ZN(n10453) );
  OAI221_X1 U11182 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_182), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_183), .A(n10453), .ZN(n10454)
         );
  NOR4_X1 U11183 ( .A1(n10457), .A2(n10456), .A3(n10455), .A4(n10454), .ZN(
        n10543) );
  AOI22_X1 U11184 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_176), .B1(
        n10459), .B2(keyinput_177), .ZN(n10458) );
  OAI221_X1 U11185 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_176), .C1(
        n10459), .C2(keyinput_177), .A(n10458), .ZN(n10537) );
  OAI22_X1 U11186 ( .A1(n10461), .A2(keyinput_175), .B1(
        P2_REG3_REG_12__SCAN_IN), .B2(keyinput_174), .ZN(n10460) );
  AOI221_X1 U11187 ( .B1(n10461), .B2(keyinput_175), .C1(keyinput_174), .C2(
        P2_REG3_REG_12__SCAN_IN), .A(n10460), .ZN(n10536) );
  AOI22_X1 U11188 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_172), .B1(n7592), 
        .B2(keyinput_171), .ZN(n10462) );
  OAI221_X1 U11189 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_172), .C1(n7592), .C2(keyinput_171), .A(n10462), .ZN(n10532) );
  INV_X1 U11190 ( .A(keyinput_165), .ZN(n10522) );
  INV_X1 U11191 ( .A(keyinput_164), .ZN(n10519) );
  OAI22_X1 U11192 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_161), .B1(
        keyinput_160), .B2(SI_0_), .ZN(n10463) );
  AOI221_X1 U11193 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_161), .C1(SI_0_), 
        .C2(keyinput_160), .A(n10463), .ZN(n10518) );
  INV_X1 U11194 ( .A(keyinput_159), .ZN(n10512) );
  OAI22_X1 U11195 ( .A1(SI_4_), .A2(keyinput_156), .B1(SI_3_), .B2(
        keyinput_157), .ZN(n10464) );
  AOI221_X1 U11196 ( .B1(SI_4_), .B2(keyinput_156), .C1(keyinput_157), .C2(
        SI_3_), .A(n10464), .ZN(n10508) );
  INV_X1 U11197 ( .A(keyinput_150), .ZN(n10499) );
  AOI22_X1 U11198 ( .A1(n10467), .A2(keyinput_148), .B1(n10466), .B2(
        keyinput_147), .ZN(n10465) );
  OAI221_X1 U11199 ( .B1(n10467), .B2(keyinput_148), .C1(n10466), .C2(
        keyinput_147), .A(n10465), .ZN(n10496) );
  OAI22_X1 U11200 ( .A1(n10469), .A2(keyinput_142), .B1(SI_17_), .B2(
        keyinput_143), .ZN(n10468) );
  AOI221_X1 U11201 ( .B1(n10469), .B2(keyinput_142), .C1(keyinput_143), .C2(
        SI_17_), .A(n10468), .ZN(n10495) );
  INV_X1 U11202 ( .A(keyinput_141), .ZN(n10488) );
  INV_X1 U11203 ( .A(keyinput_140), .ZN(n10486) );
  INV_X1 U11204 ( .A(keyinput_139), .ZN(n10483) );
  OAI22_X1 U11205 ( .A1(n10471), .A2(keyinput_136), .B1(SI_26_), .B2(
        keyinput_134), .ZN(n10470) );
  AOI221_X1 U11206 ( .B1(n10471), .B2(keyinput_136), .C1(keyinput_134), .C2(
        SI_26_), .A(n10470), .ZN(n10476) );
  OAI22_X1 U11207 ( .A1(n10474), .A2(keyinput_133), .B1(n10473), .B2(
        keyinput_137), .ZN(n10472) );
  AOI221_X1 U11208 ( .B1(n10474), .B2(keyinput_133), .C1(keyinput_137), .C2(
        n10473), .A(n10472), .ZN(n10475) );
  OAI211_X1 U11209 ( .C1(SI_25_), .C2(keyinput_135), .A(n10476), .B(n10475), 
        .ZN(n10477) );
  OAI22_X1 U11210 ( .A1(SI_31_), .A2(keyinput_129), .B1(P2_WR_REG_SCAN_IN), 
        .B2(keyinput_128), .ZN(n10478) );
  AOI221_X1 U11211 ( .B1(SI_31_), .B2(keyinput_129), .C1(keyinput_128), .C2(
        P2_WR_REG_SCAN_IN), .A(n10478), .ZN(n10480) );
  OAI21_X1 U11212 ( .B1(SI_29_), .B2(keyinput_131), .A(n5098), .ZN(n10481) );
  OAI221_X1 U11213 ( .B1(SI_19_), .B2(keyinput_141), .C1(n10489), .C2(n10488), 
        .A(n10487), .ZN(n10494) );
  XOR2_X1 U11214 ( .A(SI_16_), .B(keyinput_144), .Z(n10493) );
  AOI22_X1 U11215 ( .A1(SI_14_), .A2(keyinput_146), .B1(n10491), .B2(
        keyinput_145), .ZN(n10490) );
  OAI221_X1 U11216 ( .B1(SI_14_), .B2(keyinput_146), .C1(n10491), .C2(
        keyinput_145), .A(n10490), .ZN(n10492) );
  XNOR2_X1 U11217 ( .A(SI_9_), .B(keyinput_151), .ZN(n10505) );
  OAI22_X1 U11218 ( .A1(n10501), .A2(keyinput_152), .B1(keyinput_154), .B2(
        SI_6_), .ZN(n10500) );
  AOI221_X1 U11219 ( .B1(n10501), .B2(keyinput_152), .C1(SI_6_), .C2(
        keyinput_154), .A(n10500), .ZN(n10504) );
  OAI22_X1 U11220 ( .A1(SI_7_), .A2(keyinput_153), .B1(keyinput_155), .B2(
        SI_5_), .ZN(n10502) );
  AOI221_X1 U11221 ( .B1(SI_7_), .B2(keyinput_153), .C1(SI_5_), .C2(
        keyinput_155), .A(n10502), .ZN(n10503) );
  OAI211_X1 U11222 ( .C1(n10506), .C2(n10505), .A(n10504), .B(n10503), .ZN(
        n10507) );
  AOI22_X1 U11223 ( .A1(n10508), .A2(n10507), .B1(keyinput_158), .B2(SI_2_), 
        .ZN(n10509) );
  OAI21_X1 U11224 ( .B1(keyinput_158), .B2(SI_2_), .A(n10509), .ZN(n10510) );
  OAI221_X1 U11225 ( .B1(SI_1_), .B2(n10512), .C1(n10511), .C2(keyinput_159), 
        .A(n10510), .ZN(n10517) );
  AOI22_X1 U11226 ( .A1(P2_U3152), .A2(keyinput_162), .B1(n10514), .B2(
        keyinput_163), .ZN(n10513) );
  OAI221_X1 U11227 ( .B1(P2_U3152), .B2(keyinput_162), .C1(n10514), .C2(
        keyinput_163), .A(n10513), .ZN(n10516) );
  AOI22_X1 U11228 ( .A1(n10525), .A2(keyinput_168), .B1(keyinput_169), .B2(
        n10524), .ZN(n10523) );
  OAI221_X1 U11229 ( .B1(n10525), .B2(keyinput_168), .C1(n10524), .C2(
        keyinput_169), .A(n10523), .ZN(n10529) );
  AOI22_X1 U11230 ( .A1(n10527), .A2(keyinput_167), .B1(keyinput_166), .B2(
        n8280), .ZN(n10526) );
  OAI221_X1 U11231 ( .B1(n10527), .B2(keyinput_167), .C1(n8280), .C2(
        keyinput_166), .A(n10526), .ZN(n10528) );
  NAND2_X1 U11232 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_173), .ZN(
        n10530) );
  OAI221_X1 U11233 ( .B1(n10532), .B2(n10531), .C1(P2_REG3_REG_21__SCAN_IN), 
        .C2(keyinput_173), .A(n10530), .ZN(n10535) );
  OAI22_X1 U11234 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_178), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput_179), .ZN(n10533) );
  AOI221_X1 U11235 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_178), .C1(
        keyinput_179), .C2(P2_REG3_REG_24__SCAN_IN), .A(n10533), .ZN(n10534)
         );
  OAI221_X1 U11236 ( .B1(n10537), .B2(n10536), .C1(n10537), .C2(n10535), .A(
        n10534), .ZN(n10542) );
  AOI22_X1 U11237 ( .A1(n10540), .A2(keyinput_188), .B1(n10539), .B2(
        keyinput_189), .ZN(n10538) );
  OAI221_X1 U11238 ( .B1(n10540), .B2(keyinput_188), .C1(n10539), .C2(
        keyinput_189), .A(n10538), .ZN(n10541) );
  AOI21_X1 U11239 ( .B1(n10543), .B2(n10542), .A(n10541), .ZN(n10553) );
  AOI22_X1 U11240 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_190), .B1(
        n10545), .B2(keyinput_191), .ZN(n10544) );
  OAI221_X1 U11241 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_190), .C1(
        n10545), .C2(keyinput_191), .A(n10544), .ZN(n10552) );
  OAI22_X1 U11242 ( .A1(n10547), .A2(keyinput_192), .B1(keyinput_193), .B2(
        P2_DATAO_REG_31__SCAN_IN), .ZN(n10546) );
  AOI221_X1 U11243 ( .B1(n10547), .B2(keyinput_192), .C1(
        P2_DATAO_REG_31__SCAN_IN), .C2(keyinput_193), .A(n10546), .ZN(n10551)
         );
  OAI22_X1 U11244 ( .A1(n10549), .A2(keyinput_194), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_196), .ZN(n10548) );
  AOI221_X1 U11245 ( .B1(n10549), .B2(keyinput_194), .C1(keyinput_196), .C2(
        P2_DATAO_REG_28__SCAN_IN), .A(n10548), .ZN(n10550) );
  AOI22_X1 U11246 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(keyinput_202), .B1(
        n10555), .B2(keyinput_200), .ZN(n10554) );
  OAI221_X1 U11247 ( .B1(P2_DATAO_REG_22__SCAN_IN), .B2(keyinput_202), .C1(
        n10555), .C2(keyinput_200), .A(n10554), .ZN(n10559) );
  AOI22_X1 U11248 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(keyinput_201), .B1(
        n10557), .B2(keyinput_203), .ZN(n10556) );
  OAI221_X1 U11249 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_201), .C1(
        n10557), .C2(keyinput_203), .A(n10556), .ZN(n10558) );
  AOI22_X1 U11250 ( .A1(n10563), .A2(keyinput_205), .B1(n10562), .B2(
        keyinput_204), .ZN(n10561) );
  OAI221_X1 U11251 ( .B1(n10563), .B2(keyinput_205), .C1(n10562), .C2(
        keyinput_204), .A(n10561), .ZN(n10564) );
  AOI21_X1 U11252 ( .B1(n10566), .B2(n10565), .A(n10564), .ZN(n10578) );
  AOI22_X1 U11253 ( .A1(n10569), .A2(keyinput_208), .B1(keyinput_211), .B2(
        n10568), .ZN(n10567) );
  OAI221_X1 U11254 ( .B1(n10569), .B2(keyinput_208), .C1(n10568), .C2(
        keyinput_211), .A(n10567), .ZN(n10577) );
  AOI22_X1 U11255 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(keyinput_207), .B1(
        n10571), .B2(keyinput_206), .ZN(n10570) );
  OAI221_X1 U11256 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_207), .C1(
        n10571), .C2(keyinput_206), .A(n10570), .ZN(n10576) );
  AOI22_X1 U11257 ( .A1(n10574), .A2(keyinput_209), .B1(keyinput_210), .B2(
        n10573), .ZN(n10572) );
  OAI221_X1 U11258 ( .B1(n10574), .B2(keyinput_209), .C1(n10573), .C2(
        keyinput_210), .A(n10572), .ZN(n10575) );
  AOI22_X1 U11259 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_220), .B1(n10753), 
        .B2(keyinput_219), .ZN(n10581) );
  OAI221_X1 U11260 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_220), .C1(n10753), 
        .C2(keyinput_219), .A(n10581), .ZN(n10591) );
  AOI22_X1 U11261 ( .A1(n10584), .A2(keyinput_218), .B1(n10583), .B2(
        keyinput_221), .ZN(n10582) );
  OAI221_X1 U11262 ( .B1(n10584), .B2(keyinput_218), .C1(n10583), .C2(
        keyinput_221), .A(n10582), .ZN(n10588) );
  AOI22_X1 U11263 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput_216), .B1(
        n10586), .B2(keyinput_217), .ZN(n10585) );
  OAI221_X1 U11264 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_216), .C1(
        n10586), .C2(keyinput_217), .A(n10585), .ZN(n10587) );
  AOI211_X1 U11265 ( .C1(keyinput_215), .C2(P2_DATAO_REG_9__SCAN_IN), .A(
        n10588), .B(n10587), .ZN(n10589) );
  OAI21_X1 U11266 ( .B1(keyinput_215), .B2(P2_DATAO_REG_9__SCAN_IN), .A(n10589), .ZN(n10590) );
  XNOR2_X1 U11267 ( .A(n10593), .B(keyinput_224), .ZN(n10594) );
  NOR2_X1 U11268 ( .A1(n10595), .A2(n10594), .ZN(n10600) );
  INV_X1 U11269 ( .A(keyinput_225), .ZN(n10596) );
  MUX2_X1 U11270 ( .A(keyinput_225), .B(n10596), .S(P1_IR_REG_6__SCAN_IN), .Z(
        n10599) );
  XNOR2_X1 U11271 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_227), .ZN(n10598) );
  XNOR2_X1 U11272 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_226), .ZN(n10597) );
  OAI211_X1 U11273 ( .C1(n10600), .C2(n10599), .A(n10598), .B(n10597), .ZN(
        n10602) );
  NAND2_X1 U11274 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput_228), .ZN(n10601)
         );
  OAI211_X1 U11275 ( .C1(P1_IR_REG_9__SCAN_IN), .C2(keyinput_228), .A(n10602), 
        .B(n10601), .ZN(n10605) );
  INV_X1 U11276 ( .A(keyinput_229), .ZN(n10603) );
  MUX2_X1 U11277 ( .A(n10603), .B(keyinput_229), .S(P1_IR_REG_10__SCAN_IN), 
        .Z(n10604) );
  NAND2_X1 U11278 ( .A1(n10605), .A2(n10604), .ZN(n10612) );
  INV_X1 U11279 ( .A(keyinput_230), .ZN(n10606) );
  MUX2_X1 U11280 ( .A(n10606), .B(keyinput_230), .S(P1_IR_REG_11__SCAN_IN), 
        .Z(n10611) );
  OAI22_X1 U11281 ( .A1(n10608), .A2(keyinput_232), .B1(P1_IR_REG_12__SCAN_IN), 
        .B2(keyinput_231), .ZN(n10607) );
  AOI221_X1 U11282 ( .B1(n10608), .B2(keyinput_232), .C1(keyinput_231), .C2(
        P1_IR_REG_12__SCAN_IN), .A(n10607), .ZN(n10609) );
  INV_X1 U11283 ( .A(n10609), .ZN(n10610) );
  AOI21_X1 U11284 ( .B1(n10612), .B2(n10611), .A(n10610), .ZN(n10616) );
  XNOR2_X1 U11285 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_233), .ZN(n10615)
         );
  INV_X1 U11286 ( .A(keyinput_234), .ZN(n10613) );
  MUX2_X1 U11287 ( .A(keyinput_234), .B(n10613), .S(P1_IR_REG_15__SCAN_IN), 
        .Z(n10614) );
  OAI22_X1 U11288 ( .A1(n10619), .A2(keyinput_235), .B1(n10618), .B2(
        keyinput_237), .ZN(n10617) );
  AOI221_X1 U11289 ( .B1(n10619), .B2(keyinput_235), .C1(keyinput_237), .C2(
        n10618), .A(n10617), .ZN(n10621) );
  XNOR2_X1 U11290 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_236), .ZN(n10620)
         );
  NAND3_X1 U11291 ( .A1(n10622), .A2(n10621), .A3(n10620), .ZN(n10625) );
  XNOR2_X1 U11292 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_238), .ZN(n10624)
         );
  XNOR2_X1 U11293 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_239), .ZN(n10623)
         );
  NAND3_X1 U11294 ( .A1(n10625), .A2(n10624), .A3(n10623), .ZN(n10626) );
  OAI21_X1 U11295 ( .B1(keyinput_240), .B2(n10628), .A(n10626), .ZN(n10627) );
  AOI22_X1 U11296 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(keyinput_244), .B1(
        P1_IR_REG_23__SCAN_IN), .B2(keyinput_242), .ZN(n10631) );
  OAI221_X1 U11297 ( .B1(P1_IR_REG_25__SCAN_IN), .B2(keyinput_244), .C1(
        P1_IR_REG_23__SCAN_IN), .C2(keyinput_242), .A(n10631), .ZN(n10632) );
  XNOR2_X1 U11298 ( .A(n10633), .B(keyinput_247), .ZN(n10637) );
  XNOR2_X1 U11299 ( .A(n10634), .B(keyinput_245), .ZN(n10636) );
  XNOR2_X1 U11300 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_246), .ZN(n10635)
         );
  NOR3_X1 U11301 ( .A1(n10637), .A2(n10636), .A3(n10635), .ZN(n10640) );
  INV_X1 U11302 ( .A(keyinput_248), .ZN(n10638) );
  MUX2_X1 U11303 ( .A(keyinput_248), .B(n10638), .S(P1_IR_REG_29__SCAN_IN), 
        .Z(n10639) );
  AOI21_X1 U11304 ( .B1(n10641), .B2(n10640), .A(n10639), .ZN(n10644) );
  INV_X1 U11305 ( .A(keyinput_249), .ZN(n10642) );
  MUX2_X1 U11306 ( .A(n10642), .B(keyinput_249), .S(P1_IR_REG_30__SCAN_IN), 
        .Z(n10643) );
  NOR2_X1 U11307 ( .A1(n10644), .A2(n10643), .ZN(n10651) );
  AOI22_X1 U11308 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput_250), .B1(n10646), 
        .B2(keyinput_251), .ZN(n10645) );
  OAI221_X1 U11309 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput_250), .C1(n10646), .C2(keyinput_251), .A(n10645), .ZN(n10650) );
  XOR2_X1 U11310 ( .A(n10668), .B(keyinput_254), .Z(n10649) );
  OAI22_X1 U11311 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput_253), .B1(
        P1_D_REG_1__SCAN_IN), .B2(keyinput_252), .ZN(n10647) );
  AOI221_X1 U11312 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput_253), .C1(
        keyinput_252), .C2(P1_D_REG_1__SCAN_IN), .A(n10647), .ZN(n10648) );
  AOI21_X1 U11313 ( .B1(keyinput_255), .B2(n10653), .A(keyinput_127), .ZN(
        n10655) );
  INV_X1 U11314 ( .A(keyinput_255), .ZN(n10652) );
  AOI21_X1 U11315 ( .B1(n10653), .B2(n10652), .A(n10669), .ZN(n10654) );
  AOI22_X1 U11316 ( .A1(n10669), .A2(n10655), .B1(keyinput_127), .B2(n10654), 
        .ZN(n10656) );
  AOI222_X1 U11317 ( .A1(n10661), .A2(n10660), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10659), .C1(P2_DATAO_REG_19__SCAN_IN), .C2(n10658), .ZN(n10662) );
  XNOR2_X1 U11318 ( .A(n10663), .B(n10662), .ZN(P1_U3334) );
  MUX2_X1 U11319 ( .A(n10664), .B(n10753), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3353) );
  NOR2_X1 U11320 ( .A1(n10666), .A2(n10665), .ZN(n10698) );
  INV_X1 U11321 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10667) );
  NOR2_X1 U11322 ( .A1(n10686), .A2(n10667), .ZN(P1_U3321) );
  NOR2_X1 U11323 ( .A1(n10686), .A2(n10668), .ZN(P1_U3320) );
  NOR2_X1 U11324 ( .A1(n10686), .A2(n10669), .ZN(P1_U3319) );
  INV_X1 U11325 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10670) );
  NOR2_X1 U11326 ( .A1(n10686), .A2(n10670), .ZN(P1_U3318) );
  INV_X1 U11327 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10671) );
  NOR2_X1 U11328 ( .A1(n10686), .A2(n10671), .ZN(P1_U3317) );
  INV_X1 U11329 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10672) );
  NOR2_X1 U11330 ( .A1(n10686), .A2(n10672), .ZN(P1_U3316) );
  INV_X1 U11331 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10673) );
  NOR2_X1 U11332 ( .A1(n10686), .A2(n10673), .ZN(P1_U3315) );
  INV_X1 U11333 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10674) );
  NOR2_X1 U11334 ( .A1(n10686), .A2(n10674), .ZN(P1_U3314) );
  INV_X1 U11335 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10675) );
  NOR2_X1 U11336 ( .A1(n10686), .A2(n10675), .ZN(P1_U3313) );
  INV_X1 U11337 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10676) );
  NOR2_X1 U11338 ( .A1(n10686), .A2(n10676), .ZN(P1_U3312) );
  INV_X1 U11339 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10677) );
  NOR2_X1 U11340 ( .A1(n10686), .A2(n10677), .ZN(P1_U3311) );
  INV_X1 U11341 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10678) );
  NOR2_X1 U11342 ( .A1(n10686), .A2(n10678), .ZN(P1_U3310) );
  INV_X1 U11343 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10679) );
  NOR2_X1 U11344 ( .A1(n10686), .A2(n10679), .ZN(P1_U3309) );
  INV_X1 U11345 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10680) );
  NOR2_X1 U11346 ( .A1(n10686), .A2(n10680), .ZN(P1_U3308) );
  INV_X1 U11347 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10681) );
  NOR2_X1 U11348 ( .A1(n10686), .A2(n10681), .ZN(P1_U3307) );
  INV_X1 U11349 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10682) );
  NOR2_X1 U11350 ( .A1(n10686), .A2(n10682), .ZN(P1_U3306) );
  INV_X1 U11351 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10683) );
  NOR2_X1 U11352 ( .A1(n10686), .A2(n10683), .ZN(P1_U3305) );
  INV_X1 U11353 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10684) );
  NOR2_X1 U11354 ( .A1(n10686), .A2(n10684), .ZN(P1_U3304) );
  INV_X1 U11355 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10685) );
  NOR2_X1 U11356 ( .A1(n10686), .A2(n10685), .ZN(P1_U3303) );
  INV_X1 U11357 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10687) );
  NOR2_X1 U11358 ( .A1(n10698), .A2(n10687), .ZN(P1_U3302) );
  INV_X1 U11359 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10688) );
  NOR2_X1 U11360 ( .A1(n10698), .A2(n10688), .ZN(P1_U3301) );
  INV_X1 U11361 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10689) );
  NOR2_X1 U11362 ( .A1(n10698), .A2(n10689), .ZN(P1_U3300) );
  INV_X1 U11363 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10690) );
  NOR2_X1 U11364 ( .A1(n10698), .A2(n10690), .ZN(P1_U3299) );
  INV_X1 U11365 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10691) );
  NOR2_X1 U11366 ( .A1(n10698), .A2(n10691), .ZN(P1_U3298) );
  INV_X1 U11367 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10692) );
  NOR2_X1 U11368 ( .A1(n10698), .A2(n10692), .ZN(P1_U3297) );
  INV_X1 U11369 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10693) );
  NOR2_X1 U11370 ( .A1(n10698), .A2(n10693), .ZN(P1_U3296) );
  INV_X1 U11371 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10694) );
  NOR2_X1 U11372 ( .A1(n10698), .A2(n10694), .ZN(P1_U3295) );
  INV_X1 U11373 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10695) );
  NOR2_X1 U11374 ( .A1(n10698), .A2(n10695), .ZN(P1_U3294) );
  INV_X1 U11375 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10696) );
  NOR2_X1 U11376 ( .A1(n10698), .A2(n10696), .ZN(P1_U3293) );
  INV_X1 U11377 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10697) );
  NOR2_X1 U11378 ( .A1(n10698), .A2(n10697), .ZN(P1_U3292) );
  INV_X1 U11379 ( .A(n10699), .ZN(n10704) );
  AOI22_X1 U11380 ( .A1(n10772), .A2(n10704), .B1(n10703), .B2(n10769), .ZN(
        P2_U3438) );
  AND2_X1 U11381 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10769), .ZN(P2_U3326) );
  AND2_X1 U11382 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10769), .ZN(P2_U3325) );
  AND2_X1 U11383 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10769), .ZN(P2_U3324) );
  AND2_X1 U11384 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10769), .ZN(P2_U3323) );
  AND2_X1 U11385 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10769), .ZN(P2_U3322) );
  AND2_X1 U11386 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10769), .ZN(P2_U3321) );
  AND2_X1 U11387 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10769), .ZN(P2_U3320) );
  AND2_X1 U11388 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10769), .ZN(P2_U3319) );
  AND2_X1 U11389 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10769), .ZN(P2_U3318) );
  AND2_X1 U11390 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10769), .ZN(P2_U3317) );
  AND2_X1 U11391 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10769), .ZN(P2_U3316) );
  AND2_X1 U11392 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10769), .ZN(P2_U3315) );
  AND2_X1 U11393 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10769), .ZN(P2_U3314) );
  AND2_X1 U11394 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10769), .ZN(P2_U3313) );
  AND2_X1 U11395 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10769), .ZN(P2_U3312) );
  AND2_X1 U11396 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10769), .ZN(P2_U3311) );
  AND2_X1 U11397 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10769), .ZN(P2_U3310) );
  AND2_X1 U11398 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10769), .ZN(P2_U3309) );
  AND2_X1 U11399 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10769), .ZN(P2_U3308) );
  AND2_X1 U11400 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10769), .ZN(P2_U3307) );
  AND2_X1 U11401 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10769), .ZN(P2_U3306) );
  AND2_X1 U11402 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10769), .ZN(P2_U3305) );
  AND2_X1 U11403 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10769), .ZN(P2_U3304) );
  AND2_X1 U11404 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10769), .ZN(P2_U3303) );
  AND2_X1 U11405 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10769), .ZN(P2_U3302) );
  AND2_X1 U11406 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10769), .ZN(P2_U3301) );
  AND2_X1 U11407 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10769), .ZN(P2_U3300) );
  AND2_X1 U11408 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10769), .ZN(P2_U3299) );
  AND2_X1 U11409 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10769), .ZN(P2_U3298) );
  AND2_X1 U11410 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10769), .ZN(P2_U3297) );
  XOR2_X1 U11411 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  INV_X1 U11412 ( .A(n10705), .ZN(n10706) );
  NAND2_X1 U11413 ( .A1(n10707), .A2(n10706), .ZN(n10708) );
  XOR2_X1 U11414 ( .A(n10786), .B(n10708), .Z(ADD_1071_U5) );
  XOR2_X1 U11415 ( .A(n10710), .B(n10709), .Z(ADD_1071_U54) );
  XOR2_X1 U11416 ( .A(n10712), .B(n10711), .Z(ADD_1071_U53) );
  XNOR2_X1 U11417 ( .A(n10714), .B(n10713), .ZN(ADD_1071_U52) );
  NOR2_X1 U11418 ( .A1(n10716), .A2(n10715), .ZN(n10717) );
  XOR2_X1 U11419 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10717), .Z(ADD_1071_U51) );
  XOR2_X1 U11420 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10718), .Z(ADD_1071_U50) );
  XOR2_X1 U11421 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10719), .Z(ADD_1071_U49) );
  XOR2_X1 U11422 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10720), .Z(ADD_1071_U48) );
  XOR2_X1 U11423 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10721), .Z(ADD_1071_U47) );
  XOR2_X1 U11424 ( .A(n10723), .B(n10722), .Z(ADD_1071_U63) );
  XOR2_X1 U11425 ( .A(n10725), .B(n10724), .Z(ADD_1071_U62) );
  XNOR2_X1 U11426 ( .A(n10727), .B(n10726), .ZN(ADD_1071_U61) );
  XNOR2_X1 U11427 ( .A(n10729), .B(n10728), .ZN(ADD_1071_U60) );
  XNOR2_X1 U11428 ( .A(n10731), .B(n10730), .ZN(ADD_1071_U59) );
  XNOR2_X1 U11429 ( .A(n10733), .B(n10732), .ZN(ADD_1071_U58) );
  XNOR2_X1 U11430 ( .A(n10735), .B(n10734), .ZN(ADD_1071_U57) );
  XNOR2_X1 U11431 ( .A(n10737), .B(n10736), .ZN(ADD_1071_U56) );
  NOR2_X1 U11432 ( .A1(n10739), .A2(n10738), .ZN(n10740) );
  XOR2_X1 U11433 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(n10740), .Z(ADD_1071_U55)
         );
  AOI211_X1 U11434 ( .C1(n10753), .C2(n10741), .A(P1_U3084), .B(n5814), .ZN(
        n10743) );
  AOI22_X1 U11435 ( .A1(n10745), .A2(n10744), .B1(n10743), .B2(n10742), .ZN(
        n10748) );
  NOR3_X1 U11436 ( .A1(n10746), .A2(n10753), .A3(P1_REG1_REG_0__SCAN_IN), .ZN(
        n10747) );
  OR2_X1 U11437 ( .A1(n10748), .A2(n10747), .ZN(n10751) );
  AOI22_X1 U11438 ( .A1(n10761), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n10750) );
  OAI21_X1 U11439 ( .B1(n10752), .B2(n10751), .A(n10750), .ZN(P1_U3241) );
  NAND2_X1 U11440 ( .A1(n10753), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10757) );
  AOI211_X1 U11441 ( .C1(n10757), .C2(n10756), .A(n10755), .B(n10754), .ZN(
        n10758) );
  AOI21_X1 U11442 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(P1_U3084), .A(n10758), 
        .ZN(n10768) );
  AOI22_X1 U11443 ( .A1(n10761), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(n10760), 
        .B2(n10759), .ZN(n10767) );
  OAI211_X1 U11444 ( .C1(n10765), .C2(n10764), .A(n10763), .B(n10762), .ZN(
        n10766) );
  NAND3_X1 U11445 ( .A1(n10768), .A2(n10767), .A3(n10766), .ZN(P1_U3242) );
  AOI22_X1 U11446 ( .A1(n10772), .A2(n10771), .B1(n10770), .B2(n10769), .ZN(
        P2_U3437) );
  AOI22_X1 U11447 ( .A1(n10776), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n10809), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n10779) );
  OAI21_X1 U11448 ( .B1(n10773), .B2(P2_REG1_REG_0__SCAN_IN), .A(n10792), .ZN(
        n10774) );
  AOI21_X1 U11449 ( .B1(n10776), .B2(n10775), .A(n10774), .ZN(n10778) );
  AOI22_X1 U11450 ( .A1(n10800), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10777) );
  OAI221_X1 U11451 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n10779), .C1(n10794), .C2(
        n10778), .A(n10777), .ZN(P2_U3245) );
  NAND2_X1 U11452 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10780) );
  AND2_X1 U11453 ( .A1(n10781), .A2(n10780), .ZN(n10782) );
  OR2_X1 U11454 ( .A1(n10783), .A2(n10782), .ZN(n10784) );
  OR2_X1 U11455 ( .A1(n10801), .A2(n10784), .ZN(n10790) );
  OAI22_X1 U11456 ( .A1(n10787), .A2(n10786), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10785), .ZN(n10788) );
  INV_X1 U11457 ( .A(n10788), .ZN(n10789) );
  OAI211_X1 U11458 ( .C1(n10792), .C2(n10791), .A(n10790), .B(n10789), .ZN(
        n10793) );
  INV_X1 U11459 ( .A(n10793), .ZN(n10799) );
  INV_X1 U11460 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10835) );
  NOR2_X1 U11461 ( .A1(n10794), .A2(n10835), .ZN(n10797) );
  OAI211_X1 U11462 ( .C1(n10797), .C2(n10796), .A(n10809), .B(n10795), .ZN(
        n10798) );
  NAND2_X1 U11463 ( .A1(n10799), .A2(n10798), .ZN(P2_U3246) );
  AOI22_X1 U11464 ( .A1(n10800), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n10814) );
  AOI211_X1 U11465 ( .C1(n10804), .C2(n10803), .A(n10802), .B(n10801), .ZN(
        n10805) );
  AOI21_X1 U11466 ( .B1(n10807), .B2(n10806), .A(n10805), .ZN(n10813) );
  OAI211_X1 U11467 ( .C1(n10811), .C2(n10810), .A(n10809), .B(n10808), .ZN(
        n10812) );
  NAND3_X1 U11468 ( .A1(n10814), .A2(n10813), .A3(n10812), .ZN(P2_U3247) );
  XNOR2_X1 U11469 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  NAND2_X1 U11470 ( .A1(n10816), .A2(n10815), .ZN(n10832) );
  AOI21_X1 U11471 ( .B1(n10819), .B2(n10818), .A(n10817), .ZN(n10826) );
  AOI22_X1 U11472 ( .A1(n10832), .A2(n10822), .B1(n10821), .B2(n10820), .ZN(
        n10834) );
  OAI22_X1 U11473 ( .A1(n10834), .A2(n9303), .B1(n10824), .B2(n10823), .ZN(
        n10825) );
  AOI211_X1 U11474 ( .C1(n10827), .C2(n10832), .A(n10826), .B(n10825), .ZN(
        n10828) );
  OAI21_X1 U11475 ( .B1(n10775), .B2(n10829), .A(n10828), .ZN(P2_U3296) );
  AOI22_X1 U11476 ( .A1(n10832), .A2(n10980), .B1(n10831), .B2(n10830), .ZN(
        n10833) );
  AND2_X1 U11477 ( .A1(n10834), .A2(n10833), .ZN(n10837) );
  AOI22_X1 U11478 ( .A1(n11002), .A2(n10837), .B1(n10835), .B2(n11000), .ZN(
        P2_U3520) );
  INV_X1 U11479 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U11480 ( .A1(n11006), .A2(n10837), .B1(n10836), .B2(n11003), .ZN(
        P2_U3451) );
  INV_X1 U11481 ( .A(n10844), .ZN(n10842) );
  AOI21_X1 U11482 ( .B1(n10946), .B2(n10839), .A(n10838), .ZN(n10840) );
  OAI211_X1 U11483 ( .C1(n10923), .C2(n10842), .A(n10841), .B(n10840), .ZN(
        n10843) );
  AOI21_X1 U11484 ( .B1(n10929), .B2(n10844), .A(n10843), .ZN(n10846) );
  INV_X1 U11485 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U11486 ( .A1(n11024), .A2(n10846), .B1(n10845), .B2(n11023), .ZN(
        P1_U3524) );
  AOI22_X1 U11487 ( .A1(n11028), .A2(n10846), .B1(n5784), .B2(n11025), .ZN(
        P1_U3457) );
  NAND3_X1 U11488 ( .A1(n10848), .A2(n10847), .A3(n10881), .ZN(n10849) );
  OAI211_X1 U11489 ( .C1(n10851), .C2(n10992), .A(n10850), .B(n10849), .ZN(
        n10852) );
  AOI21_X1 U11490 ( .B1(n10980), .B2(n10853), .A(n10852), .ZN(n10855) );
  AOI22_X1 U11491 ( .A1(n11002), .A2(n10855), .B1(n6792), .B2(n11000), .ZN(
        P2_U3521) );
  INV_X1 U11492 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U11493 ( .A1(n11006), .A2(n10855), .B1(n10854), .B2(n11003), .ZN(
        P2_U3454) );
  INV_X1 U11494 ( .A(n10923), .ZN(n11014) );
  INV_X1 U11495 ( .A(n10856), .ZN(n10858) );
  OAI22_X1 U11496 ( .A1(n10858), .A2(n11009), .B1(n10857), .B2(n11018), .ZN(
        n10860) );
  AOI211_X1 U11497 ( .C1(n11014), .C2(n10861), .A(n10860), .B(n10859), .ZN(
        n10863) );
  INV_X1 U11498 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U11499 ( .A1(n11024), .A2(n10863), .B1(n10862), .B2(n11023), .ZN(
        P1_U3525) );
  AOI22_X1 U11500 ( .A1(n11028), .A2(n10863), .B1(n5805), .B2(n11025), .ZN(
        P1_U3460) );
  OAI22_X1 U11501 ( .A1(n10865), .A2(n10994), .B1(n10864), .B2(n10992), .ZN(
        n10866) );
  NOR2_X1 U11502 ( .A1(n10867), .A2(n10866), .ZN(n10869) );
  AOI22_X1 U11503 ( .A1(n11002), .A2(n10869), .B1(n6790), .B2(n11000), .ZN(
        P2_U3522) );
  INV_X1 U11504 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10868) );
  AOI22_X1 U11505 ( .A1(n11006), .A2(n10869), .B1(n10868), .B2(n11003), .ZN(
        P2_U3457) );
  OAI22_X1 U11506 ( .A1(n10871), .A2(n11009), .B1(n10870), .B2(n11018), .ZN(
        n10873) );
  AOI211_X1 U11507 ( .C1(n11014), .C2(n10874), .A(n10873), .B(n10872), .ZN(
        n10876) );
  INV_X1 U11508 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10875) );
  AOI22_X1 U11509 ( .A1(n11024), .A2(n10876), .B1(n10875), .B2(n11023), .ZN(
        P1_U3526) );
  AOI22_X1 U11510 ( .A1(n11028), .A2(n10876), .B1(n5833), .B2(n11025), .ZN(
        P1_U3463) );
  NOR2_X1 U11511 ( .A1(n10992), .A2(n10877), .ZN(n10879) );
  AOI211_X1 U11512 ( .C1(n10881), .C2(n10880), .A(n10879), .B(n10878), .ZN(
        n10883) );
  AOI22_X1 U11513 ( .A1(n11002), .A2(n10883), .B1(n6789), .B2(n11000), .ZN(
        P2_U3523) );
  INV_X1 U11514 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10882) );
  AOI22_X1 U11515 ( .A1(n11006), .A2(n10883), .B1(n10882), .B2(n11003), .ZN(
        P2_U3460) );
  OAI22_X1 U11516 ( .A1(n10884), .A2(n11009), .B1(n7411), .B2(n11018), .ZN(
        n10886) );
  AOI211_X1 U11517 ( .C1(n11014), .C2(n10887), .A(n10886), .B(n10885), .ZN(
        n10888) );
  AOI22_X1 U11518 ( .A1(n11024), .A2(n10888), .B1(n6623), .B2(n11023), .ZN(
        P1_U3527) );
  AOI22_X1 U11519 ( .A1(n11028), .A2(n10888), .B1(n5857), .B2(n11025), .ZN(
        P1_U3466) );
  OAI21_X1 U11520 ( .B1(n10890), .B2(n11018), .A(n10889), .ZN(n10892) );
  AOI211_X1 U11521 ( .C1(n10893), .C2(n10948), .A(n10892), .B(n10891), .ZN(
        n10895) );
  INV_X1 U11522 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U11523 ( .A1(n11024), .A2(n10895), .B1(n10894), .B2(n11023), .ZN(
        P1_U3528) );
  AOI22_X1 U11524 ( .A1(n11028), .A2(n10895), .B1(n5885), .B2(n11025), .ZN(
        P1_U3469) );
  OAI211_X1 U11525 ( .C1(n10898), .C2(n10992), .A(n10897), .B(n10896), .ZN(
        n10899) );
  AOI21_X1 U11526 ( .B1(n10980), .B2(n10900), .A(n10899), .ZN(n10902) );
  AOI22_X1 U11527 ( .A1(n11002), .A2(n10902), .B1(n7112), .B2(n11000), .ZN(
        P2_U3525) );
  INV_X1 U11528 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10901) );
  AOI22_X1 U11529 ( .A1(n11006), .A2(n10902), .B1(n10901), .B2(n11003), .ZN(
        P2_U3466) );
  AOI22_X1 U11530 ( .A1(n10904), .A2(n11021), .B1(n10946), .B2(n10903), .ZN(
        n10905) );
  OAI211_X1 U11531 ( .C1(n10907), .C2(n10923), .A(n10906), .B(n10905), .ZN(
        n10908) );
  INV_X1 U11532 ( .A(n10908), .ZN(n10910) );
  INV_X1 U11533 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U11534 ( .A1(n11024), .A2(n10910), .B1(n10909), .B2(n11023), .ZN(
        P1_U3529) );
  AOI22_X1 U11535 ( .A1(n11028), .A2(n10910), .B1(n5899), .B2(n11025), .ZN(
        P1_U3472) );
  NOR2_X1 U11536 ( .A1(n10911), .A2(n10990), .ZN(n10917) );
  OAI22_X1 U11537 ( .A1(n10913), .A2(n10994), .B1(n10912), .B2(n10992), .ZN(
        n10915) );
  AOI211_X1 U11538 ( .C1(n10917), .C2(n10916), .A(n10915), .B(n10914), .ZN(
        n10919) );
  AOI22_X1 U11539 ( .A1(n11002), .A2(n10919), .B1(n7121), .B2(n11000), .ZN(
        P2_U3526) );
  INV_X1 U11540 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10918) );
  AOI22_X1 U11541 ( .A1(n11006), .A2(n10919), .B1(n10918), .B2(n11003), .ZN(
        P2_U3469) );
  INV_X1 U11542 ( .A(n10924), .ZN(n10928) );
  AOI21_X1 U11543 ( .B1(n10946), .B2(n10921), .A(n10920), .ZN(n10922) );
  OAI21_X1 U11544 ( .B1(n10924), .B2(n10923), .A(n10922), .ZN(n10927) );
  INV_X1 U11545 ( .A(n10925), .ZN(n10926) );
  AOI211_X1 U11546 ( .C1(n10929), .C2(n10928), .A(n10927), .B(n10926), .ZN(
        n10930) );
  AOI22_X1 U11547 ( .A1(n11024), .A2(n10930), .B1(n6633), .B2(n11023), .ZN(
        P1_U3530) );
  AOI22_X1 U11548 ( .A1(n11028), .A2(n10930), .B1(n5930), .B2(n11025), .ZN(
        P1_U3475) );
  OAI22_X1 U11549 ( .A1(n10932), .A2(n10994), .B1(n10931), .B2(n10992), .ZN(
        n10934) );
  AOI211_X1 U11550 ( .C1(n10980), .C2(n10935), .A(n10934), .B(n10933), .ZN(
        n10937) );
  AOI22_X1 U11551 ( .A1(n11002), .A2(n10937), .B1(n7320), .B2(n11000), .ZN(
        P2_U3527) );
  INV_X1 U11552 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10936) );
  AOI22_X1 U11553 ( .A1(n11006), .A2(n10937), .B1(n10936), .B2(n11003), .ZN(
        P2_U3472) );
  INV_X1 U11554 ( .A(n10938), .ZN(n10943) );
  INV_X1 U11555 ( .A(n10939), .ZN(n10940) );
  OAI22_X1 U11556 ( .A1(n10940), .A2(n11009), .B1(n5311), .B2(n11018), .ZN(
        n10942) );
  AOI211_X1 U11557 ( .C1(n11014), .C2(n10943), .A(n10942), .B(n10941), .ZN(
        n10944) );
  AOI22_X1 U11558 ( .A1(n11024), .A2(n10944), .B1(n6635), .B2(n11023), .ZN(
        P1_U3531) );
  AOI22_X1 U11559 ( .A1(n11028), .A2(n10944), .B1(n5955), .B2(n11025), .ZN(
        P1_U3478) );
  AOI22_X1 U11560 ( .A1(n10947), .A2(n11021), .B1(n10946), .B2(n10945), .ZN(
        n10951) );
  NAND2_X1 U11561 ( .A1(n10949), .A2(n10948), .ZN(n10950) );
  AOI22_X1 U11562 ( .A1(n11024), .A2(n10954), .B1(n6622), .B2(n11023), .ZN(
        P1_U3532) );
  INV_X1 U11563 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10953) );
  AOI22_X1 U11564 ( .A1(n11028), .A2(n10954), .B1(n10953), .B2(n11025), .ZN(
        P1_U3481) );
  NOR3_X1 U11565 ( .A1(n10956), .A2(n10955), .A3(n10994), .ZN(n10958) );
  AOI211_X1 U11566 ( .C1(n10971), .C2(n10959), .A(n10958), .B(n10957), .ZN(
        n10961) );
  AOI22_X1 U11567 ( .A1(n11002), .A2(n10961), .B1(n7528), .B2(n11000), .ZN(
        P2_U3529) );
  INV_X1 U11568 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U11569 ( .A1(n11006), .A2(n10961), .B1(n10960), .B2(n11003), .ZN(
        P2_U3478) );
  OAI21_X1 U11570 ( .B1(n10963), .B2(n11018), .A(n10962), .ZN(n10965) );
  AOI211_X1 U11571 ( .C1(n11014), .C2(n10966), .A(n10965), .B(n10964), .ZN(
        n10967) );
  AOI22_X1 U11572 ( .A1(n11024), .A2(n10967), .B1(n6639), .B2(n11023), .ZN(
        P1_U3534) );
  AOI22_X1 U11573 ( .A1(n11028), .A2(n10967), .B1(n5750), .B2(n11025), .ZN(
        P1_U3487) );
  AOI211_X1 U11574 ( .C1(n10971), .C2(n10970), .A(n10969), .B(n10968), .ZN(
        n10974) );
  AOI22_X1 U11575 ( .A1(n11002), .A2(n10974), .B1(n10972), .B2(n11000), .ZN(
        P2_U3531) );
  INV_X1 U11576 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10973) );
  AOI22_X1 U11577 ( .A1(n11006), .A2(n10974), .B1(n10973), .B2(n11003), .ZN(
        P2_U3484) );
  OAI22_X1 U11578 ( .A1(n10976), .A2(n10994), .B1(n10975), .B2(n10992), .ZN(
        n10978) );
  AOI211_X1 U11579 ( .C1(n10980), .C2(n10979), .A(n10978), .B(n10977), .ZN(
        n10982) );
  AOI22_X1 U11580 ( .A1(n11002), .A2(n10982), .B1(n7791), .B2(n11000), .ZN(
        P2_U3532) );
  INV_X1 U11581 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10981) );
  AOI22_X1 U11582 ( .A1(n11006), .A2(n10982), .B1(n10981), .B2(n11003), .ZN(
        P2_U3487) );
  OAI22_X1 U11583 ( .A1(n10984), .A2(n11009), .B1(n10983), .B2(n11018), .ZN(
        n10986) );
  AOI211_X1 U11584 ( .C1(n11014), .C2(n10987), .A(n10986), .B(n10985), .ZN(
        n10989) );
  AOI22_X1 U11585 ( .A1(n11024), .A2(n10989), .B1(n10988), .B2(n11023), .ZN(
        P1_U3536) );
  AOI22_X1 U11586 ( .A1(n11028), .A2(n10989), .B1(n6054), .B2(n11025), .ZN(
        P1_U3493) );
  NOR2_X1 U11587 ( .A1(n10991), .A2(n10990), .ZN(n10999) );
  OAI22_X1 U11588 ( .A1(n10995), .A2(n10994), .B1(n10993), .B2(n10992), .ZN(
        n10997) );
  AOI211_X1 U11589 ( .C1(n10999), .C2(n10998), .A(n10997), .B(n10996), .ZN(
        n11005) );
  AOI22_X1 U11590 ( .A1(n11002), .A2(n11005), .B1(n11001), .B2(n11000), .ZN(
        P2_U3533) );
  INV_X1 U11591 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11004) );
  AOI22_X1 U11592 ( .A1(n11006), .A2(n11005), .B1(n11004), .B2(n11003), .ZN(
        P2_U3490) );
  INV_X1 U11593 ( .A(n11007), .ZN(n11013) );
  OAI22_X1 U11594 ( .A1(n11010), .A2(n11009), .B1(n11008), .B2(n11018), .ZN(
        n11012) );
  AOI211_X1 U11595 ( .C1(n11014), .C2(n11013), .A(n11012), .B(n11011), .ZN(
        n11016) );
  AOI22_X1 U11596 ( .A1(n11024), .A2(n11016), .B1(n11015), .B2(n11023), .ZN(
        P1_U3538) );
  AOI22_X1 U11597 ( .A1(n11028), .A2(n11016), .B1(n6100), .B2(n11025), .ZN(
        P1_U3499) );
  OAI21_X1 U11598 ( .B1(n11019), .B2(n11018), .A(n11017), .ZN(n11020) );
  AOI21_X1 U11599 ( .B1(n11022), .B2(n11021), .A(n11020), .ZN(n11027) );
  AOI22_X1 U11600 ( .A1(n11024), .A2(n11027), .B1(n8461), .B2(n11023), .ZN(
        P1_U3553) );
  INV_X1 U11601 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n11026) );
  AOI22_X1 U11602 ( .A1(n11028), .A2(n11027), .B1(n11026), .B2(n11025), .ZN(
        P1_U3521) );
  XNOR2_X1 U11603 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  NAND2_X2 U5131 ( .A1(n6521), .A2(n9423), .ZN(n8253) );
  AND3_X1 U5101 ( .A1(n5822), .A2(n5821), .A3(n5820), .ZN(n10857) );
endmodule

