

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598;

  MUX2_X1 U4936 ( .A(n9395), .B(n9394), .S(n9683), .Z(n9397) );
  NAND2_X1 U4937 ( .A1(n8581), .A2(n8406), .ZN(n6557) );
  NAND2_X1 U4938 ( .A1(n8153), .A2(n8152), .ZN(n9683) );
  BUF_X1 U4939 ( .A(n6693), .Z(n6838) );
  NAND2_X1 U4940 ( .A1(n5808), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9179) );
  OR2_X1 U4941 ( .A1(n9113), .A2(n7724), .ZN(n9458) );
  NAND2_X1 U4942 ( .A1(n7984), .A2(n10147), .ZN(n7616) );
  AND2_X1 U4943 ( .A1(n4954), .A2(n4955), .ZN(n4953) );
  INV_X1 U4944 ( .A(n5629), .ZN(n7762) );
  INV_X1 U4945 ( .A(n9920), .ZN(n9511) );
  INV_X1 U4946 ( .A(n8151), .ZN(n5876) );
  CLKBUF_X2 U4947 ( .A(n6225), .Z(n7973) );
  NAND2_X1 U4948 ( .A1(n6175), .A2(n6173), .ZN(n6223) );
  NOR2_X1 U4949 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4860) );
  AND2_X1 U4950 ( .A1(n6103), .A2(n4991), .ZN(n9680) );
  INV_X1 U4951 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5780) );
  OR2_X1 U4952 ( .A1(n8579), .A2(n4825), .ZN(n4824) );
  INV_X1 U4953 ( .A(n7969), .ZN(n6474) );
  NAND2_X1 U4954 ( .A1(n6547), .A2(n8144), .ZN(n6370) );
  AND2_X1 U4955 ( .A1(n8874), .A2(n8611), .ZN(n8526) );
  INV_X1 U4956 ( .A(n8570), .ZN(n8577) );
  INV_X2 U4957 ( .A(n6832), .ZN(n6837) );
  NAND2_X1 U4958 ( .A1(n5576), .A2(n10139), .ZN(n9292) );
  NAND2_X1 U4959 ( .A1(n7809), .A2(n6071), .ZN(n7365) );
  INV_X2 U4960 ( .A(n8090), .ZN(n8101) );
  INV_X1 U4961 ( .A(n6312), .ZN(n6494) );
  CLKBUF_X2 U4962 ( .A(n6665), .Z(n6843) );
  INV_X1 U4963 ( .A(n5643), .ZN(n5894) );
  AND4_X1 U4964 ( .A1(n6284), .A2(n6283), .A3(n6282), .A4(n6281), .ZN(n7851)
         );
  INV_X1 U4965 ( .A(n5359), .ZN(n6539) );
  NAND2_X1 U4966 ( .A1(n8401), .A2(n8400), .ZN(n8994) );
  NAND2_X1 U4967 ( .A1(n4550), .A2(n8554), .ZN(n8798) );
  INV_X1 U4968 ( .A(n7867), .ZN(n9145) );
  OR2_X1 U4969 ( .A1(n6599), .A2(n6594), .ZN(n7769) );
  NAND2_X1 U4970 ( .A1(n5506), .A2(n4652), .ZN(n7452) );
  INV_X1 U4971 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5456) );
  AND2_X1 U4972 ( .A1(n6255), .A2(n6254), .ZN(n7566) );
  BUF_X1 U4973 ( .A(n5416), .Z(n6994) );
  INV_X1 U4974 ( .A(n7742), .ZN(n7816) );
  NAND2_X1 U4975 ( .A1(n5915), .A2(n5914), .ZN(n9821) );
  INV_X1 U4976 ( .A(n9302), .ZN(n9557) );
  MUX2_X1 U4977 ( .A(n10020), .B(n10019), .S(n10155), .Z(n10021) );
  AND4_X2 U4978 ( .A1(n5455), .A2(n5454), .A3(n6060), .A4(n6064), .ZN(n4430)
         );
  BUF_X1 U4979 ( .A(n7027), .Z(n4431) );
  BUF_X4 U4980 ( .A(n7027), .Z(n4432) );
  INV_X2 U4981 ( .A(n5543), .ZN(n7027) );
  NAND2_X2 U4982 ( .A1(n9148), .A2(n9149), .ZN(n5086) );
  NAND2_X2 U4983 ( .A1(n9410), .A2(n7364), .ZN(n7363) );
  AND2_X2 U4984 ( .A1(n8939), .A2(n10213), .ZN(n4740) );
  NOR2_X2 U4985 ( .A1(n9506), .A2(n9505), .ZN(n9523) );
  CLKBUF_X2 U4986 ( .A(n7163), .Z(n8461) );
  MUX2_X1 U4987 ( .A(n10061), .B(n10062), .S(n5543), .Z(n7742) );
  OAI21_X2 U4988 ( .B1(n6889), .B2(n10229), .A(n5218), .ZN(n6890) );
  NAND2_X2 U4989 ( .A1(n9732), .A2(n9733), .ZN(n4864) );
  NAND2_X2 U4990 ( .A1(n6086), .A2(n9444), .ZN(n9732) );
  AOI21_X2 U4991 ( .B1(n9376), .B2(n9754), .A(n9375), .ZN(n9386) );
  NAND2_X2 U4992 ( .A1(n7046), .A2(n7045), .ZN(n9613) );
  INV_X2 U4993 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5477) );
  NAND2_X2 U4994 ( .A1(n5472), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U4995 ( .A1(n6157), .A2(n9578), .ZN(n4433) );
  NAND2_X1 U4996 ( .A1(n6157), .A2(n9578), .ZN(n4434) );
  NOR2_X2 U4997 ( .A1(n5423), .A2(n6253), .ZN(n6912) );
  NAND3_X2 U4998 ( .A1(n4935), .A2(n4936), .A3(n5538), .ZN(n5557) );
  XNOR2_X2 U4999 ( .A(n5473), .B(n5458), .ZN(n6157) );
  AOI21_X2 U5000 ( .B1(n8460), .B2(n7142), .A(n6506), .ZN(n7162) );
  OAI21_X2 U5001 ( .B1(n4858), .B2(n4498), .A(n6076), .ZN(n4855) );
  XNOR2_X1 U5002 ( .A(n5306), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U5003 ( .A1(n8798), .A2(n8561), .ZN(n5118) );
  NAND2_X2 U5004 ( .A1(n9502), .A2(n9504), .ZN(n9689) );
  NAND2_X1 U5005 ( .A1(n6144), .A2(n6143), .ZN(n6163) );
  NAND2_X1 U5006 ( .A1(n5945), .A2(n5944), .ZN(n9957) );
  NAND2_X1 U5007 ( .A1(n7473), .A2(n7474), .ZN(n7472) );
  INV_X1 U5009 ( .A(n8411), .ZN(n5129) );
  INV_X1 U5010 ( .A(n9868), .ZN(n9897) );
  NAND2_X1 U5011 ( .A1(n9556), .A2(n7762), .ZN(n9408) );
  INV_X1 U5012 ( .A(n9914), .ZN(n9280) );
  NAND2_X1 U5013 ( .A1(n9292), .A2(n9449), .ZN(n9413) );
  NAND2_X1 U5014 ( .A1(n9557), .A2(n10103), .ZN(n9415) );
  NAND2_X1 U5015 ( .A1(n7164), .A2(n6507), .ZN(n7356) );
  CLKBUF_X2 U5016 ( .A(n6619), .Z(n6693) );
  CLKBUF_X1 U5017 ( .A(n6632), .Z(n6845) );
  NAND2_X2 U5018 ( .A1(n8467), .A2(n8485), .ZN(n7355) );
  NAND2_X2 U5019 ( .A1(n6072), .A2(n9452), .ZN(n9410) );
  INV_X2 U5020 ( .A(n9394), .ZN(n9381) );
  AOI21_X1 U5021 ( .B1(n7017), .B2(n4919), .A(n4538), .ZN(n4917) );
  INV_X1 U5022 ( .A(n8617), .ZN(n7592) );
  NAND4_X1 U5023 ( .A1(n6264), .A2(n6263), .A3(n6262), .A4(n6261), .ZN(n8617)
         );
  INV_X1 U5024 ( .A(n9556), .ZN(n7984) );
  AND2_X2 U5025 ( .A1(n6105), .A2(n6062), .ZN(n6068) );
  CLKBUF_X1 U5026 ( .A(n6593), .Z(n9447) );
  CLKBUF_X2 U5027 ( .A(n6223), .Z(n6312) );
  INV_X2 U5028 ( .A(n7130), .ZN(n6530) );
  INV_X1 U5029 ( .A(n7239), .ZN(n6191) );
  CLKBUF_X1 U5030 ( .A(n5636), .Z(n6112) );
  AND2_X1 U5031 ( .A1(n4746), .A2(n5308), .ZN(n5289) );
  NAND4_X1 U5032 ( .A1(n4861), .A2(n4860), .A3(n10272), .A4(n5456), .ZN(n5457)
         );
  AND3_X1 U5033 ( .A1(n5242), .A2(n5241), .A3(n5310), .ZN(n4746) );
  NOR2_X1 U5034 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n5255) );
  CLKBUF_X2 U5035 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n10061) );
  OAI21_X1 U5036 ( .B1(n8442), .B2(n8994), .A(n5231), .ZN(n8445) );
  AND2_X1 U5037 ( .A1(n4561), .A2(n4560), .ZN(n10019) );
  XNOR2_X1 U5038 ( .A(n4539), .B(n9689), .ZN(n6161) );
  AND2_X1 U5039 ( .A1(n9935), .A2(n4630), .ZN(n10015) );
  NAND2_X1 U5040 ( .A1(n4625), .A2(n4624), .ZN(n9939) );
  NAND2_X1 U5041 ( .A1(n6152), .A2(n9501), .ZN(n4539) );
  NAND2_X1 U5042 ( .A1(n6527), .A2(n8432), .ZN(n8179) );
  NAND2_X1 U5043 ( .A1(n5118), .A2(n5117), .ZN(n6527) );
  OAI21_X1 U5044 ( .B1(n9936), .B2(n10143), .A(n9934), .ZN(n4631) );
  CLKBUF_X1 U5045 ( .A(n6524), .Z(n4632) );
  NAND2_X1 U5046 ( .A1(n4554), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8685) );
  NAND2_X1 U5047 ( .A1(n6081), .A2(n9487), .ZN(n9803) );
  NAND2_X1 U5048 ( .A1(n5080), .A2(n5079), .ZN(n9157) );
  OR2_X1 U5049 ( .A1(n6163), .A2(n6145), .ZN(n9502) );
  NAND2_X1 U5050 ( .A1(n4549), .A2(n4548), .ZN(n9851) );
  XNOR2_X1 U5051 ( .A(n8138), .B(SI_29_), .ZN(n8109) );
  NAND2_X2 U5052 ( .A1(n6042), .A2(n6041), .ZN(n6873) );
  NAND2_X1 U5053 ( .A1(n4556), .A2(n5432), .ZN(n8646) );
  AND2_X1 U5054 ( .A1(n6526), .A2(n8560), .ZN(n5117) );
  AND2_X1 U5055 ( .A1(n9740), .A2(n10022), .ZN(n9706) );
  AOI21_X1 U5056 ( .B1(n5112), .B2(n5114), .A(n5110), .ZN(n5109) );
  NAND2_X1 U5057 ( .A1(n6040), .A2(n6039), .ZN(n6138) );
  NOR2_X1 U5058 ( .A1(n9646), .A2(n9645), .ZN(n9661) );
  NAND2_X1 U5059 ( .A1(n6014), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U5060 ( .A1(n7472), .A2(n6639), .ZN(n7398) );
  NAND2_X1 U5061 ( .A1(n5428), .A2(n6973), .ZN(n5429) );
  NAND2_X1 U5062 ( .A1(n7420), .A2(n7419), .ZN(n7548) );
  NAND2_X1 U5063 ( .A1(n5890), .A2(n5889), .ZN(n9971) );
  AND2_X1 U5064 ( .A1(n5152), .A2(n7306), .ZN(n7344) );
  NAND2_X1 U5065 ( .A1(n5904), .A2(n5903), .ZN(n9966) );
  NAND2_X1 U5066 ( .A1(n5878), .A2(n5877), .ZN(n9975) );
  NAND2_X1 U5067 ( .A1(n6351), .A2(n6350), .ZN(n9055) );
  NAND2_X1 U5068 ( .A1(n5806), .A2(n5805), .ZN(n6720) );
  OAI21_X1 U5069 ( .B1(n5922), .B2(n5921), .A(n5920), .ZN(n5981) );
  NAND2_X1 U5070 ( .A1(n6322), .A2(n6321), .ZN(n7913) );
  INV_X1 U5071 ( .A(n8298), .ZN(n7966) );
  NAND2_X1 U5072 ( .A1(n6382), .A2(n6381), .ZN(n8969) );
  XNOR2_X1 U5073 ( .A(n8988), .B(n8613), .ZN(n8411) );
  NAND2_X1 U5074 ( .A1(n5835), .A2(n5834), .ZN(n9988) );
  NAND2_X1 U5075 ( .A1(n4829), .A2(n6311), .ZN(n8298) );
  XNOR2_X1 U5076 ( .A(n5801), .B(n5800), .ZN(n7372) );
  AND2_X1 U5077 ( .A1(n5722), .A2(n5721), .ZN(n7867) );
  NAND2_X2 U5078 ( .A1(n5765), .A2(n5764), .ZN(n10003) );
  NAND2_X1 U5079 ( .A1(n4623), .A2(n9554), .ZN(n9342) );
  NAND2_X1 U5080 ( .A1(n6299), .A2(n6298), .ZN(n8988) );
  NAND2_X1 U5081 ( .A1(n5693), .A2(n5692), .ZN(n9326) );
  OR2_X1 U5082 ( .A1(n7859), .A2(n7850), .ZN(n8494) );
  CLKBUF_X1 U5083 ( .A(n7859), .Z(n4644) );
  OAI21_X1 U5084 ( .B1(n5845), .B2(n5844), .A(n5843), .ZN(n5863) );
  AND2_X1 U5085 ( .A1(n5712), .A2(n5731), .ZN(n6975) );
  INV_X1 U5087 ( .A(n7783), .ZN(n7986) );
  NAND2_X1 U5088 ( .A1(n6268), .A2(n6267), .ZN(n7859) );
  OAI21_X1 U5089 ( .B1(n5759), .B2(n5758), .A(n5757), .ZN(n5777) );
  NAND2_X1 U5090 ( .A1(n6276), .A2(n6275), .ZN(n7628) );
  NAND2_X1 U5091 ( .A1(n5687), .A2(n5675), .ZN(n6956) );
  OAI211_X2 U5092 ( .C1(n4804), .C2(n4801), .A(n5705), .B(n4798), .ZN(n5759)
         );
  INV_X1 U5093 ( .A(n9412), .ZN(n4435) );
  INV_X2 U5094 ( .A(n9304), .ZN(n10139) );
  INV_X1 U5095 ( .A(n7138), .ZN(n7301) );
  INV_X1 U5096 ( .A(n10132), .ZN(n7954) );
  OAI21_X1 U5097 ( .B1(n4918), .B2(n5323), .A(n4917), .ZN(n7019) );
  AND2_X2 U5098 ( .A1(n7843), .A2(n9511), .ZN(n9394) );
  XNOR2_X1 U5099 ( .A(n5589), .B(n5588), .ZN(n6934) );
  AND2_X1 U5100 ( .A1(n6217), .A2(n6216), .ZN(n10201) );
  AND2_X2 U5101 ( .A1(n5510), .A2(n5509), .ZN(n7948) );
  INV_X1 U5102 ( .A(n9561), .ZN(n7947) );
  NAND2_X1 U5103 ( .A1(n6199), .A2(n4456), .ZN(n6207) );
  AND4_X1 U5104 ( .A1(n6230), .A2(n6229), .A3(n6228), .A4(n6227), .ZN(n7302)
         );
  CLKBUF_X1 U5105 ( .A(n6193), .Z(n8620) );
  INV_X1 U5106 ( .A(n7411), .ZN(n9448) );
  AND4_X1 U5107 ( .A1(n6273), .A2(n6272), .A3(n6271), .A4(n6270), .ZN(n7850)
         );
  OAI21_X1 U5109 ( .B1(n7065), .B2(n7064), .A(n7063), .ZN(n7274) );
  NAND4_X2 U5110 ( .A1(n5555), .A2(n5554), .A3(n5553), .A4(n5552), .ZN(n9558)
         );
  BUF_X1 U5111 ( .A(n6597), .Z(n6908) );
  AOI21_X1 U5112 ( .B1(n4984), .B2(n4982), .A(n4981), .ZN(n4980) );
  CLKBUF_X3 U5113 ( .A(n6222), .Z(n7967) );
  AND2_X1 U5114 ( .A1(n5756), .A2(n5755), .ZN(n5757) );
  AND2_X1 U5115 ( .A1(n5758), .A2(n4961), .ZN(n4959) );
  AND2_X2 U5116 ( .A1(n4669), .A2(n5465), .ZN(n5909) );
  NAND2_X1 U5117 ( .A1(n4802), .A2(n5686), .ZN(n4801) );
  NAND2_X1 U5118 ( .A1(n4946), .A2(n4458), .ZN(n4945) );
  CLKBUF_X1 U5119 ( .A(n6370), .Z(n8403) );
  INV_X1 U5120 ( .A(n6200), .ZN(n6287) );
  NAND2_X1 U5121 ( .A1(n4852), .A2(n4670), .ZN(n5467) );
  NOR2_X1 U5122 ( .A1(n5652), .A2(n4950), .ZN(n4943) );
  BUF_X1 U5123 ( .A(n9578), .Z(n4437) );
  NAND2_X1 U5124 ( .A1(n5462), .A2(n4853), .ZN(n4670) );
  NAND2_X1 U5125 ( .A1(n9075), .A2(n5352), .ZN(n6171) );
  NAND2_X1 U5126 ( .A1(n5618), .A2(SI_7_), .ZN(n5631) );
  OAI21_X1 U5127 ( .B1(n5778), .B2(n5565), .A(n5564), .ZN(n5566) );
  NAND2_X1 U5128 ( .A1(n4745), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5285) );
  NAND2_X1 U5129 ( .A1(n5778), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5564) );
  OR2_X1 U5130 ( .A1(n5274), .A2(n5246), .ZN(n5357) );
  AND3_X1 U5131 ( .A1(n5186), .A2(n5183), .A3(n5185), .ZN(n5274) );
  XNOR2_X1 U5132 ( .A(n5311), .B(P2_IR_REG_3__SCAN_IN), .ZN(n7159) );
  INV_X2 U5133 ( .A(n6929), .ZN(n5778) );
  INV_X1 U5134 ( .A(n5457), .ZN(n4684) );
  AND3_X1 U5135 ( .A1(n10400), .A2(n5762), .A3(n5451), .ZN(n5452) );
  BUF_X1 U5136 ( .A(n5308), .Z(n5412) );
  INV_X1 U5137 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5471) );
  NOR2_X1 U5138 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5237) );
  NOR2_X1 U5139 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5238) );
  BUF_X4 U5140 ( .A(P2_IR_REG_31__SCAN_IN), .Z(n5352) );
  INV_X1 U5141 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5476) );
  INV_X1 U5142 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6060) );
  NOR2_X1 U5143 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n4861) );
  NOR2_X1 U5144 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5455) );
  INV_X1 U5145 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6064) );
  NOR2_X1 U5146 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5236) );
  NOR2_X2 U5147 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5308) );
  INV_X1 U5148 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5070) );
  INV_X1 U5149 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5762) );
  INV_X4 U5150 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5151 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4436) );
  NOR2_X1 U5152 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5257) );
  INV_X4 U5153 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U5154 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5256) );
  AND2_X1 U5155 ( .A1(n6547), .A2(n6929), .ZN(n6200) );
  NAND2_X1 U5156 ( .A1(n9416), .A2(n7810), .ZN(n7809) );
  INV_X2 U5157 ( .A(n6632), .ZN(n6818) );
  NAND2_X1 U5158 ( .A1(n6632), .A2(n6646), .ZN(n6619) );
  NOR2_X2 U5159 ( .A1(n9179), .A2(n5853), .ZN(n4618) );
  XNOR2_X1 U5160 ( .A(n5475), .B(n5474), .ZN(n9578) );
  NAND2_X1 U5161 ( .A1(n9204), .A2(n7714), .ZN(n9323) );
  INV_X2 U5162 ( .A(n9204), .ZN(n4623) );
  NOR2_X2 U5163 ( .A1(n5418), .A2(n5419), .ZN(n7152) );
  NAND4_X4 U5164 ( .A1(n6214), .A2(n6215), .A3(n6213), .A4(n6212), .ZN(n6508)
         );
  NAND2_X1 U5165 ( .A1(n6541), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6215) );
  OR2_X1 U5166 ( .A1(n6544), .A2(n6211), .ZN(n6214) );
  AOI21_X2 U5167 ( .B1(n9321), .B2(n4505), .A(n4859), .ZN(n4858) );
  NOR2_X2 U5168 ( .A1(n6063), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n6066) );
  AND2_X2 U5169 ( .A1(n5208), .A2(n9815), .ZN(n9809) );
  NOR2_X2 U5170 ( .A1(n4985), .A2(n6101), .ZN(n5208) );
  AOI211_X2 U5171 ( .C1(n6163), .C2(n6147), .A(n9907), .B(n9680), .ZN(n9696)
         );
  INV_X1 U5172 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5242) );
  INV_X1 U5173 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5241) );
  AND2_X2 U5174 ( .A1(n9342), .A2(n9314), .ZN(n9321) );
  NAND2_X1 U5175 ( .A1(n6517), .A2(n4490), .ZN(n5120) );
  OR2_X1 U5176 ( .A1(n9061), .A2(n8081), .ZN(n8515) );
  OR2_X1 U5177 ( .A1(n7913), .A2(n7801), .ZN(n8507) );
  XNOR2_X1 U5178 ( .A(n8582), .B(n8607), .ZN(n8779) );
  AND2_X1 U5179 ( .A1(n9679), .A2(n9543), .ZN(n9524) );
  NAND2_X1 U5180 ( .A1(n9783), .A2(n5038), .ZN(n5034) );
  NOR2_X1 U5181 ( .A1(n5956), .A2(n5039), .ZN(n5038) );
  INV_X1 U5182 ( .A(n5935), .ZN(n5039) );
  INV_X1 U5183 ( .A(n8524), .ZN(n4565) );
  NAND2_X1 U5184 ( .A1(n4710), .A2(n6252), .ZN(n4709) );
  INV_X1 U5185 ( .A(n6251), .ZN(n4710) );
  OR2_X1 U5186 ( .A1(n8969), .A2(n8870), .ZN(n8533) );
  OR2_X1 U5187 ( .A1(n10040), .A2(n6130), .ZN(n6848) );
  AND2_X1 U5188 ( .A1(n4962), .A2(n4957), .ZN(n4956) );
  OR2_X1 U5189 ( .A1(n4957), .A2(n4960), .ZN(n4954) );
  OR2_X1 U5190 ( .A1(n4962), .A2(n5757), .ZN(n4955) );
  AND2_X1 U5191 ( .A1(n5757), .A2(n4961), .ZN(n4960) );
  INV_X1 U5192 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4796) );
  INV_X1 U5193 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4797) );
  OR2_X1 U5194 ( .A1(n8409), .A2(n8994), .ZN(n8583) );
  INV_X1 U5195 ( .A(n6174), .ZN(n6222) );
  NAND2_X1 U5196 ( .A1(n4880), .A2(n4879), .ZN(n5421) );
  INV_X1 U5197 ( .A(n7010), .ZN(n4775) );
  OR2_X1 U5198 ( .A1(n6588), .A2(n8606), .ZN(n8581) );
  OR2_X1 U5199 ( .A1(n6484), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8074) );
  NOR2_X1 U5200 ( .A1(n6424), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n4782) );
  NAND2_X1 U5201 ( .A1(n6193), .A2(n7239), .ZN(n8455) );
  NAND2_X1 U5202 ( .A1(n6192), .A2(n6191), .ZN(n8460) );
  OR2_X1 U5203 ( .A1(n6951), .A2(n6575), .ZN(n6877) );
  NAND2_X1 U5204 ( .A1(n4449), .A2(n8329), .ZN(n8547) );
  OR2_X1 U5205 ( .A1(n8329), .A2(n4449), .ZN(n8554) );
  OR2_X1 U5206 ( .A1(n8261), .A2(n8826), .ZN(n8546) );
  AND2_X1 U5207 ( .A1(n7134), .A2(n7131), .ZN(n7077) );
  AND2_X1 U5208 ( .A1(n5412), .A2(n4576), .ZN(n5183) );
  AND2_X1 U5209 ( .A1(n4746), .A2(n5243), .ZN(n4576) );
  INV_X1 U5210 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U5211 ( .A1(n10056), .A2(n5467), .ZN(n5836) );
  OR2_X1 U5212 ( .A1(n8118), .A2(n9718), .ZN(n9497) );
  INV_X1 U5213 ( .A(n9323), .ZN(n4859) );
  NAND2_X1 U5214 ( .A1(n5511), .A2(n9559), .ZN(n9451) );
  NAND2_X1 U5215 ( .A1(n9560), .A2(n10132), .ZN(n9450) );
  INV_X1 U5216 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4704) );
  AND2_X1 U5217 ( .A1(n6025), .A2(n6011), .ZN(n6023) );
  NAND2_X1 U5218 ( .A1(n4546), .A2(n4478), .ZN(n6006) );
  NAND2_X1 U5219 ( .A1(n5985), .A2(n5225), .ZN(n4546) );
  INV_X1 U5220 ( .A(n5986), .ZN(n4545) );
  AND2_X1 U5221 ( .A1(n6007), .A2(n5990), .ZN(n6005) );
  AOI22_X1 U5222 ( .A1(n4973), .A2(n4974), .B1(n4975), .B2(n4977), .ZN(n4971)
         );
  INV_X1 U5223 ( .A(n4980), .ZN(n4977) );
  NAND2_X1 U5224 ( .A1(n5865), .A2(n5864), .ZN(n5885) );
  OAI21_X1 U5225 ( .B1(n5087), .B2(n10046), .A(n5088), .ZN(n5875) );
  AOI21_X1 U5226 ( .B1(n5090), .B2(P1_IR_REG_31__SCAN_IN), .A(
        P1_IR_REG_17__SCAN_IN), .ZN(n5088) );
  NAND2_X1 U5227 ( .A1(n5861), .A2(SI_18_), .ZN(n5862) );
  NAND2_X1 U5228 ( .A1(n5751), .A2(n5753), .ZN(n5758) );
  AND2_X1 U5229 ( .A1(n4579), .A2(n5673), .ZN(n4804) );
  AOI21_X1 U5230 ( .B1(n8280), .B2(n5164), .A(n5167), .ZN(n5163) );
  INV_X1 U5231 ( .A(n5168), .ZN(n5164) );
  AND2_X1 U5232 ( .A1(n7976), .A2(n7975), .ZN(n8772) );
  AND2_X1 U5233 ( .A1(n7096), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6576) );
  AND2_X1 U5234 ( .A1(n6891), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4895) );
  NAND2_X1 U5235 ( .A1(n4757), .A2(n4761), .ZN(n4756) );
  INV_X1 U5236 ( .A(n4759), .ZN(n4757) );
  AOI21_X1 U5237 ( .B1(n5395), .B2(n5394), .A(n4760), .ZN(n4759) );
  INV_X1 U5238 ( .A(n8677), .ZN(n4760) );
  AND2_X1 U5239 ( .A1(n6366), .A2(n6365), .ZN(n8882) );
  AND2_X1 U5240 ( .A1(n5125), .A2(n8412), .ZN(n5124) );
  NAND2_X1 U5241 ( .A1(n5128), .A2(n5126), .ZN(n5125) );
  NAND2_X1 U5242 ( .A1(n6308), .A2(n5235), .ZN(n5064) );
  INV_X1 U5243 ( .A(n9074), .ZN(n7073) );
  NAND2_X1 U5244 ( .A1(n8073), .A2(n10198), .ZN(n6558) );
  NOR2_X1 U5245 ( .A1(n4457), .A2(n5061), .ZN(n5060) );
  OR2_X1 U5246 ( .A1(n9007), .A2(n8815), .ZN(n8560) );
  NAND2_X1 U5247 ( .A1(n5069), .A2(n5068), .ZN(n4731) );
  AND2_X1 U5248 ( .A1(n6432), .A2(n5223), .ZN(n5068) );
  NOR2_X1 U5249 ( .A1(n5102), .A2(n4495), .ZN(n5100) );
  NAND2_X1 U5250 ( .A1(n4743), .A2(n4741), .ZN(n7909) );
  NOR2_X1 U5251 ( .A1(n8425), .A2(n4742), .ZN(n4741) );
  INV_X1 U5252 ( .A(n6320), .ZN(n4742) );
  NOR2_X1 U5253 ( .A1(n6878), .A2(n6883), .ZN(n7107) );
  AND2_X1 U5254 ( .A1(n7097), .A2(n6576), .ZN(n7108) );
  NAND2_X1 U5255 ( .A1(n6068), .A2(n9447), .ZN(n9529) );
  NAND2_X1 U5256 ( .A1(n4689), .A2(n4690), .ZN(n9398) );
  AOI21_X1 U5257 ( .B1(n4942), .B2(n4940), .A(n9514), .ZN(n4690) );
  NOR2_X1 U5258 ( .A1(n5232), .A2(n4941), .ZN(n4940) );
  CLKBUF_X1 U5259 ( .A(n5836), .Z(n5837) );
  NAND2_X1 U5260 ( .A1(n4841), .A2(n4840), .ZN(n4839) );
  NAND2_X1 U5261 ( .A1(n9616), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4840) );
  NOR2_X1 U5262 ( .A1(n7656), .A2(n7655), .ZN(n8202) );
  NAND2_X1 U5263 ( .A1(n4844), .A2(n4843), .ZN(n9668) );
  AOI21_X1 U5264 ( .B1(n4845), .B2(n9637), .A(n4533), .ZN(n4843) );
  INV_X1 U5265 ( .A(n6016), .ZN(n6014) );
  AND2_X1 U5266 ( .A1(n9501), .A2(n9380), .ZN(n9403) );
  AOI21_X1 U5267 ( .B1(n5025), .B2(n5028), .A(n4494), .ZN(n5023) );
  INV_X1 U5268 ( .A(n6004), .ZN(n5028) );
  NOR2_X1 U5269 ( .A1(n9754), .A2(n5035), .ZN(n5033) );
  NAND2_X1 U5270 ( .A1(n7661), .A2(n5665), .ZN(n7705) );
  AND2_X1 U5271 ( .A1(n6135), .A2(n10042), .ZN(n7732) );
  NAND2_X1 U5272 ( .A1(n4804), .A2(n4803), .ZN(n5687) );
  NAND2_X1 U5273 ( .A1(n6483), .A2(n6482), .ZN(n8582) );
  NAND2_X1 U5274 ( .A1(n6479), .A2(n6478), .ZN(n8781) );
  NOR2_X1 U5275 ( .A1(n7270), .A2(n7269), .ZN(n7268) );
  NOR2_X1 U5276 ( .A1(n8155), .A2(n9907), .ZN(n9675) );
  NAND2_X1 U5277 ( .A1(n8464), .A2(n8577), .ZN(n4591) );
  AND2_X1 U5278 ( .A1(n9465), .A2(n9348), .ZN(n4679) );
  INV_X1 U5279 ( .A(n4679), .ZN(n4678) );
  AND2_X1 U5280 ( .A1(n8505), .A2(n8507), .ZN(n4813) );
  NOR2_X1 U5281 ( .A1(n9483), .A2(n4590), .ZN(n4589) );
  AND2_X1 U5282 ( .A1(n8905), .A2(n8517), .ZN(n4594) );
  AOI21_X1 U5283 ( .B1(n4821), .B2(n8530), .A(n4820), .ZN(n4819) );
  INV_X1 U5284 ( .A(n8533), .ZN(n4820) );
  OR2_X1 U5285 ( .A1(n8524), .A2(n8531), .ZN(n4821) );
  NAND2_X1 U5286 ( .A1(n8529), .A2(n4567), .ZN(n4828) );
  NOR2_X1 U5287 ( .A1(n4568), .A2(n8570), .ZN(n4567) );
  INV_X1 U5288 ( .A(n8539), .ZN(n4568) );
  NAND2_X1 U5289 ( .A1(n4638), .A2(n9381), .ZN(n4637) );
  NAND2_X1 U5290 ( .A1(n9386), .A2(n9492), .ZN(n4667) );
  OR2_X1 U5291 ( .A1(n9387), .A2(n9394), .ZN(n4665) );
  NAND2_X1 U5292 ( .A1(n9380), .A2(n9379), .ZN(n9388) );
  AND2_X1 U5293 ( .A1(n9988), .A2(n9867), .ZN(n5842) );
  AND2_X1 U5294 ( .A1(n4980), .A2(SI_20_), .ZN(n4978) );
  NAND2_X1 U5295 ( .A1(n5757), .A2(n5758), .ZN(n4963) );
  NAND2_X1 U5296 ( .A1(n5160), .A2(n5161), .ZN(n5159) );
  INV_X1 U5297 ( .A(n8350), .ZN(n5161) );
  NAND2_X1 U5298 ( .A1(n5165), .A2(n5163), .ZN(n5160) );
  NAND2_X1 U5299 ( .A1(n7124), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4916) );
  INV_X1 U5300 ( .A(n6252), .ZN(n4711) );
  AND2_X1 U5301 ( .A1(n8585), .A2(n8587), .ZN(n6577) );
  NAND2_X1 U5302 ( .A1(n4660), .A2(n9392), .ZN(n9395) );
  NAND2_X1 U5303 ( .A1(n4662), .A2(n4661), .ZN(n4660) );
  NAND2_X1 U5304 ( .A1(n4668), .A2(n4663), .ZN(n4662) );
  NOR2_X1 U5305 ( .A1(n5767), .A2(n5766), .ZN(n4617) );
  NAND2_X1 U5306 ( .A1(n5964), .A2(n5963), .ZN(n5986) );
  AOI21_X1 U5307 ( .B1(n4978), .B2(n4976), .A(n5900), .ZN(n4973) );
  AOI21_X1 U5308 ( .B1(n4980), .B2(n4976), .A(SI_20_), .ZN(n4975) );
  NAND2_X1 U5309 ( .A1(n8144), .A2(n10442), .ZN(n4645) );
  OAI21_X1 U5310 ( .B1(n8144), .B2(n4634), .A(n4633), .ZN(n5703) );
  NAND2_X1 U5311 ( .A1(n8144), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n4633) );
  NOR2_X1 U5312 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5633) );
  INV_X1 U5313 ( .A(n8092), .ZN(n5156) );
  INV_X1 U5314 ( .A(n5158), .ZN(n5157) );
  OAI21_X1 U5315 ( .B1(n5159), .B2(n5163), .A(n8348), .ZN(n5158) );
  INV_X1 U5316 ( .A(n5179), .ZN(n5178) );
  AOI21_X1 U5317 ( .B1(n4805), .B2(n8568), .A(n4646), .ZN(n8579) );
  NAND2_X1 U5318 ( .A1(n8581), .A2(n8574), .ZN(n4646) );
  AND2_X1 U5319 ( .A1(n8578), .A2(n8583), .ZN(n4823) );
  OR2_X1 U5320 ( .A1(n6223), .A2(n7172), .ZN(n6197) );
  NAND2_X1 U5321 ( .A1(n4883), .A2(n4496), .ZN(n4881) );
  OR2_X1 U5322 ( .A1(n8637), .A2(n10545), .ZN(n5427) );
  OR2_X1 U5323 ( .A1(n5330), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5298) );
  NOR2_X1 U5324 ( .A1(n6895), .A2(n4929), .ZN(n5341) );
  NOR2_X1 U5325 ( .A1(n6310), .A2(n7803), .ZN(n4929) );
  NOR2_X1 U5326 ( .A1(n8673), .A2(n8695), .ZN(n4910) );
  NAND2_X1 U5327 ( .A1(n4913), .A2(n4915), .ZN(n4908) );
  NAND2_X1 U5328 ( .A1(n8710), .A2(n4570), .ZN(n5349) );
  NAND2_X1 U5329 ( .A1(n4571), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4570) );
  AND2_X1 U5330 ( .A1(n10383), .A2(n4793), .ZN(n4792) );
  INV_X1 U5331 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n4793) );
  INV_X1 U5332 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10383) );
  INV_X1 U5333 ( .A(n6344), .ZN(n6343) );
  NOR2_X1 U5334 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n4790) );
  INV_X1 U5335 ( .A(n6314), .ZN(n6313) );
  NAND2_X1 U5336 ( .A1(n8451), .A2(n8452), .ZN(n4580) );
  NOR2_X1 U5337 ( .A1(n8483), .A2(n5134), .ZN(n5133) );
  INV_X1 U5338 ( .A(n8494), .ZN(n5134) );
  AND2_X1 U5339 ( .A1(n5140), .A2(n8496), .ZN(n5139) );
  INV_X1 U5340 ( .A(n8491), .ZN(n5141) );
  AND2_X1 U5341 ( .A1(n6507), .A2(n8462), .ZN(n7163) );
  INV_X1 U5342 ( .A(n8821), .ZN(n4725) );
  NOR2_X1 U5343 ( .A1(n4726), .A2(n4725), .ZN(n4723) );
  INV_X1 U5344 ( .A(n6401), .ZN(n4726) );
  AOI21_X1 U5345 ( .B1(n6401), .B2(n6402), .A(n4728), .ZN(n4727) );
  AND2_X1 U5346 ( .A1(n8410), .A2(n5051), .ZN(n5050) );
  NAND2_X1 U5347 ( .A1(n5052), .A2(n6349), .ZN(n5051) );
  INV_X1 U5348 ( .A(n6349), .ZN(n5053) );
  AND2_X1 U5349 ( .A1(n5050), .A2(n4717), .ZN(n4716) );
  NAND2_X1 U5350 ( .A1(n4718), .A2(n6340), .ZN(n4717) );
  INV_X1 U5351 ( .A(n6339), .ZN(n4718) );
  NAND2_X1 U5352 ( .A1(n4716), .A2(n4719), .ZN(n4714) );
  INV_X1 U5353 ( .A(n6340), .ZN(n4719) );
  NOR2_X1 U5354 ( .A1(n5260), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n5261) );
  OR2_X1 U5355 ( .A1(n5324), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5327) );
  INV_X1 U5356 ( .A(n9228), .ZN(n5078) );
  NAND2_X1 U5357 ( .A1(n4695), .A2(n6787), .ZN(n9129) );
  NOR2_X1 U5359 ( .A1(n4701), .A2(n4499), .ZN(n4700) );
  INV_X1 U5360 ( .A(n6748), .ZN(n4701) );
  OR2_X1 U5361 ( .A1(n9950), .A2(n9771), .ZN(n9444) );
  OR2_X1 U5362 ( .A1(n9957), .A2(n9231), .ZN(n9369) );
  NAND2_X1 U5363 ( .A1(n4618), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5892) );
  OR2_X1 U5364 ( .A1(n9988), .A2(n9855), .ZN(n9478) );
  NAND2_X1 U5365 ( .A1(n4617), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5810) );
  OAI21_X1 U5366 ( .B1(n9419), .B2(n5009), .A(n5702), .ZN(n5008) );
  INV_X1 U5367 ( .A(n5008), .ZN(n5007) );
  NAND2_X1 U5368 ( .A1(n5657), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5696) );
  INV_X1 U5369 ( .A(n5659), .ZN(n5657) );
  AOI21_X1 U5370 ( .B1(n4441), .B2(n5011), .A(n4497), .ZN(n5010) );
  NAND2_X1 U5371 ( .A1(n6142), .A2(n6141), .ZN(n8136) );
  NAND2_X1 U5372 ( .A1(n6138), .A2(n6137), .ZN(n6142) );
  AND2_X1 U5373 ( .A1(n6039), .A2(n6029), .ZN(n6037) );
  INV_X1 U5374 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5454) );
  OR2_X1 U5375 ( .A1(n5957), .A2(n5959), .ZN(n5982) );
  XNOR2_X1 U5376 ( .A(n6067), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6593) );
  OR2_X1 U5377 ( .A1(n6066), .A2(n10046), .ZN(n6067) );
  NAND2_X1 U5378 ( .A1(n5831), .A2(n5830), .ZN(n5843) );
  INV_X1 U5379 ( .A(n5859), .ZN(n4984) );
  XNOR2_X1 U5380 ( .A(n5860), .B(SI_18_), .ZN(n5859) );
  AND2_X1 U5381 ( .A1(n4953), .A2(n5759), .ZN(n4639) );
  NAND2_X1 U5382 ( .A1(n4952), .A2(n5819), .ZN(n4951) );
  INV_X1 U5383 ( .A(n5631), .ZN(n4950) );
  NAND2_X1 U5384 ( .A1(n4945), .A2(n4948), .ZN(n4803) );
  XNOR2_X1 U5385 ( .A(n5666), .B(n10418), .ZN(n5667) );
  AND2_X1 U5386 ( .A1(n5613), .A2(n5614), .ZN(n4540) );
  OAI211_X1 U5387 ( .C1(n4969), .C2(P2_DATAO_REG_1__SCAN_IN), .A(n4966), .B(
        n4964), .ZN(n5480) );
  NAND2_X1 U5388 ( .A1(n4965), .A2(n4970), .ZN(n4964) );
  INV_X1 U5389 ( .A(n4968), .ZN(n4965) );
  INV_X1 U5390 ( .A(n7552), .ZN(n5169) );
  XNOR2_X1 U5391 ( .A(n7258), .B(n6204), .ZN(n7259) );
  INV_X1 U5392 ( .A(n8099), .ZN(n5175) );
  INV_X1 U5393 ( .A(n8381), .ZN(n5172) );
  NAND2_X1 U5394 ( .A1(n7139), .A2(n8620), .ZN(n5147) );
  NAND2_X1 U5395 ( .A1(n7140), .A2(n7167), .ZN(n7143) );
  NOR2_X1 U5396 ( .A1(n7856), .A2(n5180), .ZN(n5179) );
  INV_X1 U5397 ( .A(n7853), .ZN(n5180) );
  NAND2_X1 U5398 ( .A1(n8280), .A2(n5166), .ZN(n5165) );
  INV_X1 U5399 ( .A(n8340), .ZN(n5166) );
  INV_X1 U5400 ( .A(n5149), .ZN(n5148) );
  OAI21_X1 U5401 ( .B1(n7306), .B2(n5151), .A(n7345), .ZN(n5149) );
  OAI21_X1 U5402 ( .B1(n8439), .B2(n8438), .A(n8437), .ZN(n8441) );
  NAND2_X1 U5403 ( .A1(n8439), .A2(n5214), .ZN(n8437) );
  AND3_X1 U5404 ( .A1(n5356), .A2(n6501), .A3(n5244), .ZN(n5245) );
  NAND2_X1 U5405 ( .A1(n6495), .A2(n6494), .ZN(n7976) );
  NAND4_X1 U5406 ( .A1(n6176), .A2(n6179), .A3(n6177), .A4(n6178), .ZN(n6193)
         );
  NAND4_X1 U5407 ( .A1(n6187), .A2(n6188), .A3(n6189), .A4(n6186), .ZN(n6505)
         );
  NAND2_X1 U5408 ( .A1(n6183), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U5409 ( .A1(n5412), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4903) );
  NAND2_X1 U5410 ( .A1(n4922), .A2(n6985), .ZN(n4920) );
  AND2_X1 U5411 ( .A1(n5309), .A2(n7159), .ZN(n4922) );
  NAND2_X1 U5412 ( .A1(n5419), .A2(n4884), .ZN(n4883) );
  AOI21_X1 U5413 ( .B1(n4772), .B2(n4774), .A(n4770), .ZN(n4769) );
  INV_X1 U5414 ( .A(n7392), .ZN(n4770) );
  INV_X1 U5415 ( .A(n6915), .ZN(n4766) );
  INV_X1 U5416 ( .A(n6916), .ZN(n4767) );
  OR2_X1 U5417 ( .A1(n6310), .A2(n10328), .ZN(n5430) );
  NOR2_X1 U5418 ( .A1(n8646), .A2(n8647), .ZN(n8665) );
  OAI21_X1 U5419 ( .B1(n8665), .B2(n8664), .A(n8663), .ZN(n8662) );
  NAND2_X1 U5420 ( .A1(n4754), .A2(n4749), .ZN(n4748) );
  INV_X1 U5421 ( .A(n8690), .ZN(n4749) );
  NAND2_X1 U5422 ( .A1(n6899), .A2(n4752), .ZN(n4755) );
  NAND2_X1 U5423 ( .A1(n5349), .A2(n8731), .ZN(n5351) );
  OR2_X1 U5424 ( .A1(n5349), .A2(n8731), .ZN(n5350) );
  OAI22_X1 U5425 ( .A1(n6491), .A2(n5057), .B1(n8182), .B2(n8998), .ZN(n5056)
         );
  NAND2_X1 U5426 ( .A1(n5059), .A2(n8569), .ZN(n5057) );
  NOR2_X1 U5427 ( .A1(n6491), .A2(n8573), .ZN(n5058) );
  INV_X1 U5428 ( .A(n6557), .ZN(n6533) );
  NAND2_X1 U5429 ( .A1(n6556), .A2(n6555), .ZN(n8397) );
  OR2_X1 U5430 ( .A1(n6458), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6472) );
  NAND2_X1 U5431 ( .A1(n4782), .A2(n6435), .ZN(n6448) );
  OR2_X1 U5432 ( .A1(n6383), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U5433 ( .A1(n5129), .A2(n5135), .ZN(n5128) );
  NOR2_X1 U5434 ( .A1(n8450), .A2(n5131), .ZN(n5130) );
  INV_X1 U5435 ( .A(n4580), .ZN(n8412) );
  AND4_X1 U5436 ( .A1(n6328), .A2(n6327), .A3(n6326), .A4(n6325), .ZN(n7801)
         );
  NAND2_X1 U5437 ( .A1(n6513), .A2(n6512), .ZN(n6514) );
  NAND2_X1 U5438 ( .A1(n5106), .A2(n8490), .ZN(n5105) );
  NAND2_X1 U5439 ( .A1(n5045), .A2(n5044), .ZN(n7456) );
  AOI21_X1 U5440 ( .B1(n8415), .B2(n5047), .A(n4460), .ZN(n5044) );
  INV_X1 U5441 ( .A(n10163), .ZN(n5047) );
  NOR2_X1 U5442 ( .A1(n4473), .A2(n4730), .ZN(n4729) );
  INV_X1 U5443 ( .A(n6443), .ZN(n4730) );
  INV_X1 U5444 ( .A(n8781), .ZN(n8793) );
  NAND2_X1 U5445 ( .A1(n6493), .A2(n6492), .ZN(n6588) );
  INV_X1 U5446 ( .A(n8783), .ZN(n4737) );
  INV_X1 U5447 ( .A(n8563), .ZN(n8790) );
  NAND2_X1 U5448 ( .A1(n6434), .A2(n6433), .ZN(n8329) );
  INV_X1 U5449 ( .A(n5113), .ZN(n5112) );
  OAI21_X1 U5450 ( .B1(n5115), .B2(n5114), .A(n8546), .ZN(n5113) );
  AND2_X1 U5451 ( .A1(n8554), .A2(n8547), .ZN(n8812) );
  AND2_X1 U5452 ( .A1(n6419), .A2(n6418), .ZN(n8543) );
  NOR2_X1 U5453 ( .A1(n6525), .A2(n5116), .ZN(n5115) );
  INV_X1 U5454 ( .A(n8541), .ZN(n5116) );
  AOI21_X1 U5455 ( .B1(n8842), .B2(n6494), .A(n6409), .ZN(n8854) );
  AND2_X1 U5456 ( .A1(n6430), .A2(n6429), .ZN(n8826) );
  OR2_X1 U5457 ( .A1(n9028), .A2(n8854), .ZN(n8541) );
  AND2_X1 U5458 ( .A1(n6518), .A2(n8523), .ZN(n5119) );
  INV_X1 U5459 ( .A(n8410), .ZN(n8905) );
  NAND2_X1 U5460 ( .A1(n4715), .A2(n6340), .ZN(n8914) );
  NAND2_X1 U5461 ( .A1(n8924), .A2(n6339), .ZN(n4715) );
  AND2_X1 U5462 ( .A1(n8577), .A2(n7127), .ZN(n10167) );
  INV_X1 U5463 ( .A(n8881), .ZN(n10168) );
  OR2_X1 U5464 ( .A1(n8570), .A2(n7127), .ZN(n8881) );
  NAND2_X1 U5465 ( .A1(n5064), .A2(n5063), .ZN(n4743) );
  AND2_X1 U5466 ( .A1(n4477), .A2(n6309), .ZN(n5063) );
  AND2_X1 U5467 ( .A1(n6884), .A2(n7073), .ZN(n7105) );
  NAND2_X1 U5468 ( .A1(n5275), .A2(n5352), .ZN(n6502) );
  INV_X1 U5469 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6501) );
  NAND2_X1 U5470 ( .A1(n5304), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U5471 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5306) );
  NAND2_X1 U5472 ( .A1(n6132), .A2(n6116), .ZN(n6597) );
  AND2_X1 U5473 ( .A1(n6118), .A2(n6117), .ZN(n6116) );
  AOI21_X1 U5474 ( .B1(n5082), .B2(n5085), .A(n4492), .ZN(n5079) );
  INV_X1 U5475 ( .A(n6712), .ZN(n5085) );
  OR2_X1 U5476 ( .A1(n5948), .A2(n5947), .ZN(n5971) );
  XNOR2_X1 U5477 ( .A(n6604), .B(n6841), .ZN(n6605) );
  AOI21_X1 U5478 ( .B1(n7411), .B2(n6818), .A(n6598), .ZN(n6606) );
  OR2_X1 U5479 ( .A1(n5892), .A2(n5891), .ZN(n5907) );
  CLKBUF_X1 U5480 ( .A(n9129), .Z(n9130) );
  NAND2_X1 U5481 ( .A1(n7398), .A2(n6643), .ZN(n6648) );
  OR2_X1 U5482 ( .A1(n6862), .A2(n10269), .ZN(n6858) );
  INV_X1 U5483 ( .A(n9529), .ZN(n7028) );
  INV_X1 U5484 ( .A(n6858), .ZN(n6866) );
  XNOR2_X1 U5485 ( .A(n6065), .B(n6064), .ZN(n6592) );
  NAND2_X1 U5486 ( .A1(n4544), .A2(n4543), .ZN(n4542) );
  INV_X1 U5487 ( .A(n9543), .ZN(n4543) );
  INV_X1 U5488 ( .A(n7035), .ZN(n4838) );
  AOI21_X1 U5489 ( .B1(n7274), .B2(n7273), .A(n7272), .ZN(n7292) );
  NOR2_X1 U5490 ( .A1(n7652), .A2(n4530), .ZN(n7656) );
  XNOR2_X1 U5491 ( .A(n8195), .B(n9628), .ZN(n9624) );
  INV_X1 U5492 ( .A(n4842), .ZN(n8204) );
  AND2_X1 U5493 ( .A1(n9653), .A2(n8207), .ZN(n4845) );
  OR2_X1 U5494 ( .A1(n9638), .A2(n9637), .ZN(n9635) );
  OR2_X1 U5495 ( .A1(n9666), .A2(n8210), .ZN(n8211) );
  OR2_X1 U5496 ( .A1(n6045), .A2(n6044), .ZN(n9693) );
  INV_X1 U5497 ( .A(n9701), .ZN(n9698) );
  AOI21_X1 U5498 ( .B1(n9708), .B2(n6047), .A(n6035), .ZN(n9718) );
  NAND2_X1 U5499 ( .A1(n5036), .A2(n5955), .ZN(n5035) );
  OR2_X1 U5500 ( .A1(n5037), .A2(n5956), .ZN(n5036) );
  NAND2_X1 U5501 ( .A1(n5936), .A2(n5935), .ZN(n5037) );
  OR2_X1 U5502 ( .A1(n9966), .A2(n9821), .ZN(n5916) );
  NAND2_X1 U5503 ( .A1(n8220), .A2(n9478), .ZN(n9853) );
  AND2_X1 U5504 ( .A1(n4441), .A2(n5774), .ZN(n5017) );
  NOR2_X1 U5505 ( .A1(n9883), .A2(n5816), .ZN(n9880) );
  NAND2_X1 U5506 ( .A1(n7862), .A2(n6078), .ZN(n9911) );
  CLKBUF_X1 U5507 ( .A(n9887), .Z(n9889) );
  INV_X1 U5508 ( .A(n9419), .ZN(n4854) );
  NAND2_X1 U5509 ( .A1(n7490), .A2(n9424), .ZN(n9460) );
  NAND2_X1 U5510 ( .A1(n7705), .A2(n9419), .ZN(n7704) );
  INV_X1 U5511 ( .A(n7615), .ZN(n5030) );
  INV_X1 U5512 ( .A(n9915), .ZN(n9898) );
  INV_X1 U5513 ( .A(n9913), .ZN(n9896) );
  OR2_X1 U5514 ( .A1(n6070), .A2(n7737), .ZN(n7814) );
  AND2_X1 U5515 ( .A1(n7028), .A2(n7030), .ZN(n9915) );
  AND2_X1 U5516 ( .A1(n8159), .A2(n9543), .ZN(n9932) );
  NAND2_X1 U5517 ( .A1(n6013), .A2(n6012), .ZN(n9723) );
  OAI21_X1 U5518 ( .B1(n5543), .B2(n4698), .A(n4696), .ZN(n4699) );
  NAND2_X1 U5519 ( .A1(n5543), .A2(n4697), .ZN(n4696) );
  AND2_X1 U5520 ( .A1(n7337), .A2(n9534), .ZN(n10148) );
  NOR2_X1 U5521 ( .A1(n7730), .A2(n6134), .ZN(n6166) );
  NAND2_X1 U5522 ( .A1(n6120), .A2(n6132), .ZN(n10040) );
  XNOR2_X1 U5523 ( .A(n6038), .B(n6037), .ZN(n9086) );
  NOR2_X1 U5524 ( .A1(n5919), .A2(SI_21_), .ZN(n5921) );
  INV_X1 U5525 ( .A(n5886), .ZN(n4983) );
  OAI211_X1 U5526 ( .C1(n5875), .C2(n5874), .A(n5873), .B(n5872), .ZN(n6594)
         );
  NAND2_X1 U5527 ( .A1(n5875), .A2(n4846), .ZN(n5873) );
  NAND2_X1 U5528 ( .A1(n5803), .A2(n5091), .ZN(n5090) );
  INV_X1 U5529 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5091) );
  NAND2_X1 U5530 ( .A1(n5632), .A2(n4943), .ZN(n4949) );
  OAI211_X1 U5531 ( .C1(n5584), .C2(P1_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n4541), .ZN(n5536) );
  INV_X1 U5532 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4651) );
  AND3_X1 U5533 ( .A1(n6348), .A2(n6347), .A3(n6346), .ZN(n8081) );
  NAND2_X1 U5534 ( .A1(n7144), .A2(n7145), .ZN(n7261) );
  INV_X1 U5535 ( .A(n5192), .ZN(n5191) );
  OAI22_X1 U5536 ( .A1(n4455), .A2(n5193), .B1(n8085), .B2(n8899), .ZN(n5192)
         );
  NAND2_X1 U5537 ( .A1(n5145), .A2(n7142), .ZN(n5146) );
  NAND2_X1 U5538 ( .A1(n7301), .A2(n7141), .ZN(n5145) );
  NAND2_X1 U5539 ( .A1(n5147), .A2(n7143), .ZN(n7236) );
  INV_X1 U5540 ( .A(n10179), .ZN(n10211) );
  AND4_X1 U5541 ( .A1(n6250), .A2(n6249), .A3(n6248), .A4(n6247), .ZN(n7555)
         );
  AND2_X1 U5542 ( .A1(n6399), .A2(n6398), .ZN(n8880) );
  AND3_X1 U5543 ( .A1(n6338), .A2(n6337), .A3(n6336), .ZN(n8056) );
  AND2_X1 U5544 ( .A1(n7110), .A2(n7109), .ZN(n8375) );
  AND2_X1 U5545 ( .A1(n6454), .A2(n6453), .ZN(n8815) );
  INV_X1 U5546 ( .A(n8373), .ZN(n8392) );
  INV_X1 U5547 ( .A(n8375), .ZN(n8395) );
  INV_X1 U5548 ( .A(n8815), .ZN(n8608) );
  INV_X1 U5549 ( .A(n4449), .ZN(n8801) );
  INV_X1 U5550 ( .A(n8882), .ZN(n8907) );
  CLKBUF_X1 U5551 ( .A(n6207), .Z(n8619) );
  OR2_X1 U5552 ( .A1(n5374), .A2(n5320), .ZN(n4777) );
  OR2_X1 U5553 ( .A1(n7178), .A2(n7177), .ZN(n4776) );
  INV_X1 U5554 ( .A(n8718), .ZN(n8755) );
  XNOR2_X1 U5555 ( .A(n5344), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8671) );
  AND2_X1 U5556 ( .A1(n4536), .A2(n4888), .ZN(n4886) );
  NAND2_X1 U5557 ( .A1(n4888), .A2(n4892), .ZN(n4887) );
  AOI21_X1 U5558 ( .B1(n8718), .B2(n8596), .A(n5410), .ZN(n4779) );
  XNOR2_X1 U5559 ( .A(n4781), .B(n5408), .ZN(n4780) );
  INV_X1 U5560 ( .A(n5407), .ZN(n4781) );
  NAND2_X1 U5561 ( .A1(n6423), .A2(n6422), .ZN(n8261) );
  INV_X1 U5562 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10293) );
  NAND2_X1 U5563 ( .A1(n4443), .A2(n6558), .ZN(n4788) );
  AND2_X1 U5564 ( .A1(n6289), .A2(n6288), .ZN(n7892) );
  AND2_X1 U5565 ( .A1(n6553), .A2(n5067), .ZN(n4657) );
  INV_X1 U5566 ( .A(n6588), .ZN(n8076) );
  INV_X1 U5567 ( .A(n8582), .ZN(n8998) );
  NOR2_X1 U5568 ( .A1(n4740), .A2(n4735), .ZN(n4734) );
  OR2_X1 U5569 ( .A1(n4737), .A2(n10229), .ZN(n4735) );
  NAND2_X1 U5570 ( .A1(n4732), .A2(n10171), .ZN(n4738) );
  INV_X1 U5571 ( .A(n8779), .ZN(n4736) );
  OR2_X1 U5572 ( .A1(n10229), .A2(n10223), .ZN(n9045) );
  XNOR2_X1 U5573 ( .A(n6107), .B(n6106), .ZN(n7029) );
  OR2_X1 U5574 ( .A1(n6956), .A2(n5676), .ZN(n5680) );
  OR2_X1 U5575 ( .A1(n8151), .A2(n6941), .ZN(n5495) );
  NAND2_X1 U5576 ( .A1(n5992), .A2(n5991), .ZN(n9741) );
  NAND2_X1 U5577 ( .A1(n6002), .A2(n6001), .ZN(n9750) );
  NAND4_X2 U5578 ( .A1(n5530), .A2(n5529), .A3(n5528), .A4(n5527), .ZN(n9561)
         );
  NAND2_X1 U5579 ( .A1(n5551), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5527) );
  OR2_X1 U5580 ( .A1(n7268), .A2(n4470), .ZN(n4837) );
  AND2_X1 U5581 ( .A1(n4837), .A2(n4836), .ZN(n10066) );
  INV_X1 U5582 ( .A(n7282), .ZN(n4836) );
  NOR2_X1 U5583 ( .A1(n9633), .A2(n9632), .ZN(n9631) );
  INV_X1 U5584 ( .A(n5803), .ZN(n5089) );
  INV_X1 U5585 ( .A(n10090), .ZN(n9663) );
  OR2_X1 U5586 ( .A1(n7118), .A2(n7030), .ZN(n10088) );
  OAI21_X1 U5587 ( .B1(n10098), .B2(n8215), .A(n9123), .ZN(n4831) );
  INV_X1 U5588 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8215) );
  XNOR2_X1 U5589 ( .A(n4574), .B(n4661), .ZN(n9690) );
  NAND2_X1 U5590 ( .A1(n9688), .A2(n9687), .ZN(n4574) );
  INV_X1 U5591 ( .A(n9926), .ZN(n10119) );
  INV_X1 U5592 ( .A(n7727), .ZN(n9948) );
  AND2_X1 U5593 ( .A1(n10161), .A2(n10148), .ZN(n7727) );
  AOI21_X2 U5594 ( .B1(n10044), .B2(n5505), .A(n8148), .ZN(n9679) );
  INV_X1 U5595 ( .A(n8241), .ZN(n4647) );
  INV_X1 U5596 ( .A(n8247), .ZN(n4649) );
  INV_X1 U5597 ( .A(n8118), .ZN(n10018) );
  INV_X1 U5598 ( .A(n9723), .ZN(n10022) );
  NAND2_X1 U5599 ( .A1(n10155), .A2(n10148), .ZN(n10026) );
  NOR2_X1 U5600 ( .A1(n8022), .A2(n8021), .ZN(n10590) );
  NOR2_X1 U5601 ( .A1(n8028), .A2(n8027), .ZN(n10267) );
  NOR2_X1 U5602 ( .A1(n10265), .A2(n10264), .ZN(n8031) );
  NOR2_X1 U5603 ( .A1(n8036), .A2(n8035), .ZN(n10259) );
  NOR2_X1 U5604 ( .A1(n10261), .A2(n10260), .ZN(n8035) );
  NOR2_X1 U5605 ( .A1(n8497), .A2(n8474), .ZN(n8493) );
  NAND2_X1 U5606 ( .A1(n8493), .A2(n4479), .ZN(n4563) );
  AND2_X1 U5607 ( .A1(n8500), .A2(n8481), .ZN(n4606) );
  INV_X1 U5608 ( .A(n9473), .ZN(n4674) );
  INV_X1 U5609 ( .A(n4676), .ZN(n4675) );
  AOI21_X1 U5610 ( .B1(n4677), .B2(n4678), .A(n4872), .ZN(n4676) );
  OAI21_X1 U5611 ( .B1(n9333), .B2(n9475), .A(n4589), .ZN(n4588) );
  MUX2_X1 U5612 ( .A(n9440), .B(n9290), .S(n9394), .Z(n9363) );
  INV_X1 U5613 ( .A(n4819), .ZN(n4815) );
  AOI21_X1 U5614 ( .B1(n4819), .B2(n4818), .A(n4817), .ZN(n4816) );
  INV_X1 U5615 ( .A(n8530), .ZN(n4818) );
  NAND2_X1 U5616 ( .A1(n8412), .A2(n8411), .ZN(n4811) );
  OAI21_X1 U5617 ( .B1(n8553), .B2(n5114), .A(n8552), .ZN(n8557) );
  INV_X1 U5618 ( .A(n4811), .ZN(n8484) );
  AOI21_X1 U5619 ( .B1(n8550), .B2(n8549), .A(n8548), .ZN(n8559) );
  NOR2_X1 U5620 ( .A1(n9388), .A2(n4665), .ZN(n4664) );
  NOR2_X1 U5621 ( .A1(n5842), .A2(n5019), .ZN(n5018) );
  INV_X1 U5622 ( .A(n5774), .ZN(n5019) );
  INV_X1 U5623 ( .A(SI_14_), .ZN(n4961) );
  NAND2_X1 U5624 ( .A1(n7616), .A2(n9319), .ZN(n9316) );
  NAND2_X1 U5625 ( .A1(n9450), .A2(n4687), .ZN(n4862) );
  OR2_X1 U5626 ( .A1(n9983), .A2(n9975), .ZN(n4987) );
  NOR2_X1 U5627 ( .A1(n5013), .A2(n5012), .ZN(n5011) );
  INV_X1 U5628 ( .A(n5775), .ZN(n5012) );
  INV_X1 U5629 ( .A(n5018), .ZN(n5013) );
  INV_X1 U5630 ( .A(n5842), .ZN(n5015) );
  INV_X1 U5631 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5451) );
  NOR2_X1 U5632 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5449) );
  INV_X1 U5633 ( .A(n4978), .ZN(n4974) );
  NAND2_X1 U5634 ( .A1(n4953), .A2(n4956), .ZN(n4952) );
  OAI21_X1 U5635 ( .B1(n8144), .B2(n4636), .A(n4635), .ZN(n5708) );
  NAND2_X1 U5636 ( .A1(n8144), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n4635) );
  NAND2_X1 U5637 ( .A1(n5456), .A2(n10476), .ZN(n5714) );
  NOR2_X1 U5638 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5716) );
  OAI21_X1 U5639 ( .B1(n5778), .B2(n4655), .A(n4654), .ZN(n5666) );
  NAND2_X1 U5640 ( .A1(n5778), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n4654) );
  INV_X1 U5641 ( .A(SI_9_), .ZN(n10418) );
  XNOR2_X1 U5642 ( .A(n7138), .B(n6191), .ZN(n7140) );
  INV_X1 U5643 ( .A(n7301), .ZN(n7258) );
  CLKBUF_X1 U5644 ( .A(n7301), .Z(n8090) );
  NAND2_X1 U5645 ( .A1(n8083), .A2(n8882), .ZN(n5201) );
  INV_X1 U5646 ( .A(n5204), .ZN(n5200) );
  NOR2_X1 U5647 ( .A1(n6981), .A2(n4640), .ZN(n5417) );
  NOR2_X1 U5648 ( .A1(n6242), .A2(n10242), .ZN(n5422) );
  NAND2_X1 U5649 ( .A1(n7019), .A2(n5326), .ZN(n5329) );
  AND2_X1 U5650 ( .A1(n6920), .A2(n5332), .ZN(n5334) );
  INV_X1 U5651 ( .A(n8676), .ZN(n4761) );
  NOR2_X1 U5652 ( .A1(n4753), .A2(n8690), .ZN(n4750) );
  NAND2_X1 U5653 ( .A1(n8702), .A2(n4877), .ZN(n5436) );
  NAND2_X1 U5654 ( .A1(n4571), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4877) );
  OR2_X1 U5655 ( .A1(n8582), .A2(n8182), .ZN(n6555) );
  AND2_X1 U5656 ( .A1(n6373), .A2(n4795), .ZN(n4794) );
  INV_X1 U5657 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n4795) );
  INV_X1 U5658 ( .A(n6392), .ZN(n6374) );
  INV_X1 U5659 ( .A(n5130), .ZN(n5126) );
  AND2_X1 U5660 ( .A1(n5128), .A2(n5133), .ZN(n5122) );
  NOR2_X1 U5661 ( .A1(n6280), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n4787) );
  AND2_X1 U5662 ( .A1(n4706), .A2(n6266), .ZN(n4705) );
  INV_X1 U5663 ( .A(n8486), .ZN(n5106) );
  NOR2_X1 U5664 ( .A1(n5107), .A2(n7432), .ZN(n5103) );
  INV_X1 U5665 ( .A(n8490), .ZN(n5107) );
  INV_X1 U5666 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n4783) );
  INV_X1 U5667 ( .A(n6577), .ZN(n7136) );
  INV_X1 U5668 ( .A(n6455), .ZN(n5061) );
  NAND2_X1 U5669 ( .A1(n8810), .A2(n8547), .ZN(n5110) );
  INV_X1 U5670 ( .A(n8510), .ZN(n5101) );
  INV_X1 U5671 ( .A(n8516), .ZN(n5102) );
  NOR2_X1 U5672 ( .A1(n5278), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n5270) );
  AND2_X1 U5673 ( .A1(n9219), .A2(n5083), .ZN(n5082) );
  NAND2_X1 U5674 ( .A1(n5084), .A2(n6712), .ZN(n5083) );
  INV_X1 U5675 ( .A(n9141), .ZN(n5084) );
  AND2_X1 U5676 ( .A1(n5076), .A2(n6790), .ZN(n4694) );
  AND2_X1 U5677 ( .A1(n5074), .A2(n9101), .ZN(n5073) );
  NAND2_X1 U5678 ( .A1(n5077), .A2(n5076), .ZN(n5074) );
  INV_X1 U5679 ( .A(n6597), .ZN(n6611) );
  NOR2_X1 U5680 ( .A1(n9683), .A2(n9381), .ZN(n4941) );
  NAND2_X1 U5681 ( .A1(n9393), .A2(n9683), .ZN(n4942) );
  NOR2_X1 U5682 ( .A1(n6163), .A2(n6873), .ZN(n4991) );
  AND2_X1 U5683 ( .A1(n9721), .A2(n5026), .ZN(n5025) );
  NAND2_X1 U5684 ( .A1(n5027), .A2(n6004), .ZN(n5026) );
  INV_X1 U5685 ( .A(n6003), .ZN(n5027) );
  AND2_X1 U5686 ( .A1(n9706), .A2(n10018), .ZN(n6103) );
  NAND2_X1 U5687 ( .A1(n5993), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6016) );
  INV_X1 U5688 ( .A(n5995), .ZN(n5993) );
  OR2_X1 U5689 ( .A1(n9741), .A2(n9717), .ZN(n9384) );
  OR2_X1 U5690 ( .A1(n5971), .A2(n10521), .ZN(n5995) );
  NAND2_X1 U5691 ( .A1(n5003), .A2(n5002), .ZN(n5000) );
  NOR2_X1 U5692 ( .A1(n9957), .A2(n9960), .ZN(n5003) );
  INV_X1 U5693 ( .A(n4618), .ZN(n5879) );
  NOR2_X1 U5694 ( .A1(n9870), .A2(n5807), .ZN(n8224) );
  INV_X1 U5695 ( .A(n4617), .ZN(n5787) );
  NOR2_X1 U5696 ( .A1(n6099), .A2(n4993), .ZN(n4992) );
  NAND2_X1 U5697 ( .A1(n4995), .A2(n4994), .ZN(n4993) );
  OR2_X1 U5698 ( .A1(n5743), .A2(n5742), .ZN(n5767) );
  INV_X1 U5699 ( .A(n9449), .ZN(n4856) );
  INV_X1 U5700 ( .A(n5630), .ZN(n5031) );
  INV_X1 U5701 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5640) );
  OR2_X1 U5702 ( .A1(n5641), .A2(n5640), .ZN(n5659) );
  NAND2_X1 U5703 ( .A1(n5601), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5641) );
  INV_X1 U5704 ( .A(n5603), .ZN(n5601) );
  AND2_X1 U5705 ( .A1(n4998), .A2(n10103), .ZN(n4997) );
  AND2_X1 U5706 ( .A1(n9304), .A2(n10116), .ZN(n4998) );
  NAND2_X1 U5707 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5549) );
  CLKBUF_X1 U5708 ( .A(n9451), .Z(n4573) );
  AND2_X1 U5709 ( .A1(n9497), .A2(n9379), .ZN(n9701) );
  NAND2_X1 U5710 ( .A1(n6102), .A2(n4986), .ZN(n4985) );
  INV_X1 U5711 ( .A(n4987), .ZN(n4986) );
  NAND2_X1 U5712 ( .A1(n4582), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4697) );
  OR2_X1 U5713 ( .A1(n6860), .A2(n6131), .ZN(n7730) );
  NOR2_X1 U5714 ( .A1(n5713), .A2(n5461), .ZN(n4682) );
  AND2_X1 U5715 ( .A1(n4430), .A2(n5460), .ZN(n4681) );
  NAND2_X1 U5716 ( .A1(n6059), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6061) );
  INV_X1 U5717 ( .A(n5825), .ZN(n5822) );
  NAND2_X1 U5718 ( .A1(n5796), .A2(n5795), .ZN(n5797) );
  NAND2_X1 U5719 ( .A1(n5733), .A2(n5732), .ZN(n5753) );
  NAND2_X1 U5720 ( .A1(n4800), .A2(n4799), .ZN(n4798) );
  NAND2_X1 U5721 ( .A1(n4599), .A2(n4598), .ZN(n5731) );
  INV_X1 U5722 ( .A(n5711), .ZN(n4598) );
  INV_X1 U5723 ( .A(n5759), .ZN(n4599) );
  OAI21_X1 U5724 ( .B1(n8144), .B2(n4601), .A(n4600), .ZN(n5669) );
  NAND2_X1 U5725 ( .A1(n8144), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n4600) );
  INV_X1 U5726 ( .A(n5566), .ZN(n5567) );
  OAI21_X1 U5727 ( .B1(n5584), .B2(n4620), .A(n4619), .ZN(n5486) );
  NAND2_X1 U5728 ( .A1(n5584), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4619) );
  NAND2_X1 U5729 ( .A1(n5584), .A2(n6948), .ZN(n4608) );
  INV_X2 U5730 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n10405) );
  AND2_X1 U5731 ( .A1(n4578), .A2(n4577), .ZN(n8265) );
  NAND2_X1 U5732 ( .A1(n8264), .A2(n8263), .ZN(n4577) );
  NAND2_X1 U5733 ( .A1(n5195), .A2(n5194), .ZN(n5193) );
  INV_X1 U5734 ( .A(n8369), .ZN(n5194) );
  NOR2_X1 U5735 ( .A1(n5193), .A2(n5199), .ZN(n5188) );
  NAND2_X1 U5736 ( .A1(n8087), .A2(n8867), .ZN(n5168) );
  INV_X1 U5737 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U5738 ( .A1(n5203), .A2(n8313), .ZN(n5202) );
  OAI21_X1 U5739 ( .B1(n5154), .B2(n5153), .A(n5155), .ZN(n8301) );
  AOI21_X1 U5740 ( .B1(n5157), .B2(n4476), .A(n5156), .ZN(n5155) );
  NAND2_X1 U5741 ( .A1(n5157), .A2(n4452), .ZN(n5153) );
  NAND2_X1 U5742 ( .A1(n5182), .A2(n4464), .ZN(n5181) );
  NAND2_X1 U5743 ( .A1(n4459), .A2(n5178), .ZN(n5177) );
  OR2_X1 U5744 ( .A1(n8322), .A2(n5196), .ZN(n5195) );
  INV_X1 U5745 ( .A(n5201), .ZN(n5196) );
  NAND2_X1 U5746 ( .A1(n8579), .A2(n4823), .ZN(n4822) );
  OR2_X1 U5747 ( .A1(n6225), .A2(n10558), .ZN(n6196) );
  NAND2_X1 U5748 ( .A1(n7152), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7218) );
  NAND2_X1 U5749 ( .A1(n5315), .A2(n7209), .ZN(n7214) );
  AOI21_X1 U5750 ( .B1(n5420), .B2(n5320), .A(n5421), .ZN(n7180) );
  NAND2_X1 U5751 ( .A1(n5322), .A2(n6930), .ZN(n7017) );
  AOI21_X1 U5752 ( .B1(n7179), .B2(n7013), .A(n7014), .ZN(n7012) );
  NAND2_X1 U5753 ( .A1(n4901), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4899) );
  NAND2_X1 U5754 ( .A1(n4569), .A2(n6253), .ZN(n5221) );
  INV_X1 U5755 ( .A(n5329), .ZN(n4569) );
  NAND2_X1 U5756 ( .A1(n5329), .A2(n7385), .ZN(n6918) );
  NAND2_X1 U5757 ( .A1(n4529), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7383) );
  OR2_X1 U5758 ( .A1(n5334), .A2(n7540), .ZN(n8638) );
  NAND2_X1 U5759 ( .A1(n4897), .A2(n7881), .ZN(n4896) );
  NAND2_X1 U5760 ( .A1(n4523), .A2(n4438), .ZN(n7882) );
  OAI21_X1 U5761 ( .B1(n4438), .B2(n6896), .A(n4928), .ZN(n6895) );
  NAND2_X1 U5762 ( .A1(n5338), .A2(n4488), .ZN(n4928) );
  OR2_X1 U5763 ( .A1(n5298), .A2(n5293), .ZN(n5339) );
  NAND2_X1 U5764 ( .A1(n4758), .A2(n5394), .ZN(n8678) );
  OR2_X1 U5765 ( .A1(n6899), .A2(n5395), .ZN(n4758) );
  OR2_X1 U5766 ( .A1(n8671), .A2(n8982), .ZN(n4586) );
  AND4_X1 U5767 ( .A1(n4909), .A2(n4905), .A3(n4906), .A4(n4908), .ZN(n8697)
         );
  NAND2_X1 U5768 ( .A1(n4912), .A2(n4907), .ZN(n4906) );
  AND2_X1 U5769 ( .A1(n8673), .A2(n8695), .ZN(n4907) );
  NAND2_X1 U5770 ( .A1(n8697), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8696) );
  NAND2_X1 U5771 ( .A1(n5440), .A2(n5441), .ZN(n4892) );
  INV_X1 U5772 ( .A(n4889), .ZN(n4888) );
  OAI21_X1 U5773 ( .B1(n8741), .B2(n4892), .A(n4890), .ZN(n4889) );
  NAND2_X1 U5774 ( .A1(n4891), .A2(n5442), .ZN(n4890) );
  INV_X1 U5775 ( .A(n5440), .ZN(n4891) );
  AND2_X1 U5776 ( .A1(n5351), .A2(n4448), .ZN(n4933) );
  AND2_X1 U5777 ( .A1(n6533), .A2(n6534), .ZN(n6538) );
  INV_X1 U5778 ( .A(n6554), .ZN(n8778) );
  NAND2_X1 U5779 ( .A1(n6471), .A2(n6470), .ZN(n6484) );
  INV_X1 U5780 ( .A(n6472), .ZN(n6471) );
  NAND2_X1 U5781 ( .A1(n6447), .A2(n6446), .ZN(n6458) );
  INV_X1 U5782 ( .A(n6448), .ZN(n6447) );
  NAND2_X1 U5783 ( .A1(n6437), .A2(n6448), .ZN(n8334) );
  INV_X1 U5784 ( .A(n4782), .ZN(n6436) );
  OR2_X1 U5785 ( .A1(n6412), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6424) );
  NAND2_X1 U5786 ( .A1(n6374), .A2(n4794), .ZN(n6405) );
  AOI21_X1 U5787 ( .B1(n8884), .B2(n6494), .A(n6387), .ZN(n8870) );
  NAND2_X1 U5788 ( .A1(n6374), .A2(n6373), .ZN(n6394) );
  INV_X1 U5789 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n4791) );
  NAND2_X1 U5790 ( .A1(n6343), .A2(n4792), .ZN(n6360) );
  NAND2_X1 U5791 ( .A1(n6343), .A2(n10383), .ZN(n6352) );
  NAND2_X1 U5792 ( .A1(n6313), .A2(n4474), .ZN(n6344) );
  INV_X1 U5793 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n4789) );
  NAND2_X1 U5794 ( .A1(n6313), .A2(n10445), .ZN(n6323) );
  NAND2_X1 U5795 ( .A1(n6313), .A2(n4790), .ZN(n6334) );
  INV_X1 U5796 ( .A(n8614), .ZN(n8288) );
  NAND2_X1 U5797 ( .A1(n4785), .A2(n4784), .ZN(n6314) );
  INV_X1 U5798 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n4784) );
  INV_X1 U5799 ( .A(n6301), .ZN(n4785) );
  OR2_X1 U5800 ( .A1(n8483), .A2(n5131), .ZN(n8423) );
  INV_X1 U5801 ( .A(n4787), .ZN(n6290) );
  NAND2_X1 U5802 ( .A1(n4787), .A2(n4786), .ZN(n6301) );
  INV_X1 U5803 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n4786) );
  AOI21_X1 U5804 ( .B1(n5139), .B2(n8474), .A(n5137), .ZN(n5136) );
  INV_X1 U5805 ( .A(n8477), .ZN(n5137) );
  OR2_X1 U5806 ( .A1(n6278), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U5807 ( .A1(n6257), .A2(n6256), .ZN(n6278) );
  INV_X1 U5808 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6256) );
  INV_X1 U5809 ( .A(n6258), .ZN(n6257) );
  NAND2_X1 U5810 ( .A1(n7464), .A2(n8416), .ZN(n7598) );
  OR2_X1 U5811 ( .A1(n6245), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6258) );
  NAND2_X1 U5812 ( .A1(n10293), .A2(n4783), .ZN(n6233) );
  NAND2_X1 U5813 ( .A1(n6509), .A2(n8467), .ZN(n7427) );
  INV_X1 U5814 ( .A(n7432), .ZN(n8465) );
  NAND2_X1 U5815 ( .A1(n7427), .A2(n8465), .ZN(n7426) );
  AND2_X1 U5816 ( .A1(n8585), .A2(n8596), .ZN(n7171) );
  NAND2_X1 U5817 ( .A1(n7162), .A2(n7163), .ZN(n7164) );
  OR2_X1 U5818 ( .A1(n8570), .A2(n7136), .ZN(n6879) );
  OR2_X1 U5819 ( .A1(n8877), .A2(n8833), .ZN(n8864) );
  AND2_X1 U5820 ( .A1(n6878), .A2(n6578), .ZN(n7075) );
  AND2_X1 U5821 ( .A1(n10189), .A2(n7171), .ZN(n7078) );
  NOR2_X1 U5822 ( .A1(n8772), .A2(n8771), .ZN(n8991) );
  INV_X1 U5823 ( .A(n6528), .ZN(n5059) );
  AND2_X1 U5824 ( .A1(n8569), .A2(n6528), .ZN(n8567) );
  INV_X1 U5825 ( .A(n4721), .ZN(n4720) );
  OAI21_X1 U5826 ( .B1(n4727), .B2(n4725), .A(n8542), .ZN(n4721) );
  NAND2_X1 U5827 ( .A1(n4724), .A2(n4727), .ZN(n8836) );
  NAND2_X1 U5828 ( .A1(n8878), .A2(n6401), .ZN(n4724) );
  CLKBUF_X1 U5829 ( .A(n8845), .Z(n8861) );
  NAND2_X1 U5830 ( .A1(n5120), .A2(n8523), .ZN(n8890) );
  AND2_X1 U5831 ( .A1(n4714), .A2(n5048), .ZN(n4713) );
  AOI21_X1 U5832 ( .B1(n5050), .B2(n5053), .A(n4491), .ZN(n5048) );
  OR2_X1 U5833 ( .A1(n9055), .A2(n8313), .ZN(n8519) );
  AND2_X1 U5834 ( .A1(n8511), .A2(n8510), .ZN(n8923) );
  INV_X1 U5835 ( .A(n6539), .ZN(n5404) );
  AND2_X1 U5836 ( .A1(n5267), .A2(n5281), .ZN(n6563) );
  INV_X1 U5837 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5356) );
  INV_X1 U5838 ( .A(n5260), .ZN(n5185) );
  INV_X1 U5839 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5288) );
  INV_X1 U5840 ( .A(n5184), .ZN(n5317) );
  NAND2_X1 U5841 ( .A1(n6061), .A2(n6060), .ZN(n6105) );
  OR2_X1 U5842 ( .A1(n6795), .A2(n5078), .ZN(n5076) );
  AND2_X1 U5843 ( .A1(n6795), .A2(n5078), .ZN(n5077) );
  NAND2_X1 U5844 ( .A1(n5905), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5948) );
  CLKBUF_X2 U5845 ( .A(n6837), .Z(n6665) );
  NAND2_X1 U5846 ( .A1(n9157), .A2(n4469), .ZN(n6749) );
  INV_X1 U5847 ( .A(n4451), .ZN(n5095) );
  AOI21_X1 U5848 ( .B1(n9613), .B2(n7048), .A(n7047), .ZN(n7065) );
  NOR2_X1 U5849 ( .A1(n10066), .A2(n4551), .ZN(n10063) );
  OR2_X1 U5850 ( .A1(n10064), .A2(n10065), .ZN(n4551) );
  NOR2_X1 U5851 ( .A1(n10071), .A2(n10072), .ZN(n10070) );
  NOR2_X1 U5852 ( .A1(n10086), .A2(n10087), .ZN(n10085) );
  OR2_X1 U5853 ( .A1(n8202), .A2(n4531), .ZN(n4842) );
  OAI21_X1 U5854 ( .B1(n8194), .B2(n8193), .A(n8192), .ZN(n8195) );
  NAND2_X1 U5855 ( .A1(n9624), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9623) );
  NOR3_X1 U5856 ( .A1(n9661), .A2(n9660), .A3(n9659), .ZN(n9658) );
  NAND2_X1 U5857 ( .A1(n4989), .A2(n6103), .ZN(n9681) );
  NOR2_X1 U5858 ( .A1(n9683), .A2(n4990), .ZN(n4989) );
  INV_X1 U5859 ( .A(n4991), .ZN(n4990) );
  AND2_X1 U5860 ( .A1(n9809), .A2(n4999), .ZN(n9740) );
  NOR2_X1 U5861 ( .A1(n5000), .A2(n9741), .ZN(n4999) );
  AND2_X1 U5862 ( .A1(n9384), .A2(n9492), .ZN(n9733) );
  NAND2_X1 U5863 ( .A1(n9809), .A2(n5001), .ZN(n9756) );
  INV_X1 U5864 ( .A(n5000), .ZN(n5001) );
  NAND2_X1 U5865 ( .A1(n9809), .A2(n5003), .ZN(n9772) );
  NAND2_X1 U5866 ( .A1(n9809), .A2(n9789), .ZN(n9784) );
  OR2_X1 U5867 ( .A1(n9971), .A2(n9124), .ZN(n9802) );
  OR2_X1 U5868 ( .A1(n9975), .A2(n9820), .ZN(n4597) );
  AND2_X1 U5869 ( .A1(n9335), .A2(n9487), .ZN(n9834) );
  INV_X1 U5870 ( .A(n9860), .ZN(n4548) );
  INV_X1 U5871 ( .A(n5810), .ZN(n5808) );
  NAND3_X1 U5872 ( .A1(n7706), .A2(n4992), .A3(n9288), .ZN(n9870) );
  NAND2_X1 U5873 ( .A1(n5021), .A2(n5774), .ZN(n9879) );
  AND2_X1 U5874 ( .A1(n4992), .A2(n7706), .ZN(n9890) );
  NAND2_X1 U5875 ( .A1(n7706), .A2(n4996), .ZN(n9905) );
  NOR2_X1 U5876 ( .A1(n6099), .A2(n9326), .ZN(n4996) );
  NAND2_X1 U5877 ( .A1(n4616), .A2(n4486), .ZN(n5723) );
  INV_X1 U5878 ( .A(n5696), .ZN(n4616) );
  NAND2_X1 U5879 ( .A1(n4615), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5743) );
  INV_X1 U5880 ( .A(n5723), .ZN(n4615) );
  INV_X1 U5881 ( .A(n5005), .ZN(n5004) );
  OAI21_X1 U5882 ( .B1(n5008), .B2(n5685), .A(n4503), .ZN(n5005) );
  OR2_X1 U5883 ( .A1(n6932), .A2(n5676), .ZN(n5628) );
  AND2_X1 U5884 ( .A1(n4997), .A2(n6098), .ZN(n7758) );
  NAND2_X1 U5885 ( .A1(n6098), .A2(n4998), .ZN(n7774) );
  NAND2_X1 U5886 ( .A1(n6098), .A2(n10116), .ZN(n7776) );
  NOR2_X1 U5887 ( .A1(n7448), .A2(n4687), .ZN(n4686) );
  CLKBUF_X1 U5888 ( .A(n7442), .Z(n7443) );
  NOR2_X1 U5889 ( .A1(n7815), .A2(n6097), .ZN(n7951) );
  NOR2_X1 U5890 ( .A1(n9689), .A2(n10143), .ZN(n6150) );
  NAND2_X1 U5891 ( .A1(n5656), .A2(n5655), .ZN(n9204) );
  NAND2_X1 U5892 ( .A1(n7611), .A2(n7615), .ZN(n7610) );
  NAND2_X1 U5893 ( .A1(n7748), .A2(n5630), .ZN(n7611) );
  OR2_X1 U5894 ( .A1(n8136), .A2(n8135), .ZN(n8137) );
  XNOR2_X1 U5895 ( .A(n8150), .B(n8149), .ZN(n8398) );
  INV_X1 U5896 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5474) );
  XNOR2_X1 U5897 ( .A(n6110), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U5898 ( .A1(n6056), .A2(n4430), .ZN(n6111) );
  XNOR2_X1 U5899 ( .A(n5968), .B(n5967), .ZN(n7998) );
  NAND2_X1 U5900 ( .A1(n5962), .A2(n5983), .ZN(n5968) );
  OR2_X1 U5901 ( .A1(n6061), .A2(n6060), .ZN(n6062) );
  INV_X1 U5902 ( .A(n5885), .ZN(n4981) );
  OAI21_X1 U5903 ( .B1(n5863), .B2(n4984), .A(n5862), .ZN(n5887) );
  AND2_X1 U5904 ( .A1(n5849), .A2(n5848), .ZN(n8209) );
  INV_X1 U5905 ( .A(n5480), .ZN(n5482) );
  NOR2_X1 U5906 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5531) );
  NAND2_X1 U5907 ( .A1(n7548), .A2(n7547), .ZN(n7553) );
  NAND2_X1 U5908 ( .A1(n8384), .A2(n8099), .ZN(n8252) );
  NAND2_X1 U5909 ( .A1(n8384), .A2(n5173), .ZN(n8253) );
  AOI21_X1 U5910 ( .B1(n5173), .B2(n5172), .A(n4493), .ZN(n5171) );
  OAI21_X1 U5911 ( .B1(n8341), .B2(n8340), .A(n5168), .ZN(n8281) );
  NAND2_X1 U5912 ( .A1(n8079), .A2(n5204), .ZN(n8316) );
  NAND2_X1 U5913 ( .A1(n5197), .A2(n5202), .ZN(n8323) );
  INV_X1 U5914 ( .A(n7308), .ZN(n5152) );
  NAND2_X1 U5915 ( .A1(n7854), .A2(n7853), .ZN(n7855) );
  OR2_X1 U5916 ( .A1(n7106), .A2(n7127), .ZN(n8373) );
  INV_X1 U5917 ( .A(n5162), .ZN(n8347) );
  AND2_X1 U5918 ( .A1(n6202), .A2(n6201), .ZN(n4607) );
  INV_X1 U5919 ( .A(n5189), .ZN(n8370) );
  AOI21_X1 U5920 ( .B1(n5197), .B2(n4455), .A(n5190), .ZN(n5189) );
  INV_X1 U5921 ( .A(n5195), .ZN(n5190) );
  AND2_X1 U5922 ( .A1(n7418), .A2(n7417), .ZN(n7420) );
  INV_X1 U5923 ( .A(n8618), .ZN(n7421) );
  NOR2_X1 U5924 ( .A1(n8059), .A2(n8058), .ZN(n8061) );
  AND2_X1 U5925 ( .A1(n8057), .A2(n8056), .ZN(n8058) );
  INV_X1 U5926 ( .A(n8378), .ZN(n8385) );
  NAND2_X1 U5927 ( .A1(n7103), .A2(n7102), .ZN(n8388) );
  NOR2_X1 U5928 ( .A1(n8441), .A2(n8585), .ZN(n8444) );
  NAND2_X1 U5929 ( .A1(n4564), .A2(n8434), .ZN(n8586) );
  NAND2_X1 U5930 ( .A1(n8594), .A2(n8593), .ZN(n4564) );
  XNOR2_X1 U5931 ( .A(n5279), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U5932 ( .A1(n8590), .A2(n4762), .ZN(n8591) );
  NOR2_X1 U5933 ( .A1(n5409), .A2(n6539), .ZN(n4762) );
  INV_X1 U5934 ( .A(n8772), .ZN(n8593) );
  NAND2_X1 U5935 ( .A1(n6490), .A2(n6489), .ZN(n8607) );
  INV_X1 U5936 ( .A(n8543), .ZN(n8839) );
  INV_X1 U5937 ( .A(n8880), .ZN(n8611) );
  INV_X1 U5938 ( .A(n7801), .ZN(n8925) );
  CLKBUF_X1 U5939 ( .A(n6505), .Z(n8621) );
  NAND2_X1 U5940 ( .A1(n4902), .A2(n4903), .ZN(n7001) );
  AND2_X1 U5941 ( .A1(n7210), .A2(n4920), .ZN(n7154) );
  OR2_X1 U5942 ( .A1(P2_U3150), .A2(n5363), .ZN(n8759) );
  OAI21_X1 U5943 ( .B1(n7178), .B2(n4771), .A(n4769), .ZN(n7391) );
  NAND2_X1 U5944 ( .A1(n4772), .A2(n6916), .ZN(n4768) );
  INV_X1 U5945 ( .A(n4765), .ZN(n4764) );
  OAI21_X1 U5946 ( .B1(n4769), .B2(n4767), .A(n4766), .ZN(n4765) );
  NOR2_X1 U5947 ( .A1(n4876), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4875) );
  AND2_X1 U5948 ( .A1(n4874), .A2(n5426), .ZN(n4876) );
  XNOR2_X1 U5949 ( .A(n5303), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8637) );
  AOI21_X1 U5950 ( .B1(n8640), .B2(n8638), .A(n8639), .ZN(n8642) );
  AND3_X1 U5951 ( .A1(n4896), .A2(n5429), .A3(P2_REG1_REG_11__SCAN_IN), .ZN(
        n7872) );
  NAND2_X1 U5952 ( .A1(n4896), .A2(n5429), .ZN(n7873) );
  AND2_X1 U5953 ( .A1(n4894), .A2(n4893), .ZN(n6894) );
  NAND2_X1 U5954 ( .A1(n4557), .A2(n8656), .ZN(n4556) );
  INV_X1 U5955 ( .A(n5431), .ZN(n4557) );
  CLKBUF_X1 U5956 ( .A(n8665), .Z(n4575) );
  NAND2_X1 U5957 ( .A1(n8674), .A2(n8672), .ZN(n4911) );
  AND2_X1 U5958 ( .A1(n4755), .A2(n4751), .ZN(n8691) );
  NOR2_X1 U5959 ( .A1(n8725), .A2(n10471), .ZN(n8749) );
  AND2_X1 U5960 ( .A1(n5443), .A2(n6539), .ZN(n8750) );
  INV_X1 U5961 ( .A(n5056), .ZN(n5055) );
  INV_X1 U5962 ( .A(n5123), .ZN(n7798) );
  AOI21_X1 U5963 ( .B1(n5132), .B2(n5130), .A(n5127), .ZN(n5123) );
  INV_X1 U5964 ( .A(n5128), .ZN(n5127) );
  NAND2_X1 U5965 ( .A1(n5064), .A2(n6309), .ZN(n7799) );
  NAND2_X1 U5966 ( .A1(n7456), .A2(n6251), .ZN(n4708) );
  NAND2_X1 U5967 ( .A1(n7108), .A2(n7078), .ZN(n8885) );
  INV_X1 U5968 ( .A(n8873), .ZN(n10178) );
  INV_X1 U5969 ( .A(n8885), .ZN(n10175) );
  NAND2_X1 U5970 ( .A1(n5062), .A2(n6455), .ZN(n8791) );
  NAND2_X1 U5971 ( .A1(n6469), .A2(n6468), .ZN(n8571) );
  NAND2_X1 U5972 ( .A1(n6457), .A2(n6456), .ZN(n9001) );
  NAND2_X1 U5973 ( .A1(n5118), .A2(n8560), .ZN(n8789) );
  NAND2_X1 U5974 ( .A1(n6445), .A2(n6444), .ZN(n9007) );
  NAND2_X1 U5975 ( .A1(n4731), .A2(n6443), .ZN(n8800) );
  NAND2_X1 U5976 ( .A1(n5069), .A2(n6432), .ZN(n8813) );
  OAI21_X1 U5977 ( .B1(n4632), .B2(n5114), .A(n5112), .ZN(n8809) );
  NAND2_X1 U5978 ( .A1(n5111), .A2(n8551), .ZN(n8172) );
  NAND2_X1 U5979 ( .A1(n4632), .A2(n5115), .ZN(n5111) );
  NAND2_X1 U5980 ( .A1(n6411), .A2(n6410), .ZN(n9023) );
  NAND2_X1 U5981 ( .A1(n4632), .A2(n8541), .ZN(n8820) );
  NAND2_X1 U5982 ( .A1(n6404), .A2(n6403), .ZN(n9028) );
  NAND2_X1 U5983 ( .A1(n6359), .A2(n6358), .ZN(n9049) );
  NAND2_X1 U5984 ( .A1(n5049), .A2(n6349), .ZN(n8906) );
  NAND2_X1 U5985 ( .A1(n8914), .A2(n8513), .ZN(n5049) );
  NAND2_X1 U5986 ( .A1(n6342), .A2(n6341), .ZN(n9061) );
  NAND2_X1 U5987 ( .A1(n8922), .A2(n8510), .ZN(n5099) );
  NAND2_X1 U5988 ( .A1(n6331), .A2(n6330), .ZN(n9067) );
  NAND2_X1 U5989 ( .A1(n4743), .A2(n6320), .ZN(n7907) );
  INV_X1 U5990 ( .A(n7892), .ZN(n8167) );
  INV_X1 U5991 ( .A(n9045), .ZN(n9066) );
  NAND2_X1 U5992 ( .A1(n7108), .A2(n6951), .ZN(n6961) );
  INV_X1 U5993 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9076) );
  AND2_X1 U5994 ( .A1(n5143), .A2(n6172), .ZN(n5142) );
  INV_X1 U5995 ( .A(n5281), .ZN(n5283) );
  INV_X1 U5996 ( .A(n6563), .ZN(n8068) );
  NAND2_X1 U5997 ( .A1(n5254), .A2(n5352), .ZN(n5251) );
  INV_X1 U5998 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8054) );
  INV_X1 U5999 ( .A(n8592), .ZN(n7841) );
  INV_X1 U6000 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7675) );
  NAND2_X1 U6001 ( .A1(n5276), .A2(n5352), .ZN(n5277) );
  INV_X1 U6002 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7501) );
  INV_X1 U6003 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10411) );
  INV_X1 U6004 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7342) );
  INV_X1 U6005 ( .A(n7159), .ZN(n6928) );
  NAND2_X1 U6006 ( .A1(n7573), .A2(n4702), .ZN(n7643) );
  INV_X1 U6007 ( .A(n6661), .ZN(n4703) );
  NAND2_X1 U6008 ( .A1(n7573), .A2(n6661), .ZN(n7639) );
  NAND2_X1 U6009 ( .A1(n4691), .A2(n4487), .ZN(n4692) );
  NAND2_X1 U6010 ( .A1(n5086), .A2(n4444), .ZN(n4691) );
  NAND2_X1 U6011 ( .A1(n6031), .A2(n6030), .ZN(n8118) );
  NAND2_X1 U6012 ( .A1(n5072), .A2(n5076), .ZN(n9100) );
  OR2_X1 U6013 ( .A1(n4440), .A2(n5077), .ZN(n5072) );
  AND2_X1 U6014 ( .A1(n6855), .A2(n9276), .ZN(n6856) );
  CLKBUF_X1 U6015 ( .A(n9139), .Z(n9140) );
  AND2_X1 U6016 ( .A1(n6022), .A2(n6021), .ZN(n9736) );
  OR2_X1 U6017 ( .A1(n9725), .A2(n6094), .ZN(n6022) );
  NAND2_X1 U6018 ( .A1(n6651), .A2(n6650), .ZN(n7505) );
  INV_X1 U6019 ( .A(n6649), .ZN(n6650) );
  NAND2_X1 U6020 ( .A1(n6749), .A2(n6748), .ZN(n9173) );
  CLKBUF_X1 U6021 ( .A(n9186), .Z(n9187) );
  AND2_X1 U6022 ( .A1(n9174), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9267) );
  NAND2_X1 U6023 ( .A1(n5093), .A2(n5094), .ZN(n9211) );
  NOR2_X1 U6024 ( .A1(n5095), .A2(n4462), .ZN(n5094) );
  NAND2_X1 U6025 ( .A1(n5081), .A2(n6712), .ZN(n9218) );
  NAND2_X1 U6026 ( .A1(n9140), .A2(n9141), .ZN(n5081) );
  NAND2_X1 U6027 ( .A1(n4440), .A2(n6795), .ZN(n9227) );
  OR2_X1 U6028 ( .A1(n4440), .A2(n6795), .ZN(n9226) );
  NAND2_X1 U6029 ( .A1(n6866), .A2(n6865), .ZN(n9250) );
  NAND2_X1 U6030 ( .A1(n5086), .A2(n6823), .ZN(n9264) );
  INV_X1 U6031 ( .A(n9262), .ZN(n9276) );
  OR2_X1 U6032 ( .A1(n9447), .A2(n9920), .ZN(n4937) );
  INV_X1 U6033 ( .A(n9402), .ZN(n4939) );
  NAND2_X1 U6034 ( .A1(n9513), .A2(n4542), .ZN(n9526) );
  INV_X1 U6035 ( .A(n6595), .ZN(n9534) );
  INV_X1 U6036 ( .A(n9771), .ZN(n9549) );
  NAND2_X1 U6037 ( .A1(n5909), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4851) );
  NAND2_X1 U6038 ( .A1(n5909), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U6039 ( .A1(n9588), .A2(n9587), .ZN(n9586) );
  INV_X1 U6040 ( .A(n4839), .ZN(n7036) );
  NOR2_X1 U6041 ( .A1(n7190), .A2(n4463), .ZN(n7270) );
  NAND2_X1 U6042 ( .A1(n7322), .A2(n7321), .ZN(n10081) );
  XNOR2_X1 U6043 ( .A(n5691), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7517) );
  OR2_X1 U6044 ( .A1(n7054), .A2(n7053), .ZN(n10098) );
  NOR2_X1 U6045 ( .A1(n7518), .A2(n7519), .ZN(n7652) );
  NOR3_X1 U6046 ( .A1(n10085), .A2(n7525), .A3(n7527), .ZN(n7650) );
  XNOR2_X1 U6047 ( .A(n4842), .B(n8205), .ZN(n9622) );
  NAND2_X1 U6048 ( .A1(n9635), .A2(n4845), .ZN(n9652) );
  NOR2_X1 U6049 ( .A1(n9631), .A2(n8200), .ZN(n9646) );
  AND2_X1 U6050 ( .A1(n6046), .A2(n9693), .ZN(n8242) );
  INV_X1 U6051 ( .A(n9719), .ZN(n4624) );
  NAND2_X1 U6052 ( .A1(n4626), .A2(n9918), .ZN(n4625) );
  NAND2_X1 U6053 ( .A1(n5024), .A2(n6004), .ZN(n9720) );
  NAND2_X1 U6054 ( .A1(n5034), .A2(n5032), .ZN(n9755) );
  INV_X1 U6055 ( .A(n5035), .ZN(n5032) );
  CLKBUF_X1 U6056 ( .A(n9752), .Z(n9753) );
  OAI21_X1 U6057 ( .B1(n9783), .B2(n5936), .A(n5935), .ZN(n9763) );
  AND2_X1 U6058 ( .A1(n5016), .A2(n5020), .ZN(n8219) );
  NAND2_X1 U6059 ( .A1(n5017), .A2(n5021), .ZN(n5016) );
  NAND2_X1 U6060 ( .A1(n9911), .A2(n9466), .ZN(n9894) );
  INV_X1 U6061 ( .A(n9922), .ZN(n10110) );
  NAND2_X1 U6062 ( .A1(n7704), .A2(n5685), .ZN(n7719) );
  NAND2_X1 U6063 ( .A1(n9460), .A2(n9457), .ZN(n7712) );
  OR2_X1 U6064 ( .A1(n6857), .A2(n10269), .ZN(n9922) );
  OR2_X1 U6065 ( .A1(n10112), .A2(n7740), .ZN(n10115) );
  NAND2_X1 U6066 ( .A1(n6072), .A2(n4688), .ZN(n7945) );
  OR2_X1 U6067 ( .A1(n10112), .A2(n7770), .ZN(n9926) );
  OR2_X1 U6068 ( .A1(n8151), .A2(n4970), .ZN(n4850) );
  INV_X1 U6069 ( .A(n4849), .ZN(n4848) );
  INV_X1 U6070 ( .A(n10115), .ZN(n9929) );
  NAND2_X1 U6071 ( .A1(n4868), .A2(n4656), .ZN(n5041) );
  AND2_X1 U6072 ( .A1(n4867), .A2(n6162), .ZN(n4656) );
  INV_X1 U6073 ( .A(n4631), .ZN(n4630) );
  CLKBUF_X1 U6074 ( .A(n9204), .Z(n4572) );
  AND2_X2 U6075 ( .A1(n5639), .A2(n5638), .ZN(n7783) );
  OR2_X1 U6076 ( .A1(n5676), .A2(n6943), .ZN(n5506) );
  INV_X1 U6077 ( .A(n4653), .ZN(n4652) );
  CLKBUF_X1 U6078 ( .A(n6157), .Z(n6158) );
  INV_X1 U6079 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10550) );
  XNOR2_X1 U6080 ( .A(n5943), .B(n5942), .ZN(n7934) );
  INV_X1 U6081 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10416) );
  INV_X1 U6082 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7503) );
  OAI21_X1 U6083 ( .B1(n5802), .B2(n5090), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5846) );
  NAND2_X1 U6084 ( .A1(n4944), .A2(n4650), .ZN(n5675) );
  AND2_X1 U6085 ( .A1(n4945), .A2(n5674), .ZN(n4650) );
  NAND2_X1 U6086 ( .A1(n4949), .A2(n4947), .ZN(n4944) );
  INV_X1 U6087 ( .A(n5557), .ZN(n5489) );
  NOR2_X1 U6088 ( .A1(n8025), .A2(n8024), .ZN(n10586) );
  NOR2_X1 U6089 ( .A1(n10590), .A2(n10589), .ZN(n8024) );
  NOR2_X1 U6090 ( .A1(n8030), .A2(n8029), .ZN(n10265) );
  NOR2_X1 U6091 ( .A1(n10267), .A2(n10266), .ZN(n8029) );
  NOR2_X1 U6092 ( .A1(n8034), .A2(n8033), .ZN(n10261) );
  NOR2_X1 U6093 ( .A1(n8038), .A2(n8037), .ZN(n10257) );
  NOR2_X1 U6094 ( .A1(n10259), .A2(n10258), .ZN(n8037) );
  NAND2_X1 U6095 ( .A1(n7261), .A2(n7260), .ZN(n7264) );
  INV_X1 U6096 ( .A(n5146), .ZN(n7237) );
  NAND2_X1 U6097 ( .A1(n4776), .A2(n4777), .ZN(n7011) );
  OR2_X1 U6098 ( .A1(n4780), .A2(n8760), .ZN(n4596) );
  AND2_X1 U6099 ( .A1(n5446), .A2(n4779), .ZN(n4778) );
  OAI21_X1 U6100 ( .B1(n4788), .B2(n5066), .A(n6587), .ZN(n6589) );
  NAND2_X1 U6101 ( .A1(n4642), .A2(n4641), .ZN(n8940) );
  NAND2_X1 U6102 ( .A1(n6586), .A2(n10477), .ZN(n4641) );
  NAND2_X1 U6103 ( .A1(n4739), .A2(n4447), .ZN(n8997) );
  INV_X1 U6104 ( .A(n4837), .ZN(n7283) );
  INV_X1 U6105 ( .A(n4831), .ZN(n4830) );
  INV_X1 U6106 ( .A(n9697), .ZN(n4584) );
  MUX2_X1 U6107 ( .A(n8217), .B(n8216), .S(n10161), .Z(n8218) );
  AND2_X1 U6108 ( .A1(n5234), .A2(n6136), .ZN(n5042) );
  NAND2_X1 U6109 ( .A1(n6169), .A2(n10161), .ZN(n5043) );
  INV_X1 U6110 ( .A(n4628), .ZN(n4627) );
  OAI22_X1 U6111 ( .A1(n10022), .A2(n9948), .B1(n10161), .B2(n9942), .ZN(n4628) );
  MUX2_X1 U6112 ( .A(n8160), .B(n8216), .S(n10155), .Z(n8161) );
  INV_X1 U6113 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10046) );
  OR2_X1 U6114 ( .A1(n5337), .A2(n7881), .ZN(n4438) );
  INV_X1 U6115 ( .A(n7540), .ZN(n4923) );
  INV_X1 U6116 ( .A(n5584), .ZN(n4582) );
  AND2_X1 U6117 ( .A1(n7854), .A2(n5179), .ZN(n4439) );
  INV_X1 U6118 ( .A(n8314), .ZN(n5203) );
  AND2_X1 U6119 ( .A1(n9130), .A2(n6790), .ZN(n4440) );
  NOR2_X1 U6120 ( .A1(n9878), .A2(n5817), .ZN(n4441) );
  AND2_X1 U6121 ( .A1(n6828), .A2(n6823), .ZN(n4442) );
  AND2_X1 U6122 ( .A1(n5067), .A2(n10245), .ZN(n4443) );
  INV_X1 U6123 ( .A(n8500), .ZN(n5131) );
  INV_X1 U6124 ( .A(n8513), .ZN(n5052) );
  AND2_X1 U6125 ( .A1(n8113), .A2(n4442), .ZN(n4444) );
  AND2_X1 U6126 ( .A1(n4983), .A2(n5862), .ZN(n4982) );
  INV_X1 U6127 ( .A(n4982), .ZN(n4976) );
  AND2_X1 U6128 ( .A1(n4510), .A2(n4862), .ZN(n4445) );
  INV_X1 U6129 ( .A(n5685), .ZN(n5009) );
  AND2_X1 U6130 ( .A1(n5169), .A2(n7547), .ZN(n4446) );
  INV_X1 U6131 ( .A(n10112), .ZN(n9776) );
  INV_X1 U6132 ( .A(n8695), .ZN(n4915) );
  INV_X1 U6133 ( .A(n9326), .ZN(n4994) );
  OR2_X1 U6134 ( .A1(n10230), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n4447) );
  INV_X2 U6135 ( .A(n10161), .ZN(n10159) );
  AND2_X1 U6136 ( .A1(n8747), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4448) );
  INV_X1 U6137 ( .A(n7302), .ZN(n7255) );
  INV_X1 U6138 ( .A(n6204), .ZN(n6208) );
  AND2_X1 U6139 ( .A1(n6442), .A2(n6441), .ZN(n4449) );
  NAND2_X2 U6140 ( .A1(n5741), .A2(n5740), .ZN(n10008) );
  NAND2_X1 U6141 ( .A1(n5542), .A2(n4699), .ZN(n6097) );
  OR2_X1 U6142 ( .A1(n7612), .A2(n7986), .ZN(n4450) );
  OR2_X1 U6143 ( .A1(n6770), .A2(n6769), .ZN(n4451) );
  AND2_X1 U6144 ( .A1(n7643), .A2(n7638), .ZN(n7978) );
  NOR2_X2 U6145 ( .A1(n9679), .A2(n9543), .ZN(n9514) );
  XNOR2_X1 U6146 ( .A(n6138), .B(n6137), .ZN(n6480) );
  OR2_X1 U6147 ( .A1(n8263), .A2(n8609), .ZN(n4452) );
  AND2_X1 U6148 ( .A1(n4871), .A2(n9911), .ZN(n4453) );
  INV_X1 U6149 ( .A(n8551), .ZN(n5114) );
  XNOR2_X1 U6150 ( .A(n5325), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6242) );
  AND2_X1 U6151 ( .A1(n4839), .A2(n4838), .ZN(n4454) );
  AND2_X1 U6152 ( .A1(n7597), .A2(n8476), .ZN(n8416) );
  AND2_X1 U6153 ( .A1(n5202), .A2(n5201), .ZN(n4455) );
  OR2_X1 U6154 ( .A1(n7969), .A2(n10234), .ZN(n4456) );
  NOR2_X1 U6155 ( .A1(n9001), .A2(n8802), .ZN(n4457) );
  OR2_X1 U6156 ( .A1(n5666), .A2(SI_9_), .ZN(n4458) );
  INV_X1 U6157 ( .A(n9683), .ZN(n10014) );
  AND4_X1 U6158 ( .A1(n4464), .A2(n8359), .A3(n7891), .A4(n8000), .ZN(n4459)
         );
  AND2_X1 U6159 ( .A1(n7421), .A2(n10211), .ZN(n4460) );
  AND4_X1 U6160 ( .A1(n5868), .A2(n5448), .A3(n5780), .A4(n5447), .ZN(n4461)
         );
  NAND2_X1 U6161 ( .A1(n5254), .A2(n5253), .ZN(n6559) );
  AND2_X1 U6162 ( .A1(n6774), .A2(n6773), .ZN(n4462) );
  AND2_X1 U6163 ( .A1(n7197), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4463) );
  NAND2_X1 U6164 ( .A1(n7137), .A2(n7136), .ZN(n7138) );
  OR2_X1 U6165 ( .A1(n7888), .A2(n8363), .ZN(n4464) );
  INV_X1 U6166 ( .A(n9689), .ZN(n4661) );
  INV_X1 U6167 ( .A(n10103), .ZN(n7497) );
  INV_X1 U6168 ( .A(n9466), .ZN(n4872) );
  INV_X1 U6169 ( .A(n9554), .ZN(n7714) );
  NOR3_X1 U6170 ( .A1(n8567), .A2(n8433), .A3(n8563), .ZN(n4465) );
  AND2_X1 U6171 ( .A1(n8214), .A2(n10093), .ZN(n4466) );
  AND2_X1 U6172 ( .A1(n9888), .A2(n9468), .ZN(n4467) );
  AND2_X1 U6173 ( .A1(n9690), .A2(n10119), .ZN(n4468) );
  AND2_X1 U6174 ( .A1(n6738), .A2(n6737), .ZN(n4469) );
  AND2_X1 U6175 ( .A1(n7198), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4470) );
  AND2_X1 U6176 ( .A1(n9681), .A2(n4614), .ZN(n4471) );
  INV_X1 U6177 ( .A(n9407), .ZN(n4621) );
  AND3_X1 U6178 ( .A1(n8492), .A2(n8491), .A3(n8490), .ZN(n4472) );
  AND2_X1 U6179 ( .A1(n9007), .A2(n8608), .ZN(n4473) );
  AND2_X1 U6180 ( .A1(n4790), .A2(n4789), .ZN(n4474) );
  OR2_X1 U6181 ( .A1(n4973), .A2(n4975), .ZN(n4475) );
  NAND2_X1 U6182 ( .A1(n5928), .A2(n5927), .ZN(n9960) );
  AND2_X1 U6183 ( .A1(n5159), .A2(n4452), .ZN(n4476) );
  NAND2_X1 U6184 ( .A1(n8298), .A2(n8612), .ZN(n4477) );
  INV_X1 U6185 ( .A(n8257), .ZN(n8802) );
  AND2_X1 U6186 ( .A1(n6464), .A2(n6463), .ZN(n8257) );
  NOR2_X1 U6187 ( .A1(n5224), .A2(n4545), .ZN(n4478) );
  INV_X1 U6188 ( .A(n8534), .ZN(n4817) );
  NAND2_X1 U6189 ( .A1(n7461), .A2(n7555), .ZN(n4479) );
  AND2_X1 U6190 ( .A1(n8405), .A2(n8404), .ZN(n8993) );
  AND2_X1 U6191 ( .A1(n4884), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4480) );
  AND2_X1 U6192 ( .A1(n4909), .A2(n4908), .ZN(n4481) );
  INV_X1 U6193 ( .A(n4774), .ZN(n4773) );
  NAND2_X1 U6194 ( .A1(n4775), .A2(n4777), .ZN(n4774) );
  AND2_X1 U6195 ( .A1(n9382), .A2(n4637), .ZN(n4482) );
  NAND2_X1 U6196 ( .A1(n9346), .A2(n9458), .ZN(n4483) );
  AND2_X1 U6197 ( .A1(n9444), .A2(n9491), .ZN(n9754) );
  INV_X1 U6198 ( .A(n4988), .ZN(n9850) );
  NOR2_X1 U6199 ( .A1(n6101), .A2(n9983), .ZN(n4988) );
  NAND2_X1 U6200 ( .A1(n4932), .A2(n4931), .ZN(n4484) );
  AND2_X1 U6201 ( .A1(n8411), .A2(n8577), .ZN(n4485) );
  AND2_X1 U6202 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n4486) );
  OR2_X1 U6203 ( .A1(n4693), .A2(n6831), .ZN(n4487) );
  AND2_X1 U6204 ( .A1(n4930), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4488) );
  AND2_X1 U6205 ( .A1(n9432), .A2(n9384), .ZN(n4489) );
  AND2_X1 U6206 ( .A1(n6367), .A2(n8519), .ZN(n4490) );
  INV_X1 U6207 ( .A(n8450), .ZN(n5135) );
  AND2_X1 U6208 ( .A1(n9055), .A2(n8916), .ZN(n4491) );
  INV_X1 U6209 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5284) );
  AND2_X1 U6210 ( .A1(n8560), .A2(n8561), .ZN(n8799) );
  AND2_X1 U6211 ( .A1(n6719), .A2(n6718), .ZN(n4492) );
  NOR2_X1 U6212 ( .A1(n8100), .A2(n8793), .ZN(n4493) );
  INV_X1 U6213 ( .A(n4948), .ZN(n4947) );
  NAND2_X1 U6214 ( .A1(n4458), .A2(n5651), .ZN(n4948) );
  AND2_X1 U6215 ( .A1(n8507), .A2(n8506), .ZN(n8425) );
  AND2_X1 U6216 ( .A1(n9723), .A2(n9548), .ZN(n4494) );
  AND2_X1 U6217 ( .A1(n5101), .A2(n8511), .ZN(n4495) );
  INV_X1 U6218 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n10272) );
  OR2_X1 U6219 ( .A1(n6219), .A2(n10238), .ZN(n4496) );
  NOR2_X1 U6220 ( .A1(n9988), .A2(n9867), .ZN(n4497) );
  INV_X1 U6221 ( .A(n8113), .ZN(n4693) );
  INV_X1 U6222 ( .A(n4772), .ZN(n4771) );
  AOI21_X1 U6223 ( .B1(n4773), .B2(n7177), .A(n7393), .ZN(n4772) );
  AND2_X1 U6224 ( .A1(n6075), .A2(n4856), .ZN(n4498) );
  AND2_X1 U6225 ( .A1(n9171), .A2(n9170), .ZN(n4499) );
  INV_X1 U6226 ( .A(n5199), .ZN(n5198) );
  OR2_X1 U6227 ( .A1(n8082), .A2(n5200), .ZN(n5199) );
  AND2_X1 U6228 ( .A1(n5186), .A2(n5185), .ZN(n4500) );
  NAND2_X1 U6229 ( .A1(n5093), .A2(n4451), .ZN(n4501) );
  AND3_X1 U6230 ( .A1(n8576), .A2(n8585), .A3(n8584), .ZN(n4502) );
  INV_X1 U6231 ( .A(n5144), .ZN(n5143) );
  NAND2_X1 U6232 ( .A1(n5282), .A2(n5284), .ZN(n5144) );
  OR2_X1 U6233 ( .A1(n9326), .A2(n9552), .ZN(n4503) );
  INV_X1 U6234 ( .A(n4913), .ZN(n4912) );
  OAI21_X1 U6235 ( .B1(n8672), .B2(n8673), .A(n4916), .ZN(n4913) );
  INV_X1 U6236 ( .A(n9514), .ZN(n4544) );
  OR2_X1 U6237 ( .A1(n9067), .A2(n8056), .ZN(n8511) );
  OR2_X1 U6238 ( .A1(n8503), .A2(n8570), .ZN(n4504) );
  OR2_X1 U6239 ( .A1(n8571), .A2(n8781), .ZN(n8569) );
  AND2_X1 U6240 ( .A1(n9408), .A2(n9415), .ZN(n4505) );
  AND2_X1 U6241 ( .A1(n6679), .A2(n7638), .ZN(n4506) );
  AND2_X1 U6242 ( .A1(n8474), .A2(n4709), .ZN(n4507) );
  AND2_X1 U6243 ( .A1(n9452), .A2(n9450), .ZN(n4508) );
  AND2_X1 U6244 ( .A1(n8487), .A2(n5105), .ZN(n4509) );
  AND2_X1 U6245 ( .A1(n7447), .A2(n9291), .ZN(n4510) );
  AND2_X1 U6246 ( .A1(n7783), .A2(n9202), .ZN(n4511) );
  AND2_X1 U6247 ( .A1(n4693), .A2(n6831), .ZN(n4512) );
  AND2_X1 U6248 ( .A1(n5556), .A2(n5559), .ZN(n4513) );
  AND2_X1 U6249 ( .A1(n4441), .A2(n5018), .ZN(n4514) );
  AND2_X1 U6250 ( .A1(n5014), .A2(n5010), .ZN(n4515) );
  OR2_X1 U6251 ( .A1(n8264), .A2(n8263), .ZN(n4578) );
  AND2_X1 U6252 ( .A1(n8511), .A2(n8507), .ZN(n4516) );
  AND2_X1 U6253 ( .A1(n7199), .A2(n7200), .ZN(n4517) );
  AND2_X1 U6254 ( .A1(n8480), .A2(n4606), .ZN(n4518) );
  AND2_X1 U6255 ( .A1(n8508), .A2(n8923), .ZN(n4519) );
  AND2_X1 U6256 ( .A1(n9635), .A2(n8207), .ZN(n4520) );
  OR2_X1 U6257 ( .A1(n5802), .A2(n5089), .ZN(n4521) );
  INV_X1 U6258 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7087) );
  INV_X1 U6259 ( .A(n5174), .ZN(n5173) );
  OR2_X1 U6260 ( .A1(n8251), .A2(n5175), .ZN(n5174) );
  NAND2_X1 U6261 ( .A1(n6514), .A2(n5133), .ZN(n5132) );
  NAND2_X1 U6262 ( .A1(n10181), .A2(n7354), .ZN(n8934) );
  XNOR2_X1 U6263 ( .A(n5251), .B(n5250), .ZN(n6560) );
  NAND2_X1 U6264 ( .A1(n7706), .A2(n4994), .ZN(n7720) );
  INV_X1 U6265 ( .A(n8673), .ZN(n4914) );
  NAND2_X1 U6266 ( .A1(n4707), .A2(n4705), .ZN(n7600) );
  NAND2_X1 U6267 ( .A1(n6074), .A2(n9449), .ZN(n7490) );
  NAND2_X1 U6268 ( .A1(n7430), .A2(n6231), .ZN(n7431) );
  INV_X1 U6269 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4970) );
  AND2_X1 U6270 ( .A1(n6594), .A2(n6592), .ZN(n6595) );
  OR2_X1 U6271 ( .A1(n6101), .A2(n4987), .ZN(n4522) );
  INV_X1 U6272 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n4919) );
  AOI21_X1 U6273 ( .B1(n7686), .B2(n6297), .A(n5212), .ZN(n7698) );
  NAND2_X1 U6274 ( .A1(n6515), .A2(n8507), .ZN(n8922) );
  NAND2_X1 U6275 ( .A1(n5132), .A2(n8500), .ZN(n7697) );
  NAND2_X1 U6276 ( .A1(n4708), .A2(n6252), .ZN(n7468) );
  NAND2_X1 U6277 ( .A1(n6517), .A2(n8519), .ZN(n8896) );
  NAND2_X1 U6278 ( .A1(n5099), .A2(n8511), .ZN(n8913) );
  NAND2_X1 U6279 ( .A1(n6514), .A2(n8494), .ZN(n7684) );
  NAND2_X1 U6280 ( .A1(n5970), .A2(n5969), .ZN(n9950) );
  INV_X1 U6281 ( .A(n9950), .ZN(n5002) );
  INV_X1 U6282 ( .A(n8834), .ZN(n4728) );
  NAND2_X1 U6283 ( .A1(n7589), .A2(n7588), .ZN(n7854) );
  INV_X1 U6284 ( .A(n5259), .ZN(n5186) );
  NAND2_X1 U6285 ( .A1(n6562), .A2(n5206), .ZN(n7134) );
  INV_X1 U6286 ( .A(n8313), .ZN(n8916) );
  INV_X1 U6287 ( .A(n8867), .ZN(n8838) );
  AND2_X1 U6288 ( .A1(n6380), .A2(n6379), .ZN(n8867) );
  INV_X1 U6289 ( .A(n6896), .ZN(n4930) );
  INV_X1 U6290 ( .A(n4753), .ZN(n4752) );
  NAND2_X1 U6291 ( .A1(n4761), .A2(n5394), .ZN(n4753) );
  AND2_X1 U6292 ( .A1(n5338), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4523) );
  INV_X1 U6293 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10445) );
  NAND3_X1 U6294 ( .A1(n5186), .A2(n5184), .A3(n5185), .ZN(n4524) );
  INV_X1 U6295 ( .A(n4847), .ZN(n5847) );
  INV_X1 U6296 ( .A(n4754), .ZN(n4751) );
  NAND2_X1 U6297 ( .A1(n4756), .A2(n5398), .ZN(n4754) );
  AND2_X1 U6298 ( .A1(n4438), .A2(n5338), .ZN(n4525) );
  INV_X1 U6299 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n4927) );
  INV_X1 U6300 ( .A(SI_20_), .ZN(n10446) );
  AND2_X1 U6301 ( .A1(n4794), .A2(n10502), .ZN(n4526) );
  AND2_X1 U6302 ( .A1(n4792), .A2(n4791), .ZN(n4527) );
  AND2_X1 U6303 ( .A1(n4911), .A2(n4914), .ZN(n4528) );
  NAND2_X1 U6304 ( .A1(n6503), .A2(n6880), .ZN(n10171) );
  AND2_X1 U6305 ( .A1(n5221), .A2(n6918), .ZN(n4529) );
  NAND2_X1 U6306 ( .A1(n9402), .A2(n9399), .ZN(n9918) );
  INV_X1 U6307 ( .A(n10155), .ZN(n10154) );
  AND2_X2 U6308 ( .A1(n6166), .A2(n6165), .ZN(n10155) );
  NOR2_X1 U6309 ( .A1(n6912), .A2(n4899), .ZN(n6910) );
  INV_X1 U6310 ( .A(n10003), .ZN(n4995) );
  AND2_X1 U6311 ( .A1(n7653), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4530) );
  NAND2_X1 U6312 ( .A1(n7426), .A2(n8486), .ZN(n10162) );
  AND2_X2 U6313 ( .A1(n7075), .A2(n6585), .ZN(n10245) );
  INV_X1 U6314 ( .A(n7343), .ZN(n5151) );
  INV_X1 U6315 ( .A(n6601), .ZN(n7378) );
  AND2_X1 U6316 ( .A1(n8203), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4531) );
  AND2_X1 U6317 ( .A1(n4776), .A2(n4773), .ZN(n4532) );
  INV_X1 U6318 ( .A(n10067), .ZN(n10093) );
  INV_X1 U6319 ( .A(n4763), .ZN(n7536) );
  NOR2_X1 U6320 ( .A1(n9651), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4533) );
  AND2_X1 U6321 ( .A1(n5323), .A2(n7017), .ZN(n4534) );
  AND2_X1 U6322 ( .A1(n10154), .A2(n6590), .ZN(n4535) );
  NAND2_X1 U6323 ( .A1(n8741), .A2(n5442), .ZN(n4536) );
  INV_X1 U6324 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4853) );
  NAND2_X1 U6325 ( .A1(n4921), .A2(n6928), .ZN(n7210) );
  XNOR2_X1 U6326 ( .A(n6502), .B(n6501), .ZN(n8585) );
  XOR2_X1 U6327 ( .A(n6274), .B(P2_REG2_REG_8__SCAN_IN), .Z(n4537) );
  XOR2_X1 U6328 ( .A(n6242), .B(P2_REG2_REG_6__SCAN_IN), .Z(n4538) );
  NAND2_X1 U6329 ( .A1(n9606), .A2(n9607), .ZN(n4841) );
  INV_X2 U6330 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5071) );
  INV_X1 U6331 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4967) );
  NAND2_X1 U6332 ( .A1(n5713), .A2(n5534), .ZN(n9580) );
  INV_X1 U6333 ( .A(n9580), .ZN(n4698) );
  INV_X1 U6334 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n4634) );
  INV_X1 U6335 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4620) );
  INV_X1 U6336 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n4601) );
  INV_X1 U6337 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n4655) );
  INV_X1 U6338 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n4636) );
  INV_X1 U6339 ( .A(n8717), .ZN(n4571) );
  NAND2_X1 U6340 ( .A1(n9129), .A2(n4694), .ZN(n5075) );
  NAND2_X2 U6341 ( .A1(n9803), .A2(n9440), .ZN(n9790) );
  NAND2_X1 U6342 ( .A1(n5615), .A2(n4540), .ZN(n5616) );
  NAND2_X1 U6343 ( .A1(n5075), .A2(n5073), .ZN(n6804) );
  NAND2_X1 U6344 ( .A1(n4934), .A2(n5563), .ZN(n5615) );
  INV_X1 U6345 ( .A(n4553), .ZN(n4552) );
  NAND2_X1 U6346 ( .A1(n5584), .A2(n4651), .ZN(n4541) );
  NAND2_X1 U6347 ( .A1(n7906), .A2(n8506), .ZN(n6515) );
  NAND2_X1 U6348 ( .A1(n6026), .A2(n6025), .ZN(n6038) );
  NAND2_X1 U6349 ( .A1(n4547), .A2(n6007), .ZN(n6024) );
  NAND2_X1 U6350 ( .A1(n4972), .A2(n4971), .ZN(n5922) );
  NAND2_X1 U6351 ( .A1(n6006), .A2(n6005), .ZN(n4547) );
  OAI21_X1 U6352 ( .B1(n5610), .B2(n5611), .A(n5609), .ZN(n5612) );
  NAND2_X1 U6353 ( .A1(n5566), .A2(SI_5_), .ZN(n5610) );
  OAI211_X1 U6354 ( .C1(n4857), .C2(n6074), .A(n4855), .B(n4854), .ZN(n7710)
         );
  NAND2_X2 U6355 ( .A1(n4864), .A2(n4489), .ZN(n9716) );
  OAI21_X2 U6356 ( .B1(n7862), .B2(n4870), .A(n4552), .ZN(n8234) );
  INV_X1 U6357 ( .A(n9853), .ZN(n4549) );
  NAND2_X2 U6358 ( .A1(n4848), .A2(n4850), .ZN(n6601) );
  NAND2_X2 U6359 ( .A1(n6157), .A2(n9578), .ZN(n5543) );
  XNOR2_X2 U6360 ( .A(n5466), .B(P1_IR_REG_29__SCAN_IN), .ZN(n10056) );
  NAND2_X1 U6361 ( .A1(n4622), .A2(n4621), .ZN(n7862) );
  NAND2_X1 U6362 ( .A1(n7710), .A2(n9344), .ZN(n7722) );
  NAND2_X1 U6363 ( .A1(n6077), .A2(n9348), .ZN(n7863) );
  AOI21_X1 U6364 ( .B1(n9688), .B2(n6146), .A(n6160), .ZN(n4867) );
  AOI21_X1 U6365 ( .B1(n4609), .B2(n7441), .A(n4435), .ZN(n5546) );
  NAND2_X1 U6366 ( .A1(n9752), .A2(n5980), .ZN(n9731) );
  NAND2_X1 U6367 ( .A1(n7662), .A2(n7668), .ZN(n7661) );
  OAI21_X1 U6368 ( .B1(n9861), .B2(n5858), .A(n5857), .ZN(n9839) );
  NAND2_X1 U6369 ( .A1(n5468), .A2(n5469), .ZN(n9560) );
  INV_X2 U6370 ( .A(n9560), .ZN(n8129) );
  NAND2_X1 U6371 ( .A1(n7797), .A2(n8451), .ZN(n7906) );
  NAND2_X1 U6372 ( .A1(n5108), .A2(n5109), .ZN(n4550) );
  NAND2_X1 U6373 ( .A1(n5104), .A2(n4509), .ZN(n7455) );
  NAND2_X2 U6374 ( .A1(n7574), .A2(n7575), .ZN(n7573) );
  NOR2_X1 U6375 ( .A1(n7012), .A2(n5422), .ZN(n5423) );
  NOR2_X1 U6376 ( .A1(n6982), .A2(n6983), .ZN(n6981) );
  NAND3_X1 U6377 ( .A1(n4778), .A2(n4596), .A3(n5445), .ZN(P2_U3201) );
  NOR2_X1 U6378 ( .A1(n5417), .A2(n7159), .ZN(n5419) );
  NAND2_X1 U6379 ( .A1(n9611), .A2(n9610), .ZN(n7046) );
  NAND2_X1 U6380 ( .A1(n7043), .A2(n7042), .ZN(n9611) );
  OAI21_X1 U6381 ( .B1(n7292), .B2(n7285), .A(n4517), .ZN(n7290) );
  NAND2_X1 U6382 ( .A1(n9585), .A2(n9584), .ZN(n9599) );
  NAND2_X1 U6383 ( .A1(n9566), .A2(n9567), .ZN(n9565) );
  NAND2_X1 U6384 ( .A1(n4833), .A2(n9920), .ZN(n4832) );
  NAND2_X1 U6385 ( .A1(n8212), .A2(n9663), .ZN(n4834) );
  XNOR2_X1 U6386 ( .A(n5522), .B(n5521), .ZN(n7037) );
  NOR2_X1 U6387 ( .A1(n4466), .A2(n8213), .ZN(n4835) );
  OR2_X1 U6388 ( .A1(n8191), .A2(n8190), .ZN(n8192) );
  NAND2_X1 U6389 ( .A1(n9592), .A2(n7033), .ZN(n9606) );
  NOR2_X1 U6390 ( .A1(n9622), .A2(n10368), .ZN(n9621) );
  OAI21_X1 U6391 ( .B1(n8214), .B2(n10067), .A(n4834), .ZN(n4833) );
  XNOR2_X1 U6392 ( .A(n8201), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n8212) );
  NOR3_X1 U6393 ( .A1(n10070), .A2(n7202), .A3(n7204), .ZN(n7316) );
  NAND2_X1 U6394 ( .A1(n9833), .A2(n9834), .ZN(n6081) );
  OR2_X2 U6395 ( .A1(n10008), .A2(n9899), .ZN(n9468) );
  OAI21_X1 U6396 ( .B1(n4870), .B2(n6078), .A(n6079), .ZN(n4553) );
  NAND2_X1 U6397 ( .A1(n9851), .A2(n9479), .ZN(n9833) );
  NAND2_X1 U6398 ( .A1(n8221), .A2(n9428), .ZN(n8220) );
  NAND2_X1 U6399 ( .A1(n6089), .A2(n9403), .ZN(n6152) );
  INV_X1 U6400 ( .A(n8687), .ZN(n4554) );
  NAND2_X1 U6401 ( .A1(n4558), .A2(n5434), .ZN(n8687) );
  NOR2_X1 U6402 ( .A1(n6996), .A2(n10232), .ZN(n6995) );
  NAND2_X1 U6403 ( .A1(n6914), .A2(n5207), .ZN(n5425) );
  NAND2_X1 U6404 ( .A1(n4873), .A2(n7540), .ZN(n4874) );
  NAND2_X1 U6405 ( .A1(n4436), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4555) );
  NAND2_X1 U6406 ( .A1(n6180), .A2(n4555), .ZN(n5413) );
  NAND2_X1 U6407 ( .A1(n4559), .A2(n8695), .ZN(n4558) );
  INV_X1 U6408 ( .A(n5433), .ZN(n4559) );
  NAND2_X2 U6409 ( .A1(n5484), .A2(n5478), .ZN(n5539) );
  NAND2_X1 U6410 ( .A1(n5567), .A2(n10294), .ZN(n5613) );
  NAND2_X1 U6411 ( .A1(n4513), .A2(n5557), .ZN(n4934) );
  NAND2_X1 U6412 ( .A1(n9941), .A2(n10136), .ZN(n4560) );
  NOR2_X1 U6413 ( .A1(n9939), .A2(n9940), .ZN(n4561) );
  NAND2_X1 U6414 ( .A1(n4562), .A2(n4813), .ZN(n8509) );
  NAND3_X1 U6415 ( .A1(n8502), .A2(n4812), .A3(n4810), .ZN(n4562) );
  OAI21_X1 U6416 ( .B1(n4472), .B2(n4563), .A(n8499), .ZN(n8501) );
  NAND2_X1 U6417 ( .A1(n4566), .A2(n4565), .ZN(n8532) );
  INV_X1 U6418 ( .A(n8525), .ZN(n4566) );
  AOI21_X1 U6419 ( .B1(n5341), .B2(n8656), .A(n5342), .ZN(n8657) );
  NAND2_X1 U6420 ( .A1(n4863), .A2(n4445), .ZN(n6073) );
  INV_X1 U6421 ( .A(n6072), .ZN(n4687) );
  NAND2_X1 U6422 ( .A1(n6088), .A2(n9497), .ZN(n6089) );
  NAND2_X2 U6424 ( .A1(n4744), .A2(n5262), .ZN(n5281) );
  AND2_X2 U6425 ( .A1(n5261), .A2(n5289), .ZN(n4744) );
  OAI21_X2 U6426 ( .B1(n8179), .B2(n8567), .A(n6529), .ZN(n6554) );
  NAND2_X1 U6427 ( .A1(n8416), .A2(n5141), .ZN(n5140) );
  NOR2_X2 U6428 ( .A1(n5259), .A2(n5263), .ZN(n5262) );
  BUF_X4 U6429 ( .A(n6174), .Z(n6544) );
  NAND2_X1 U6430 ( .A1(n8832), .A2(n8539), .ZN(n6524) );
  NAND2_X1 U6431 ( .A1(n5431), .A2(n7086), .ZN(n5432) );
  NAND3_X1 U6432 ( .A1(n4894), .A2(n4893), .A3(n5430), .ZN(n5431) );
  INV_X1 U6433 ( .A(n7307), .ZN(n7306) );
  AOI22_X2 U6434 ( .A1(n8273), .A2(n8272), .B1(n8880), .B2(n8086), .ZN(n8341)
         );
  NAND3_X1 U6435 ( .A1(n5632), .A2(n4945), .A3(n4943), .ZN(n4579) );
  NAND2_X1 U6436 ( .A1(n7966), .A2(n8612), .ZN(n8451) );
  NAND2_X1 U6437 ( .A1(n6975), .A2(n8402), .ZN(n4829) );
  NAND2_X1 U6438 ( .A1(n5616), .A2(n5617), .ZN(n5622) );
  NOR3_X1 U6439 ( .A1(n8600), .A2(n8596), .A3(n8595), .ZN(n8597) );
  MUX2_X1 U6440 ( .A(n8473), .B(n8472), .S(n8570), .Z(n8497) );
  NAND2_X1 U6441 ( .A1(n4608), .A2(n4581), .ZN(n5484) );
  NOR2_X1 U6442 ( .A1(n4580), .A2(n8483), .ZN(n4604) );
  NAND2_X1 U6443 ( .A1(n4582), .A2(n6926), .ZN(n4581) );
  NAND2_X2 U6444 ( .A1(n5622), .A2(n5621), .ZN(n5632) );
  NAND2_X1 U6445 ( .A1(n5501), .A2(n5500), .ZN(n5559) );
  INV_X2 U6446 ( .A(n5584), .ZN(n6929) );
  OAI21_X2 U6447 ( .B1(n9824), .B2(n5898), .A(n5899), .ZN(n9808) );
  NAND2_X1 U6448 ( .A1(n7488), .A2(n5600), .ZN(n7746) );
  NAND2_X1 U6449 ( .A1(n4605), .A2(n4603), .ZN(n4812) );
  NAND2_X1 U6450 ( .A1(n4585), .A2(n4583), .ZN(P1_U3356) );
  NOR2_X1 U6451 ( .A1(n4468), .A2(n4584), .ZN(n4583) );
  NAND2_X1 U6452 ( .A1(n4587), .A2(n9776), .ZN(n4585) );
  NAND2_X2 U6453 ( .A1(n10008), .A2(n9899), .ZN(n9466) );
  NOR2_X1 U6454 ( .A1(n8112), .A2(n4692), .ZN(n8120) );
  NAND2_X1 U6455 ( .A1(n9716), .A2(n9715), .ZN(n4626) );
  NAND2_X1 U6456 ( .A1(n6892), .A2(n6891), .ZN(n4894) );
  NAND2_X1 U6457 ( .A1(n4898), .A2(n6911), .ZN(n6914) );
  NAND2_X1 U6458 ( .A1(n8662), .A2(n4586), .ZN(n5433) );
  NAND2_X1 U6459 ( .A1(n8622), .A2(n5427), .ZN(n5428) );
  NOR2_X1 U6460 ( .A1(n6995), .A2(n5415), .ZN(n6982) );
  AND2_X4 U6461 ( .A1(n10056), .A2(n4669), .ZN(n5551) );
  INV_X1 U6462 ( .A(n7948), .ZN(n9559) );
  NAND2_X1 U6463 ( .A1(n4868), .A2(n4869), .ZN(n4587) );
  NAND2_X1 U6464 ( .A1(n7771), .A2(n9292), .ZN(n6074) );
  NAND2_X1 U6465 ( .A1(n4667), .A2(n9496), .ZN(n4666) );
  NAND3_X1 U6466 ( .A1(n4588), .A2(n9361), .A3(n9360), .ZN(n9362) );
  NAND2_X1 U6467 ( .A1(n9478), .A2(n9381), .ZN(n4590) );
  INV_X1 U6468 ( .A(n4871), .ZN(n4870) );
  NAND2_X1 U6469 ( .A1(n8482), .A2(n4518), .ZN(n4605) );
  NAND2_X1 U6470 ( .A1(n4593), .A2(n8570), .ZN(n4592) );
  NAND2_X1 U6471 ( .A1(n4592), .A2(n4591), .ZN(n8466) );
  NAND3_X1 U6472 ( .A1(n8457), .A2(n8456), .A3(n8467), .ZN(n4593) );
  NAND2_X1 U6473 ( .A1(n4595), .A2(n4594), .ZN(n8522) );
  NAND2_X1 U6474 ( .A1(n8514), .A2(n5052), .ZN(n4595) );
  AOI21_X1 U6475 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n7653), .A(n7650), .ZN(
        n8191) );
  AOI21_X1 U6476 ( .B1(n6918), .B2(n4927), .A(n4537), .ZN(n4925) );
  INV_X1 U6477 ( .A(n5221), .ZN(n4924) );
  NAND3_X1 U6478 ( .A1(n7210), .A2(n4920), .A3(P2_REG2_REG_3__SCAN_IN), .ZN(
        n7212) );
  NAND2_X1 U6479 ( .A1(n4933), .A2(n5350), .ZN(n4932) );
  NAND2_X1 U6480 ( .A1(n6605), .A2(n6606), .ZN(n8125) );
  INV_X1 U6481 ( .A(n9132), .ZN(n4695) );
  NAND2_X1 U6482 ( .A1(n4963), .A2(SI_14_), .ZN(n4962) );
  OAI21_X2 U6483 ( .B1(n9839), .B2(n5884), .A(n4597), .ZN(n9824) );
  OAI21_X2 U6484 ( .B1(n4951), .B2(n4639), .A(n5828), .ZN(n5845) );
  NAND3_X1 U6485 ( .A1(n4649), .A2(n4648), .A3(n4647), .ZN(n6169) );
  OAI21_X1 U6486 ( .B1(n8527), .B2(n8526), .A(n8538), .ZN(n8528) );
  NAND3_X1 U6487 ( .A1(n8470), .A2(n8487), .A3(n4479), .ZN(n8475) );
  NAND2_X1 U6488 ( .A1(n4602), .A2(n8512), .ZN(n8514) );
  NAND2_X1 U6489 ( .A1(n8509), .A2(n4519), .ZN(n4602) );
  AND2_X1 U6490 ( .A1(n4485), .A2(n4604), .ZN(n4603) );
  NAND2_X2 U6491 ( .A1(n6203), .A2(n4607), .ZN(n6204) );
  AOI21_X1 U6492 ( .B1(n8522), .B2(n8521), .A(n8520), .ZN(n8525) );
  XNOR2_X2 U6493 ( .A(n5496), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9596) );
  OAI211_X1 U6494 ( .C1(n4835), .C2(n9920), .A(n4832), .B(n4830), .ZN(P1_U3262) );
  NAND2_X2 U6495 ( .A1(n9468), .A2(n9466), .ZN(n9925) );
  OAI21_X2 U6496 ( .B1(n9699), .B2(n9701), .A(n6036), .ZN(n6054) );
  OAI21_X2 U6497 ( .B1(n7748), .B2(n5030), .A(n5029), .ZN(n7662) );
  AOI21_X1 U6498 ( .B1(n4866), .B2(n9893), .A(n4535), .ZN(n4865) );
  NAND2_X1 U6499 ( .A1(n5034), .A2(n5033), .ZN(n9752) );
  INV_X1 U6500 ( .A(n9414), .ZN(n4609) );
  NAND2_X1 U6501 ( .A1(n4865), .A2(n4610), .ZN(n6591) );
  NAND2_X1 U6502 ( .A1(n4866), .A2(n4611), .ZN(n4610) );
  INV_X1 U6503 ( .A(n6161), .ZN(n4611) );
  AND3_X2 U6504 ( .A1(n4867), .A2(n6162), .A3(n10155), .ZN(n4866) );
  NAND2_X1 U6505 ( .A1(n4515), .A2(n4612), .ZN(n9861) );
  OAI21_X2 U6506 ( .B1(n9808), .B2(n5917), .A(n5916), .ZN(n9783) );
  NAND2_X1 U6507 ( .A1(n9887), .A2(n4514), .ZN(n4612) );
  NAND2_X1 U6508 ( .A1(n5043), .A2(n5042), .ZN(P1_U3550) );
  NAND2_X1 U6509 ( .A1(n4613), .A2(n10136), .ZN(n4648) );
  INV_X1 U6510 ( .A(n8249), .ZN(n4613) );
  NAND2_X1 U6511 ( .A1(n9688), .A2(n6055), .ZN(n8249) );
  AOI21_X1 U6512 ( .B1(n9682), .B2(n9683), .A(n9907), .ZN(n4614) );
  NAND2_X1 U6513 ( .A1(n9397), .A2(n9396), .ZN(n4689) );
  NAND2_X1 U6514 ( .A1(n5577), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U6515 ( .A1(n9398), .A2(n4939), .ZN(n4938) );
  NAND2_X1 U6516 ( .A1(n9390), .A2(n9391), .ZN(n4668) );
  INV_X1 U6517 ( .A(n7863), .ZN(n4622) );
  NAND2_X2 U6518 ( .A1(n9316), .A2(n9321), .ZN(n6076) );
  NAND2_X1 U6519 ( .A1(n4629), .A2(n4627), .ZN(P1_U3548) );
  OR2_X1 U6520 ( .A1(n10019), .A2(n10159), .ZN(n4629) );
  INV_X4 U6521 ( .A(n5676), .ZN(n5505) );
  INV_X1 U6522 ( .A(n4801), .ZN(n4799) );
  NAND2_X1 U6523 ( .A1(n5281), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6524 ( .A1(n6558), .A2(n4657), .ZN(n6889) );
  INV_X1 U6525 ( .A(n5706), .ZN(n4802) );
  NAND2_X1 U6526 ( .A1(n4938), .A2(n4937), .ZN(n9439) );
  NAND2_X1 U6527 ( .A1(n5757), .A2(n4959), .ZN(n4958) );
  NAND2_X1 U6528 ( .A1(n9383), .A2(n4482), .ZN(n9389) );
  INV_X1 U6529 ( .A(n9501), .ZN(n4638) );
  NAND2_X2 U6530 ( .A1(n8744), .A2(n8743), .ZN(n5439) );
  AND2_X1 U6531 ( .A1(n6994), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4640) );
  AND3_X4 U6532 ( .A1(n4461), .A2(n5453), .A3(n5452), .ZN(n6056) );
  NAND4_X2 U6533 ( .A1(n6056), .A2(n4643), .A3(n4684), .A4(n4430), .ZN(n10045)
         );
  OAI21_X2 U6534 ( .B1(n5281), .B2(n5144), .A(n5352), .ZN(n5065) );
  NAND2_X1 U6535 ( .A1(n5121), .A2(n5124), .ZN(n7797) );
  NAND2_X1 U6536 ( .A1(n5138), .A2(n5136), .ZN(n7626) );
  NAND3_X1 U6537 ( .A1(n4733), .A2(n10245), .A3(n4738), .ZN(n4642) );
  NAND2_X1 U6538 ( .A1(n7746), .A2(n9299), .ZN(n7748) );
  AND2_X2 U6539 ( .A1(n4683), .A2(n5460), .ZN(n4643) );
  AND3_X4 U6540 ( .A1(n5495), .A2(n5494), .A3(n5493), .ZN(n10132) );
  NAND2_X4 U6541 ( .A1(n4969), .A2(n4968), .ZN(n5584) );
  XNOR2_X2 U6542 ( .A(n5668), .B(n5667), .ZN(n6958) );
  NAND2_X1 U6543 ( .A1(n4958), .A2(n5776), .ZN(n4957) );
  OAI21_X1 U6544 ( .B1(n8144), .B2(P1_DATAO_REG_13__SCAN_IN), .A(n4645), .ZN(
        n5733) );
  NOR2_X1 U6545 ( .A1(n8594), .A2(n8593), .ZN(n8600) );
  NAND2_X2 U6546 ( .A1(n9458), .A2(n9344), .ZN(n9419) );
  OAI22_X1 U6547 ( .A1(n8151), .A2(n6944), .B1(n5543), .B2(n9608), .ZN(n4653)
         );
  INV_X1 U6548 ( .A(n4803), .ZN(n4800) );
  NAND2_X1 U6549 ( .A1(n4864), .A2(n9384), .ZN(n9714) );
  NAND2_X1 U6550 ( .A1(n5687), .A2(n5686), .ZN(n5707) );
  NAND2_X1 U6551 ( .A1(n5599), .A2(n5598), .ZN(n7488) );
  NAND2_X1 U6552 ( .A1(n9343), .A2(n9342), .ZN(n9345) );
  NAND2_X1 U6553 ( .A1(n4658), .A2(n9322), .ZN(n9343) );
  NAND2_X1 U6554 ( .A1(n4659), .A2(n9318), .ZN(n4658) );
  NAND4_X1 U6555 ( .A1(n9311), .A2(n9310), .A3(n9313), .A4(n9312), .ZN(n4659)
         );
  AOI21_X1 U6556 ( .B1(n4666), .B2(n4664), .A(n9389), .ZN(n4663) );
  INV_X2 U6557 ( .A(n5467), .ZN(n4669) );
  NAND2_X1 U6558 ( .A1(n4673), .A2(n4671), .ZN(n9352) );
  NAND2_X1 U6559 ( .A1(n9347), .A2(n4672), .ZN(n4671) );
  AND2_X1 U6560 ( .A1(n4467), .A2(n4677), .ZN(n4672) );
  AOI21_X1 U6561 ( .B1(n4675), .B2(n4467), .A(n4674), .ZN(n4673) );
  AOI21_X1 U6562 ( .B1(n4679), .B2(n4483), .A(n9909), .ZN(n4677) );
  NAND2_X1 U6563 ( .A1(n4680), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5463) );
  NAND4_X1 U6564 ( .A1(n4681), .A2(n4682), .A3(n4684), .A4(n6056), .ZN(n4680)
         );
  NOR2_X2 U6565 ( .A1(n5457), .A2(n5713), .ZN(n5470) );
  INV_X2 U6566 ( .A(n5713), .ZN(n4683) );
  NAND2_X1 U6567 ( .A1(n7365), .A2(n9452), .ZN(n4688) );
  NAND2_X1 U6568 ( .A1(n4688), .A2(n4686), .ZN(n4685) );
  NAND2_X1 U6569 ( .A1(n4685), .A2(n9450), .ZN(n9296) );
  NAND2_X1 U6570 ( .A1(n5086), .A2(n4442), .ZN(n9265) );
  AND2_X2 U6571 ( .A1(n9265), .A2(n4512), .ZN(n8112) );
  NAND2_X4 U6572 ( .A1(n4434), .A2(n6929), .ZN(n8151) );
  NAND2_X1 U6573 ( .A1(n6749), .A2(n4700), .ZN(n9117) );
  NAND2_X1 U6574 ( .A1(n9117), .A2(n6771), .ZN(n5096) );
  NOR2_X1 U6575 ( .A1(n7640), .A2(n4703), .ZN(n4702) );
  NAND2_X1 U6576 ( .A1(n7643), .A2(n4506), .ZN(n6685) );
  NAND3_X1 U6577 ( .A1(n6056), .A2(n5470), .A3(n4430), .ZN(n6114) );
  AND4_X2 U6578 ( .A1(n6056), .A2(n5470), .A3(n4430), .A4(n4704), .ZN(n6108)
         );
  NAND3_X1 U6579 ( .A1(n8474), .A2(n4709), .A3(n4711), .ZN(n4706) );
  NAND2_X1 U6580 ( .A1(n7456), .A2(n4507), .ZN(n4707) );
  NAND2_X1 U6581 ( .A1(n8924), .A2(n4716), .ZN(n4712) );
  NAND2_X1 U6582 ( .A1(n4712), .A2(n4713), .ZN(n8898) );
  NAND2_X1 U6583 ( .A1(n4722), .A2(n4720), .ZN(n8824) );
  NAND2_X1 U6584 ( .A1(n8878), .A2(n4723), .ZN(n4722) );
  NAND2_X1 U6585 ( .A1(n4731), .A2(n4729), .ZN(n5062) );
  XNOR2_X1 U6586 ( .A(n8780), .B(n4736), .ZN(n4732) );
  NOR2_X1 U6587 ( .A1(n4740), .A2(n4737), .ZN(n4733) );
  NAND2_X1 U6588 ( .A1(n4738), .A2(n8783), .ZN(n8938) );
  NAND2_X1 U6589 ( .A1(n4738), .A2(n4734), .ZN(n4739) );
  NAND3_X1 U6590 ( .A1(n4744), .A2(n5262), .A3(n5282), .ZN(n4745) );
  NAND2_X1 U6591 ( .A1(n4747), .A2(n4748), .ZN(n8689) );
  NAND2_X1 U6592 ( .A1(n6899), .A2(n4750), .ZN(n4747) );
  NAND2_X1 U6593 ( .A1(n4755), .A2(n4756), .ZN(n8680) );
  MUX2_X1 U6594 ( .A(P2_REG1_REG_1__SCAN_IN), .B(P2_REG2_REG_1__SCAN_IN), .S(
        n6539), .Z(n5367) );
  MUX2_X1 U6595 ( .A(n5411), .B(n6185), .S(n6539), .Z(n5366) );
  MUX2_X1 U6596 ( .A(P2_REG1_REG_2__SCAN_IN), .B(P2_REG2_REG_2__SCAN_IN), .S(
        n6539), .Z(n5368) );
  MUX2_X1 U6597 ( .A(P2_REG1_REG_3__SCAN_IN), .B(P2_REG2_REG_3__SCAN_IN), .S(
        n6539), .Z(n5371) );
  MUX2_X1 U6598 ( .A(P2_REG1_REG_4__SCAN_IN), .B(P2_REG2_REG_4__SCAN_IN), .S(
        n6539), .Z(n5372) );
  MUX2_X1 U6599 ( .A(P2_REG1_REG_5__SCAN_IN), .B(P2_REG2_REG_5__SCAN_IN), .S(
        n6539), .Z(n5373) );
  MUX2_X1 U6600 ( .A(n10242), .B(n7458), .S(n6539), .Z(n5375) );
  MUX2_X1 U6601 ( .A(n7563), .B(n4927), .S(n6539), .Z(n5377) );
  MUX2_X1 U6602 ( .A(P2_REG1_REG_0__SCAN_IN), .B(P2_REG2_REG_0__SCAN_IN), .S(
        n6539), .Z(n6965) );
  OAI21_X1 U6603 ( .B1(n7178), .B2(n4768), .A(n4764), .ZN(n4763) );
  NAND3_X1 U6604 ( .A1(n10293), .A2(n4783), .A3(n6232), .ZN(n6245) );
  INV_X1 U6605 ( .A(n5110), .ZN(n8556) );
  NAND2_X1 U6606 ( .A1(n6343), .A2(n4527), .ZN(n6383) );
  NAND2_X1 U6607 ( .A1(n6374), .A2(n4526), .ZN(n6412) );
  NAND3_X2 U6608 ( .A1(n5477), .A2(n4796), .A3(n4797), .ZN(n4969) );
  NAND2_X1 U6609 ( .A1(n4806), .A2(n8790), .ZN(n4805) );
  NAND2_X1 U6610 ( .A1(n4807), .A2(n8562), .ZN(n4806) );
  NAND3_X1 U6611 ( .A1(n4809), .A2(n4808), .A3(n8799), .ZN(n4807) );
  NAND2_X1 U6612 ( .A1(n8559), .A2(n8570), .ZN(n4808) );
  NAND2_X1 U6613 ( .A1(n8558), .A2(n8577), .ZN(n4809) );
  NAND2_X1 U6614 ( .A1(n4504), .A2(n4811), .ZN(n4810) );
  OR2_X1 U6615 ( .A1(n8525), .A2(n4815), .ZN(n4814) );
  NAND2_X1 U6616 ( .A1(n4814), .A2(n4816), .ZN(n8537) );
  NAND3_X1 U6617 ( .A1(n4824), .A2(n4822), .A3(n4502), .ZN(n8594) );
  NAND3_X1 U6618 ( .A1(n8575), .A2(n8583), .A3(n8581), .ZN(n4825) );
  NAND3_X1 U6619 ( .A1(n4828), .A2(n8822), .A3(n4826), .ZN(n8545) );
  NAND3_X1 U6620 ( .A1(n4827), .A2(n8570), .A3(n8541), .ZN(n4826) );
  NAND3_X1 U6621 ( .A1(n8540), .A2(n8538), .A3(n8539), .ZN(n4827) );
  NAND2_X1 U6622 ( .A1(n9638), .A2(n4845), .ZN(n4844) );
  NAND2_X1 U6623 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n10061), .ZN(n5521) );
  NAND2_X1 U6624 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5464) );
  NAND2_X1 U6625 ( .A1(n5761), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U6626 ( .A1(n6112), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U6627 ( .A1(n6114), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6115) );
  OAI21_X1 U6628 ( .B1(n6112), .B2(n6111), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6113) );
  NAND2_X1 U6629 ( .A1(n5677), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U6630 ( .A1(n5802), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5781) );
  NOR2_X1 U6631 ( .A1(n10046), .A2(n5871), .ZN(n4846) );
  NAND2_X1 U6632 ( .A1(n5875), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4847) );
  NAND2_X1 U6633 ( .A1(n5678), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U6634 ( .A1(n5782), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U6635 ( .A1(n5690), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5691) );
  XNOR2_X2 U6636 ( .A(n7411), .B(n6601), .ZN(n9416) );
  OAI22_X1 U6637 ( .A1(n5676), .A2(n6936), .B1(n5543), .B2(n7037), .ZN(n4849)
         );
  NAND2_X2 U6638 ( .A1(n4433), .A2(n8144), .ZN(n5676) );
  NAND4_X2 U6639 ( .A1(n5519), .A2(n4851), .A3(n5518), .A4(n5520), .ZN(n7411)
         );
  NAND2_X1 U6640 ( .A1(n5463), .A2(P1_IR_REG_30__SCAN_IN), .ZN(n4852) );
  XNOR2_X2 U6641 ( .A(n5466), .B(n10047), .ZN(n5465) );
  NAND2_X2 U6642 ( .A1(n10045), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5475) );
  NAND2_X2 U6643 ( .A1(n5475), .A2(n5464), .ZN(n5466) );
  NAND2_X1 U6644 ( .A1(n6076), .A2(n6075), .ZN(n4857) );
  NAND2_X1 U6645 ( .A1(n4858), .A2(n6076), .ZN(n9457) );
  INV_X1 U6646 ( .A(n4857), .ZN(n9424) );
  INV_X1 U6647 ( .A(n9321), .ZN(n9420) );
  NAND2_X2 U6648 ( .A1(n9794), .A2(n6084), .ZN(n9765) );
  NAND2_X2 U6649 ( .A1(n9790), .A2(n6082), .ZN(n9794) );
  NAND2_X1 U6650 ( .A1(n7365), .A2(n4508), .ZN(n4863) );
  INV_X1 U6651 ( .A(n6073), .ZN(n9309) );
  NAND2_X1 U6652 ( .A1(n6161), .A2(n9918), .ZN(n4868) );
  INV_X1 U6653 ( .A(n6160), .ZN(n4869) );
  NOR2_X2 U6654 ( .A1(n9895), .A2(n4872), .ZN(n4871) );
  AND3_X2 U6655 ( .A1(n4874), .A2(n5426), .A3(P2_REG1_REG_9__SCAN_IN), .ZN(
        n8625) );
  INV_X1 U6656 ( .A(n5425), .ZN(n4873) );
  NOR2_X1 U6657 ( .A1(n8625), .A2(n4875), .ZN(n7545) );
  INV_X1 U6658 ( .A(n5436), .ZN(n5435) );
  NAND2_X1 U6659 ( .A1(n8703), .A2(n8704), .ZN(n8702) );
  NAND2_X1 U6660 ( .A1(n8685), .A2(n5434), .ZN(n8703) );
  NOR2_X1 U6661 ( .A1(n4881), .A2(n4878), .ZN(n5420) );
  INV_X1 U6662 ( .A(n4882), .ZN(n4878) );
  NAND2_X1 U6663 ( .A1(n4480), .A2(n7152), .ZN(n4882) );
  NAND3_X1 U6664 ( .A1(n4480), .A2(n7152), .A3(n6930), .ZN(n4879) );
  NAND2_X1 U6665 ( .A1(n4881), .A2(n6930), .ZN(n4880) );
  NAND2_X1 U6666 ( .A1(n4882), .A2(n4883), .ZN(n7220) );
  INV_X1 U6667 ( .A(n7217), .ZN(n4884) );
  NAND2_X1 U6668 ( .A1(n5439), .A2(n4886), .ZN(n4885) );
  OAI211_X1 U6669 ( .C1(n5439), .C2(n4887), .A(n5444), .B(n4885), .ZN(n5445)
         );
  NAND2_X1 U6670 ( .A1(n5439), .A2(n8741), .ZN(n8746) );
  NAND3_X1 U6671 ( .A1(n4896), .A2(n5429), .A3(n4895), .ZN(n4893) );
  INV_X1 U6672 ( .A(n5428), .ZN(n4897) );
  NAND2_X1 U6673 ( .A1(n4900), .A2(n4899), .ZN(n4898) );
  NAND2_X1 U6674 ( .A1(n5423), .A2(n6253), .ZN(n4901) );
  NAND2_X1 U6675 ( .A1(n4900), .A2(n4901), .ZN(n7386) );
  INV_X1 U6676 ( .A(n6912), .ZN(n4900) );
  NAND3_X1 U6677 ( .A1(n4903), .A2(n4902), .A3(P2_REG2_REG_1__SCAN_IN), .ZN(
        n6999) );
  NAND2_X1 U6678 ( .A1(n6999), .A2(n4903), .ZN(n6986) );
  NAND2_X1 U6679 ( .A1(n5307), .A2(n6180), .ZN(n4902) );
  INV_X1 U6680 ( .A(n8674), .ZN(n4904) );
  NAND2_X1 U6681 ( .A1(n4904), .A2(n4910), .ZN(n4909) );
  NAND3_X1 U6682 ( .A1(n8674), .A2(n4912), .A3(n8695), .ZN(n4905) );
  INV_X1 U6683 ( .A(n7017), .ZN(n4918) );
  NAND3_X1 U6684 ( .A1(n5323), .A2(n7017), .A3(P2_REG2_REG_5__SCAN_IN), .ZN(
        n7181) );
  NAND2_X1 U6685 ( .A1(n6985), .A2(n5309), .ZN(n4921) );
  XNOR2_X1 U6686 ( .A(n5334), .B(n4923), .ZN(n7541) );
  NAND2_X1 U6687 ( .A1(n4924), .A2(n6918), .ZN(n4926) );
  NAND2_X1 U6688 ( .A1(n4926), .A2(n4925), .ZN(n6920) );
  NAND2_X1 U6689 ( .A1(n8748), .A2(n8747), .ZN(n4931) );
  NAND3_X1 U6690 ( .A1(n4932), .A2(n5355), .A3(n4931), .ZN(n5358) );
  NAND2_X1 U6691 ( .A1(n5350), .A2(n5351), .ZN(n8725) );
  NAND2_X1 U6692 ( .A1(n5413), .A2(n5414), .ZN(n6996) );
  AOI21_X2 U6693 ( .B1(n9866), .B2(n9883), .A(n9475), .ZN(n8221) );
  OAI21_X2 U6694 ( .B1(n8625), .B2(n8624), .A(n8623), .ZN(n8622) );
  NAND2_X1 U6695 ( .A1(n8234), .A2(n9351), .ZN(n9866) );
  NAND2_X1 U6696 ( .A1(n5040), .A2(n5205), .ZN(P1_U3551) );
  NAND3_X1 U6697 ( .A1(n5481), .A2(n5523), .A3(n5539), .ZN(n4935) );
  NAND2_X1 U6698 ( .A1(n5483), .A2(n5539), .ZN(n4936) );
  INV_X1 U6699 ( .A(n5667), .ZN(n4946) );
  NAND2_X1 U6700 ( .A1(n5632), .A2(n5631), .ZN(n5653) );
  NAND2_X1 U6701 ( .A1(n4949), .A2(n5651), .ZN(n5668) );
  OAI21_X2 U6702 ( .B1(n5759), .B2(n4956), .A(n4953), .ZN(n5820) );
  NAND3_X2 U6703 ( .A1(n5476), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4968) );
  NAND3_X1 U6704 ( .A1(n4969), .A2(n4968), .A3(n4967), .ZN(n4966) );
  NAND2_X1 U6705 ( .A1(n5863), .A2(n4475), .ZN(n4972) );
  NAND2_X1 U6706 ( .A1(n5863), .A2(n4982), .ZN(n4979) );
  NAND2_X1 U6707 ( .A1(n4979), .A2(n4980), .ZN(n5901) );
  INV_X1 U6708 ( .A(n6101), .ZN(n9849) );
  NAND2_X1 U6709 ( .A1(n6103), .A2(n8245), .ZN(n6147) );
  XNOR2_X1 U6710 ( .A(n9681), .B(n8154), .ZN(n8155) );
  NAND3_X1 U6711 ( .A1(n4997), .A2(n7762), .A3(n6098), .ZN(n7612) );
  NAND2_X1 U6712 ( .A1(n5006), .A2(n5004), .ZN(n7861) );
  NAND2_X1 U6713 ( .A1(n7705), .A2(n5007), .ZN(n5006) );
  INV_X1 U6714 ( .A(n5818), .ZN(n5020) );
  OR2_X1 U6715 ( .A1(n9889), .A2(n5775), .ZN(n5021) );
  NAND2_X1 U6716 ( .A1(n5818), .A2(n5015), .ZN(n5014) );
  NAND2_X1 U6717 ( .A1(n9731), .A2(n5025), .ZN(n5022) );
  NAND2_X1 U6718 ( .A1(n5022), .A2(n5023), .ZN(n9699) );
  NAND2_X1 U6719 ( .A1(n9731), .A2(n6003), .ZN(n5024) );
  AOI21_X1 U6720 ( .B1(n7615), .B2(n5031), .A(n4511), .ZN(n5029) );
  NAND2_X1 U6721 ( .A1(n5041), .A2(n10161), .ZN(n5040) );
  NAND3_X1 U6722 ( .A1(n7430), .A2(n6231), .A3(n8415), .ZN(n5045) );
  NAND2_X1 U6723 ( .A1(n5046), .A2(n8415), .ZN(n10166) );
  NAND2_X1 U6724 ( .A1(n7431), .A2(n10163), .ZN(n5046) );
  NAND2_X1 U6725 ( .A1(n8180), .A2(n5058), .ZN(n5054) );
  OAI21_X1 U6726 ( .B1(n8180), .B2(n5059), .A(n8569), .ZN(n8780) );
  NAND2_X1 U6727 ( .A1(n5054), .A2(n5055), .ZN(n6500) );
  NAND2_X1 U6728 ( .A1(n5062), .A2(n5060), .ZN(n6466) );
  NAND2_X1 U6730 ( .A1(n6504), .A2(n10171), .ZN(n5067) );
  INV_X1 U6731 ( .A(n6553), .ZN(n5066) );
  AND2_X1 U6732 ( .A1(n5067), .A2(n6553), .ZN(n8072) );
  NAND2_X1 U6733 ( .A1(n8173), .A2(n6431), .ZN(n5069) );
  NAND3_X2 U6734 ( .A1(n10405), .A2(n5071), .A3(n5070), .ZN(n5713) );
  NAND2_X1 U6735 ( .A1(n9139), .A2(n5082), .ZN(n5080) );
  INV_X1 U6736 ( .A(n5802), .ZN(n5087) );
  NAND2_X1 U6737 ( .A1(n5096), .A2(n5092), .ZN(n5097) );
  NOR3_X1 U6738 ( .A1(n5095), .A2(n9208), .A3(n4462), .ZN(n5092) );
  CLKBUF_X1 U6739 ( .A(n5096), .Z(n5093) );
  NAND2_X1 U6740 ( .A1(n5097), .A2(n9207), .ZN(n9132) );
  NAND2_X1 U6741 ( .A1(n5098), .A2(n5100), .ZN(n6516) );
  NAND2_X1 U6742 ( .A1(n6515), .A2(n4516), .ZN(n5098) );
  NAND2_X1 U6743 ( .A1(n7427), .A2(n5103), .ZN(n5104) );
  NAND2_X1 U6744 ( .A1(n6524), .A2(n5112), .ZN(n5108) );
  NAND2_X1 U6745 ( .A1(n5120), .A2(n5119), .ZN(n8888) );
  NAND2_X1 U6746 ( .A1(n6514), .A2(n5122), .ZN(n5121) );
  NAND2_X1 U6747 ( .A1(n6511), .A2(n5139), .ZN(n5138) );
  NAND2_X1 U6748 ( .A1(n6511), .A2(n8491), .ZN(n7464) );
  NAND2_X1 U6749 ( .A1(n5283), .A2(n5142), .ZN(n9075) );
  NAND3_X1 U6750 ( .A1(n5147), .A2(n7143), .A3(n5146), .ZN(n7234) );
  NAND2_X1 U6751 ( .A1(n5150), .A2(n5148), .ZN(n7418) );
  NAND2_X1 U6752 ( .A1(n7308), .A2(n7343), .ZN(n5150) );
  NAND3_X1 U6753 ( .A1(n7262), .A2(n7260), .A3(n7261), .ZN(n7300) );
  INV_X1 U6754 ( .A(n8341), .ZN(n5154) );
  OAI21_X1 U6755 ( .B1(n8341), .B2(n5159), .A(n5157), .ZN(n8262) );
  OAI21_X1 U6756 ( .B1(n8341), .B2(n5165), .A(n5163), .ZN(n5162) );
  AND2_X1 U6757 ( .A1(n8088), .A2(n8854), .ZN(n5167) );
  NAND2_X1 U6758 ( .A1(n7548), .A2(n4446), .ZN(n7587) );
  OR2_X1 U6759 ( .A1(n8097), .A2(n5174), .ZN(n5170) );
  NAND2_X1 U6760 ( .A1(n5170), .A2(n5171), .ZN(n8103) );
  NAND2_X1 U6761 ( .A1(n8097), .A2(n8381), .ZN(n8384) );
  NAND3_X1 U6762 ( .A1(n7589), .A2(n7588), .A3(n4459), .ZN(n5176) );
  NAND3_X1 U6763 ( .A1(n5176), .A2(n5181), .A3(n5177), .ZN(n7899) );
  INV_X1 U6764 ( .A(n7898), .ZN(n5182) );
  CLKBUF_X1 U6765 ( .A(n5289), .Z(n5184) );
  NAND2_X1 U6766 ( .A1(n8079), .A2(n5188), .ZN(n5187) );
  NAND2_X1 U6767 ( .A1(n8079), .A2(n5198), .ZN(n5197) );
  NAND2_X1 U6768 ( .A1(n5187), .A2(n5191), .ZN(n8273) );
  OR2_X1 U6769 ( .A1(n8080), .A2(n8081), .ZN(n5204) );
  NAND4_X4 U6770 ( .A1(n5515), .A2(n5514), .A3(n5513), .A4(n5512), .ZN(n7808)
         );
  NAND2_X1 U6771 ( .A1(n8129), .A2(n7954), .ZN(n7447) );
  NAND2_X1 U6772 ( .A1(n6038), .A2(n6037), .ZN(n6040) );
  INV_X1 U6773 ( .A(n5622), .ZN(n5619) );
  NAND2_X1 U6774 ( .A1(n8224), .A2(n6100), .ZN(n6101) );
  INV_X1 U6775 ( .A(n6873), .ZN(n8245) );
  INV_X1 U6776 ( .A(n7452), .ZN(n5511) );
  AOI21_X2 U6777 ( .B1(n6151), .B2(n6150), .A(n6149), .ZN(n6162) );
  INV_X1 U6778 ( .A(n7445), .ZN(n6098) );
  INV_X1 U6781 ( .A(n6648), .ZN(n6651) );
  NAND2_X1 U6782 ( .A1(n6369), .A2(n6368), .ZN(n8878) );
  INV_X1 U6783 ( .A(n6057), .ZN(n5677) );
  OR2_X4 U6784 ( .A1(n6599), .A2(n6611), .ZN(n6832) );
  INV_X1 U6785 ( .A(n6175), .ZN(n8110) );
  AND2_X1 U6786 ( .A1(n5215), .A2(n6164), .ZN(n5205) );
  AND2_X1 U6787 ( .A1(n6563), .A2(n6953), .ZN(n5206) );
  OR2_X1 U6788 ( .A1(n6274), .A2(n5424), .ZN(n5207) );
  INV_X1 U6789 ( .A(n9971), .ZN(n6102) );
  AND2_X1 U6790 ( .A1(n8422), .A2(n5211), .ZN(n5209) );
  AND2_X1 U6791 ( .A1(n4432), .A2(n7197), .ZN(n5210) );
  OR2_X1 U6792 ( .A1(n10224), .A2(n7851), .ZN(n5211) );
  AND2_X1 U6793 ( .A1(n8167), .A2(n8614), .ZN(n5212) );
  OR2_X1 U6794 ( .A1(n6508), .A2(n7360), .ZN(n5213) );
  AND2_X1 U6795 ( .A1(n8436), .A2(n6530), .ZN(n5214) );
  OR2_X1 U6796 ( .A1(n9691), .A2(n9948), .ZN(n5215) );
  OR2_X1 U6797 ( .A1(n8076), .A2(n8974), .ZN(n5216) );
  AND2_X1 U6798 ( .A1(n9117), .A2(n9116), .ZN(n5217) );
  OR2_X1 U6799 ( .A1(P2_REG0_REG_29__SCAN_IN), .A2(n10230), .ZN(n5218) );
  OR2_X1 U6800 ( .A1(n8076), .A2(n9045), .ZN(n5219) );
  OR2_X1 U6801 ( .A1(n9691), .A2(n10026), .ZN(n5220) );
  AND2_X1 U6802 ( .A1(n5456), .A2(n10272), .ZN(n5222) );
  OR2_X1 U6803 ( .A1(n8329), .A2(n8801), .ZN(n5223) );
  INV_X1 U6804 ( .A(n8768), .ZN(n5444) );
  INV_X1 U6805 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6172) );
  INV_X1 U6806 ( .A(n9754), .ZN(n5979) );
  NOR2_X1 U6807 ( .A1(n5984), .A2(n5983), .ZN(n5224) );
  NOR2_X1 U6808 ( .A1(n5982), .A2(n5984), .ZN(n5225) );
  INV_X1 U6809 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5565) );
  AND2_X1 U6810 ( .A1(n7486), .A2(n7485), .ZN(n5226) );
  INV_X1 U6811 ( .A(n9988), .ZN(n6100) );
  AND2_X1 U6812 ( .A1(n6557), .A2(n6555), .ZN(n5227) );
  NAND2_X1 U6813 ( .A1(n6537), .A2(n6536), .ZN(n5228) );
  OR3_X1 U6814 ( .A1(n9689), .A2(n10143), .A3(n9687), .ZN(n5229) );
  AND2_X1 U6815 ( .A1(n8583), .A2(n6530), .ZN(n5230) );
  AND2_X1 U6816 ( .A1(n8993), .A2(n6530), .ZN(n5231) );
  OR2_X1 U6817 ( .A1(n9679), .A2(n9435), .ZN(n5232) );
  AND2_X1 U6818 ( .A1(n9687), .A2(n10136), .ZN(n5233) );
  NAND2_X1 U6819 ( .A1(n6873), .A2(n7727), .ZN(n5234) );
  NAND2_X1 U6820 ( .A1(n7951), .A2(n10132), .ZN(n7445) );
  OR2_X1 U6821 ( .A1(n8988), .A2(n8613), .ZN(n5235) );
  AND2_X1 U6822 ( .A1(n8535), .A2(n8846), .ZN(n8536) );
  INV_X1 U6823 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5448) );
  INV_X1 U6824 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10400) );
  AND2_X1 U6825 ( .A1(n5417), .A2(n7159), .ZN(n5418) );
  INV_X1 U6826 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5282) );
  INV_X1 U6827 ( .A(n5579), .ZN(n5577) );
  NOR2_X1 U6828 ( .A1(n8151), .A2(n6950), .ZN(n5592) );
  INV_X1 U6829 ( .A(SI_11_), .ZN(n10559) );
  OR2_X1 U6830 ( .A1(n8571), .A2(n8793), .ZN(n6529) );
  INV_X1 U6831 ( .A(n5918), .ZN(n5919) );
  NAND2_X1 U6832 ( .A1(n8098), .A2(n8257), .ZN(n8099) );
  INV_X1 U6833 ( .A(n7265), .ZN(n7262) );
  NAND2_X1 U6834 ( .A1(n5337), .A2(n7881), .ZN(n5338) );
  INV_X1 U6835 ( .A(n6549), .ZN(n6550) );
  INV_X1 U6836 ( .A(n6877), .ZN(n6883) );
  AND2_X1 U6837 ( .A1(n6601), .A2(n6837), .ZN(n6598) );
  INV_X1 U6838 ( .A(n7376), .ZN(n6617) );
  NAND2_X1 U6839 ( .A1(n5547), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5579) );
  INV_X1 U6840 ( .A(n9679), .ZN(n8154) );
  AND2_X1 U6841 ( .A1(n9689), .A2(n5233), .ZN(n6146) );
  NAND2_X1 U6842 ( .A1(n5594), .A2(n5593), .ZN(n5595) );
  AND2_X1 U6843 ( .A1(n5961), .A2(n5960), .ZN(n5983) );
  INV_X1 U6844 ( .A(n8612), .ZN(n8363) );
  INV_X1 U6845 ( .A(n8371), .ZN(n8390) );
  INV_X1 U6846 ( .A(n8967), .ZN(n8874) );
  INV_X1 U6847 ( .A(n8607), .ZN(n8182) );
  INV_X1 U6848 ( .A(n10167), .ZN(n8883) );
  INV_X1 U6849 ( .A(n10171), .ZN(n10185) );
  INV_X1 U6850 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U6851 ( .A1(n6685), .A2(n6684), .ZN(n9240) );
  INV_X1 U6852 ( .A(n9750), .ZN(n9717) );
  INV_X1 U6853 ( .A(n9267), .ZN(n9282) );
  INV_X1 U6854 ( .A(n9966), .ZN(n9815) );
  OR2_X1 U6855 ( .A1(n10040), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6135) );
  INV_X1 U6856 ( .A(n9916), .ZN(n9251) );
  NOR2_X2 U6857 ( .A1(n4450), .A2(n4572), .ZN(n7707) );
  INV_X1 U6858 ( .A(n9976), .ZN(n9907) );
  INV_X1 U6859 ( .A(n9918), .ZN(n9893) );
  XNOR2_X1 U6860 ( .A(n5703), .B(SI_11_), .ZN(n5706) );
  XNOR2_X1 U6861 ( .A(n5648), .B(SI_8_), .ZN(n5652) );
  AND2_X1 U6862 ( .A1(n7128), .A2(n7127), .ZN(n8371) );
  AND2_X1 U6863 ( .A1(n7976), .A2(n6499), .ZN(n8606) );
  AND3_X1 U6864 ( .A1(n6356), .A2(n6355), .A3(n6354), .ZN(n8313) );
  INV_X1 U6865 ( .A(n8587), .ZN(n8596) );
  AND2_X1 U6866 ( .A1(n8546), .A2(n8810), .ZN(n8552) );
  INV_X1 U6867 ( .A(n8974), .ZN(n8983) );
  AND2_X1 U6868 ( .A1(n6584), .A2(n6583), .ZN(n6585) );
  AND2_X1 U6869 ( .A1(n7171), .A2(n7841), .ZN(n10198) );
  AND2_X1 U6870 ( .A1(n7130), .A2(n7841), .ZN(n10189) );
  OR2_X1 U6871 ( .A1(n6951), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6565) );
  INV_X1 U6872 ( .A(n9279), .ZN(n9247) );
  INV_X1 U6873 ( .A(n9287), .ZN(n9236) );
  INV_X1 U6874 ( .A(n9250), .ZN(n9284) );
  AND2_X1 U6875 ( .A1(n5978), .A2(n5977), .ZN(n9771) );
  OR2_X1 U6876 ( .A1(n7118), .A2(n7034), .ZN(n10067) );
  INV_X1 U6877 ( .A(n10088), .ZN(n9650) );
  AND2_X1 U6878 ( .A1(n9478), .A2(n9480), .ZN(n9428) );
  INV_X1 U6879 ( .A(n9876), .ZN(n10108) );
  AND2_X1 U6880 ( .A1(n7028), .A2(n4437), .ZN(n9913) );
  OAI21_X1 U6881 ( .B1(n8245), .B2(n10026), .A(n6167), .ZN(n6168) );
  AND2_X1 U6882 ( .A1(n7814), .A2(n10151), .ZN(n10143) );
  INV_X1 U6883 ( .A(n10143), .ZN(n10136) );
  AND2_X1 U6884 ( .A1(n7843), .A2(n7674), .ZN(n7337) );
  NAND2_X1 U6885 ( .A1(n7029), .A2(n6850), .ZN(n10269) );
  INV_X1 U6886 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10414) );
  NOR2_X1 U6887 ( .A1(n10588), .A2(n10587), .ZN(n8021) );
  NOR2_X1 U6888 ( .A1(n10586), .A2(n10585), .ZN(n8027) );
  NOR2_X1 U6889 ( .A1(n10263), .A2(n10262), .ZN(n8033) );
  OR3_X1 U6890 ( .A1(n7093), .A2(n7092), .A3(n9073), .ZN(n8378) );
  INV_X1 U6891 ( .A(n8388), .ZN(n8336) );
  INV_X1 U6892 ( .A(n8826), .ZN(n8609) );
  INV_X1 U6893 ( .A(n8081), .ZN(n8926) );
  OR2_X1 U6894 ( .A1(n7097), .A2(n5273), .ZN(n8756) );
  OR2_X1 U6895 ( .A1(n8756), .A2(n8589), .ZN(n8760) );
  OR2_X1 U6896 ( .A1(n6967), .A2(n6539), .ZN(n8768) );
  INV_X1 U6897 ( .A(n10181), .ZN(n10183) );
  NAND2_X2 U6898 ( .A1(n7079), .A2(n8885), .ZN(n10181) );
  NAND2_X1 U6899 ( .A1(n10245), .A2(n10189), .ZN(n8974) );
  OR2_X1 U6900 ( .A1(n10229), .A2(n10225), .ZN(n9070) );
  AND2_X1 U6901 ( .A1(n6888), .A2(n6887), .ZN(n10229) );
  INV_X2 U6902 ( .A(n10229), .ZN(n10230) );
  INV_X1 U6903 ( .A(n6961), .ZN(n6962) );
  AND2_X1 U6904 ( .A1(n6565), .A2(n6564), .ZN(n9074) );
  INV_X1 U6905 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n10474) );
  INV_X1 U6906 ( .A(n6253), .ZN(n7385) );
  INV_X1 U6907 ( .A(n10098), .ZN(n9671) );
  NAND2_X1 U6908 ( .A1(n6866), .A2(n6851), .ZN(n9262) );
  INV_X1 U6909 ( .A(n9223), .ZN(n9287) );
  INV_X1 U6910 ( .A(n9736), .ZN(n9548) );
  OR2_X1 U6911 ( .A1(n7118), .A2(n9535), .ZN(n10090) );
  AND2_X2 U6912 ( .A1(n7741), .A2(n9922), .ZN(n10112) );
  AND2_X2 U6913 ( .A1(n6166), .A2(n7732), .ZN(n10161) );
  AOI21_X1 U6914 ( .B1(n6169), .B2(n10155), .A(n6168), .ZN(n6170) );
  INV_X1 U6915 ( .A(n10122), .ZN(n10270) );
  OR2_X1 U6916 ( .A1(n10269), .A2(n10041), .ZN(n10122) );
  OR2_X1 U6917 ( .A1(n7029), .A2(P1_U3086), .ZN(n9538) );
  INV_X1 U6918 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7482) );
  INV_X1 U6919 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10442) );
  NOR2_X1 U6920 ( .A1(n8020), .A2(n8019), .ZN(n10588) );
  NOR2_X1 U6921 ( .A1(n8032), .A2(n8031), .ZN(n10263) );
  INV_X1 U6922 ( .A(n8756), .ZN(P2_U3893) );
  INV_X1 U6923 ( .A(n6170), .ZN(P1_U3518) );
  NAND4_X1 U6924 ( .A1(n5238), .A2(n5237), .A3(n5236), .A4(n5335), .ZN(n5259)
         );
  NOR2_X2 U6925 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5294) );
  NOR2_X1 U6926 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5240) );
  NOR2_X1 U6927 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5239) );
  NAND3_X1 U6928 ( .A1(n5294), .A2(n5240), .A3(n5239), .ZN(n5260) );
  INV_X1 U6929 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5244) );
  NAND2_X1 U6930 ( .A1(n5274), .A2(n5245), .ZN(n5278) );
  INV_X1 U6931 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5247) );
  INV_X1 U6932 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5246) );
  AOI21_X1 U6933 ( .B1(n5270), .B2(n5247), .A(n5246), .ZN(n5252) );
  INV_X1 U6934 ( .A(n5252), .ZN(n5249) );
  INV_X1 U6935 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U6936 ( .A1(n5249), .A2(n5248), .ZN(n5254) );
  INV_X1 U6937 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5250) );
  INV_X1 U6938 ( .A(n6560), .ZN(n5269) );
  NAND2_X1 U6939 ( .A1(n5252), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n5253) );
  NOR2_X1 U6940 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5258) );
  NAND4_X1 U6941 ( .A1(n5258), .A2(n5257), .A3(n5256), .A4(n5255), .ZN(n5263)
         );
  INV_X1 U6942 ( .A(n5263), .ZN(n5264) );
  NAND3_X1 U6943 ( .A1(n4500), .A2(n5184), .A3(n5264), .ZN(n5265) );
  NAND2_X1 U6944 ( .A1(n5265), .A2(n5352), .ZN(n5266) );
  MUX2_X1 U6945 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5266), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5267) );
  NOR2_X1 U6946 ( .A1(n6559), .A2(n8068), .ZN(n5268) );
  NAND2_X1 U6947 ( .A1(n5269), .A2(n5268), .ZN(n7097) );
  INV_X1 U6948 ( .A(n5270), .ZN(n5271) );
  NAND2_X1 U6949 ( .A1(n5271), .A2(n5352), .ZN(n5272) );
  XNOR2_X1 U6950 ( .A(n5272), .B(n5247), .ZN(n7096) );
  INV_X1 U6951 ( .A(n6576), .ZN(n5273) );
  NAND2_X1 U6952 ( .A1(n5357), .A2(n5356), .ZN(n5275) );
  NAND2_X1 U6953 ( .A1(n6502), .A2(n6501), .ZN(n5276) );
  XNOR2_X2 U6954 ( .A(n5277), .B(n5244), .ZN(n7130) );
  NAND2_X1 U6955 ( .A1(n5278), .A2(n5352), .ZN(n5279) );
  NAND2_X2 U6956 ( .A1(n6530), .A2(n8592), .ZN(n8570) );
  NAND2_X1 U6957 ( .A1(n7097), .A2(n8570), .ZN(n5280) );
  NAND2_X1 U6958 ( .A1(n5280), .A2(n7096), .ZN(n5361) );
  XNOR2_X2 U6959 ( .A(n5285), .B(n5284), .ZN(n5409) );
  XNOR2_X1 U6960 ( .A(n5286), .B(n5282), .ZN(n5359) );
  NAND2_X2 U6961 ( .A1(n5409), .A2(n5359), .ZN(n6547) );
  NAND2_X1 U6962 ( .A1(n5361), .A2(n6547), .ZN(n5287) );
  NAND2_X1 U6963 ( .A1(n5287), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U6964 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8909) );
  NAND2_X1 U6965 ( .A1(n5289), .A2(n5288), .ZN(n5324) );
  INV_X1 U6966 ( .A(n5327), .ZN(n5291) );
  INV_X1 U6967 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U6968 ( .A1(n5291), .A2(n5290), .ZN(n5330) );
  INV_X1 U6969 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5301) );
  INV_X1 U6970 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n10298) );
  INV_X1 U6971 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5292) );
  NAND4_X1 U6972 ( .A1(n5335), .A2(n5301), .A3(n10298), .A4(n5292), .ZN(n5293)
         );
  OAI21_X1 U6973 ( .B1(n5339), .B2(P2_IR_REG_13__SCAN_IN), .A(n5352), .ZN(
        n5344) );
  INV_X1 U6974 ( .A(n5294), .ZN(n5295) );
  NAND2_X1 U6975 ( .A1(n5295), .A2(n5352), .ZN(n5296) );
  NAND2_X1 U6976 ( .A1(n5344), .A2(n5296), .ZN(n5347) );
  INV_X1 U6977 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5297) );
  XNOR2_X1 U6978 ( .A(n5347), .B(n5297), .ZN(n8717) );
  INV_X1 U6979 ( .A(n8671), .ZN(n7124) );
  NAND2_X1 U6980 ( .A1(n5298), .A2(n5352), .ZN(n5333) );
  OAI21_X1 U6981 ( .B1(P2_IR_REG_9__SCAN_IN), .B2(P2_IR_REG_10__SCAN_IN), .A(
        n5352), .ZN(n5299) );
  NAND2_X1 U6982 ( .A1(n5333), .A2(n5299), .ZN(n5336) );
  OAI21_X1 U6983 ( .B1(n5336), .B2(P2_IR_REG_11__SCAN_IN), .A(n5352), .ZN(
        n5300) );
  XNOR2_X1 U6984 ( .A(n5300), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6310) );
  INV_X1 U6985 ( .A(n6310), .ZN(n6978) );
  NAND2_X1 U6986 ( .A1(n5333), .A2(n5301), .ZN(n5302) );
  NAND2_X1 U6987 ( .A1(n5302), .A2(n5352), .ZN(n5303) );
  INV_X1 U6988 ( .A(n8637), .ZN(n6957) );
  INV_X1 U6989 ( .A(n5308), .ZN(n5304) );
  INV_X2 U6990 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5310) );
  XNOR2_X1 U6991 ( .A(n5305), .B(n5310), .ZN(n5416) );
  INV_X1 U6992 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10558) );
  XNOR2_X1 U6993 ( .A(n5416), .B(n10558), .ZN(n6987) );
  NAND2_X1 U6994 ( .A1(n4436), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5307) );
  INV_X1 U6995 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7249) );
  NAND2_X1 U6996 ( .A1(n6987), .A2(n6986), .ZN(n6985) );
  NAND2_X1 U6997 ( .A1(n6994), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U6998 ( .A1(n5412), .A2(n5310), .ZN(n5312) );
  NAND2_X1 U6999 ( .A1(n5312), .A2(n5352), .ZN(n5311) );
  NAND2_X1 U7000 ( .A1(n7212), .A2(n7210), .ZN(n5315) );
  OAI21_X1 U7001 ( .B1(n5312), .B2(P2_IR_REG_3__SCAN_IN), .A(n5352), .ZN(n5313) );
  MUX2_X1 U7002 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5313), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5314) );
  AND2_X1 U7003 ( .A1(n5314), .A2(n5317), .ZN(n6219) );
  XNOR2_X1 U7004 ( .A(n6219), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n7209) );
  INV_X1 U7005 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6226) );
  OR2_X1 U7006 ( .A1(n6219), .A2(n6226), .ZN(n5316) );
  NAND2_X1 U7007 ( .A1(n7214), .A2(n5316), .ZN(n5322) );
  INV_X1 U7008 ( .A(n5322), .ZN(n5321) );
  NAND2_X1 U7009 ( .A1(n5317), .A2(n5352), .ZN(n5318) );
  MUX2_X1 U7010 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5318), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5319) );
  NAND2_X1 U7011 ( .A1(n5319), .A2(n5324), .ZN(n6930) );
  INV_X1 U7012 ( .A(n6930), .ZN(n5320) );
  NAND2_X1 U7013 ( .A1(n5321), .A2(n5320), .ZN(n5323) );
  NAND2_X1 U7014 ( .A1(n5324), .A2(n5352), .ZN(n5325) );
  INV_X1 U7015 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7458) );
  OR2_X1 U7016 ( .A1(n6242), .A2(n7458), .ZN(n5326) );
  NAND2_X1 U7017 ( .A1(n5327), .A2(n5352), .ZN(n5328) );
  XNOR2_X1 U7018 ( .A(n5328), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7019 ( .A1(n5330), .A2(n5352), .ZN(n5331) );
  XNOR2_X1 U7020 ( .A(n5331), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6274) );
  INV_X1 U7021 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7602) );
  OR2_X1 U7022 ( .A1(n6274), .A2(n7602), .ZN(n5332) );
  XNOR2_X1 U7023 ( .A(n5333), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7540) );
  NAND2_X1 U7024 ( .A1(n7541), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8640) );
  INV_X1 U7025 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8164) );
  XNOR2_X1 U7026 ( .A(n8637), .B(n8164), .ZN(n8639) );
  AOI21_X1 U7027 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n6957), .A(n8642), .ZN(
        n5337) );
  XNOR2_X1 U7028 ( .A(n5336), .B(n5335), .ZN(n7881) );
  INV_X1 U7029 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7803) );
  XNOR2_X1 U7030 ( .A(n6310), .B(n7803), .ZN(n6896) );
  NAND2_X1 U7031 ( .A1(n5339), .A2(n5352), .ZN(n5340) );
  XNOR2_X1 U7032 ( .A(n5340), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8656) );
  NOR2_X1 U7033 ( .A1(n5341), .A2(n8656), .ZN(n5342) );
  NAND2_X1 U7034 ( .A1(n8657), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8674) );
  INV_X1 U7035 ( .A(n5342), .ZN(n8672) );
  INV_X1 U7036 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n10356) );
  XNOR2_X1 U7037 ( .A(n8671), .B(n10356), .ZN(n8673) );
  INV_X1 U7038 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U7039 ( .A1(n5344), .A2(n5343), .ZN(n5345) );
  NAND2_X1 U7040 ( .A1(n5345), .A2(n5352), .ZN(n5346) );
  XNOR2_X1 U7041 ( .A(n5346), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8695) );
  NAND2_X1 U7042 ( .A1(n8696), .A2(n4481), .ZN(n8711) );
  XNOR2_X1 U7043 ( .A(n8717), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n8712) );
  NAND2_X1 U7044 ( .A1(n8711), .A2(n8712), .ZN(n8710) );
  OAI21_X1 U7045 ( .B1(n5347), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5348) );
  XNOR2_X1 U7046 ( .A(n5348), .B(P2_IR_REG_17__SCAN_IN), .ZN(n6357) );
  INV_X1 U7047 ( .A(n6357), .ZN(n8731) );
  INV_X1 U7048 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n10471) );
  INV_X1 U7049 ( .A(n5351), .ZN(n8748) );
  NAND2_X1 U7050 ( .A1(n4524), .A2(n5352), .ZN(n5353) );
  XNOR2_X1 U7051 ( .A(n5353), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8765) );
  INV_X1 U7052 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8887) );
  OR2_X1 U7053 ( .A1(n8765), .A2(n8887), .ZN(n5355) );
  NAND2_X1 U7054 ( .A1(n8765), .A2(n8887), .ZN(n5354) );
  AND2_X1 U7055 ( .A1(n5355), .A2(n5354), .ZN(n8747) );
  XNOR2_X1 U7056 ( .A(n5357), .B(n5356), .ZN(n8587) );
  XNOR2_X1 U7057 ( .A(n8596), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n5364) );
  XNOR2_X1 U7058 ( .A(n5358), .B(n5364), .ZN(n5360) );
  NOR2_X1 U7059 ( .A1(n5409), .A2(P2_U3151), .ZN(n9083) );
  AND2_X1 U7060 ( .A1(n5361), .A2(n9083), .ZN(n5443) );
  NAND2_X1 U7061 ( .A1(n5360), .A2(n8750), .ZN(n5446) );
  NOR2_X1 U7062 ( .A1(n5404), .A2(P2_U3151), .ZN(n9087) );
  AND2_X1 U7063 ( .A1(n5361), .A2(n9087), .ZN(n5362) );
  MUX2_X1 U7064 ( .A(P2_U3893), .B(n5362), .S(n5409), .Z(n8718) );
  INV_X1 U7065 ( .A(n7096), .ZN(n7935) );
  NOR2_X1 U7066 ( .A1(n7097), .A2(n7935), .ZN(n5363) );
  NAND2_X1 U7067 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8274) );
  OAI21_X1 U7068 ( .B1(n8759), .B2(n5477), .A(n8274), .ZN(n5410) );
  XNOR2_X1 U7069 ( .A(n8587), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n5441) );
  INV_X1 U7070 ( .A(n5364), .ZN(n5365) );
  MUX2_X1 U7071 ( .A(n5441), .B(n5365), .S(n6539), .Z(n5408) );
  MUX2_X1 U7072 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n5404), .Z(n5399) );
  INV_X1 U7073 ( .A(n5399), .ZN(n5400) );
  INV_X1 U7074 ( .A(n6219), .ZN(n7233) );
  XNOR2_X1 U7075 ( .A(n5367), .B(n6180), .ZN(n7003) );
  INV_X1 U7076 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6185) );
  INV_X1 U7077 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U7078 ( .A1(n5366), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7002) );
  INV_X1 U7079 ( .A(n6180), .ZN(n7009) );
  AOI22_X1 U7080 ( .A1(n7003), .A2(n7002), .B1(n5367), .B2(n7009), .ZN(n6979)
         );
  XNOR2_X1 U7081 ( .A(n5368), .B(n6994), .ZN(n6980) );
  INV_X1 U7082 ( .A(n6994), .ZN(n5370) );
  INV_X1 U7083 ( .A(n5368), .ZN(n5369) );
  OAI22_X1 U7084 ( .A1(n6979), .A2(n6980), .B1(n5370), .B2(n5369), .ZN(n7150)
         );
  XOR2_X1 U7085 ( .A(n7159), .B(n5371), .Z(n7151) );
  NOR2_X1 U7086 ( .A1(n7150), .A2(n7151), .ZN(n7228) );
  NOR2_X1 U7087 ( .A1(n5371), .A2(n6928), .ZN(n7227) );
  XNOR2_X1 U7088 ( .A(n5372), .B(n7233), .ZN(n7226) );
  NOR3_X1 U7089 ( .A1(n7228), .A2(n7227), .A3(n7226), .ZN(n7225) );
  AOI21_X1 U7090 ( .B1(n5372), .B2(n7233), .A(n7225), .ZN(n7178) );
  XNOR2_X1 U7091 ( .A(n5373), .B(n6930), .ZN(n7177) );
  INV_X1 U7092 ( .A(n5373), .ZN(n5374) );
  INV_X1 U7093 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10242) );
  NAND2_X1 U7094 ( .A1(n5375), .A2(n6242), .ZN(n5376) );
  OAI21_X1 U7095 ( .B1(n5375), .B2(n6242), .A(n5376), .ZN(n7010) );
  INV_X1 U7096 ( .A(n5376), .ZN(n7393) );
  INV_X1 U7097 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7563) );
  NAND2_X1 U7098 ( .A1(n5377), .A2(n6253), .ZN(n6916) );
  INV_X1 U7099 ( .A(n5377), .ZN(n5378) );
  NAND2_X1 U7100 ( .A1(n5378), .A2(n7385), .ZN(n5379) );
  AND2_X1 U7101 ( .A1(n6916), .A2(n5379), .ZN(n7392) );
  INV_X1 U7102 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5424) );
  MUX2_X1 U7103 ( .A(n7602), .B(n5424), .S(n5404), .Z(n5380) );
  NAND2_X1 U7104 ( .A1(n5380), .A2(n6274), .ZN(n5383) );
  INV_X1 U7105 ( .A(n5380), .ZN(n5381) );
  INV_X1 U7106 ( .A(n6274), .ZN(n6938) );
  NAND2_X1 U7107 ( .A1(n5381), .A2(n6938), .ZN(n5382) );
  NAND2_X1 U7108 ( .A1(n5383), .A2(n5382), .ZN(n6915) );
  INV_X1 U7109 ( .A(n5383), .ZN(n7535) );
  INV_X1 U7110 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7679) );
  INV_X1 U7111 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10500) );
  MUX2_X1 U7112 ( .A(n7679), .B(n10500), .S(n5404), .Z(n5384) );
  NAND2_X1 U7113 ( .A1(n7540), .A2(n5384), .ZN(n8631) );
  OR2_X1 U7114 ( .A1(n7540), .A2(n5384), .ZN(n5385) );
  AND2_X1 U7115 ( .A1(n8631), .A2(n5385), .ZN(n7534) );
  OAI21_X1 U7116 ( .B1(n7536), .B2(n7535), .A(n7534), .ZN(n8632) );
  INV_X1 U7117 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10545) );
  MUX2_X1 U7118 ( .A(n8164), .B(n10545), .S(n5404), .Z(n5386) );
  NAND2_X1 U7119 ( .A1(n8637), .A2(n5386), .ZN(n5388) );
  OR2_X1 U7120 ( .A1(n8637), .A2(n5386), .ZN(n5387) );
  NAND2_X1 U7121 ( .A1(n5388), .A2(n5387), .ZN(n8630) );
  AOI21_X1 U7122 ( .B1(n8632), .B2(n8631), .A(n8630), .ZN(n8629) );
  INV_X1 U7123 ( .A(n5388), .ZN(n7876) );
  INV_X1 U7124 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7701) );
  INV_X1 U7125 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10547) );
  MUX2_X1 U7126 ( .A(n7701), .B(n10547), .S(n5404), .Z(n5389) );
  NAND2_X1 U7127 ( .A1(n7881), .A2(n5389), .ZN(n6901) );
  OR2_X1 U7128 ( .A1(n7881), .A2(n5389), .ZN(n5390) );
  AND2_X1 U7129 ( .A1(n6901), .A2(n5390), .ZN(n7875) );
  OAI21_X1 U7130 ( .B1(n8629), .B2(n7876), .A(n7875), .ZN(n7878) );
  INV_X1 U7131 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10328) );
  MUX2_X1 U7132 ( .A(n7803), .B(n10328), .S(n5404), .Z(n5391) );
  NAND2_X1 U7133 ( .A1(n6310), .A2(n5391), .ZN(n8651) );
  OR2_X1 U7134 ( .A1(n6310), .A2(n5391), .ZN(n5392) );
  NAND2_X1 U7135 ( .A1(n8651), .A2(n5392), .ZN(n6900) );
  AOI21_X1 U7136 ( .B1(n7878), .B2(n6901), .A(n6900), .ZN(n6899) );
  INV_X1 U7137 ( .A(n8651), .ZN(n5395) );
  INV_X1 U7138 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10350) );
  INV_X1 U7139 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8647) );
  MUX2_X1 U7140 ( .A(n10350), .B(n8647), .S(n5404), .Z(n5393) );
  NAND2_X1 U7141 ( .A1(n8656), .A2(n5393), .ZN(n8677) );
  OAI21_X1 U7142 ( .B1(n8656), .B2(n5393), .A(n8677), .ZN(n8650) );
  INV_X1 U7143 ( .A(n8650), .ZN(n5394) );
  INV_X1 U7144 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8982) );
  MUX2_X1 U7145 ( .A(n10356), .B(n8982), .S(n5404), .Z(n5396) );
  NAND2_X1 U7146 ( .A1(n8671), .A2(n5396), .ZN(n5398) );
  OR2_X1 U7147 ( .A1(n8671), .A2(n5396), .ZN(n5397) );
  NAND2_X1 U7148 ( .A1(n5398), .A2(n5397), .ZN(n8676) );
  XOR2_X1 U7149 ( .A(n5399), .B(n8695), .Z(n8690) );
  AOI21_X1 U7150 ( .B1(n8695), .B2(n5400), .A(n8689), .ZN(n8709) );
  INV_X1 U7151 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n10563) );
  MUX2_X1 U7152 ( .A(n8909), .B(n10563), .S(n5404), .Z(n5401) );
  NOR2_X1 U7153 ( .A1(n8717), .A2(n5401), .ZN(n8707) );
  NAND2_X1 U7154 ( .A1(n8717), .A2(n5401), .ZN(n8705) );
  OAI21_X1 U7155 ( .B1(n8709), .B2(n8707), .A(n8705), .ZN(n8727) );
  MUX2_X1 U7156 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n5404), .Z(n5402) );
  XNOR2_X1 U7157 ( .A(n6357), .B(n5402), .ZN(n8726) );
  INV_X1 U7158 ( .A(n5402), .ZN(n5403) );
  AOI22_X1 U7159 ( .A1(n8727), .A2(n8726), .B1(n6357), .B2(n5403), .ZN(n5406)
         );
  MUX2_X1 U7160 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n5404), .Z(n5405) );
  NOR2_X1 U7161 ( .A1(n5406), .A2(n5405), .ZN(n8754) );
  NAND2_X1 U7162 ( .A1(n5406), .A2(n5405), .ZN(n8752) );
  OAI21_X1 U7163 ( .B1(n8754), .B2(n8765), .A(n8752), .ZN(n5407) );
  INV_X1 U7164 ( .A(n5409), .ZN(n8589) );
  NAND2_X1 U7165 ( .A1(n5412), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5414) );
  INV_X1 U7166 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10232) );
  INV_X1 U7167 ( .A(n5414), .ZN(n5415) );
  XNOR2_X1 U7168 ( .A(n5416), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n6983) );
  INV_X1 U7169 ( .A(n5419), .ZN(n7216) );
  INV_X1 U7170 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10238) );
  XNOR2_X1 U7171 ( .A(n6219), .B(n10238), .ZN(n7217) );
  NAND2_X1 U7172 ( .A1(n7180), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7179) );
  INV_X1 U7173 ( .A(n5421), .ZN(n7013) );
  XNOR2_X1 U7174 ( .A(n6242), .B(n10242), .ZN(n7014) );
  INV_X1 U7175 ( .A(n6242), .ZN(n7021) );
  XNOR2_X1 U7176 ( .A(n6274), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n6911) );
  NAND2_X1 U7177 ( .A1(n5425), .A2(n4923), .ZN(n5426) );
  INV_X1 U7178 ( .A(n5426), .ZN(n8624) );
  XNOR2_X1 U7179 ( .A(n8637), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n8623) );
  INV_X1 U7180 ( .A(n7881), .ZN(n6973) );
  INV_X1 U7181 ( .A(n5429), .ZN(n6892) );
  XNOR2_X1 U7182 ( .A(n6310), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n6891) );
  INV_X1 U7183 ( .A(n8656), .ZN(n7086) );
  INV_X1 U7184 ( .A(n5432), .ZN(n8664) );
  XNOR2_X1 U7185 ( .A(n8671), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n8663) );
  NAND2_X1 U7186 ( .A1(n5433), .A2(n4915), .ZN(n5434) );
  INV_X1 U7187 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10373) );
  XNOR2_X1 U7188 ( .A(n8717), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U7189 ( .A1(n5435), .A2(n6357), .ZN(n5437) );
  NAND2_X2 U7190 ( .A1(n5436), .A2(n8731), .ZN(n8743) );
  AND2_X2 U7191 ( .A1(n5437), .A2(n8743), .ZN(n8735) );
  NAND2_X2 U7192 ( .A1(n8735), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8744) );
  INV_X1 U7193 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n10504) );
  OR2_X1 U7194 ( .A1(n8765), .A2(n10504), .ZN(n5440) );
  NAND2_X1 U7195 ( .A1(n8765), .A2(n10504), .ZN(n5438) );
  AND2_X1 U7196 ( .A1(n5440), .A2(n5438), .ZN(n8741) );
  INV_X1 U7197 ( .A(n5441), .ZN(n5442) );
  INV_X1 U7198 ( .A(n5443), .ZN(n6967) );
  INV_X2 U7199 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5868) );
  INV_X1 U7200 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5447) );
  NOR2_X1 U7201 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5450) );
  AND2_X1 U7202 ( .A1(n5450), .A2(n5449), .ZN(n5453) );
  INV_X1 U7203 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U7204 ( .A1(n5458), .A2(n5471), .ZN(n5459) );
  NOR2_X1 U7205 ( .A1(n5459), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n5460) );
  INV_X1 U7206 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n10047) );
  NAND2_X1 U7207 ( .A1(n10047), .A2(n5474), .ZN(n5461) );
  INV_X1 U7208 ( .A(n5463), .ZN(n5462) );
  NAND2_X2 U7209 ( .A1(n5467), .A2(n5465), .ZN(n6094) );
  INV_X1 U7210 ( .A(n6094), .ZN(n5517) );
  INV_X1 U7211 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7475) );
  AOI22_X1 U7212 ( .A1(n5517), .A2(n7475), .B1(n5909), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n5469) );
  INV_X4 U7213 ( .A(n5836), .ZN(n5895) );
  AOI22_X1 U7214 ( .A1(n5895), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n5551), .B2(
        P1_REG0_REG_3__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U7215 ( .A1(n6108), .A2(n5471), .ZN(n5472) );
  INV_X1 U7216 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6941) );
  INV_X8 U7217 ( .A(n6929), .ZN(n8144) );
  INV_X1 U7218 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6926) );
  INV_X1 U7219 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6948) );
  INV_X1 U7220 ( .A(SI_2_), .ZN(n5478) );
  INV_X1 U7221 ( .A(SI_1_), .ZN(n5479) );
  NAND2_X1 U7222 ( .A1(n5480), .A2(n5479), .ZN(n5523) );
  INV_X1 U7223 ( .A(n5536), .ZN(n5481) );
  NAND2_X1 U7224 ( .A1(n5482), .A2(SI_1_), .ZN(n5535) );
  INV_X1 U7225 ( .A(n5535), .ZN(n5483) );
  INV_X1 U7226 ( .A(n5484), .ZN(n5485) );
  NAND2_X1 U7227 ( .A1(n5485), .A2(SI_2_), .ZN(n5538) );
  NAND2_X1 U7228 ( .A1(n5486), .A2(SI_3_), .ZN(n5558) );
  INV_X1 U7229 ( .A(n5486), .ZN(n5488) );
  INV_X1 U7230 ( .A(SI_3_), .ZN(n5487) );
  NAND2_X1 U7231 ( .A1(n5488), .A2(n5487), .ZN(n5556) );
  NAND2_X1 U7232 ( .A1(n5558), .A2(n5556), .ZN(n5490) );
  NAND2_X1 U7233 ( .A1(n5489), .A2(n5490), .ZN(n5492) );
  INV_X1 U7234 ( .A(n5490), .ZN(n5491) );
  NAND2_X1 U7235 ( .A1(n5557), .A2(n5491), .ZN(n5499) );
  NAND2_X1 U7236 ( .A1(n5492), .A2(n5499), .ZN(n6942) );
  OR2_X1 U7237 ( .A1(n5676), .A2(n6942), .ZN(n5494) );
  OR2_X1 U7238 ( .A1(n4683), .A2(n10046), .ZN(n5496) );
  NAND2_X1 U7239 ( .A1(n4431), .A2(n9596), .ZN(n5493) );
  NAND2_X1 U7240 ( .A1(n7447), .A2(n9450), .ZN(n9414) );
  NAND2_X1 U7241 ( .A1(n8129), .A2(n10132), .ZN(n7441) );
  NAND2_X1 U7242 ( .A1(n5496), .A2(n10272), .ZN(n5497) );
  NAND2_X1 U7243 ( .A1(n5497), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5498) );
  XNOR2_X1 U7244 ( .A(n5498), .B(n5456), .ZN(n9608) );
  NAND2_X1 U7245 ( .A1(n5499), .A2(n5558), .ZN(n5504) );
  INV_X1 U7246 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6927) );
  INV_X1 U7247 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6944) );
  MUX2_X1 U7248 ( .A(n6927), .B(n6944), .S(n5584), .Z(n5501) );
  INV_X1 U7249 ( .A(SI_4_), .ZN(n5500) );
  INV_X1 U7250 ( .A(n5501), .ZN(n5502) );
  NAND2_X1 U7251 ( .A1(n5502), .A2(SI_4_), .ZN(n5561) );
  AND2_X1 U7252 ( .A1(n5559), .A2(n5561), .ZN(n5503) );
  XNOR2_X1 U7253 ( .A(n5504), .B(n5503), .ZN(n6943) );
  AOI22_X1 U7254 ( .A1(n5895), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n5909), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n5510) );
  OAI21_X1 U7255 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5549), .ZN(n7401) );
  NAND2_X1 U7256 ( .A1(n5551), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5507) );
  OAI21_X1 U7257 ( .B1(n7401), .B2(n6094), .A(n5507), .ZN(n5508) );
  INV_X1 U7258 ( .A(n5508), .ZN(n5509) );
  NAND2_X1 U7259 ( .A1(n7948), .A2(n7452), .ZN(n9291) );
  NAND2_X2 U7260 ( .A1(n9451), .A2(n9291), .ZN(n9412) );
  NAND2_X1 U7261 ( .A1(n5895), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5515) );
  NAND2_X1 U7262 ( .A1(n5517), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U7263 ( .A1(n5769), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U7264 ( .A1(n8144), .A2(SI_0_), .ZN(n5516) );
  XNOR2_X1 U7265 ( .A(n5516), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10062) );
  NAND2_X1 U7266 ( .A1(n7808), .A2(n7742), .ZN(n7807) );
  NAND2_X1 U7267 ( .A1(n5517), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7268 ( .A1(n5895), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7269 ( .A1(n5551), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5518) );
  INV_X1 U7270 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7271 ( .A1(n5535), .A2(n5523), .ZN(n5537) );
  XNOR2_X1 U7272 ( .A(n5536), .B(n5537), .ZN(n6936) );
  NAND2_X1 U7273 ( .A1(n7411), .A2(n6601), .ZN(n5524) );
  NAND2_X1 U7274 ( .A1(n7807), .A2(n5524), .ZN(n5526) );
  NAND2_X1 U7275 ( .A1(n9448), .A2(n7378), .ZN(n5525) );
  NAND2_X1 U7276 ( .A1(n5526), .A2(n5525), .ZN(n7364) );
  NAND2_X1 U7277 ( .A1(n5895), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U7278 ( .A1(n5517), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U7279 ( .A1(n5909), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5528) );
  NOR2_X1 U7280 ( .A1(n5531), .A2(n10046), .ZN(n5532) );
  MUX2_X1 U7281 ( .A(n10046), .B(n5532), .S(P1_IR_REG_2__SCAN_IN), .Z(n5533)
         );
  INV_X1 U7282 ( .A(n5533), .ZN(n5534) );
  OAI21_X1 U7283 ( .B1(n5537), .B2(n5536), .A(n5535), .ZN(n5541) );
  AND2_X1 U7284 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  XNOR2_X1 U7285 ( .A(n5541), .B(n5540), .ZN(n6947) );
  OR2_X1 U7286 ( .A1(n5676), .A2(n6947), .ZN(n5542) );
  NAND2_X1 U7287 ( .A1(n7947), .A2(n6097), .ZN(n6072) );
  INV_X1 U7288 ( .A(n6097), .ZN(n8131) );
  NAND2_X1 U7289 ( .A1(n9561), .A2(n8131), .ZN(n9452) );
  NAND2_X1 U7290 ( .A1(n7947), .A2(n8131), .ZN(n7440) );
  AND2_X1 U7291 ( .A1(n7441), .A2(n7440), .ZN(n5544) );
  NAND2_X1 U7292 ( .A1(n7363), .A2(n5544), .ZN(n5545) );
  NAND2_X1 U7293 ( .A1(n5546), .A2(n5545), .ZN(n7442) );
  INV_X2 U7294 ( .A(n6094), .ZN(n6047) );
  INV_X1 U7295 ( .A(n5549), .ZN(n5547) );
  INV_X1 U7296 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U7297 ( .A1(n5549), .A2(n5548), .ZN(n5550) );
  AND2_X1 U7298 ( .A1(n5579), .A2(n5550), .ZN(n7509) );
  NAND2_X1 U7299 ( .A1(n6047), .A2(n7509), .ZN(n5555) );
  NAND2_X1 U7300 ( .A1(n5895), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5554) );
  INV_X1 U7301 ( .A(n5551), .ZN(n5789) );
  NAND2_X1 U7302 ( .A1(n5551), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5553) );
  INV_X1 U7303 ( .A(n5909), .ZN(n5643) );
  NAND2_X1 U7304 ( .A1(n5909), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5552) );
  INV_X1 U7305 ( .A(n9558), .ZN(n5576) );
  INV_X1 U7306 ( .A(n5558), .ZN(n5560) );
  NAND2_X1 U7307 ( .A1(n5560), .A2(n5559), .ZN(n5562) );
  AND2_X1 U7308 ( .A1(n5562), .A2(n5561), .ZN(n5563) );
  INV_X1 U7309 ( .A(n5615), .ZN(n5568) );
  INV_X1 U7310 ( .A(SI_5_), .ZN(n10294) );
  NAND2_X1 U7311 ( .A1(n5610), .A2(n5613), .ZN(n5569) );
  NAND2_X1 U7312 ( .A1(n5568), .A2(n5569), .ZN(n5571) );
  INV_X1 U7313 ( .A(n5569), .ZN(n5570) );
  NAND2_X1 U7314 ( .A1(n5615), .A2(n5570), .ZN(n5583) );
  NAND2_X1 U7315 ( .A1(n5571), .A2(n5583), .ZN(n6239) );
  OR2_X1 U7316 ( .A1(n6239), .A2(n5676), .ZN(n5575) );
  INV_X1 U7317 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6954) );
  OR2_X1 U7318 ( .A1(n8151), .A2(n6954), .ZN(n5574) );
  NAND2_X1 U7319 ( .A1(n4683), .A2(n5222), .ZN(n5590) );
  NAND2_X1 U7320 ( .A1(n5590), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5572) );
  XNOR2_X1 U7321 ( .A(n5572), .B(P1_IR_REG_5__SCAN_IN), .ZN(n7058) );
  NAND2_X1 U7322 ( .A1(n4432), .A2(n7058), .ZN(n5573) );
  AND3_X2 U7323 ( .A1(n5575), .A2(n5574), .A3(n5573), .ZN(n9304) );
  NAND2_X1 U7324 ( .A1(n5576), .A2(n9304), .ZN(n7486) );
  NAND2_X1 U7325 ( .A1(n7948), .A2(n10116), .ZN(n7485) );
  NAND2_X1 U7326 ( .A1(n7442), .A2(n5226), .ZN(n5599) );
  NAND2_X1 U7327 ( .A1(n9558), .A2(n9304), .ZN(n9449) );
  INV_X1 U7328 ( .A(n7486), .ZN(n5596) );
  INV_X1 U7329 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7330 ( .A1(n5579), .A2(n5578), .ZN(n5580) );
  AND2_X1 U7331 ( .A1(n5603), .A2(n5580), .ZN(n10100) );
  AOI22_X1 U7332 ( .A1(n6047), .A2(n10100), .B1(n5909), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n5582) );
  AOI22_X1 U7333 ( .A1(n5895), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n5551), .B2(
        P1_REG0_REG_6__SCAN_IN), .ZN(n5581) );
  AND2_X2 U7334 ( .A1(n5582), .A2(n5581), .ZN(n9302) );
  NAND2_X1 U7335 ( .A1(n5583), .A2(n5610), .ZN(n5589) );
  INV_X1 U7336 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6935) );
  INV_X1 U7337 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6950) );
  MUX2_X1 U7338 ( .A(n6935), .B(n6950), .S(n5584), .Z(n5586) );
  INV_X1 U7339 ( .A(SI_6_), .ZN(n5585) );
  NAND2_X1 U7340 ( .A1(n5586), .A2(n5585), .ZN(n5614) );
  INV_X1 U7341 ( .A(n5586), .ZN(n5587) );
  NAND2_X1 U7342 ( .A1(n5587), .A2(SI_6_), .ZN(n5609) );
  NAND2_X1 U7343 ( .A1(n5614), .A2(n5609), .ZN(n5588) );
  NAND2_X1 U7344 ( .A1(n6934), .A2(n5505), .ZN(n5594) );
  NOR2_X2 U7345 ( .A1(n5590), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5634) );
  INV_X1 U7346 ( .A(n5634), .ZN(n5591) );
  NAND2_X1 U7347 ( .A1(n5591), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5624) );
  XNOR2_X1 U7348 ( .A(n5624), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7197) );
  NOR2_X1 U7349 ( .A1(n5210), .A2(n5592), .ZN(n5593) );
  NAND2_X1 U7350 ( .A1(n9302), .A2(n5595), .ZN(n9293) );
  INV_X2 U7351 ( .A(n5595), .ZN(n10103) );
  NAND2_X1 U7352 ( .A1(n9293), .A2(n9415), .ZN(n7491) );
  OAI21_X1 U7353 ( .B1(n9413), .B2(n5596), .A(n7491), .ZN(n5597) );
  INV_X1 U7354 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U7355 ( .A1(n9302), .A2(n10103), .ZN(n5600) );
  INV_X1 U7356 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5602) );
  NAND2_X1 U7357 ( .A1(n5603), .A2(n5602), .ZN(n5604) );
  AND2_X1 U7358 ( .A1(n5641), .A2(n5604), .ZN(n7645) );
  NAND2_X1 U7359 ( .A1(n6047), .A2(n7645), .ZN(n5608) );
  NAND2_X1 U7360 ( .A1(n5895), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U7361 ( .A1(n5551), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7362 ( .A1(n5909), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5605) );
  NAND4_X1 U7363 ( .A1(n5608), .A2(n5607), .A3(n5606), .A4(n5605), .ZN(n9556)
         );
  INV_X1 U7364 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6933) );
  INV_X1 U7365 ( .A(n5614), .ZN(n5611) );
  INV_X1 U7366 ( .A(n5612), .ZN(n5617) );
  MUX2_X1 U7367 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5778), .Z(n5618) );
  OAI21_X1 U7368 ( .B1(n5618), .B2(SI_7_), .A(n5631), .ZN(n5620) );
  NAND2_X1 U7369 ( .A1(n5619), .A2(n5620), .ZN(n5623) );
  INV_X1 U7370 ( .A(n5620), .ZN(n5621) );
  NAND2_X1 U7371 ( .A1(n5623), .A2(n5632), .ZN(n6932) );
  INV_X1 U7372 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n10476) );
  NAND2_X1 U7373 ( .A1(n5624), .A2(n10476), .ZN(n5625) );
  NAND2_X1 U7374 ( .A1(n5625), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5626) );
  XNOR2_X1 U7375 ( .A(n5626), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7198) );
  NAND2_X1 U7376 ( .A1(n4432), .A2(n7198), .ZN(n5627) );
  OAI211_X1 U7377 ( .C1(n8151), .C2(n6933), .A(n5628), .B(n5627), .ZN(n5629)
         );
  NAND2_X1 U7378 ( .A1(n7616), .A2(n9408), .ZN(n9299) );
  NAND2_X1 U7379 ( .A1(n7984), .A2(n7762), .ZN(n5630) );
  MUX2_X1 U7380 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n5778), .Z(n5648) );
  XNOR2_X1 U7381 ( .A(n5653), .B(n5652), .ZN(n6937) );
  NAND2_X1 U7382 ( .A1(n6937), .A2(n5505), .ZN(n5639) );
  NAND2_X1 U7383 ( .A1(n5634), .A2(n5633), .ZN(n5636) );
  MUX2_X1 U7384 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5635), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5637) );
  NOR2_X2 U7385 ( .A1(n5636), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6057) );
  AND2_X1 U7386 ( .A1(n5637), .A2(n5677), .ZN(n7286) );
  AOI22_X1 U7387 ( .A1(n5876), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n4432), .B2(
        n7286), .ZN(n5638) );
  NAND2_X1 U7388 ( .A1(n5895), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5647) );
  NAND2_X1 U7389 ( .A1(n5641), .A2(n5640), .ZN(n5642) );
  AND2_X1 U7390 ( .A1(n5659), .A2(n5642), .ZN(n7981) );
  NAND2_X1 U7391 ( .A1(n6047), .A2(n7981), .ZN(n5646) );
  NAND2_X1 U7392 ( .A1(n5909), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U7393 ( .A1(n5769), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5644) );
  NAND4_X1 U7394 ( .A1(n5647), .A2(n5646), .A3(n5645), .A4(n5644), .ZN(n9555)
         );
  NAND2_X1 U7395 ( .A1(n7783), .A2(n9555), .ZN(n9314) );
  INV_X1 U7396 ( .A(n9555), .ZN(n9202) );
  NAND2_X1 U7397 ( .A1(n9202), .A2(n7986), .ZN(n9319) );
  NAND2_X1 U7398 ( .A1(n9314), .A2(n9319), .ZN(n7615) );
  INV_X1 U7399 ( .A(n5648), .ZN(n5650) );
  INV_X1 U7400 ( .A(SI_8_), .ZN(n5649) );
  NAND2_X1 U7401 ( .A1(n5650), .A2(n5649), .ZN(n5651) );
  NAND2_X1 U7402 ( .A1(n6958), .A2(n5505), .ZN(n5656) );
  XNOR2_X1 U7403 ( .A(n5654), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7201) );
  AOI22_X1 U7404 ( .A1(n5876), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n4432), .B2(
        n7201), .ZN(n5655) );
  INV_X1 U7405 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U7406 ( .A1(n5659), .A2(n5658), .ZN(n5660) );
  AND2_X1 U7407 ( .A1(n5696), .A2(n5660), .ZN(n9200) );
  NAND2_X1 U7408 ( .A1(n6047), .A2(n9200), .ZN(n5664) );
  NAND2_X1 U7409 ( .A1(n5895), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U7410 ( .A1(n5769), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7411 ( .A1(n5909), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5661) );
  NAND4_X1 U7412 ( .A1(n5664), .A2(n5663), .A3(n5662), .A4(n5661), .ZN(n9554)
         );
  NAND2_X1 U7413 ( .A1(n9342), .A2(n9323), .ZN(n7668) );
  OR2_X1 U7414 ( .A1(n4572), .A2(n9554), .ZN(n5665) );
  NAND2_X1 U7415 ( .A1(n5669), .A2(SI_10_), .ZN(n5686) );
  INV_X1 U7416 ( .A(n5669), .ZN(n5671) );
  INV_X1 U7417 ( .A(SI_10_), .ZN(n5670) );
  NAND2_X1 U7418 ( .A1(n5671), .A2(n5670), .ZN(n5672) );
  NAND2_X1 U7419 ( .A1(n5686), .A2(n5672), .ZN(n5674) );
  INV_X1 U7420 ( .A(n5674), .ZN(n5673) );
  OR2_X1 U7421 ( .A1(n5677), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5678) );
  XNOR2_X1 U7422 ( .A(n5689), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7317) );
  AOI22_X1 U7423 ( .A1(n5876), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n4432), .B2(
        n7317), .ZN(n5679) );
  NAND2_X2 U7424 ( .A1(n5680), .A2(n5679), .ZN(n9113) );
  XNOR2_X1 U7425 ( .A(n5696), .B(P1_REG3_REG_10__SCAN_IN), .ZN(n9109) );
  NAND2_X1 U7426 ( .A1(n6047), .A2(n9109), .ZN(n5684) );
  NAND2_X1 U7427 ( .A1(n5895), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U7428 ( .A1(n5909), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U7429 ( .A1(n5769), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5681) );
  NAND4_X1 U7430 ( .A1(n5684), .A2(n5683), .A3(n5682), .A4(n5681), .ZN(n9553)
         );
  INV_X1 U7431 ( .A(n9553), .ZN(n7724) );
  NAND2_X1 U7432 ( .A1(n9113), .A2(n7724), .ZN(n9344) );
  OR2_X1 U7433 ( .A1(n9113), .A2(n9553), .ZN(n5685) );
  XNOR2_X1 U7434 ( .A(n5707), .B(n5706), .ZN(n6963) );
  NAND2_X1 U7435 ( .A1(n6963), .A2(n5505), .ZN(n5693) );
  INV_X1 U7436 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U7437 ( .A1(n5689), .A2(n5688), .ZN(n5690) );
  AOI22_X1 U7438 ( .A1(n5876), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n4432), .B2(
        n7517), .ZN(n5692) );
  INV_X1 U7439 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5695) );
  INV_X1 U7440 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5694) );
  OAI21_X1 U7441 ( .B1(n5696), .B2(n5695), .A(n5694), .ZN(n5697) );
  AND2_X1 U7442 ( .A1(n5697), .A2(n5723), .ZN(n9246) );
  NAND2_X1 U7443 ( .A1(n6047), .A2(n9246), .ZN(n5701) );
  NAND2_X1 U7444 ( .A1(n5895), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7445 ( .A1(n5551), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U7446 ( .A1(n5894), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5698) );
  NAND4_X1 U7447 ( .A1(n5701), .A2(n5700), .A3(n5699), .A4(n5698), .ZN(n9552)
         );
  NAND2_X1 U7448 ( .A1(n9326), .A2(n9552), .ZN(n5702) );
  INV_X1 U7449 ( .A(n5703), .ZN(n5704) );
  NAND2_X1 U7450 ( .A1(n5704), .A2(n10559), .ZN(n5705) );
  NAND2_X1 U7451 ( .A1(n5708), .A2(SI_12_), .ZN(n5752) );
  INV_X1 U7452 ( .A(n5708), .ZN(n5710) );
  INV_X1 U7453 ( .A(SI_12_), .ZN(n5709) );
  NAND2_X1 U7454 ( .A1(n5710), .A2(n5709), .ZN(n5751) );
  NAND2_X1 U7455 ( .A1(n5752), .A2(n5751), .ZN(n5711) );
  NAND2_X1 U7456 ( .A1(n5759), .A2(n5711), .ZN(n5712) );
  NAND2_X1 U7457 ( .A1(n6975), .A2(n5505), .ZN(n5722) );
  NOR2_X1 U7458 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5719) );
  NOR2_X1 U7459 ( .A1(n5714), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5718) );
  NOR2_X1 U7460 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5715) );
  AND2_X1 U7461 ( .A1(n5716), .A2(n5715), .ZN(n5717) );
  NAND4_X1 U7462 ( .A1(n4683), .A2(n5719), .A3(n5718), .A4(n5717), .ZN(n5737)
         );
  NAND2_X1 U7463 ( .A1(n5737), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5720) );
  XNOR2_X1 U7464 ( .A(n5720), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7524) );
  AOI22_X1 U7465 ( .A1(n5876), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n4432), .B2(
        n7524), .ZN(n5721) );
  INV_X1 U7466 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10384) );
  NAND2_X1 U7467 ( .A1(n5723), .A2(n10384), .ZN(n5724) );
  AND2_X1 U7468 ( .A1(n5743), .A2(n5724), .ZN(n9142) );
  NAND2_X1 U7469 ( .A1(n6047), .A2(n9142), .ZN(n5728) );
  NAND2_X1 U7470 ( .A1(n5895), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5727) );
  NAND2_X1 U7471 ( .A1(n6153), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U7472 ( .A1(n5894), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5725) );
  NAND4_X1 U7473 ( .A1(n5728), .A2(n5727), .A3(n5726), .A4(n5725), .ZN(n9916)
         );
  NAND2_X1 U7474 ( .A1(n7867), .A2(n9916), .ZN(n9349) );
  NAND2_X1 U7475 ( .A1(n9145), .A2(n9251), .ZN(n9465) );
  NAND2_X1 U7476 ( .A1(n9349), .A2(n9465), .ZN(n9407) );
  NAND2_X1 U7477 ( .A1(n7861), .A2(n9407), .ZN(n5730) );
  NAND2_X1 U7478 ( .A1(n7867), .A2(n9251), .ZN(n5729) );
  NAND2_X1 U7479 ( .A1(n5730), .A2(n5729), .ZN(n9924) );
  NAND2_X1 U7480 ( .A1(n5731), .A2(n5752), .ZN(n5736) );
  INV_X1 U7481 ( .A(SI_13_), .ZN(n5732) );
  INV_X1 U7482 ( .A(n5733), .ZN(n5734) );
  NAND2_X1 U7483 ( .A1(n5734), .A2(SI_13_), .ZN(n5755) );
  NAND2_X1 U7484 ( .A1(n5753), .A2(n5755), .ZN(n5735) );
  XNOR2_X2 U7485 ( .A(n5736), .B(n5735), .ZN(n7085) );
  NAND2_X1 U7486 ( .A1(n7085), .A2(n5505), .ZN(n5741) );
  INV_X1 U7487 ( .A(n5737), .ZN(n5738) );
  NAND2_X1 U7488 ( .A1(n5738), .A2(n10400), .ZN(n5761) );
  XNOR2_X1 U7489 ( .A(n5739), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7653) );
  AOI22_X1 U7490 ( .A1(n5876), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n4432), .B2(
        n7653), .ZN(n5740) );
  INV_X1 U7491 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5742) );
  NAND2_X1 U7492 ( .A1(n5743), .A2(n5742), .ZN(n5744) );
  AND2_X1 U7493 ( .A1(n5767), .A2(n5744), .ZN(n9921) );
  NAND2_X1 U7494 ( .A1(n6047), .A2(n9921), .ZN(n5748) );
  NAND2_X1 U7495 ( .A1(n5895), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5747) );
  INV_X1 U7496 ( .A(n5789), .ZN(n6153) );
  NAND2_X1 U7497 ( .A1(n6153), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U7498 ( .A1(n5894), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5745) );
  NAND4_X1 U7499 ( .A1(n5748), .A2(n5747), .A3(n5746), .A4(n5745), .ZN(n9551)
         );
  INV_X1 U7500 ( .A(n9551), .ZN(n9899) );
  NAND2_X1 U7501 ( .A1(n9924), .A2(n9925), .ZN(n5750) );
  OR2_X1 U7502 ( .A1(n10008), .A2(n9551), .ZN(n5749) );
  NAND2_X1 U7503 ( .A1(n5750), .A2(n5749), .ZN(n9887) );
  INV_X1 U7504 ( .A(n5752), .ZN(n5754) );
  NAND2_X1 U7505 ( .A1(n5754), .A2(n5753), .ZN(n5756) );
  MUX2_X1 U7506 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n8144), .Z(n5776) );
  XNOR2_X1 U7507 ( .A(n5776), .B(SI_14_), .ZN(n5760) );
  XNOR2_X1 U7508 ( .A(n5777), .B(n5760), .ZN(n7122) );
  NAND2_X1 U7509 ( .A1(n7122), .A2(n5505), .ZN(n5765) );
  INV_X1 U7510 ( .A(n5761), .ZN(n5763) );
  NAND2_X1 U7511 ( .A1(n5763), .A2(n5762), .ZN(n5802) );
  XNOR2_X1 U7512 ( .A(n5781), .B(P1_IR_REG_14__SCAN_IN), .ZN(n8203) );
  AOI22_X1 U7513 ( .A1(n5876), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n4432), .B2(
        n8203), .ZN(n5764) );
  INV_X1 U7514 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5766) );
  NAND2_X1 U7515 ( .A1(n5767), .A2(n5766), .ZN(n5768) );
  AND2_X1 U7516 ( .A1(n5787), .A2(n5768), .ZN(n9891) );
  NAND2_X1 U7517 ( .A1(n6047), .A2(n9891), .ZN(n5773) );
  NAND2_X1 U7518 ( .A1(n5895), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5772) );
  INV_X1 U7519 ( .A(n5789), .ZN(n5769) );
  NAND2_X1 U7520 ( .A1(n5769), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5771) );
  NAND2_X1 U7521 ( .A1(n5894), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5770) );
  NAND4_X1 U7522 ( .A1(n5773), .A2(n5772), .A3(n5771), .A4(n5770), .ZN(n9914)
         );
  NOR2_X1 U7523 ( .A1(n10003), .A2(n9914), .ZN(n5775) );
  NAND2_X1 U7524 ( .A1(n10003), .A2(n9914), .ZN(n5774) );
  MUX2_X1 U7525 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n8144), .Z(n5825) );
  XNOR2_X1 U7526 ( .A(n5825), .B(SI_15_), .ZN(n5779) );
  XNOR2_X1 U7527 ( .A(n5820), .B(n5779), .ZN(n7331) );
  NAND2_X1 U7528 ( .A1(n7331), .A2(n5505), .ZN(n5785) );
  NAND2_X1 U7529 ( .A1(n5781), .A2(n5780), .ZN(n5782) );
  XNOR2_X1 U7530 ( .A(n5783), .B(P1_IR_REG_15__SCAN_IN), .ZN(n8205) );
  AOI22_X1 U7531 ( .A1(n5876), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n4432), .B2(
        n8205), .ZN(n5784) );
  NAND2_X2 U7532 ( .A1(n5785), .A2(n5784), .ZN(n9998) );
  NAND2_X1 U7533 ( .A1(n5895), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5793) );
  INV_X1 U7534 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5786) );
  NAND2_X1 U7535 ( .A1(n5787), .A2(n5786), .ZN(n5788) );
  AND2_X1 U7536 ( .A1(n5810), .A2(n5788), .ZN(n9278) );
  NAND2_X1 U7537 ( .A1(n5517), .A2(n9278), .ZN(n5792) );
  NAND2_X1 U7538 ( .A1(n5894), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5791) );
  NAND2_X1 U7539 ( .A1(n6153), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5790) );
  NAND4_X1 U7540 ( .A1(n5793), .A2(n5792), .A3(n5791), .A4(n5790), .ZN(n9868)
         );
  AND2_X1 U7541 ( .A1(n9998), .A2(n9868), .ZN(n9878) );
  NAND2_X1 U7542 ( .A1(n5820), .A2(SI_15_), .ZN(n5794) );
  NAND2_X1 U7543 ( .A1(n5794), .A2(n5822), .ZN(n5798) );
  INV_X1 U7544 ( .A(n5820), .ZN(n5796) );
  INV_X1 U7545 ( .A(SI_15_), .ZN(n5795) );
  NAND2_X1 U7546 ( .A1(n5798), .A2(n5797), .ZN(n5801) );
  INV_X1 U7547 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5799) );
  INV_X1 U7548 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7408) );
  MUX2_X1 U7549 ( .A(n5799), .B(n7408), .S(n8144), .Z(n5823) );
  XNOR2_X1 U7550 ( .A(n5823), .B(SI_16_), .ZN(n5800) );
  NAND2_X1 U7551 ( .A1(n7372), .A2(n5505), .ZN(n5806) );
  NOR2_X1 U7552 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5803) );
  NAND2_X1 U7553 ( .A1(n4521), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5804) );
  XNOR2_X1 U7554 ( .A(n5804), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9641) );
  AOI22_X1 U7555 ( .A1(n5876), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n4432), .B2(
        n9641), .ZN(n5805) );
  INV_X1 U7556 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5809) );
  NAND2_X1 U7557 ( .A1(n5810), .A2(n5809), .ZN(n5811) );
  AND2_X1 U7558 ( .A1(n9179), .A2(n5811), .ZN(n9873) );
  NAND2_X1 U7559 ( .A1(n6047), .A2(n9873), .ZN(n5815) );
  NAND2_X1 U7560 ( .A1(n5895), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7561 ( .A1(n5894), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7562 ( .A1(n6153), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5812) );
  NAND4_X1 U7563 ( .A1(n5815), .A2(n5814), .A3(n5813), .A4(n5812), .ZN(n9550)
         );
  AND2_X1 U7564 ( .A1(n5807), .A2(n9550), .ZN(n5817) );
  INV_X1 U7565 ( .A(n9550), .ZN(n9177) );
  OR2_X1 U7566 ( .A1(n6720), .A2(n9177), .ZN(n9476) );
  NAND2_X1 U7567 ( .A1(n6720), .A2(n9177), .ZN(n6080) );
  AND2_X2 U7568 ( .A1(n9476), .A2(n6080), .ZN(n9883) );
  OR2_X1 U7569 ( .A1(n9998), .A2(n9868), .ZN(n9881) );
  INV_X1 U7570 ( .A(n9881), .ZN(n5816) );
  NOR2_X1 U7571 ( .A1(n5817), .A2(n9880), .ZN(n5818) );
  INV_X1 U7572 ( .A(SI_16_), .ZN(n5821) );
  AOI22_X1 U7573 ( .A1(n5795), .A2(n5822), .B1(n5823), .B2(n5821), .ZN(n5819)
         );
  OAI21_X1 U7574 ( .B1(n5822), .B2(n5795), .A(n5821), .ZN(n5827) );
  INV_X1 U7575 ( .A(n5823), .ZN(n5826) );
  AND2_X1 U7576 ( .A1(SI_16_), .A2(SI_15_), .ZN(n5824) );
  AOI22_X1 U7577 ( .A1(n5827), .A2(n5826), .B1(n5825), .B2(n5824), .ZN(n5828)
         );
  INV_X1 U7578 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5829) );
  MUX2_X1 U7579 ( .A(n7342), .B(n5829), .S(n8144), .Z(n5831) );
  INV_X1 U7580 ( .A(SI_17_), .ZN(n5830) );
  INV_X1 U7581 ( .A(n5831), .ZN(n5832) );
  NAND2_X1 U7582 ( .A1(n5832), .A2(SI_17_), .ZN(n5833) );
  NAND2_X1 U7583 ( .A1(n5843), .A2(n5833), .ZN(n5844) );
  XNOR2_X1 U7584 ( .A(n5845), .B(n5844), .ZN(n7328) );
  NAND2_X1 U7585 ( .A1(n7328), .A2(n5505), .ZN(n5835) );
  XNOR2_X1 U7586 ( .A(n5846), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9651) );
  AOI22_X1 U7587 ( .A1(n5876), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n4432), .B2(
        n9651), .ZN(n5834) );
  INV_X1 U7588 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8208) );
  XNOR2_X1 U7589 ( .A(n9179), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n8225) );
  NAND2_X1 U7590 ( .A1(n8225), .A2(n6047), .ZN(n5841) );
  NAND2_X1 U7591 ( .A1(n5551), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U7592 ( .A1(n5894), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5838) );
  AND2_X1 U7593 ( .A1(n5839), .A2(n5838), .ZN(n5840) );
  OAI211_X1 U7594 ( .C1(n5837), .C2(n8208), .A(n5841), .B(n5840), .ZN(n9867)
         );
  MUX2_X1 U7595 ( .A(n10411), .B(n7482), .S(n8144), .Z(n5860) );
  XNOR2_X1 U7596 ( .A(n5863), .B(n5859), .ZN(n7481) );
  NAND2_X1 U7597 ( .A1(n7481), .A2(n5505), .ZN(n5851) );
  INV_X1 U7598 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n10488) );
  NAND2_X1 U7599 ( .A1(n5847), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U7600 ( .A1(n4847), .A2(n5868), .ZN(n5848) );
  AOI22_X1 U7601 ( .A1(n5876), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n4432), .B2(
        n8209), .ZN(n5850) );
  NAND2_X2 U7602 ( .A1(n5851), .A2(n5850), .ZN(n9983) );
  INV_X1 U7603 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9859) );
  INV_X1 U7604 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9647) );
  INV_X1 U7605 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5852) );
  OAI21_X1 U7606 ( .B1(n9179), .B2(n9647), .A(n5852), .ZN(n5854) );
  NAND2_X1 U7607 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n5853) );
  AND2_X1 U7608 ( .A1(n5854), .A2(n5879), .ZN(n9857) );
  NAND2_X1 U7609 ( .A1(n9857), .A2(n6047), .ZN(n5856) );
  AOI22_X1 U7610 ( .A1(n5909), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n6153), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5855) );
  OAI211_X1 U7611 ( .C1(n5837), .C2(n9859), .A(n5856), .B(n5855), .ZN(n9835)
         );
  NOR2_X1 U7612 ( .A1(n9983), .A2(n9835), .ZN(n5858) );
  NAND2_X1 U7613 ( .A1(n9983), .A2(n9835), .ZN(n5857) );
  INV_X1 U7614 ( .A(n5860), .ZN(n5861) );
  MUX2_X1 U7615 ( .A(n7501), .B(n7503), .S(n8144), .Z(n5865) );
  INV_X1 U7616 ( .A(SI_19_), .ZN(n5864) );
  INV_X1 U7617 ( .A(n5865), .ZN(n5866) );
  NAND2_X1 U7618 ( .A1(n5866), .A2(SI_19_), .ZN(n5867) );
  NAND2_X1 U7619 ( .A1(n5885), .A2(n5867), .ZN(n5886) );
  XNOR2_X1 U7620 ( .A(n5887), .B(n5886), .ZN(n7500) );
  NAND2_X1 U7621 ( .A1(n7500), .A2(n5505), .ZN(n5878) );
  INV_X1 U7622 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U7623 ( .A1(n5868), .A2(n5871), .ZN(n5874) );
  NAND2_X1 U7624 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n5869) );
  NAND2_X1 U7625 ( .A1(n5869), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5870) );
  OAI21_X1 U7626 ( .B1(n5871), .B2(P1_IR_REG_31__SCAN_IN), .A(n5870), .ZN(
        n5872) );
  AOI22_X1 U7627 ( .A1(n5876), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9511), .B2(
        n4432), .ZN(n5877) );
  INV_X1 U7628 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n5883) );
  INV_X1 U7629 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n10376) );
  NAND2_X1 U7630 ( .A1(n5879), .A2(n10376), .ZN(n5880) );
  NAND2_X1 U7631 ( .A1(n5892), .A2(n5880), .ZN(n9841) );
  OR2_X1 U7632 ( .A1(n9841), .A2(n6094), .ZN(n5882) );
  AOI22_X1 U7633 ( .A1(n5909), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n5551), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5881) );
  OAI211_X1 U7634 ( .C1(n5837), .C2(n5883), .A(n5882), .B(n5881), .ZN(n9820)
         );
  AND2_X1 U7635 ( .A1(n9975), .A2(n9820), .ZN(n5884) );
  MUX2_X1 U7636 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n8144), .Z(n5900) );
  XNOR2_X1 U7637 ( .A(n5900), .B(n10446), .ZN(n5888) );
  XNOR2_X1 U7638 ( .A(n5901), .B(n5888), .ZN(n7607) );
  NAND2_X1 U7639 ( .A1(n7607), .A2(n5505), .ZN(n5890) );
  INV_X1 U7640 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10480) );
  OR2_X1 U7641 ( .A1(n8151), .A2(n10480), .ZN(n5889) );
  INV_X1 U7642 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U7643 ( .A1(n5892), .A2(n5891), .ZN(n5893) );
  NAND2_X1 U7644 ( .A1(n5907), .A2(n5893), .ZN(n9212) );
  AOI22_X1 U7645 ( .A1(n5894), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n6153), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U7646 ( .A1(n5895), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5896) );
  OAI211_X1 U7647 ( .C1(n9212), .C2(n6094), .A(n5897), .B(n5896), .ZN(n9836)
         );
  NOR2_X1 U7648 ( .A1(n9971), .A2(n9836), .ZN(n5898) );
  NAND2_X1 U7649 ( .A1(n9971), .A2(n9836), .ZN(n5899) );
  MUX2_X1 U7650 ( .A(n7675), .B(n10416), .S(n8144), .Z(n5918) );
  XNOR2_X1 U7651 ( .A(n5918), .B(SI_21_), .ZN(n5902) );
  XNOR2_X1 U7652 ( .A(n5922), .B(n5902), .ZN(n7673) );
  NAND2_X1 U7653 ( .A1(n7673), .A2(n5505), .ZN(n5904) );
  OR2_X1 U7654 ( .A1(n8151), .A2(n10416), .ZN(n5903) );
  INV_X1 U7655 ( .A(n5907), .ZN(n5905) );
  INV_X1 U7656 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7657 ( .A1(n5907), .A2(n5906), .ZN(n5908) );
  NAND2_X1 U7658 ( .A1(n5948), .A2(n5908), .ZN(n9811) );
  OR2_X1 U7659 ( .A1(n9811), .A2(n6094), .ZN(n5915) );
  INV_X1 U7660 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U7661 ( .A1(n5909), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5911) );
  NAND2_X1 U7662 ( .A1(n5551), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5910) );
  OAI211_X1 U7663 ( .C1(n5837), .C2(n5912), .A(n5911), .B(n5910), .ZN(n5913)
         );
  INV_X1 U7664 ( .A(n5913), .ZN(n5914) );
  AND2_X1 U7665 ( .A1(n9966), .A2(n9821), .ZN(n5917) );
  NAND2_X1 U7666 ( .A1(n5919), .A2(SI_21_), .ZN(n5920) );
  INV_X1 U7667 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7842) );
  INV_X1 U7668 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7845) );
  MUX2_X1 U7669 ( .A(n7842), .B(n7845), .S(n8144), .Z(n5924) );
  INV_X1 U7670 ( .A(SI_22_), .ZN(n5923) );
  NAND2_X1 U7671 ( .A1(n5924), .A2(n5923), .ZN(n5958) );
  INV_X1 U7672 ( .A(n5924), .ZN(n5925) );
  NAND2_X1 U7673 ( .A1(n5925), .A2(SI_22_), .ZN(n5926) );
  NAND2_X1 U7674 ( .A1(n5958), .A2(n5926), .ZN(n5957) );
  XNOR2_X1 U7675 ( .A(n5981), .B(n5957), .ZN(n7840) );
  NAND2_X1 U7676 ( .A1(n7840), .A2(n5505), .ZN(n5928) );
  OR2_X1 U7677 ( .A1(n8151), .A2(n7845), .ZN(n5927) );
  XNOR2_X1 U7678 ( .A(n5948), .B(P1_REG3_REG_22__SCAN_IN), .ZN(n9787) );
  NAND2_X1 U7679 ( .A1(n9787), .A2(n6047), .ZN(n5934) );
  INV_X1 U7680 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7681 ( .A1(n6153), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5930) );
  NAND2_X1 U7682 ( .A1(n5894), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5929) );
  OAI211_X1 U7683 ( .C1(n5931), .C2(n5837), .A(n5930), .B(n5929), .ZN(n5932)
         );
  INV_X1 U7684 ( .A(n5932), .ZN(n5933) );
  NAND2_X1 U7685 ( .A1(n5934), .A2(n5933), .ZN(n9805) );
  NOR2_X1 U7686 ( .A1(n9960), .A2(n9805), .ZN(n5936) );
  NAND2_X1 U7687 ( .A1(n9960), .A2(n9805), .ZN(n5935) );
  OR2_X1 U7688 ( .A1(n5981), .A2(n5957), .ZN(n5937) );
  NAND2_X1 U7689 ( .A1(n5937), .A2(n5958), .ZN(n5943) );
  INV_X1 U7690 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7937) );
  INV_X1 U7691 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7933) );
  MUX2_X1 U7692 ( .A(n7937), .B(n7933), .S(n8144), .Z(n5939) );
  INV_X1 U7693 ( .A(SI_23_), .ZN(n5938) );
  NAND2_X1 U7694 ( .A1(n5939), .A2(n5938), .ZN(n5961) );
  INV_X1 U7695 ( .A(n5939), .ZN(n5940) );
  NAND2_X1 U7696 ( .A1(n5940), .A2(SI_23_), .ZN(n5941) );
  NAND2_X1 U7697 ( .A1(n5961), .A2(n5941), .ZN(n5959) );
  INV_X1 U7698 ( .A(n5959), .ZN(n5942) );
  NAND2_X1 U7699 ( .A1(n7934), .A2(n5505), .ZN(n5945) );
  OR2_X1 U7700 ( .A1(n8151), .A2(n7933), .ZN(n5944) );
  INV_X1 U7701 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9230) );
  INV_X1 U7702 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5946) );
  OAI21_X1 U7703 ( .B1(n5948), .B2(n9230), .A(n5946), .ZN(n5949) );
  NAND2_X1 U7704 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n5947) );
  NAND2_X1 U7705 ( .A1(n5949), .A2(n5971), .ZN(n9777) );
  OR2_X1 U7706 ( .A1(n9777), .A2(n6094), .ZN(n5954) );
  INV_X1 U7707 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U7708 ( .A1(n6153), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U7709 ( .A1(n5894), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5950) );
  OAI211_X1 U7710 ( .C1(n9775), .C2(n5837), .A(n5951), .B(n5950), .ZN(n5952)
         );
  INV_X1 U7711 ( .A(n5952), .ZN(n5953) );
  NAND2_X1 U7712 ( .A1(n5954), .A2(n5953), .ZN(n9796) );
  AND2_X1 U7713 ( .A1(n9957), .A2(n9796), .ZN(n5956) );
  OR2_X1 U7714 ( .A1(n9957), .A2(n9796), .ZN(n5955) );
  OR2_X1 U7715 ( .A1(n5981), .A2(n5982), .ZN(n5962) );
  OR2_X1 U7716 ( .A1(n5959), .A2(n5958), .ZN(n5960) );
  MUX2_X1 U7717 ( .A(n8054), .B(n10550), .S(n8144), .Z(n5964) );
  INV_X1 U7718 ( .A(SI_24_), .ZN(n5963) );
  INV_X1 U7719 ( .A(n5964), .ZN(n5965) );
  NAND2_X1 U7720 ( .A1(n5965), .A2(SI_24_), .ZN(n5966) );
  NAND2_X1 U7721 ( .A1(n5986), .A2(n5966), .ZN(n5984) );
  INV_X1 U7722 ( .A(n5984), .ZN(n5967) );
  NAND2_X1 U7723 ( .A1(n7998), .A2(n5505), .ZN(n5970) );
  OR2_X1 U7724 ( .A1(n8151), .A2(n10550), .ZN(n5969) );
  INV_X1 U7725 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n10521) );
  NAND2_X1 U7726 ( .A1(n5971), .A2(n10521), .ZN(n5972) );
  AND2_X1 U7727 ( .A1(n5995), .A2(n5972), .ZN(n9758) );
  NAND2_X1 U7728 ( .A1(n9758), .A2(n5517), .ZN(n5978) );
  INV_X1 U7729 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U7730 ( .A1(n6153), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U7731 ( .A1(n5894), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5973) );
  OAI211_X1 U7732 ( .C1(n5975), .C2(n5837), .A(n5974), .B(n5973), .ZN(n5976)
         );
  INV_X1 U7733 ( .A(n5976), .ZN(n5977) );
  NAND2_X1 U7734 ( .A1(n9950), .A2(n9771), .ZN(n9491) );
  NAND2_X1 U7735 ( .A1(n9950), .A2(n9549), .ZN(n5980) );
  INV_X1 U7736 ( .A(n5981), .ZN(n5985) );
  INV_X1 U7737 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8121) );
  INV_X1 U7738 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8052) );
  MUX2_X1 U7739 ( .A(n8121), .B(n8052), .S(n8144), .Z(n5988) );
  INV_X1 U7740 ( .A(SI_25_), .ZN(n5987) );
  NAND2_X1 U7741 ( .A1(n5988), .A2(n5987), .ZN(n6007) );
  INV_X1 U7742 ( .A(n5988), .ZN(n5989) );
  NAND2_X1 U7743 ( .A1(n5989), .A2(SI_25_), .ZN(n5990) );
  XNOR2_X1 U7744 ( .A(n6006), .B(n6005), .ZN(n8051) );
  NAND2_X1 U7745 ( .A1(n8051), .A2(n5505), .ZN(n5992) );
  OR2_X1 U7746 ( .A1(n8151), .A2(n8052), .ZN(n5991) );
  INV_X1 U7747 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U7748 ( .A1(n5995), .A2(n5994), .ZN(n5996) );
  AND2_X1 U7749 ( .A1(n6016), .A2(n5996), .ZN(n9742) );
  NAND2_X1 U7750 ( .A1(n9742), .A2(n6047), .ZN(n6002) );
  INV_X1 U7751 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U7752 ( .A1(n6153), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7753 ( .A1(n5894), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5997) );
  OAI211_X1 U7754 ( .C1(n5999), .C2(n5837), .A(n5998), .B(n5997), .ZN(n6000)
         );
  INV_X1 U7755 ( .A(n6000), .ZN(n6001) );
  OR2_X1 U7756 ( .A1(n9741), .A2(n9750), .ZN(n6003) );
  NAND2_X1 U7757 ( .A1(n9741), .A2(n9750), .ZN(n6004) );
  INV_X1 U7758 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8069) );
  MUX2_X1 U7759 ( .A(n10474), .B(n8069), .S(n8144), .Z(n6009) );
  INV_X1 U7760 ( .A(SI_26_), .ZN(n6008) );
  NAND2_X1 U7761 ( .A1(n6009), .A2(n6008), .ZN(n6025) );
  INV_X1 U7762 ( .A(n6009), .ZN(n6010) );
  NAND2_X1 U7763 ( .A1(n6010), .A2(SI_26_), .ZN(n6011) );
  XNOR2_X1 U7764 ( .A(n6024), .B(n6023), .ZN(n8067) );
  NAND2_X1 U7765 ( .A1(n8067), .A2(n5505), .ZN(n6013) );
  OR2_X1 U7766 ( .A1(n8151), .A2(n8069), .ZN(n6012) );
  INV_X1 U7767 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7768 ( .A1(n6016), .A2(n6015), .ZN(n6017) );
  NAND2_X1 U7769 ( .A1(n6045), .A2(n6017), .ZN(n9725) );
  INV_X1 U7770 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9724) );
  NAND2_X1 U7771 ( .A1(n6153), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7772 ( .A1(n5894), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6018) );
  OAI211_X1 U7773 ( .C1(n9724), .C2(n5837), .A(n6019), .B(n6018), .ZN(n6020)
         );
  INV_X1 U7774 ( .A(n6020), .ZN(n6021) );
  OR2_X1 U7775 ( .A1(n9723), .A2(n9736), .ZN(n9385) );
  NAND2_X1 U7776 ( .A1(n9723), .A2(n9736), .ZN(n9700) );
  NAND2_X1 U7777 ( .A1(n9385), .A2(n9700), .ZN(n9721) );
  NAND2_X1 U7778 ( .A1(n6024), .A2(n6023), .ZN(n6026) );
  INV_X1 U7779 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6467) );
  INV_X1 U7780 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10059) );
  MUX2_X1 U7781 ( .A(n6467), .B(n10059), .S(n8144), .Z(n6027) );
  INV_X1 U7782 ( .A(SI_27_), .ZN(n10533) );
  NAND2_X1 U7783 ( .A1(n6027), .A2(n10533), .ZN(n6039) );
  INV_X1 U7784 ( .A(n6027), .ZN(n6028) );
  NAND2_X1 U7785 ( .A1(n6028), .A2(SI_27_), .ZN(n6029) );
  NAND2_X1 U7786 ( .A1(n9086), .A2(n5505), .ZN(n6031) );
  OR2_X1 U7787 ( .A1(n8151), .A2(n10059), .ZN(n6030) );
  XNOR2_X1 U7788 ( .A(n6045), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9708) );
  INV_X1 U7789 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7790 ( .A1(n6153), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U7791 ( .A1(n5894), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6032) );
  OAI211_X1 U7792 ( .C1(n6034), .C2(n5837), .A(n6033), .B(n6032), .ZN(n6035)
         );
  NAND2_X1 U7793 ( .A1(n8118), .A2(n9718), .ZN(n9379) );
  INV_X1 U7794 ( .A(n9718), .ZN(n9547) );
  OR2_X1 U7795 ( .A1(n8118), .A2(n9547), .ZN(n6036) );
  INV_X1 U7796 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6481) );
  INV_X1 U7797 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8250) );
  MUX2_X1 U7798 ( .A(n6481), .B(n8250), .S(n8144), .Z(n6140) );
  XNOR2_X1 U7799 ( .A(n6140), .B(SI_28_), .ZN(n6137) );
  NAND2_X1 U7800 ( .A1(n6480), .A2(n5505), .ZN(n6042) );
  OR2_X1 U7801 ( .A1(n8151), .A2(n8250), .ZN(n6041) );
  INV_X1 U7802 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8114) );
  INV_X1 U7803 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6043) );
  OAI21_X1 U7804 ( .B1(n6045), .B2(n8114), .A(n6043), .ZN(n6046) );
  NAND2_X1 U7805 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6044) );
  NAND2_X1 U7806 ( .A1(n8242), .A2(n6047), .ZN(n6053) );
  INV_X1 U7807 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7808 ( .A1(n6153), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7809 ( .A1(n5894), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6048) );
  OAI211_X1 U7810 ( .C1(n6050), .C2(n5837), .A(n6049), .B(n6048), .ZN(n6051)
         );
  INV_X1 U7811 ( .A(n6051), .ZN(n6052) );
  AND2_X2 U7812 ( .A1(n6053), .A2(n6052), .ZN(n9703) );
  OR2_X2 U7813 ( .A1(n6873), .A2(n9703), .ZN(n9501) );
  NAND2_X1 U7814 ( .A1(n6873), .A2(n9703), .ZN(n9380) );
  OR2_X2 U7815 ( .A1(n6054), .A2(n9403), .ZN(n9688) );
  NAND2_X1 U7816 ( .A1(n6054), .A2(n9403), .ZN(n6055) );
  NAND2_X1 U7817 ( .A1(n6057), .A2(n6056), .ZN(n6063) );
  INV_X1 U7818 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7819 ( .A1(n6066), .A2(n6058), .ZN(n6059) );
  NAND2_X1 U7820 ( .A1(n6068), .A2(n6594), .ZN(n6600) );
  NAND2_X1 U7821 ( .A1(n6063), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6065) );
  AND2_X1 U7822 ( .A1(n6600), .A2(n9534), .ZN(n6070) );
  INV_X1 U7823 ( .A(n6068), .ZN(n7843) );
  INV_X1 U7824 ( .A(n9447), .ZN(n7674) );
  INV_X1 U7825 ( .A(n7337), .ZN(n6069) );
  OAI21_X1 U7826 ( .B1(n9529), .B2(n9534), .A(n6069), .ZN(n7737) );
  NAND2_X1 U7827 ( .A1(n9394), .A2(n6592), .ZN(n10151) );
  NOR2_X1 U7828 ( .A1(n7808), .A2(n7816), .ZN(n7810) );
  NAND2_X1 U7829 ( .A1(n9448), .A2(n6601), .ZN(n6071) );
  NAND2_X1 U7830 ( .A1(n6073), .A2(n4573), .ZN(n7771) );
  AND2_X1 U7831 ( .A1(n9323), .A2(n9293), .ZN(n6075) );
  XNOR2_X1 U7832 ( .A(n9326), .B(n9552), .ZN(n9422) );
  NAND2_X1 U7833 ( .A1(n7722), .A2(n9422), .ZN(n6077) );
  INV_X1 U7834 ( .A(n9552), .ZN(n9325) );
  NAND2_X1 U7835 ( .A1(n9326), .A2(n9325), .ZN(n9348) );
  INV_X1 U7836 ( .A(n9349), .ZN(n9909) );
  NOR2_X1 U7837 ( .A1(n9925), .A2(n9909), .ZN(n6078) );
  OR2_X2 U7838 ( .A1(n10003), .A2(n9280), .ZN(n9467) );
  NAND2_X1 U7839 ( .A1(n10003), .A2(n9280), .ZN(n9350) );
  NAND2_X1 U7840 ( .A1(n9467), .A2(n9350), .ZN(n9895) );
  OR2_X1 U7841 ( .A1(n9998), .A2(n9897), .ZN(n9471) );
  NAND2_X1 U7842 ( .A1(n9998), .A2(n9897), .ZN(n9351) );
  NAND2_X1 U7843 ( .A1(n9471), .A2(n9351), .ZN(n9426) );
  INV_X1 U7844 ( .A(n9467), .ZN(n8233) );
  NOR2_X1 U7845 ( .A1(n9426), .A2(n8233), .ZN(n6079) );
  INV_X1 U7846 ( .A(n6080), .ZN(n9475) );
  INV_X1 U7847 ( .A(n9867), .ZN(n9855) );
  NAND2_X1 U7848 ( .A1(n9988), .A2(n9855), .ZN(n9480) );
  INV_X1 U7849 ( .A(n9835), .ZN(n9178) );
  OR2_X1 U7850 ( .A1(n9983), .A2(n9178), .ZN(n9353) );
  NAND2_X1 U7851 ( .A1(n9983), .A2(n9178), .ZN(n9479) );
  NAND2_X1 U7852 ( .A1(n9353), .A2(n9479), .ZN(n9860) );
  INV_X1 U7853 ( .A(n9820), .ZN(n9856) );
  OR2_X1 U7854 ( .A1(n9975), .A2(n9856), .ZN(n9335) );
  NAND2_X1 U7855 ( .A1(n9975), .A2(n9856), .ZN(n9487) );
  INV_X1 U7856 ( .A(n9821), .ZN(n9233) );
  OR2_X1 U7857 ( .A1(n9966), .A2(n9233), .ZN(n9405) );
  INV_X1 U7858 ( .A(n9836), .ZN(n9124) );
  AND2_X1 U7859 ( .A1(n9405), .A2(n9802), .ZN(n9440) );
  INV_X1 U7860 ( .A(n9805), .ZN(n9770) );
  OR2_X1 U7861 ( .A1(n9960), .A2(n9770), .ZN(n9764) );
  NAND2_X1 U7862 ( .A1(n9960), .A2(n9770), .ZN(n9367) );
  NAND2_X1 U7863 ( .A1(n9764), .A2(n9367), .ZN(n9791) );
  NAND2_X1 U7864 ( .A1(n9966), .A2(n9233), .ZN(n9404) );
  NAND2_X1 U7865 ( .A1(n9971), .A2(n9124), .ZN(n9406) );
  NAND2_X1 U7866 ( .A1(n9404), .A2(n9406), .ZN(n9289) );
  AND2_X1 U7867 ( .A1(n9289), .A2(n9405), .ZN(n9792) );
  NOR2_X1 U7868 ( .A1(n9791), .A2(n9792), .ZN(n6082) );
  INV_X1 U7869 ( .A(n9796), .ZN(n9231) );
  NAND2_X1 U7870 ( .A1(n9957), .A2(n9231), .ZN(n9748) );
  NAND2_X1 U7871 ( .A1(n9369), .A2(n9748), .ZN(n9768) );
  INV_X1 U7872 ( .A(n9764), .ZN(n6083) );
  NOR2_X1 U7873 ( .A1(n9768), .A2(n6083), .ZN(n6084) );
  INV_X1 U7874 ( .A(n9748), .ZN(n9370) );
  NOR2_X1 U7875 ( .A1(n5979), .A2(n9370), .ZN(n6085) );
  NAND2_X1 U7876 ( .A1(n9765), .A2(n6085), .ZN(n6086) );
  NAND2_X1 U7877 ( .A1(n9741), .A2(n9717), .ZN(n9492) );
  INV_X1 U7878 ( .A(n9700), .ZN(n9387) );
  NOR2_X1 U7879 ( .A1(n9698), .A2(n9387), .ZN(n6087) );
  NAND2_X1 U7880 ( .A1(n9716), .A2(n6087), .ZN(n6088) );
  NAND2_X1 U7881 ( .A1(n6068), .A2(n9511), .ZN(n9402) );
  INV_X1 U7882 ( .A(n6592), .ZN(n9527) );
  NAND2_X1 U7883 ( .A1(n9447), .A2(n9527), .ZN(n9399) );
  OAI211_X1 U7884 ( .C1(n6089), .C2(n9403), .A(n6152), .B(n9918), .ZN(n6096)
         );
  INV_X1 U7885 ( .A(n4437), .ZN(n7030) );
  INV_X1 U7886 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9692) );
  NAND2_X1 U7887 ( .A1(n5894), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7888 ( .A1(n6153), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6090) );
  OAI211_X1 U7889 ( .C1(n9692), .C2(n5837), .A(n6091), .B(n6090), .ZN(n6092)
         );
  INV_X1 U7890 ( .A(n6092), .ZN(n6093) );
  OAI21_X1 U7891 ( .B1(n9693), .B2(n6094), .A(n6093), .ZN(n9545) );
  AOI22_X1 U7892 ( .A1(n9547), .A2(n9915), .B1(n9545), .B2(n9913), .ZN(n6095)
         );
  NAND2_X1 U7893 ( .A1(n6096), .A2(n6095), .ZN(n8247) );
  NAND2_X1 U7894 ( .A1(n7378), .A2(n7816), .ZN(n7815) );
  INV_X1 U7895 ( .A(n9113), .ZN(n7709) );
  AND2_X2 U7896 ( .A1(n7707), .A2(n7709), .ZN(n7706) );
  OR2_X1 U7897 ( .A1(n10008), .A2(n9145), .ZN(n6099) );
  INV_X1 U7898 ( .A(n9998), .ZN(n9288) );
  INV_X1 U7899 ( .A(n9960), .ZN(n9789) );
  INV_X1 U7900 ( .A(n6103), .ZN(n9707) );
  AND2_X1 U7901 ( .A1(n7337), .A2(n6592), .ZN(n9976) );
  AOI21_X1 U7902 ( .B1(n9707), .B2(n6873), .A(n9907), .ZN(n6104) );
  AND2_X1 U7903 ( .A1(n6147), .A2(n6104), .ZN(n8241) );
  NAND2_X1 U7904 ( .A1(n6105), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6107) );
  INV_X1 U7905 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6106) );
  INV_X1 U7906 ( .A(n6108), .ZN(n6109) );
  NAND2_X1 U7907 ( .A1(n6109), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6110) );
  XNOR2_X1 U7908 ( .A(n6113), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6118) );
  XNOR2_X1 U7909 ( .A(n6115), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6117) );
  OAI211_X1 U7910 ( .C1(n9529), .C2(n6595), .A(n7029), .B(n6908), .ZN(n6860)
         );
  INV_X1 U7911 ( .A(n6117), .ZN(n8053) );
  NAND2_X1 U7912 ( .A1(n8053), .A2(P1_B_REG_SCAN_IN), .ZN(n6119) );
  MUX2_X1 U7913 ( .A(n6119), .B(P1_B_REG_SCAN_IN), .S(n6118), .Z(n6120) );
  NOR4_X1 U7914 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6121) );
  INV_X1 U7915 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10518) );
  INV_X1 U7916 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10522) );
  NAND3_X1 U7917 ( .A1(n6121), .A2(n10518), .A3(n10522), .ZN(n6127) );
  NOR4_X1 U7918 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n6125) );
  NOR4_X1 U7919 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6124) );
  NOR4_X1 U7920 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6123) );
  NOR4_X1 U7921 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6122) );
  NAND4_X1 U7922 ( .A1(n6125), .A2(n6124), .A3(n6123), .A4(n6122), .ZN(n6126)
         );
  NOR4_X1 U7923 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        n6127), .A4(n6126), .ZN(n6129) );
  INV_X1 U7924 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10486) );
  INV_X1 U7925 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10345) );
  INV_X1 U7926 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10358) );
  INV_X1 U7927 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10365) );
  NAND4_X1 U7928 ( .A1(n10486), .A2(n10345), .A3(n10358), .A4(n10365), .ZN(
        n6128) );
  NOR3_X1 U7929 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6128), .ZN(n10284) );
  AND2_X1 U7930 ( .A1(n6129), .A2(n10284), .ZN(n6130) );
  NAND2_X1 U7931 ( .A1(n6848), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7932 ( .A1(n9976), .A2(n9511), .ZN(n6857) );
  OR2_X1 U7933 ( .A1(n10040), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6133) );
  INV_X1 U7934 ( .A(n6132), .ZN(n8071) );
  NAND2_X1 U7935 ( .A1(n8071), .A2(n8053), .ZN(n10268) );
  NAND2_X1 U7936 ( .A1(n6133), .A2(n10268), .ZN(n7731) );
  NAND2_X1 U7937 ( .A1(n6857), .A2(n7731), .ZN(n6134) );
  INV_X1 U7938 ( .A(n6118), .ZN(n7999) );
  NAND2_X1 U7939 ( .A1(n7999), .A2(n8071), .ZN(n10042) );
  NAND2_X1 U7940 ( .A1(n10159), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6136) );
  INV_X1 U7941 ( .A(SI_28_), .ZN(n6139) );
  NAND2_X1 U7942 ( .A1(n6140), .A2(n6139), .ZN(n6141) );
  INV_X1 U7943 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8111) );
  INV_X1 U7944 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10428) );
  MUX2_X1 U7945 ( .A(n8111), .B(n10428), .S(n8144), .Z(n8135) );
  XNOR2_X2 U7946 ( .A(n8136), .B(n8135), .ZN(n8138) );
  NAND2_X1 U7947 ( .A1(n8109), .A2(n5505), .ZN(n6144) );
  OR2_X1 U7948 ( .A1(n8151), .A2(n10428), .ZN(n6143) );
  INV_X1 U7949 ( .A(n9545), .ZN(n6145) );
  NAND2_X1 U7950 ( .A1(n6163), .A2(n6145), .ZN(n9504) );
  INV_X1 U7951 ( .A(n9703), .ZN(n9546) );
  NAND2_X1 U7952 ( .A1(n6873), .A2(n9546), .ZN(n9687) );
  INV_X1 U7953 ( .A(n9688), .ZN(n6151) );
  INV_X1 U7954 ( .A(n9696), .ZN(n6148) );
  NAND2_X1 U7955 ( .A1(n6148), .A2(n5229), .ZN(n6149) );
  INV_X1 U7956 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U7957 ( .A1(n5894), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7958 ( .A1(n6153), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6154) );
  OAI211_X1 U7959 ( .C1(n5837), .C2(n6156), .A(n6155), .B(n6154), .ZN(n9544)
         );
  INV_X1 U7960 ( .A(n9544), .ZN(n9435) );
  INV_X1 U7961 ( .A(n6158), .ZN(n9535) );
  NAND2_X1 U7962 ( .A1(n9535), .A2(P1_B_REG_SCAN_IN), .ZN(n6159) );
  NAND2_X1 U7963 ( .A1(n9913), .A2(n6159), .ZN(n8156) );
  OAI22_X1 U7964 ( .A1(n9703), .A2(n9898), .B1(n9435), .B2(n8156), .ZN(n6160)
         );
  INV_X1 U7965 ( .A(n6163), .ZN(n9691) );
  NAND2_X1 U7966 ( .A1(n10159), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6164) );
  INV_X1 U7967 ( .A(n7732), .ZN(n6165) );
  NAND2_X1 U7968 ( .A1(n10154), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6167) );
  XNOR2_X2 U7969 ( .A(n6171), .B(n9076), .ZN(n8240) );
  INV_X1 U7970 ( .A(n8240), .ZN(n6173) );
  INV_X1 U7971 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6997) );
  OR2_X1 U7972 ( .A1(n6223), .A2(n6997), .ZN(n6179) );
  NAND2_X1 U7973 ( .A1(n6222), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6178) );
  OR2_X2 U7974 ( .A1(n8240), .A2(n6175), .ZN(n6225) );
  OR2_X1 U7975 ( .A1(n6225), .A2(n7249), .ZN(n6177) );
  NAND2_X1 U7977 ( .A1(n6183), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7978 ( .A1(n6200), .A2(n6936), .ZN(n6182) );
  OR2_X1 U7979 ( .A1(n6547), .A2(n6180), .ZN(n6181) );
  OAI211_X1 U7980 ( .C1(n6370), .C2(P1_DATAO_REG_1__SCAN_IN), .A(n6182), .B(
        n6181), .ZN(n7239) );
  OR2_X1 U7981 ( .A1(n8620), .A2(n6191), .ZN(n6195) );
  INV_X1 U7982 ( .A(n7969), .ZN(n6183) );
  NAND2_X1 U7983 ( .A1(n6222), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6188) );
  INV_X1 U7984 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6184) );
  OR2_X1 U7985 ( .A1(n6223), .A2(n6184), .ZN(n6187) );
  OR2_X1 U7986 ( .A1(n6225), .A2(n6185), .ZN(n6186) );
  NOR2_X1 U7987 ( .A1(n8144), .A2(n10538), .ZN(n6190) );
  XNOR2_X1 U7988 ( .A(n6190), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9091) );
  MUX2_X1 U7989 ( .A(n4436), .B(n9091), .S(n6547), .Z(n7141) );
  INV_X1 U7990 ( .A(n7141), .ZN(n10188) );
  NAND2_X1 U7991 ( .A1(n8621), .A2(n10188), .ZN(n7245) );
  INV_X1 U7992 ( .A(n6193), .ZN(n6192) );
  NAND2_X1 U7993 ( .A1(n8460), .A2(n8455), .ZN(n7244) );
  NAND2_X1 U7994 ( .A1(n7245), .A2(n7244), .ZN(n6194) );
  NAND2_X1 U7995 ( .A1(n6195), .A2(n6194), .ZN(n7165) );
  NAND2_X1 U7996 ( .A1(n6222), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6198) );
  INV_X1 U7997 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7172) );
  AND3_X1 U7998 ( .A1(n6198), .A2(n6197), .A3(n6196), .ZN(n6199) );
  INV_X1 U7999 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10234) );
  INV_X1 U8000 ( .A(n6207), .ZN(n6205) );
  OR2_X1 U8001 ( .A1(n6947), .A2(n6287), .ZN(n6203) );
  OR2_X1 U8002 ( .A1(n6370), .A2(n6926), .ZN(n6202) );
  OR2_X1 U8003 ( .A1(n6547), .A2(n6994), .ZN(n6201) );
  NAND2_X1 U8004 ( .A1(n6205), .A2(n6204), .ZN(n6507) );
  NAND2_X1 U8005 ( .A1(n6208), .A2(n6207), .ZN(n8462) );
  INV_X1 U8006 ( .A(n8461), .ZN(n6206) );
  NAND2_X1 U8007 ( .A1(n7165), .A2(n6206), .ZN(n6210) );
  OR2_X1 U8008 ( .A1(n8619), .A2(n6204), .ZN(n6209) );
  NAND2_X1 U8009 ( .A1(n6210), .A2(n6209), .ZN(n7357) );
  INV_X1 U8010 ( .A(n7357), .ZN(n6218) );
  INV_X2 U8011 ( .A(n6225), .ZN(n6541) );
  INV_X1 U8012 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6211) );
  OR2_X1 U8013 ( .A1(n6223), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6213) );
  INV_X1 U8014 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10236) );
  OR2_X1 U8015 ( .A1(n7969), .A2(n10236), .ZN(n6212) );
  OR2_X1 U8016 ( .A1(n6942), .A2(n6287), .ZN(n6217) );
  INV_X2 U8017 ( .A(n6370), .ZN(n6389) );
  INV_X2 U8018 ( .A(n6547), .ZN(n6388) );
  AOI22_X1 U8019 ( .A1(n6389), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n6388), .B2(
        n7159), .ZN(n6216) );
  INV_X1 U8020 ( .A(n10201), .ZN(n7360) );
  NAND2_X1 U8021 ( .A1(n6218), .A2(n5213), .ZN(n7430) );
  OR2_X1 U8022 ( .A1(n6943), .A2(n6287), .ZN(n6221) );
  AOI22_X1 U8023 ( .A1(n6389), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n6388), .B2(
        n6219), .ZN(n6220) );
  NAND2_X1 U8024 ( .A1(n6221), .A2(n6220), .ZN(n7309) );
  INV_X1 U8025 ( .A(n7309), .ZN(n10205) );
  NAND2_X1 U8026 ( .A1(n7967), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6230) );
  OR2_X1 U8027 ( .A1(n7969), .A2(n10238), .ZN(n6229) );
  NAND2_X1 U8028 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6224) );
  AND2_X1 U8029 ( .A1(n6233), .A2(n6224), .ZN(n7428) );
  OR2_X1 U8030 ( .A1(n6312), .A2(n7428), .ZN(n6228) );
  OR2_X1 U8031 ( .A1(n7973), .A2(n6226), .ZN(n6227) );
  NAND2_X1 U8032 ( .A1(n10205), .A2(n7255), .ZN(n8468) );
  NAND2_X1 U8033 ( .A1(n7302), .A2(n7309), .ZN(n8486) );
  NAND2_X1 U8034 ( .A1(n8468), .A2(n8486), .ZN(n7432) );
  NAND2_X1 U8035 ( .A1(n6508), .A2(n7360), .ZN(n7429) );
  AND2_X1 U8036 ( .A1(n7432), .A2(n7429), .ZN(n6231) );
  NAND2_X1 U8037 ( .A1(n7302), .A2(n10205), .ZN(n10163) );
  NAND2_X1 U8038 ( .A1(n7967), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6238) );
  OR2_X1 U8039 ( .A1(n7973), .A2(n4919), .ZN(n6237) );
  INV_X1 U8040 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10240) );
  OR2_X1 U8041 ( .A1(n7969), .A2(n10240), .ZN(n6236) );
  NAND2_X1 U8042 ( .A1(n6233), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6234) );
  AND2_X1 U8043 ( .A1(n6245), .A2(n6234), .ZN(n10174) );
  OR2_X1 U8044 ( .A1(n6312), .A2(n10174), .ZN(n6235) );
  NAND4_X1 U8045 ( .A1(n6238), .A2(n6237), .A3(n6236), .A4(n6235), .ZN(n8618)
         );
  OR2_X1 U8046 ( .A1(n6239), .A2(n6287), .ZN(n6241) );
  AOI22_X1 U8047 ( .A1(n6389), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6388), .B2(
        n5320), .ZN(n6240) );
  NAND2_X1 U8048 ( .A1(n6241), .A2(n6240), .ZN(n10179) );
  NAND2_X1 U8049 ( .A1(n7421), .A2(n10179), .ZN(n8487) );
  NAND2_X1 U8050 ( .A1(n10211), .A2(n8618), .ZN(n8490) );
  NAND2_X1 U8051 ( .A1(n8487), .A2(n8490), .ZN(n8415) );
  INV_X2 U8052 ( .A(n6287), .ZN(n8402) );
  NAND2_X1 U8053 ( .A1(n6934), .A2(n8402), .ZN(n6244) );
  AOI22_X1 U8054 ( .A1(n6389), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6388), .B2(
        n6242), .ZN(n6243) );
  NAND2_X1 U8055 ( .A1(n6244), .A2(n6243), .ZN(n7461) );
  NAND2_X1 U8056 ( .A1(n7967), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6250) );
  OR2_X1 U8057 ( .A1(n7969), .A2(n10242), .ZN(n6249) );
  NAND2_X1 U8058 ( .A1(n6245), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6246) );
  AND2_X1 U8059 ( .A1(n6258), .A2(n6246), .ZN(n7459) );
  OR2_X1 U8060 ( .A1(n6312), .A2(n7459), .ZN(n6248) );
  OR2_X1 U8061 ( .A1(n7973), .A2(n7458), .ZN(n6247) );
  INV_X1 U8062 ( .A(n7555), .ZN(n10169) );
  NAND2_X1 U8063 ( .A1(n7461), .A2(n10169), .ZN(n6251) );
  OR2_X1 U8064 ( .A1(n7461), .A2(n10169), .ZN(n6252) );
  OR2_X1 U8065 ( .A1(n6932), .A2(n6287), .ZN(n6255) );
  AOI22_X1 U8066 ( .A1(n6389), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6388), .B2(
        n6253), .ZN(n6254) );
  NAND2_X1 U8067 ( .A1(n6541), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6264) );
  OR2_X1 U8068 ( .A1(n7969), .A2(n7563), .ZN(n6263) );
  NAND2_X1 U8069 ( .A1(n6258), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6259) );
  AND2_X1 U8070 ( .A1(n6278), .A2(n6259), .ZN(n7565) );
  OR2_X1 U8071 ( .A1(n6312), .A2(n7565), .ZN(n6262) );
  INV_X1 U8072 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6260) );
  OR2_X1 U8073 ( .A1(n6544), .A2(n6260), .ZN(n6261) );
  NAND2_X1 U8074 ( .A1(n7566), .A2(n8617), .ZN(n7597) );
  INV_X1 U8075 ( .A(n7566), .ZN(n6265) );
  NAND2_X1 U8076 ( .A1(n6265), .A2(n7592), .ZN(n8476) );
  INV_X1 U8077 ( .A(n8416), .ZN(n8474) );
  NAND2_X1 U8078 ( .A1(n7566), .A2(n7592), .ZN(n6266) );
  NAND2_X1 U8079 ( .A1(n6958), .A2(n8402), .ZN(n6268) );
  AOI22_X1 U8080 ( .A1(n6389), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7540), .B2(
        n6388), .ZN(n6267) );
  NAND2_X1 U8081 ( .A1(n7967), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6273) );
  OR2_X1 U8082 ( .A1(n7969), .A2(n10500), .ZN(n6272) );
  NAND2_X1 U8083 ( .A1(n6280), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6269) );
  AND2_X1 U8084 ( .A1(n6290), .A2(n6269), .ZN(n7680) );
  OR2_X1 U8085 ( .A1(n6312), .A2(n7680), .ZN(n6271) );
  OR2_X1 U8086 ( .A1(n7973), .A2(n7679), .ZN(n6270) );
  NAND2_X1 U8087 ( .A1(n7859), .A2(n7850), .ZN(n8481) );
  NAND2_X1 U8088 ( .A1(n8494), .A2(n8481), .ZN(n8422) );
  NAND2_X1 U8089 ( .A1(n6937), .A2(n8402), .ZN(n6276) );
  AOI22_X1 U8090 ( .A1(n6389), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6388), .B2(
        n6274), .ZN(n6275) );
  INV_X1 U8091 ( .A(n7628), .ZN(n10224) );
  NAND2_X1 U8092 ( .A1(n6474), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6284) );
  INV_X1 U8093 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6277) );
  OR2_X1 U8094 ( .A1(n6544), .A2(n6277), .ZN(n6283) );
  NAND2_X1 U8095 ( .A1(n6278), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6279) );
  AND2_X1 U8096 ( .A1(n6280), .A2(n6279), .ZN(n7603) );
  OR2_X1 U8097 ( .A1(n6312), .A2(n7603), .ZN(n6282) );
  OR2_X1 U8098 ( .A1(n7973), .A2(n7602), .ZN(n6281) );
  NAND2_X1 U8099 ( .A1(n7600), .A2(n5209), .ZN(n7686) );
  INV_X1 U8100 ( .A(n7851), .ZN(n8616) );
  NOR2_X1 U8101 ( .A1(n7628), .A2(n8616), .ZN(n6286) );
  INV_X1 U8102 ( .A(n7850), .ZN(n8615) );
  NOR2_X1 U8103 ( .A1(n4644), .A2(n8615), .ZN(n6285) );
  AOI21_X1 U8104 ( .B1(n8422), .B2(n6286), .A(n6285), .ZN(n7685) );
  OR2_X1 U8105 ( .A1(n6956), .A2(n6287), .ZN(n6289) );
  AOI22_X1 U8106 ( .A1(n8637), .A2(n6388), .B1(n6389), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U8107 ( .A1(n7967), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6295) );
  OR2_X1 U8108 ( .A1(n7969), .A2(n10545), .ZN(n6294) );
  NAND2_X1 U8109 ( .A1(n6290), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6291) );
  AND2_X1 U8110 ( .A1(n6301), .A2(n6291), .ZN(n8165) );
  OR2_X1 U8111 ( .A1(n6312), .A2(n8165), .ZN(n6293) );
  OR2_X1 U8112 ( .A1(n7973), .A2(n8164), .ZN(n6292) );
  NAND4_X1 U8113 ( .A1(n6295), .A2(n6294), .A3(n6293), .A4(n6292), .ZN(n8614)
         );
  OR2_X1 U8114 ( .A1(n8167), .A2(n8614), .ZN(n6296) );
  AND2_X1 U8115 ( .A1(n7685), .A2(n6296), .ZN(n6297) );
  INV_X1 U8116 ( .A(n7698), .ZN(n6308) );
  NAND2_X1 U8117 ( .A1(n6963), .A2(n8402), .ZN(n6299) );
  AOI22_X1 U8118 ( .A1(n7881), .A2(n6388), .B1(n6389), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n6298) );
  NAND2_X1 U8119 ( .A1(n6541), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6307) );
  OR2_X1 U8120 ( .A1(n7969), .A2(n10547), .ZN(n6306) );
  INV_X1 U8121 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n6300) );
  OR2_X1 U8122 ( .A1(n6544), .A2(n6300), .ZN(n6305) );
  NAND2_X1 U8123 ( .A1(n6301), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U8124 ( .A1(n6314), .A2(n6302), .ZN(n8365) );
  INV_X1 U8125 ( .A(n8365), .ZN(n6303) );
  OR2_X1 U8126 ( .A1(n6312), .A2(n6303), .ZN(n6304) );
  NAND4_X1 U8127 ( .A1(n6307), .A2(n6306), .A3(n6305), .A4(n6304), .ZN(n8613)
         );
  NAND2_X1 U8128 ( .A1(n8988), .A2(n8613), .ZN(n6309) );
  AOI22_X1 U8129 ( .A1(n6310), .A2(n6388), .B1(n6389), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U8130 ( .A1(n6314), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U8131 ( .A1(n6323), .A2(n6315), .ZN(n8292) );
  NAND2_X1 U8132 ( .A1(n6494), .A2(n8292), .ZN(n6319) );
  OR2_X1 U8133 ( .A1(n7973), .A2(n7803), .ZN(n6318) );
  OR2_X1 U8134 ( .A1(n7969), .A2(n10328), .ZN(n6317) );
  INV_X1 U8135 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7964) );
  OR2_X1 U8136 ( .A1(n6544), .A2(n7964), .ZN(n6316) );
  NAND4_X1 U8137 ( .A1(n6319), .A2(n6318), .A3(n6317), .A4(n6316), .ZN(n8612)
         );
  NAND2_X1 U8138 ( .A1(n7966), .A2(n8363), .ZN(n6320) );
  NAND2_X1 U8139 ( .A1(n7085), .A2(n8402), .ZN(n6322) );
  AOI22_X1 U8140 ( .A1(n8656), .A2(n6388), .B1(n6389), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n6321) );
  NAND2_X1 U8141 ( .A1(n6323), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6324) );
  NAND2_X1 U8142 ( .A1(n6334), .A2(n6324), .ZN(n7919) );
  NAND2_X1 U8143 ( .A1(n6494), .A2(n7919), .ZN(n6328) );
  OR2_X1 U8144 ( .A1(n7969), .A2(n8647), .ZN(n6327) );
  OR2_X1 U8145 ( .A1(n7973), .A2(n10350), .ZN(n6326) );
  INV_X1 U8146 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10377) );
  OR2_X1 U8147 ( .A1(n6544), .A2(n10377), .ZN(n6325) );
  NAND2_X1 U8148 ( .A1(n7913), .A2(n7801), .ZN(n8506) );
  NAND2_X1 U8149 ( .A1(n7913), .A2(n8925), .ZN(n6329) );
  NAND2_X1 U8150 ( .A1(n7909), .A2(n6329), .ZN(n8924) );
  NAND2_X1 U8151 ( .A1(n7122), .A2(n8402), .ZN(n6331) );
  AOI22_X1 U8152 ( .A1(n8671), .A2(n6388), .B1(n6389), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6330) );
  OR2_X1 U8153 ( .A1(n7973), .A2(n10356), .ZN(n6333) );
  OR2_X1 U8154 ( .A1(n7969), .A2(n8982), .ZN(n6332) );
  AND2_X1 U8155 ( .A1(n6333), .A2(n6332), .ZN(n6338) );
  NAND2_X1 U8156 ( .A1(n6334), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U8157 ( .A1(n6344), .A2(n6335), .ZN(n8931) );
  NAND2_X1 U8158 ( .A1(n8931), .A2(n6494), .ZN(n6337) );
  INV_X1 U8159 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10517) );
  OR2_X1 U8160 ( .A1(n6544), .A2(n10517), .ZN(n6336) );
  INV_X1 U8161 ( .A(n8056), .ZN(n8915) );
  OR2_X1 U8162 ( .A1(n9067), .A2(n8915), .ZN(n6339) );
  NAND2_X1 U8163 ( .A1(n9067), .A2(n8915), .ZN(n6340) );
  NAND2_X1 U8164 ( .A1(n7331), .A2(n8402), .ZN(n6342) );
  AOI22_X1 U8165 ( .A1(n8695), .A2(n6388), .B1(n6389), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6341) );
  NAND2_X1 U8166 ( .A1(n6344), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6345) );
  NAND2_X1 U8167 ( .A1(n6352), .A2(n6345), .ZN(n8919) );
  NAND2_X1 U8168 ( .A1(n8919), .A2(n6494), .ZN(n6348) );
  AOI22_X1 U8169 ( .A1(n7967), .A2(P2_REG0_REG_15__SCAN_IN), .B1(n6474), .B2(
        P2_REG1_REG_15__SCAN_IN), .ZN(n6347) );
  NAND2_X1 U8170 ( .A1(n6541), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U8171 ( .A1(n9061), .A2(n8081), .ZN(n8516) );
  NAND2_X1 U8172 ( .A1(n8515), .A2(n8516), .ZN(n8513) );
  NAND2_X1 U8173 ( .A1(n9061), .A2(n8926), .ZN(n6349) );
  NAND2_X1 U8174 ( .A1(n7372), .A2(n8402), .ZN(n6351) );
  AOI22_X1 U8175 ( .A1(n8717), .A2(n6388), .B1(n6389), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n6350) );
  NAND2_X1 U8176 ( .A1(n6352), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6353) );
  NAND2_X1 U8177 ( .A1(n6360), .A2(n6353), .ZN(n8910) );
  NAND2_X1 U8178 ( .A1(n8910), .A2(n6494), .ZN(n6356) );
  AOI22_X1 U8179 ( .A1(n6541), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n6474), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U8180 ( .A1(n7967), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U8181 ( .A1(n9055), .A2(n8313), .ZN(n8518) );
  NAND2_X1 U8182 ( .A1(n8519), .A2(n8518), .ZN(n8410) );
  NAND2_X1 U8183 ( .A1(n7328), .A2(n8402), .ZN(n6359) );
  AOI22_X1 U8184 ( .A1(n6357), .A2(n6388), .B1(n6389), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U8185 ( .A1(n6360), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6361) );
  NAND2_X1 U8186 ( .A1(n6383), .A2(n6361), .ZN(n8901) );
  NAND2_X1 U8187 ( .A1(n8901), .A2(n6494), .ZN(n6366) );
  NAND2_X1 U8188 ( .A1(n6474), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6363) );
  NAND2_X1 U8189 ( .A1(n7967), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6362) );
  OAI211_X1 U8190 ( .C1(n10471), .C2(n7973), .A(n6363), .B(n6362), .ZN(n6364)
         );
  INV_X1 U8191 ( .A(n6364), .ZN(n6365) );
  NOR2_X1 U8192 ( .A1(n9049), .A2(n8882), .ZN(n8531) );
  INV_X1 U8193 ( .A(n8531), .ZN(n6367) );
  NAND2_X1 U8194 ( .A1(n9049), .A2(n8882), .ZN(n8523) );
  NAND2_X1 U8195 ( .A1(n6367), .A2(n8523), .ZN(n8520) );
  NAND2_X1 U8196 ( .A1(n8898), .A2(n8520), .ZN(n6369) );
  NAND2_X1 U8197 ( .A1(n9049), .A2(n8907), .ZN(n6368) );
  NAND2_X1 U8198 ( .A1(n7607), .A2(n8402), .ZN(n6372) );
  INV_X1 U8199 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7608) );
  OR2_X1 U8200 ( .A1(n8403), .A2(n7608), .ZN(n6371) );
  NAND2_X2 U8201 ( .A1(n6372), .A2(n6371), .ZN(n9034) );
  INV_X1 U8202 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U8203 ( .A1(n6394), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6375) );
  NAND2_X1 U8204 ( .A1(n6405), .A2(n6375), .ZN(n8856) );
  NAND2_X1 U8205 ( .A1(n8856), .A2(n6494), .ZN(n6380) );
  INV_X1 U8206 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9033) );
  NAND2_X1 U8207 ( .A1(n6541), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6377) );
  NAND2_X1 U8208 ( .A1(n6474), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6376) );
  OAI211_X1 U8209 ( .C1(n9033), .C2(n6544), .A(n6377), .B(n6376), .ZN(n6378)
         );
  INV_X1 U8210 ( .A(n6378), .ZN(n6379) );
  OR2_X1 U8211 ( .A1(n9034), .A2(n8867), .ZN(n8535) );
  NAND2_X1 U8212 ( .A1(n9034), .A2(n8867), .ZN(n8538) );
  NAND2_X1 U8213 ( .A1(n8535), .A2(n8538), .ZN(n8849) );
  NAND2_X1 U8214 ( .A1(n7481), .A2(n8402), .ZN(n6382) );
  AOI22_X1 U8215 ( .A1(n6389), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6388), .B2(
        n8765), .ZN(n6381) );
  NAND2_X1 U8216 ( .A1(n6383), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6384) );
  NAND2_X1 U8217 ( .A1(n6392), .A2(n6384), .ZN(n8884) );
  NAND2_X1 U8218 ( .A1(n6541), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U8219 ( .A1(n7967), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6385) );
  OAI211_X1 U8220 ( .C1(n7969), .C2(n10504), .A(n6386), .B(n6385), .ZN(n6387)
         );
  NAND2_X1 U8221 ( .A1(n8969), .A2(n8870), .ZN(n8530) );
  NAND2_X1 U8222 ( .A1(n8533), .A2(n8530), .ZN(n8889) );
  NAND2_X1 U8223 ( .A1(n7500), .A2(n8402), .ZN(n6391) );
  AOI22_X1 U8224 ( .A1(n6389), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6388), .B2(
        n8596), .ZN(n6390) );
  NAND2_X2 U8225 ( .A1(n6391), .A2(n6390), .ZN(n8967) );
  NAND2_X1 U8226 ( .A1(n6392), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U8227 ( .A1(n6394), .A2(n6393), .ZN(n8871) );
  NAND2_X1 U8228 ( .A1(n8871), .A2(n6494), .ZN(n6399) );
  INV_X1 U8229 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n10505) );
  NAND2_X1 U8230 ( .A1(n7967), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6396) );
  INV_X1 U8231 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n10532) );
  OR2_X1 U8232 ( .A1(n7969), .A2(n10532), .ZN(n6395) );
  OAI211_X1 U8233 ( .C1(n7973), .C2(n10505), .A(n6396), .B(n6395), .ZN(n6397)
         );
  INV_X1 U8234 ( .A(n6397), .ZN(n6398) );
  NAND2_X1 U8235 ( .A1(n8967), .A2(n8611), .ZN(n8850) );
  NAND3_X1 U8236 ( .A1(n8849), .A2(n8889), .A3(n8850), .ZN(n6402) );
  INV_X2 U8237 ( .A(n8526), .ZN(n8846) );
  NAND2_X1 U8238 ( .A1(n8967), .A2(n8880), .ZN(n8534) );
  NAND2_X1 U8239 ( .A1(n8846), .A2(n8534), .ZN(n8865) );
  INV_X1 U8240 ( .A(n8870), .ZN(n8899) );
  OR2_X1 U8241 ( .A1(n8969), .A2(n8899), .ZN(n8862) );
  NAND2_X1 U8242 ( .A1(n8865), .A2(n8862), .ZN(n8833) );
  NAND3_X1 U8243 ( .A1(n8849), .A2(n8850), .A3(n8833), .ZN(n6400) );
  OR2_X1 U8244 ( .A1(n9034), .A2(n8838), .ZN(n8835) );
  AND2_X1 U8245 ( .A1(n6400), .A2(n8835), .ZN(n6401) );
  NAND2_X1 U8246 ( .A1(n7673), .A2(n8402), .ZN(n6404) );
  OR2_X1 U8247 ( .A1(n8403), .A2(n7675), .ZN(n6403) );
  INV_X1 U8248 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10502) );
  NAND2_X1 U8249 ( .A1(n6405), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U8250 ( .A1(n6412), .A2(n6406), .ZN(n8842) );
  INV_X1 U8251 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9027) );
  NAND2_X1 U8252 ( .A1(n6541), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6408) );
  NAND2_X1 U8253 ( .A1(n6474), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6407) );
  OAI211_X1 U8254 ( .C1(n9027), .C2(n6544), .A(n6408), .B(n6407), .ZN(n6409)
         );
  NAND2_X1 U8255 ( .A1(n9028), .A2(n8854), .ZN(n8539) );
  NAND2_X1 U8256 ( .A1(n8541), .A2(n8539), .ZN(n8834) );
  INV_X1 U8257 ( .A(n8854), .ZN(n8610) );
  OR2_X1 U8258 ( .A1(n9028), .A2(n8610), .ZN(n8821) );
  NAND2_X1 U8259 ( .A1(n7840), .A2(n8402), .ZN(n6411) );
  OR2_X1 U8260 ( .A1(n8403), .A2(n7842), .ZN(n6410) );
  NAND2_X1 U8261 ( .A1(n6412), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U8262 ( .A1(n6424), .A2(n6413), .ZN(n8829) );
  NAND2_X1 U8263 ( .A1(n8829), .A2(n6494), .ZN(n6419) );
  INV_X1 U8264 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n6416) );
  NAND2_X1 U8265 ( .A1(n6541), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6415) );
  NAND2_X1 U8266 ( .A1(n6474), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6414) );
  OAI211_X1 U8267 ( .C1(n6416), .C2(n6544), .A(n6415), .B(n6414), .ZN(n6417)
         );
  INV_X1 U8268 ( .A(n6417), .ZN(n6418) );
  NOR2_X1 U8269 ( .A1(n9023), .A2(n8543), .ZN(n6525) );
  INV_X1 U8270 ( .A(n6525), .ZN(n6420) );
  NAND2_X1 U8271 ( .A1(n9023), .A2(n8543), .ZN(n8551) );
  NAND2_X1 U8272 ( .A1(n6420), .A2(n8551), .ZN(n8542) );
  OR2_X1 U8273 ( .A1(n9023), .A2(n8839), .ZN(n6421) );
  NAND2_X1 U8274 ( .A1(n8824), .A2(n6421), .ZN(n8173) );
  NAND2_X1 U8275 ( .A1(n7934), .A2(n8402), .ZN(n6423) );
  OR2_X1 U8276 ( .A1(n8403), .A2(n7937), .ZN(n6422) );
  NAND2_X1 U8277 ( .A1(n6424), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6425) );
  NAND2_X1 U8278 ( .A1(n6436), .A2(n6425), .ZN(n8269) );
  NAND2_X1 U8279 ( .A1(n8269), .A2(n6494), .ZN(n6430) );
  INV_X1 U8280 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n10564) );
  NAND2_X1 U8281 ( .A1(n6541), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6427) );
  NAND2_X1 U8282 ( .A1(n6474), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6426) );
  OAI211_X1 U8283 ( .C1(n10564), .C2(n6544), .A(n6427), .B(n6426), .ZN(n6428)
         );
  INV_X1 U8284 ( .A(n6428), .ZN(n6429) );
  NAND2_X1 U8285 ( .A1(n8261), .A2(n8609), .ZN(n6431) );
  OR2_X1 U8286 ( .A1(n8261), .A2(n8609), .ZN(n6432) );
  NAND2_X1 U8287 ( .A1(n7998), .A2(n8402), .ZN(n6434) );
  OR2_X1 U8288 ( .A1(n8403), .A2(n8054), .ZN(n6433) );
  INV_X1 U8289 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6435) );
  NAND2_X1 U8290 ( .A1(n6436), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6437) );
  NAND2_X1 U8291 ( .A1(n8334), .A2(n6494), .ZN(n6442) );
  INV_X1 U8292 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n10520) );
  NAND2_X1 U8293 ( .A1(n6474), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U8294 ( .A1(n6541), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6438) );
  OAI211_X1 U8295 ( .C1(n10520), .C2(n6544), .A(n6439), .B(n6438), .ZN(n6440)
         );
  INV_X1 U8296 ( .A(n6440), .ZN(n6441) );
  NAND2_X1 U8297 ( .A1(n8329), .A2(n8801), .ZN(n6443) );
  NAND2_X1 U8298 ( .A1(n8051), .A2(n8402), .ZN(n6445) );
  OR2_X1 U8299 ( .A1(n8403), .A2(n8121), .ZN(n6444) );
  INV_X1 U8300 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6446) );
  NAND2_X1 U8301 ( .A1(n6448), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6449) );
  NAND2_X1 U8302 ( .A1(n6458), .A2(n6449), .ZN(n8804) );
  NAND2_X1 U8303 ( .A1(n8804), .A2(n6494), .ZN(n6454) );
  INV_X1 U8304 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9006) );
  NAND2_X1 U8305 ( .A1(n6474), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6451) );
  NAND2_X1 U8306 ( .A1(n6541), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6450) );
  OAI211_X1 U8307 ( .C1(n6544), .C2(n9006), .A(n6451), .B(n6450), .ZN(n6452)
         );
  INV_X1 U8308 ( .A(n6452), .ZN(n6453) );
  OR2_X1 U8309 ( .A1(n9007), .A2(n8608), .ZN(n6455) );
  NAND2_X1 U8310 ( .A1(n8067), .A2(n8402), .ZN(n6457) );
  OR2_X1 U8311 ( .A1(n8403), .A2(n10474), .ZN(n6456) );
  NAND2_X1 U8312 ( .A1(n6458), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U8313 ( .A1(n6472), .A2(n6459), .ZN(n8795) );
  NAND2_X1 U8314 ( .A1(n8795), .A2(n6494), .ZN(n6464) );
  INV_X1 U8315 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9000) );
  NAND2_X1 U8316 ( .A1(n6541), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6461) );
  NAND2_X1 U8317 ( .A1(n6474), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6460) );
  OAI211_X1 U8318 ( .C1(n9000), .C2(n6544), .A(n6461), .B(n6460), .ZN(n6462)
         );
  INV_X1 U8319 ( .A(n6462), .ZN(n6463) );
  NAND2_X1 U8320 ( .A1(n9001), .A2(n8802), .ZN(n6465) );
  NAND2_X1 U8321 ( .A1(n6466), .A2(n6465), .ZN(n8180) );
  NAND2_X1 U8322 ( .A1(n9086), .A2(n8402), .ZN(n6469) );
  OR2_X1 U8323 ( .A1(n8403), .A2(n6467), .ZN(n6468) );
  INV_X1 U8324 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U8325 ( .A1(n6472), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U8326 ( .A1(n6484), .A2(n6473), .ZN(n8255) );
  NAND2_X1 U8327 ( .A1(n8255), .A2(n6494), .ZN(n6479) );
  INV_X1 U8328 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8183) );
  NAND2_X1 U8329 ( .A1(n6541), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6476) );
  NAND2_X1 U8330 ( .A1(n6474), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6475) );
  OAI211_X1 U8331 ( .C1(n8183), .C2(n6544), .A(n6476), .B(n6475), .ZN(n6477)
         );
  INV_X1 U8332 ( .A(n6477), .ZN(n6478) );
  NAND2_X1 U8333 ( .A1(n8571), .A2(n8781), .ZN(n6528) );
  NAND2_X1 U8334 ( .A1(n6480), .A2(n8402), .ZN(n6483) );
  OR2_X1 U8335 ( .A1(n8403), .A2(n6481), .ZN(n6482) );
  NAND2_X1 U8336 ( .A1(n6484), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6485) );
  NAND2_X1 U8337 ( .A1(n8074), .A2(n6485), .ZN(n8784) );
  NAND2_X1 U8338 ( .A1(n8784), .A2(n6494), .ZN(n6490) );
  INV_X1 U8339 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10477) );
  NAND2_X1 U8340 ( .A1(n7967), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U8341 ( .A1(n6541), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6486) );
  OAI211_X1 U8342 ( .C1(n7969), .C2(n10477), .A(n6487), .B(n6486), .ZN(n6488)
         );
  INV_X1 U8343 ( .A(n6488), .ZN(n6489) );
  NOR2_X1 U8344 ( .A1(n8582), .A2(n8607), .ZN(n6491) );
  NAND2_X1 U8345 ( .A1(n8109), .A2(n8402), .ZN(n6493) );
  OR2_X1 U8346 ( .A1(n8403), .A2(n8111), .ZN(n6492) );
  INV_X1 U8347 ( .A(n8074), .ZN(n6495) );
  INV_X1 U8348 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10367) );
  NAND2_X1 U8349 ( .A1(n6541), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6497) );
  NAND2_X1 U8350 ( .A1(n7967), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6496) );
  OAI211_X1 U8351 ( .C1(n7969), .C2(n10367), .A(n6497), .B(n6496), .ZN(n6498)
         );
  INV_X1 U8352 ( .A(n6498), .ZN(n6499) );
  NAND2_X1 U8353 ( .A1(n6588), .A2(n8606), .ZN(n8406) );
  XNOR2_X1 U8354 ( .A(n6500), .B(n6533), .ZN(n6504) );
  INV_X1 U8355 ( .A(n8585), .ZN(n8440) );
  NAND2_X1 U8356 ( .A1(n6530), .A2(n8440), .ZN(n6503) );
  NAND2_X1 U8357 ( .A1(n8592), .A2(n8596), .ZN(n6880) );
  OR2_X1 U8358 ( .A1(n6505), .A2(n7141), .ZN(n7142) );
  INV_X1 U8359 ( .A(n8455), .ZN(n6506) );
  OR2_X2 U8360 ( .A1(n10201), .A2(n6508), .ZN(n8467) );
  NAND2_X1 U8361 ( .A1(n6508), .A2(n10201), .ZN(n8485) );
  INV_X1 U8362 ( .A(n7355), .ZN(n8414) );
  NAND2_X1 U8363 ( .A1(n7356), .A2(n8414), .ZN(n6509) );
  INV_X1 U8364 ( .A(n7455), .ZN(n6510) );
  NAND2_X1 U8365 ( .A1(n6510), .A2(n4479), .ZN(n6511) );
  OR2_X1 U8366 ( .A1(n7461), .A2(n7555), .ZN(n8491) );
  OR2_X1 U8367 ( .A1(n7628), .A2(n7851), .ZN(n8471) );
  AND2_X1 U8368 ( .A1(n8471), .A2(n7597), .ZN(n8496) );
  NAND2_X1 U8369 ( .A1(n7628), .A2(n7851), .ZN(n8477) );
  INV_X1 U8370 ( .A(n7626), .ZN(n6513) );
  INV_X1 U8371 ( .A(n8422), .ZN(n6512) );
  AND2_X1 U8372 ( .A1(n7892), .A2(n8614), .ZN(n8483) );
  NAND2_X1 U8373 ( .A1(n8167), .A2(n8288), .ZN(n8500) );
  INV_X1 U8374 ( .A(n8613), .ZN(n8296) );
  AND2_X1 U8375 ( .A1(n8988), .A2(n8296), .ZN(n8450) );
  NAND2_X1 U8376 ( .A1(n8298), .A2(n8363), .ZN(n8452) );
  NAND2_X1 U8377 ( .A1(n9067), .A2(n8056), .ZN(n8510) );
  NAND2_X1 U8378 ( .A1(n6516), .A2(n8515), .ZN(n8904) );
  NAND2_X1 U8379 ( .A1(n8904), .A2(n8518), .ZN(n6517) );
  INV_X1 U8380 ( .A(n8889), .ZN(n6518) );
  NAND2_X1 U8381 ( .A1(n8888), .A2(n8533), .ZN(n8845) );
  INV_X1 U8382 ( .A(n8538), .ZN(n6519) );
  NOR2_X1 U8383 ( .A1(n6519), .A2(n4817), .ZN(n6520) );
  NAND2_X1 U8384 ( .A1(n8845), .A2(n6520), .ZN(n6523) );
  INV_X1 U8385 ( .A(n9034), .ZN(n8963) );
  NAND2_X1 U8386 ( .A1(n8846), .A2(n8867), .ZN(n6521) );
  AOI22_X1 U8387 ( .A1(n8963), .A2(n6521), .B1(n8526), .B2(n8838), .ZN(n6522)
         );
  NAND2_X1 U8388 ( .A1(n6523), .A2(n6522), .ZN(n8832) );
  NAND2_X1 U8389 ( .A1(n8261), .A2(n8826), .ZN(n8810) );
  NAND2_X1 U8390 ( .A1(n9007), .A2(n8815), .ZN(n8561) );
  NOR2_X1 U8391 ( .A1(n9001), .A2(n8257), .ZN(n8565) );
  INV_X1 U8392 ( .A(n8565), .ZN(n6526) );
  NAND2_X1 U8393 ( .A1(n9001), .A2(n8257), .ZN(n8432) );
  NAND2_X1 U8394 ( .A1(n8582), .A2(n8182), .ZN(n6534) );
  INV_X1 U8395 ( .A(n6555), .ZN(n6532) );
  NAND2_X1 U8396 ( .A1(n6530), .A2(n8585), .ZN(n7133) );
  AOI21_X1 U8397 ( .B1(n7133), .B2(n7841), .A(n8596), .ZN(n6531) );
  NAND2_X1 U8398 ( .A1(n6531), .A2(n6879), .ZN(n7691) );
  AOI21_X1 U8399 ( .B1(n6533), .B2(n6532), .A(n7691), .ZN(n6537) );
  INV_X1 U8400 ( .A(n6534), .ZN(n6535) );
  NAND2_X1 U8401 ( .A1(n6557), .A2(n6535), .ZN(n6536) );
  AOI21_X1 U8402 ( .B1(n6554), .B2(n6538), .A(n5228), .ZN(n6552) );
  NAND2_X1 U8403 ( .A1(n8778), .A2(n5227), .ZN(n6551) );
  NAND2_X1 U8404 ( .A1(n8589), .A2(n6539), .ZN(n6540) );
  AND2_X1 U8405 ( .A1(n6547), .A2(n6540), .ZN(n7127) );
  INV_X1 U8406 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n10561) );
  NAND2_X1 U8407 ( .A1(n6541), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6543) );
  INV_X1 U8408 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n10426) );
  OR2_X1 U8409 ( .A1(n7969), .A2(n10426), .ZN(n6542) );
  OAI211_X1 U8410 ( .C1(n10561), .C2(n6544), .A(n6543), .B(n6542), .ZN(n6545)
         );
  INV_X1 U8411 ( .A(n6545), .ZN(n6546) );
  NAND2_X1 U8412 ( .A1(n7976), .A2(n6546), .ZN(n8605) );
  AND2_X1 U8413 ( .A1(n6547), .A2(P2_B_REG_SCAN_IN), .ZN(n6548) );
  NOR2_X1 U8414 ( .A1(n8881), .A2(n6548), .ZN(n8770) );
  AOI22_X1 U8415 ( .A1(n10167), .A2(n8607), .B1(n8605), .B2(n8770), .ZN(n6549)
         );
  AOI21_X2 U8416 ( .B1(n6551), .B2(n6552), .A(n6550), .ZN(n6553) );
  NAND2_X1 U8417 ( .A1(n6554), .A2(n8779), .ZN(n6556) );
  XNOR2_X1 U8418 ( .A(n8397), .B(n6557), .ZN(n8073) );
  XNOR2_X1 U8419 ( .A(n6559), .B(P2_B_REG_SCAN_IN), .ZN(n6561) );
  NAND2_X1 U8420 ( .A1(n6561), .A2(n6560), .ZN(n6562) );
  INV_X1 U8421 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6953) );
  NAND2_X1 U8422 ( .A1(n6559), .A2(n8068), .ZN(n7131) );
  NAND2_X1 U8423 ( .A1(n6562), .A2(n6563), .ZN(n6951) );
  NAND2_X1 U8424 ( .A1(n6560), .A2(n8068), .ZN(n6564) );
  NAND2_X1 U8425 ( .A1(n7077), .A2(n9074), .ZN(n6878) );
  NOR4_X1 U8426 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n6574) );
  INV_X1 U8427 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10531) );
  INV_X1 U8428 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10461) );
  INV_X1 U8429 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10465) );
  INV_X1 U8430 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10499) );
  NAND4_X1 U8431 ( .A1(n10531), .A2(n10461), .A3(n10465), .A4(n10499), .ZN(
        n6571) );
  NOR4_X1 U8432 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6569) );
  NOR4_X1 U8433 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6568) );
  NOR4_X1 U8434 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6567) );
  NOR4_X1 U8435 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6566) );
  NAND4_X1 U8436 ( .A1(n6569), .A2(n6568), .A3(n6567), .A4(n6566), .ZN(n6570)
         );
  NOR4_X1 U8437 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        n6571), .A4(n6570), .ZN(n6573) );
  NOR4_X1 U8438 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6572) );
  AND3_X1 U8439 ( .A1(n6574), .A2(n6573), .A3(n6572), .ZN(n6575) );
  OR2_X1 U8440 ( .A1(n8570), .A2(n6577), .ZN(n7095) );
  AND3_X1 U8441 ( .A1(n6877), .A2(n7108), .A3(n7095), .ZN(n6578) );
  INV_X1 U8442 ( .A(n7077), .ZN(n6581) );
  NAND2_X1 U8443 ( .A1(n8440), .A2(n8587), .ZN(n6579) );
  NAND2_X1 U8444 ( .A1(n7130), .A2(n6579), .ZN(n6580) );
  NAND2_X1 U8445 ( .A1(n6580), .A2(n8592), .ZN(n7076) );
  OAI21_X1 U8446 ( .B1(n6581), .B2(n7078), .A(n7076), .ZN(n6584) );
  INV_X1 U8447 ( .A(n7076), .ZN(n6582) );
  NAND2_X1 U8448 ( .A1(n7073), .A2(n6582), .ZN(n6583) );
  INV_X1 U8449 ( .A(n10245), .ZN(n6586) );
  NAND2_X1 U8450 ( .A1(n6586), .A2(n10367), .ZN(n6587) );
  NAND2_X1 U8451 ( .A1(n6589), .A2(n5216), .ZN(P2_U3488) );
  INV_X1 U8452 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6590) );
  NAND2_X1 U8453 ( .A1(n6591), .A2(n5220), .ZN(P1_U3519) );
  NAND2_X1 U8454 ( .A1(n7843), .A2(n6595), .ZN(n6596) );
  NAND3_X2 U8455 ( .A1(n7769), .A2(n6596), .A3(n6908), .ZN(n6632) );
  NAND2_X1 U8456 ( .A1(n6619), .A2(n6601), .ZN(n6603) );
  NAND2_X1 U8457 ( .A1(n7411), .A2(n6837), .ZN(n6602) );
  NAND2_X1 U8458 ( .A1(n6603), .A2(n6602), .ZN(n6604) );
  INV_X4 U8459 ( .A(n6646), .ZN(n6841) );
  OAI21_X1 U8460 ( .B1(n6606), .B2(n6605), .A(n8125), .ZN(n7375) );
  INV_X1 U8461 ( .A(n7375), .ZN(n6618) );
  NAND2_X1 U8462 ( .A1(n7808), .A2(n6837), .ZN(n6608) );
  NAND2_X1 U8463 ( .A1(n6619), .A2(n7742), .ZN(n6607) );
  AND2_X1 U8464 ( .A1(n6608), .A2(n6607), .ZN(n6614) );
  INV_X1 U8465 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6609) );
  OR2_X1 U8466 ( .A1(n6908), .A2(n6609), .ZN(n6610) );
  NAND2_X1 U8467 ( .A1(n6614), .A2(n6610), .ZN(n7409) );
  NAND2_X1 U8468 ( .A1(n7808), .A2(n6818), .ZN(n6613) );
  AOI22_X1 U8469 ( .A1(n7742), .A2(n6837), .B1(n10061), .B2(n6611), .ZN(n6612)
         );
  NAND2_X1 U8470 ( .A1(n6613), .A2(n6612), .ZN(n7410) );
  NAND2_X1 U8471 ( .A1(n7409), .A2(n7410), .ZN(n6616) );
  NAND2_X1 U8472 ( .A1(n6614), .A2(n6841), .ZN(n6615) );
  NAND2_X1 U8473 ( .A1(n6616), .A2(n6615), .ZN(n7376) );
  NAND2_X1 U8474 ( .A1(n6618), .A2(n6617), .ZN(n8126) );
  NAND2_X1 U8475 ( .A1(n8126), .A2(n8125), .ZN(n6629) );
  NAND2_X1 U8476 ( .A1(n9561), .A2(n6665), .ZN(n6621) );
  NAND2_X1 U8477 ( .A1(n6693), .A2(n6097), .ZN(n6620) );
  NAND2_X1 U8478 ( .A1(n6621), .A2(n6620), .ZN(n6622) );
  XNOR2_X1 U8479 ( .A(n6622), .B(n6841), .ZN(n6627) );
  INV_X1 U8480 ( .A(n6627), .ZN(n6625) );
  AND2_X1 U8481 ( .A1(n6097), .A2(n6665), .ZN(n6623) );
  AOI21_X1 U8482 ( .B1(n9561), .B2(n6818), .A(n6623), .ZN(n6626) );
  INV_X1 U8483 ( .A(n6626), .ZN(n6624) );
  NAND2_X1 U8484 ( .A1(n6625), .A2(n6624), .ZN(n6628) );
  NAND2_X1 U8485 ( .A1(n6627), .A2(n6626), .ZN(n6630) );
  AND2_X1 U8486 ( .A1(n6628), .A2(n6630), .ZN(n8124) );
  NAND2_X1 U8487 ( .A1(n6629), .A2(n8124), .ZN(n8123) );
  NAND2_X1 U8488 ( .A1(n8123), .A2(n6630), .ZN(n7473) );
  INV_X1 U8489 ( .A(n6693), .ZN(n6707) );
  OAI22_X1 U8490 ( .A1(n8129), .A2(n6832), .B1(n10132), .B2(n6707), .ZN(n6631)
         );
  XNOR2_X1 U8491 ( .A(n6631), .B(n6841), .ZN(n6638) );
  OR2_X1 U8492 ( .A1(n8129), .A2(n6845), .ZN(n6634) );
  NAND2_X1 U8493 ( .A1(n7954), .A2(n6665), .ZN(n6633) );
  NAND2_X1 U8494 ( .A1(n6634), .A2(n6633), .ZN(n6636) );
  XNOR2_X1 U8495 ( .A(n6638), .B(n6636), .ZN(n7474) );
  OAI22_X1 U8496 ( .A1(n7948), .A2(n6832), .B1(n10116), .B2(n6707), .ZN(n6635)
         );
  XNOR2_X1 U8497 ( .A(n6635), .B(n6841), .ZN(n6640) );
  INV_X1 U8498 ( .A(n7452), .ZN(n10116) );
  OAI22_X1 U8499 ( .A1(n7948), .A2(n6845), .B1(n10116), .B2(n6832), .ZN(n6641)
         );
  XNOR2_X1 U8500 ( .A(n6640), .B(n6641), .ZN(n7399) );
  INV_X1 U8501 ( .A(n6636), .ZN(n6637) );
  NAND2_X1 U8502 ( .A1(n6638), .A2(n6637), .ZN(n7400) );
  AND2_X1 U8503 ( .A1(n7399), .A2(n7400), .ZN(n6639) );
  INV_X1 U8504 ( .A(n6640), .ZN(n6642) );
  NAND2_X1 U8505 ( .A1(n6642), .A2(n6641), .ZN(n6643) );
  NAND2_X1 U8506 ( .A1(n9558), .A2(n6843), .ZN(n6645) );
  NAND2_X1 U8507 ( .A1(n10139), .A2(n6838), .ZN(n6644) );
  NAND2_X1 U8508 ( .A1(n6645), .A2(n6644), .ZN(n6647) );
  XNOR2_X1 U8509 ( .A(n6647), .B(n6816), .ZN(n6649) );
  NAND2_X1 U8510 ( .A1(n6648), .A2(n6649), .ZN(n7504) );
  AOI22_X1 U8511 ( .A1(n9558), .A2(n6818), .B1(n10139), .B2(n6665), .ZN(n7506)
         );
  NAND2_X1 U8512 ( .A1(n7504), .A2(n7506), .ZN(n6652) );
  NAND2_X1 U8513 ( .A1(n6652), .A2(n7505), .ZN(n7574) );
  OAI22_X1 U8514 ( .A1(n9302), .A2(n6832), .B1(n10103), .B2(n6707), .ZN(n6653)
         );
  XNOR2_X1 U8515 ( .A(n6653), .B(n6841), .ZN(n6656) );
  OR2_X1 U8516 ( .A1(n9302), .A2(n6845), .ZN(n6655) );
  NAND2_X1 U8517 ( .A1(n7497), .A2(n6665), .ZN(n6654) );
  AND2_X1 U8518 ( .A1(n6655), .A2(n6654), .ZN(n6657) );
  NAND2_X1 U8519 ( .A1(n6656), .A2(n6657), .ZN(n6661) );
  INV_X1 U8520 ( .A(n6656), .ZN(n6659) );
  INV_X1 U8521 ( .A(n6657), .ZN(n6658) );
  NAND2_X1 U8522 ( .A1(n6659), .A2(n6658), .ZN(n6660) );
  AND2_X1 U8523 ( .A1(n6661), .A2(n6660), .ZN(n7575) );
  NAND2_X1 U8524 ( .A1(n9556), .A2(n6843), .ZN(n6663) );
  NAND2_X1 U8525 ( .A1(n6693), .A2(n10147), .ZN(n6662) );
  NAND2_X1 U8526 ( .A1(n6663), .A2(n6662), .ZN(n6664) );
  XNOR2_X1 U8527 ( .A(n6664), .B(n6841), .ZN(n6666) );
  AOI22_X1 U8528 ( .A1(n9556), .A2(n6818), .B1(n6665), .B2(n10147), .ZN(n6667)
         );
  AND2_X1 U8529 ( .A1(n6666), .A2(n6667), .ZN(n7640) );
  INV_X1 U8530 ( .A(n6666), .ZN(n6669) );
  INV_X1 U8531 ( .A(n6667), .ZN(n6668) );
  NAND2_X1 U8532 ( .A1(n6669), .A2(n6668), .ZN(n7638) );
  NAND2_X1 U8533 ( .A1(n4572), .A2(n6693), .ZN(n6671) );
  NAND2_X1 U8534 ( .A1(n9554), .A2(n6843), .ZN(n6670) );
  NAND2_X1 U8535 ( .A1(n6671), .A2(n6670), .ZN(n6672) );
  XNOR2_X1 U8536 ( .A(n6672), .B(n6816), .ZN(n6680) );
  NAND2_X1 U8537 ( .A1(n4572), .A2(n6843), .ZN(n6674) );
  NAND2_X1 U8538 ( .A1(n9554), .A2(n6818), .ZN(n6673) );
  NAND2_X1 U8539 ( .A1(n6674), .A2(n6673), .ZN(n9196) );
  NAND2_X1 U8540 ( .A1(n9555), .A2(n6843), .ZN(n6675) );
  OAI21_X1 U8541 ( .B1(n7783), .B2(n6707), .A(n6675), .ZN(n6676) );
  XNOR2_X1 U8542 ( .A(n6676), .B(n6816), .ZN(n6681) );
  OR2_X1 U8543 ( .A1(n7783), .A2(n6832), .ZN(n6678) );
  NAND2_X1 U8544 ( .A1(n9555), .A2(n6818), .ZN(n6677) );
  NAND2_X1 U8545 ( .A1(n6678), .A2(n6677), .ZN(n7980) );
  AOI22_X1 U8546 ( .A1(n6680), .A2(n9196), .B1(n6681), .B2(n7980), .ZN(n6679)
         );
  OAI21_X1 U8547 ( .B1(n6681), .B2(n7980), .A(n9196), .ZN(n6683) );
  INV_X1 U8548 ( .A(n6680), .ZN(n9197) );
  INV_X1 U8549 ( .A(n6681), .ZN(n9195) );
  NOR2_X1 U8550 ( .A1(n9196), .A2(n7980), .ZN(n6682) );
  AOI22_X1 U8551 ( .A1(n6683), .A2(n9197), .B1(n9195), .B2(n6682), .ZN(n6684)
         );
  NAND2_X1 U8552 ( .A1(n9326), .A2(n6693), .ZN(n6687) );
  NAND2_X1 U8553 ( .A1(n9552), .A2(n6843), .ZN(n6686) );
  NAND2_X1 U8554 ( .A1(n6687), .A2(n6686), .ZN(n6688) );
  XNOR2_X1 U8555 ( .A(n6688), .B(n6816), .ZN(n9243) );
  NAND2_X1 U8556 ( .A1(n9326), .A2(n6843), .ZN(n6690) );
  NAND2_X1 U8557 ( .A1(n9552), .A2(n6818), .ZN(n6689) );
  NAND2_X1 U8558 ( .A1(n6690), .A2(n6689), .ZN(n6701) );
  NAND2_X1 U8559 ( .A1(n9113), .A2(n6843), .ZN(n6692) );
  NAND2_X1 U8560 ( .A1(n9553), .A2(n6818), .ZN(n6691) );
  NAND2_X1 U8561 ( .A1(n6692), .A2(n6691), .ZN(n9107) );
  NAND2_X1 U8562 ( .A1(n9113), .A2(n6693), .ZN(n6695) );
  NAND2_X1 U8563 ( .A1(n9553), .A2(n6843), .ZN(n6694) );
  NAND2_X1 U8564 ( .A1(n6695), .A2(n6694), .ZN(n6696) );
  XNOR2_X1 U8565 ( .A(n6696), .B(n6816), .ZN(n6698) );
  AOI22_X1 U8566 ( .A1(n9243), .A2(n6701), .B1(n9107), .B2(n6698), .ZN(n6697)
         );
  NAND2_X1 U8567 ( .A1(n9240), .A2(n6697), .ZN(n6706) );
  INV_X1 U8568 ( .A(n9243), .ZN(n6704) );
  INV_X1 U8569 ( .A(n6698), .ZN(n9241) );
  INV_X1 U8570 ( .A(n9107), .ZN(n6699) );
  NAND2_X1 U8571 ( .A1(n9241), .A2(n6699), .ZN(n6700) );
  NAND2_X1 U8572 ( .A1(n6700), .A2(n6701), .ZN(n6703) );
  INV_X1 U8573 ( .A(n6700), .ZN(n6702) );
  INV_X1 U8574 ( .A(n6701), .ZN(n9242) );
  AOI22_X1 U8575 ( .A1(n6704), .A2(n6703), .B1(n6702), .B2(n9242), .ZN(n6705)
         );
  NAND2_X1 U8576 ( .A1(n6706), .A2(n6705), .ZN(n9139) );
  OAI22_X1 U8577 ( .A1(n7867), .A2(n6707), .B1(n9251), .B2(n6832), .ZN(n6708)
         );
  XNOR2_X1 U8578 ( .A(n6708), .B(n6841), .ZN(n6711) );
  OAI22_X1 U8579 ( .A1(n7867), .A2(n6832), .B1(n9251), .B2(n6845), .ZN(n6709)
         );
  XNOR2_X1 U8580 ( .A(n6711), .B(n6709), .ZN(n9141) );
  INV_X1 U8581 ( .A(n6709), .ZN(n6710) );
  NAND2_X1 U8582 ( .A1(n6711), .A2(n6710), .ZN(n6712) );
  NAND2_X1 U8583 ( .A1(n10008), .A2(n6838), .ZN(n6714) );
  NAND2_X1 U8584 ( .A1(n9551), .A2(n6843), .ZN(n6713) );
  NAND2_X1 U8585 ( .A1(n6714), .A2(n6713), .ZN(n6715) );
  XNOR2_X1 U8586 ( .A(n6715), .B(n6816), .ZN(n6717) );
  AND2_X1 U8587 ( .A1(n9551), .A2(n6818), .ZN(n6716) );
  AOI21_X1 U8588 ( .B1(n10008), .B2(n6843), .A(n6716), .ZN(n6718) );
  XNOR2_X1 U8589 ( .A(n6717), .B(n6718), .ZN(n9219) );
  INV_X1 U8590 ( .A(n6717), .ZN(n6719) );
  NAND2_X1 U8591 ( .A1(n6720), .A2(n6838), .ZN(n6722) );
  NAND2_X1 U8592 ( .A1(n9550), .A2(n6843), .ZN(n6721) );
  NAND2_X1 U8593 ( .A1(n6722), .A2(n6721), .ZN(n6723) );
  XNOR2_X1 U8594 ( .A(n6723), .B(n6816), .ZN(n9163) );
  NAND2_X1 U8595 ( .A1(n5807), .A2(n6843), .ZN(n6725) );
  NAND2_X1 U8596 ( .A1(n9550), .A2(n6818), .ZN(n6724) );
  NAND2_X1 U8597 ( .A1(n6725), .A2(n6724), .ZN(n9162) );
  NAND2_X1 U8598 ( .A1(n9998), .A2(n6838), .ZN(n6727) );
  NAND2_X1 U8599 ( .A1(n9868), .A2(n6843), .ZN(n6726) );
  NAND2_X1 U8600 ( .A1(n6727), .A2(n6726), .ZN(n6728) );
  XNOR2_X1 U8601 ( .A(n6728), .B(n6816), .ZN(n9160) );
  NAND2_X1 U8602 ( .A1(n9998), .A2(n6843), .ZN(n6730) );
  NAND2_X1 U8603 ( .A1(n9868), .A2(n6818), .ZN(n6729) );
  NAND2_X1 U8604 ( .A1(n6730), .A2(n6729), .ZN(n6740) );
  AND2_X1 U8605 ( .A1(n9160), .A2(n6740), .ZN(n6731) );
  AOI21_X1 U8606 ( .B1(n9163), .B2(n9162), .A(n6731), .ZN(n6738) );
  NAND2_X1 U8607 ( .A1(n10003), .A2(n6838), .ZN(n6733) );
  NAND2_X1 U8608 ( .A1(n9914), .A2(n6843), .ZN(n6732) );
  NAND2_X1 U8609 ( .A1(n6733), .A2(n6732), .ZN(n6734) );
  XNOR2_X1 U8610 ( .A(n6734), .B(n6816), .ZN(n9155) );
  NAND2_X1 U8611 ( .A1(n10003), .A2(n6843), .ZN(n6736) );
  NAND2_X1 U8612 ( .A1(n9914), .A2(n6818), .ZN(n6735) );
  NAND2_X1 U8613 ( .A1(n6736), .A2(n6735), .ZN(n9093) );
  NAND2_X1 U8614 ( .A1(n9155), .A2(n9093), .ZN(n6737) );
  INV_X1 U8615 ( .A(n6738), .ZN(n6739) );
  OR3_X1 U8616 ( .A1(n6739), .A2(n9093), .A3(n9155), .ZN(n6747) );
  INV_X1 U8617 ( .A(n9163), .ZN(n6745) );
  INV_X1 U8618 ( .A(n9160), .ZN(n9159) );
  INV_X1 U8619 ( .A(n6740), .ZN(n9275) );
  NAND2_X1 U8620 ( .A1(n9159), .A2(n9275), .ZN(n6741) );
  NAND2_X1 U8621 ( .A1(n6741), .A2(n9162), .ZN(n6744) );
  INV_X1 U8622 ( .A(n6741), .ZN(n6743) );
  INV_X1 U8623 ( .A(n9162), .ZN(n6742) );
  AOI22_X1 U8624 ( .A1(n6745), .A2(n6744), .B1(n6743), .B2(n6742), .ZN(n6746)
         );
  AND2_X1 U8625 ( .A1(n6747), .A2(n6746), .ZN(n6748) );
  NAND2_X1 U8626 ( .A1(n9988), .A2(n6838), .ZN(n6751) );
  NAND2_X1 U8627 ( .A1(n9867), .A2(n6843), .ZN(n6750) );
  NAND2_X1 U8628 ( .A1(n6751), .A2(n6750), .ZN(n6752) );
  XNOR2_X1 U8629 ( .A(n6752), .B(n6841), .ZN(n9171) );
  AND2_X1 U8630 ( .A1(n9867), .A2(n6818), .ZN(n6753) );
  AOI21_X1 U8631 ( .B1(n9988), .B2(n6843), .A(n6753), .ZN(n9170) );
  INV_X1 U8632 ( .A(n9171), .ZN(n6755) );
  INV_X1 U8633 ( .A(n9170), .ZN(n6754) );
  NAND2_X1 U8634 ( .A1(n6755), .A2(n6754), .ZN(n9116) );
  NAND2_X1 U8635 ( .A1(n9975), .A2(n6838), .ZN(n6757) );
  NAND2_X1 U8636 ( .A1(n9820), .A2(n6843), .ZN(n6756) );
  NAND2_X1 U8637 ( .A1(n6757), .A2(n6756), .ZN(n6758) );
  XNOR2_X1 U8638 ( .A(n6758), .B(n6816), .ZN(n6772) );
  AND2_X1 U8639 ( .A1(n9820), .A2(n6818), .ZN(n6759) );
  AOI21_X1 U8640 ( .B1(n9975), .B2(n6843), .A(n6759), .ZN(n6773) );
  XNOR2_X1 U8641 ( .A(n6772), .B(n6773), .ZN(n9121) );
  NAND2_X1 U8642 ( .A1(n9983), .A2(n6838), .ZN(n6761) );
  NAND2_X1 U8643 ( .A1(n9835), .A2(n6843), .ZN(n6760) );
  NAND2_X1 U8644 ( .A1(n6761), .A2(n6760), .ZN(n6762) );
  XNOR2_X1 U8645 ( .A(n6762), .B(n6841), .ZN(n9118) );
  INV_X1 U8646 ( .A(n9118), .ZN(n6765) );
  NAND2_X1 U8647 ( .A1(n9983), .A2(n6843), .ZN(n6764) );
  NAND2_X1 U8648 ( .A1(n9835), .A2(n6818), .ZN(n6763) );
  AND2_X1 U8649 ( .A1(n6764), .A2(n6763), .ZN(n6768) );
  INV_X1 U8650 ( .A(n6768), .ZN(n9257) );
  NAND2_X1 U8651 ( .A1(n6765), .A2(n9257), .ZN(n6766) );
  AND2_X1 U8652 ( .A1(n9121), .A2(n6766), .ZN(n6767) );
  AND2_X1 U8653 ( .A1(n9116), .A2(n6767), .ZN(n6771) );
  INV_X1 U8654 ( .A(n6767), .ZN(n6770) );
  NAND2_X1 U8655 ( .A1(n9118), .A2(n6768), .ZN(n6769) );
  INV_X1 U8656 ( .A(n6772), .ZN(n6774) );
  NAND2_X1 U8657 ( .A1(n9971), .A2(n6838), .ZN(n6776) );
  NAND2_X1 U8658 ( .A1(n9836), .A2(n6843), .ZN(n6775) );
  NAND2_X1 U8659 ( .A1(n6776), .A2(n6775), .ZN(n6777) );
  XNOR2_X1 U8660 ( .A(n6777), .B(n6841), .ZN(n6779) );
  AND2_X1 U8661 ( .A1(n9836), .A2(n6818), .ZN(n6778) );
  AOI21_X1 U8662 ( .B1(n9971), .B2(n6843), .A(n6778), .ZN(n6780) );
  AND2_X1 U8663 ( .A1(n6779), .A2(n6780), .ZN(n9208) );
  INV_X1 U8664 ( .A(n6779), .ZN(n6782) );
  INV_X1 U8665 ( .A(n6780), .ZN(n6781) );
  NAND2_X1 U8666 ( .A1(n6782), .A2(n6781), .ZN(n9207) );
  NAND2_X1 U8667 ( .A1(n9966), .A2(n6838), .ZN(n6784) );
  NAND2_X1 U8668 ( .A1(n9821), .A2(n6843), .ZN(n6783) );
  NAND2_X1 U8669 ( .A1(n6784), .A2(n6783), .ZN(n6785) );
  XNOR2_X1 U8670 ( .A(n6785), .B(n6841), .ZN(n6789) );
  AND2_X1 U8671 ( .A1(n9821), .A2(n6818), .ZN(n6786) );
  AOI21_X1 U8672 ( .B1(n9966), .B2(n6837), .A(n6786), .ZN(n6788) );
  XNOR2_X1 U8673 ( .A(n6789), .B(n6788), .ZN(n9133) );
  INV_X1 U8674 ( .A(n9133), .ZN(n6787) );
  NAND2_X1 U8675 ( .A1(n6789), .A2(n6788), .ZN(n6790) );
  NAND2_X1 U8676 ( .A1(n9960), .A2(n6838), .ZN(n6792) );
  NAND2_X1 U8677 ( .A1(n9805), .A2(n6843), .ZN(n6791) );
  NAND2_X1 U8678 ( .A1(n6792), .A2(n6791), .ZN(n6793) );
  XNOR2_X1 U8679 ( .A(n6793), .B(n6816), .ZN(n6795) );
  AND2_X1 U8680 ( .A1(n9805), .A2(n6818), .ZN(n6794) );
  AOI21_X1 U8681 ( .B1(n9960), .B2(n6843), .A(n6794), .ZN(n9228) );
  NAND2_X1 U8682 ( .A1(n9957), .A2(n6838), .ZN(n6797) );
  NAND2_X1 U8683 ( .A1(n9796), .A2(n6843), .ZN(n6796) );
  NAND2_X1 U8684 ( .A1(n6797), .A2(n6796), .ZN(n6798) );
  XNOR2_X1 U8685 ( .A(n6798), .B(n6816), .ZN(n6800) );
  AND2_X1 U8686 ( .A1(n9796), .A2(n6818), .ZN(n6799) );
  AOI21_X1 U8687 ( .B1(n9957), .B2(n6843), .A(n6799), .ZN(n6801) );
  XNOR2_X1 U8688 ( .A(n6800), .B(n6801), .ZN(n9101) );
  INV_X1 U8689 ( .A(n6800), .ZN(n6802) );
  NAND2_X1 U8690 ( .A1(n6802), .A2(n6801), .ZN(n6803) );
  NAND2_X1 U8691 ( .A1(n6804), .A2(n6803), .ZN(n9186) );
  NAND2_X1 U8692 ( .A1(n9950), .A2(n6838), .ZN(n6806) );
  NAND2_X1 U8693 ( .A1(n9549), .A2(n6843), .ZN(n6805) );
  NAND2_X1 U8694 ( .A1(n6806), .A2(n6805), .ZN(n6807) );
  XNOR2_X1 U8695 ( .A(n6807), .B(n6816), .ZN(n6809) );
  NOR2_X1 U8696 ( .A1(n9771), .A2(n6845), .ZN(n6808) );
  AOI21_X1 U8697 ( .B1(n9950), .B2(n6837), .A(n6808), .ZN(n6810) );
  XNOR2_X1 U8698 ( .A(n6809), .B(n6810), .ZN(n9188) );
  NAND2_X1 U8699 ( .A1(n9186), .A2(n9188), .ZN(n6813) );
  INV_X1 U8700 ( .A(n6809), .ZN(n6811) );
  NAND2_X1 U8701 ( .A1(n6811), .A2(n6810), .ZN(n6812) );
  NAND2_X1 U8702 ( .A1(n6813), .A2(n6812), .ZN(n9148) );
  NAND2_X1 U8703 ( .A1(n9741), .A2(n6838), .ZN(n6815) );
  NAND2_X1 U8704 ( .A1(n9750), .A2(n6843), .ZN(n6814) );
  NAND2_X1 U8705 ( .A1(n6815), .A2(n6814), .ZN(n6817) );
  XNOR2_X1 U8706 ( .A(n6817), .B(n6816), .ZN(n6820) );
  AND2_X1 U8707 ( .A1(n9750), .A2(n6818), .ZN(n6819) );
  AOI21_X1 U8708 ( .B1(n9741), .B2(n6843), .A(n6819), .ZN(n6821) );
  XNOR2_X1 U8709 ( .A(n6820), .B(n6821), .ZN(n9149) );
  INV_X1 U8710 ( .A(n6820), .ZN(n6822) );
  NAND2_X1 U8711 ( .A1(n6822), .A2(n6821), .ZN(n6823) );
  NAND2_X1 U8712 ( .A1(n9723), .A2(n6838), .ZN(n6825) );
  NAND2_X1 U8713 ( .A1(n9548), .A2(n6843), .ZN(n6824) );
  NAND2_X1 U8714 ( .A1(n6825), .A2(n6824), .ZN(n6826) );
  XNOR2_X1 U8715 ( .A(n6826), .B(n6841), .ZN(n6830) );
  NOR2_X1 U8716 ( .A1(n9736), .A2(n6845), .ZN(n6827) );
  AOI21_X1 U8717 ( .B1(n9723), .B2(n6837), .A(n6827), .ZN(n6829) );
  XNOR2_X1 U8718 ( .A(n6830), .B(n6829), .ZN(n9263) );
  INV_X1 U8719 ( .A(n9263), .ZN(n6828) );
  OR2_X1 U8720 ( .A1(n6830), .A2(n6829), .ZN(n6831) );
  NAND2_X1 U8721 ( .A1(n8118), .A2(n6838), .ZN(n6834) );
  OR2_X1 U8722 ( .A1(n9718), .A2(n6832), .ZN(n6833) );
  NAND2_X1 U8723 ( .A1(n6834), .A2(n6833), .ZN(n6835) );
  XNOR2_X1 U8724 ( .A(n6835), .B(n6841), .ZN(n6853) );
  NOR2_X1 U8725 ( .A1(n9718), .A2(n6845), .ZN(n6836) );
  AOI21_X1 U8726 ( .B1(n8118), .B2(n6837), .A(n6836), .ZN(n6852) );
  XNOR2_X1 U8727 ( .A(n6853), .B(n6852), .ZN(n8113) );
  NAND2_X1 U8728 ( .A1(n6873), .A2(n6838), .ZN(n6840) );
  NAND2_X1 U8729 ( .A1(n9546), .A2(n6843), .ZN(n6839) );
  NAND2_X1 U8730 ( .A1(n6840), .A2(n6839), .ZN(n6842) );
  XNOR2_X1 U8731 ( .A(n6842), .B(n6841), .ZN(n6847) );
  NAND2_X1 U8732 ( .A1(n6873), .A2(n6843), .ZN(n6844) );
  OAI21_X1 U8733 ( .B1(n9703), .B2(n6845), .A(n6844), .ZN(n6846) );
  XNOR2_X1 U8734 ( .A(n6847), .B(n6846), .ZN(n6855) );
  INV_X1 U8735 ( .A(n6855), .ZN(n6870) );
  INV_X1 U8736 ( .A(n7731), .ZN(n6849) );
  NAND3_X1 U8737 ( .A1(n6849), .A2(n7732), .A3(n6848), .ZN(n6862) );
  AND2_X1 U8738 ( .A1(n6908), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6850) );
  NOR2_X1 U8739 ( .A1(n10148), .A2(n7028), .ZN(n6851) );
  NAND2_X1 U8740 ( .A1(n6853), .A2(n6852), .ZN(n6869) );
  NAND3_X1 U8741 ( .A1(n6870), .A2(n9276), .A3(n6869), .ZN(n6854) );
  OR2_X2 U8742 ( .A1(n8112), .A2(n6854), .ZN(n6876) );
  NAND2_X1 U8743 ( .A1(n8112), .A2(n6856), .ZN(n6875) );
  NAND2_X1 U8744 ( .A1(n7337), .A2(n9527), .ZN(n7740) );
  OAI21_X1 U8745 ( .B1(n6858), .B2(n7740), .A(n9922), .ZN(n9223) );
  AND2_X1 U8746 ( .A1(n9915), .A2(n6595), .ZN(n6859) );
  NAND2_X1 U8747 ( .A1(n6866), .A2(n6859), .ZN(n9279) );
  INV_X1 U8748 ( .A(n6860), .ZN(n6864) );
  NAND2_X1 U8749 ( .A1(n9527), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7582) );
  NAND2_X1 U8750 ( .A1(n10148), .A2(n7582), .ZN(n6861) );
  NAND2_X1 U8751 ( .A1(n6862), .A2(n6861), .ZN(n6863) );
  NAND2_X1 U8752 ( .A1(n6864), .A2(n6863), .ZN(n9174) );
  AOI22_X1 U8753 ( .A1(n8242), .A2(n9267), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6868) );
  AND2_X1 U8754 ( .A1(n9913), .A2(n6595), .ZN(n6865) );
  NAND2_X1 U8755 ( .A1(n9545), .A2(n9284), .ZN(n6867) );
  OAI211_X1 U8756 ( .C1(n9718), .C2(n9279), .A(n6868), .B(n6867), .ZN(n6872)
         );
  NOR3_X1 U8757 ( .A1(n6870), .A2(n9262), .A3(n6869), .ZN(n6871) );
  AOI211_X1 U8758 ( .C1(n6873), .C2(n9236), .A(n6872), .B(n6871), .ZN(n6874)
         );
  NAND3_X1 U8759 ( .A1(n6876), .A2(n6875), .A3(n6874), .ZN(P1_U3220) );
  INV_X1 U8760 ( .A(n6879), .ZN(n7081) );
  NAND2_X1 U8761 ( .A1(n7108), .A2(n7081), .ZN(n7104) );
  OR3_X1 U8762 ( .A1(n6530), .A2(n8585), .A3(n6880), .ZN(n7089) );
  INV_X1 U8763 ( .A(n7089), .ZN(n7090) );
  NAND2_X1 U8764 ( .A1(n7108), .A2(n7090), .ZN(n6881) );
  NAND2_X1 U8765 ( .A1(n7104), .A2(n6881), .ZN(n6882) );
  NAND2_X1 U8766 ( .A1(n7107), .A2(n6882), .ZN(n6888) );
  NOR2_X1 U8767 ( .A1(n7077), .A2(n6883), .ZN(n6884) );
  NAND2_X1 U8768 ( .A1(n8570), .A2(n7089), .ZN(n6886) );
  INV_X1 U8769 ( .A(n7171), .ZN(n6885) );
  NAND2_X1 U8770 ( .A1(n10189), .A2(n6885), .ZN(n8928) );
  OAI21_X1 U8771 ( .B1(n6886), .B2(n10189), .A(n8928), .ZN(n7094) );
  NAND3_X1 U8772 ( .A1(n7105), .A2(n7108), .A3(n7094), .ZN(n6887) );
  INV_X1 U8773 ( .A(n10189), .ZN(n10223) );
  NAND2_X1 U8774 ( .A1(n6890), .A2(n5219), .ZN(P2_U3456) );
  OR3_X1 U8775 ( .A1(n7872), .A2(n6892), .A3(n6891), .ZN(n6893) );
  AOI21_X1 U8776 ( .B1(n6894), .B2(n6893), .A(n8768), .ZN(n6907) );
  INV_X1 U8777 ( .A(n6895), .ZN(n6898) );
  NAND3_X1 U8778 ( .A1(n7882), .A2(n6896), .A3(n4438), .ZN(n6897) );
  INV_X1 U8779 ( .A(n8750), .ZN(n8739) );
  AOI21_X1 U8780 ( .B1(n6898), .B2(n6897), .A(n8739), .ZN(n6906) );
  INV_X1 U8781 ( .A(n6899), .ZN(n8652) );
  NAND3_X1 U8782 ( .A1(n7878), .A2(n6901), .A3(n6900), .ZN(n6902) );
  AOI21_X1 U8783 ( .B1(n8652), .B2(n6902), .A(n8760), .ZN(n6905) );
  INV_X1 U8784 ( .A(n8759), .ZN(n8728) );
  NOR2_X1 U8785 ( .A1(n10445), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8293) );
  AOI21_X1 U8786 ( .B1(n8728), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8293), .ZN(
        n6903) );
  OAI21_X1 U8787 ( .B1(n8755), .B2(n6978), .A(n6903), .ZN(n6904) );
  OR4_X1 U8788 ( .A1(n6907), .A2(n6906), .A3(n6905), .A4(n6904), .ZN(P2_U3194)
         );
  NOR2_X1 U8789 ( .A1(n6908), .A2(P1_U3086), .ZN(n6909) );
  AND2_X2 U8790 ( .A1(n7029), .A2(n6909), .ZN(P1_U3973) );
  OR3_X1 U8791 ( .A1(n6912), .A2(n6910), .A3(n6911), .ZN(n6913) );
  AOI21_X1 U8792 ( .B1(n6914), .B2(n6913), .A(n8768), .ZN(n6925) );
  NAND3_X1 U8793 ( .A1(n7391), .A2(n6916), .A3(n6915), .ZN(n6917) );
  AOI21_X1 U8794 ( .B1(n4763), .B2(n6917), .A(n8760), .ZN(n6924) );
  NAND3_X1 U8795 ( .A1(n7383), .A2(n4537), .A3(n6918), .ZN(n6919) );
  AOI21_X1 U8796 ( .B1(n6920), .B2(n6919), .A(n8739), .ZN(n6923) );
  AND2_X1 U8797 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7594) );
  AOI21_X1 U8798 ( .B1(n8728), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7594), .ZN(
        n6921) );
  OAI21_X1 U8799 ( .B1(n8755), .B2(n6938), .A(n6921), .ZN(n6922) );
  OR4_X1 U8800 ( .A1(n6925), .A2(n6924), .A3(n6923), .A4(n6922), .ZN(P2_U3190)
         );
  AND2_X1 U8801 ( .A1(n8144), .A2(P2_U3151), .ZN(n9088) );
  INV_X2 U8802 ( .A(n9088), .ZN(n9077) );
  NOR2_X1 U8803 ( .A1(n8144), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9081) );
  INV_X2 U8804 ( .A(n9081), .ZN(n9090) );
  OAI222_X1 U8805 ( .A1(n9077), .A2(n6926), .B1(n9090), .B2(n6947), .C1(
        P2_U3151), .C2(n6994), .ZN(P2_U3293) );
  OAI222_X1 U8806 ( .A1(n9077), .A2(n6927), .B1(n9090), .B2(n6943), .C1(
        P2_U3151), .C2(n7233), .ZN(P2_U3291) );
  OAI222_X1 U8807 ( .A1(P2_U3151), .A2(n6928), .B1(n9090), .B2(n6942), .C1(
        n4620), .C2(n9077), .ZN(P2_U3292) );
  AND2_X1 U8808 ( .A1(n8144), .A2(P1_U3086), .ZN(n10043) );
  INV_X2 U8809 ( .A(n10043), .ZN(n10058) );
  AND2_X1 U8810 ( .A1(n6929), .A2(P1_U3086), .ZN(n7329) );
  INV_X2 U8811 ( .A(n7329), .ZN(n10060) );
  OAI222_X1 U8812 ( .A1(n10058), .A2(n6936), .B1(n10060), .B2(n4970), .C1(
        P1_U3086), .C2(n7037), .ZN(P1_U3354) );
  OAI222_X1 U8813 ( .A1(P2_U3151), .A2(n6930), .B1(n9090), .B2(n6239), .C1(
        n5565), .C2(n9077), .ZN(P2_U3290) );
  INV_X1 U8814 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6931) );
  OAI222_X1 U8815 ( .A1(P2_U3151), .A2(n7385), .B1(n9090), .B2(n6932), .C1(
        n6931), .C2(n9077), .ZN(P2_U3288) );
  INV_X1 U8816 ( .A(n7198), .ZN(n7279) );
  OAI222_X1 U8817 ( .A1(n10060), .A2(n6933), .B1(n10058), .B2(n6932), .C1(
        n7279), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U8818 ( .A(n6934), .ZN(n6949) );
  OAI222_X1 U8819 ( .A1(n9077), .A2(n6935), .B1(n9090), .B2(n6949), .C1(
        P2_U3151), .C2(n7021), .ZN(P2_U3289) );
  OAI222_X1 U8820 ( .A1(P2_U3151), .A2(n7009), .B1(n9077), .B2(n4967), .C1(
        n6936), .C2(n9090), .ZN(P2_U3294) );
  INV_X1 U8821 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6939) );
  INV_X1 U8822 ( .A(n6937), .ZN(n6945) );
  OAI222_X1 U8823 ( .A1(n9077), .A2(n6939), .B1(n9090), .B2(n6945), .C1(
        P2_U3151), .C2(n6938), .ZN(P2_U3287) );
  INV_X1 U8824 ( .A(n9596), .ZN(n6940) );
  OAI222_X1 U8825 ( .A1(n10058), .A2(n6942), .B1(n10060), .B2(n6941), .C1(
        P1_U3086), .C2(n6940), .ZN(P1_U3352) );
  OAI222_X1 U8826 ( .A1(n10060), .A2(n6944), .B1(n10058), .B2(n6943), .C1(
        P1_U3086), .C2(n9608), .ZN(P1_U3351) );
  INV_X1 U8827 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6946) );
  INV_X1 U8828 ( .A(n7286), .ZN(n7295) );
  OAI222_X1 U8829 ( .A1(n10060), .A2(n6946), .B1(n10058), .B2(n6945), .C1(
        P1_U3086), .C2(n7295), .ZN(P1_U3347) );
  OAI222_X1 U8830 ( .A1(n10060), .A2(n6948), .B1(n10058), .B2(n6947), .C1(
        P1_U3086), .C2(n9580), .ZN(P1_U3353) );
  INV_X1 U8831 ( .A(n7197), .ZN(n7072) );
  OAI222_X1 U8832 ( .A1(n10060), .A2(n6950), .B1(n10058), .B2(n6949), .C1(
        P1_U3086), .C2(n7072), .ZN(P1_U3349) );
  NOR3_X1 U8833 ( .A1(n7131), .A2(n7935), .A3(P2_U3151), .ZN(n6952) );
  AOI21_X1 U8834 ( .B1(n6961), .B2(n6953), .A(n6952), .ZN(P2_U3376) );
  AND2_X1 U8835 ( .A1(n6961), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8836 ( .A1(n6961), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8837 ( .A1(n6961), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8838 ( .A1(n6961), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8839 ( .A1(n6961), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8840 ( .A1(n6961), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8841 ( .A1(n6961), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8842 ( .A1(n6961), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8843 ( .A1(n6961), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8844 ( .A1(n6961), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8845 ( .A1(n6961), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8846 ( .A1(n6961), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8847 ( .A1(n6961), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8848 ( .A1(n6961), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8849 ( .A1(n6961), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8850 ( .A1(n6961), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8851 ( .A1(n6961), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8852 ( .A1(n6961), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8853 ( .A1(n6961), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8854 ( .A1(n6961), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8855 ( .A1(n6961), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  INV_X1 U8856 ( .A(n7058), .ZN(n7061) );
  OAI222_X1 U8857 ( .A1(n10060), .A2(n6954), .B1(n10058), .B2(n6239), .C1(
        n7061), .C2(P1_U3086), .ZN(P1_U3350) );
  INV_X1 U8858 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6955) );
  INV_X1 U8859 ( .A(n7317), .ZN(n7319) );
  OAI222_X1 U8860 ( .A1(n10060), .A2(n6955), .B1(n10058), .B2(n6956), .C1(
        n7319), .C2(P1_U3086), .ZN(P1_U3345) );
  OAI222_X1 U8861 ( .A1(P2_U3151), .A2(n6957), .B1(n9090), .B2(n6956), .C1(
        n4601), .C2(n9077), .ZN(P2_U3285) );
  INV_X1 U8862 ( .A(n6958), .ZN(n6959) );
  OAI222_X1 U8863 ( .A1(P2_U3151), .A2(n4923), .B1(n9090), .B2(n6959), .C1(
        n4655), .C2(n9077), .ZN(P2_U3286) );
  INV_X1 U8864 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6960) );
  INV_X1 U8865 ( .A(n7201), .ZN(n10073) );
  OAI222_X1 U8866 ( .A1(n10060), .A2(n6960), .B1(n10058), .B2(n6959), .C1(
        n10073), .C2(P1_U3086), .ZN(P1_U3346) );
  NOR2_X1 U8867 ( .A1(n6962), .A2(n10461), .ZN(P2_U3254) );
  NOR2_X1 U8868 ( .A1(n6962), .A2(n10499), .ZN(P2_U3238) );
  INV_X1 U8869 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10406) );
  NOR2_X1 U8870 ( .A1(n6962), .A2(n10406), .ZN(P2_U3258) );
  NOR2_X1 U8871 ( .A1(n6962), .A2(n10531), .ZN(P2_U3245) );
  INV_X1 U8872 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10396) );
  NOR2_X1 U8873 ( .A1(n6962), .A2(n10396), .ZN(P2_U3237) );
  INV_X1 U8874 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n10430) );
  NOR2_X1 U8875 ( .A1(n6962), .A2(n10430), .ZN(P2_U3257) );
  INV_X1 U8876 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10334) );
  NOR2_X1 U8877 ( .A1(n6962), .A2(n10334), .ZN(P2_U3240) );
  INV_X1 U8878 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n10347) );
  NOR2_X1 U8879 ( .A1(n6962), .A2(n10347), .ZN(P2_U3234) );
  NOR2_X1 U8880 ( .A1(n6962), .A2(n10465), .ZN(P2_U3244) );
  INV_X1 U8881 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6964) );
  INV_X1 U8882 ( .A(n6963), .ZN(n6972) );
  INV_X1 U8883 ( .A(n7517), .ZN(n7521) );
  OAI222_X1 U8884 ( .A1(n10060), .A2(n6964), .B1(n10058), .B2(n6972), .C1(
        P1_U3086), .C2(n7521), .ZN(P1_U3344) );
  INV_X1 U8885 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6971) );
  NAND2_X1 U8886 ( .A1(n6965), .A2(n4436), .ZN(n6966) );
  AOI22_X1 U8887 ( .A1(n6967), .A2(n8760), .B1(n7002), .B2(n6966), .ZN(n6968)
         );
  AOI21_X1 U8888 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n6968), .ZN(
        n6970) );
  NAND2_X1 U8889 ( .A1(n8718), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6969) );
  OAI211_X1 U8890 ( .C1(n8759), .C2(n6971), .A(n6970), .B(n6969), .ZN(P2_U3182) );
  OAI222_X1 U8891 ( .A1(n4634), .A2(n9077), .B1(P2_U3151), .B2(n6973), .C1(
        n9090), .C2(n6972), .ZN(P2_U3284) );
  NAND2_X1 U8892 ( .A1(n7411), .A2(P1_U3973), .ZN(n6974) );
  OAI21_X1 U8893 ( .B1(P1_U3973), .B2(n4967), .A(n6974), .ZN(P1_U3555) );
  INV_X1 U8894 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6976) );
  INV_X1 U8895 ( .A(n6975), .ZN(n6977) );
  INV_X1 U8896 ( .A(n7524), .ZN(n10089) );
  OAI222_X1 U8897 ( .A1(n10060), .A2(n6976), .B1(n10058), .B2(n6977), .C1(
        n10089), .C2(P1_U3086), .ZN(P1_U3343) );
  OAI222_X1 U8898 ( .A1(P2_U3151), .A2(n6978), .B1(n9090), .B2(n6977), .C1(
        n4636), .C2(n9077), .ZN(P2_U3283) );
  INV_X1 U8899 ( .A(n8760), .ZN(n8733) );
  XOR2_X1 U8900 ( .A(n6980), .B(n6979), .Z(n6992) );
  AOI21_X1 U8901 ( .B1(n6983), .B2(n6982), .A(n6981), .ZN(n6984) );
  OAI22_X1 U8902 ( .A1(n8768), .A2(n6984), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7172), .ZN(n6991) );
  OAI21_X1 U8903 ( .B1(n6987), .B2(n6986), .A(n6985), .ZN(n6988) );
  AOI22_X1 U8904 ( .A1(n8728), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n8750), .B2(
        n6988), .ZN(n6989) );
  INV_X1 U8905 ( .A(n6989), .ZN(n6990) );
  AOI211_X1 U8906 ( .C1(n8733), .C2(n6992), .A(n6991), .B(n6990), .ZN(n6993)
         );
  OAI21_X1 U8907 ( .B1(n6994), .B2(n8755), .A(n6993), .ZN(P2_U3184) );
  AOI21_X1 U8908 ( .B1(n10232), .B2(n6996), .A(n6995), .ZN(n6998) );
  OAI22_X1 U8909 ( .A1(n8768), .A2(n6998), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6997), .ZN(n7007) );
  INV_X1 U8910 ( .A(n6999), .ZN(n7000) );
  AOI21_X1 U8911 ( .B1(n7249), .B2(n7001), .A(n7000), .ZN(n7005) );
  XNOR2_X1 U8912 ( .A(n7003), .B(n7002), .ZN(n7004) );
  OAI22_X1 U8913 ( .A1(n8739), .A2(n7005), .B1(n8760), .B2(n7004), .ZN(n7006)
         );
  AOI211_X1 U8914 ( .C1(n8728), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n7007), .B(
        n7006), .ZN(n7008) );
  OAI21_X1 U8915 ( .B1(n7009), .B2(n8755), .A(n7008), .ZN(P2_U3183) );
  AOI21_X1 U8916 ( .B1(n7011), .B2(n7010), .A(n4532), .ZN(n7026) );
  INV_X1 U8917 ( .A(n7012), .ZN(n7016) );
  NAND3_X1 U8918 ( .A1(n7179), .A2(n7014), .A3(n7013), .ZN(n7015) );
  AOI21_X1 U8919 ( .B1(n7016), .B2(n7015), .A(n8768), .ZN(n7024) );
  NAND3_X1 U8920 ( .A1(n7181), .A2(n4538), .A3(n7017), .ZN(n7018) );
  AOI21_X1 U8921 ( .B1(n7019), .B2(n7018), .A(n8739), .ZN(n7023) );
  AND2_X1 U8922 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7423) );
  AOI21_X1 U8923 ( .B1(n8728), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7423), .ZN(
        n7020) );
  OAI21_X1 U8924 ( .B1(n8755), .B2(n7021), .A(n7020), .ZN(n7022) );
  NOR3_X1 U8925 ( .A1(n7024), .A2(n7023), .A3(n7022), .ZN(n7025) );
  OAI21_X1 U8926 ( .B1(n7026), .B2(n8760), .A(n7025), .ZN(P2_U3188) );
  AOI21_X1 U8927 ( .B1(n7028), .B2(n7029), .A(n4432), .ZN(n7053) );
  NAND2_X1 U8928 ( .A1(n9538), .A2(n10269), .ZN(n7052) );
  NAND2_X1 U8929 ( .A1(n7053), .A2(n7052), .ZN(n7118) );
  INV_X1 U8930 ( .A(n9608), .ZN(n9616) );
  XNOR2_X1 U8931 ( .A(n9580), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n9588) );
  XNOR2_X1 U8932 ( .A(n7037), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9570) );
  NAND2_X1 U8933 ( .A1(n10061), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9575) );
  INV_X1 U8934 ( .A(n9575), .ZN(n9569) );
  NAND2_X1 U8935 ( .A1(n9570), .A2(n9569), .ZN(n9568) );
  INV_X1 U8936 ( .A(n7037), .ZN(n9564) );
  NAND2_X1 U8937 ( .A1(n9564), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7031) );
  NAND2_X1 U8938 ( .A1(n9568), .A2(n7031), .ZN(n9587) );
  INV_X1 U8939 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10359) );
  OR2_X1 U8940 ( .A1(n9580), .A2(n10359), .ZN(n7032) );
  NAND2_X1 U8941 ( .A1(n9586), .A2(n7032), .ZN(n9593) );
  INV_X1 U8942 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7952) );
  XNOR2_X1 U8943 ( .A(n9596), .B(n7952), .ZN(n9594) );
  NAND2_X1 U8944 ( .A1(n9593), .A2(n9594), .ZN(n9592) );
  NAND2_X1 U8945 ( .A1(n9596), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7033) );
  XNOR2_X1 U8946 ( .A(n9608), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9607) );
  INV_X1 U8947 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7773) );
  MUX2_X1 U8948 ( .A(n7773), .B(P1_REG2_REG_5__SCAN_IN), .S(n7058), .Z(n7035)
         );
  OR2_X1 U8949 ( .A1(n4437), .A2(n6158), .ZN(n7034) );
  AOI211_X1 U8950 ( .C1(n7036), .C2(n7035), .A(n4454), .B(n10067), .ZN(n7051)
         );
  INV_X1 U8951 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7040) );
  MUX2_X1 U8952 ( .A(n7040), .B(P1_REG1_REG_2__SCAN_IN), .S(n9580), .Z(n9585)
         );
  INV_X1 U8953 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7038) );
  MUX2_X1 U8954 ( .A(n7038), .B(P1_REG1_REG_1__SCAN_IN), .S(n7037), .Z(n9566)
         );
  AND2_X1 U8955 ( .A1(n10061), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9567) );
  NAND2_X1 U8956 ( .A1(n9564), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7039) );
  NAND2_X1 U8957 ( .A1(n9565), .A2(n7039), .ZN(n9584) );
  OR2_X1 U8958 ( .A1(n9580), .A2(n7040), .ZN(n9598) );
  NAND2_X1 U8959 ( .A1(n9599), .A2(n9598), .ZN(n7043) );
  INV_X1 U8960 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7041) );
  MUX2_X1 U8961 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n7041), .S(n9596), .Z(n7042)
         );
  NAND2_X1 U8962 ( .A1(n9596), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9610) );
  INV_X1 U8963 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7044) );
  MUX2_X1 U8964 ( .A(n7044), .B(P1_REG1_REG_4__SCAN_IN), .S(n9608), .Z(n7045)
         );
  NAND2_X1 U8965 ( .A1(n9616), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7048) );
  INV_X1 U8966 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10425) );
  MUX2_X1 U8967 ( .A(n10425), .B(P1_REG1_REG_5__SCAN_IN), .S(n7058), .Z(n7047)
         );
  AND3_X1 U8968 ( .A1(n9613), .A2(n7048), .A3(n7047), .ZN(n7049) );
  NOR3_X1 U8969 ( .A1(n10090), .A2(n7065), .A3(n7049), .ZN(n7050) );
  NOR2_X1 U8970 ( .A1(n7051), .A2(n7050), .ZN(n7057) );
  INV_X1 U8971 ( .A(n7052), .ZN(n7054) );
  NAND2_X1 U8972 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n7508) );
  INV_X1 U8973 ( .A(n7508), .ZN(n7055) );
  AOI21_X1 U8974 ( .B1(n9671), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n7055), .ZN(
        n7056) );
  OAI211_X1 U8975 ( .C1(n7061), .C2(n10088), .A(n7057), .B(n7056), .ZN(
        P1_U3248) );
  AOI21_X1 U8976 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n7058), .A(n4454), .ZN(
        n7060) );
  XNOR2_X1 U8977 ( .A(n7197), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n7059) );
  NOR2_X1 U8978 ( .A1(n7060), .A2(n7059), .ZN(n7190) );
  AOI211_X1 U8979 ( .C1(n7060), .C2(n7059), .A(n10067), .B(n7190), .ZN(n7069)
         );
  NOR2_X1 U8980 ( .A1(n7061), .A2(n10425), .ZN(n7064) );
  INV_X1 U8981 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7062) );
  MUX2_X1 U8982 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n7062), .S(n7197), .Z(n7063)
         );
  INV_X1 U8983 ( .A(n7274), .ZN(n7067) );
  NOR3_X1 U8984 ( .A1(n7065), .A2(n7064), .A3(n7063), .ZN(n7066) );
  NOR3_X1 U8985 ( .A1(n10090), .A2(n7067), .A3(n7066), .ZN(n7068) );
  NOR2_X1 U8986 ( .A1(n7069), .A2(n7068), .ZN(n7071) );
  AND2_X1 U8987 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7576) );
  AOI21_X1 U8988 ( .B1(n9671), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n7576), .ZN(
        n7070) );
  OAI211_X1 U8989 ( .C1(n7072), .C2(n10088), .A(n7071), .B(n7070), .ZN(
        P1_U3249) );
  NAND2_X1 U8990 ( .A1(n7073), .A2(n7076), .ZN(n7074) );
  OAI211_X1 U8991 ( .C1(n7077), .C2(n7076), .A(n7075), .B(n7074), .ZN(n7079)
         );
  INV_X1 U8992 ( .A(n7079), .ZN(n7080) );
  INV_X1 U8993 ( .A(n8928), .ZN(n8805) );
  NAND2_X1 U8994 ( .A1(n7080), .A2(n8805), .ZN(n8873) );
  AOI22_X1 U8995 ( .A1(n10178), .A2(n10188), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n10175), .ZN(n7084) );
  INV_X1 U8996 ( .A(n8620), .ZN(n7167) );
  NOR2_X1 U8997 ( .A1(n7167), .A2(n8881), .ZN(n10187) );
  NAND2_X1 U8998 ( .A1(n8621), .A2(n7141), .ZN(n8454) );
  AND2_X1 U8999 ( .A1(n7142), .A2(n8454), .ZN(n10184) );
  NOR3_X1 U9000 ( .A1(n10184), .A2(n7081), .A3(n10189), .ZN(n7082) );
  OAI21_X1 U9001 ( .B1(n10187), .B2(n7082), .A(n10181), .ZN(n7083) );
  OAI211_X1 U9002 ( .C1(n6185), .C2(n10181), .A(n7084), .B(n7083), .ZN(
        P2_U3233) );
  INV_X1 U9003 ( .A(n7085), .ZN(n7088) );
  OAI222_X1 U9004 ( .A1(n9077), .A2(n7087), .B1(n9090), .B2(n7088), .C1(
        P2_U3151), .C2(n7086), .ZN(P2_U3282) );
  INV_X1 U9005 ( .A(n7653), .ZN(n7529) );
  OAI222_X1 U9006 ( .A1(n10060), .A2(n10442), .B1(n10058), .B2(n7088), .C1(
        P1_U3086), .C2(n7529), .ZN(P1_U3342) );
  OR2_X1 U9007 ( .A1(n7105), .A2(n7089), .ZN(n7099) );
  INV_X1 U9008 ( .A(n7099), .ZN(n7093) );
  NOR2_X1 U9009 ( .A1(n8577), .A2(n10189), .ZN(n7091) );
  AOI21_X1 U9010 ( .B1(n7107), .B2(n7091), .A(n7090), .ZN(n7092) );
  INV_X1 U9011 ( .A(n7108), .ZN(n9073) );
  INV_X1 U9012 ( .A(n7094), .ZN(n7100) );
  AND3_X1 U9013 ( .A1(n7097), .A2(n7096), .A3(n7095), .ZN(n7098) );
  OAI211_X1 U9014 ( .C1(n7100), .C2(n7107), .A(n7099), .B(n7098), .ZN(n7101)
         );
  NAND2_X1 U9015 ( .A1(n7101), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7103) );
  OR2_X1 U9016 ( .A1(n7105), .A2(n7104), .ZN(n7102) );
  NAND2_X1 U9017 ( .A1(n8336), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7241) );
  NAND2_X1 U9018 ( .A1(n7241), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7112) );
  INV_X1 U9019 ( .A(n7104), .ZN(n8590) );
  AND2_X1 U9020 ( .A1(n7105), .A2(n8590), .ZN(n7128) );
  INV_X1 U9021 ( .A(n7128), .ZN(n7106) );
  OR2_X1 U9022 ( .A1(n7107), .A2(n7171), .ZN(n7110) );
  AND2_X1 U9023 ( .A1(n7108), .A2(n10189), .ZN(n7109) );
  AOI22_X1 U9024 ( .A1(n8392), .A2(n8620), .B1(n8375), .B2(n10188), .ZN(n7111)
         );
  OAI211_X1 U9025 ( .C1(n10184), .C2(n8378), .A(n7112), .B(n7111), .ZN(
        P2_U3172) );
  NOR2_X1 U9026 ( .A1(n6158), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7113) );
  OR2_X1 U9027 ( .A1(n4437), .A2(n7113), .ZN(n9576) );
  INV_X1 U9028 ( .A(n9576), .ZN(n7114) );
  OAI21_X1 U9029 ( .B1(n9535), .B2(P1_REG1_REG_0__SCAN_IN), .A(n7114), .ZN(
        n7115) );
  MUX2_X1 U9030 ( .A(n7115), .B(n7114), .S(n10061), .Z(n7117) );
  INV_X1 U9031 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7116) );
  OAI22_X1 U9032 ( .A1(n7118), .A2(n7117), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7116), .ZN(n7120) );
  NOR3_X1 U9033 ( .A1(n10090), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n5071), .ZN(
        n7119) );
  AOI211_X1 U9034 ( .C1(n9671), .C2(P1_ADDR_REG_0__SCAN_IN), .A(n7120), .B(
        n7119), .ZN(n7121) );
  INV_X1 U9035 ( .A(n7121), .ZN(P1_U3243) );
  INV_X1 U9036 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7123) );
  INV_X1 U9037 ( .A(n7122), .ZN(n7125) );
  INV_X1 U9038 ( .A(n8203), .ZN(n8193) );
  OAI222_X1 U9039 ( .A1(n10060), .A2(n7123), .B1(n10058), .B2(n7125), .C1(
        P1_U3086), .C2(n8193), .ZN(P1_U3341) );
  INV_X1 U9040 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7126) );
  OAI222_X1 U9041 ( .A1(n9077), .A2(n7126), .B1(n9090), .B2(n7125), .C1(
        P2_U3151), .C2(n7124), .ZN(P2_U3281) );
  INV_X1 U9042 ( .A(n7241), .ZN(n7149) );
  INV_X1 U9043 ( .A(n6508), .ZN(n7166) );
  OAI22_X1 U9044 ( .A1(n8390), .A2(n7167), .B1(n7166), .B2(n8373), .ZN(n7129)
         );
  AOI21_X1 U9045 ( .B1(n8375), .B2(n6204), .A(n7129), .ZN(n7148) );
  NAND3_X1 U9046 ( .A1(n7131), .A2(n8440), .A3(n7130), .ZN(n7132) );
  NAND2_X1 U9047 ( .A1(n7133), .A2(n7132), .ZN(n7135) );
  NAND2_X1 U9048 ( .A1(n7135), .A2(n7134), .ZN(n7137) );
  XNOR2_X1 U9049 ( .A(n7259), .B(n8619), .ZN(n7145) );
  INV_X1 U9050 ( .A(n7140), .ZN(n7139) );
  NAND2_X1 U9051 ( .A1(n7234), .A2(n7143), .ZN(n7144) );
  OAI21_X1 U9052 ( .B1(n7145), .B2(n7144), .A(n7261), .ZN(n7146) );
  NAND2_X1 U9053 ( .A1(n7146), .A2(n8385), .ZN(n7147) );
  OAI211_X1 U9054 ( .C1(n7149), .C2(n7172), .A(n7148), .B(n7147), .ZN(P2_U3177) );
  AOI21_X1 U9055 ( .B1(n7151), .B2(n7150), .A(n7228), .ZN(n7161) );
  INV_X1 U9056 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10344) );
  OAI21_X1 U9057 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n7152), .A(n7218), .ZN(
        n7153) );
  AOI22_X1 U9058 ( .A1(n5444), .A2(n7153), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3151), .ZN(n7157) );
  OAI21_X1 U9059 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n7154), .A(n7212), .ZN(
        n7155) );
  NAND2_X1 U9060 ( .A1(n8750), .A2(n7155), .ZN(n7156) );
  OAI211_X1 U9061 ( .C1(n10344), .C2(n8759), .A(n7157), .B(n7156), .ZN(n7158)
         );
  AOI21_X1 U9062 ( .B1(n7159), .B2(n8718), .A(n7158), .ZN(n7160) );
  OAI21_X1 U9063 ( .B1(n7161), .B2(n8760), .A(n7160), .ZN(P2_U3185) );
  AND2_X1 U9064 ( .A1(n7171), .A2(n6530), .ZN(n7352) );
  AND2_X1 U9065 ( .A1(n10181), .A2(n7352), .ZN(n10177) );
  INV_X1 U9066 ( .A(n10177), .ZN(n8170) );
  OAI21_X1 U9067 ( .B1(n7162), .B2(n8461), .A(n7164), .ZN(n10197) );
  INV_X1 U9068 ( .A(n10197), .ZN(n7176) );
  XNOR2_X1 U9069 ( .A(n7165), .B(n8461), .ZN(n7170) );
  INV_X1 U9070 ( .A(n7691), .ZN(n10173) );
  OAI22_X1 U9071 ( .A1(n7167), .A2(n8883), .B1(n7166), .B2(n8881), .ZN(n7168)
         );
  AOI21_X1 U9072 ( .B1(n10197), .B2(n10173), .A(n7168), .ZN(n7169) );
  OAI21_X1 U9073 ( .B1(n10185), .B2(n7170), .A(n7169), .ZN(n10195) );
  NAND2_X1 U9074 ( .A1(n6204), .A2(n10189), .ZN(n10194) );
  OAI22_X1 U9075 ( .A1(n8885), .A2(n7172), .B1(n7171), .B2(n10194), .ZN(n7173)
         );
  NOR2_X1 U9076 ( .A1(n10195), .A2(n7173), .ZN(n7174) );
  MUX2_X1 U9077 ( .A(n10558), .B(n7174), .S(n10181), .Z(n7175) );
  OAI21_X1 U9078 ( .B1(n8170), .B2(n7176), .A(n7175), .ZN(P2_U3231) );
  XNOR2_X1 U9079 ( .A(n7178), .B(n7177), .ZN(n7189) );
  INV_X1 U9080 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7186) );
  OAI21_X1 U9081 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n7180), .A(n7179), .ZN(
        n7183) );
  OAI21_X1 U9082 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n4534), .A(n7181), .ZN(
        n7182) );
  AOI22_X1 U9083 ( .A1(n7183), .A2(n5444), .B1(n8750), .B2(n7182), .ZN(n7185)
         );
  NOR2_X1 U9084 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6232), .ZN(n7349) );
  INV_X1 U9085 ( .A(n7349), .ZN(n7184) );
  OAI211_X1 U9086 ( .C1(n7186), .C2(n8759), .A(n7185), .B(n7184), .ZN(n7187)
         );
  AOI21_X1 U9087 ( .B1(n5320), .B2(n8718), .A(n7187), .ZN(n7188) );
  OAI21_X1 U9088 ( .B1(n8760), .B2(n7189), .A(n7188), .ZN(P2_U3187) );
  INV_X1 U9089 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7193) );
  INV_X1 U9090 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7191) );
  MUX2_X1 U9091 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7191), .S(n7198), .Z(n7192)
         );
  INV_X1 U9092 ( .A(n7192), .ZN(n7269) );
  XNOR2_X1 U9093 ( .A(n7286), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n7282) );
  AND2_X1 U9094 ( .A1(n7286), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10065) );
  XNOR2_X1 U9095 ( .A(n7201), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n10064) );
  AOI21_X1 U9096 ( .B1(n7193), .B2(n10073), .A(n10063), .ZN(n7195) );
  XOR2_X1 U9097 ( .A(n7317), .B(P1_REG2_REG_10__SCAN_IN), .Z(n7194) );
  NAND2_X1 U9098 ( .A1(n7195), .A2(n7194), .ZN(n7318) );
  OAI211_X1 U9099 ( .C1(n7195), .C2(n7194), .A(n7318), .B(n10093), .ZN(n7208)
         );
  INV_X1 U9100 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7196) );
  NAND2_X1 U9101 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9110) );
  OAI21_X1 U9102 ( .B1(n10098), .B2(n7196), .A(n9110), .ZN(n7206) );
  XNOR2_X1 U9103 ( .A(n7317), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n7204) );
  NAND2_X1 U9104 ( .A1(n7197), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7273) );
  INV_X1 U9105 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10489) );
  MUX2_X1 U9106 ( .A(n10489), .B(P1_REG1_REG_7__SCAN_IN), .S(n7198), .Z(n7272)
         );
  NOR2_X1 U9107 ( .A1(n7279), .A2(n10489), .ZN(n7285) );
  NAND2_X1 U9108 ( .A1(n7286), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7200) );
  INV_X1 U9109 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7287) );
  NAND2_X1 U9110 ( .A1(n7295), .A2(n7287), .ZN(n7199) );
  NAND2_X1 U9111 ( .A1(n7290), .A2(n7200), .ZN(n10071) );
  XNOR2_X1 U9112 ( .A(n7201), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n10072) );
  NOR2_X1 U9113 ( .A1(n7201), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7202) );
  OR2_X1 U9114 ( .A1(n10070), .A2(n7202), .ZN(n7203) );
  AOI211_X1 U9115 ( .C1(n7204), .C2(n7203), .A(n10090), .B(n7316), .ZN(n7205)
         );
  AOI211_X1 U9116 ( .C1(n9650), .C2(n7317), .A(n7206), .B(n7205), .ZN(n7207)
         );
  NAND2_X1 U9117 ( .A1(n7208), .A2(n7207), .ZN(P1_U3253) );
  INV_X1 U9118 ( .A(n7209), .ZN(n7211) );
  NAND3_X1 U9119 ( .A1(n7212), .A2(n7211), .A3(n7210), .ZN(n7213) );
  NAND2_X1 U9120 ( .A1(n7214), .A2(n7213), .ZN(n7224) );
  INV_X1 U9121 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7215) );
  NOR2_X1 U9122 ( .A1(n8759), .A2(n7215), .ZN(n7223) );
  AND3_X1 U9123 ( .A1(n7218), .A2(n7217), .A3(n7216), .ZN(n7219) );
  OAI21_X1 U9124 ( .B1(n7220), .B2(n7219), .A(n5444), .ZN(n7221) );
  NAND2_X1 U9125 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7310) );
  NAND2_X1 U9126 ( .A1(n7221), .A2(n7310), .ZN(n7222) );
  AOI211_X1 U9127 ( .C1(n8750), .C2(n7224), .A(n7223), .B(n7222), .ZN(n7232)
         );
  INV_X1 U9128 ( .A(n7225), .ZN(n7230) );
  OAI21_X1 U9129 ( .B1(n7228), .B2(n7227), .A(n7226), .ZN(n7229) );
  NAND3_X1 U9130 ( .A1(n7230), .A2(n8733), .A3(n7229), .ZN(n7231) );
  OAI211_X1 U9131 ( .C1(n8755), .C2(n7233), .A(n7232), .B(n7231), .ZN(P2_U3186) );
  INV_X1 U9132 ( .A(n7234), .ZN(n7235) );
  AOI21_X1 U9133 ( .B1(n7237), .B2(n7236), .A(n7235), .ZN(n7243) );
  AOI22_X1 U9134 ( .A1(n8392), .A2(n8619), .B1(n8371), .B2(n8621), .ZN(n7238)
         );
  OAI21_X1 U9135 ( .B1(n7239), .B2(n8395), .A(n7238), .ZN(n7240) );
  AOI21_X1 U9136 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7241), .A(n7240), .ZN(
        n7242) );
  OAI21_X1 U9137 ( .B1(n7243), .B2(n8378), .A(n7242), .ZN(P2_U3162) );
  NOR2_X1 U9138 ( .A1(n9671), .A2(P1_U3973), .ZN(P1_U3085) );
  XNOR2_X1 U9139 ( .A(n7142), .B(n7244), .ZN(n10190) );
  INV_X1 U9140 ( .A(n10190), .ZN(n7252) );
  AOI22_X1 U9141 ( .A1(n10178), .A2(n6191), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n10175), .ZN(n7251) );
  INV_X1 U9142 ( .A(n7244), .ZN(n8413) );
  XNOR2_X1 U9143 ( .A(n8413), .B(n7245), .ZN(n7247) );
  AOI22_X1 U9144 ( .A1(n10167), .A2(n8621), .B1(n8619), .B2(n10168), .ZN(n7246) );
  OAI21_X1 U9145 ( .B1(n7247), .B2(n10185), .A(n7246), .ZN(n7248) );
  AOI21_X1 U9146 ( .B1(n10173), .B2(n10190), .A(n7248), .ZN(n10192) );
  MUX2_X1 U9147 ( .A(n7249), .B(n10192), .S(n10181), .Z(n7250) );
  OAI211_X1 U9148 ( .C1(n7252), .C2(n8170), .A(n7251), .B(n7250), .ZN(P2_U3232) );
  INV_X1 U9149 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n7254) );
  NAND2_X1 U9150 ( .A1(n7808), .A2(P1_U3973), .ZN(n7253) );
  OAI21_X1 U9151 ( .B1(P1_U3973), .B2(n7254), .A(n7253), .ZN(P1_U3554) );
  MUX2_X1 U9152 ( .A(P2_STATE_REG_SCAN_IN), .B(n8336), .S(n10293), .Z(n7257)
         );
  AOI22_X1 U9153 ( .A1(n8392), .A2(n7255), .B1(n8371), .B2(n8619), .ZN(n7256)
         );
  OAI211_X1 U9154 ( .C1(n10201), .C2(n8395), .A(n7257), .B(n7256), .ZN(n7267)
         );
  XNOR2_X1 U9155 ( .A(n7258), .B(n10201), .ZN(n7298) );
  XNOR2_X1 U9156 ( .A(n7298), .B(n6508), .ZN(n7265) );
  NAND2_X1 U9157 ( .A1(n7259), .A2(n6205), .ZN(n7260) );
  INV_X1 U9158 ( .A(n7300), .ZN(n7263) );
  AOI211_X1 U9159 ( .C1(n7265), .C2(n7264), .A(n8378), .B(n7263), .ZN(n7266)
         );
  OR2_X1 U9160 ( .A1(n7267), .A2(n7266), .ZN(P2_U3158) );
  AOI211_X1 U9161 ( .C1(n7270), .C2(n7269), .A(n10067), .B(n7268), .ZN(n7281)
         );
  NAND2_X1 U9162 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n7644) );
  INV_X1 U9163 ( .A(n7644), .ZN(n7271) );
  AOI21_X1 U9164 ( .B1(n9671), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n7271), .ZN(
        n7278) );
  INV_X1 U9165 ( .A(n7292), .ZN(n7276) );
  NAND3_X1 U9166 ( .A1(n7274), .A2(n7273), .A3(n7272), .ZN(n7275) );
  NAND3_X1 U9167 ( .A1(n9663), .A2(n7276), .A3(n7275), .ZN(n7277) );
  OAI211_X1 U9168 ( .C1(n10088), .C2(n7279), .A(n7278), .B(n7277), .ZN(n7280)
         );
  OR2_X1 U9169 ( .A1(n7281), .A2(n7280), .ZN(P1_U3250) );
  AOI211_X1 U9170 ( .C1(n7283), .C2(n7282), .A(n10067), .B(n10066), .ZN(n7297)
         );
  NAND2_X1 U9171 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n7982) );
  INV_X1 U9172 ( .A(n7982), .ZN(n7284) );
  AOI21_X1 U9173 ( .B1(n9671), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n7284), .ZN(
        n7294) );
  INV_X1 U9174 ( .A(n7285), .ZN(n7289) );
  MUX2_X1 U9175 ( .A(n7287), .B(P1_REG1_REG_8__SCAN_IN), .S(n7286), .Z(n7288)
         );
  NAND2_X1 U9176 ( .A1(n7289), .A2(n7288), .ZN(n7291) );
  OAI211_X1 U9177 ( .C1(n7292), .C2(n7291), .A(n9663), .B(n7290), .ZN(n7293)
         );
  OAI211_X1 U9178 ( .C1(n10088), .C2(n7295), .A(n7294), .B(n7293), .ZN(n7296)
         );
  OR2_X1 U9179 ( .A1(n7297), .A2(n7296), .ZN(P1_U3251) );
  NAND2_X1 U9180 ( .A1(n7298), .A2(n6508), .ZN(n7299) );
  NAND2_X1 U9181 ( .A1(n7300), .A2(n7299), .ZN(n7308) );
  XNOR2_X1 U9182 ( .A(n7258), .B(n7309), .ZN(n7303) );
  NAND2_X1 U9183 ( .A1(n7303), .A2(n7302), .ZN(n7343) );
  INV_X1 U9184 ( .A(n7303), .ZN(n7304) );
  NAND2_X1 U9185 ( .A1(n7304), .A2(n7255), .ZN(n7305) );
  NAND2_X1 U9186 ( .A1(n7343), .A2(n7305), .ZN(n7307) );
  AOI21_X1 U9187 ( .B1(n7308), .B2(n7307), .A(n7344), .ZN(n7315) );
  INV_X1 U9188 ( .A(n7428), .ZN(n7313) );
  AOI22_X1 U9189 ( .A1(n8371), .A2(n6508), .B1(n8375), .B2(n7309), .ZN(n7311)
         );
  OAI211_X1 U9190 ( .C1(n7421), .C2(n8373), .A(n7311), .B(n7310), .ZN(n7312)
         );
  AOI21_X1 U9191 ( .B1(n7313), .B2(n8388), .A(n7312), .ZN(n7314) );
  OAI21_X1 U9192 ( .B1(n7315), .B2(n8378), .A(n7314), .ZN(P2_U3170) );
  AOI21_X1 U9193 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n7317), .A(n7316), .ZN(
        n7523) );
  XNOR2_X1 U9194 ( .A(n7517), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n7522) );
  XNOR2_X1 U9195 ( .A(n7523), .B(n7522), .ZN(n7327) );
  INV_X1 U9196 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7320) );
  OAI21_X1 U9197 ( .B1(n7320), .B2(n7319), .A(n7318), .ZN(n7322) );
  XOR2_X1 U9198 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n7517), .Z(n7321) );
  OAI211_X1 U9199 ( .C1(n7322), .C2(n7321), .A(n10081), .B(n10093), .ZN(n7326)
         );
  INV_X1 U9200 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7323) );
  NAND2_X1 U9201 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9248) );
  OAI21_X1 U9202 ( .B1(n10098), .B2(n7323), .A(n9248), .ZN(n7324) );
  AOI21_X1 U9203 ( .B1(n7517), .B2(n9650), .A(n7324), .ZN(n7325) );
  OAI211_X1 U9204 ( .C1(n7327), .C2(n10090), .A(n7326), .B(n7325), .ZN(
        P1_U3254) );
  INV_X1 U9205 ( .A(n7328), .ZN(n7341) );
  AOI22_X1 U9206 ( .A1(n9651), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n7329), .ZN(n7330) );
  OAI21_X1 U9207 ( .B1(n7341), .B2(n10058), .A(n7330), .ZN(P1_U3338) );
  INV_X1 U9208 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7332) );
  INV_X1 U9209 ( .A(n7331), .ZN(n7333) );
  OAI222_X1 U9210 ( .A1(n9077), .A2(n7332), .B1(n9090), .B2(n7333), .C1(
        P2_U3151), .C2(n4915), .ZN(P2_U3280) );
  INV_X1 U9211 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7334) );
  INV_X1 U9212 ( .A(n8205), .ZN(n9628) );
  OAI222_X1 U9213 ( .A1(n10060), .A2(n7334), .B1(n10058), .B2(n7333), .C1(
        P1_U3086), .C2(n9628), .ZN(P1_U3340) );
  NOR2_X1 U9214 ( .A1(n9448), .A2(n9896), .ZN(n7735) );
  INV_X1 U9215 ( .A(n7810), .ZN(n7335) );
  NAND2_X1 U9216 ( .A1(n7808), .A2(n7816), .ZN(n9446) );
  NAND2_X1 U9217 ( .A1(n7335), .A2(n9446), .ZN(n9411) );
  INV_X1 U9218 ( .A(n9411), .ZN(n7738) );
  AOI21_X1 U9219 ( .B1(n9893), .B2(n10143), .A(n7738), .ZN(n7336) );
  AOI211_X1 U9220 ( .C1(n7337), .C2(n7742), .A(n7735), .B(n7336), .ZN(n7340)
         );
  NAND2_X1 U9221 ( .A1(n10159), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7338) );
  OAI21_X1 U9222 ( .B1(n7340), .B2(n10159), .A(n7338), .ZN(P1_U3522) );
  INV_X1 U9223 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10374) );
  NAND2_X1 U9224 ( .A1(n10154), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n7339) );
  OAI21_X1 U9225 ( .B1(n7340), .B2(n10154), .A(n7339), .ZN(P1_U3453) );
  OAI222_X1 U9226 ( .A1(n9077), .A2(n7342), .B1(n9090), .B2(n7341), .C1(
        P2_U3151), .C2(n8731), .ZN(P2_U3278) );
  XNOR2_X1 U9227 ( .A(n7138), .B(n10211), .ZN(n7415) );
  XNOR2_X1 U9228 ( .A(n7415), .B(n7421), .ZN(n7345) );
  NOR3_X1 U9229 ( .A1(n7344), .A2(n5151), .A3(n7345), .ZN(n7347) );
  INV_X1 U9230 ( .A(n7418), .ZN(n7346) );
  OAI21_X1 U9231 ( .B1(n7347), .B2(n7346), .A(n8385), .ZN(n7351) );
  OAI22_X1 U9232 ( .A1(n8395), .A2(n10211), .B1(n7555), .B2(n8373), .ZN(n7348)
         );
  AOI211_X1 U9233 ( .C1(n8371), .C2(n7255), .A(n7349), .B(n7348), .ZN(n7350)
         );
  OAI211_X1 U9234 ( .C1(n10174), .C2(n8336), .A(n7351), .B(n7350), .ZN(
        P2_U3167) );
  INV_X1 U9235 ( .A(n7352), .ZN(n7353) );
  NAND2_X1 U9236 ( .A1(n7691), .A2(n7353), .ZN(n7354) );
  XNOR2_X1 U9237 ( .A(n7356), .B(n7355), .ZN(n10202) );
  INV_X1 U9238 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7359) );
  XNOR2_X1 U9239 ( .A(n7355), .B(n7357), .ZN(n7358) );
  AOI222_X1 U9240 ( .A1(n10171), .A2(n7358), .B1(n7255), .B2(n10168), .C1(
        n8619), .C2(n10167), .ZN(n10200) );
  MUX2_X1 U9241 ( .A(n7359), .B(n10200), .S(n10181), .Z(n7362) );
  AOI22_X1 U9242 ( .A1(n10178), .A2(n7360), .B1(n10175), .B2(n10293), .ZN(
        n7361) );
  OAI211_X1 U9243 ( .C1(n8934), .C2(n10202), .A(n7362), .B(n7361), .ZN(
        P2_U3230) );
  OAI21_X1 U9244 ( .B1(n9410), .B2(n7364), .A(n7363), .ZN(n7830) );
  AOI211_X1 U9245 ( .C1(n6097), .C2(n7815), .A(n9907), .B(n7951), .ZN(n7831)
         );
  XNOR2_X1 U9246 ( .A(n9410), .B(n7365), .ZN(n7366) );
  OAI222_X1 U9247 ( .A1(n9896), .A2(n8129), .B1(n9898), .B2(n9448), .C1(n7366), 
        .C2(n9893), .ZN(n7834) );
  AOI211_X1 U9248 ( .C1(n10136), .C2(n7830), .A(n7831), .B(n7834), .ZN(n7371)
         );
  AOI22_X1 U9249 ( .A1(n7727), .A2(n6097), .B1(n10159), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n7367) );
  OAI21_X1 U9250 ( .B1(n7371), .B2(n10159), .A(n7367), .ZN(P1_U3524) );
  INV_X1 U9251 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7368) );
  OAI22_X1 U9252 ( .A1(n10026), .A2(n8131), .B1(n10155), .B2(n7368), .ZN(n7369) );
  INV_X1 U9253 ( .A(n7369), .ZN(n7370) );
  OAI21_X1 U9254 ( .B1(n7371), .B2(n10154), .A(n7370), .ZN(P1_U3459) );
  INV_X1 U9255 ( .A(n7372), .ZN(n7407) );
  AOI22_X1 U9256 ( .A1(n8717), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n9088), .ZN(n7373) );
  OAI21_X1 U9257 ( .B1(n7407), .B2(n9090), .A(n7373), .ZN(P2_U3279) );
  INV_X1 U9258 ( .A(n8126), .ZN(n7374) );
  AOI21_X1 U9259 ( .B1(n7376), .B2(n7375), .A(n7374), .ZN(n7382) );
  NOR2_X1 U9260 ( .A1(n9174), .A2(P1_U3086), .ZN(n8130) );
  INV_X1 U9261 ( .A(n8130), .ZN(n7412) );
  INV_X1 U9262 ( .A(n7808), .ZN(n7377) );
  OAI22_X1 U9263 ( .A1(n7377), .A2(n9279), .B1(n9250), .B2(n7947), .ZN(n7380)
         );
  NOR2_X1 U9264 ( .A1(n9287), .A2(n7378), .ZN(n7379) );
  AOI211_X1 U9265 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n7412), .A(n7380), .B(
        n7379), .ZN(n7381) );
  OAI21_X1 U9266 ( .B1(n7382), .B2(n9262), .A(n7381), .ZN(P1_U3222) );
  OAI21_X1 U9267 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n4529), .A(n7383), .ZN(
        n7390) );
  NAND2_X1 U9268 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7554) );
  NAND2_X1 U9269 ( .A1(n8728), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7384) );
  OAI211_X1 U9270 ( .C1(n8755), .C2(n7385), .A(n7554), .B(n7384), .ZN(n7389)
         );
  AOI21_X1 U9271 ( .B1(n7563), .B2(n7386), .A(n6910), .ZN(n7387) );
  NOR2_X1 U9272 ( .A1(n7387), .A2(n8768), .ZN(n7388) );
  AOI211_X1 U9273 ( .C1(n8750), .C2(n7390), .A(n7389), .B(n7388), .ZN(n7397)
         );
  INV_X1 U9274 ( .A(n7391), .ZN(n7395) );
  NOR3_X1 U9275 ( .A1(n4532), .A2(n7393), .A3(n7392), .ZN(n7394) );
  OAI21_X1 U9276 ( .B1(n7395), .B2(n7394), .A(n8733), .ZN(n7396) );
  NAND2_X1 U9277 ( .A1(n7397), .A2(n7396), .ZN(P2_U3189) );
  NAND2_X1 U9278 ( .A1(n7398), .A2(n9276), .ZN(n7406) );
  AOI21_X1 U9279 ( .B1(n7472), .B2(n7400), .A(n7399), .ZN(n7405) );
  INV_X1 U9280 ( .A(n7401), .ZN(n10111) );
  AOI22_X1 U9281 ( .A1(n9284), .A2(n9558), .B1(n9267), .B2(n10111), .ZN(n7404)
         );
  INV_X1 U9282 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10548) );
  NOR2_X1 U9283 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10548), .ZN(n9605) );
  NOR2_X1 U9284 ( .A1(n9279), .A2(n8129), .ZN(n7402) );
  AOI211_X1 U9285 ( .C1(n7452), .C2(n9236), .A(n9605), .B(n7402), .ZN(n7403)
         );
  OAI211_X1 U9286 ( .C1(n7406), .C2(n7405), .A(n7404), .B(n7403), .ZN(P1_U3230) );
  INV_X1 U9287 ( .A(n9641), .ZN(n8198) );
  OAI222_X1 U9288 ( .A1(n10060), .A2(n7408), .B1(n10058), .B2(n7407), .C1(
        n8198), .C2(P1_U3086), .ZN(P1_U3339) );
  XOR2_X1 U9289 ( .A(n7410), .B(n7409), .Z(n9574) );
  NAND2_X1 U9290 ( .A1(n9574), .A2(n9276), .ZN(n7414) );
  AOI22_X1 U9291 ( .A1(n7412), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n9284), .B2(
        n7411), .ZN(n7413) );
  OAI211_X1 U9292 ( .C1(n9287), .C2(n7816), .A(n7414), .B(n7413), .ZN(P1_U3232) );
  INV_X1 U9293 ( .A(n7415), .ZN(n7416) );
  NAND2_X1 U9294 ( .A1(n7416), .A2(n7421), .ZN(n7417) );
  XNOR2_X1 U9295 ( .A(n8101), .B(n7461), .ZN(n7546) );
  XNOR2_X1 U9296 ( .A(n7546), .B(n10169), .ZN(n7419) );
  OAI211_X1 U9297 ( .C1(n7420), .C2(n7419), .A(n7548), .B(n8385), .ZN(n7425)
         );
  INV_X1 U9298 ( .A(n7461), .ZN(n10217) );
  OAI22_X1 U9299 ( .A1(n8390), .A2(n7421), .B1(n8395), .B2(n10217), .ZN(n7422)
         );
  AOI211_X1 U9300 ( .C1(n8392), .C2(n8617), .A(n7423), .B(n7422), .ZN(n7424)
         );
  OAI211_X1 U9301 ( .C1(n7459), .C2(n8336), .A(n7425), .B(n7424), .ZN(P2_U3179) );
  INV_X1 U9302 ( .A(n8934), .ZN(n7570) );
  OAI21_X1 U9303 ( .B1(n7427), .B2(n8465), .A(n7426), .ZN(n10208) );
  OAI22_X1 U9304 ( .A1(n8873), .A2(n10205), .B1(n7428), .B2(n8885), .ZN(n7438)
         );
  AND2_X1 U9305 ( .A1(n7430), .A2(n7429), .ZN(n7433) );
  OAI21_X1 U9306 ( .B1(n7433), .B2(n7432), .A(n7431), .ZN(n7434) );
  NAND2_X1 U9307 ( .A1(n7434), .A2(n10171), .ZN(n7436) );
  AOI22_X1 U9308 ( .A1(n10167), .A2(n6508), .B1(n8618), .B2(n10168), .ZN(n7435) );
  NAND2_X1 U9309 ( .A1(n7436), .A2(n7435), .ZN(n10206) );
  MUX2_X1 U9310 ( .A(n10206), .B(P2_REG2_REG_4__SCAN_IN), .S(n10183), .Z(n7437) );
  AOI211_X1 U9311 ( .C1(n7570), .C2(n10208), .A(n7438), .B(n7437), .ZN(n7439)
         );
  INV_X1 U9312 ( .A(n7439), .ZN(P2_U3229) );
  NAND2_X1 U9313 ( .A1(n7363), .A2(n7440), .ZN(n7950) );
  NAND2_X1 U9314 ( .A1(n7950), .A2(n9414), .ZN(n7949) );
  NAND3_X1 U9315 ( .A1(n7949), .A2(n4435), .A3(n7441), .ZN(n7444) );
  NAND2_X1 U9316 ( .A1(n7444), .A2(n7443), .ZN(n10118) );
  INV_X1 U9317 ( .A(n7776), .ZN(n7446) );
  AOI211_X1 U9318 ( .C1(n7452), .C2(n7445), .A(n9907), .B(n7446), .ZN(n10109)
         );
  INV_X1 U9319 ( .A(n7447), .ZN(n7448) );
  XNOR2_X1 U9320 ( .A(n9412), .B(n9296), .ZN(n7449) );
  AOI222_X1 U9321 ( .A1(n9918), .A2(n7449), .B1(n9560), .B2(n9915), .C1(n9558), 
        .C2(n9913), .ZN(n10121) );
  INV_X1 U9322 ( .A(n10121), .ZN(n7450) );
  AOI211_X1 U9323 ( .C1(n10136), .C2(n10118), .A(n10109), .B(n7450), .ZN(n7454) );
  INV_X1 U9324 ( .A(n10026), .ZN(n7725) );
  AOI22_X1 U9325 ( .A1(n7725), .A2(n7452), .B1(n10154), .B2(
        P1_REG0_REG_4__SCAN_IN), .ZN(n7451) );
  OAI21_X1 U9326 ( .B1(n7454), .B2(n10154), .A(n7451), .ZN(P1_U3465) );
  AOI22_X1 U9327 ( .A1(n7727), .A2(n7452), .B1(n10159), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n7453) );
  OAI21_X1 U9328 ( .B1(n7454), .B2(n10159), .A(n7453), .ZN(P1_U3526) );
  AND2_X1 U9329 ( .A1(n4479), .A2(n8491), .ZN(n8418) );
  XOR2_X1 U9330 ( .A(n7455), .B(n8418), .Z(n10218) );
  XOR2_X1 U9331 ( .A(n7456), .B(n8418), .Z(n7457) );
  AOI222_X1 U9332 ( .A1(n10171), .A2(n7457), .B1(n8617), .B2(n10168), .C1(
        n8618), .C2(n10167), .ZN(n10216) );
  MUX2_X1 U9333 ( .A(n7458), .B(n10216), .S(n10181), .Z(n7463) );
  INV_X1 U9334 ( .A(n7459), .ZN(n7460) );
  AOI22_X1 U9335 ( .A1(n10178), .A2(n7461), .B1(n10175), .B2(n7460), .ZN(n7462) );
  OAI211_X1 U9336 ( .C1(n8934), .C2(n10218), .A(n7463), .B(n7462), .ZN(
        P2_U3227) );
  INV_X1 U9337 ( .A(n7464), .ZN(n7466) );
  INV_X1 U9338 ( .A(n7598), .ZN(n7465) );
  AOI21_X1 U9339 ( .B1(n7466), .B2(n8474), .A(n7465), .ZN(n7571) );
  INV_X1 U9340 ( .A(n10198), .ZN(n7467) );
  NAND2_X1 U9341 ( .A1(n7691), .A2(n7467), .ZN(n10213) );
  XNOR2_X1 U9342 ( .A(n7468), .B(n8416), .ZN(n7469) );
  OAI222_X1 U9343 ( .A1(n8881), .A2(n7851), .B1(n8883), .B2(n7555), .C1(n10185), .C2(n7469), .ZN(n7567) );
  AOI21_X1 U9344 ( .B1(n7571), .B2(n10213), .A(n7567), .ZN(n7562) );
  OAI22_X1 U9345 ( .A1(n7566), .A2(n9045), .B1(n10230), .B2(n6260), .ZN(n7470)
         );
  INV_X1 U9346 ( .A(n7470), .ZN(n7471) );
  OAI21_X1 U9347 ( .B1(n7562), .B2(n10229), .A(n7471), .ZN(P2_U3411) );
  OAI21_X1 U9348 ( .B1(n7474), .B2(n7473), .A(n7472), .ZN(n7479) );
  AOI22_X1 U9349 ( .A1(n9284), .A2(n9559), .B1(n9267), .B2(n7475), .ZN(n7477)
         );
  AND2_X1 U9350 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9595) );
  AOI21_X1 U9351 ( .B1(n9247), .B2(n9561), .A(n9595), .ZN(n7476) );
  OAI211_X1 U9352 ( .C1(n10132), .C2(n9287), .A(n7477), .B(n7476), .ZN(n7478)
         );
  AOI21_X1 U9353 ( .B1(n7479), .B2(n9276), .A(n7478), .ZN(n7480) );
  INV_X1 U9354 ( .A(n7480), .ZN(P1_U3218) );
  INV_X1 U9355 ( .A(n7481), .ZN(n7483) );
  INV_X1 U9356 ( .A(n8209), .ZN(n9674) );
  OAI222_X1 U9357 ( .A1(n10060), .A2(n7482), .B1(n10058), .B2(n7483), .C1(
        n9674), .C2(P1_U3086), .ZN(P1_U3337) );
  INV_X1 U9358 ( .A(n8765), .ZN(n7484) );
  OAI222_X1 U9359 ( .A1(P2_U3151), .A2(n7484), .B1(n9090), .B2(n7483), .C1(
        n10411), .C2(n9077), .ZN(P2_U3277) );
  NAND2_X1 U9360 ( .A1(n7443), .A2(n7485), .ZN(n7767) );
  NAND2_X1 U9361 ( .A1(n7767), .A2(n9413), .ZN(n7766) );
  INV_X1 U9362 ( .A(n7491), .ZN(n7487) );
  NAND3_X1 U9363 ( .A1(n7766), .A2(n7487), .A3(n7486), .ZN(n7489) );
  NAND2_X1 U9364 ( .A1(n7489), .A2(n7488), .ZN(n10105) );
  AOI211_X1 U9365 ( .C1(n7497), .C2(n7774), .A(n9907), .B(n7758), .ZN(n10099)
         );
  XNOR2_X1 U9366 ( .A(n7490), .B(n7491), .ZN(n7492) );
  AOI222_X1 U9367 ( .A1(n9918), .A2(n7492), .B1(n9556), .B2(n9913), .C1(n9558), 
        .C2(n9915), .ZN(n10107) );
  INV_X1 U9368 ( .A(n10107), .ZN(n7493) );
  AOI211_X1 U9369 ( .C1(n10136), .C2(n10105), .A(n10099), .B(n7493), .ZN(n7499) );
  INV_X1 U9370 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7494) );
  OAI22_X1 U9371 ( .A1(n10026), .A2(n10103), .B1(n10155), .B2(n7494), .ZN(
        n7495) );
  INV_X1 U9372 ( .A(n7495), .ZN(n7496) );
  OAI21_X1 U9373 ( .B1(n7499), .B2(n10154), .A(n7496), .ZN(P1_U3471) );
  AOI22_X1 U9374 ( .A1(n7727), .A2(n7497), .B1(n10159), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n7498) );
  OAI21_X1 U9375 ( .B1(n7499), .B2(n10159), .A(n7498), .ZN(P1_U3528) );
  INV_X1 U9376 ( .A(n7500), .ZN(n7502) );
  OAI222_X1 U9377 ( .A1(n9077), .A2(n7501), .B1(n9090), .B2(n7502), .C1(
        P2_U3151), .C2(n8587), .ZN(P2_U3276) );
  OAI222_X1 U9378 ( .A1(n10060), .A2(n7503), .B1(n10058), .B2(n7502), .C1(
        n9920), .C2(P1_U3086), .ZN(P1_U3336) );
  NAND2_X1 U9379 ( .A1(n7505), .A2(n7504), .ZN(n7507) );
  XNOR2_X1 U9380 ( .A(n7507), .B(n7506), .ZN(n7513) );
  OAI21_X1 U9381 ( .B1(n9279), .B2(n7948), .A(n7508), .ZN(n7511) );
  INV_X1 U9382 ( .A(n7509), .ZN(n7777) );
  OAI22_X1 U9383 ( .A1(n9282), .A2(n7777), .B1(n9302), .B2(n9250), .ZN(n7510)
         );
  AOI211_X1 U9384 ( .C1(n10139), .C2(n9236), .A(n7511), .B(n7510), .ZN(n7512)
         );
  OAI21_X1 U9385 ( .B1(n7513), .B2(n9262), .A(n7512), .ZN(P1_U3227) );
  INV_X1 U9386 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7514) );
  MUX2_X1 U9387 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n7514), .S(n7653), .Z(n7515)
         );
  INV_X1 U9388 ( .A(n7515), .ZN(n7519) );
  INV_X1 U9389 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7516) );
  XNOR2_X1 U9390 ( .A(n7524), .B(n7516), .ZN(n10083) );
  NAND2_X1 U9391 ( .A1(n7517), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10080) );
  NAND3_X1 U9392 ( .A1(n10081), .A2(n10083), .A3(n10080), .ZN(n10082) );
  OAI21_X1 U9393 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7524), .A(n10082), .ZN(
        n7518) );
  AOI211_X1 U9394 ( .C1(n7519), .C2(n7518), .A(n10067), .B(n7652), .ZN(n7532)
         );
  XNOR2_X1 U9395 ( .A(n7653), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n7527) );
  INV_X1 U9396 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7520) );
  OAI22_X1 U9397 ( .A1(n7523), .A2(n7522), .B1(n7521), .B2(n7520), .ZN(n10086)
         );
  XNOR2_X1 U9398 ( .A(n7524), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n10087) );
  NOR2_X1 U9399 ( .A1(n7524), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7525) );
  OR2_X1 U9400 ( .A1(n10085), .A2(n7525), .ZN(n7526) );
  AOI211_X1 U9401 ( .C1(n7527), .C2(n7526), .A(n10090), .B(n7650), .ZN(n7531)
         );
  NAND2_X1 U9402 ( .A1(n9671), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n7528) );
  NAND2_X1 U9403 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9220) );
  OAI211_X1 U9404 ( .C1(n10088), .C2(n7529), .A(n7528), .B(n9220), .ZN(n7530)
         );
  OR3_X1 U9405 ( .A1(n7532), .A2(n7531), .A3(n7530), .ZN(P1_U3256) );
  INV_X1 U9406 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n8026) );
  AND2_X1 U9407 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7847) );
  INV_X1 U9408 ( .A(n7847), .ZN(n7533) );
  OAI21_X1 U9409 ( .B1(n8759), .B2(n8026), .A(n7533), .ZN(n7539) );
  OR3_X1 U9410 ( .A1(n7536), .A2(n7535), .A3(n7534), .ZN(n7537) );
  AOI21_X1 U9411 ( .B1(n8632), .B2(n7537), .A(n8760), .ZN(n7538) );
  AOI211_X1 U9412 ( .C1(n8718), .C2(n7540), .A(n7539), .B(n7538), .ZN(n7544)
         );
  OAI21_X1 U9413 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n7541), .A(n8640), .ZN(
        n7542) );
  NAND2_X1 U9414 ( .A1(n7542), .A2(n8750), .ZN(n7543) );
  OAI211_X1 U9415 ( .C1(n7545), .C2(n8768), .A(n7544), .B(n7543), .ZN(P2_U3191) );
  OR2_X1 U9416 ( .A1(n7546), .A2(n7555), .ZN(n7547) );
  XNOR2_X1 U9417 ( .A(n8090), .B(n7566), .ZN(n7549) );
  NAND2_X1 U9418 ( .A1(n7549), .A2(n7592), .ZN(n7586) );
  INV_X1 U9419 ( .A(n7549), .ZN(n7550) );
  NAND2_X1 U9420 ( .A1(n7550), .A2(n8617), .ZN(n7551) );
  NAND2_X1 U9421 ( .A1(n7586), .A2(n7551), .ZN(n7552) );
  INV_X1 U9422 ( .A(n7587), .ZN(n7585) );
  AOI21_X1 U9423 ( .B1(n7553), .B2(n7552), .A(n7585), .ZN(n7561) );
  INV_X1 U9424 ( .A(n7554), .ZN(n7557) );
  OAI22_X1 U9425 ( .A1(n8390), .A2(n7555), .B1(n8395), .B2(n7566), .ZN(n7556)
         );
  AOI211_X1 U9426 ( .C1(n8392), .C2(n8616), .A(n7557), .B(n7556), .ZN(n7560)
         );
  INV_X1 U9427 ( .A(n7565), .ZN(n7558) );
  NAND2_X1 U9428 ( .A1(n8388), .A2(n7558), .ZN(n7559) );
  OAI211_X1 U9429 ( .C1(n7561), .C2(n8378), .A(n7560), .B(n7559), .ZN(P2_U3153) );
  MUX2_X1 U9430 ( .A(n7563), .B(n7562), .S(n10245), .Z(n7564) );
  OAI21_X1 U9431 ( .B1(n7566), .B2(n8974), .A(n7564), .ZN(P2_U3466) );
  OAI22_X1 U9432 ( .A1(n8873), .A2(n7566), .B1(n7565), .B2(n8885), .ZN(n7569)
         );
  MUX2_X1 U9433 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7567), .S(n10181), .Z(n7568)
         );
  AOI211_X1 U9434 ( .C1(n7571), .C2(n7570), .A(n7569), .B(n7568), .ZN(n7572)
         );
  INV_X1 U9435 ( .A(n7572), .ZN(P2_U3226) );
  OAI21_X1 U9436 ( .B1(n7575), .B2(n7574), .A(n7573), .ZN(n7580) );
  AOI22_X1 U9437 ( .A1(n9284), .A2(n9556), .B1(n9267), .B2(n10100), .ZN(n7578)
         );
  AOI21_X1 U9438 ( .B1(n9247), .B2(n9558), .A(n7576), .ZN(n7577) );
  OAI211_X1 U9439 ( .C1(n10103), .C2(n9287), .A(n7578), .B(n7577), .ZN(n7579)
         );
  AOI21_X1 U9440 ( .B1(n7580), .B2(n9276), .A(n7579), .ZN(n7581) );
  INV_X1 U9441 ( .A(n7581), .ZN(P1_U3239) );
  NAND2_X1 U9442 ( .A1(n7607), .A2(n10043), .ZN(n7583) );
  OAI211_X1 U9443 ( .C1(n10480), .C2(n10060), .A(n7583), .B(n7582), .ZN(
        P1_U3335) );
  INV_X1 U9444 ( .A(n7586), .ZN(n7584) );
  XNOR2_X1 U9445 ( .A(n7628), .B(n8101), .ZN(n7852) );
  XNOR2_X1 U9446 ( .A(n7852), .B(n8616), .ZN(n7588) );
  NOR3_X1 U9447 ( .A1(n7585), .A2(n7584), .A3(n7588), .ZN(n7591) );
  NAND2_X1 U9448 ( .A1(n7587), .A2(n7586), .ZN(n7589) );
  INV_X1 U9449 ( .A(n7854), .ZN(n7590) );
  OAI21_X1 U9450 ( .B1(n7591), .B2(n7590), .A(n8385), .ZN(n7596) );
  OAI22_X1 U9451 ( .A1(n8390), .A2(n7592), .B1(n8395), .B2(n10224), .ZN(n7593)
         );
  AOI211_X1 U9452 ( .C1(n8392), .C2(n8615), .A(n7594), .B(n7593), .ZN(n7595)
         );
  OAI211_X1 U9453 ( .C1(n7603), .C2(n8336), .A(n7596), .B(n7595), .ZN(P2_U3161) );
  NAND2_X1 U9454 ( .A1(n7598), .A2(n7597), .ZN(n7599) );
  AND2_X1 U9455 ( .A1(n8471), .A2(n8477), .ZN(n8419) );
  XNOR2_X1 U9456 ( .A(n7599), .B(n8419), .ZN(n10226) );
  INV_X1 U9457 ( .A(n7600), .ZN(n7629) );
  XNOR2_X1 U9458 ( .A(n7629), .B(n8419), .ZN(n7601) );
  AOI222_X1 U9459 ( .A1(n10171), .A2(n7601), .B1(n8615), .B2(n10168), .C1(
        n8617), .C2(n10167), .ZN(n10222) );
  MUX2_X1 U9460 ( .A(n7602), .B(n10222), .S(n10181), .Z(n7606) );
  INV_X1 U9461 ( .A(n7603), .ZN(n7604) );
  AOI22_X1 U9462 ( .A1(n10178), .A2(n7628), .B1(n10175), .B2(n7604), .ZN(n7605) );
  OAI211_X1 U9463 ( .C1(n10226), .C2(n8934), .A(n7606), .B(n7605), .ZN(
        P2_U3225) );
  INV_X1 U9464 ( .A(n7607), .ZN(n7609) );
  OAI222_X1 U9465 ( .A1(P2_U3151), .A2(n8585), .B1(n9090), .B2(n7609), .C1(
        n7608), .C2(n9077), .ZN(P2_U3275) );
  INV_X1 U9466 ( .A(n10151), .ZN(n10128) );
  OAI21_X1 U9467 ( .B1(n7611), .B2(n7615), .A(n7610), .ZN(n7620) );
  INV_X1 U9468 ( .A(n4450), .ZN(n7663) );
  AOI211_X1 U9469 ( .C1(n7986), .C2(n7612), .A(n9907), .B(n7663), .ZN(n7785)
         );
  INV_X1 U9470 ( .A(n7620), .ZN(n7788) );
  INV_X1 U9471 ( .A(n9415), .ZN(n7613) );
  OR2_X1 U9472 ( .A1(n7490), .A2(n7613), .ZN(n7614) );
  NAND2_X1 U9473 ( .A1(n7614), .A2(n9293), .ZN(n7750) );
  INV_X1 U9474 ( .A(n9299), .ZN(n7751) );
  NAND2_X1 U9475 ( .A1(n7750), .A2(n7751), .ZN(n7749) );
  AOI21_X1 U9476 ( .B1(n7749), .B2(n7616), .A(n7615), .ZN(n7666) );
  AND3_X1 U9477 ( .A1(n7749), .A2(n7616), .A3(n7615), .ZN(n7617) );
  OAI21_X1 U9478 ( .B1(n7666), .B2(n7617), .A(n9918), .ZN(n7619) );
  AOI22_X1 U9479 ( .A1(n9915), .A2(n9556), .B1(n9554), .B2(n9913), .ZN(n7618)
         );
  OAI211_X1 U9480 ( .C1(n7788), .C2(n7814), .A(n7619), .B(n7618), .ZN(n7781)
         );
  AOI211_X1 U9481 ( .C1(n10128), .C2(n7620), .A(n7785), .B(n7781), .ZN(n7625)
         );
  AOI22_X1 U9482 ( .A1(n7727), .A2(n7986), .B1(n10159), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n7621) );
  OAI21_X1 U9483 ( .B1(n7625), .B2(n10159), .A(n7621), .ZN(P1_U3530) );
  INV_X1 U9484 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7622) );
  OAI22_X1 U9485 ( .A1(n10026), .A2(n7783), .B1(n10155), .B2(n7622), .ZN(n7623) );
  INV_X1 U9486 ( .A(n7623), .ZN(n7624) );
  OAI21_X1 U9487 ( .B1(n7625), .B2(n10154), .A(n7624), .ZN(P1_U3477) );
  XNOR2_X1 U9488 ( .A(n7626), .B(n8422), .ZN(n7683) );
  INV_X1 U9489 ( .A(n7683), .ZN(n7634) );
  AOI21_X1 U9490 ( .B1(n7600), .B2(n10224), .A(n7851), .ZN(n7627) );
  AOI21_X1 U9491 ( .B1(n7629), .B2(n7628), .A(n7627), .ZN(n7630) );
  XNOR2_X1 U9492 ( .A(n7630), .B(n8422), .ZN(n7631) );
  NAND2_X1 U9493 ( .A1(n7631), .A2(n10171), .ZN(n7633) );
  AOI22_X1 U9494 ( .A1(n8616), .A2(n10167), .B1(n10168), .B2(n8614), .ZN(n7632) );
  OAI211_X1 U9495 ( .C1(n7683), .C2(n7691), .A(n7633), .B(n7632), .ZN(n7677)
         );
  AOI21_X1 U9496 ( .B1(n10198), .B2(n7634), .A(n7677), .ZN(n7694) );
  INV_X1 U9497 ( .A(n4644), .ZN(n7696) );
  INV_X1 U9498 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7635) );
  OAI22_X1 U9499 ( .A1(n7696), .A2(n9045), .B1(n10230), .B2(n7635), .ZN(n7636)
         );
  INV_X1 U9500 ( .A(n7636), .ZN(n7637) );
  OAI21_X1 U9501 ( .B1(n7694), .B2(n10229), .A(n7637), .ZN(P2_U3417) );
  INV_X1 U9502 ( .A(n7638), .ZN(n7642) );
  OAI21_X1 U9503 ( .B1(n7642), .B2(n7640), .A(n7639), .ZN(n7641) );
  OAI211_X1 U9504 ( .C1(n7643), .C2(n7642), .A(n9276), .B(n7641), .ZN(n7649)
         );
  OAI21_X1 U9505 ( .B1(n9279), .B2(n9302), .A(n7644), .ZN(n7647) );
  INV_X1 U9506 ( .A(n7645), .ZN(n7761) );
  OAI22_X1 U9507 ( .A1(n9282), .A2(n7761), .B1(n9202), .B2(n9250), .ZN(n7646)
         );
  AOI211_X1 U9508 ( .C1(n10147), .C2(n9223), .A(n7647), .B(n7646), .ZN(n7648)
         );
  NAND2_X1 U9509 ( .A1(n7649), .A2(n7648), .ZN(P1_U3213) );
  XNOR2_X1 U9510 ( .A(n8203), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n8190) );
  XOR2_X1 U9511 ( .A(n8190), .B(n8191), .Z(n7659) );
  NAND2_X1 U9512 ( .A1(n9671), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n7651) );
  NAND2_X1 U9513 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9095) );
  OAI211_X1 U9514 ( .C1(n10088), .C2(n8193), .A(n7651), .B(n9095), .ZN(n7658)
         );
  NAND2_X1 U9515 ( .A1(n8203), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7654) );
  OAI21_X1 U9516 ( .B1(n8203), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7654), .ZN(
        n7655) );
  AOI211_X1 U9517 ( .C1(n7656), .C2(n7655), .A(n10067), .B(n8202), .ZN(n7657)
         );
  AOI211_X1 U9518 ( .C1(n9663), .C2(n7659), .A(n7658), .B(n7657), .ZN(n7660)
         );
  INV_X1 U9519 ( .A(n7660), .ZN(P1_U3257) );
  OAI21_X1 U9520 ( .B1(n7662), .B2(n7668), .A(n7661), .ZN(n7827) );
  OAI21_X1 U9521 ( .B1(n7663), .B2(n4623), .A(n9976), .ZN(n7664) );
  OAI22_X1 U9522 ( .A1(n7664), .A2(n7707), .B1(n7724), .B2(n9896), .ZN(n7823)
         );
  INV_X1 U9523 ( .A(n9319), .ZN(n7665) );
  NOR2_X1 U9524 ( .A1(n7666), .A2(n7665), .ZN(n7667) );
  XOR2_X1 U9525 ( .A(n7668), .B(n7667), .Z(n7669) );
  OAI22_X1 U9526 ( .A1(n7669), .A2(n9893), .B1(n9202), .B2(n9898), .ZN(n7822)
         );
  AOI211_X1 U9527 ( .C1(n10136), .C2(n7827), .A(n7823), .B(n7822), .ZN(n7672)
         );
  AOI22_X1 U9528 ( .A1(n7725), .A2(n4572), .B1(P1_REG0_REG_9__SCAN_IN), .B2(
        n10154), .ZN(n7670) );
  OAI21_X1 U9529 ( .B1(n7672), .B2(n10154), .A(n7670), .ZN(P1_U3480) );
  AOI22_X1 U9530 ( .A1(n7727), .A2(n4572), .B1(n10159), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7671) );
  OAI21_X1 U9531 ( .B1(n7672), .B2(n10159), .A(n7671), .ZN(P1_U3531) );
  INV_X1 U9532 ( .A(n7673), .ZN(n7676) );
  OAI222_X1 U9533 ( .A1(P1_U3086), .A2(n7674), .B1(n10058), .B2(n7676), .C1(
        n10416), .C2(n10060), .ZN(P1_U3334) );
  OAI222_X1 U9534 ( .A1(P2_U3151), .A2(n7130), .B1(n9090), .B2(n7676), .C1(
        n7675), .C2(n9077), .ZN(P2_U3274) );
  INV_X1 U9535 ( .A(n7677), .ZN(n7678) );
  MUX2_X1 U9536 ( .A(n7679), .B(n7678), .S(n10181), .Z(n7682) );
  INV_X1 U9537 ( .A(n7680), .ZN(n7846) );
  AOI22_X1 U9538 ( .A1(n10178), .A2(n4644), .B1(n10175), .B2(n7846), .ZN(n7681) );
  OAI211_X1 U9539 ( .C1(n7683), .C2(n8170), .A(n7682), .B(n7681), .ZN(P2_U3224) );
  XOR2_X1 U9540 ( .A(n7684), .B(n8423), .Z(n8171) );
  INV_X1 U9541 ( .A(n8171), .ZN(n7692) );
  NAND2_X1 U9542 ( .A1(n7686), .A2(n7685), .ZN(n7687) );
  XNOR2_X1 U9543 ( .A(n7687), .B(n8423), .ZN(n7689) );
  OAI22_X1 U9544 ( .A1(n8296), .A2(n8881), .B1(n7850), .B2(n8883), .ZN(n7688)
         );
  AOI21_X1 U9545 ( .B1(n7689), .B2(n10171), .A(n7688), .ZN(n7690) );
  OAI21_X1 U9546 ( .B1(n8171), .B2(n7691), .A(n7690), .ZN(n8162) );
  AOI21_X1 U9547 ( .B1(n10198), .B2(n7692), .A(n8162), .ZN(n7838) );
  AOI22_X1 U9548 ( .A1(n9066), .A2(n8167), .B1(P2_REG0_REG_10__SCAN_IN), .B2(
        n10229), .ZN(n7693) );
  OAI21_X1 U9549 ( .B1(n7838), .B2(n10229), .A(n7693), .ZN(P2_U3420) );
  MUX2_X1 U9550 ( .A(n10500), .B(n7694), .S(n10245), .Z(n7695) );
  OAI21_X1 U9551 ( .B1(n7696), .B2(n8974), .A(n7695), .ZN(P2_U3468) );
  XNOR2_X1 U9552 ( .A(n7697), .B(n5129), .ZN(n8990) );
  XNOR2_X1 U9553 ( .A(n7698), .B(n8411), .ZN(n7699) );
  OAI222_X1 U9554 ( .A1(n8881), .A2(n8363), .B1(n8883), .B2(n8288), .C1(n7699), 
        .C2(n10185), .ZN(n8987) );
  INV_X1 U9555 ( .A(n8987), .ZN(n7700) );
  MUX2_X1 U9556 ( .A(n7701), .B(n7700), .S(n10181), .Z(n7703) );
  AOI22_X1 U9557 ( .A1(n10178), .A2(n8988), .B1(n10175), .B2(n8365), .ZN(n7702) );
  OAI211_X1 U9558 ( .C1(n8990), .C2(n8934), .A(n7703), .B(n7702), .ZN(P2_U3222) );
  OAI21_X1 U9559 ( .B1(n7705), .B2(n9419), .A(n7704), .ZN(n7929) );
  NOR2_X1 U9560 ( .A1(n7707), .A2(n7709), .ZN(n7708) );
  OR2_X1 U9561 ( .A1(n7706), .A2(n7708), .ZN(n7927) );
  INV_X1 U9562 ( .A(n10148), .ZN(n10131) );
  OAI22_X1 U9563 ( .A1(n7927), .A2(n9907), .B1(n7709), .B2(n10131), .ZN(n7715)
         );
  INV_X1 U9564 ( .A(n7710), .ZN(n7711) );
  AOI21_X1 U9565 ( .B1(n9419), .B2(n7712), .A(n7711), .ZN(n7713) );
  OAI222_X1 U9566 ( .A1(n9898), .A2(n7714), .B1(n9896), .B2(n9325), .C1(n9893), 
        .C2(n7713), .ZN(n7923) );
  AOI211_X1 U9567 ( .C1(n10136), .C2(n7929), .A(n7715), .B(n7923), .ZN(n7718)
         );
  NAND2_X1 U9568 ( .A1(n10154), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7716) );
  OAI21_X1 U9569 ( .B1(n7718), .B2(n10154), .A(n7716), .ZN(P1_U3483) );
  NAND2_X1 U9570 ( .A1(n10159), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7717) );
  OAI21_X1 U9571 ( .B1(n7718), .B2(n10159), .A(n7717), .ZN(P1_U3532) );
  XOR2_X1 U9572 ( .A(n7719), .B(n9422), .Z(n7794) );
  OR2_X1 U9573 ( .A1(n7706), .A2(n4994), .ZN(n7721) );
  AND3_X1 U9574 ( .A1(n7720), .A2(n7721), .A3(n9976), .ZN(n7790) );
  XOR2_X1 U9575 ( .A(n7722), .B(n9422), .Z(n7723) );
  OAI222_X1 U9576 ( .A1(n9896), .A2(n9251), .B1(n9898), .B2(n7724), .C1(n9893), 
        .C2(n7723), .ZN(n7789) );
  AOI211_X1 U9577 ( .C1(n7794), .C2(n10136), .A(n7790), .B(n7789), .ZN(n7729)
         );
  AOI22_X1 U9578 ( .A1(n9326), .A2(n7725), .B1(P1_REG0_REG_11__SCAN_IN), .B2(
        n10154), .ZN(n7726) );
  OAI21_X1 U9579 ( .B1(n7729), .B2(n10154), .A(n7726), .ZN(P1_U3486) );
  AOI22_X1 U9580 ( .A1(n9326), .A2(n7727), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n10159), .ZN(n7728) );
  OAI21_X1 U9581 ( .B1(n7729), .B2(n10159), .A(n7728), .ZN(P1_U3533) );
  INV_X1 U9582 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7745) );
  INV_X1 U9583 ( .A(n7730), .ZN(n7734) );
  NOR2_X1 U9584 ( .A1(n7732), .A2(n7731), .ZN(n7733) );
  NAND2_X1 U9585 ( .A1(n7734), .A2(n7733), .ZN(n7741) );
  AOI21_X1 U9586 ( .B1(n10110), .B2(P1_REG3_REG_0__SCAN_IN), .A(n7735), .ZN(
        n7736) );
  OAI21_X1 U9587 ( .B1(n7738), .B2(n7737), .A(n7736), .ZN(n7739) );
  NAND2_X1 U9588 ( .A1(n7739), .A2(n9776), .ZN(n7744) );
  OR2_X1 U9589 ( .A1(n7741), .A2(n9511), .ZN(n9876) );
  NOR2_X1 U9590 ( .A1(n9876), .A2(n9907), .ZN(n9844) );
  OAI21_X1 U9591 ( .B1(n9929), .B2(n9844), .A(n7742), .ZN(n7743) );
  OAI211_X1 U9592 ( .C1(n7745), .C2(n9776), .A(n7744), .B(n7743), .ZN(P1_U3293) );
  OR2_X1 U9593 ( .A1(n7746), .A2(n9299), .ZN(n7747) );
  NAND2_X1 U9594 ( .A1(n7748), .A2(n7747), .ZN(n7753) );
  INV_X1 U9595 ( .A(n7753), .ZN(n10152) );
  OR2_X1 U9596 ( .A1(n10112), .A2(n7769), .ZN(n7821) );
  OAI21_X1 U9597 ( .B1(n7751), .B2(n7750), .A(n7749), .ZN(n7757) );
  INV_X1 U9598 ( .A(n7814), .ZN(n7752) );
  NAND2_X1 U9599 ( .A1(n7753), .A2(n7752), .ZN(n7755) );
  AOI22_X1 U9600 ( .A1(n9557), .A2(n9915), .B1(n9913), .B2(n9555), .ZN(n7754)
         );
  NAND2_X1 U9601 ( .A1(n7755), .A2(n7754), .ZN(n7756) );
  AOI21_X1 U9602 ( .B1(n7757), .B2(n9918), .A(n7756), .ZN(n10150) );
  MUX2_X1 U9603 ( .A(n7191), .B(n10150), .S(n9776), .Z(n7765) );
  INV_X1 U9604 ( .A(n7758), .ZN(n7760) );
  INV_X1 U9605 ( .A(n7612), .ZN(n7759) );
  AOI211_X1 U9606 ( .C1(n10147), .C2(n7760), .A(n9907), .B(n7759), .ZN(n10146)
         );
  OAI22_X1 U9607 ( .A1(n10115), .A2(n7762), .B1(n9922), .B2(n7761), .ZN(n7763)
         );
  AOI21_X1 U9608 ( .B1(n10146), .B2(n10108), .A(n7763), .ZN(n7764) );
  OAI211_X1 U9609 ( .C1(n10152), .C2(n7821), .A(n7765), .B(n7764), .ZN(
        P1_U3286) );
  OAI21_X1 U9610 ( .B1(n7767), .B2(n9413), .A(n7766), .ZN(n7768) );
  INV_X1 U9611 ( .A(n7768), .ZN(n10142) );
  AND2_X1 U9612 ( .A1(n7814), .A2(n7769), .ZN(n7770) );
  XNOR2_X1 U9613 ( .A(n7771), .B(n9413), .ZN(n7772) );
  AOI222_X1 U9614 ( .A1(n9918), .A2(n7772), .B1(n9559), .B2(n9915), .C1(n9557), 
        .C2(n9913), .ZN(n10141) );
  MUX2_X1 U9615 ( .A(n7773), .B(n10141), .S(n9776), .Z(n7780) );
  INV_X1 U9616 ( .A(n7774), .ZN(n7775) );
  AOI211_X1 U9617 ( .C1(n10139), .C2(n7776), .A(n9907), .B(n7775), .ZN(n10138)
         );
  OAI22_X1 U9618 ( .A1(n10115), .A2(n9304), .B1(n9922), .B2(n7777), .ZN(n7778)
         );
  AOI21_X1 U9619 ( .B1(n10138), .B2(n10108), .A(n7778), .ZN(n7779) );
  OAI211_X1 U9620 ( .C1(n10142), .C2(n9926), .A(n7780), .B(n7779), .ZN(
        P1_U3288) );
  NAND2_X1 U9621 ( .A1(n7781), .A2(n9776), .ZN(n7787) );
  AOI22_X1 U9622 ( .A1(n10112), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7981), .B2(
        n10110), .ZN(n7782) );
  OAI21_X1 U9623 ( .B1(n10115), .B2(n7783), .A(n7782), .ZN(n7784) );
  AOI21_X1 U9624 ( .B1(n7785), .B2(n10108), .A(n7784), .ZN(n7786) );
  OAI211_X1 U9625 ( .C1(n7788), .C2(n7821), .A(n7787), .B(n7786), .ZN(P1_U3285) );
  INV_X1 U9626 ( .A(n7789), .ZN(n7796) );
  NAND2_X1 U9627 ( .A1(n7790), .A2(n10108), .ZN(n7792) );
  AOI22_X1 U9628 ( .A1(n10112), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9246), .B2(
        n10110), .ZN(n7791) );
  OAI211_X1 U9629 ( .C1(n4994), .C2(n10115), .A(n7792), .B(n7791), .ZN(n7793)
         );
  AOI21_X1 U9630 ( .B1(n7794), .B2(n10119), .A(n7793), .ZN(n7795) );
  OAI21_X1 U9631 ( .B1(n7796), .B2(n10112), .A(n7795), .ZN(P1_U3282) );
  OAI21_X1 U9632 ( .B1(n7798), .B2(n8412), .A(n7797), .ZN(n7959) );
  XOR2_X1 U9633 ( .A(n7799), .B(n8412), .Z(n7800) );
  OAI222_X1 U9634 ( .A1(n8881), .A2(n7801), .B1(n8883), .B2(n8296), .C1(n7800), 
        .C2(n10185), .ZN(n7960) );
  NAND2_X1 U9635 ( .A1(n7960), .A2(n10181), .ZN(n7806) );
  INV_X1 U9636 ( .A(n8292), .ZN(n7802) );
  OAI22_X1 U9637 ( .A1(n10181), .A2(n7803), .B1(n7802), .B2(n8885), .ZN(n7804)
         );
  AOI21_X1 U9638 ( .B1(n8298), .B2(n10178), .A(n7804), .ZN(n7805) );
  OAI211_X1 U9639 ( .C1(n7959), .C2(n8934), .A(n7806), .B(n7805), .ZN(P2_U3221) );
  XNOR2_X1 U9640 ( .A(n9416), .B(n7807), .ZN(n10123) );
  AOI22_X1 U9641 ( .A1(n9915), .A2(n7808), .B1(n9561), .B2(n9913), .ZN(n7813)
         );
  OAI21_X1 U9642 ( .B1(n7810), .B2(n9416), .A(n7809), .ZN(n7811) );
  NAND2_X1 U9643 ( .A1(n7811), .A2(n9918), .ZN(n7812) );
  OAI211_X1 U9644 ( .C1(n10123), .C2(n7814), .A(n7813), .B(n7812), .ZN(n10125)
         );
  NAND2_X1 U9645 ( .A1(n10125), .A2(n9776), .ZN(n7820) );
  OAI211_X1 U9646 ( .C1(n7378), .C2(n7816), .A(n9976), .B(n7815), .ZN(n10124)
         );
  INV_X1 U9647 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U9648 ( .A1(n10112), .A2(P1_REG2_REG_1__SCAN_IN), .B1(n10110), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7817) );
  OAI21_X1 U9649 ( .B1(n9876), .B2(n10124), .A(n7817), .ZN(n7818) );
  AOI21_X1 U9650 ( .B1(n9929), .B2(n6601), .A(n7818), .ZN(n7819) );
  OAI211_X1 U9651 ( .C1(n10123), .C2(n7821), .A(n7820), .B(n7819), .ZN(
        P1_U3292) );
  INV_X1 U9652 ( .A(n7822), .ZN(n7829) );
  NAND2_X1 U9653 ( .A1(n7823), .A2(n10108), .ZN(n7825) );
  AOI22_X1 U9654 ( .A1(n10112), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n9200), .B2(
        n10110), .ZN(n7824) );
  OAI211_X1 U9655 ( .C1(n4623), .C2(n10115), .A(n7825), .B(n7824), .ZN(n7826)
         );
  AOI21_X1 U9656 ( .B1(n10119), .B2(n7827), .A(n7826), .ZN(n7828) );
  OAI21_X1 U9657 ( .B1(n7829), .B2(n10112), .A(n7828), .ZN(P1_U3284) );
  INV_X1 U9658 ( .A(n7830), .ZN(n7837) );
  INV_X1 U9659 ( .A(n7831), .ZN(n7832) );
  INV_X1 U9660 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9581) );
  OAI22_X1 U9661 ( .A1(n7832), .A2(n9511), .B1(n9922), .B2(n9581), .ZN(n7833)
         );
  OAI21_X1 U9662 ( .B1(n7834), .B2(n7833), .A(n9776), .ZN(n7836) );
  AOI22_X1 U9663 ( .A1(n9929), .A2(n6097), .B1(n10112), .B2(
        P1_REG2_REG_2__SCAN_IN), .ZN(n7835) );
  OAI211_X1 U9664 ( .C1(n7837), .C2(n9926), .A(n7836), .B(n7835), .ZN(P1_U3291) );
  MUX2_X1 U9665 ( .A(n10545), .B(n7838), .S(n10245), .Z(n7839) );
  OAI21_X1 U9666 ( .B1(n7892), .B2(n8974), .A(n7839), .ZN(P2_U3469) );
  INV_X1 U9667 ( .A(n7840), .ZN(n7844) );
  OAI222_X1 U9668 ( .A1(n9077), .A2(n7842), .B1(n9090), .B2(n7844), .C1(
        P2_U3151), .C2(n7841), .ZN(P2_U3273) );
  OAI222_X1 U9669 ( .A1(n10060), .A2(n7845), .B1(n10058), .B2(n7844), .C1(
        n7843), .C2(P1_U3086), .ZN(P1_U3333) );
  NAND2_X1 U9670 ( .A1(n8388), .A2(n7846), .ZN(n7849) );
  AOI21_X1 U9671 ( .B1(n8392), .B2(n8614), .A(n7847), .ZN(n7848) );
  OAI211_X1 U9672 ( .C1(n8390), .C2(n7851), .A(n7849), .B(n7848), .ZN(n7858)
         );
  XNOR2_X1 U9673 ( .A(n4644), .B(n8101), .ZN(n7889) );
  XNOR2_X1 U9674 ( .A(n7889), .B(n7850), .ZN(n7856) );
  NAND2_X1 U9675 ( .A1(n7852), .A2(n7851), .ZN(n7853) );
  AOI211_X1 U9676 ( .C1(n7856), .C2(n7855), .A(n8378), .B(n4439), .ZN(n7857)
         );
  AOI211_X1 U9677 ( .C1(n8375), .C2(n4644), .A(n7858), .B(n7857), .ZN(n7860)
         );
  INV_X1 U9678 ( .A(n7860), .ZN(P2_U3171) );
  XNOR2_X1 U9679 ( .A(n7861), .B(n9407), .ZN(n7942) );
  INV_X1 U9680 ( .A(n7862), .ZN(n9910) );
  AOI211_X1 U9681 ( .C1(n9407), .C2(n7863), .A(n9893), .B(n9910), .ZN(n7865)
         );
  OAI22_X1 U9682 ( .A1(n9325), .A2(n9898), .B1(n9899), .B2(n9896), .ZN(n7864)
         );
  NOR2_X1 U9683 ( .A1(n7865), .A2(n7864), .ZN(n7944) );
  AOI21_X1 U9684 ( .B1(n7720), .B2(n9145), .A(n9907), .ZN(n7866) );
  OR2_X1 U9685 ( .A1(n7720), .A2(n9145), .ZN(n9908) );
  NAND2_X1 U9686 ( .A1(n7866), .A2(n9908), .ZN(n7940) );
  OAI211_X1 U9687 ( .C1(n7867), .C2(n10131), .A(n7944), .B(n7940), .ZN(n7868)
         );
  AOI21_X1 U9688 ( .B1(n10136), .B2(n7942), .A(n7868), .ZN(n7871) );
  NAND2_X1 U9689 ( .A1(n10154), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7869) );
  OAI21_X1 U9690 ( .B1(n7871), .B2(n10154), .A(n7869), .ZN(P1_U3489) );
  NAND2_X1 U9691 ( .A1(n10159), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7870) );
  OAI21_X1 U9692 ( .B1(n7871), .B2(n10159), .A(n7870), .ZN(P1_U3534) );
  AOI21_X1 U9693 ( .B1(n10547), .B2(n7873), .A(n7872), .ZN(n7886) );
  INV_X1 U9694 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7874) );
  NAND2_X1 U9695 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8361) );
  OAI21_X1 U9696 ( .B1(n8759), .B2(n7874), .A(n8361), .ZN(n7880) );
  OR3_X1 U9697 ( .A1(n8629), .A2(n7876), .A3(n7875), .ZN(n7877) );
  AOI21_X1 U9698 ( .B1(n7878), .B2(n7877), .A(n8760), .ZN(n7879) );
  AOI211_X1 U9699 ( .C1(n8718), .C2(n7881), .A(n7880), .B(n7879), .ZN(n7885)
         );
  OAI21_X1 U9700 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n4525), .A(n7882), .ZN(
        n7883) );
  NAND2_X1 U9701 ( .A1(n7883), .A2(n8750), .ZN(n7884) );
  OAI211_X1 U9702 ( .C1(n7886), .C2(n8768), .A(n7885), .B(n7884), .ZN(P2_U3193) );
  INV_X1 U9703 ( .A(n7913), .ZN(n7917) );
  XNOR2_X1 U9704 ( .A(n7913), .B(n8090), .ZN(n7887) );
  NOR2_X1 U9705 ( .A1(n7887), .A2(n8925), .ZN(n7989) );
  AOI21_X1 U9706 ( .B1(n7887), .B2(n8925), .A(n7989), .ZN(n7900) );
  XNOR2_X1 U9707 ( .A(n7966), .B(n8101), .ZN(n7895) );
  INV_X1 U9708 ( .A(n7895), .ZN(n7888) );
  XNOR2_X1 U9709 ( .A(n8411), .B(n8101), .ZN(n8359) );
  XNOR2_X1 U9710 ( .A(n7892), .B(n8101), .ZN(n8003) );
  NAND2_X1 U9711 ( .A1(n8003), .A2(n8614), .ZN(n7891) );
  INV_X1 U9712 ( .A(n7889), .ZN(n7890) );
  NAND2_X1 U9713 ( .A1(n7890), .A2(n8615), .ZN(n8000) );
  NAND3_X1 U9714 ( .A1(n7892), .A2(n8288), .A3(n8090), .ZN(n7893) );
  OAI211_X1 U9715 ( .C1(n8090), .C2(n8613), .A(n5129), .B(n7893), .ZN(n7897)
         );
  NAND3_X1 U9716 ( .A1(n8167), .A2(n8288), .A3(n8101), .ZN(n7894) );
  OAI211_X1 U9717 ( .C1(n8613), .C2(n8101), .A(n8411), .B(n7894), .ZN(n7896)
         );
  XNOR2_X1 U9718 ( .A(n7895), .B(n8612), .ZN(n8291) );
  AOI21_X1 U9719 ( .B1(n7897), .B2(n7896), .A(n8291), .ZN(n7898) );
  NAND2_X1 U9720 ( .A1(n7899), .A2(n7900), .ZN(n7992) );
  OAI21_X1 U9721 ( .B1(n7900), .B2(n7899), .A(n7992), .ZN(n7901) );
  NAND2_X1 U9722 ( .A1(n7901), .A2(n8385), .ZN(n7905) );
  NAND2_X1 U9723 ( .A1(n8371), .A2(n8612), .ZN(n7902) );
  NAND2_X1 U9724 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8648) );
  OAI211_X1 U9725 ( .C1(n8056), .C2(n8373), .A(n7902), .B(n8648), .ZN(n7903)
         );
  AOI21_X1 U9726 ( .B1(n7919), .B2(n8388), .A(n7903), .ZN(n7904) );
  OAI211_X1 U9727 ( .C1(n7917), .C2(n8395), .A(n7905), .B(n7904), .ZN(P2_U3174) );
  XNOR2_X1 U9728 ( .A(n7906), .B(n8425), .ZN(n7922) );
  NAND2_X1 U9729 ( .A1(n10245), .A2(n10213), .ZN(n8986) );
  AOI21_X1 U9730 ( .B1(n7907), .B2(n8425), .A(n10185), .ZN(n7910) );
  OAI22_X1 U9731 ( .A1(n8056), .A2(n8881), .B1(n8363), .B2(n8883), .ZN(n7908)
         );
  AOI21_X1 U9732 ( .B1(n7910), .B2(n7909), .A(n7908), .ZN(n7916) );
  MUX2_X1 U9733 ( .A(n7916), .B(n8647), .S(n6586), .Z(n7912) );
  NAND2_X1 U9734 ( .A1(n7913), .A2(n8983), .ZN(n7911) );
  OAI211_X1 U9735 ( .C1(n7922), .C2(n8986), .A(n7912), .B(n7911), .ZN(P2_U3472) );
  INV_X1 U9736 ( .A(n10213), .ZN(n10225) );
  MUX2_X1 U9737 ( .A(n7916), .B(n10377), .S(n10229), .Z(n7915) );
  NAND2_X1 U9738 ( .A1(n7913), .A2(n9066), .ZN(n7914) );
  OAI211_X1 U9739 ( .C1(n7922), .C2(n9070), .A(n7915), .B(n7914), .ZN(P2_U3429) );
  OAI21_X1 U9740 ( .B1(n7917), .B2(n8928), .A(n7916), .ZN(n7918) );
  NAND2_X1 U9741 ( .A1(n7918), .A2(n10181), .ZN(n7921) );
  AOI22_X1 U9742 ( .A1(n10183), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n10175), 
        .B2(n7919), .ZN(n7920) );
  OAI211_X1 U9743 ( .C1(n7922), .C2(n8934), .A(n7921), .B(n7920), .ZN(P2_U3220) );
  INV_X1 U9744 ( .A(n7923), .ZN(n7931) );
  INV_X1 U9745 ( .A(n9844), .ZN(n7926) );
  AOI22_X1 U9746 ( .A1(n10112), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n9109), .B2(
        n10110), .ZN(n7925) );
  NAND2_X1 U9747 ( .A1(n9929), .A2(n9113), .ZN(n7924) );
  OAI211_X1 U9748 ( .C1(n7927), .C2(n7926), .A(n7925), .B(n7924), .ZN(n7928)
         );
  AOI21_X1 U9749 ( .B1(n7929), .B2(n10119), .A(n7928), .ZN(n7930) );
  OAI21_X1 U9750 ( .B1(n7931), .B2(n10112), .A(n7930), .ZN(P1_U3283) );
  NAND2_X1 U9751 ( .A1(n7934), .A2(n10043), .ZN(n7932) );
  OAI211_X1 U9752 ( .C1(n7933), .C2(n10060), .A(n7932), .B(n9538), .ZN(
        P1_U3332) );
  NAND2_X1 U9753 ( .A1(n7934), .A2(n9081), .ZN(n7936) );
  NAND2_X1 U9754 ( .A1(n7935), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8595) );
  OAI211_X1 U9755 ( .C1(n7937), .C2(n9077), .A(n7936), .B(n8595), .ZN(P2_U3272) );
  AOI22_X1 U9756 ( .A1(n10112), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9142), .B2(
        n10110), .ZN(n7939) );
  NAND2_X1 U9757 ( .A1(n9145), .A2(n9929), .ZN(n7938) );
  OAI211_X1 U9758 ( .C1(n7940), .C2(n9876), .A(n7939), .B(n7938), .ZN(n7941)
         );
  AOI21_X1 U9759 ( .B1(n7942), .B2(n10119), .A(n7941), .ZN(n7943) );
  OAI21_X1 U9760 ( .B1(n7944), .B2(n10112), .A(n7943), .ZN(P1_U3281) );
  XNOR2_X1 U9761 ( .A(n9414), .B(n7945), .ZN(n7946) );
  OAI222_X1 U9762 ( .A1(n9896), .A2(n7948), .B1(n9898), .B2(n7947), .C1(n7946), 
        .C2(n9893), .ZN(n10133) );
  INV_X1 U9763 ( .A(n10133), .ZN(n7958) );
  OAI21_X1 U9764 ( .B1(n7950), .B2(n9414), .A(n7949), .ZN(n10135) );
  OAI211_X1 U9765 ( .C1(n7951), .C2(n10132), .A(n7445), .B(n9976), .ZN(n10130)
         );
  OAI22_X1 U9766 ( .A1(n9776), .A2(n7952), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9922), .ZN(n7953) );
  AOI21_X1 U9767 ( .B1(n9929), .B2(n7954), .A(n7953), .ZN(n7955) );
  OAI21_X1 U9768 ( .B1(n9876), .B2(n10130), .A(n7955), .ZN(n7956) );
  AOI21_X1 U9769 ( .B1(n10119), .B2(n10135), .A(n7956), .ZN(n7957) );
  OAI21_X1 U9770 ( .B1(n7958), .B2(n10112), .A(n7957), .ZN(P1_U3290) );
  INV_X1 U9771 ( .A(n7959), .ZN(n7961) );
  AOI21_X1 U9772 ( .B1(n7961), .B2(n10213), .A(n7960), .ZN(n7963) );
  MUX2_X1 U9773 ( .A(n10328), .B(n7963), .S(n10245), .Z(n7962) );
  OAI21_X1 U9774 ( .B1(n7966), .B2(n8974), .A(n7962), .ZN(P2_U3471) );
  MUX2_X1 U9775 ( .A(n7964), .B(n7963), .S(n10230), .Z(n7965) );
  OAI21_X1 U9776 ( .B1(n7966), .B2(n9045), .A(n7965), .ZN(P2_U3426) );
  INV_X1 U9777 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10440) );
  INV_X1 U9778 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7972) );
  NAND2_X1 U9779 ( .A1(n7967), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7971) );
  INV_X1 U9780 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7968) );
  OR2_X1 U9781 ( .A1(n7969), .A2(n7968), .ZN(n7970) );
  OAI211_X1 U9782 ( .C1(n7973), .C2(n7972), .A(n7971), .B(n7970), .ZN(n7974)
         );
  INV_X1 U9783 ( .A(n7974), .ZN(n7975) );
  NAND2_X1 U9784 ( .A1(n8593), .A2(P2_U3893), .ZN(n7977) );
  OAI21_X1 U9785 ( .B1(P2_U3893), .B2(n10440), .A(n7977), .ZN(P2_U3522) );
  XNOR2_X1 U9786 ( .A(n7978), .B(n9195), .ZN(n7979) );
  NOR2_X1 U9787 ( .A1(n7979), .A2(n7980), .ZN(n9194) );
  AOI21_X1 U9788 ( .B1(n7980), .B2(n7979), .A(n9194), .ZN(n7988) );
  AOI22_X1 U9789 ( .A1(n9284), .A2(n9554), .B1(n9267), .B2(n7981), .ZN(n7983)
         );
  OAI211_X1 U9790 ( .C1(n7984), .C2(n9279), .A(n7983), .B(n7982), .ZN(n7985)
         );
  AOI21_X1 U9791 ( .B1(n7986), .B2(n9223), .A(n7985), .ZN(n7987) );
  OAI21_X1 U9792 ( .B1(n7988), .B2(n9262), .A(n7987), .ZN(P1_U3221) );
  INV_X1 U9793 ( .A(n9067), .ZN(n8929) );
  INV_X1 U9794 ( .A(n7989), .ZN(n7990) );
  XNOR2_X1 U9795 ( .A(n9067), .B(n8101), .ZN(n8057) );
  XNOR2_X1 U9796 ( .A(n8057), .B(n8056), .ZN(n7991) );
  AOI21_X1 U9797 ( .B1(n7992), .B2(n7990), .A(n7991), .ZN(n8059) );
  AND3_X1 U9798 ( .A1(n7992), .A2(n7991), .A3(n7990), .ZN(n7993) );
  OAI21_X1 U9799 ( .B1(n8059), .B2(n7993), .A(n8385), .ZN(n7997) );
  NAND2_X1 U9800 ( .A1(n8371), .A2(n8925), .ZN(n7994) );
  NAND2_X1 U9801 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8668) );
  OAI211_X1 U9802 ( .C1(n8081), .C2(n8373), .A(n7994), .B(n8668), .ZN(n7995)
         );
  AOI21_X1 U9803 ( .B1(n8931), .B2(n8388), .A(n7995), .ZN(n7996) );
  OAI211_X1 U9804 ( .C1(n8929), .C2(n8395), .A(n7997), .B(n7996), .ZN(P2_U3155) );
  INV_X1 U9805 ( .A(n7998), .ZN(n8055) );
  OAI222_X1 U9806 ( .A1(n7999), .A2(P1_U3086), .B1(n10058), .B2(n8055), .C1(
        n10550), .C2(n10060), .ZN(P1_U3331) );
  INV_X1 U9807 ( .A(n8000), .ZN(n8001) );
  NOR2_X1 U9808 ( .A1(n4439), .A2(n8001), .ZN(n8289) );
  XNOR2_X1 U9809 ( .A(n8289), .B(n8288), .ZN(n8002) );
  NOR2_X1 U9810 ( .A1(n8002), .A2(n8003), .ZN(n8287) );
  AOI21_X1 U9811 ( .B1(n8003), .B2(n8002), .A(n8287), .ZN(n8008) );
  NAND2_X1 U9812 ( .A1(n8371), .A2(n8615), .ZN(n8004) );
  NAND2_X1 U9813 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8628) );
  OAI211_X1 U9814 ( .C1(n8296), .C2(n8373), .A(n8004), .B(n8628), .ZN(n8006)
         );
  NOR2_X1 U9815 ( .A1(n8336), .A2(n8165), .ZN(n8005) );
  AOI211_X1 U9816 ( .C1(n8375), .C2(n8167), .A(n8006), .B(n8005), .ZN(n8007)
         );
  OAI21_X1 U9817 ( .B1(n8008), .B2(n8378), .A(n8007), .ZN(P2_U3157) );
  NOR2_X1 U9818 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n8046) );
  NOR2_X1 U9819 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8044) );
  NOR2_X1 U9820 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n8041) );
  NOR2_X1 U9821 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8038) );
  NOR2_X1 U9822 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8036) );
  NOR2_X1 U9823 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8034) );
  NOR2_X1 U9824 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n8032) );
  NOR2_X1 U9825 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n8030) );
  NOR2_X1 U9826 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n8028) );
  NOR2_X1 U9827 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n8025) );
  NOR2_X1 U9828 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n8022) );
  NOR2_X1 U9829 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n8020) );
  NOR2_X1 U9830 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n8018) );
  NOR2_X1 U9831 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n8016) );
  NAND2_X1 U9832 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n8014) );
  AOI22_X1 U9833 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .B1(n10344), .B2(n10414), .ZN(n10596) );
  NAND2_X1 U9834 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n8012) );
  AOI21_X1 U9835 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10247) );
  INV_X1 U9836 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9562) );
  NAND2_X1 U9837 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n8009) );
  NOR2_X1 U9838 ( .A1(n9562), .A2(n8009), .ZN(n10246) );
  NOR2_X1 U9839 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10246), .ZN(n8010) );
  NOR2_X1 U9840 ( .A1(n10247), .A2(n8010), .ZN(n10594) );
  XOR2_X1 U9841 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10593) );
  NAND2_X1 U9842 ( .A1(n10594), .A2(n10593), .ZN(n8011) );
  NAND2_X1 U9843 ( .A1(n8012), .A2(n8011), .ZN(n10595) );
  NAND2_X1 U9844 ( .A1(n10596), .A2(n10595), .ZN(n8013) );
  NAND2_X1 U9845 ( .A1(n8014), .A2(n8013), .ZN(n10598) );
  XNOR2_X1 U9846 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10597) );
  NOR2_X1 U9847 ( .A1(n10598), .A2(n10597), .ZN(n8015) );
  NOR2_X1 U9848 ( .A1(n8016), .A2(n8015), .ZN(n10584) );
  XNOR2_X1 U9849 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10583) );
  NOR2_X1 U9850 ( .A1(n10584), .A2(n10583), .ZN(n8017) );
  NOR2_X1 U9851 ( .A1(n8018), .A2(n8017), .ZN(n10592) );
  XNOR2_X1 U9852 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10591) );
  NOR2_X1 U9853 ( .A1(n10592), .A2(n10591), .ZN(n8019) );
  XNOR2_X1 U9854 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10587) );
  INV_X1 U9855 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n8023) );
  INV_X1 U9856 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10342) );
  AOI22_X1 U9857 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n8023), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n10342), .ZN(n10589) );
  INV_X1 U9858 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10079) );
  AOI22_X1 U9859 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10079), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n8026), .ZN(n10585) );
  INV_X1 U9860 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U9861 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n7196), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n10357), .ZN(n10266) );
  XNOR2_X1 U9862 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10264) );
  XNOR2_X1 U9863 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10262) );
  XNOR2_X1 U9864 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10260) );
  XNOR2_X1 U9865 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10258) );
  INV_X1 U9866 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n8039) );
  INV_X1 U9867 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8688) );
  AOI22_X1 U9868 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n8039), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n8688), .ZN(n10256) );
  NOR2_X1 U9869 ( .A1(n10257), .A2(n10256), .ZN(n8040) );
  NOR2_X1 U9870 ( .A1(n8041), .A2(n8040), .ZN(n10255) );
  INV_X1 U9871 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n8042) );
  INV_X1 U9872 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8715) );
  AOI22_X1 U9873 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n8042), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n8715), .ZN(n10254) );
  NOR2_X1 U9874 ( .A1(n10255), .A2(n10254), .ZN(n8043) );
  NOR2_X1 U9875 ( .A1(n8044), .A2(n8043), .ZN(n10253) );
  XNOR2_X1 U9876 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10252) );
  NOR2_X1 U9877 ( .A1(n10253), .A2(n10252), .ZN(n8045) );
  NOR2_X1 U9878 ( .A1(n8046), .A2(n8045), .ZN(n8047) );
  AND2_X1 U9879 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n8047), .ZN(n10250) );
  NOR2_X1 U9880 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10250), .ZN(n8048) );
  NOR2_X1 U9881 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n8047), .ZN(n10249) );
  NOR2_X1 U9882 ( .A1(n8048), .A2(n10249), .ZN(n8050) );
  XNOR2_X1 U9883 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8049) );
  XNOR2_X1 U9884 ( .A(n8050), .B(n8049), .ZN(ADD_1068_U4) );
  INV_X1 U9885 ( .A(n8051), .ZN(n8122) );
  OAI222_X1 U9886 ( .A1(n8053), .A2(P1_U3086), .B1(n10058), .B2(n8122), .C1(
        n8052), .C2(n10060), .ZN(P1_U3330) );
  OAI222_X1 U9887 ( .A1(P2_U3151), .A2(n6559), .B1(n9090), .B2(n8055), .C1(
        n8054), .C2(n9077), .ZN(P2_U3271) );
  INV_X1 U9888 ( .A(n9061), .ZN(n8066) );
  XNOR2_X1 U9889 ( .A(n9061), .B(n8101), .ZN(n8080) );
  XNOR2_X1 U9890 ( .A(n8080), .B(n8926), .ZN(n8060) );
  NAND2_X1 U9891 ( .A1(n8061), .A2(n8060), .ZN(n8079) );
  OAI211_X1 U9892 ( .C1(n8061), .C2(n8060), .A(n8079), .B(n8385), .ZN(n8065)
         );
  NAND2_X1 U9893 ( .A1(n8371), .A2(n8915), .ZN(n8062) );
  NAND2_X1 U9894 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n10277) );
  OAI211_X1 U9895 ( .C1(n8313), .C2(n8373), .A(n8062), .B(n10277), .ZN(n8063)
         );
  AOI21_X1 U9896 ( .B1(n8919), .B2(n8388), .A(n8063), .ZN(n8064) );
  OAI211_X1 U9897 ( .C1(n8066), .C2(n8395), .A(n8065), .B(n8064), .ZN(P2_U3181) );
  INV_X1 U9898 ( .A(n8067), .ZN(n8070) );
  OAI222_X1 U9899 ( .A1(P2_U3151), .A2(n8068), .B1(n9090), .B2(n8070), .C1(
        n10474), .C2(n9077), .ZN(P2_U3269) );
  OAI222_X1 U9900 ( .A1(n8071), .A2(P1_U3086), .B1(n10058), .B2(n8070), .C1(
        n8069), .C2(n10060), .ZN(P1_U3329) );
  NOR2_X1 U9901 ( .A1(n8074), .A2(n8885), .ZN(n8773) );
  AOI21_X1 U9902 ( .B1(n10183), .B2(P2_REG2_REG_29__SCAN_IN), .A(n8773), .ZN(
        n8075) );
  OAI21_X1 U9903 ( .B1(n8076), .B2(n8873), .A(n8075), .ZN(n8077) );
  AOI21_X1 U9904 ( .B1(n8073), .B2(n10177), .A(n8077), .ZN(n8078) );
  OAI21_X1 U9905 ( .B1(n8072), .B2(n10183), .A(n8078), .ZN(P2_U3204) );
  XOR2_X1 U9906 ( .A(n8101), .B(n9055), .Z(n8314) );
  NOR2_X1 U9907 ( .A1(n5203), .A2(n8313), .ZN(n8082) );
  XNOR2_X1 U9908 ( .A(n9049), .B(n8101), .ZN(n8083) );
  XNOR2_X1 U9909 ( .A(n8083), .B(n8907), .ZN(n8322) );
  XNOR2_X1 U9910 ( .A(n8969), .B(n8101), .ZN(n8084) );
  XNOR2_X1 U9911 ( .A(n8084), .B(n8870), .ZN(n8369) );
  INV_X1 U9912 ( .A(n8084), .ZN(n8085) );
  XNOR2_X1 U9913 ( .A(n8967), .B(n8101), .ZN(n8086) );
  XNOR2_X1 U9914 ( .A(n8086), .B(n8611), .ZN(n8272) );
  XNOR2_X1 U9915 ( .A(n9034), .B(n8101), .ZN(n8087) );
  XNOR2_X1 U9916 ( .A(n8087), .B(n8867), .ZN(n8340) );
  XNOR2_X1 U9917 ( .A(n9028), .B(n8101), .ZN(n8088) );
  XNOR2_X1 U9918 ( .A(n8088), .B(n8610), .ZN(n8280) );
  XNOR2_X1 U9919 ( .A(n9023), .B(n8101), .ZN(n8089) );
  NOR2_X1 U9920 ( .A1(n8089), .A2(n8543), .ZN(n8350) );
  NAND2_X1 U9921 ( .A1(n8089), .A2(n8543), .ZN(n8348) );
  XNOR2_X1 U9922 ( .A(n8261), .B(n8090), .ZN(n8263) );
  XNOR2_X1 U9923 ( .A(n8329), .B(n8101), .ZN(n8091) );
  NAND2_X1 U9924 ( .A1(n8091), .A2(n4449), .ZN(n8302) );
  OAI21_X1 U9925 ( .B1(n8091), .B2(n4449), .A(n8302), .ZN(n8330) );
  AOI21_X1 U9926 ( .B1(n8263), .B2(n8609), .A(n8330), .ZN(n8092) );
  NAND2_X1 U9927 ( .A1(n8301), .A2(n8302), .ZN(n8096) );
  XNOR2_X1 U9928 ( .A(n9007), .B(n8101), .ZN(n8093) );
  NAND2_X1 U9929 ( .A1(n8093), .A2(n8815), .ZN(n8380) );
  INV_X1 U9930 ( .A(n8093), .ZN(n8094) );
  NAND2_X1 U9931 ( .A1(n8094), .A2(n8608), .ZN(n8095) );
  AND2_X1 U9932 ( .A1(n8380), .A2(n8095), .ZN(n8303) );
  NAND2_X1 U9933 ( .A1(n8096), .A2(n8303), .ZN(n8305) );
  NAND2_X1 U9934 ( .A1(n8305), .A2(n8380), .ZN(n8097) );
  XNOR2_X1 U9935 ( .A(n9001), .B(n8101), .ZN(n8098) );
  XNOR2_X1 U9936 ( .A(n8098), .B(n8802), .ZN(n8381) );
  XNOR2_X1 U9937 ( .A(n8571), .B(n8101), .ZN(n8100) );
  XNOR2_X1 U9938 ( .A(n8100), .B(n8793), .ZN(n8251) );
  XNOR2_X1 U9939 ( .A(n8779), .B(n8101), .ZN(n8102) );
  XNOR2_X1 U9940 ( .A(n8103), .B(n8102), .ZN(n8108) );
  AOI22_X1 U9941 ( .A1(n8784), .A2(n8388), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8105) );
  NAND2_X1 U9942 ( .A1(n8781), .A2(n8371), .ZN(n8104) );
  OAI211_X1 U9943 ( .C1(n8606), .C2(n8373), .A(n8105), .B(n8104), .ZN(n8106)
         );
  AOI21_X1 U9944 ( .B1(n8582), .B2(n8375), .A(n8106), .ZN(n8107) );
  OAI21_X1 U9945 ( .B1(n8108), .B2(n8378), .A(n8107), .ZN(P2_U3160) );
  INV_X1 U9946 ( .A(n8109), .ZN(n10055) );
  OAI222_X1 U9947 ( .A1(n9077), .A2(n8111), .B1(n9090), .B2(n10055), .C1(n8110), .C2(P2_U3151), .ZN(P2_U3266) );
  OAI22_X1 U9948 ( .A1(n9736), .A2(n9279), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8114), .ZN(n8115) );
  AOI21_X1 U9949 ( .B1(n9708), .B2(n9267), .A(n8115), .ZN(n8116) );
  OAI21_X1 U9950 ( .B1(n9703), .B2(n9250), .A(n8116), .ZN(n8117) );
  AOI21_X1 U9951 ( .B1(n8118), .B2(n9236), .A(n8117), .ZN(n8119) );
  OAI21_X1 U9952 ( .B1(n8120), .B2(n9262), .A(n8119), .ZN(P1_U3214) );
  OAI222_X1 U9953 ( .A1(P2_U3151), .A2(n6560), .B1(n9090), .B2(n8122), .C1(
        n8121), .C2(n9077), .ZN(P2_U3270) );
  INV_X1 U9954 ( .A(n8124), .ZN(n8127) );
  NAND3_X1 U9955 ( .A1(n8127), .A2(n8126), .A3(n8125), .ZN(n8128) );
  AOI21_X1 U9956 ( .B1(n8123), .B2(n8128), .A(n9262), .ZN(n8134) );
  OAI22_X1 U9957 ( .A1(n9448), .A2(n9279), .B1(n9250), .B2(n8129), .ZN(n8133)
         );
  OAI22_X1 U9958 ( .A1(n9287), .A2(n8131), .B1(n8130), .B2(n9581), .ZN(n8132)
         );
  OR3_X1 U9959 ( .A1(n8134), .A2(n8133), .A3(n8132), .ZN(P1_U3237) );
  INV_X1 U9960 ( .A(SI_29_), .ZN(n10419) );
  OAI21_X2 U9961 ( .B1(n8138), .B2(n10419), .A(n8137), .ZN(n8150) );
  INV_X1 U9962 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8399) );
  INV_X1 U9963 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10054) );
  MUX2_X1 U9964 ( .A(n8399), .B(n10054), .S(n8144), .Z(n8140) );
  INV_X1 U9965 ( .A(SI_30_), .ZN(n8139) );
  NAND2_X1 U9966 ( .A1(n8140), .A2(n8139), .ZN(n8143) );
  INV_X1 U9967 ( .A(n8140), .ZN(n8141) );
  NAND2_X1 U9968 ( .A1(n8141), .A2(SI_30_), .ZN(n8142) );
  NAND2_X1 U9969 ( .A1(n8143), .A2(n8142), .ZN(n8149) );
  OAI21_X2 U9970 ( .B1(n8150), .B2(n8149), .A(n8143), .ZN(n8147) );
  INV_X1 U9971 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9078) );
  MUX2_X1 U9972 ( .A(n9078), .B(n10440), .S(n8144), .Z(n8145) );
  XNOR2_X1 U9973 ( .A(n8145), .B(SI_31_), .ZN(n8146) );
  XNOR2_X2 U9974 ( .A(n8147), .B(n8146), .ZN(n10044) );
  NOR2_X1 U9975 ( .A1(n8151), .A2(n10440), .ZN(n8148) );
  INV_X1 U9976 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8160) );
  NAND2_X1 U9977 ( .A1(n8398), .A2(n5505), .ZN(n8153) );
  OR2_X1 U9978 ( .A1(n8151), .A2(n10054), .ZN(n8152) );
  INV_X1 U9979 ( .A(n8156), .ZN(n8159) );
  INV_X1 U9980 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n10271) );
  NAND2_X1 U9981 ( .A1(n5894), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8158) );
  NAND2_X1 U9982 ( .A1(n6153), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8157) );
  OAI211_X1 U9983 ( .C1(n5837), .C2(n10271), .A(n8158), .B(n8157), .ZN(n9543)
         );
  NOR2_X1 U9984 ( .A1(n9675), .A2(n9932), .ZN(n8216) );
  OAI21_X1 U9985 ( .B1(n9679), .B2(n10026), .A(n8161), .ZN(P1_U3521) );
  INV_X1 U9986 ( .A(n8162), .ZN(n8163) );
  MUX2_X1 U9987 ( .A(n8164), .B(n8163), .S(n10181), .Z(n8169) );
  INV_X1 U9988 ( .A(n8165), .ZN(n8166) );
  AOI22_X1 U9989 ( .A1(n10178), .A2(n8167), .B1(n10175), .B2(n8166), .ZN(n8168) );
  OAI211_X1 U9990 ( .C1(n8171), .C2(n8170), .A(n8169), .B(n8168), .ZN(P2_U3223) );
  XOR2_X1 U9991 ( .A(n8172), .B(n8552), .Z(n9017) );
  INV_X1 U9992 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8176) );
  XNOR2_X1 U9993 ( .A(n8173), .B(n8552), .ZN(n8174) );
  OAI222_X1 U9994 ( .A1(n8881), .A2(n4449), .B1(n8883), .B2(n8543), .C1(n10185), .C2(n8174), .ZN(n9018) );
  INV_X1 U9995 ( .A(n9018), .ZN(n8175) );
  MUX2_X1 U9996 ( .A(n8176), .B(n8175), .S(n10181), .Z(n8178) );
  AOI22_X1 U9997 ( .A1(n8261), .A2(n10178), .B1(n10175), .B2(n8269), .ZN(n8177) );
  OAI211_X1 U9998 ( .C1(n9017), .C2(n8934), .A(n8178), .B(n8177), .ZN(P2_U3210) );
  XNOR2_X1 U9999 ( .A(n8179), .B(n8567), .ZN(n8943) );
  XNOR2_X1 U10000 ( .A(n8180), .B(n8567), .ZN(n8181) );
  OAI222_X1 U10001 ( .A1(n8881), .A2(n8182), .B1(n8883), .B2(n8257), .C1(
        n10185), .C2(n8181), .ZN(n8941) );
  INV_X1 U10002 ( .A(n8941), .ZN(n8186) );
  MUX2_X1 U10003 ( .A(n8183), .B(n8186), .S(n10230), .Z(n8185) );
  NAND2_X1 U10004 ( .A1(n8571), .A2(n9066), .ZN(n8184) );
  OAI211_X1 U10005 ( .C1(n8943), .C2(n9070), .A(n8185), .B(n8184), .ZN(
        P2_U3454) );
  INV_X1 U10006 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8187) );
  MUX2_X1 U10007 ( .A(n8187), .B(n8186), .S(n10181), .Z(n8189) );
  AOI22_X1 U10008 ( .A1(n8571), .A2(n10178), .B1(n10175), .B2(n8255), .ZN(
        n8188) );
  OAI211_X1 U10009 ( .C1(n8943), .C2(n8934), .A(n8189), .B(n8188), .ZN(
        P2_U3206) );
  INV_X1 U10010 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8194) );
  NAND2_X1 U10011 ( .A1(n8205), .A2(n8195), .ZN(n8196) );
  NAND2_X1 U10012 ( .A1(n8196), .A2(n9623), .ZN(n9633) );
  INV_X1 U10013 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U10014 ( .A1(n8198), .A2(n8197), .ZN(n8199) );
  OAI21_X1 U10015 ( .B1(n8198), .B2(n8197), .A(n8199), .ZN(n9632) );
  INV_X1 U10016 ( .A(n8199), .ZN(n8200) );
  XNOR2_X1 U10017 ( .A(n9651), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9645) );
  NOR2_X1 U10018 ( .A1(n9651), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9660) );
  XNOR2_X1 U10019 ( .A(n8209), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9659) );
  AOI21_X1 U10020 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n8209), .A(n9658), .ZN(
        n8201) );
  NOR2_X1 U10021 ( .A1(n8204), .A2(n9628), .ZN(n8206) );
  INV_X1 U10022 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10368) );
  NOR2_X1 U10023 ( .A1(n8206), .A2(n9621), .ZN(n9638) );
  XNOR2_X1 U10024 ( .A(n9641), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9637) );
  NAND2_X1 U10025 ( .A1(n9641), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8207) );
  XNOR2_X1 U10026 ( .A(n9651), .B(n8208), .ZN(n9653) );
  MUX2_X1 U10027 ( .A(n9859), .B(P1_REG2_REG_18__SCAN_IN), .S(n8209), .Z(n9667) );
  NOR2_X1 U10028 ( .A1(n9668), .A2(n9667), .ZN(n9666) );
  AND2_X1 U10029 ( .A1(n8209), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8210) );
  XNOR2_X1 U10030 ( .A(n8211), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n8214) );
  OAI21_X1 U10031 ( .B1(n8212), .B2(n10090), .A(n10088), .ZN(n8213) );
  NAND2_X1 U10032 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9123) );
  INV_X1 U10033 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8217) );
  OAI21_X1 U10034 ( .B1(n9679), .B2(n9948), .A(n8218), .ZN(P1_U3553) );
  XOR2_X1 U10035 ( .A(n9428), .B(n8219), .Z(n9990) );
  OAI211_X1 U10036 ( .C1(n8221), .C2(n9428), .A(n8220), .B(n9918), .ZN(n8223)
         );
  AOI22_X1 U10037 ( .A1(n9835), .A2(n9913), .B1(n9915), .B2(n9550), .ZN(n8222)
         );
  NAND2_X1 U10038 ( .A1(n8223), .A2(n8222), .ZN(n9986) );
  INV_X1 U10039 ( .A(n8224), .ZN(n9871) );
  AOI211_X1 U10040 ( .C1(n9988), .C2(n9871), .A(n9907), .B(n9849), .ZN(n9987)
         );
  NAND2_X1 U10041 ( .A1(n9987), .A2(n10108), .ZN(n8227) );
  AOI22_X1 U10042 ( .A1(n10112), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n8225), 
        .B2(n10110), .ZN(n8226) );
  OAI211_X1 U10043 ( .C1(n6100), .C2(n10115), .A(n8227), .B(n8226), .ZN(n8228)
         );
  AOI21_X1 U10044 ( .B1(n9776), .B2(n9986), .A(n8228), .ZN(n8229) );
  OAI21_X1 U10045 ( .B1(n9990), .B2(n9926), .A(n8229), .ZN(P1_U3276) );
  XNOR2_X1 U10046 ( .A(n9879), .B(n9426), .ZN(n10001) );
  INV_X1 U10047 ( .A(n9890), .ZN(n8231) );
  INV_X1 U10048 ( .A(n9870), .ZN(n8230) );
  AOI211_X1 U10049 ( .C1(n9998), .C2(n8231), .A(n9907), .B(n8230), .ZN(n9997)
         );
  AOI22_X1 U10050 ( .A1(n10112), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9278), 
        .B2(n10110), .ZN(n8232) );
  OAI21_X1 U10051 ( .B1(n9288), .B2(n10115), .A(n8232), .ZN(n8238) );
  OAI21_X1 U10052 ( .B1(n4453), .B2(n8233), .A(n9426), .ZN(n8235) );
  NAND2_X1 U10053 ( .A1(n8235), .A2(n8234), .ZN(n8236) );
  AOI222_X1 U10054 ( .A1(n9918), .A2(n8236), .B1(n9550), .B2(n9913), .C1(n9914), .C2(n9915), .ZN(n10000) );
  NOR2_X1 U10055 ( .A1(n10000), .A2(n10112), .ZN(n8237) );
  AOI211_X1 U10056 ( .C1(n9997), .C2(n10108), .A(n8238), .B(n8237), .ZN(n8239)
         );
  OAI21_X1 U10057 ( .B1(n9926), .B2(n10001), .A(n8239), .ZN(P1_U3278) );
  INV_X1 U10058 ( .A(n8398), .ZN(n10053) );
  OAI222_X1 U10059 ( .A1(P2_U3151), .A2(n8240), .B1(n9090), .B2(n10053), .C1(
        n8399), .C2(n9077), .ZN(P2_U3265) );
  NAND2_X1 U10060 ( .A1(n8241), .A2(n10108), .ZN(n8244) );
  AOI22_X1 U10061 ( .A1(n8242), .A2(n10110), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10112), .ZN(n8243) );
  OAI211_X1 U10062 ( .C1(n8245), .C2(n10115), .A(n8244), .B(n8243), .ZN(n8246)
         );
  AOI21_X1 U10063 ( .B1(n8247), .B2(n9776), .A(n8246), .ZN(n8248) );
  OAI21_X1 U10064 ( .B1(n8249), .B2(n9926), .A(n8248), .ZN(P1_U3265) );
  INV_X1 U10065 ( .A(n6480), .ZN(n9085) );
  OAI222_X1 U10066 ( .A1(n10060), .A2(n8250), .B1(P1_U3086), .B2(n4437), .C1(
        n10058), .C2(n9085), .ZN(P1_U3327) );
  INV_X1 U10067 ( .A(n8571), .ZN(n8942) );
  AOI21_X1 U10068 ( .B1(n8252), .B2(n8251), .A(n8378), .ZN(n8254) );
  NAND2_X1 U10069 ( .A1(n8254), .A2(n8253), .ZN(n8260) );
  AOI22_X1 U10070 ( .A1(n8255), .A2(n8388), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8256) );
  OAI21_X1 U10071 ( .B1(n8257), .B2(n8390), .A(n8256), .ZN(n8258) );
  AOI21_X1 U10072 ( .B1(n8392), .B2(n8607), .A(n8258), .ZN(n8259) );
  OAI211_X1 U10073 ( .C1(n8942), .C2(n8395), .A(n8260), .B(n8259), .ZN(
        P2_U3154) );
  INV_X1 U10074 ( .A(n8261), .ZN(n9016) );
  INV_X1 U10075 ( .A(n8262), .ZN(n8264) );
  NAND2_X1 U10076 ( .A1(n8265), .A2(n8826), .ZN(n8331) );
  OAI21_X1 U10077 ( .B1(n8826), .B2(n8265), .A(n8331), .ZN(n8266) );
  NAND2_X1 U10078 ( .A1(n8266), .A2(n8385), .ZN(n8271) );
  AOI22_X1 U10079 ( .A1(n8839), .A2(n8371), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8267) );
  OAI21_X1 U10080 ( .B1(n4449), .B2(n8373), .A(n8267), .ZN(n8268) );
  AOI21_X1 U10081 ( .B1(n8269), .B2(n8388), .A(n8268), .ZN(n8270) );
  OAI211_X1 U10082 ( .C1(n9016), .C2(n8395), .A(n8271), .B(n8270), .ZN(
        P2_U3156) );
  XOR2_X1 U10083 ( .A(n8273), .B(n8272), .Z(n8279) );
  NAND2_X1 U10084 ( .A1(n8371), .A2(n8899), .ZN(n8275) );
  OAI211_X1 U10085 ( .C1(n8867), .C2(n8373), .A(n8275), .B(n8274), .ZN(n8277)
         );
  NOR2_X1 U10086 ( .A1(n8874), .A2(n8395), .ZN(n8276) );
  AOI211_X1 U10087 ( .C1(n8871), .C2(n8388), .A(n8277), .B(n8276), .ZN(n8278)
         );
  OAI21_X1 U10088 ( .B1(n8279), .B2(n8378), .A(n8278), .ZN(P2_U3159) );
  XOR2_X1 U10089 ( .A(n8281), .B(n8280), .Z(n8286) );
  AOI22_X1 U10090 ( .A1(n8839), .A2(n8392), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8283) );
  NAND2_X1 U10091 ( .A1(n8388), .A2(n8842), .ZN(n8282) );
  OAI211_X1 U10092 ( .C1(n8867), .C2(n8390), .A(n8283), .B(n8282), .ZN(n8284)
         );
  AOI21_X1 U10093 ( .B1(n9028), .B2(n8375), .A(n8284), .ZN(n8285) );
  OAI21_X1 U10094 ( .B1(n8286), .B2(n8378), .A(n8285), .ZN(P2_U3163) );
  AOI21_X1 U10095 ( .B1(n8289), .B2(n8288), .A(n8287), .ZN(n8360) );
  NAND2_X1 U10096 ( .A1(n8360), .A2(n8359), .ZN(n8358) );
  OAI21_X1 U10097 ( .B1(n8296), .B2(n8359), .A(n8358), .ZN(n8290) );
  XOR2_X1 U10098 ( .A(n8291), .B(n8290), .Z(n8300) );
  NAND2_X1 U10099 ( .A1(n8388), .A2(n8292), .ZN(n8295) );
  AOI21_X1 U10100 ( .B1(n8392), .B2(n8925), .A(n8293), .ZN(n8294) );
  OAI211_X1 U10101 ( .C1(n8390), .C2(n8296), .A(n8295), .B(n8294), .ZN(n8297)
         );
  AOI21_X1 U10102 ( .B1(n8298), .B2(n8375), .A(n8297), .ZN(n8299) );
  OAI21_X1 U10103 ( .B1(n8300), .B2(n8378), .A(n8299), .ZN(P2_U3164) );
  INV_X1 U10104 ( .A(n9007), .ZN(n8312) );
  INV_X1 U10105 ( .A(n8301), .ZN(n8332) );
  INV_X1 U10106 ( .A(n8302), .ZN(n8304) );
  NOR3_X1 U10107 ( .A1(n8332), .A2(n8304), .A3(n8303), .ZN(n8306) );
  INV_X1 U10108 ( .A(n8305), .ZN(n8383) );
  OAI21_X1 U10109 ( .B1(n8306), .B2(n8383), .A(n8385), .ZN(n8311) );
  INV_X1 U10110 ( .A(n8804), .ZN(n8308) );
  AOI22_X1 U10111 ( .A1(n8801), .A2(n8371), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8307) );
  OAI21_X1 U10112 ( .B1(n8308), .B2(n8336), .A(n8307), .ZN(n8309) );
  AOI21_X1 U10113 ( .B1(n8392), .B2(n8802), .A(n8309), .ZN(n8310) );
  OAI211_X1 U10114 ( .C1(n8312), .C2(n8395), .A(n8311), .B(n8310), .ZN(
        P2_U3165) );
  XNOR2_X1 U10115 ( .A(n8314), .B(n8313), .ZN(n8315) );
  XNOR2_X1 U10116 ( .A(n8316), .B(n8315), .ZN(n8321) );
  NAND2_X1 U10117 ( .A1(n8371), .A2(n8926), .ZN(n8317) );
  NAND2_X1 U10118 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8714) );
  OAI211_X1 U10119 ( .C1(n8882), .C2(n8373), .A(n8317), .B(n8714), .ZN(n8318)
         );
  AOI21_X1 U10120 ( .B1(n8910), .B2(n8388), .A(n8318), .ZN(n8320) );
  NAND2_X1 U10121 ( .A1(n9055), .A2(n8375), .ZN(n8319) );
  OAI211_X1 U10122 ( .C1(n8321), .C2(n8378), .A(n8320), .B(n8319), .ZN(
        P2_U3166) );
  XOR2_X1 U10123 ( .A(n8323), .B(n8322), .Z(n8328) );
  NAND2_X1 U10124 ( .A1(n8371), .A2(n8916), .ZN(n8324) );
  NAND2_X1 U10125 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8730) );
  OAI211_X1 U10126 ( .C1(n8870), .C2(n8373), .A(n8324), .B(n8730), .ZN(n8325)
         );
  AOI21_X1 U10127 ( .B1(n8901), .B2(n8388), .A(n8325), .ZN(n8327) );
  NAND2_X1 U10128 ( .A1(n9049), .A2(n8375), .ZN(n8326) );
  OAI211_X1 U10129 ( .C1(n8328), .C2(n8378), .A(n8327), .B(n8326), .ZN(
        P2_U3168) );
  INV_X1 U10130 ( .A(n8329), .ZN(n9011) );
  AND3_X1 U10131 ( .A1(n8331), .A2(n8330), .A3(n4578), .ZN(n8333) );
  OAI21_X1 U10132 ( .B1(n8333), .B2(n8332), .A(n8385), .ZN(n8339) );
  INV_X1 U10133 ( .A(n8334), .ZN(n8816) );
  AOI22_X1 U10134 ( .A1(n8609), .A2(n8371), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8335) );
  OAI21_X1 U10135 ( .B1(n8816), .B2(n8336), .A(n8335), .ZN(n8337) );
  AOI21_X1 U10136 ( .B1(n8392), .B2(n8608), .A(n8337), .ZN(n8338) );
  OAI211_X1 U10137 ( .C1(n9011), .C2(n8395), .A(n8339), .B(n8338), .ZN(
        P2_U3169) );
  XOR2_X1 U10138 ( .A(n8341), .B(n8340), .Z(n8346) );
  AOI22_X1 U10139 ( .A1(n8610), .A2(n8392), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8343) );
  NAND2_X1 U10140 ( .A1(n8388), .A2(n8856), .ZN(n8342) );
  OAI211_X1 U10141 ( .C1(n8880), .C2(n8390), .A(n8343), .B(n8342), .ZN(n8344)
         );
  AOI21_X1 U10142 ( .B1(n9034), .B2(n8375), .A(n8344), .ZN(n8345) );
  OAI21_X1 U10143 ( .B1(n8346), .B2(n8378), .A(n8345), .ZN(P2_U3173) );
  INV_X1 U10144 ( .A(n8348), .ZN(n8349) );
  NOR2_X1 U10145 ( .A1(n8350), .A2(n8349), .ZN(n8351) );
  XNOR2_X1 U10146 ( .A(n8347), .B(n8351), .ZN(n8357) );
  INV_X1 U10147 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8352) );
  OAI22_X1 U10148 ( .A1(n8854), .A2(n8390), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8352), .ZN(n8354) );
  NOR2_X1 U10149 ( .A1(n8826), .A2(n8373), .ZN(n8353) );
  AOI211_X1 U10150 ( .C1(n8829), .C2(n8388), .A(n8354), .B(n8353), .ZN(n8356)
         );
  NAND2_X1 U10151 ( .A1(n9023), .A2(n8375), .ZN(n8355) );
  OAI211_X1 U10152 ( .C1(n8357), .C2(n8378), .A(n8356), .B(n8355), .ZN(
        P2_U3175) );
  INV_X1 U10153 ( .A(n8988), .ZN(n8368) );
  OAI211_X1 U10154 ( .C1(n8360), .C2(n8359), .A(n8358), .B(n8385), .ZN(n8367)
         );
  NAND2_X1 U10155 ( .A1(n8371), .A2(n8614), .ZN(n8362) );
  OAI211_X1 U10156 ( .C1(n8363), .C2(n8373), .A(n8362), .B(n8361), .ZN(n8364)
         );
  AOI21_X1 U10157 ( .B1(n8365), .B2(n8388), .A(n8364), .ZN(n8366) );
  OAI211_X1 U10158 ( .C1(n8368), .C2(n8395), .A(n8367), .B(n8366), .ZN(
        P2_U3176) );
  XOR2_X1 U10159 ( .A(n8370), .B(n8369), .Z(n8379) );
  NAND2_X1 U10160 ( .A1(n8371), .A2(n8907), .ZN(n8372) );
  NAND2_X1 U10161 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8758) );
  OAI211_X1 U10162 ( .C1(n8880), .C2(n8373), .A(n8372), .B(n8758), .ZN(n8374)
         );
  AOI21_X1 U10163 ( .B1(n8884), .B2(n8388), .A(n8374), .ZN(n8377) );
  NAND2_X1 U10164 ( .A1(n8969), .A2(n8375), .ZN(n8376) );
  OAI211_X1 U10165 ( .C1(n8379), .C2(n8378), .A(n8377), .B(n8376), .ZN(
        P2_U3178) );
  INV_X1 U10166 ( .A(n9001), .ZN(n8947) );
  INV_X1 U10167 ( .A(n8380), .ZN(n8382) );
  NOR3_X1 U10168 ( .A1(n8383), .A2(n8382), .A3(n8381), .ZN(n8387) );
  INV_X1 U10169 ( .A(n8384), .ZN(n8386) );
  OAI21_X1 U10170 ( .B1(n8387), .B2(n8386), .A(n8385), .ZN(n8394) );
  AOI22_X1 U10171 ( .A1(n8795), .A2(n8388), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8389) );
  OAI21_X1 U10172 ( .B1(n8815), .B2(n8390), .A(n8389), .ZN(n8391) );
  AOI21_X1 U10173 ( .B1(n8781), .B2(n8392), .A(n8391), .ZN(n8393) );
  OAI211_X1 U10174 ( .C1(n8947), .C2(n8395), .A(n8394), .B(n8393), .ZN(
        P2_U3180) );
  INV_X1 U10175 ( .A(n8581), .ZN(n8396) );
  NOR2_X2 U10176 ( .A1(n8397), .A2(n8396), .ZN(n8442) );
  NAND2_X1 U10177 ( .A1(n8398), .A2(n8402), .ZN(n8401) );
  OR2_X1 U10178 ( .A1(n8403), .A2(n8399), .ZN(n8400) );
  NAND2_X1 U10179 ( .A1(n10044), .A2(n8402), .ZN(n8405) );
  OR2_X1 U10180 ( .A1(n8403), .A2(n9078), .ZN(n8404) );
  INV_X1 U10181 ( .A(n8993), .ZN(n8434) );
  OR2_X1 U10182 ( .A1(n8434), .A2(n8772), .ZN(n8408) );
  INV_X1 U10183 ( .A(n8605), .ZN(n8409) );
  NAND2_X1 U10184 ( .A1(n8994), .A2(n8409), .ZN(n8407) );
  AND2_X1 U10185 ( .A1(n8407), .A2(n8406), .ZN(n8446) );
  NAND2_X1 U10186 ( .A1(n8408), .A2(n8446), .ZN(n8439) );
  INV_X1 U10187 ( .A(n8520), .ZN(n8897) );
  AND4_X1 U10188 ( .A1(n8414), .A2(n8413), .A3(n10184), .A4(n7130), .ZN(n8417)
         );
  INV_X1 U10189 ( .A(n8415), .ZN(n10164) );
  AND4_X1 U10190 ( .A1(n8417), .A2(n8416), .A3(n8461), .A4(n10164), .ZN(n8420)
         );
  NAND4_X1 U10191 ( .A1(n8420), .A2(n8419), .A3(n8465), .A4(n8418), .ZN(n8421)
         );
  NOR3_X1 U10192 ( .A1(n8423), .A2(n8422), .A3(n8421), .ZN(n8424) );
  NAND4_X1 U10193 ( .A1(n8425), .A2(n8484), .A3(n8923), .A4(n8424), .ZN(n8426)
         );
  NOR2_X1 U10194 ( .A1(n8513), .A2(n8426), .ZN(n8427) );
  NAND3_X1 U10195 ( .A1(n8905), .A2(n8897), .A3(n8427), .ZN(n8428) );
  OR3_X1 U10196 ( .A1(n8865), .A2(n8428), .A3(n8889), .ZN(n8429) );
  OR3_X1 U10197 ( .A1(n8834), .A2(n8429), .A3(n8849), .ZN(n8430) );
  NOR2_X1 U10198 ( .A1(n8542), .A2(n8430), .ZN(n8431) );
  NAND4_X1 U10199 ( .A1(n8799), .A2(n8552), .A3(n8812), .A4(n8431), .ZN(n8433)
         );
  INV_X1 U10200 ( .A(n8432), .ZN(n8564) );
  OR2_X1 U10201 ( .A1(n8565), .A2(n8564), .ZN(n8563) );
  NAND4_X1 U10202 ( .A1(n8583), .A2(n4465), .A3(n8779), .A4(n8581), .ZN(n8438)
         );
  INV_X1 U10203 ( .A(n8583), .ZN(n8435) );
  NAND2_X1 U10204 ( .A1(n8435), .A2(n8434), .ZN(n8436) );
  NAND2_X1 U10205 ( .A1(n8442), .A2(n5230), .ZN(n8443) );
  NAND3_X1 U10206 ( .A1(n8445), .A2(n8444), .A3(n8443), .ZN(n8598) );
  INV_X1 U10207 ( .A(n8446), .ZN(n8447) );
  NAND2_X1 U10208 ( .A1(n8447), .A2(n8583), .ZN(n8576) );
  OR2_X1 U10209 ( .A1(n8582), .A2(n8577), .ZN(n8448) );
  NAND2_X1 U10210 ( .A1(n8448), .A2(n8607), .ZN(n8580) );
  INV_X1 U10211 ( .A(n8580), .ZN(n8449) );
  AOI21_X1 U10212 ( .B1(n8449), .B2(n8998), .A(n8570), .ZN(n8575) );
  NAND2_X1 U10213 ( .A1(n8451), .A2(n8450), .ZN(n8453) );
  NAND2_X1 U10214 ( .A1(n8453), .A2(n8452), .ZN(n8503) );
  INV_X1 U10215 ( .A(n7356), .ZN(n8457) );
  AND2_X1 U10216 ( .A1(n8455), .A2(n8454), .ZN(n8458) );
  NAND3_X1 U10217 ( .A1(n8461), .A2(n6530), .A3(n8458), .ZN(n8456) );
  INV_X1 U10218 ( .A(n8458), .ZN(n8459) );
  NAND3_X1 U10219 ( .A1(n8461), .A2(n8460), .A3(n8459), .ZN(n8463) );
  NAND3_X1 U10220 ( .A1(n8463), .A2(n8462), .A3(n8485), .ZN(n8464) );
  NAND2_X1 U10221 ( .A1(n8466), .A2(n8465), .ZN(n8489) );
  INV_X1 U10222 ( .A(n8467), .ZN(n8469) );
  OAI211_X1 U10223 ( .C1(n8489), .C2(n8469), .A(n8490), .B(n8468), .ZN(n8470)
         );
  NAND2_X1 U10224 ( .A1(n8494), .A2(n8471), .ZN(n8473) );
  NAND2_X1 U10225 ( .A1(n8481), .A2(n8477), .ZN(n8472) );
  NAND3_X1 U10226 ( .A1(n8475), .A2(n8493), .A3(n8491), .ZN(n8482) );
  INV_X1 U10227 ( .A(n8497), .ZN(n8479) );
  NAND2_X1 U10228 ( .A1(n8477), .A2(n8476), .ZN(n8478) );
  NAND2_X1 U10229 ( .A1(n8479), .A2(n8478), .ZN(n8480) );
  INV_X1 U10230 ( .A(n8483), .ZN(n8495) );
  INV_X1 U10231 ( .A(n8485), .ZN(n8488) );
  OAI211_X1 U10232 ( .C1(n8489), .C2(n8488), .A(n8487), .B(n8486), .ZN(n8492)
         );
  OAI211_X1 U10233 ( .C1(n8497), .C2(n8496), .A(n8495), .B(n8494), .ZN(n8498)
         );
  INV_X1 U10234 ( .A(n8498), .ZN(n8499) );
  NAND3_X1 U10235 ( .A1(n8501), .A2(n8500), .A3(n8570), .ZN(n8502) );
  INV_X1 U10236 ( .A(n8506), .ZN(n8504) );
  OAI21_X1 U10237 ( .B1(n8504), .B2(n8503), .A(n8570), .ZN(n8505) );
  MUX2_X1 U10238 ( .A(n8507), .B(n8506), .S(n8577), .Z(n8508) );
  MUX2_X1 U10239 ( .A(n8511), .B(n8510), .S(n8570), .Z(n8512) );
  MUX2_X1 U10240 ( .A(n8516), .B(n8515), .S(n8577), .Z(n8517) );
  MUX2_X1 U10241 ( .A(n8519), .B(n8518), .S(n8577), .Z(n8521) );
  AOI21_X1 U10242 ( .B1(n8530), .B2(n8523), .A(n8570), .ZN(n8524) );
  AOI21_X1 U10243 ( .B1(n8532), .B2(n8533), .A(n4817), .ZN(n8527) );
  NAND3_X1 U10244 ( .A1(n8528), .A2(n8541), .A3(n8535), .ZN(n8529) );
  NAND2_X1 U10245 ( .A1(n8537), .A2(n8536), .ZN(n8540) );
  INV_X1 U10246 ( .A(n8542), .ZN(n8822) );
  OR3_X1 U10247 ( .A1(n9023), .A2(n8543), .A3(n8577), .ZN(n8544) );
  NAND2_X1 U10248 ( .A1(n8545), .A2(n8544), .ZN(n8553) );
  NAND2_X1 U10249 ( .A1(n8553), .A2(n8552), .ZN(n8550) );
  AND2_X1 U10250 ( .A1(n8554), .A2(n8546), .ZN(n8549) );
  INV_X1 U10251 ( .A(n8547), .ZN(n8548) );
  INV_X1 U10252 ( .A(n8554), .ZN(n8555) );
  AOI21_X1 U10253 ( .B1(n8557), .B2(n8556), .A(n8555), .ZN(n8558) );
  MUX2_X1 U10254 ( .A(n8561), .B(n8560), .S(n8577), .Z(n8562) );
  MUX2_X1 U10255 ( .A(n8565), .B(n8564), .S(n8570), .Z(n8566) );
  NOR2_X1 U10256 ( .A1(n8567), .A2(n8566), .ZN(n8568) );
  INV_X1 U10257 ( .A(n8569), .ZN(n8573) );
  MUX2_X1 U10258 ( .A(n8781), .B(n8571), .S(n8570), .Z(n8572) );
  OR2_X1 U10259 ( .A1(n8573), .A2(n8572), .ZN(n8574) );
  AOI21_X1 U10260 ( .B1(n8580), .B2(n8607), .A(n8577), .ZN(n8578) );
  NAND4_X1 U10261 ( .A1(n8583), .A2(n8582), .A3(n8581), .A4(n8580), .ZN(n8584)
         );
  NAND2_X1 U10262 ( .A1(n8598), .A2(n8586), .ZN(n8588) );
  NOR2_X1 U10263 ( .A1(n8595), .A2(n8587), .ZN(n8599) );
  NAND2_X1 U10264 ( .A1(n8588), .A2(n8599), .ZN(n8604) );
  OAI211_X1 U10265 ( .C1(n8592), .C2(n8595), .A(n8591), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8603) );
  NAND3_X1 U10266 ( .A1(n8598), .A2(n8597), .A3(n8586), .ZN(n8602) );
  NAND2_X1 U10267 ( .A1(n8600), .A2(n8599), .ZN(n8601) );
  NAND4_X1 U10268 ( .A1(n8602), .A2(n8603), .A3(n8604), .A4(n8601), .ZN(
        P2_U3296) );
  MUX2_X1 U10269 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8605), .S(P2_U3893), .Z(
        P2_U3521) );
  INV_X1 U10270 ( .A(n8606), .ZN(n8782) );
  MUX2_X1 U10271 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8782), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10272 ( .A(n8607), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8756), .Z(
        P2_U3519) );
  MUX2_X1 U10273 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8781), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10274 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8802), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10275 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8608), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10276 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8801), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10277 ( .A(n8609), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8756), .Z(
        P2_U3514) );
  MUX2_X1 U10278 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8839), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10279 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8610), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10280 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8838), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10281 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8611), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10282 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8899), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10283 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8907), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10284 ( .A(n8916), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8756), .Z(
        P2_U3507) );
  MUX2_X1 U10285 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8926), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10286 ( .A(n8915), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8756), .Z(
        P2_U3505) );
  MUX2_X1 U10287 ( .A(n8925), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8756), .Z(
        P2_U3504) );
  MUX2_X1 U10288 ( .A(n8612), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8756), .Z(
        P2_U3503) );
  MUX2_X1 U10289 ( .A(n8613), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8756), .Z(
        P2_U3502) );
  MUX2_X1 U10290 ( .A(n8614), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8756), .Z(
        P2_U3501) );
  MUX2_X1 U10291 ( .A(n8615), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8756), .Z(
        P2_U3500) );
  MUX2_X1 U10292 ( .A(n8616), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8756), .Z(
        P2_U3499) );
  MUX2_X1 U10293 ( .A(n8617), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8756), .Z(
        P2_U3498) );
  MUX2_X1 U10294 ( .A(n10169), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8756), .Z(
        P2_U3497) );
  MUX2_X1 U10295 ( .A(n8618), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8756), .Z(
        P2_U3496) );
  MUX2_X1 U10296 ( .A(n7255), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8756), .Z(
        P2_U3495) );
  MUX2_X1 U10297 ( .A(n6508), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8756), .Z(
        P2_U3494) );
  MUX2_X1 U10298 ( .A(n8619), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8756), .Z(
        P2_U3493) );
  MUX2_X1 U10299 ( .A(n8620), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8756), .Z(
        P2_U3492) );
  MUX2_X1 U10300 ( .A(n8621), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8756), .Z(
        P2_U3491) );
  INV_X1 U10301 ( .A(n8622), .ZN(n8627) );
  NOR3_X1 U10302 ( .A1(n8625), .A2(n8624), .A3(n8623), .ZN(n8626) );
  OAI21_X1 U10303 ( .B1(n8627), .B2(n8626), .A(n5444), .ZN(n8645) );
  OAI21_X1 U10304 ( .B1(n8759), .B2(n10357), .A(n8628), .ZN(n8636) );
  INV_X1 U10305 ( .A(n8629), .ZN(n8634) );
  NAND3_X1 U10306 ( .A1(n8632), .A2(n8631), .A3(n8630), .ZN(n8633) );
  AOI21_X1 U10307 ( .B1(n8634), .B2(n8633), .A(n8760), .ZN(n8635) );
  AOI211_X1 U10308 ( .C1(n8718), .C2(n8637), .A(n8636), .B(n8635), .ZN(n8644)
         );
  AND3_X1 U10309 ( .A1(n8640), .A2(n8639), .A3(n8638), .ZN(n8641) );
  OAI21_X1 U10310 ( .B1(n8642), .B2(n8641), .A(n8750), .ZN(n8643) );
  NAND3_X1 U10311 ( .A1(n8645), .A2(n8644), .A3(n8643), .ZN(P2_U3192) );
  AOI21_X1 U10312 ( .B1(n8647), .B2(n8646), .A(n4575), .ZN(n8661) );
  INV_X1 U10313 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8649) );
  OAI21_X1 U10314 ( .B1(n8759), .B2(n8649), .A(n8648), .ZN(n8655) );
  NAND3_X1 U10315 ( .A1(n8652), .A2(n8651), .A3(n8650), .ZN(n8653) );
  AOI21_X1 U10316 ( .B1(n8678), .B2(n8653), .A(n8760), .ZN(n8654) );
  AOI211_X1 U10317 ( .C1(n8718), .C2(n8656), .A(n8655), .B(n8654), .ZN(n8660)
         );
  OAI21_X1 U10318 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n8657), .A(n8674), .ZN(
        n8658) );
  NAND2_X1 U10319 ( .A1(n8658), .A2(n8750), .ZN(n8659) );
  OAI211_X1 U10320 ( .C1(n8661), .C2(n8768), .A(n8660), .B(n8659), .ZN(
        P2_U3195) );
  INV_X1 U10321 ( .A(n8662), .ZN(n8667) );
  NOR3_X1 U10322 ( .A1(n4575), .A2(n8664), .A3(n8663), .ZN(n8666) );
  OAI21_X1 U10323 ( .B1(n8667), .B2(n8666), .A(n5444), .ZN(n8684) );
  INV_X1 U10324 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8669) );
  OAI21_X1 U10325 ( .B1(n8759), .B2(n8669), .A(n8668), .ZN(n8670) );
  AOI21_X1 U10326 ( .B1(n8671), .B2(n8718), .A(n8670), .ZN(n8683) );
  AND3_X1 U10327 ( .A1(n8674), .A2(n8673), .A3(n8672), .ZN(n8675) );
  OAI21_X1 U10328 ( .B1(n4528), .B2(n8675), .A(n8750), .ZN(n8682) );
  AND3_X1 U10329 ( .A1(n8678), .A2(n8677), .A3(n8676), .ZN(n8679) );
  OAI21_X1 U10330 ( .B1(n8680), .B2(n8679), .A(n8733), .ZN(n8681) );
  NAND4_X1 U10331 ( .A1(n8684), .A2(n8683), .A3(n8682), .A4(n8681), .ZN(
        P2_U3196) );
  INV_X1 U10332 ( .A(n8685), .ZN(n8686) );
  AOI21_X1 U10333 ( .B1(n10373), .B2(n8687), .A(n8686), .ZN(n8701) );
  OAI21_X1 U10334 ( .B1(n8759), .B2(n8688), .A(n10277), .ZN(n8694) );
  AOI21_X1 U10335 ( .B1(n8691), .B2(n8690), .A(n8689), .ZN(n8692) );
  NOR2_X1 U10336 ( .A1(n8692), .A2(n8760), .ZN(n8693) );
  AOI211_X1 U10337 ( .C1(n8718), .C2(n8695), .A(n8694), .B(n8693), .ZN(n8700)
         );
  OAI21_X1 U10338 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n8697), .A(n8696), .ZN(
        n8698) );
  NAND2_X1 U10339 ( .A1(n8698), .A2(n8750), .ZN(n8699) );
  OAI211_X1 U10340 ( .C1(n8701), .C2(n8768), .A(n8700), .B(n8699), .ZN(
        P2_U3197) );
  OAI21_X1 U10341 ( .B1(n8704), .B2(n8703), .A(n8702), .ZN(n8723) );
  INV_X1 U10342 ( .A(n8705), .ZN(n8706) );
  NOR2_X1 U10343 ( .A1(n8707), .A2(n8706), .ZN(n8708) );
  XNOR2_X1 U10344 ( .A(n8709), .B(n8708), .ZN(n8721) );
  OAI21_X1 U10345 ( .B1(n8712), .B2(n8711), .A(n8710), .ZN(n8713) );
  NAND2_X1 U10346 ( .A1(n8713), .A2(n8750), .ZN(n8720) );
  OAI21_X1 U10347 ( .B1(n8759), .B2(n8715), .A(n8714), .ZN(n8716) );
  AOI21_X1 U10348 ( .B1(n8718), .B2(n8717), .A(n8716), .ZN(n8719) );
  OAI211_X1 U10349 ( .C1(n8760), .C2(n8721), .A(n8720), .B(n8719), .ZN(n8722)
         );
  AOI21_X1 U10350 ( .B1(n5444), .B2(n8723), .A(n8722), .ZN(n8724) );
  INV_X1 U10351 ( .A(n8724), .ZN(P2_U3198) );
  AOI21_X1 U10352 ( .B1(n10471), .B2(n8725), .A(n8749), .ZN(n8740) );
  XNOR2_X1 U10353 ( .A(n8727), .B(n8726), .ZN(n8734) );
  NAND2_X1 U10354 ( .A1(n8728), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8729) );
  OAI211_X1 U10355 ( .C1(n8755), .C2(n8731), .A(n8730), .B(n8729), .ZN(n8732)
         );
  AOI21_X1 U10356 ( .B1(n8734), .B2(n8733), .A(n8732), .ZN(n8738) );
  OAI21_X1 U10357 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8735), .A(n8744), .ZN(
        n8736) );
  NAND2_X1 U10358 ( .A1(n8736), .A2(n5444), .ZN(n8737) );
  OAI211_X1 U10359 ( .C1(n8740), .C2(n8739), .A(n8738), .B(n8737), .ZN(
        P2_U3199) );
  INV_X1 U10360 ( .A(n8741), .ZN(n8742) );
  NAND3_X1 U10361 ( .A1(n8744), .A2(n8743), .A3(n8742), .ZN(n8745) );
  AND2_X1 U10362 ( .A1(n8746), .A2(n8745), .ZN(n8769) );
  NOR3_X1 U10363 ( .A1(n8749), .A2(n8748), .A3(n8747), .ZN(n8751) );
  OAI21_X1 U10364 ( .B1(n4484), .B2(n8751), .A(n8750), .ZN(n8767) );
  INV_X1 U10365 ( .A(n8752), .ZN(n8753) );
  NOR2_X1 U10366 ( .A1(n8754), .A2(n8753), .ZN(n8761) );
  INV_X1 U10367 ( .A(n8761), .ZN(n8757) );
  OAI21_X1 U10368 ( .B1(n8757), .B2(n8756), .A(n8755), .ZN(n8764) );
  INV_X1 U10369 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10333) );
  OAI21_X1 U10370 ( .B1(n8759), .B2(n10333), .A(n8758), .ZN(n8763) );
  NOR3_X1 U10371 ( .A1(n8761), .A2(n8765), .A3(n8760), .ZN(n8762) );
  AOI211_X1 U10372 ( .C1(n8765), .C2(n8764), .A(n8763), .B(n8762), .ZN(n8766)
         );
  OAI211_X1 U10373 ( .C1(n8769), .C2(n8768), .A(n8767), .B(n8766), .ZN(
        P2_U3200) );
  INV_X1 U10374 ( .A(n8770), .ZN(n8771) );
  AOI21_X1 U10375 ( .B1(n8991), .B2(n10181), .A(n8773), .ZN(n8776) );
  NAND2_X1 U10376 ( .A1(n10183), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8774) );
  OAI211_X1 U10377 ( .C1(n8993), .C2(n8873), .A(n8776), .B(n8774), .ZN(
        P2_U3202) );
  INV_X1 U10378 ( .A(n8994), .ZN(n8777) );
  NAND2_X1 U10379 ( .A1(n10183), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8775) );
  OAI211_X1 U10380 ( .C1(n8777), .C2(n8873), .A(n8776), .B(n8775), .ZN(
        P2_U3203) );
  XNOR2_X1 U10381 ( .A(n8778), .B(n8779), .ZN(n8939) );
  INV_X1 U10382 ( .A(n8939), .ZN(n8788) );
  AOI22_X1 U10383 ( .A1(n8782), .A2(n10168), .B1(n10167), .B2(n8781), .ZN(
        n8783) );
  AOI22_X1 U10384 ( .A1(n8784), .A2(n10175), .B1(n10183), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8785) );
  OAI21_X1 U10385 ( .B1(n8998), .B2(n8873), .A(n8785), .ZN(n8786) );
  AOI21_X1 U10386 ( .B1(n8938), .B2(n10181), .A(n8786), .ZN(n8787) );
  OAI21_X1 U10387 ( .B1(n8788), .B2(n8934), .A(n8787), .ZN(P2_U3205) );
  XNOR2_X1 U10388 ( .A(n8789), .B(n8790), .ZN(n9004) );
  INV_X1 U10389 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8794) );
  XNOR2_X1 U10390 ( .A(n8791), .B(n8790), .ZN(n8792) );
  OAI222_X1 U10391 ( .A1(n8881), .A2(n8793), .B1(n8883), .B2(n8815), .C1(
        n10185), .C2(n8792), .ZN(n8946) );
  INV_X1 U10392 ( .A(n8946), .ZN(n8999) );
  MUX2_X1 U10393 ( .A(n8794), .B(n8999), .S(n10181), .Z(n8797) );
  AOI22_X1 U10394 ( .A1(n9001), .A2(n10178), .B1(n10175), .B2(n8795), .ZN(
        n8796) );
  OAI211_X1 U10395 ( .C1(n9004), .C2(n8934), .A(n8797), .B(n8796), .ZN(
        P2_U3207) );
  XNOR2_X1 U10396 ( .A(n8798), .B(n8799), .ZN(n9010) );
  XNOR2_X1 U10397 ( .A(n8800), .B(n8799), .ZN(n8803) );
  AOI222_X1 U10398 ( .A1(n10171), .A2(n8803), .B1(n8802), .B2(n10168), .C1(
        n8801), .C2(n10167), .ZN(n9005) );
  AOI22_X1 U10399 ( .A1(n9007), .A2(n8805), .B1(n10175), .B2(n8804), .ZN(n8806) );
  AOI21_X1 U10400 ( .B1(n9005), .B2(n8806), .A(n10183), .ZN(n8807) );
  AOI21_X1 U10401 ( .B1(n10183), .B2(P2_REG2_REG_25__SCAN_IN), .A(n8807), .ZN(
        n8808) );
  OAI21_X1 U10402 ( .B1(n9010), .B2(n8934), .A(n8808), .ZN(P2_U3208) );
  NAND2_X1 U10403 ( .A1(n8809), .A2(n8810), .ZN(n8811) );
  XOR2_X1 U10404 ( .A(n8812), .B(n8811), .Z(n9012) );
  XNOR2_X1 U10405 ( .A(n8813), .B(n8812), .ZN(n8814) );
  OAI222_X1 U10406 ( .A1(n8881), .A2(n8815), .B1(n8883), .B2(n8826), .C1(
        n10185), .C2(n8814), .ZN(n9013) );
  OAI22_X1 U10407 ( .A1(n9011), .A2(n8928), .B1(n8816), .B2(n8885), .ZN(n8817)
         );
  OAI21_X1 U10408 ( .B1(n9013), .B2(n8817), .A(n10181), .ZN(n8819) );
  NAND2_X1 U10409 ( .A1(n10183), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8818) );
  OAI211_X1 U10410 ( .C1(n9012), .C2(n8934), .A(n8819), .B(n8818), .ZN(
        P2_U3209) );
  XNOR2_X1 U10411 ( .A(n8820), .B(n8822), .ZN(n9025) );
  INV_X1 U10412 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8828) );
  NAND3_X1 U10413 ( .A1(n8836), .A2(n8822), .A3(n8821), .ZN(n8823) );
  AND2_X1 U10414 ( .A1(n8824), .A2(n8823), .ZN(n8825) );
  OAI222_X1 U10415 ( .A1(n8881), .A2(n8826), .B1(n8883), .B2(n8854), .C1(
        n10185), .C2(n8825), .ZN(n9021) );
  INV_X1 U10416 ( .A(n9021), .ZN(n8827) );
  MUX2_X1 U10417 ( .A(n8828), .B(n8827), .S(n10181), .Z(n8831) );
  AOI22_X1 U10418 ( .A1(n9023), .A2(n10178), .B1(n10175), .B2(n8829), .ZN(
        n8830) );
  OAI211_X1 U10419 ( .C1(n9025), .C2(n8934), .A(n8831), .B(n8830), .ZN(
        P2_U3211) );
  XOR2_X1 U10420 ( .A(n8832), .B(n8834), .Z(n9031) );
  INV_X1 U10421 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8841) );
  NOR2_X1 U10422 ( .A1(n8878), .A2(n6518), .ZN(n8877) );
  NAND3_X1 U10423 ( .A1(n8864), .A2(n8849), .A3(n8850), .ZN(n8848) );
  NAND3_X1 U10424 ( .A1(n8848), .A2(n4728), .A3(n8835), .ZN(n8837) );
  NAND2_X1 U10425 ( .A1(n8837), .A2(n8836), .ZN(n8840) );
  AOI222_X1 U10426 ( .A1(n10171), .A2(n8840), .B1(n8839), .B2(n10168), .C1(
        n8838), .C2(n10167), .ZN(n9026) );
  MUX2_X1 U10427 ( .A(n8841), .B(n9026), .S(n10181), .Z(n8844) );
  AOI22_X1 U10428 ( .A1(n9028), .A2(n10178), .B1(n10175), .B2(n8842), .ZN(
        n8843) );
  OAI211_X1 U10429 ( .C1(n9031), .C2(n8934), .A(n8844), .B(n8843), .ZN(
        P2_U3212) );
  INV_X1 U10430 ( .A(n8865), .ZN(n8860) );
  NAND2_X1 U10431 ( .A1(n8861), .A2(n8860), .ZN(n8859) );
  NAND2_X1 U10432 ( .A1(n8859), .A2(n8846), .ZN(n8847) );
  XOR2_X1 U10433 ( .A(n8849), .B(n8847), .Z(n9037) );
  INV_X1 U10434 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8855) );
  INV_X1 U10435 ( .A(n8848), .ZN(n8852) );
  AOI21_X1 U10436 ( .B1(n8864), .B2(n8850), .A(n8849), .ZN(n8851) );
  NOR2_X1 U10437 ( .A1(n8852), .A2(n8851), .ZN(n8853) );
  OAI222_X1 U10438 ( .A1(n8881), .A2(n8854), .B1(n8883), .B2(n8880), .C1(
        n10185), .C2(n8853), .ZN(n8962) );
  INV_X1 U10439 ( .A(n8962), .ZN(n9032) );
  MUX2_X1 U10440 ( .A(n8855), .B(n9032), .S(n10181), .Z(n8858) );
  AOI22_X1 U10441 ( .A1(n9034), .A2(n10178), .B1(n10175), .B2(n8856), .ZN(
        n8857) );
  OAI211_X1 U10442 ( .C1(n9037), .C2(n8934), .A(n8858), .B(n8857), .ZN(
        P2_U3213) );
  OAI21_X1 U10443 ( .B1(n8861), .B2(n8860), .A(n8859), .ZN(n9041) );
  INV_X1 U10444 ( .A(n8862), .ZN(n8863) );
  NOR2_X1 U10445 ( .A1(n8877), .A2(n8863), .ZN(n8866) );
  OAI211_X1 U10446 ( .C1(n8866), .C2(n8865), .A(n10171), .B(n8864), .ZN(n8869)
         );
  OR2_X1 U10447 ( .A1(n8867), .A2(n8881), .ZN(n8868) );
  OAI211_X1 U10448 ( .C1(n8870), .C2(n8883), .A(n8869), .B(n8868), .ZN(n8966)
         );
  AOI22_X1 U10449 ( .A1(n10183), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n10175), 
        .B2(n8871), .ZN(n8872) );
  OAI21_X1 U10450 ( .B1(n8874), .B2(n8873), .A(n8872), .ZN(n8875) );
  AOI21_X1 U10451 ( .B1(n8966), .B2(n10181), .A(n8875), .ZN(n8876) );
  OAI21_X1 U10452 ( .B1(n8934), .B2(n9041), .A(n8876), .ZN(P2_U3214) );
  AOI21_X1 U10453 ( .B1(n6518), .B2(n8878), .A(n8877), .ZN(n8879) );
  OAI222_X1 U10454 ( .A1(n8883), .A2(n8882), .B1(n8881), .B2(n8880), .C1(
        n10185), .C2(n8879), .ZN(n8971) );
  INV_X1 U10455 ( .A(n8971), .ZN(n8895) );
  INV_X1 U10456 ( .A(n8884), .ZN(n8886) );
  OAI22_X1 U10457 ( .A1(n10181), .A2(n8887), .B1(n8886), .B2(n8885), .ZN(n8893) );
  INV_X1 U10458 ( .A(n8888), .ZN(n8891) );
  AND2_X1 U10459 ( .A1(n8890), .A2(n8889), .ZN(n8970) );
  NOR3_X1 U10460 ( .A1(n8891), .A2(n8970), .A3(n8934), .ZN(n8892) );
  AOI211_X1 U10461 ( .C1(n10178), .C2(n8969), .A(n8893), .B(n8892), .ZN(n8894)
         );
  OAI21_X1 U10462 ( .B1(n8895), .B2(n10183), .A(n8894), .ZN(P2_U3215) );
  XNOR2_X1 U10463 ( .A(n8896), .B(n8897), .ZN(n9052) );
  XNOR2_X1 U10464 ( .A(n8898), .B(n8897), .ZN(n8900) );
  AOI222_X1 U10465 ( .A1(n10171), .A2(n8900), .B1(n8899), .B2(n10168), .C1(
        n8916), .C2(n10167), .ZN(n9047) );
  MUX2_X1 U10466 ( .A(n10471), .B(n9047), .S(n10181), .Z(n8903) );
  AOI22_X1 U10467 ( .A1(n9049), .A2(n10178), .B1(n10175), .B2(n8901), .ZN(
        n8902) );
  OAI211_X1 U10468 ( .C1(n9052), .C2(n8934), .A(n8903), .B(n8902), .ZN(
        P2_U3216) );
  XNOR2_X1 U10469 ( .A(n8904), .B(n8905), .ZN(n9058) );
  XNOR2_X1 U10470 ( .A(n8906), .B(n8905), .ZN(n8908) );
  AOI222_X1 U10471 ( .A1(n10171), .A2(n8908), .B1(n8907), .B2(n10168), .C1(
        n8926), .C2(n10167), .ZN(n9053) );
  MUX2_X1 U10472 ( .A(n8909), .B(n9053), .S(n10181), .Z(n8912) );
  AOI22_X1 U10473 ( .A1(n9055), .A2(n10178), .B1(n10175), .B2(n8910), .ZN(
        n8911) );
  OAI211_X1 U10474 ( .C1(n9058), .C2(n8934), .A(n8912), .B(n8911), .ZN(
        P2_U3217) );
  XNOR2_X1 U10475 ( .A(n8913), .B(n5052), .ZN(n9064) );
  INV_X1 U10476 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8918) );
  XNOR2_X1 U10477 ( .A(n8914), .B(n5052), .ZN(n8917) );
  AOI222_X1 U10478 ( .A1(n10171), .A2(n8917), .B1(n8916), .B2(n10168), .C1(
        n8915), .C2(n10167), .ZN(n9059) );
  MUX2_X1 U10479 ( .A(n8918), .B(n9059), .S(n10181), .Z(n8921) );
  AOI22_X1 U10480 ( .A1(n9061), .A2(n10178), .B1(n10175), .B2(n8919), .ZN(
        n8920) );
  OAI211_X1 U10481 ( .C1(n9064), .C2(n8934), .A(n8921), .B(n8920), .ZN(
        P2_U3218) );
  XNOR2_X1 U10482 ( .A(n8922), .B(n8923), .ZN(n9071) );
  XNOR2_X1 U10483 ( .A(n8924), .B(n8923), .ZN(n8927) );
  AOI222_X1 U10484 ( .A1(n10171), .A2(n8927), .B1(n8926), .B2(n10168), .C1(
        n8925), .C2(n10167), .ZN(n9065) );
  OAI21_X1 U10485 ( .B1(n8929), .B2(n8928), .A(n9065), .ZN(n8930) );
  NAND2_X1 U10486 ( .A1(n8930), .A2(n10181), .ZN(n8933) );
  AOI22_X1 U10487 ( .A1(n10183), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n10175), 
        .B2(n8931), .ZN(n8932) );
  OAI211_X1 U10488 ( .C1(n9071), .C2(n8934), .A(n8933), .B(n8932), .ZN(
        P2_U3219) );
  NAND2_X1 U10489 ( .A1(n6586), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8935) );
  NAND2_X1 U10490 ( .A1(n8991), .A2(n10245), .ZN(n8936) );
  OAI211_X1 U10491 ( .C1(n8993), .C2(n8974), .A(n8935), .B(n8936), .ZN(
        P2_U3490) );
  NAND2_X1 U10492 ( .A1(n8994), .A2(n8983), .ZN(n8937) );
  OAI211_X1 U10493 ( .C1(n10245), .C2(n10426), .A(n8937), .B(n8936), .ZN(
        P2_U3489) );
  OAI21_X1 U10494 ( .B1(n8998), .B2(n8974), .A(n8940), .ZN(P2_U3487) );
  MUX2_X1 U10495 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8941), .S(n10245), .Z(
        n8945) );
  OAI22_X1 U10496 ( .A1(n8943), .A2(n8986), .B1(n8942), .B2(n8974), .ZN(n8944)
         );
  OR2_X1 U10497 ( .A1(n8945), .A2(n8944), .ZN(P2_U3486) );
  MUX2_X1 U10498 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8946), .S(n10245), .Z(
        n8949) );
  OAI22_X1 U10499 ( .A1(n9004), .A2(n8986), .B1(n8947), .B2(n8974), .ZN(n8948)
         );
  OR2_X1 U10500 ( .A1(n8949), .A2(n8948), .ZN(P2_U3485) );
  INV_X1 U10501 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8950) );
  MUX2_X1 U10502 ( .A(n8950), .B(n9005), .S(n10245), .Z(n8952) );
  NAND2_X1 U10503 ( .A1(n9007), .A2(n8983), .ZN(n8951) );
  OAI211_X1 U10504 ( .C1(n9010), .C2(n8986), .A(n8952), .B(n8951), .ZN(
        P2_U3484) );
  OAI22_X1 U10505 ( .A1(n9012), .A2(n8986), .B1(n9011), .B2(n8974), .ZN(n8954)
         );
  MUX2_X1 U10506 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9013), .S(n10245), .Z(
        n8953) );
  OR2_X1 U10507 ( .A1(n8954), .A2(n8953), .ZN(P2_U3483) );
  OAI22_X1 U10508 ( .A1(n9017), .A2(n8986), .B1(n9016), .B2(n8974), .ZN(n8956)
         );
  MUX2_X1 U10509 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9018), .S(n10245), .Z(
        n8955) );
  OR2_X1 U10510 ( .A1(n8956), .A2(n8955), .ZN(P2_U3482) );
  MUX2_X1 U10511 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9021), .S(n10245), .Z(
        n8957) );
  AOI21_X1 U10512 ( .B1(n8983), .B2(n9023), .A(n8957), .ZN(n8958) );
  OAI21_X1 U10513 ( .B1(n9025), .B2(n8986), .A(n8958), .ZN(P2_U3481) );
  INV_X1 U10514 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8959) );
  MUX2_X1 U10515 ( .A(n8959), .B(n9026), .S(n10245), .Z(n8961) );
  NAND2_X1 U10516 ( .A1(n9028), .A2(n8983), .ZN(n8960) );
  OAI211_X1 U10517 ( .C1(n9031), .C2(n8986), .A(n8961), .B(n8960), .ZN(
        P2_U3480) );
  MUX2_X1 U10518 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8962), .S(n10245), .Z(
        n8965) );
  OAI22_X1 U10519 ( .A1(n9037), .A2(n8986), .B1(n8963), .B2(n8974), .ZN(n8964)
         );
  OR2_X1 U10520 ( .A1(n8965), .A2(n8964), .ZN(P2_U3479) );
  AOI21_X1 U10521 ( .B1(n10189), .B2(n8967), .A(n8966), .ZN(n9038) );
  MUX2_X1 U10522 ( .A(n10532), .B(n9038), .S(n10245), .Z(n8968) );
  OAI21_X1 U10523 ( .B1(n8986), .B2(n9041), .A(n8968), .ZN(P2_U3478) );
  INV_X1 U10524 ( .A(n8969), .ZN(n9046) );
  NOR2_X1 U10525 ( .A1(n8970), .A2(n10225), .ZN(n8972) );
  AOI21_X1 U10526 ( .B1(n8972), .B2(n8888), .A(n8971), .ZN(n9042) );
  MUX2_X1 U10527 ( .A(n10504), .B(n9042), .S(n10245), .Z(n8973) );
  OAI21_X1 U10528 ( .B1(n9046), .B2(n8974), .A(n8973), .ZN(P2_U3477) );
  INV_X1 U10529 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8975) );
  MUX2_X1 U10530 ( .A(n8975), .B(n9047), .S(n10245), .Z(n8977) );
  NAND2_X1 U10531 ( .A1(n9049), .A2(n8983), .ZN(n8976) );
  OAI211_X1 U10532 ( .C1(n9052), .C2(n8986), .A(n8977), .B(n8976), .ZN(
        P2_U3476) );
  MUX2_X1 U10533 ( .A(n10563), .B(n9053), .S(n10245), .Z(n8979) );
  NAND2_X1 U10534 ( .A1(n9055), .A2(n8983), .ZN(n8978) );
  OAI211_X1 U10535 ( .C1(n9058), .C2(n8986), .A(n8979), .B(n8978), .ZN(
        P2_U3475) );
  MUX2_X1 U10536 ( .A(n10373), .B(n9059), .S(n10245), .Z(n8981) );
  NAND2_X1 U10537 ( .A1(n9061), .A2(n8983), .ZN(n8980) );
  OAI211_X1 U10538 ( .C1(n9064), .C2(n8986), .A(n8981), .B(n8980), .ZN(
        P2_U3474) );
  MUX2_X1 U10539 ( .A(n8982), .B(n9065), .S(n10245), .Z(n8985) );
  NAND2_X1 U10540 ( .A1(n9067), .A2(n8983), .ZN(n8984) );
  OAI211_X1 U10541 ( .C1(n9071), .C2(n8986), .A(n8985), .B(n8984), .ZN(
        P2_U3473) );
  AOI21_X1 U10542 ( .B1(n10189), .B2(n8988), .A(n8987), .ZN(n8989) );
  OAI21_X1 U10543 ( .B1(n10225), .B2(n8990), .A(n8989), .ZN(n9072) );
  MUX2_X1 U10544 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9072), .S(n10245), .Z(
        P2_U3470) );
  NAND2_X1 U10545 ( .A1(n10229), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8992) );
  NAND2_X1 U10546 ( .A1(n8991), .A2(n10230), .ZN(n8995) );
  OAI211_X1 U10547 ( .C1(n8993), .C2(n9045), .A(n8992), .B(n8995), .ZN(
        P2_U3458) );
  NAND2_X1 U10548 ( .A1(n8994), .A2(n9066), .ZN(n8996) );
  OAI211_X1 U10549 ( .C1(n10230), .C2(n10561), .A(n8996), .B(n8995), .ZN(
        P2_U3457) );
  OAI21_X1 U10550 ( .B1(n8998), .B2(n9045), .A(n8997), .ZN(P2_U3455) );
  MUX2_X1 U10551 ( .A(n9000), .B(n8999), .S(n10230), .Z(n9003) );
  NAND2_X1 U10552 ( .A1(n9001), .A2(n9066), .ZN(n9002) );
  OAI211_X1 U10553 ( .C1(n9004), .C2(n9070), .A(n9003), .B(n9002), .ZN(
        P2_U3453) );
  MUX2_X1 U10554 ( .A(n9006), .B(n9005), .S(n10230), .Z(n9009) );
  NAND2_X1 U10555 ( .A1(n9007), .A2(n9066), .ZN(n9008) );
  OAI211_X1 U10556 ( .C1(n9010), .C2(n9070), .A(n9009), .B(n9008), .ZN(
        P2_U3452) );
  OAI22_X1 U10557 ( .A1(n9012), .A2(n9070), .B1(n9011), .B2(n9045), .ZN(n9015)
         );
  MUX2_X1 U10558 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9013), .S(n10230), .Z(
        n9014) );
  OR2_X1 U10559 ( .A1(n9015), .A2(n9014), .ZN(P2_U3451) );
  OAI22_X1 U10560 ( .A1(n9017), .A2(n9070), .B1(n9016), .B2(n9045), .ZN(n9020)
         );
  MUX2_X1 U10561 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9018), .S(n10230), .Z(
        n9019) );
  OR2_X1 U10562 ( .A1(n9020), .A2(n9019), .ZN(P2_U3450) );
  MUX2_X1 U10563 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9021), .S(n10230), .Z(
        n9022) );
  AOI21_X1 U10564 ( .B1(n9066), .B2(n9023), .A(n9022), .ZN(n9024) );
  OAI21_X1 U10565 ( .B1(n9025), .B2(n9070), .A(n9024), .ZN(P2_U3449) );
  MUX2_X1 U10566 ( .A(n9027), .B(n9026), .S(n10230), .Z(n9030) );
  NAND2_X1 U10567 ( .A1(n9028), .A2(n9066), .ZN(n9029) );
  OAI211_X1 U10568 ( .C1(n9031), .C2(n9070), .A(n9030), .B(n9029), .ZN(
        P2_U3448) );
  MUX2_X1 U10569 ( .A(n9033), .B(n9032), .S(n10230), .Z(n9036) );
  NAND2_X1 U10570 ( .A1(n9034), .A2(n9066), .ZN(n9035) );
  OAI211_X1 U10571 ( .C1(n9037), .C2(n9070), .A(n9036), .B(n9035), .ZN(
        P2_U3447) );
  INV_X1 U10572 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9039) );
  MUX2_X1 U10573 ( .A(n9039), .B(n9038), .S(n10230), .Z(n9040) );
  OAI21_X1 U10574 ( .B1(n9041), .B2(n9070), .A(n9040), .ZN(P2_U3446) );
  INV_X1 U10575 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9043) );
  MUX2_X1 U10576 ( .A(n9043), .B(n9042), .S(n10230), .Z(n9044) );
  OAI21_X1 U10577 ( .B1(n9046), .B2(n9045), .A(n9044), .ZN(P2_U3444) );
  INV_X1 U10578 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9048) );
  MUX2_X1 U10579 ( .A(n9048), .B(n9047), .S(n10230), .Z(n9051) );
  NAND2_X1 U10580 ( .A1(n9049), .A2(n9066), .ZN(n9050) );
  OAI211_X1 U10581 ( .C1(n9052), .C2(n9070), .A(n9051), .B(n9050), .ZN(
        P2_U3441) );
  INV_X1 U10582 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9054) );
  MUX2_X1 U10583 ( .A(n9054), .B(n9053), .S(n10230), .Z(n9057) );
  NAND2_X1 U10584 ( .A1(n9055), .A2(n9066), .ZN(n9056) );
  OAI211_X1 U10585 ( .C1(n9058), .C2(n9070), .A(n9057), .B(n9056), .ZN(
        P2_U3438) );
  INV_X1 U10586 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9060) );
  MUX2_X1 U10587 ( .A(n9060), .B(n9059), .S(n10230), .Z(n9063) );
  NAND2_X1 U10588 ( .A1(n9061), .A2(n9066), .ZN(n9062) );
  OAI211_X1 U10589 ( .C1(n9064), .C2(n9070), .A(n9063), .B(n9062), .ZN(
        P2_U3435) );
  MUX2_X1 U10590 ( .A(n10517), .B(n9065), .S(n10230), .Z(n9069) );
  NAND2_X1 U10591 ( .A1(n9067), .A2(n9066), .ZN(n9068) );
  OAI211_X1 U10592 ( .C1(n9071), .C2(n9070), .A(n9069), .B(n9068), .ZN(
        P2_U3432) );
  MUX2_X1 U10593 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n9072), .S(n10230), .Z(
        P2_U3423) );
  MUX2_X1 U10594 ( .A(n9074), .B(P2_D_REG_1__SCAN_IN), .S(n9073), .Z(P2_U3377)
         );
  NAND3_X1 U10595 ( .A1(n9076), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n9079) );
  OAI22_X1 U10596 ( .A1(n9075), .A2(n9079), .B1(n9078), .B2(n9077), .ZN(n9080)
         );
  AOI21_X1 U10597 ( .B1(n10044), .B2(n9081), .A(n9080), .ZN(n9082) );
  INV_X1 U10598 ( .A(n9082), .ZN(P2_U3264) );
  AOI21_X1 U10599 ( .B1(n9088), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n9083), .ZN(
        n9084) );
  OAI21_X1 U10600 ( .B1(n9085), .B2(n9090), .A(n9084), .ZN(P2_U3267) );
  INV_X1 U10601 ( .A(n9086), .ZN(n10057) );
  AOI21_X1 U10602 ( .B1(n9088), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n9087), .ZN(
        n9089) );
  OAI21_X1 U10603 ( .B1(n10057), .B2(n9090), .A(n9089), .ZN(P2_U3268) );
  INV_X1 U10604 ( .A(n9091), .ZN(n9092) );
  MUX2_X1 U10605 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9092), .S(P2_U3151), .Z(
        P2_U3295) );
  XOR2_X1 U10606 ( .A(n9155), .B(n9157), .Z(n9094) );
  NOR2_X1 U10607 ( .A1(n9094), .A2(n9093), .ZN(n9156) );
  AOI21_X1 U10608 ( .B1(n9094), .B2(n9093), .A(n9156), .ZN(n9099) );
  AOI22_X1 U10609 ( .A1(n9247), .A2(n9551), .B1(n9267), .B2(n9891), .ZN(n9096)
         );
  OAI211_X1 U10610 ( .C1(n9897), .C2(n9250), .A(n9096), .B(n9095), .ZN(n9097)
         );
  AOI21_X1 U10611 ( .B1(n10003), .B2(n9236), .A(n9097), .ZN(n9098) );
  OAI21_X1 U10612 ( .B1(n9099), .B2(n9262), .A(n9098), .ZN(P1_U3215) );
  XOR2_X1 U10613 ( .A(n9101), .B(n9100), .Z(n9106) );
  AOI22_X1 U10614 ( .A1(n9549), .A2(n9284), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9103) );
  NAND2_X1 U10615 ( .A1(n9805), .A2(n9247), .ZN(n9102) );
  OAI211_X1 U10616 ( .C1(n9282), .C2(n9777), .A(n9103), .B(n9102), .ZN(n9104)
         );
  AOI21_X1 U10617 ( .B1(n9957), .B2(n9236), .A(n9104), .ZN(n9105) );
  OAI21_X1 U10618 ( .B1(n9106), .B2(n9262), .A(n9105), .ZN(P1_U3216) );
  XNOR2_X1 U10619 ( .A(n9240), .B(n9241), .ZN(n9108) );
  NOR2_X1 U10620 ( .A1(n9108), .A2(n9107), .ZN(n9239) );
  AOI21_X1 U10621 ( .B1(n9108), .B2(n9107), .A(n9239), .ZN(n9115) );
  AOI22_X1 U10622 ( .A1(n9247), .A2(n9554), .B1(n9267), .B2(n9109), .ZN(n9111)
         );
  OAI211_X1 U10623 ( .C1(n9325), .C2(n9250), .A(n9111), .B(n9110), .ZN(n9112)
         );
  AOI21_X1 U10624 ( .B1(n9113), .B2(n9223), .A(n9112), .ZN(n9114) );
  OAI21_X1 U10625 ( .B1(n9115), .B2(n9262), .A(n9114), .ZN(P1_U3217) );
  INV_X1 U10626 ( .A(n9975), .ZN(n9334) );
  NAND2_X1 U10627 ( .A1(n5217), .A2(n9118), .ZN(n9119) );
  OAI21_X1 U10628 ( .B1(n5217), .B2(n9118), .A(n9119), .ZN(n9256) );
  NOR2_X1 U10629 ( .A1(n9256), .A2(n9257), .ZN(n9255) );
  INV_X1 U10630 ( .A(n9119), .ZN(n9120) );
  NOR3_X1 U10631 ( .A1(n9255), .A2(n9121), .A3(n9120), .ZN(n9122) );
  OAI21_X1 U10632 ( .B1(n9122), .B2(n4501), .A(n9276), .ZN(n9128) );
  INV_X1 U10633 ( .A(n9123), .ZN(n9126) );
  OAI22_X1 U10634 ( .A1(n9124), .A2(n9250), .B1(n9282), .B2(n9841), .ZN(n9125)
         );
  AOI211_X1 U10635 ( .C1(n9247), .C2(n9835), .A(n9126), .B(n9125), .ZN(n9127)
         );
  OAI211_X1 U10636 ( .C1(n9334), .C2(n9287), .A(n9128), .B(n9127), .ZN(
        P1_U3219) );
  INV_X1 U10637 ( .A(n9130), .ZN(n9131) );
  AOI21_X1 U10638 ( .B1(n9133), .B2(n9132), .A(n9131), .ZN(n9138) );
  NAND2_X1 U10639 ( .A1(n9805), .A2(n9284), .ZN(n9135) );
  AOI22_X1 U10640 ( .A1(n9836), .A2(n9247), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9134) );
  OAI211_X1 U10641 ( .C1(n9282), .C2(n9811), .A(n9135), .B(n9134), .ZN(n9136)
         );
  AOI21_X1 U10642 ( .B1(n9966), .B2(n9236), .A(n9136), .ZN(n9137) );
  OAI21_X1 U10643 ( .B1(n9138), .B2(n9262), .A(n9137), .ZN(P1_U3223) );
  XOR2_X1 U10644 ( .A(n9140), .B(n9141), .Z(n9147) );
  AOI22_X1 U10645 ( .A1(n9247), .A2(n9552), .B1(n9267), .B2(n9142), .ZN(n9143)
         );
  NAND2_X1 U10646 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10095)
         );
  OAI211_X1 U10647 ( .C1(n9899), .C2(n9250), .A(n9143), .B(n10095), .ZN(n9144)
         );
  AOI21_X1 U10648 ( .B1(n9145), .B2(n9223), .A(n9144), .ZN(n9146) );
  OAI21_X1 U10649 ( .B1(n9147), .B2(n9262), .A(n9146), .ZN(P1_U3224) );
  XOR2_X1 U10650 ( .A(n9149), .B(n9148), .Z(n9154) );
  AOI22_X1 U10651 ( .A1(n9549), .A2(n9247), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9151) );
  NAND2_X1 U10652 ( .A1(n9742), .A2(n9267), .ZN(n9150) );
  OAI211_X1 U10653 ( .C1(n9736), .C2(n9250), .A(n9151), .B(n9150), .ZN(n9152)
         );
  AOI21_X1 U10654 ( .B1(n9741), .B2(n9223), .A(n9152), .ZN(n9153) );
  OAI21_X1 U10655 ( .B1(n9154), .B2(n9262), .A(n9153), .ZN(P1_U3225) );
  INV_X1 U10656 ( .A(n9155), .ZN(n9158) );
  AOI21_X1 U10657 ( .B1(n9158), .B2(n9157), .A(n9156), .ZN(n9161) );
  XNOR2_X1 U10658 ( .A(n9161), .B(n9159), .ZN(n9274) );
  NAND2_X1 U10659 ( .A1(n9274), .A2(n9275), .ZN(n9273) );
  OAI21_X1 U10660 ( .B1(n9161), .B2(n9160), .A(n9273), .ZN(n9165) );
  XNOR2_X1 U10661 ( .A(n9163), .B(n9162), .ZN(n9164) );
  XNOR2_X1 U10662 ( .A(n9165), .B(n9164), .ZN(n9169) );
  AOI22_X1 U10663 ( .A1(n9247), .A2(n9868), .B1(n9267), .B2(n9873), .ZN(n9166)
         );
  NAND2_X1 U10664 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9634) );
  OAI211_X1 U10665 ( .C1(n9855), .C2(n9250), .A(n9166), .B(n9634), .ZN(n9167)
         );
  AOI21_X1 U10666 ( .B1(n5807), .B2(n9223), .A(n9167), .ZN(n9168) );
  OAI21_X1 U10667 ( .B1(n9169), .B2(n9262), .A(n9168), .ZN(P1_U3226) );
  XNOR2_X1 U10668 ( .A(n9171), .B(n9170), .ZN(n9172) );
  XNOR2_X1 U10669 ( .A(n9173), .B(n9172), .ZN(n9185) );
  INV_X1 U10670 ( .A(n9174), .ZN(n9176) );
  INV_X1 U10671 ( .A(n9179), .ZN(n9175) );
  OAI21_X1 U10672 ( .B1(n9176), .B2(n9175), .A(P1_STATE_REG_SCAN_IN), .ZN(
        n9182) );
  OAI22_X1 U10673 ( .A1(n9178), .A2(n9250), .B1(n9279), .B2(n9177), .ZN(n9181)
         );
  NOR3_X1 U10674 ( .A1(n9282), .A2(P1_REG3_REG_17__SCAN_IN), .A3(n9179), .ZN(
        n9180) );
  AOI211_X1 U10675 ( .C1(P1_REG3_REG_17__SCAN_IN), .C2(n9182), .A(n9181), .B(
        n9180), .ZN(n9184) );
  NAND2_X1 U10676 ( .A1(n9988), .A2(n9236), .ZN(n9183) );
  OAI211_X1 U10677 ( .C1(n9185), .C2(n9262), .A(n9184), .B(n9183), .ZN(
        P1_U3228) );
  XOR2_X1 U10678 ( .A(n9188), .B(n9187), .Z(n9193) );
  AOI22_X1 U10679 ( .A1(n9796), .A2(n9247), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9190) );
  NAND2_X1 U10680 ( .A1(n9758), .A2(n9267), .ZN(n9189) );
  OAI211_X1 U10681 ( .C1(n9717), .C2(n9250), .A(n9190), .B(n9189), .ZN(n9191)
         );
  AOI21_X1 U10682 ( .B1(n9950), .B2(n9223), .A(n9191), .ZN(n9192) );
  OAI21_X1 U10683 ( .B1(n9193), .B2(n9262), .A(n9192), .ZN(P1_U3229) );
  AOI21_X1 U10684 ( .B1(n9195), .B2(n7978), .A(n9194), .ZN(n9199) );
  XNOR2_X1 U10685 ( .A(n9197), .B(n9196), .ZN(n9198) );
  XNOR2_X1 U10686 ( .A(n9199), .B(n9198), .ZN(n9206) );
  AOI22_X1 U10687 ( .A1(n9284), .A2(n9553), .B1(n9267), .B2(n9200), .ZN(n9201)
         );
  NAND2_X1 U10688 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n10077) );
  OAI211_X1 U10689 ( .C1(n9202), .C2(n9279), .A(n9201), .B(n10077), .ZN(n9203)
         );
  AOI21_X1 U10690 ( .B1(n4572), .B2(n9223), .A(n9203), .ZN(n9205) );
  OAI21_X1 U10691 ( .B1(n9206), .B2(n9262), .A(n9205), .ZN(P1_U3231) );
  INV_X1 U10692 ( .A(n9207), .ZN(n9209) );
  NOR2_X1 U10693 ( .A1(n9209), .A2(n9208), .ZN(n9210) );
  XNOR2_X1 U10694 ( .A(n9211), .B(n9210), .ZN(n9216) );
  AOI22_X1 U10695 ( .A1(n9247), .A2(n9820), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9214) );
  INV_X1 U10696 ( .A(n9212), .ZN(n9827) );
  AOI22_X1 U10697 ( .A1(n9821), .A2(n9284), .B1(n9827), .B2(n9267), .ZN(n9213)
         );
  OAI211_X1 U10698 ( .C1(n6102), .C2(n9287), .A(n9214), .B(n9213), .ZN(n9215)
         );
  AOI21_X1 U10699 ( .B1(n9216), .B2(n9276), .A(n9215), .ZN(n9217) );
  INV_X1 U10700 ( .A(n9217), .ZN(P1_U3233) );
  XOR2_X1 U10701 ( .A(n9219), .B(n9218), .Z(n9225) );
  AOI22_X1 U10702 ( .A1(n9247), .A2(n9916), .B1(n9267), .B2(n9921), .ZN(n9221)
         );
  OAI211_X1 U10703 ( .C1(n9280), .C2(n9250), .A(n9221), .B(n9220), .ZN(n9222)
         );
  AOI21_X1 U10704 ( .B1(n10008), .B2(n9223), .A(n9222), .ZN(n9224) );
  OAI21_X1 U10705 ( .B1(n9225), .B2(n9262), .A(n9224), .ZN(P1_U3234) );
  NAND2_X1 U10706 ( .A1(n9227), .A2(n9226), .ZN(n9229) );
  XNOR2_X1 U10707 ( .A(n9229), .B(n9228), .ZN(n9238) );
  OAI22_X1 U10708 ( .A1(n9231), .A2(n9250), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9230), .ZN(n9235) );
  INV_X1 U10709 ( .A(n9787), .ZN(n9232) );
  OAI22_X1 U10710 ( .A1(n9233), .A2(n9279), .B1(n9232), .B2(n9282), .ZN(n9234)
         );
  AOI211_X1 U10711 ( .C1(n9960), .C2(n9236), .A(n9235), .B(n9234), .ZN(n9237)
         );
  OAI21_X1 U10712 ( .B1(n9238), .B2(n9262), .A(n9237), .ZN(P1_U3235) );
  AOI21_X1 U10713 ( .B1(n9241), .B2(n9240), .A(n9239), .ZN(n9245) );
  XNOR2_X1 U10714 ( .A(n9243), .B(n9242), .ZN(n9244) );
  XNOR2_X1 U10715 ( .A(n9245), .B(n9244), .ZN(n9254) );
  AOI22_X1 U10716 ( .A1(n9247), .A2(n9553), .B1(n9267), .B2(n9246), .ZN(n9249)
         );
  OAI211_X1 U10717 ( .C1(n9251), .C2(n9250), .A(n9249), .B(n9248), .ZN(n9252)
         );
  AOI21_X1 U10718 ( .B1(n9326), .B2(n9223), .A(n9252), .ZN(n9253) );
  OAI21_X1 U10719 ( .B1(n9254), .B2(n9262), .A(n9253), .ZN(P1_U3236) );
  AOI21_X1 U10720 ( .B1(n9257), .B2(n9256), .A(n9255), .ZN(n9261) );
  AOI22_X1 U10721 ( .A1(n9284), .A2(n9820), .B1(n9267), .B2(n9857), .ZN(n9258)
         );
  NAND2_X1 U10722 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9665) );
  OAI211_X1 U10723 ( .C1(n9855), .C2(n9279), .A(n9258), .B(n9665), .ZN(n9259)
         );
  AOI21_X1 U10724 ( .B1(n9983), .B2(n9236), .A(n9259), .ZN(n9260) );
  OAI21_X1 U10725 ( .B1(n9261), .B2(n9262), .A(n9260), .ZN(P1_U3238) );
  AOI21_X1 U10726 ( .B1(n9264), .B2(n9263), .A(n9262), .ZN(n9266) );
  NAND2_X1 U10727 ( .A1(n9266), .A2(n9265), .ZN(n9272) );
  INV_X1 U10728 ( .A(n9725), .ZN(n9268) );
  AOI22_X1 U10729 ( .A1(n9268), .A2(n9267), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9269) );
  OAI21_X1 U10730 ( .B1(n9717), .B2(n9279), .A(n9269), .ZN(n9270) );
  AOI21_X1 U10731 ( .B1(n9547), .B2(n9284), .A(n9270), .ZN(n9271) );
  OAI211_X1 U10732 ( .C1(n10022), .C2(n9287), .A(n9272), .B(n9271), .ZN(
        P1_U3240) );
  OAI21_X1 U10733 ( .B1(n9275), .B2(n9274), .A(n9273), .ZN(n9277) );
  NAND2_X1 U10734 ( .A1(n9277), .A2(n9276), .ZN(n9286) );
  AND2_X1 U10735 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9625) );
  INV_X1 U10736 ( .A(n9278), .ZN(n9281) );
  OAI22_X1 U10737 ( .A1(n9282), .A2(n9281), .B1(n9280), .B2(n9279), .ZN(n9283)
         );
  AOI211_X1 U10738 ( .C1(n9284), .C2(n9550), .A(n9625), .B(n9283), .ZN(n9285)
         );
  OAI211_X1 U10739 ( .C1(n9288), .C2(n9287), .A(n9286), .B(n9285), .ZN(
        P1_U3241) );
  INV_X1 U10740 ( .A(n9524), .ZN(n9436) );
  AND4_X1 U10741 ( .A1(n9501), .A2(n9394), .A3(n9385), .A4(n9497), .ZN(n9391)
         );
  INV_X1 U10742 ( .A(n9289), .ZN(n9290) );
  NAND2_X1 U10743 ( .A1(n9335), .A2(n9353), .ZN(n9483) );
  INV_X1 U10744 ( .A(n4573), .ZN(n9295) );
  AND4_X1 U10745 ( .A1(n9291), .A2(n9292), .A3(n9293), .A4(n9381), .ZN(n9294)
         );
  OAI21_X1 U10746 ( .B1(n9296), .B2(n9295), .A(n9294), .ZN(n9313) );
  NOR2_X1 U10747 ( .A1(n9558), .A2(n9381), .ZN(n9303) );
  NAND2_X1 U10748 ( .A1(n9303), .A2(n9302), .ZN(n9297) );
  NAND2_X1 U10749 ( .A1(n9297), .A2(n10139), .ZN(n9301) );
  AND2_X1 U10750 ( .A1(n9558), .A2(n9381), .ZN(n9305) );
  INV_X1 U10751 ( .A(n9305), .ZN(n9298) );
  OAI21_X1 U10752 ( .B1(n9298), .B2(n9302), .A(n9304), .ZN(n9300) );
  AOI21_X1 U10753 ( .B1(n9301), .B2(n9300), .A(n9299), .ZN(n9312) );
  AOI22_X1 U10754 ( .A1(n9303), .A2(n10139), .B1(n9394), .B2(n9302), .ZN(n9307) );
  AOI22_X1 U10755 ( .A1(n9557), .A2(n9381), .B1(n9305), .B2(n9304), .ZN(n9306)
         );
  MUX2_X1 U10756 ( .A(n9307), .B(n9306), .S(n10103), .Z(n9311) );
  NAND4_X1 U10757 ( .A1(n4573), .A2(n9415), .A3(n9449), .A4(n9394), .ZN(n9308)
         );
  OR2_X1 U10758 ( .A1(n9309), .A2(n9308), .ZN(n9310) );
  NAND2_X1 U10759 ( .A1(n9314), .A2(n9408), .ZN(n9315) );
  MUX2_X1 U10760 ( .A(n9316), .B(n9315), .S(n9394), .Z(n9317) );
  INV_X1 U10761 ( .A(n9317), .ZN(n9318) );
  AND2_X1 U10762 ( .A1(n9323), .A2(n9319), .ZN(n9320) );
  MUX2_X1 U10763 ( .A(n9321), .B(n9320), .S(n9394), .Z(n9322) );
  NAND2_X1 U10764 ( .A1(n9343), .A2(n9323), .ZN(n9324) );
  NAND2_X1 U10765 ( .A1(n9348), .A2(n9344), .ZN(n9461) );
  AOI21_X1 U10766 ( .B1(n9324), .B2(n9458), .A(n9461), .ZN(n9327) );
  OR2_X1 U10767 ( .A1(n9326), .A2(n9325), .ZN(n9346) );
  NAND2_X1 U10768 ( .A1(n9349), .A2(n9346), .ZN(n9462) );
  OAI21_X1 U10769 ( .B1(n9327), .B2(n9462), .A(n9465), .ZN(n9328) );
  NAND2_X1 U10770 ( .A1(n9328), .A2(n9468), .ZN(n9329) );
  INV_X1 U10771 ( .A(n9895), .ZN(n9888) );
  NAND3_X1 U10772 ( .A1(n9329), .A2(n9888), .A3(n9466), .ZN(n9330) );
  NAND3_X1 U10773 ( .A1(n9330), .A2(n9471), .A3(n9467), .ZN(n9332) );
  INV_X1 U10774 ( .A(n9476), .ZN(n9331) );
  AOI21_X1 U10775 ( .B1(n9332), .B2(n9351), .A(n9331), .ZN(n9333) );
  AOI21_X1 U10776 ( .B1(n9406), .B2(n9334), .A(n9394), .ZN(n9338) );
  NAND2_X1 U10777 ( .A1(n9802), .A2(n9335), .ZN(n9337) );
  NAND3_X1 U10778 ( .A1(n9406), .A2(n9381), .A3(n9820), .ZN(n9336) );
  OAI21_X1 U10779 ( .B1(n9338), .B2(n9337), .A(n9336), .ZN(n9361) );
  NAND2_X1 U10780 ( .A1(n9483), .A2(n9381), .ZN(n9359) );
  INV_X1 U10781 ( .A(n9479), .ZN(n9340) );
  NOR2_X1 U10782 ( .A1(n9480), .A2(n9381), .ZN(n9339) );
  AOI22_X1 U10783 ( .A1(n9340), .A2(n9394), .B1(n9353), .B2(n9339), .ZN(n9341)
         );
  AND2_X1 U10784 ( .A1(n9341), .A2(n9487), .ZN(n9358) );
  NAND2_X1 U10785 ( .A1(n9345), .A2(n9344), .ZN(n9347) );
  AND2_X1 U10786 ( .A1(n9351), .A2(n9350), .ZN(n9473) );
  AOI21_X1 U10787 ( .B1(n9352), .B2(n9471), .A(n9475), .ZN(n9355) );
  NAND4_X1 U10788 ( .A1(n9353), .A2(n9394), .A3(n9476), .A4(n9478), .ZN(n9354)
         );
  OR2_X1 U10789 ( .A1(n9355), .A2(n9354), .ZN(n9357) );
  NAND3_X1 U10790 ( .A1(n9479), .A2(n9381), .A3(n9480), .ZN(n9356) );
  NAND4_X1 U10791 ( .A1(n9359), .A2(n9358), .A3(n9357), .A4(n9356), .ZN(n9360)
         );
  NAND2_X1 U10792 ( .A1(n9363), .A2(n9362), .ZN(n9365) );
  MUX2_X1 U10793 ( .A(n9404), .B(n9405), .S(n9394), .Z(n9364) );
  NAND2_X1 U10794 ( .A1(n9365), .A2(n9364), .ZN(n9366) );
  INV_X1 U10795 ( .A(n9791), .ZN(n9782) );
  NAND2_X1 U10796 ( .A1(n9366), .A2(n9782), .ZN(n9371) );
  AND2_X1 U10797 ( .A1(n9748), .A2(n9367), .ZN(n9489) );
  INV_X1 U10798 ( .A(n9369), .ZN(n9368) );
  AOI21_X1 U10799 ( .B1(n9371), .B2(n9489), .A(n9368), .ZN(n9373) );
  AND2_X1 U10800 ( .A1(n9369), .A2(n9764), .ZN(n9441) );
  AOI21_X1 U10801 ( .B1(n9371), .B2(n9441), .A(n9370), .ZN(n9372) );
  MUX2_X1 U10802 ( .A(n9373), .B(n9372), .S(n9394), .Z(n9376) );
  MUX2_X1 U10803 ( .A(n9444), .B(n9491), .S(n9381), .Z(n9374) );
  INV_X1 U10804 ( .A(n9374), .ZN(n9375) );
  INV_X1 U10805 ( .A(n9386), .ZN(n9378) );
  INV_X1 U10806 ( .A(n9384), .ZN(n9377) );
  OAI211_X1 U10807 ( .C1(n9378), .C2(n9377), .A(n9492), .B(n9700), .ZN(n9390)
         );
  INV_X1 U10808 ( .A(n9388), .ZN(n9499) );
  INV_X1 U10809 ( .A(n9497), .ZN(n9516) );
  NAND3_X1 U10810 ( .A1(n9499), .A2(n9516), .A3(n9381), .ZN(n9383) );
  NAND3_X1 U10811 ( .A1(n9388), .A2(n9394), .A3(n9501), .ZN(n9382) );
  NAND2_X1 U10812 ( .A1(n9385), .A2(n9384), .ZN(n9488) );
  MUX2_X1 U10813 ( .A(n9502), .B(n9504), .S(n9394), .Z(n9392) );
  INV_X1 U10814 ( .A(n9395), .ZN(n9393) );
  AOI21_X1 U10815 ( .B1(n9543), .B2(n9544), .A(n9524), .ZN(n9396) );
  OAI21_X1 U10816 ( .B1(n4544), .B2(n9920), .A(n9398), .ZN(n9401) );
  NOR3_X1 U10817 ( .A1(n9538), .A2(n6068), .A3(n9399), .ZN(n9400) );
  OAI211_X1 U10818 ( .C1(n9436), .C2(n9920), .A(n9401), .B(n9400), .ZN(n9542)
         );
  INV_X1 U10819 ( .A(n9538), .ZN(n9438) );
  AOI21_X1 U10820 ( .B1(n10014), .B2(n9544), .A(n9514), .ZN(n9512) );
  INV_X1 U10821 ( .A(n9403), .ZN(n9434) );
  INV_X1 U10822 ( .A(n9721), .ZN(n9432) );
  NAND2_X1 U10823 ( .A1(n9405), .A2(n9404), .ZN(n9807) );
  NAND2_X1 U10824 ( .A1(n9802), .A2(n9406), .ZN(n9823) );
  INV_X1 U10825 ( .A(n9834), .ZN(n9838) );
  INV_X1 U10826 ( .A(n9408), .ZN(n9409) );
  NOR4_X1 U10827 ( .A1(n9411), .A2(n9410), .A3(n9409), .A4(n9447), .ZN(n9418)
         );
  NOR3_X1 U10828 ( .A1(n9414), .A2(n9413), .A3(n9412), .ZN(n9417) );
  NAND4_X1 U10829 ( .A1(n9418), .A2(n9417), .A3(n9416), .A4(n9415), .ZN(n9421)
         );
  NOR3_X1 U10830 ( .A1(n9421), .A2(n9420), .A3(n9419), .ZN(n9423) );
  NAND4_X1 U10831 ( .A1(n4621), .A2(n9424), .A3(n9423), .A4(n9422), .ZN(n9425)
         );
  NOR4_X1 U10832 ( .A1(n9426), .A2(n9425), .A3(n9895), .A4(n9925), .ZN(n9427)
         );
  NAND3_X1 U10833 ( .A1(n9883), .A2(n9428), .A3(n9427), .ZN(n9429) );
  OR4_X1 U10834 ( .A1(n9823), .A2(n9838), .A3(n9860), .A4(n9429), .ZN(n9430)
         );
  NOR4_X1 U10835 ( .A1(n9768), .A2(n9791), .A3(n9807), .A4(n9430), .ZN(n9431)
         );
  NAND4_X1 U10836 ( .A1(n9432), .A2(n9754), .A3(n9733), .A4(n9431), .ZN(n9433)
         );
  NOR4_X1 U10837 ( .A1(n9689), .A2(n9434), .A3(n9698), .A4(n9433), .ZN(n9437)
         );
  NAND2_X1 U10838 ( .A1(n9683), .A2(n9435), .ZN(n9503) );
  NAND4_X1 U10839 ( .A1(n9512), .A2(n9437), .A3(n9436), .A4(n9503), .ZN(n9528)
         );
  NAND4_X1 U10840 ( .A1(n9439), .A2(n9527), .A3(n9438), .A4(n9528), .ZN(n9541)
         );
  INV_X1 U10841 ( .A(n9440), .ZN(n9445) );
  INV_X1 U10842 ( .A(n9441), .ZN(n9442) );
  NAND2_X1 U10843 ( .A1(n9442), .A2(n9748), .ZN(n9443) );
  NAND2_X1 U10844 ( .A1(n9444), .A2(n9443), .ZN(n9494) );
  NOR3_X1 U10845 ( .A1(n9488), .A2(n9445), .A3(n9494), .ZN(n9515) );
  INV_X1 U10846 ( .A(n9446), .ZN(n9456) );
  OAI21_X1 U10847 ( .B1(n9448), .B2(n6601), .A(n9447), .ZN(n9455) );
  NAND3_X1 U10848 ( .A1(n4573), .A2(n9450), .A3(n9449), .ZN(n9454) );
  INV_X1 U10849 ( .A(n9452), .ZN(n9453) );
  NOR4_X1 U10850 ( .A1(n9456), .A2(n9455), .A3(n9454), .A4(n9453), .ZN(n9459)
         );
  OAI211_X1 U10851 ( .C1(n9460), .C2(n9459), .A(n9458), .B(n9457), .ZN(n9464)
         );
  INV_X1 U10852 ( .A(n9461), .ZN(n9463) );
  AOI21_X1 U10853 ( .B1(n9464), .B2(n9463), .A(n9462), .ZN(n9470) );
  NAND2_X1 U10854 ( .A1(n9466), .A2(n9465), .ZN(n9469) );
  OAI211_X1 U10855 ( .C1(n9470), .C2(n9469), .A(n9468), .B(n9467), .ZN(n9474)
         );
  INV_X1 U10856 ( .A(n9471), .ZN(n9472) );
  AOI21_X1 U10857 ( .B1(n9474), .B2(n9473), .A(n9472), .ZN(n9477) );
  AOI21_X1 U10858 ( .B1(n9477), .B2(n9476), .A(n9475), .ZN(n9482) );
  INV_X1 U10859 ( .A(n9478), .ZN(n9481) );
  OAI211_X1 U10860 ( .C1(n9482), .C2(n9481), .A(n9480), .B(n9479), .ZN(n9485)
         );
  INV_X1 U10861 ( .A(n9483), .ZN(n9484) );
  NAND2_X1 U10862 ( .A1(n9485), .A2(n9484), .ZN(n9486) );
  AOI21_X1 U10863 ( .B1(n9487), .B2(n9486), .A(n9516), .ZN(n9500) );
  INV_X1 U10864 ( .A(n9488), .ZN(n9496) );
  INV_X1 U10865 ( .A(n9489), .ZN(n9490) );
  NOR2_X1 U10866 ( .A1(n9490), .A2(n9792), .ZN(n9493) );
  OAI211_X1 U10867 ( .C1(n9494), .C2(n9493), .A(n9492), .B(n9491), .ZN(n9495)
         );
  NAND3_X1 U10868 ( .A1(n9497), .A2(n9496), .A3(n9495), .ZN(n9498) );
  OAI211_X1 U10869 ( .C1(n9516), .C2(n9700), .A(n9499), .B(n9498), .ZN(n9520)
         );
  AOI21_X1 U10870 ( .B1(n9515), .B2(n9500), .A(n9520), .ZN(n9507) );
  NAND2_X1 U10871 ( .A1(n9502), .A2(n9501), .ZN(n9518) );
  INV_X1 U10872 ( .A(n9503), .ZN(n9506) );
  INV_X1 U10873 ( .A(n9504), .ZN(n9505) );
  OAI21_X1 U10874 ( .B1(n9507), .B2(n9518), .A(n9523), .ZN(n9508) );
  AOI21_X1 U10875 ( .B1(n9512), .B2(n9508), .A(n9524), .ZN(n9509) );
  INV_X1 U10876 ( .A(n9509), .ZN(n9533) );
  NOR2_X1 U10877 ( .A1(n9509), .A2(n9920), .ZN(n9510) );
  AOI211_X1 U10878 ( .C1(n9527), .C2(n9511), .A(n9538), .B(n9510), .ZN(n9532)
         );
  INV_X1 U10879 ( .A(n9512), .ZN(n9513) );
  INV_X1 U10880 ( .A(n9515), .ZN(n9517) );
  INV_X1 U10881 ( .A(n9803), .ZN(n9819) );
  NOR3_X1 U10882 ( .A1(n9517), .A2(n9516), .A3(n9819), .ZN(n9521) );
  INV_X1 U10883 ( .A(n9518), .ZN(n9519) );
  OAI21_X1 U10884 ( .B1(n9521), .B2(n9520), .A(n9519), .ZN(n9522) );
  OAI211_X1 U10885 ( .C1(n10014), .C2(n9543), .A(n9523), .B(n9522), .ZN(n9525)
         );
  AOI21_X1 U10886 ( .B1(n9526), .B2(n9525), .A(n9524), .ZN(n9530) );
  OAI211_X1 U10887 ( .C1(n9530), .C2(n9529), .A(n9528), .B(n9527), .ZN(n9531)
         );
  OAI211_X1 U10888 ( .C1(n9534), .C2(n9533), .A(n9532), .B(n9531), .ZN(n9540)
         );
  INV_X1 U10889 ( .A(n10269), .ZN(n9536) );
  NAND4_X1 U10890 ( .A1(n9536), .A2(n9915), .A3(n9535), .A4(n6595), .ZN(n9537)
         );
  OAI211_X1 U10891 ( .C1(n6068), .C2(n9538), .A(n9537), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9539) );
  NAND4_X1 U10892 ( .A1(n9540), .A2(n9541), .A3(n9542), .A4(n9539), .ZN(
        P1_U3242) );
  MUX2_X1 U10893 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9543), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10894 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9544), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10895 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9545), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10896 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9546), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10897 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9547), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10898 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9548), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10899 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9750), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10900 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9549), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10901 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9796), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10902 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9805), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10903 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9821), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10904 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9836), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10905 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9820), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10906 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9835), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10907 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9867), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10908 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9550), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10909 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9868), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10910 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9914), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10911 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9551), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10912 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9916), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10913 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9552), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10914 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9553), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10915 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9554), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10916 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9555), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10917 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9556), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10918 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9557), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10919 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9558), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10920 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9559), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10921 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9560), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10922 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9561), .S(P1_U3973), .Z(
        P1_U3556) );
  OAI22_X1 U10923 ( .A1(n10098), .A2(n9562), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10283), .ZN(n9563) );
  AOI21_X1 U10924 ( .B1(n9564), .B2(n9650), .A(n9563), .ZN(n9573) );
  OAI211_X1 U10925 ( .C1(n9567), .C2(n9566), .A(n9663), .B(n9565), .ZN(n9572)
         );
  OAI211_X1 U10926 ( .C1(n9570), .C2(n9569), .A(n10093), .B(n9568), .ZN(n9571)
         );
  NAND3_X1 U10927 ( .A1(n9573), .A2(n9572), .A3(n9571), .ZN(P1_U3244) );
  MUX2_X1 U10928 ( .A(n9575), .B(n9574), .S(n6158), .Z(n9579) );
  NAND2_X1 U10929 ( .A1(n9576), .A2(n5071), .ZN(n9577) );
  OAI211_X1 U10930 ( .C1(n9579), .C2(n4437), .A(P1_U3973), .B(n9577), .ZN(
        n9620) );
  INV_X1 U10931 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9582) );
  OAI22_X1 U10932 ( .A1(n10098), .A2(n9582), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9581), .ZN(n9583) );
  AOI21_X1 U10933 ( .B1(n4698), .B2(n9650), .A(n9583), .ZN(n9591) );
  OAI211_X1 U10934 ( .C1(n9585), .C2(n9584), .A(n9663), .B(n9599), .ZN(n9590)
         );
  OAI211_X1 U10935 ( .C1(n9588), .C2(n9587), .A(n10093), .B(n9586), .ZN(n9589)
         );
  NAND4_X1 U10936 ( .A1(n9620), .A2(n9591), .A3(n9590), .A4(n9589), .ZN(
        P1_U3245) );
  OAI211_X1 U10937 ( .C1(n9594), .C2(n9593), .A(n10093), .B(n9592), .ZN(n9604)
         );
  AOI21_X1 U10938 ( .B1(n9671), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n9595), .ZN(
        n9603) );
  NAND2_X1 U10939 ( .A1(n9650), .A2(n9596), .ZN(n9602) );
  MUX2_X1 U10940 ( .A(n7041), .B(P1_REG1_REG_3__SCAN_IN), .S(n9596), .Z(n9597)
         );
  NAND3_X1 U10941 ( .A1(n9599), .A2(n9598), .A3(n9597), .ZN(n9600) );
  NAND3_X1 U10942 ( .A1(n9663), .A2(n9611), .A3(n9600), .ZN(n9601) );
  NAND4_X1 U10943 ( .A1(n9604), .A2(n9603), .A3(n9602), .A4(n9601), .ZN(
        P1_U3246) );
  AOI21_X1 U10944 ( .B1(n9671), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n9605), .ZN(
        n9619) );
  OAI211_X1 U10945 ( .C1(n9607), .C2(n9606), .A(n10093), .B(n4841), .ZN(n9615)
         );
  MUX2_X1 U10946 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n7044), .S(n9608), .Z(n9609)
         );
  NAND3_X1 U10947 ( .A1(n9611), .A2(n9610), .A3(n9609), .ZN(n9612) );
  NAND3_X1 U10948 ( .A1(n9663), .A2(n9613), .A3(n9612), .ZN(n9614) );
  AND2_X1 U10949 ( .A1(n9615), .A2(n9614), .ZN(n9618) );
  NAND2_X1 U10950 ( .A1(n9650), .A2(n9616), .ZN(n9617) );
  NAND4_X1 U10951 ( .A1(n9620), .A2(n9619), .A3(n9618), .A4(n9617), .ZN(
        P1_U3247) );
  AOI211_X1 U10952 ( .C1(n10368), .C2(n9622), .A(n9621), .B(n10067), .ZN(n9630) );
  OAI211_X1 U10953 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9624), .A(n9663), .B(
        n9623), .ZN(n9627) );
  AOI21_X1 U10954 ( .B1(n9671), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n9625), .ZN(
        n9626) );
  OAI211_X1 U10955 ( .C1(n10088), .C2(n9628), .A(n9627), .B(n9626), .ZN(n9629)
         );
  OR2_X1 U10956 ( .A1(n9630), .A2(n9629), .ZN(P1_U3258) );
  AOI21_X1 U10957 ( .B1(n9633), .B2(n9632), .A(n9631), .ZN(n9644) );
  INV_X1 U10958 ( .A(n9634), .ZN(n9640) );
  INV_X1 U10959 ( .A(n9635), .ZN(n9636) );
  AOI211_X1 U10960 ( .C1(n9638), .C2(n9637), .A(n9636), .B(n10067), .ZN(n9639)
         );
  AOI211_X1 U10961 ( .C1(n9671), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9640), .B(
        n9639), .ZN(n9643) );
  NAND2_X1 U10962 ( .A1(n9650), .A2(n9641), .ZN(n9642) );
  OAI211_X1 U10963 ( .C1(n9644), .C2(n10090), .A(n9643), .B(n9642), .ZN(
        P1_U3259) );
  AOI21_X1 U10964 ( .B1(n9646), .B2(n9645), .A(n9661), .ZN(n9657) );
  INV_X1 U10965 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9648) );
  OAI22_X1 U10966 ( .A1(n10098), .A2(n9648), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9647), .ZN(n9649) );
  AOI21_X1 U10967 ( .B1(n9651), .B2(n9650), .A(n9649), .ZN(n9656) );
  OAI21_X1 U10968 ( .B1(n9653), .B2(n4520), .A(n9652), .ZN(n9654) );
  NAND2_X1 U10969 ( .A1(n9654), .A2(n10093), .ZN(n9655) );
  OAI211_X1 U10970 ( .C1(n9657), .C2(n10090), .A(n9656), .B(n9655), .ZN(
        P1_U3260) );
  INV_X1 U10971 ( .A(n9658), .ZN(n9664) );
  OAI21_X1 U10972 ( .B1(n9661), .B2(n9660), .A(n9659), .ZN(n9662) );
  NAND3_X1 U10973 ( .A1(n9664), .A2(n9663), .A3(n9662), .ZN(n9673) );
  INV_X1 U10974 ( .A(n9665), .ZN(n9670) );
  AOI211_X1 U10975 ( .C1(n9668), .C2(n9667), .A(n9666), .B(n10067), .ZN(n9669)
         );
  AOI211_X1 U10976 ( .C1(n9671), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9670), .B(
        n9669), .ZN(n9672) );
  OAI211_X1 U10977 ( .C1(n10088), .C2(n9674), .A(n9673), .B(n9672), .ZN(
        P1_U3261) );
  NAND2_X1 U10978 ( .A1(n9675), .A2(n10108), .ZN(n9678) );
  INV_X1 U10979 ( .A(n9932), .ZN(n9676) );
  NOR2_X1 U10980 ( .A1(n10112), .A2(n9676), .ZN(n9684) );
  AOI21_X1 U10981 ( .B1(n10112), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9684), .ZN(
        n9677) );
  OAI211_X1 U10982 ( .C1(n9679), .C2(n10115), .A(n9678), .B(n9677), .ZN(
        P1_U3263) );
  INV_X1 U10983 ( .A(n9680), .ZN(n9682) );
  NAND2_X1 U10984 ( .A1(n4471), .A2(n10108), .ZN(n9686) );
  AOI21_X1 U10985 ( .B1(n10112), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9684), .ZN(
        n9685) );
  OAI211_X1 U10986 ( .C1(n10014), .C2(n10115), .A(n9686), .B(n9685), .ZN(
        P1_U3264) );
  NOR2_X1 U10987 ( .A1(n9691), .A2(n10115), .ZN(n9695) );
  OAI22_X1 U10988 ( .A1(n9693), .A2(n9922), .B1(n9692), .B2(n9776), .ZN(n9694)
         );
  AOI211_X1 U10989 ( .C1(n9696), .C2(n10108), .A(n9695), .B(n9694), .ZN(n9697)
         );
  XNOR2_X1 U10990 ( .A(n9699), .B(n9698), .ZN(n9936) );
  NAND2_X1 U10991 ( .A1(n9716), .A2(n9700), .ZN(n9702) );
  XNOR2_X1 U10992 ( .A(n9702), .B(n9701), .ZN(n9705) );
  OAI22_X1 U10993 ( .A1(n9703), .A2(n9896), .B1(n9736), .B2(n9898), .ZN(n9704)
         );
  AOI21_X1 U10994 ( .B1(n9705), .B2(n9918), .A(n9704), .ZN(n9935) );
  INV_X1 U10995 ( .A(n9935), .ZN(n9712) );
  OAI211_X1 U10996 ( .C1(n10018), .C2(n9706), .A(n9707), .B(n9976), .ZN(n9934)
         );
  NOR2_X1 U10997 ( .A1(n9934), .A2(n9876), .ZN(n9711) );
  AOI22_X1 U10998 ( .A1(n9708), .A2(n10110), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10112), .ZN(n9709) );
  OAI21_X1 U10999 ( .B1(n10018), .B2(n10115), .A(n9709), .ZN(n9710) );
  AOI211_X1 U11000 ( .C1(n9712), .C2(n9776), .A(n9711), .B(n9710), .ZN(n9713)
         );
  OAI21_X1 U11001 ( .B1(n9936), .B2(n9926), .A(n9713), .ZN(P1_U3266) );
  NAND2_X1 U11002 ( .A1(n9714), .A2(n9721), .ZN(n9715) );
  OAI22_X1 U11003 ( .A1(n9718), .A2(n9896), .B1(n9717), .B2(n9898), .ZN(n9719)
         );
  INV_X1 U11004 ( .A(n9939), .ZN(n9730) );
  XOR2_X1 U11005 ( .A(n9721), .B(n9720), .Z(n9941) );
  NAND2_X1 U11006 ( .A1(n9941), .A2(n10119), .ZN(n9729) );
  INV_X1 U11007 ( .A(n9740), .ZN(n9722) );
  AOI211_X1 U11008 ( .C1(n9723), .C2(n9722), .A(n9907), .B(n9706), .ZN(n9940)
         );
  NOR2_X1 U11009 ( .A1(n10022), .A2(n10115), .ZN(n9727) );
  OAI22_X1 U11010 ( .A1(n9725), .A2(n9922), .B1(n9724), .B2(n9776), .ZN(n9726)
         );
  AOI211_X1 U11011 ( .C1(n9940), .C2(n10108), .A(n9727), .B(n9726), .ZN(n9728)
         );
  OAI211_X1 U11012 ( .C1(n10112), .C2(n9730), .A(n9729), .B(n9728), .ZN(
        P1_U3267) );
  XNOR2_X1 U11013 ( .A(n9731), .B(n9733), .ZN(n9945) );
  INV_X1 U11014 ( .A(n9945), .ZN(n9747) );
  INV_X1 U11015 ( .A(n9733), .ZN(n9734) );
  XNOR2_X1 U11016 ( .A(n9732), .B(n9734), .ZN(n9735) );
  NAND2_X1 U11017 ( .A1(n9735), .A2(n9918), .ZN(n9739) );
  OAI22_X1 U11018 ( .A1(n9736), .A2(n9896), .B1(n9771), .B2(n9898), .ZN(n9737)
         );
  INV_X1 U11019 ( .A(n9737), .ZN(n9738) );
  NAND2_X1 U11020 ( .A1(n9739), .A2(n9738), .ZN(n9943) );
  INV_X1 U11021 ( .A(n9741), .ZN(n10027) );
  AOI211_X1 U11022 ( .C1(n9741), .C2(n9756), .A(n9907), .B(n9740), .ZN(n9944)
         );
  NAND2_X1 U11023 ( .A1(n9944), .A2(n10108), .ZN(n9744) );
  AOI22_X1 U11024 ( .A1(n9742), .A2(n10110), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10112), .ZN(n9743) );
  OAI211_X1 U11025 ( .C1(n10027), .C2(n10115), .A(n9744), .B(n9743), .ZN(n9745) );
  AOI21_X1 U11026 ( .B1(n9776), .B2(n9943), .A(n9745), .ZN(n9746) );
  OAI21_X1 U11027 ( .B1(n9747), .B2(n9926), .A(n9746), .ZN(P1_U3268) );
  NAND2_X1 U11028 ( .A1(n9765), .A2(n9748), .ZN(n9749) );
  XNOR2_X1 U11029 ( .A(n9749), .B(n9754), .ZN(n9751) );
  AOI222_X1 U11030 ( .A1(n9918), .A2(n9751), .B1(n9750), .B2(n9913), .C1(n9796), .C2(n9915), .ZN(n9953) );
  NAND2_X1 U11031 ( .A1(n9755), .A2(n9754), .ZN(n9949) );
  NAND3_X1 U11032 ( .A1(n9753), .A2(n9949), .A3(n10119), .ZN(n9762) );
  INV_X1 U11033 ( .A(n9756), .ZN(n9757) );
  AOI21_X1 U11034 ( .B1(n9950), .B2(n9772), .A(n9757), .ZN(n9951) );
  AOI22_X1 U11035 ( .A1(n9758), .A2(n10110), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10112), .ZN(n9759) );
  OAI21_X1 U11036 ( .B1(n5002), .B2(n10115), .A(n9759), .ZN(n9760) );
  AOI21_X1 U11037 ( .B1(n9951), .B2(n9844), .A(n9760), .ZN(n9761) );
  OAI211_X1 U11038 ( .C1(n10112), .C2(n9953), .A(n9762), .B(n9761), .ZN(
        P1_U3269) );
  XNOR2_X1 U11039 ( .A(n9763), .B(n9768), .ZN(n9959) );
  NAND2_X1 U11040 ( .A1(n9794), .A2(n9764), .ZN(n9767) );
  INV_X1 U11041 ( .A(n9765), .ZN(n9766) );
  AOI21_X1 U11042 ( .B1(n9768), .B2(n9767), .A(n9766), .ZN(n9769) );
  OAI222_X1 U11043 ( .A1(n9896), .A2(n9771), .B1(n9898), .B2(n9770), .C1(n9893), .C2(n9769), .ZN(n9955) );
  NAND2_X1 U11044 ( .A1(n9955), .A2(n9776), .ZN(n9781) );
  INV_X1 U11045 ( .A(n9772), .ZN(n9773) );
  AOI211_X1 U11046 ( .C1(n9957), .C2(n9784), .A(n9907), .B(n9773), .ZN(n9956)
         );
  INV_X1 U11047 ( .A(n9957), .ZN(n9774) );
  NOR2_X1 U11048 ( .A1(n9774), .A2(n10115), .ZN(n9779) );
  OAI22_X1 U11049 ( .A1(n9777), .A2(n9922), .B1(n9776), .B2(n9775), .ZN(n9778)
         );
  AOI211_X1 U11050 ( .C1(n9956), .C2(n10108), .A(n9779), .B(n9778), .ZN(n9780)
         );
  OAI211_X1 U11051 ( .C1(n9959), .C2(n9926), .A(n9781), .B(n9780), .ZN(
        P1_U3270) );
  XNOR2_X1 U11052 ( .A(n9783), .B(n9782), .ZN(n9964) );
  INV_X1 U11053 ( .A(n9809), .ZN(n9786) );
  INV_X1 U11054 ( .A(n9784), .ZN(n9785) );
  AOI21_X1 U11055 ( .B1(n9960), .B2(n9786), .A(n9785), .ZN(n9961) );
  AOI22_X1 U11056 ( .A1(n9787), .A2(n10110), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10112), .ZN(n9788) );
  OAI21_X1 U11057 ( .B1(n9789), .B2(n10115), .A(n9788), .ZN(n9800) );
  INV_X1 U11058 ( .A(n9790), .ZN(n9793) );
  OAI21_X1 U11059 ( .B1(n9793), .B2(n9792), .A(n9791), .ZN(n9795) );
  NAND3_X1 U11060 ( .A1(n9795), .A2(n9918), .A3(n9794), .ZN(n9798) );
  AOI22_X1 U11061 ( .A1(n9796), .A2(n9913), .B1(n9915), .B2(n9821), .ZN(n9797)
         );
  AND2_X1 U11062 ( .A1(n9798), .A2(n9797), .ZN(n9963) );
  NOR2_X1 U11063 ( .A1(n9963), .A2(n10112), .ZN(n9799) );
  AOI211_X1 U11064 ( .C1(n9844), .C2(n9961), .A(n9800), .B(n9799), .ZN(n9801)
         );
  OAI21_X1 U11065 ( .B1(n9964), .B2(n9926), .A(n9801), .ZN(P1_U3271) );
  OAI21_X1 U11066 ( .B1(n9803), .B2(n9823), .A(n9802), .ZN(n9804) );
  XNOR2_X1 U11067 ( .A(n9804), .B(n9807), .ZN(n9806) );
  AOI222_X1 U11068 ( .A1(n9918), .A2(n9806), .B1(n9805), .B2(n9913), .C1(n9836), .C2(n9915), .ZN(n9968) );
  XNOR2_X1 U11069 ( .A(n9808), .B(n9807), .ZN(n9969) );
  INV_X1 U11070 ( .A(n9969), .ZN(n9817) );
  OAI21_X1 U11071 ( .B1(n5208), .B2(n9815), .A(n9976), .ZN(n9810) );
  NOR2_X1 U11072 ( .A1(n9810), .A2(n9809), .ZN(n9965) );
  NAND2_X1 U11073 ( .A1(n9965), .A2(n10108), .ZN(n9814) );
  INV_X1 U11074 ( .A(n9811), .ZN(n9812) );
  AOI22_X1 U11075 ( .A1(n9812), .A2(n10110), .B1(n10112), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9813) );
  OAI211_X1 U11076 ( .C1(n9815), .C2(n10115), .A(n9814), .B(n9813), .ZN(n9816)
         );
  AOI21_X1 U11077 ( .B1(n9817), .B2(n10119), .A(n9816), .ZN(n9818) );
  OAI21_X1 U11078 ( .B1(n9968), .B2(n10112), .A(n9818), .ZN(P1_U3272) );
  XNOR2_X1 U11079 ( .A(n9819), .B(n9823), .ZN(n9822) );
  AOI222_X1 U11080 ( .A1(n9918), .A2(n9822), .B1(n9821), .B2(n9913), .C1(n9820), .C2(n9915), .ZN(n9973) );
  XOR2_X1 U11081 ( .A(n9824), .B(n9823), .Z(n9974) );
  INV_X1 U11082 ( .A(n9974), .ZN(n9831) );
  NAND2_X1 U11083 ( .A1(n4522), .A2(n9971), .ZN(n9825) );
  NAND2_X1 U11084 ( .A1(n9825), .A2(n9976), .ZN(n9826) );
  NOR2_X1 U11085 ( .A1(n5208), .A2(n9826), .ZN(n9970) );
  NAND2_X1 U11086 ( .A1(n9970), .A2(n10108), .ZN(n9829) );
  AOI22_X1 U11087 ( .A1(n10112), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9827), 
        .B2(n10110), .ZN(n9828) );
  OAI211_X1 U11088 ( .C1(n6102), .C2(n10115), .A(n9829), .B(n9828), .ZN(n9830)
         );
  AOI21_X1 U11089 ( .B1(n9831), .B2(n10119), .A(n9830), .ZN(n9832) );
  OAI21_X1 U11090 ( .B1(n10112), .B2(n9973), .A(n9832), .ZN(P1_U3273) );
  XNOR2_X1 U11091 ( .A(n9833), .B(n9834), .ZN(n9837) );
  AOI222_X1 U11092 ( .A1(n9918), .A2(n9837), .B1(n9836), .B2(n9913), .C1(n9835), .C2(n9915), .ZN(n9979) );
  XNOR2_X1 U11093 ( .A(n9839), .B(n9838), .ZN(n9980) );
  NAND2_X1 U11094 ( .A1(n10112), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9840) );
  OAI21_X1 U11095 ( .B1(n9922), .B2(n9841), .A(n9840), .ZN(n9842) );
  AOI21_X1 U11096 ( .B1(n9975), .B2(n9929), .A(n9842), .ZN(n9846) );
  NAND2_X1 U11097 ( .A1(n9850), .A2(n9975), .ZN(n9843) );
  AND2_X1 U11098 ( .A1(n4522), .A2(n9843), .ZN(n9977) );
  NAND2_X1 U11099 ( .A1(n9977), .A2(n9844), .ZN(n9845) );
  OAI211_X1 U11100 ( .C1(n9980), .C2(n9926), .A(n9846), .B(n9845), .ZN(n9847)
         );
  INV_X1 U11101 ( .A(n9847), .ZN(n9848) );
  OAI21_X1 U11102 ( .B1(n9979), .B2(n10112), .A(n9848), .ZN(P1_U3274) );
  AOI211_X1 U11103 ( .C1(n9983), .C2(n6101), .A(n9907), .B(n4988), .ZN(n9982)
         );
  INV_X1 U11104 ( .A(n9851), .ZN(n9852) );
  AOI21_X1 U11105 ( .B1(n9860), .B2(n9853), .A(n9852), .ZN(n9854) );
  OAI222_X1 U11106 ( .A1(n9896), .A2(n9856), .B1(n9898), .B2(n9855), .C1(n9893), .C2(n9854), .ZN(n9981) );
  AOI21_X1 U11107 ( .B1(n9982), .B2(n9920), .A(n9981), .ZN(n9865) );
  INV_X1 U11108 ( .A(n9857), .ZN(n9858) );
  OAI22_X1 U11109 ( .A1(n9776), .A2(n9859), .B1(n9858), .B2(n9922), .ZN(n9863)
         );
  XOR2_X1 U11110 ( .A(n9861), .B(n9860), .Z(n9985) );
  NOR2_X1 U11111 ( .A1(n9985), .A2(n9926), .ZN(n9862) );
  AOI211_X1 U11112 ( .C1(n9929), .C2(n9983), .A(n9863), .B(n9862), .ZN(n9864)
         );
  OAI21_X1 U11113 ( .B1(n10112), .B2(n9865), .A(n9864), .ZN(P1_U3275) );
  XNOR2_X1 U11114 ( .A(n9866), .B(n9883), .ZN(n9869) );
  AOI222_X1 U11115 ( .A1(n9918), .A2(n9869), .B1(n9868), .B2(n9915), .C1(n9867), .C2(n9913), .ZN(n9996) );
  AOI21_X1 U11116 ( .B1(n9870), .B2(n5807), .A(n9907), .ZN(n9872) );
  NAND2_X1 U11117 ( .A1(n9872), .A2(n9871), .ZN(n9995) );
  AOI22_X1 U11118 ( .A1(n10112), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9873), 
        .B2(n10110), .ZN(n9875) );
  NAND2_X1 U11119 ( .A1(n5807), .A2(n9929), .ZN(n9874) );
  OAI211_X1 U11120 ( .C1(n9995), .C2(n9876), .A(n9875), .B(n9874), .ZN(n9877)
         );
  INV_X1 U11121 ( .A(n9877), .ZN(n9886) );
  OR2_X1 U11122 ( .A1(n9879), .A2(n9878), .ZN(n9882) );
  NAND2_X1 U11123 ( .A1(n9882), .A2(n9880), .ZN(n9992) );
  NAND2_X1 U11124 ( .A1(n9882), .A2(n9881), .ZN(n9884) );
  NAND2_X1 U11125 ( .A1(n9884), .A2(n9883), .ZN(n9991) );
  NAND3_X1 U11126 ( .A1(n9992), .A2(n9991), .A3(n10119), .ZN(n9885) );
  OAI211_X1 U11127 ( .C1(n9996), .C2(n10112), .A(n9886), .B(n9885), .ZN(
        P1_U3277) );
  XNOR2_X1 U11128 ( .A(n9889), .B(n9888), .ZN(n10006) );
  AOI211_X1 U11129 ( .C1(n10003), .C2(n9905), .A(n9907), .B(n9890), .ZN(n10002) );
  AOI22_X1 U11130 ( .A1(n10112), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9891), 
        .B2(n10110), .ZN(n9892) );
  OAI21_X1 U11131 ( .B1(n4995), .B2(n10115), .A(n9892), .ZN(n9903) );
  AOI211_X1 U11132 ( .C1(n9895), .C2(n9894), .A(n9893), .B(n4453), .ZN(n9901)
         );
  OAI22_X1 U11133 ( .A1(n9899), .A2(n9898), .B1(n9897), .B2(n9896), .ZN(n9900)
         );
  NOR2_X1 U11134 ( .A1(n9901), .A2(n9900), .ZN(n10005) );
  NOR2_X1 U11135 ( .A1(n10005), .A2(n10112), .ZN(n9902) );
  AOI211_X1 U11136 ( .C1(n10002), .C2(n10108), .A(n9903), .B(n9902), .ZN(n9904) );
  OAI21_X1 U11137 ( .B1(n10006), .B2(n9926), .A(n9904), .ZN(P1_U3279) );
  INV_X1 U11138 ( .A(n9905), .ZN(n9906) );
  AOI211_X1 U11139 ( .C1(n10008), .C2(n9908), .A(n9907), .B(n9906), .ZN(n10007) );
  OAI21_X1 U11140 ( .B1(n9910), .B2(n9909), .A(n9925), .ZN(n9912) );
  NAND2_X1 U11141 ( .A1(n9912), .A2(n9911), .ZN(n9917) );
  AOI222_X1 U11142 ( .A1(n9918), .A2(n9917), .B1(n9916), .B2(n9915), .C1(n9914), .C2(n9913), .ZN(n10010) );
  INV_X1 U11143 ( .A(n10010), .ZN(n9919) );
  AOI21_X1 U11144 ( .B1(n10007), .B2(n9920), .A(n9919), .ZN(n9931) );
  INV_X1 U11145 ( .A(n9921), .ZN(n9923) );
  OAI22_X1 U11146 ( .A1(n9776), .A2(n7514), .B1(n9923), .B2(n9922), .ZN(n9928)
         );
  XOR2_X1 U11147 ( .A(n9924), .B(n9925), .Z(n10011) );
  NOR2_X1 U11148 ( .A1(n10011), .A2(n9926), .ZN(n9927) );
  AOI211_X1 U11149 ( .C1(n9929), .C2(n10008), .A(n9928), .B(n9927), .ZN(n9930)
         );
  OAI21_X1 U11150 ( .B1(n9931), .B2(n10112), .A(n9930), .ZN(P1_U3280) );
  INV_X1 U11151 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10566) );
  NOR2_X1 U11152 ( .A1(n4471), .A2(n9932), .ZN(n10012) );
  MUX2_X1 U11153 ( .A(n10566), .B(n10012), .S(n10161), .Z(n9933) );
  OAI21_X1 U11154 ( .B1(n10014), .B2(n9948), .A(n9933), .ZN(P1_U3552) );
  INV_X1 U11155 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9937) );
  MUX2_X1 U11156 ( .A(n9937), .B(n10015), .S(n10161), .Z(n9938) );
  OAI21_X1 U11157 ( .B1(n10018), .B2(n9948), .A(n9938), .ZN(P1_U3549) );
  INV_X1 U11158 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9942) );
  INV_X1 U11159 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9946) );
  AOI211_X1 U11160 ( .C1(n9945), .C2(n10136), .A(n9944), .B(n9943), .ZN(n10023) );
  MUX2_X1 U11161 ( .A(n9946), .B(n10023), .S(n10161), .Z(n9947) );
  OAI21_X1 U11162 ( .B1(n10027), .B2(n9948), .A(n9947), .ZN(P1_U3547) );
  NAND3_X1 U11163 ( .A1(n9753), .A2(n10136), .A3(n9949), .ZN(n9954) );
  AOI22_X1 U11164 ( .A1(n9951), .A2(n9976), .B1(n10148), .B2(n9950), .ZN(n9952) );
  NAND3_X1 U11165 ( .A1(n9954), .A2(n9953), .A3(n9952), .ZN(n10028) );
  MUX2_X1 U11166 ( .A(n10028), .B(P1_REG1_REG_24__SCAN_IN), .S(n10159), .Z(
        P1_U3546) );
  AOI211_X1 U11167 ( .C1(n10148), .C2(n9957), .A(n9956), .B(n9955), .ZN(n9958)
         );
  OAI21_X1 U11168 ( .B1(n10143), .B2(n9959), .A(n9958), .ZN(n10029) );
  MUX2_X1 U11169 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10029), .S(n10161), .Z(
        P1_U3545) );
  AOI22_X1 U11170 ( .A1(n9961), .A2(n9976), .B1(n10148), .B2(n9960), .ZN(n9962) );
  OAI211_X1 U11171 ( .C1(n9964), .C2(n10143), .A(n9963), .B(n9962), .ZN(n10030) );
  MUX2_X1 U11172 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10030), .S(n10161), .Z(
        P1_U3544) );
  AOI21_X1 U11173 ( .B1(n10148), .B2(n9966), .A(n9965), .ZN(n9967) );
  OAI211_X1 U11174 ( .C1(n10143), .C2(n9969), .A(n9968), .B(n9967), .ZN(n10031) );
  MUX2_X1 U11175 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10031), .S(n10161), .Z(
        P1_U3543) );
  AOI21_X1 U11176 ( .B1(n10148), .B2(n9971), .A(n9970), .ZN(n9972) );
  OAI211_X1 U11177 ( .C1(n10143), .C2(n9974), .A(n9973), .B(n9972), .ZN(n10032) );
  MUX2_X1 U11178 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10032), .S(n10161), .Z(
        P1_U3542) );
  AOI22_X1 U11179 ( .A1(n9977), .A2(n9976), .B1(n10148), .B2(n9975), .ZN(n9978) );
  OAI211_X1 U11180 ( .C1(n10143), .C2(n9980), .A(n9979), .B(n9978), .ZN(n10033) );
  MUX2_X1 U11181 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10033), .S(n10161), .Z(
        P1_U3541) );
  AOI211_X1 U11182 ( .C1(n10148), .C2(n9983), .A(n9982), .B(n9981), .ZN(n9984)
         );
  OAI21_X1 U11183 ( .B1(n10143), .B2(n9985), .A(n9984), .ZN(n10034) );
  MUX2_X1 U11184 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10034), .S(n10161), .Z(
        P1_U3540) );
  AOI211_X1 U11185 ( .C1(n10148), .C2(n9988), .A(n9987), .B(n9986), .ZN(n9989)
         );
  OAI21_X1 U11186 ( .B1(n10143), .B2(n9990), .A(n9989), .ZN(n10035) );
  MUX2_X1 U11187 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10035), .S(n10161), .Z(
        P1_U3539) );
  NAND3_X1 U11188 ( .A1(n9992), .A2(n9991), .A3(n10136), .ZN(n9994) );
  NAND2_X1 U11189 ( .A1(n5807), .A2(n10148), .ZN(n9993) );
  NAND4_X1 U11190 ( .A1(n9996), .A2(n9995), .A3(n9994), .A4(n9993), .ZN(n10036) );
  MUX2_X1 U11191 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10036), .S(n10161), .Z(
        P1_U3538) );
  AOI21_X1 U11192 ( .B1(n10148), .B2(n9998), .A(n9997), .ZN(n9999) );
  OAI211_X1 U11193 ( .C1(n10143), .C2(n10001), .A(n10000), .B(n9999), .ZN(
        n10037) );
  MUX2_X1 U11194 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10037), .S(n10161), .Z(
        P1_U3537) );
  AOI21_X1 U11195 ( .B1(n10148), .B2(n10003), .A(n10002), .ZN(n10004) );
  OAI211_X1 U11196 ( .C1(n10143), .C2(n10006), .A(n10005), .B(n10004), .ZN(
        n10038) );
  MUX2_X1 U11197 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10038), .S(n10161), .Z(
        P1_U3536) );
  AOI21_X1 U11198 ( .B1(n10148), .B2(n10008), .A(n10007), .ZN(n10009) );
  OAI211_X1 U11199 ( .C1(n10143), .C2(n10011), .A(n10010), .B(n10009), .ZN(
        n10039) );
  MUX2_X1 U11200 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10039), .S(n10161), .Z(
        P1_U3535) );
  INV_X1 U11201 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10398) );
  MUX2_X1 U11202 ( .A(n10398), .B(n10012), .S(n10155), .Z(n10013) );
  OAI21_X1 U11203 ( .B1(n10014), .B2(n10026), .A(n10013), .ZN(P1_U3520) );
  INV_X1 U11204 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10016) );
  MUX2_X1 U11205 ( .A(n10016), .B(n10015), .S(n10155), .Z(n10017) );
  OAI21_X1 U11206 ( .B1(n10018), .B2(n10026), .A(n10017), .ZN(P1_U3517) );
  INV_X1 U11207 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10020) );
  OAI21_X1 U11208 ( .B1(n10022), .B2(n10026), .A(n10021), .ZN(P1_U3516) );
  INV_X1 U11209 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10024) );
  MUX2_X1 U11210 ( .A(n10024), .B(n10023), .S(n10155), .Z(n10025) );
  OAI21_X1 U11211 ( .B1(n10027), .B2(n10026), .A(n10025), .ZN(P1_U3515) );
  MUX2_X1 U11212 ( .A(n10028), .B(P1_REG0_REG_24__SCAN_IN), .S(n10154), .Z(
        P1_U3514) );
  MUX2_X1 U11213 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10029), .S(n10155), .Z(
        P1_U3513) );
  MUX2_X1 U11214 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10030), .S(n10155), .Z(
        P1_U3512) );
  MUX2_X1 U11215 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10031), .S(n10155), .Z(
        P1_U3511) );
  MUX2_X1 U11216 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10032), .S(n10155), .Z(
        P1_U3510) );
  MUX2_X1 U11217 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10033), .S(n10155), .Z(
        P1_U3509) );
  MUX2_X1 U11218 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10034), .S(n10155), .Z(
        P1_U3507) );
  MUX2_X1 U11219 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10035), .S(n10155), .Z(
        P1_U3504) );
  MUX2_X1 U11220 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10036), .S(n10155), .Z(
        P1_U3501) );
  MUX2_X1 U11221 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10037), .S(n10155), .Z(
        P1_U3498) );
  MUX2_X1 U11222 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10038), .S(n10155), .Z(
        P1_U3495) );
  MUX2_X1 U11223 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n10039), .S(n10155), .Z(
        P1_U3492) );
  INV_X1 U11224 ( .A(n10040), .ZN(n10041) );
  MUX2_X1 U11225 ( .A(n10042), .B(P1_D_REG_0__SCAN_IN), .S(n10122), .Z(
        P1_U3439) );
  NAND2_X1 U11226 ( .A1(n10044), .A2(n10043), .ZN(n10051) );
  INV_X1 U11227 ( .A(n10045), .ZN(n10049) );
  NOR3_X1 U11228 ( .A1(n10046), .A2(P1_IR_REG_28__SCAN_IN), .A3(
        P1_IR_REG_30__SCAN_IN), .ZN(n10048) );
  NAND4_X1 U11229 ( .A1(n10049), .A2(P1_STATE_REG_SCAN_IN), .A3(n10048), .A4(
        n10047), .ZN(n10050) );
  OAI211_X1 U11230 ( .C1(n10440), .C2(n10060), .A(n10051), .B(n10050), .ZN(
        P1_U3324) );
  OAI222_X1 U11231 ( .A1(n10054), .A2(n10060), .B1(n10058), .B2(n10053), .C1(
        P1_U3086), .C2(n4669), .ZN(P1_U3325) );
  OAI222_X1 U11232 ( .A1(n10060), .A2(n10428), .B1(P1_U3086), .B2(n10056), 
        .C1(n10055), .C2(n10058), .ZN(P1_U3326) );
  OAI222_X1 U11233 ( .A1(n10060), .A2(n10059), .B1(P1_U3086), .B2(n6158), .C1(
        n10058), .C2(n10057), .ZN(P1_U3328) );
  MUX2_X1 U11234 ( .A(n10062), .B(n10061), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  INV_X1 U11235 ( .A(n10063), .ZN(n10069) );
  OAI21_X1 U11236 ( .B1(n10066), .B2(n10065), .A(n10064), .ZN(n10068) );
  AOI21_X1 U11237 ( .B1(n10069), .B2(n10068), .A(n10067), .ZN(n10076) );
  AOI21_X1 U11238 ( .B1(n10072), .B2(n10071), .A(n10070), .ZN(n10074) );
  OAI22_X1 U11239 ( .A1(n10074), .A2(n10090), .B1(n10073), .B2(n10088), .ZN(
        n10075) );
  NOR2_X1 U11240 ( .A1(n10076), .A2(n10075), .ZN(n10078) );
  OAI211_X1 U11241 ( .C1(n10098), .C2(n10079), .A(n10078), .B(n10077), .ZN(
        P1_U3252) );
  XNOR2_X1 U11242 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11243 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11244 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10097) );
  AND2_X1 U11245 ( .A1(n10081), .A2(n10080), .ZN(n10084) );
  OAI21_X1 U11246 ( .B1(n10084), .B2(n10083), .A(n10082), .ZN(n10094) );
  AOI21_X1 U11247 ( .B1(n10087), .B2(n10086), .A(n10085), .ZN(n10091) );
  OAI22_X1 U11248 ( .A1(n10091), .A2(n10090), .B1(n10089), .B2(n10088), .ZN(
        n10092) );
  AOI21_X1 U11249 ( .B1(n10094), .B2(n10093), .A(n10092), .ZN(n10096) );
  OAI211_X1 U11250 ( .C1(n10098), .C2(n10097), .A(n10096), .B(n10095), .ZN(
        P1_U3255) );
  NAND2_X1 U11251 ( .A1(n10099), .A2(n10108), .ZN(n10102) );
  AOI22_X1 U11252 ( .A1(n10112), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n10100), 
        .B2(n10110), .ZN(n10101) );
  OAI211_X1 U11253 ( .C1(n10103), .C2(n10115), .A(n10102), .B(n10101), .ZN(
        n10104) );
  AOI21_X1 U11254 ( .B1(n10119), .B2(n10105), .A(n10104), .ZN(n10106) );
  OAI21_X1 U11255 ( .B1(n10112), .B2(n10107), .A(n10106), .ZN(P1_U3287) );
  NAND2_X1 U11256 ( .A1(n10109), .A2(n10108), .ZN(n10114) );
  AOI22_X1 U11257 ( .A1(n10112), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n10111), 
        .B2(n10110), .ZN(n10113) );
  OAI211_X1 U11258 ( .C1(n10116), .C2(n10115), .A(n10114), .B(n10113), .ZN(
        n10117) );
  AOI21_X1 U11259 ( .B1(n10119), .B2(n10118), .A(n10117), .ZN(n10120) );
  OAI21_X1 U11260 ( .B1(n10112), .B2(n10121), .A(n10120), .ZN(P1_U3289) );
  AND2_X1 U11261 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10122), .ZN(P1_U3294) );
  INV_X1 U11262 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10381) );
  NOR2_X1 U11263 ( .A1(n10270), .A2(n10381), .ZN(P1_U3295) );
  AND2_X1 U11264 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10122), .ZN(P1_U3296) );
  AND2_X1 U11265 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10122), .ZN(P1_U3297) );
  AND2_X1 U11266 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10122), .ZN(P1_U3298) );
  AND2_X1 U11267 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10122), .ZN(P1_U3299) );
  AND2_X1 U11268 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10122), .ZN(P1_U3300) );
  AND2_X1 U11269 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10122), .ZN(P1_U3301) );
  INV_X1 U11270 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10399) );
  NOR2_X1 U11271 ( .A1(n10270), .A2(n10399), .ZN(P1_U3302) );
  NOR2_X1 U11272 ( .A1(n10270), .A2(n10345), .ZN(P1_U3303) );
  NOR2_X1 U11273 ( .A1(n10270), .A2(n10522), .ZN(P1_U3304) );
  NOR2_X1 U11274 ( .A1(n10270), .A2(n10486), .ZN(P1_U3305) );
  INV_X1 U11275 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10364) );
  NOR2_X1 U11276 ( .A1(n10270), .A2(n10364), .ZN(P1_U3306) );
  NOR2_X1 U11277 ( .A1(n10270), .A2(n10365), .ZN(P1_U3307) );
  AND2_X1 U11278 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10122), .ZN(P1_U3308) );
  AND2_X1 U11279 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10122), .ZN(P1_U3309) );
  NOR2_X1 U11280 ( .A1(n10270), .A2(n10358), .ZN(P1_U3310) );
  AND2_X1 U11281 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10122), .ZN(P1_U3311) );
  AND2_X1 U11282 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10122), .ZN(P1_U3312) );
  AND2_X1 U11283 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10122), .ZN(P1_U3313) );
  AND2_X1 U11284 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10122), .ZN(P1_U3314) );
  AND2_X1 U11285 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10122), .ZN(P1_U3315) );
  AND2_X1 U11286 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10122), .ZN(P1_U3316) );
  NOR2_X1 U11287 ( .A1(n10270), .A2(n10518), .ZN(P1_U3317) );
  AND2_X1 U11288 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10122), .ZN(P1_U3318) );
  AND2_X1 U11289 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10122), .ZN(P1_U3319) );
  AND2_X1 U11290 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10122), .ZN(P1_U3320) );
  AND2_X1 U11291 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10122), .ZN(P1_U3321) );
  AND2_X1 U11292 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10122), .ZN(P1_U3322) );
  AND2_X1 U11293 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10122), .ZN(P1_U3323) );
  INV_X1 U11294 ( .A(n10123), .ZN(n10127) );
  OAI21_X1 U11295 ( .B1(n7378), .B2(n10131), .A(n10124), .ZN(n10126) );
  AOI211_X1 U11296 ( .C1(n10128), .C2(n10127), .A(n10126), .B(n10125), .ZN(
        n10156) );
  INV_X1 U11297 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10129) );
  AOI22_X1 U11298 ( .A1(n10155), .A2(n10156), .B1(n10129), .B2(n10154), .ZN(
        P1_U3456) );
  OAI21_X1 U11299 ( .B1(n10132), .B2(n10131), .A(n10130), .ZN(n10134) );
  AOI211_X1 U11300 ( .C1(n10136), .C2(n10135), .A(n10134), .B(n10133), .ZN(
        n10157) );
  INV_X1 U11301 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10137) );
  AOI22_X1 U11302 ( .A1(n10155), .A2(n10157), .B1(n10137), .B2(n10154), .ZN(
        P1_U3462) );
  AOI21_X1 U11303 ( .B1(n10148), .B2(n10139), .A(n10138), .ZN(n10140) );
  OAI211_X1 U11304 ( .C1(n10143), .C2(n10142), .A(n10141), .B(n10140), .ZN(
        n10144) );
  INV_X1 U11305 ( .A(n10144), .ZN(n10158) );
  INV_X1 U11306 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10145) );
  AOI22_X1 U11307 ( .A1(n10155), .A2(n10158), .B1(n10145), .B2(n10154), .ZN(
        P1_U3468) );
  AOI21_X1 U11308 ( .B1(n10148), .B2(n10147), .A(n10146), .ZN(n10149) );
  OAI211_X1 U11309 ( .C1(n10152), .C2(n10151), .A(n10150), .B(n10149), .ZN(
        n10153) );
  INV_X1 U11310 ( .A(n10153), .ZN(n10160) );
  INV_X1 U11311 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U11312 ( .A1(n10155), .A2(n10160), .B1(n10458), .B2(n10154), .ZN(
        P1_U3474) );
  AOI22_X1 U11313 ( .A1(n10161), .A2(n10156), .B1(n7038), .B2(n10159), .ZN(
        P1_U3523) );
  AOI22_X1 U11314 ( .A1(n10161), .A2(n10157), .B1(n7041), .B2(n10159), .ZN(
        P1_U3525) );
  AOI22_X1 U11315 ( .A1(n10161), .A2(n10158), .B1(n10425), .B2(n10159), .ZN(
        P1_U3527) );
  AOI22_X1 U11316 ( .A1(n10161), .A2(n10160), .B1(n10489), .B2(n10159), .ZN(
        P1_U3529) );
  XNOR2_X1 U11317 ( .A(n10162), .B(n10164), .ZN(n10214) );
  NAND3_X1 U11318 ( .A1(n7431), .A2(n10164), .A3(n10163), .ZN(n10165) );
  NAND2_X1 U11319 ( .A1(n10166), .A2(n10165), .ZN(n10170) );
  AOI222_X1 U11320 ( .A1(n10171), .A2(n10170), .B1(n10169), .B2(n10168), .C1(
        n7255), .C2(n10167), .ZN(n10210) );
  INV_X1 U11321 ( .A(n10210), .ZN(n10172) );
  AOI21_X1 U11322 ( .B1(n10173), .B2(n10214), .A(n10172), .ZN(n10182) );
  INV_X1 U11323 ( .A(n10174), .ZN(n10176) );
  AOI222_X1 U11324 ( .A1(n10179), .A2(n10178), .B1(n10214), .B2(n10177), .C1(
        n10176), .C2(n10175), .ZN(n10180) );
  OAI221_X1 U11325 ( .B1(n10183), .B2(n10182), .C1(n10181), .C2(n4919), .A(
        n10180), .ZN(P2_U3228) );
  AOI21_X1 U11326 ( .B1(n10185), .B2(n10225), .A(n10184), .ZN(n10186) );
  AOI211_X1 U11327 ( .C1(n10189), .C2(n10188), .A(n10187), .B(n10186), .ZN(
        n10231) );
  INV_X1 U11328 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U11329 ( .A1(n10230), .A2(n10231), .B1(n10330), .B2(n10229), .ZN(
        P2_U3390) );
  AOI22_X1 U11330 ( .A1(n10190), .A2(n10198), .B1(n6191), .B2(n10189), .ZN(
        n10191) );
  AND2_X1 U11331 ( .A1(n10192), .A2(n10191), .ZN(n10233) );
  INV_X1 U11332 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10193) );
  AOI22_X1 U11333 ( .A1(n10230), .A2(n10233), .B1(n10193), .B2(n10229), .ZN(
        P2_U3393) );
  INV_X1 U11334 ( .A(n10194), .ZN(n10196) );
  AOI211_X1 U11335 ( .C1(n10198), .C2(n10197), .A(n10196), .B(n10195), .ZN(
        n10235) );
  INV_X1 U11336 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10199) );
  AOI22_X1 U11337 ( .A1(n10230), .A2(n10235), .B1(n10199), .B2(n10229), .ZN(
        P2_U3396) );
  INV_X1 U11338 ( .A(n10200), .ZN(n10204) );
  OAI22_X1 U11339 ( .A1(n10202), .A2(n10225), .B1(n10201), .B2(n10223), .ZN(
        n10203) );
  NOR2_X1 U11340 ( .A1(n10204), .A2(n10203), .ZN(n10237) );
  AOI22_X1 U11341 ( .A1(n10230), .A2(n10237), .B1(n6211), .B2(n10229), .ZN(
        P2_U3399) );
  NOR2_X1 U11342 ( .A1(n10205), .A2(n10223), .ZN(n10207) );
  AOI211_X1 U11343 ( .C1(n10213), .C2(n10208), .A(n10207), .B(n10206), .ZN(
        n10239) );
  INV_X1 U11344 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10209) );
  AOI22_X1 U11345 ( .A1(n10230), .A2(n10239), .B1(n10209), .B2(n10229), .ZN(
        P2_U3402) );
  OAI21_X1 U11346 ( .B1(n10211), .B2(n10223), .A(n10210), .ZN(n10212) );
  AOI21_X1 U11347 ( .B1(n10214), .B2(n10213), .A(n10212), .ZN(n10241) );
  INV_X1 U11348 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10215) );
  AOI22_X1 U11349 ( .A1(n10230), .A2(n10241), .B1(n10215), .B2(n10229), .ZN(
        P2_U3405) );
  INV_X1 U11350 ( .A(n10216), .ZN(n10220) );
  OAI22_X1 U11351 ( .A1(n10218), .A2(n10225), .B1(n10217), .B2(n10223), .ZN(
        n10219) );
  NOR2_X1 U11352 ( .A1(n10220), .A2(n10219), .ZN(n10243) );
  INV_X1 U11353 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10221) );
  AOI22_X1 U11354 ( .A1(n10230), .A2(n10243), .B1(n10221), .B2(n10229), .ZN(
        P2_U3408) );
  INV_X1 U11355 ( .A(n10222), .ZN(n10228) );
  OAI22_X1 U11356 ( .A1(n10226), .A2(n10225), .B1(n10224), .B2(n10223), .ZN(
        n10227) );
  NOR2_X1 U11357 ( .A1(n10228), .A2(n10227), .ZN(n10244) );
  AOI22_X1 U11358 ( .A1(n10230), .A2(n10244), .B1(n6277), .B2(n10229), .ZN(
        P2_U3414) );
  AOI22_X1 U11359 ( .A1(n10245), .A2(n10231), .B1(n5411), .B2(n6586), .ZN(
        P2_U3459) );
  AOI22_X1 U11360 ( .A1(n10245), .A2(n10233), .B1(n10232), .B2(n6586), .ZN(
        P2_U3460) );
  AOI22_X1 U11361 ( .A1(n10245), .A2(n10235), .B1(n10234), .B2(n6586), .ZN(
        P2_U3461) );
  AOI22_X1 U11362 ( .A1(n10245), .A2(n10237), .B1(n10236), .B2(n6586), .ZN(
        P2_U3462) );
  AOI22_X1 U11363 ( .A1(n10245), .A2(n10239), .B1(n10238), .B2(n6586), .ZN(
        P2_U3463) );
  AOI22_X1 U11364 ( .A1(n10245), .A2(n10241), .B1(n10240), .B2(n6586), .ZN(
        P2_U3464) );
  AOI22_X1 U11365 ( .A1(n10245), .A2(n10243), .B1(n10242), .B2(n6586), .ZN(
        P2_U3465) );
  AOI22_X1 U11366 ( .A1(n10245), .A2(n10244), .B1(n5424), .B2(n6586), .ZN(
        P2_U3467) );
  NOR2_X1 U11367 ( .A1(n10247), .A2(n10246), .ZN(n10248) );
  XOR2_X1 U11368 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10248), .Z(ADD_1068_U5) );
  XOR2_X1 U11369 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11370 ( .A1(n10250), .A2(n10249), .ZN(n10251) );
  XNOR2_X1 U11371 ( .A(n10251), .B(n10333), .ZN(ADD_1068_U55) );
  XNOR2_X1 U11372 ( .A(n10253), .B(n10252), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11373 ( .A(n10255), .B(n10254), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11374 ( .A(n10257), .B(n10256), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11375 ( .A(n10259), .B(n10258), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11376 ( .A(n10261), .B(n10260), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11377 ( .A(n10263), .B(n10262), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11378 ( .A(n10265), .B(n10264), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11379 ( .A(n10267), .B(n10266), .ZN(ADD_1068_U63) );
  OAI22_X1 U11380 ( .A1(n10270), .A2(P1_D_REG_1__SCAN_IN), .B1(n10269), .B2(
        n10268), .ZN(n10582) );
  INV_X1 U11381 ( .A(SI_0_), .ZN(n10538) );
  NOR4_X1 U11382 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(n10538), .A3(n10517), .A4(
        n10518), .ZN(n10282) );
  NOR4_X1 U11383 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(P2_DATAO_REG_13__SCAN_IN), 
        .A3(P2_IR_REG_30__SCAN_IN), .A4(P2_REG0_REG_22__SCAN_IN), .ZN(n10281)
         );
  INV_X1 U11384 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10273) );
  NOR4_X1 U11385 ( .A1(n10273), .A2(n10272), .A3(n10271), .A4(
        P2_REG0_REG_30__SCAN_IN), .ZN(n10280) );
  NOR4_X1 U11386 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .A3(P1_ADDR_REG_3__SCAN_IN), .A4(n10344), .ZN(n10276) );
  NOR4_X1 U11387 ( .A1(P2_REG1_REG_19__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .A3(P1_ADDR_REG_5__SCAN_IN), .A4(n10342), .ZN(n10275) );
  AND4_X1 U11388 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_24__SCAN_IN), 
        .A3(P1_REG1_REG_27__SCAN_IN), .A4(n10520), .ZN(n10274) );
  NAND4_X1 U11389 ( .A1(n10533), .A2(n10276), .A3(n10275), .A4(n10274), .ZN(
        n10278) );
  NOR4_X1 U11390 ( .A1(n10531), .A2(n10278), .A3(n10277), .A4(n10522), .ZN(
        n10279) );
  AND4_X1 U11391 ( .A1(n10282), .A2(n10281), .A3(n10280), .A4(n10279), .ZN(
        n10325) );
  NAND4_X1 U11392 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n10426), .A3(n10425), 
        .A4(n7773), .ZN(n10287) );
  INV_X1 U11393 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10431) );
  NAND4_X1 U11394 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), 
        .A3(n10431), .A4(n10283), .ZN(n10286) );
  INV_X1 U11395 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10439) );
  NAND4_X1 U11396 ( .A1(SI_20_), .A2(n10284), .A3(n10439), .A4(n10440), .ZN(
        n10285) );
  NOR4_X1 U11397 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(n10287), .A3(n10286), 
        .A4(n10285), .ZN(n10323) );
  NAND4_X1 U11398 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .A3(
        P1_IR_REG_2__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n10291) );
  NAND4_X1 U11399 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .A3(P1_REG0_REG_4__SCAN_IN), .A4(n10396), .ZN(n10290) );
  NAND4_X1 U11400 ( .A1(SI_29_), .A2(SI_9_), .A3(n10416), .A4(n9859), .ZN(
        n10289) );
  INV_X1 U11401 ( .A(P1_B_REG_SCAN_IN), .ZN(n10412) );
  NAND4_X1 U11402 ( .A1(P1_REG2_REG_23__SCAN_IN), .A2(n10411), .A3(n10412), 
        .A4(n10398), .ZN(n10288) );
  NOR4_X1 U11403 ( .A1(n10291), .A2(n10290), .A3(n10289), .A4(n10288), .ZN(
        n10322) );
  NAND4_X1 U11404 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .A3(P2_REG0_REG_3__SCAN_IN), .A4(P1_IR_REG_21__SCAN_IN), .ZN(n10292)
         );
  NOR3_X1 U11405 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .A3(
        n10292), .ZN(n10321) );
  NAND4_X1 U11406 ( .A1(n10294), .A2(n10293), .A3(P2_REG2_REG_13__SCAN_IN), 
        .A4(P2_REG1_REG_0__SCAN_IN), .ZN(n10297) );
  INV_X1 U11407 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10295) );
  NAND4_X1 U11408 ( .A1(n10295), .A2(P1_IR_REG_17__SCAN_IN), .A3(
        P2_REG1_REG_12__SCAN_IN), .A4(P2_REG0_REG_0__SCAN_IN), .ZN(n10296) );
  NOR2_X1 U11409 ( .A1(n10297), .A2(n10296), .ZN(n10306) );
  NAND2_X1 U11410 ( .A1(n10298), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n10304) );
  NAND4_X1 U11411 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P1_DATAO_REG_23__SCAN_IN), 
        .A3(P1_REG0_REG_19__SCAN_IN), .A4(P1_REG0_REG_15__SCAN_IN), .ZN(n10300) );
  NAND4_X1 U11412 ( .A1(P2_REG0_REG_13__SCAN_IN), .A2(P2_REG1_REG_15__SCAN_IN), 
        .A3(P1_REG0_REG_0__SCAN_IN), .A4(n10376), .ZN(n10299) );
  NOR2_X1 U11413 ( .A1(n10300), .A2(n10299), .ZN(n10302) );
  AND4_X1 U11414 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(n10564), .A3(n10563), .A4(
        n10547), .ZN(n10301) );
  NAND4_X1 U11415 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(n10302), .A3(n10458), .A4(
        n10301), .ZN(n10303) );
  NOR2_X1 U11416 ( .A1(n10304), .A2(n10303), .ZN(n10305) );
  INV_X1 U11417 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10459) );
  NAND4_X1 U11418 ( .A1(n10306), .A2(P2_D_REG_31__SCAN_IN), .A3(n10305), .A4(
        n10459), .ZN(n10308) );
  NAND4_X1 U11419 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n10367), .A3(n10356), 
        .A4(n10368), .ZN(n10307) );
  NOR2_X1 U11420 ( .A1(n10308), .A2(n10307), .ZN(n10319) );
  INV_X1 U11421 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n10473) );
  NAND4_X1 U11422 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(
        P2_DATAO_REG_24__SCAN_IN), .A3(P2_REG2_REG_17__SCAN_IN), .A4(n10473), 
        .ZN(n10310) );
  INV_X1 U11423 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10544) );
  NAND4_X1 U11424 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(n6232), .A3(n10545), .A4(
        n10544), .ZN(n10309) );
  NOR2_X1 U11425 ( .A1(n10310), .A2(n10309), .ZN(n10318) );
  NAND4_X1 U11426 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), 
        .A3(n10477), .A4(n4853), .ZN(n10312) );
  NAND4_X1 U11427 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(P1_REG1_REG_30__SCAN_IN), 
        .A3(n10559), .A4(n9692), .ZN(n10311) );
  NOR2_X1 U11428 ( .A1(n10312), .A2(n10311), .ZN(n10317) );
  INV_X1 U11429 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10327) );
  NAND4_X1 U11430 ( .A1(P1_REG1_REG_1__SCAN_IN), .A2(P2_ADDR_REG_18__SCAN_IN), 
        .A3(n10334), .A4(n10327), .ZN(n10315) );
  NAND4_X1 U11431 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_REG1_REG_9__SCAN_IN), 
        .A3(n10504), .A4(n10505), .ZN(n10314) );
  NAND4_X1 U11432 ( .A1(n10359), .A2(P1_REG1_REG_7__SCAN_IN), .A3(
        P1_IR_REG_4__SCAN_IN), .A4(P1_REG2_REG_17__SCAN_IN), .ZN(n10313) );
  NOR3_X1 U11433 ( .A1(n10315), .A2(n10314), .A3(n10313), .ZN(n10316) );
  AND4_X1 U11434 ( .A1(n10319), .A2(n10318), .A3(n10317), .A4(n10316), .ZN(
        n10320) );
  AND4_X1 U11435 ( .A1(n10323), .A2(n10322), .A3(n10321), .A4(n10320), .ZN(
        n10324) );
  AOI21_X1 U11436 ( .B1(n10325), .B2(n10324), .A(P2_IR_REG_23__SCAN_IN), .ZN(
        n10580) );
  AOI22_X1 U11437 ( .A1(n10328), .A2(keyinput62), .B1(keyinput98), .B2(n10327), 
        .ZN(n10326) );
  OAI221_X1 U11438 ( .B1(n10328), .B2(keyinput62), .C1(n10327), .C2(keyinput98), .A(n10326), .ZN(n10340) );
  INV_X1 U11439 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10331) );
  AOI22_X1 U11440 ( .A1(n10331), .A2(keyinput96), .B1(n10330), .B2(keyinput65), 
        .ZN(n10329) );
  OAI221_X1 U11441 ( .B1(n10331), .B2(keyinput96), .C1(n10330), .C2(keyinput65), .A(n10329), .ZN(n10339) );
  AOI22_X1 U11442 ( .A1(n10334), .A2(keyinput67), .B1(keyinput16), .B2(n10333), 
        .ZN(n10332) );
  OAI221_X1 U11443 ( .B1(n10334), .B2(keyinput67), .C1(n10333), .C2(keyinput16), .A(n10332), .ZN(n10338) );
  XNOR2_X1 U11444 ( .A(P1_REG2_REG_17__SCAN_IN), .B(keyinput40), .ZN(n10336)
         );
  XNOR2_X1 U11445 ( .A(SI_5_), .B(keyinput101), .ZN(n10335) );
  NAND2_X1 U11446 ( .A1(n10336), .A2(n10335), .ZN(n10337) );
  NOR4_X1 U11447 ( .A1(n10340), .A2(n10339), .A3(n10338), .A4(n10337), .ZN(
        n10393) );
  AOI22_X1 U11448 ( .A1(n10342), .A2(keyinput31), .B1(P2_U3151), .B2(
        keyinput28), .ZN(n10341) );
  OAI221_X1 U11449 ( .B1(n10342), .B2(keyinput31), .C1(P2_U3151), .C2(
        keyinput28), .A(n10341), .ZN(n10354) );
  AOI22_X1 U11450 ( .A1(n10345), .A2(keyinput15), .B1(keyinput54), .B2(n10344), 
        .ZN(n10343) );
  OAI221_X1 U11451 ( .B1(n10345), .B2(keyinput15), .C1(n10344), .C2(keyinput54), .A(n10343), .ZN(n10353) );
  AOI22_X1 U11452 ( .A1(n7038), .A2(keyinput112), .B1(n10347), .B2(keyinput12), 
        .ZN(n10346) );
  OAI221_X1 U11453 ( .B1(n7038), .B2(keyinput112), .C1(n10347), .C2(keyinput12), .A(n10346), .ZN(n10352) );
  INV_X1 U11454 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U11455 ( .A1(n10350), .A2(keyinput55), .B1(n10349), .B2(keyinput66), 
        .ZN(n10348) );
  OAI221_X1 U11456 ( .B1(n10350), .B2(keyinput55), .C1(n10349), .C2(keyinput66), .A(n10348), .ZN(n10351) );
  NOR4_X1 U11457 ( .A1(n10354), .A2(n10353), .A3(n10352), .A4(n10351), .ZN(
        n10392) );
  AOI22_X1 U11458 ( .A1(n10357), .A2(keyinput118), .B1(n10356), .B2(keyinput99), .ZN(n10355) );
  OAI221_X1 U11459 ( .B1(n10357), .B2(keyinput118), .C1(n10356), .C2(
        keyinput99), .A(n10355), .ZN(n10362) );
  XNOR2_X1 U11460 ( .A(n10358), .B(keyinput75), .ZN(n10361) );
  XNOR2_X1 U11461 ( .A(n10359), .B(keyinput111), .ZN(n10360) );
  OR3_X1 U11462 ( .A1(n10362), .A2(n10361), .A3(n10360), .ZN(n10371) );
  AOI22_X1 U11463 ( .A1(n10365), .A2(keyinput42), .B1(n10364), .B2(keyinput114), .ZN(n10363) );
  OAI221_X1 U11464 ( .B1(n10365), .B2(keyinput42), .C1(n10364), .C2(
        keyinput114), .A(n10363), .ZN(n10370) );
  AOI22_X1 U11465 ( .A1(n10368), .A2(keyinput41), .B1(n10367), .B2(keyinput124), .ZN(n10366) );
  OAI221_X1 U11466 ( .B1(n10368), .B2(keyinput41), .C1(n10367), .C2(
        keyinput124), .A(n10366), .ZN(n10369) );
  NOR3_X1 U11467 ( .A1(n10371), .A2(n10370), .A3(n10369), .ZN(n10391) );
  AOI22_X1 U11468 ( .A1(n10374), .A2(keyinput46), .B1(n10373), .B2(keyinput72), 
        .ZN(n10372) );
  OAI221_X1 U11469 ( .B1(n10374), .B2(keyinput46), .C1(n10373), .C2(keyinput72), .A(n10372), .ZN(n10379) );
  AOI22_X1 U11470 ( .A1(n10377), .A2(keyinput47), .B1(keyinput73), .B2(n10376), 
        .ZN(n10375) );
  OAI221_X1 U11471 ( .B1(n10377), .B2(keyinput47), .C1(n10376), .C2(keyinput73), .A(n10375), .ZN(n10378) );
  NOR2_X1 U11472 ( .A1(n10379), .A2(n10378), .ZN(n10389) );
  INV_X1 U11473 ( .A(keyinput126), .ZN(n10380) );
  XNOR2_X1 U11474 ( .A(n10381), .B(n10380), .ZN(n10388) );
  XNOR2_X1 U11475 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput80), .ZN(n10387)
         );
  AOI22_X1 U11476 ( .A1(n10384), .A2(keyinput38), .B1(n10383), .B2(keyinput52), 
        .ZN(n10382) );
  OAI221_X1 U11477 ( .B1(n10384), .B2(keyinput38), .C1(n10383), .C2(keyinput52), .A(n10382), .ZN(n10385) );
  INV_X1 U11478 ( .A(n10385), .ZN(n10386) );
  AND4_X1 U11479 ( .A1(n10389), .A2(n10388), .A3(n10387), .A4(n10386), .ZN(
        n10390) );
  NAND4_X1 U11480 ( .A1(n10393), .A2(n10392), .A3(n10391), .A4(n10390), .ZN(
        n10578) );
  INV_X1 U11481 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10395) );
  AOI22_X1 U11482 ( .A1(n10396), .A2(keyinput25), .B1(keyinput36), .B2(n10395), 
        .ZN(n10394) );
  OAI221_X1 U11483 ( .B1(n10396), .B2(keyinput25), .C1(n10395), .C2(keyinput36), .A(n10394), .ZN(n10409) );
  AOI22_X1 U11484 ( .A1(n5356), .A2(keyinput95), .B1(keyinput105), .B2(n10398), 
        .ZN(n10397) );
  OAI221_X1 U11485 ( .B1(n5356), .B2(keyinput95), .C1(n10398), .C2(keyinput105), .A(n10397), .ZN(n10403) );
  XNOR2_X1 U11486 ( .A(n10399), .B(keyinput35), .ZN(n10402) );
  XNOR2_X1 U11487 ( .A(n10400), .B(keyinput9), .ZN(n10401) );
  OR3_X1 U11488 ( .A1(n10403), .A2(n10402), .A3(n10401), .ZN(n10408) );
  AOI22_X1 U11489 ( .A1(n10406), .A2(keyinput14), .B1(keyinput82), .B2(n10405), 
        .ZN(n10404) );
  OAI221_X1 U11490 ( .B1(n10406), .B2(keyinput14), .C1(n10405), .C2(keyinput82), .A(n10404), .ZN(n10407) );
  NOR3_X1 U11491 ( .A1(n10409), .A2(n10408), .A3(n10407), .ZN(n10456) );
  AOI22_X1 U11492 ( .A1(n10412), .A2(keyinput120), .B1(n10411), .B2(
        keyinput109), .ZN(n10410) );
  OAI221_X1 U11493 ( .B1(n10412), .B2(keyinput120), .C1(n10411), .C2(
        keyinput109), .A(n10410), .ZN(n10423) );
  AOI22_X1 U11494 ( .A1(n9775), .A2(keyinput102), .B1(keyinput121), .B2(n10414), .ZN(n10413) );
  OAI221_X1 U11495 ( .B1(n9775), .B2(keyinput102), .C1(n10414), .C2(
        keyinput121), .A(n10413), .ZN(n10422) );
  AOI22_X1 U11496 ( .A1(n9859), .A2(keyinput113), .B1(n10416), .B2(keyinput18), 
        .ZN(n10415) );
  OAI221_X1 U11497 ( .B1(n9859), .B2(keyinput113), .C1(n10416), .C2(keyinput18), .A(n10415), .ZN(n10421) );
  AOI22_X1 U11498 ( .A1(n10419), .A2(keyinput6), .B1(keyinput1), .B2(n10418), 
        .ZN(n10417) );
  OAI221_X1 U11499 ( .B1(n10419), .B2(keyinput6), .C1(n10418), .C2(keyinput1), 
        .A(n10417), .ZN(n10420) );
  NOR4_X1 U11500 ( .A1(n10423), .A2(n10422), .A3(n10421), .A4(n10420), .ZN(
        n10455) );
  AOI22_X1 U11501 ( .A1(n10426), .A2(keyinput86), .B1(keyinput5), .B2(n10425), 
        .ZN(n10424) );
  OAI221_X1 U11502 ( .B1(n10426), .B2(keyinput86), .C1(n10425), .C2(keyinput5), 
        .A(n10424), .ZN(n10437) );
  AOI22_X1 U11503 ( .A1(n10428), .A2(keyinput90), .B1(keyinput24), .B2(n7773), 
        .ZN(n10427) );
  OAI221_X1 U11504 ( .B1(n10428), .B2(keyinput90), .C1(n7773), .C2(keyinput24), 
        .A(n10427), .ZN(n10436) );
  AOI22_X1 U11505 ( .A1(n10431), .A2(keyinput87), .B1(n10430), .B2(keyinput115), .ZN(n10429) );
  OAI221_X1 U11506 ( .B1(n10431), .B2(keyinput87), .C1(n10430), .C2(
        keyinput115), .A(n10429), .ZN(n10435) );
  XNOR2_X1 U11507 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput11), .ZN(n10433)
         );
  XNOR2_X1 U11508 ( .A(keyinput8), .B(P1_REG3_REG_1__SCAN_IN), .ZN(n10432) );
  NAND2_X1 U11509 ( .A1(n10433), .A2(n10432), .ZN(n10434) );
  NOR4_X1 U11510 ( .A1(n10437), .A2(n10436), .A3(n10435), .A4(n10434), .ZN(
        n10454) );
  AOI22_X1 U11511 ( .A1(n10440), .A2(keyinput110), .B1(n10439), .B2(keyinput74), .ZN(n10438) );
  OAI221_X1 U11512 ( .B1(n10440), .B2(keyinput110), .C1(n10439), .C2(
        keyinput74), .A(n10438), .ZN(n10452) );
  INV_X1 U11513 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U11514 ( .A1(n10443), .A2(keyinput4), .B1(n10442), .B2(keyinput50), 
        .ZN(n10441) );
  OAI221_X1 U11515 ( .B1(n10443), .B2(keyinput4), .C1(n10442), .C2(keyinput50), 
        .A(n10441), .ZN(n10451) );
  AOI22_X1 U11516 ( .A1(n10446), .A2(keyinput53), .B1(n10445), .B2(keyinput68), 
        .ZN(n10444) );
  OAI221_X1 U11517 ( .B1(n10446), .B2(keyinput53), .C1(n10445), .C2(keyinput68), .A(n10444), .ZN(n10450) );
  XNOR2_X1 U11518 ( .A(P2_REG0_REG_22__SCAN_IN), .B(keyinput117), .ZN(n10448)
         );
  XNOR2_X1 U11519 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput21), .ZN(n10447) );
  NAND2_X1 U11520 ( .A1(n10448), .A2(n10447), .ZN(n10449) );
  NOR4_X1 U11521 ( .A1(n10452), .A2(n10451), .A3(n10450), .A4(n10449), .ZN(
        n10453) );
  NAND4_X1 U11522 ( .A1(n10456), .A2(n10455), .A3(n10454), .A4(n10453), .ZN(
        n10577) );
  AOI22_X1 U11523 ( .A1(n10459), .A2(keyinput60), .B1(keyinput77), .B2(n10458), 
        .ZN(n10457) );
  OAI221_X1 U11524 ( .B1(n10459), .B2(keyinput60), .C1(n10458), .C2(keyinput77), .A(n10457), .ZN(n10469) );
  AOI22_X1 U11525 ( .A1(n10461), .A2(keyinput23), .B1(keyinput123), .B2(n10047), .ZN(n10460) );
  OAI221_X1 U11526 ( .B1(n10461), .B2(keyinput23), .C1(n10047), .C2(
        keyinput123), .A(n10460), .ZN(n10468) );
  XNOR2_X1 U11527 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput44), .ZN(n10464) );
  XNOR2_X1 U11528 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput79), .ZN(n10463) );
  XNOR2_X1 U11529 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput26), .ZN(n10462) );
  NAND3_X1 U11530 ( .A1(n10464), .A2(n10463), .A3(n10462), .ZN(n10467) );
  XNOR2_X1 U11531 ( .A(n10465), .B(keyinput88), .ZN(n10466) );
  NOR4_X1 U11532 ( .A1(n10469), .A2(n10468), .A3(n10467), .A4(n10466), .ZN(
        n10515) );
  AOI22_X1 U11533 ( .A1(n10471), .A2(keyinput107), .B1(keyinput78), .B2(n4853), 
        .ZN(n10470) );
  OAI221_X1 U11534 ( .B1(n10471), .B2(keyinput107), .C1(n4853), .C2(keyinput78), .A(n10470), .ZN(n10484) );
  AOI22_X1 U11535 ( .A1(n10474), .A2(keyinput125), .B1(n10473), .B2(keyinput92), .ZN(n10472) );
  OAI221_X1 U11536 ( .B1(n10474), .B2(keyinput125), .C1(n10473), .C2(
        keyinput92), .A(n10472), .ZN(n10483) );
  AOI22_X1 U11537 ( .A1(n10477), .A2(keyinput58), .B1(keyinput69), .B2(n10476), 
        .ZN(n10475) );
  OAI221_X1 U11538 ( .B1(n10477), .B2(keyinput58), .C1(n10476), .C2(keyinput69), .A(n10475), .ZN(n10482) );
  INV_X1 U11539 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U11540 ( .A1(n10480), .A2(keyinput32), .B1(keyinput89), .B2(n10479), 
        .ZN(n10478) );
  OAI221_X1 U11541 ( .B1(n10480), .B2(keyinput32), .C1(n10479), .C2(keyinput89), .A(n10478), .ZN(n10481) );
  NOR4_X1 U11542 ( .A1(n10484), .A2(n10483), .A3(n10482), .A4(n10481), .ZN(
        n10514) );
  INV_X1 U11543 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U11544 ( .A1(n10487), .A2(keyinput43), .B1(n10486), .B2(keyinput61), 
        .ZN(n10485) );
  OAI221_X1 U11545 ( .B1(n10487), .B2(keyinput43), .C1(n10486), .C2(keyinput61), .A(n10485), .ZN(n10497) );
  XNOR2_X1 U11546 ( .A(keyinput39), .B(n10488), .ZN(n10496) );
  XNOR2_X1 U11547 ( .A(keyinput84), .B(n10489), .ZN(n10495) );
  XNOR2_X1 U11548 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput103), .ZN(n10493) );
  XNOR2_X1 U11549 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput10), .ZN(n10492) );
  XNOR2_X1 U11550 ( .A(P2_IR_REG_0__SCAN_IN), .B(keyinput127), .ZN(n10491) );
  XNOR2_X1 U11551 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(keyinput33), .ZN(n10490)
         );
  NAND4_X1 U11552 ( .A1(n10493), .A2(n10492), .A3(n10491), .A4(n10490), .ZN(
        n10494) );
  NOR4_X1 U11553 ( .A1(n10497), .A2(n10496), .A3(n10495), .A4(n10494), .ZN(
        n10513) );
  AOI22_X1 U11554 ( .A1(n10500), .A2(keyinput20), .B1(n10499), .B2(keyinput34), 
        .ZN(n10498) );
  OAI221_X1 U11555 ( .B1(n10500), .B2(keyinput20), .C1(n10499), .C2(keyinput34), .A(n10498), .ZN(n10511) );
  AOI22_X1 U11556 ( .A1(n6211), .A2(keyinput27), .B1(n10502), .B2(keyinput59), 
        .ZN(n10501) );
  OAI221_X1 U11557 ( .B1(n6211), .B2(keyinput27), .C1(n10502), .C2(keyinput59), 
        .A(n10501), .ZN(n10510) );
  AOI22_X1 U11558 ( .A1(n10505), .A2(keyinput97), .B1(keyinput93), .B2(n10504), 
        .ZN(n10503) );
  OAI221_X1 U11559 ( .B1(n10505), .B2(keyinput97), .C1(n10504), .C2(keyinput93), .A(n10503), .ZN(n10509) );
  XOR2_X1 U11560 ( .A(n5411), .B(keyinput13), .Z(n10507) );
  XNOR2_X1 U11561 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput122), .ZN(n10506) );
  NAND2_X1 U11562 ( .A1(n10507), .A2(n10506), .ZN(n10508) );
  NOR4_X1 U11563 ( .A1(n10511), .A2(n10510), .A3(n10509), .A4(n10508), .ZN(
        n10512) );
  NAND4_X1 U11564 ( .A1(n10515), .A2(n10514), .A3(n10513), .A4(n10512), .ZN(
        n10576) );
  AOI22_X1 U11565 ( .A1(n10518), .A2(keyinput17), .B1(n10517), .B2(keyinput106), .ZN(n10516) );
  OAI221_X1 U11566 ( .B1(n10518), .B2(keyinput17), .C1(n10517), .C2(
        keyinput106), .A(n10516), .ZN(n10529) );
  AOI22_X1 U11567 ( .A1(n10521), .A2(keyinput81), .B1(n10520), .B2(keyinput70), 
        .ZN(n10519) );
  OAI221_X1 U11568 ( .B1(n10521), .B2(keyinput81), .C1(n10520), .C2(keyinput70), .A(n10519), .ZN(n10528) );
  XOR2_X1 U11569 ( .A(n10522), .B(keyinput76), .Z(n10526) );
  XNOR2_X1 U11570 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput22), .ZN(n10525)
         );
  XNOR2_X1 U11571 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput49), .ZN(n10524) );
  XNOR2_X1 U11572 ( .A(P1_REG1_REG_27__SCAN_IN), .B(keyinput0), .ZN(n10523) );
  NAND4_X1 U11573 ( .A1(n10526), .A2(n10525), .A3(n10524), .A4(n10523), .ZN(
        n10527) );
  NOR3_X1 U11574 ( .A1(n10529), .A2(n10528), .A3(n10527), .ZN(n10574) );
  AOI22_X1 U11575 ( .A1(n10532), .A2(keyinput57), .B1(n10531), .B2(keyinput116), .ZN(n10530) );
  OAI221_X1 U11576 ( .B1(n10532), .B2(keyinput57), .C1(n10531), .C2(
        keyinput116), .A(n10530), .ZN(n10542) );
  XNOR2_X1 U11577 ( .A(n10533), .B(keyinput83), .ZN(n10534) );
  AOI21_X1 U11578 ( .B1(keyinput85), .B2(n5247), .A(n10534), .ZN(n10537) );
  XNOR2_X1 U11579 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput51), .ZN(n10536) );
  XNOR2_X1 U11580 ( .A(P1_REG2_REG_1__SCAN_IN), .B(keyinput63), .ZN(n10535) );
  NAND3_X1 U11581 ( .A1(n10537), .A2(n10536), .A3(n10535), .ZN(n10541) );
  XNOR2_X1 U11582 ( .A(keyinput91), .B(n9076), .ZN(n10540) );
  XNOR2_X1 U11583 ( .A(keyinput29), .B(n10538), .ZN(n10539) );
  NOR4_X1 U11584 ( .A1(n10542), .A2(n10541), .A3(n10540), .A4(n10539), .ZN(
        n10573) );
  AOI22_X1 U11585 ( .A1(n10545), .A2(keyinput64), .B1(keyinput45), .B2(n10544), 
        .ZN(n10543) );
  OAI221_X1 U11586 ( .B1(n10545), .B2(keyinput64), .C1(n10544), .C2(keyinput45), .A(n10543), .ZN(n10556) );
  AOI22_X1 U11587 ( .A1(n10548), .A2(keyinput119), .B1(n10547), .B2(keyinput37), .ZN(n10546) );
  OAI221_X1 U11588 ( .B1(n10548), .B2(keyinput119), .C1(n10547), .C2(
        keyinput37), .A(n10546), .ZN(n10555) );
  AOI22_X1 U11589 ( .A1(n10550), .A2(keyinput100), .B1(n6501), .B2(keyinput48), 
        .ZN(n10549) );
  OAI221_X1 U11590 ( .B1(n10550), .B2(keyinput100), .C1(n6501), .C2(keyinput48), .A(n10549), .ZN(n10554) );
  INV_X1 U11591 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n10552) );
  AOI22_X1 U11592 ( .A1(n6232), .A2(keyinput71), .B1(keyinput2), .B2(n10552), 
        .ZN(n10551) );
  OAI221_X1 U11593 ( .B1(n6232), .B2(keyinput71), .C1(n10552), .C2(keyinput2), 
        .A(n10551), .ZN(n10553) );
  NOR4_X1 U11594 ( .A1(n10556), .A2(n10555), .A3(n10554), .A4(n10553), .ZN(
        n10572) );
  AOI22_X1 U11595 ( .A1(n10559), .A2(keyinput94), .B1(keyinput7), .B2(n10558), 
        .ZN(n10557) );
  OAI221_X1 U11596 ( .B1(n10559), .B2(keyinput94), .C1(n10558), .C2(keyinput7), 
        .A(n10557), .ZN(n10570) );
  AOI22_X1 U11597 ( .A1(n10271), .A2(keyinput30), .B1(n10561), .B2(keyinput108), .ZN(n10560) );
  OAI221_X1 U11598 ( .B1(n10271), .B2(keyinput30), .C1(n10561), .C2(
        keyinput108), .A(n10560), .ZN(n10569) );
  AOI22_X1 U11599 ( .A1(n10564), .A2(keyinput56), .B1(keyinput19), .B2(n10563), 
        .ZN(n10562) );
  OAI221_X1 U11600 ( .B1(n10564), .B2(keyinput56), .C1(n10563), .C2(keyinput19), .A(n10562), .ZN(n10568) );
  AOI22_X1 U11601 ( .A1(n10566), .A2(keyinput3), .B1(n9692), .B2(keyinput104), 
        .ZN(n10565) );
  OAI221_X1 U11602 ( .B1(n10566), .B2(keyinput3), .C1(n9692), .C2(keyinput104), 
        .A(n10565), .ZN(n10567) );
  NOR4_X1 U11603 ( .A1(n10570), .A2(n10569), .A3(n10568), .A4(n10567), .ZN(
        n10571) );
  NAND4_X1 U11604 ( .A1(n10574), .A2(n10573), .A3(n10572), .A4(n10571), .ZN(
        n10575) );
  NOR4_X1 U11605 ( .A1(n10578), .A2(n10577), .A3(n10576), .A4(n10575), .ZN(
        n10579) );
  OAI21_X1 U11606 ( .B1(keyinput85), .B2(n10580), .A(n10579), .ZN(n10581) );
  XOR2_X1 U11607 ( .A(n10582), .B(n10581), .Z(P1_U3440) );
  XNOR2_X1 U11608 ( .A(n10584), .B(n10583), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11609 ( .A(n10586), .B(n10585), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11610 ( .A(n10588), .B(n10587), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11611 ( .A(n10590), .B(n10589), .ZN(ADD_1068_U48) );
  XNOR2_X1 U11612 ( .A(n10592), .B(n10591), .ZN(ADD_1068_U50) );
  XOR2_X1 U11613 ( .A(n10594), .B(n10593), .Z(ADD_1068_U54) );
  XOR2_X1 U11614 ( .A(n10596), .B(n10595), .Z(ADD_1068_U53) );
  XNOR2_X1 U11615 ( .A(n10598), .B(n10597), .ZN(ADD_1068_U52) );
  XNOR2_X1 U6729 ( .A(n5065), .B(P2_IR_REG_29__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U6779 ( .A1(n6593), .A2(n6592), .ZN(n6599) );
  CLKBUF_X1 U5086 ( .A(n5629), .Z(n10147) );
  CLKBUF_X2 U5008 ( .A(n6594), .Z(n9920) );
  NAND3_X1 U5108 ( .A1(n6599), .A2(n6908), .A3(n6600), .ZN(n6646) );
  NAND2_X1 U5358 ( .A1(n8240), .A2(n8110), .ZN(n6174) );
  CLKBUF_X1 U6423 ( .A(n6646), .Z(n6816) );
  NAND2_X2 U6780 ( .A1(n8240), .A2(n6175), .ZN(n7969) );
  CLKBUF_X1 U7976 ( .A(n6720), .Z(n5807) );
endmodule

