

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10060;

  AND2_X1 U4751 ( .A1(n5488), .A2(n5487), .ZN(n8158) );
  OAI211_X1 U4752 ( .C1(n5668), .C2(n9655), .A(n5743), .B(n5742), .ZN(n6892)
         );
  BUF_X2 U4753 ( .A(n4904), .Z(n7624) );
  CLKBUF_X2 U4755 ( .A(n4941), .Z(n6405) );
  INV_X2 U4756 ( .A(n4903), .ZN(n5548) );
  AND4_X1 U4757 ( .A1(n4877), .A2(n4878), .A3(n4876), .A4(n4875), .ZN(n6593)
         );
  AND2_X1 U4758 ( .A1(n5614), .A2(n7850), .ZN(n5711) );
  INV_X1 U4759 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4854) );
  NAND2_X1 U4760 ( .A1(n4680), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5627) );
  INV_X1 U4761 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9458) );
  INV_X1 U4762 ( .A(n5659), .ZN(n5621) );
  INV_X1 U4763 ( .A(n7850), .ZN(n5616) );
  INV_X1 U4764 ( .A(n8608), .ZN(n6018) );
  INV_X1 U4765 ( .A(n4904), .ZN(n5420) );
  NAND2_X1 U4766 ( .A1(n4880), .A2(n8594), .ZN(n4957) );
  NAND2_X1 U4767 ( .A1(n7655), .A2(n7653), .ZN(n8329) );
  INV_X1 U4768 ( .A(n6855), .ZN(n6240) );
  INV_X1 U4769 ( .A(n9713), .ZN(n9784) );
  OAI21_X1 U4770 ( .B1(n5304), .B2(n4567), .A(n4564), .ZN(n5339) );
  NAND2_X1 U4771 ( .A1(n4639), .A2(n4637), .ZN(n4641) );
  NAND4_X1 U4773 ( .A1(n5667), .A2(n5666), .A3(n5665), .A4(n5664), .ZN(n9755)
         );
  AOI21_X4 U4774 ( .B1(n4695), .B2(n4697), .A(n4295), .ZN(n4692) );
  XNOR2_X1 U4775 ( .A(n5582), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6205) );
  AOI211_X2 U4776 ( .C1(n9954), .C2(n8362), .A(n8361), .B(n8360), .ZN(n8363)
         );
  AOI21_X2 U4777 ( .B1(n6653), .B2(n6527), .A(n6652), .ZN(n6694) );
  XNOR2_X2 U4778 ( .A(n5358), .B(n5356), .ZN(n7916) );
  NAND2_X2 U4779 ( .A1(n4757), .A2(n4756), .ZN(n5358) );
  AOI21_X2 U4780 ( .B1(n7185), .B2(n7184), .A(n7183), .ZN(n7327) );
  INV_X4 U4781 ( .A(n5695), .ZN(n8605) );
  AND2_X2 U4782 ( .A1(n4831), .A2(n4829), .ZN(n4873) );
  XNOR2_X2 U4783 ( .A(n4846), .B(n4845), .ZN(n4866) );
  XNOR2_X2 U4784 ( .A(n5581), .B(n4369), .ZN(n5638) );
  INV_X1 U4785 ( .A(n4641), .ZN(n6246) );
  OR2_X1 U4786 ( .A1(n8530), .A2(n8528), .ZN(n4361) );
  NAND2_X1 U4787 ( .A1(n9051), .A2(n9058), .ZN(n9050) );
  NAND2_X1 U4788 ( .A1(n7914), .A2(n5359), .ZN(n5397) );
  AOI21_X1 U4789 ( .B1(n9066), .B2(n9727), .A(n9065), .ZN(n9309) );
  XNOR2_X1 U4790 ( .A(n9034), .B(n9033), .ZN(n9040) );
  AOI21_X1 U4791 ( .B1(n9091), .B2(n9727), .A(n4328), .ZN(n9319) );
  CLKBUF_X1 U4792 ( .A(n7859), .Z(n4341) );
  NAND2_X1 U4793 ( .A1(n8998), .A2(n8997), .ZN(n9095) );
  NAND2_X1 U4794 ( .A1(n4733), .A2(n4732), .ZN(n7862) );
  NAND2_X1 U4795 ( .A1(n9117), .A2(n9025), .ZN(n9103) );
  NAND2_X1 U4796 ( .A1(n4656), .A2(n4654), .ZN(n9154) );
  NOR2_X1 U4797 ( .A1(n8391), .A2(n4698), .ZN(n8250) );
  OAI21_X1 U4798 ( .B1(n4613), .B2(n4299), .A(n4348), .ZN(n5937) );
  AOI21_X1 U4799 ( .B1(n9078), .B2(n9739), .A(n9038), .ZN(n9039) );
  NAND2_X1 U4800 ( .A1(n4676), .A2(n4674), .ZN(n9212) );
  NAND2_X1 U4801 ( .A1(n5965), .A2(n5964), .ZN(n9511) );
  INV_X2 U4802 ( .A(n8336), .ZN(n4247) );
  OR2_X1 U4803 ( .A1(n5248), .A2(n5247), .ZN(n5268) );
  NAND2_X1 U4804 ( .A1(n6324), .A2(n6811), .ZN(n9749) );
  NAND2_X1 U4805 ( .A1(n4959), .A2(n4488), .ZN(n9953) );
  INV_X1 U4806 ( .A(n9945), .ZN(n6759) );
  INV_X1 U4807 ( .A(n9755), .ZN(n9725) );
  INV_X1 U4808 ( .A(n7960), .ZN(n8333) );
  NAND2_X1 U4809 ( .A1(n4867), .A2(n6719), .ZN(n4902) );
  INV_X2 U4810 ( .A(n6039), .ZN(n8600) );
  NAND4_X1 U4811 ( .A1(n4909), .A2(n4908), .A3(n4907), .A4(n4906), .ZN(n7960)
         );
  AND2_X2 U4812 ( .A1(n6448), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  INV_X1 U4813 ( .A(n6488), .ZN(n6343) );
  INV_X1 U4814 ( .A(n6708), .ZN(n4248) );
  AND2_X2 U4815 ( .A1(n5641), .A2(n6340), .ZN(n6855) );
  INV_X2 U4816 ( .A(n4957), .ZN(n7742) );
  BUF_X2 U4817 ( .A(n4958), .Z(n7616) );
  NAND2_X1 U4818 ( .A1(n5672), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U4819 ( .A1(n4258), .A2(n4277), .ZN(n6488) );
  INV_X1 U4820 ( .A(n5614), .ZN(n5615) );
  NAND2_X1 U4821 ( .A1(n4866), .A2(n7839), .ZN(n5543) );
  NAND2_X1 U4822 ( .A1(n6205), .A2(n8877), .ZN(n5640) );
  NAND2_X1 U4823 ( .A1(n5609), .A2(n5608), .ZN(n5614) );
  NAND2_X1 U4824 ( .A1(n5502), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U4825 ( .A1(n4853), .A2(n4852), .ZN(n7844) );
  XNOR2_X1 U4826 ( .A(n4841), .B(n4838), .ZN(n7827) );
  NAND2_X2 U4827 ( .A1(n6209), .A2(n6280), .ZN(n5668) );
  NAND2_X1 U4828 ( .A1(n4844), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4846) );
  OAI21_X1 U4829 ( .B1(n5580), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U4830 ( .A1(n8458), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4824) );
  NAND2_X1 U4831 ( .A1(n9545), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5613) );
  OAI21_X1 U4832 ( .B1(n5597), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U4833 ( .A1(n5627), .A2(n5604), .ZN(n5625) );
  OR2_X1 U4834 ( .A1(n4842), .A2(n4854), .ZN(n4847) );
  INV_X2 U4835 ( .A(n7567), .ZN(n4249) );
  NAND2_X2 U4836 ( .A1(n4817), .A2(n4731), .ZN(n4836) );
  NOR2_X1 U4837 ( .A1(n4682), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4681) );
  INV_X1 U4838 ( .A(n5756), .ZN(n5570) );
  NAND2_X1 U4839 ( .A1(n4716), .A2(n4715), .ZN(n4895) );
  AND2_X1 U4840 ( .A1(n5601), .A2(n4794), .ZN(n4793) );
  CLKBUF_X1 U4841 ( .A(n4859), .Z(n4860) );
  NOR2_X1 U4842 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5601) );
  INV_X1 U4843 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5586) );
  INV_X1 U4844 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5800) );
  INV_X1 U4845 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5565) );
  INV_X1 U4846 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5997) );
  INV_X2 U4847 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U4848 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n4811) );
  NOR2_X1 U4849 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n4812) );
  NOR2_X1 U4850 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5569) );
  INV_X1 U4851 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4720) );
  NOR2_X1 U4852 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5568) );
  NOR2_X1 U4853 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4859) );
  INV_X1 U4854 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5939) );
  OAI21_X2 U4855 ( .B1(n9247), .B2(n4770), .A(n4769), .ZN(n9219) );
  OAI22_X2 U4856 ( .A1(n9261), .A2(n8988), .B1(n9285), .B2(n9274), .ZN(n9247)
         );
  AOI21_X2 U4857 ( .B1(n7078), .B2(n7077), .A(n5104), .ZN(n7217) );
  AOI21_X2 U4858 ( .B1(n4750), .B2(n4748), .A(n4294), .ZN(n7078) );
  INV_X1 U4859 ( .A(n5489), .ZN(n4250) );
  INV_X2 U4860 ( .A(n5643), .ZN(n5635) );
  INV_X1 U4861 ( .A(n4957), .ZN(n4251) );
  INV_X1 U4862 ( .A(n5668), .ZN(n4252) );
  NAND2_X1 U4863 ( .A1(n7596), .A2(n8468), .ZN(n4904) );
  INV_X1 U4864 ( .A(n8992), .ZN(n4787) );
  OR2_X1 U4865 ( .A1(n5188), .A2(n5187), .ZN(n4547) );
  INV_X1 U4866 ( .A(n9882), .ZN(n7846) );
  NAND2_X1 U4867 ( .A1(n4560), .A2(n8830), .ZN(n4559) );
  NAND2_X1 U4868 ( .A1(n4563), .A2(n4561), .ZN(n4560) );
  OAI21_X1 U4869 ( .B1(n8834), .B2(n9299), .A(n8705), .ZN(n4563) );
  AND2_X1 U4870 ( .A1(n8711), .A2(n4562), .ZN(n4561) );
  OR2_X1 U4871 ( .A1(n6144), .A2(n8572), .ZN(n6211) );
  NAND2_X1 U4872 ( .A1(n5668), .A2(n7613), .ZN(n5695) );
  AND2_X1 U4873 ( .A1(n8630), .A2(n4335), .ZN(n4334) );
  OR2_X1 U4874 ( .A1(n4287), .A2(n8631), .ZN(n4335) );
  NAND2_X1 U4875 ( .A1(n8663), .A2(n8705), .ZN(n4339) );
  INV_X1 U4876 ( .A(n8664), .ZN(n4340) );
  NAND2_X1 U4877 ( .A1(n4464), .A2(n4461), .ZN(n7720) );
  NAND2_X1 U4878 ( .A1(n4466), .A2(n4465), .ZN(n4464) );
  NAND2_X1 U4879 ( .A1(n4462), .A2(n7754), .ZN(n4461) );
  NAND2_X1 U4880 ( .A1(n7714), .A2(n4283), .ZN(n4466) );
  AND2_X1 U4881 ( .A1(n7817), .A2(n8171), .ZN(n7820) );
  AOI21_X1 U4882 ( .B1(n5239), .B2(n4544), .A(n4543), .ZN(n4542) );
  INV_X1 U4883 ( .A(n5241), .ZN(n4543) );
  INV_X1 U4884 ( .A(n5213), .ZN(n4544) );
  INV_X1 U4885 ( .A(n5239), .ZN(n4545) );
  AOI21_X1 U4886 ( .B1(n4759), .B2(n4761), .A(n4315), .ZN(n4756) );
  NAND2_X1 U4887 ( .A1(n7859), .A2(n4759), .ZN(n4757) );
  OR2_X1 U4888 ( .A1(n6392), .A2(n6513), .ZN(n4888) );
  OR2_X1 U4889 ( .A1(n8346), .A2(n8134), .ZN(n7747) );
  OAI21_X1 U4890 ( .B1(n8156), .B2(n4288), .A(n4607), .ZN(n8114) );
  INV_X1 U4891 ( .A(n4608), .ZN(n4607) );
  OAI21_X1 U4892 ( .B1(n8137), .B2(n7825), .A(n7826), .ZN(n4608) );
  INV_X1 U4893 ( .A(n4378), .ZN(n4377) );
  OAI21_X1 U4894 ( .B1(n4713), .B2(n4379), .A(n8095), .ZN(n4378) );
  OR2_X1 U4895 ( .A1(n8093), .A2(n7926), .ZN(n7804) );
  OR2_X1 U4896 ( .A1(n8419), .A2(n7525), .ZN(n7704) );
  INV_X1 U4897 ( .A(n4396), .ZN(n4395) );
  OAI21_X1 U4898 ( .B1(n4398), .B2(n4397), .A(n4685), .ZN(n4396) );
  OR2_X1 U4899 ( .A1(n7488), .A2(n7517), .ZN(n7699) );
  XNOR2_X1 U4900 ( .A(n4370), .B(P2_IR_REG_28__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U4901 ( .A1(n8973), .A2(n8977), .ZN(n8873) );
  OR2_X1 U4902 ( .A1(n9321), .A2(n8999), .ZN(n9027) );
  INV_X1 U4903 ( .A(n9019), .ZN(n4659) );
  NAND2_X1 U4904 ( .A1(n6322), .A2(n6488), .ZN(n6325) );
  OAI21_X1 U4905 ( .B1(n7741), .B2(n7604), .A(n7606), .ZN(n7610) );
  INV_X1 U4906 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5572) );
  NOR2_X1 U4907 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4353) );
  NAND2_X1 U4908 ( .A1(n5161), .A2(n5160), .ZN(n5188) );
  AOI21_X1 U4909 ( .B1(n4551), .B2(n4273), .A(n4550), .ZN(n4549) );
  INV_X1 U4910 ( .A(n4552), .ZN(n4551) );
  OAI21_X1 U4911 ( .B1(n4555), .B2(n4273), .A(n5135), .ZN(n4552) );
  NOR2_X1 U4912 ( .A1(n5013), .A2(n5012), .ZN(n4754) );
  AND4_X1 U4913 ( .A1(n4927), .A2(n4926), .A3(n4925), .A4(n4924), .ZN(n9862)
         );
  OR2_X1 U4914 ( .A1(n5419), .A2(n6757), .ZN(n4924) );
  NAND2_X1 U4915 ( .A1(n8111), .A2(n8176), .ZN(n8112) );
  OR2_X1 U4916 ( .A1(n5417), .A2(n5416), .ZN(n5436) );
  OR2_X1 U4917 ( .A1(n8366), .A2(n8210), .ZN(n8171) );
  AOI21_X1 U4918 ( .B1(n8250), .B2(n4383), .A(n4381), .ZN(n4380) );
  NAND2_X1 U4919 ( .A1(n4382), .A2(n8104), .ZN(n4381) );
  NAND2_X1 U4920 ( .A1(n4383), .A2(n4385), .ZN(n4382) );
  INV_X1 U4921 ( .A(n8102), .ZN(n8269) );
  AND3_X1 U4922 ( .A1(n5294), .A2(n5293), .A3(n5292), .ZN(n8268) );
  NOR2_X1 U4923 ( .A1(n7766), .A2(n7765), .ZN(n8279) );
  OR2_X1 U4924 ( .A1(n7450), .A2(n7686), .ZN(n4687) );
  OR2_X1 U4925 ( .A1(n5049), .A2(n5048), .ZN(n5073) );
  OR2_X1 U4926 ( .A1(n4404), .A2(n4400), .ZN(n4403) );
  NAND2_X1 U4927 ( .A1(n6911), .A2(n4406), .ZN(n4405) );
  NOR2_X1 U4928 ( .A1(n4407), .A2(n6945), .ZN(n4406) );
  INV_X1 U4929 ( .A(n6910), .ZN(n4407) );
  AND2_X1 U4930 ( .A1(n7797), .A2(n7841), .ZN(n8292) );
  INV_X1 U4931 ( .A(n8312), .ZN(n9863) );
  AND2_X1 U4932 ( .A1(n4880), .A2(n7613), .ZN(n4958) );
  NAND2_X1 U4933 ( .A1(n6532), .A2(n6560), .ZN(n9861) );
  NAND2_X2 U4934 ( .A1(n7844), .A2(n5556), .ZN(n4880) );
  AND2_X1 U4935 ( .A1(n5527), .A2(n9915), .ZN(n7063) );
  AND2_X1 U4936 ( .A1(n7761), .A2(n4866), .ZN(n9946) );
  NAND2_X1 U4937 ( .A1(n5525), .A2(n9917), .ZN(n7061) );
  INV_X1 U4938 ( .A(n4624), .ZN(n4623) );
  OAI21_X1 U4939 ( .B1(n4627), .B2(n4625), .A(n6102), .ZN(n4624) );
  INV_X1 U4940 ( .A(n4629), .ZN(n4625) );
  NAND2_X1 U4941 ( .A1(n5679), .A2(n5678), .ZN(n5681) );
  OR2_X1 U4942 ( .A1(n9001), .A2(n8693), .ZN(n9089) );
  OR2_X1 U4943 ( .A1(n9114), .A2(n8996), .ZN(n4798) );
  INV_X1 U4944 ( .A(n4786), .ZN(n4785) );
  OAI21_X1 U4945 ( .B1(n8991), .B2(n4787), .A(n4285), .ZN(n4786) );
  NAND2_X1 U4946 ( .A1(n6864), .A2(n6854), .ZN(n7001) );
  OR2_X1 U4947 ( .A1(n5639), .A2(n9744), .ZN(n5641) );
  NAND2_X1 U4948 ( .A1(n6886), .A2(n4766), .ZN(n6864) );
  NOR2_X1 U4949 ( .A1(n8729), .A2(n4767), .ZN(n4766) );
  INV_X1 U4950 ( .A(n6853), .ZN(n4767) );
  INV_X1 U4951 ( .A(n9751), .ZN(n9727) );
  NAND2_X1 U4952 ( .A1(n6143), .A2(n6142), .ZN(n9316) );
  AND3_X1 U4953 ( .A1(n6187), .A2(n6185), .A3(n6184), .ZN(n9764) );
  AOI21_X1 U4954 ( .B1(n5580), .B2(P1_IR_REG_31__SCAN_IN), .A(n4366), .ZN(
        n4365) );
  NAND2_X1 U4955 ( .A1(n4367), .A2(n5586), .ZN(n4366) );
  NAND2_X1 U4956 ( .A1(n4368), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4367) );
  NAND2_X1 U4957 ( .A1(n5541), .A2(n8272), .ZN(n7929) );
  INV_X1 U4958 ( .A(n9120), .ZN(n8999) );
  NAND2_X1 U4959 ( .A1(n6171), .A2(n6170), .ZN(n9090) );
  AND2_X1 U4960 ( .A1(n8965), .A2(n6285), .ZN(n9707) );
  NAND2_X1 U4961 ( .A1(n8598), .A2(n8597), .ZN(n9585) );
  AND2_X1 U4962 ( .A1(n7663), .A2(n4400), .ZN(n4458) );
  NAND2_X1 U4963 ( .A1(n4336), .A2(n4334), .ZN(n8632) );
  OR2_X1 U4964 ( .A1(n7691), .A2(n7690), .ZN(n4492) );
  NAND2_X1 U4965 ( .A1(n4452), .A2(n4451), .ZN(n7715) );
  NOR2_X1 U4966 ( .A1(n7712), .A2(n7806), .ZN(n4451) );
  MUX2_X1 U4967 ( .A(n8673), .B(n8672), .S(n8705), .Z(n8674) );
  NOR2_X1 U4968 ( .A1(n8104), .A2(n7719), .ZN(n7724) );
  NAND2_X1 U4969 ( .A1(n4460), .A2(n4459), .ZN(n7718) );
  AND2_X1 U4970 ( .A1(n7814), .A2(n7764), .ZN(n4459) );
  INV_X1 U4971 ( .A(n4793), .ZN(n4682) );
  INV_X1 U4972 ( .A(n4760), .ZN(n4759) );
  OAI21_X1 U4973 ( .B1(n4278), .B2(n4761), .A(n7869), .ZN(n4760) );
  OR2_X1 U4974 ( .A1(n7424), .A2(n4636), .ZN(n4635) );
  INV_X1 U4975 ( .A(n5899), .ZN(n4636) );
  INV_X1 U4976 ( .A(n5874), .ZN(n4350) );
  INV_X1 U4977 ( .A(n5980), .ZN(n4347) );
  NOR2_X1 U4978 ( .A1(n4775), .A2(n4772), .ZN(n4771) );
  NOR2_X1 U4979 ( .A1(n9504), .A2(n9214), .ZN(n4775) );
  NOR2_X1 U4980 ( .A1(n9249), .A2(n4773), .ZN(n4772) );
  AND2_X1 U4981 ( .A1(n4569), .A2(n5320), .ZN(n4568) );
  NAND2_X1 U4982 ( .A1(n5303), .A2(n5305), .ZN(n4569) );
  NAND2_X1 U4983 ( .A1(n5139), .A2(n5138), .ZN(n5160) );
  INV_X1 U4984 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4718) );
  INV_X1 U4985 ( .A(n7861), .ZN(n5300) );
  AND2_X1 U4986 ( .A1(n9922), .A2(n7827), .ZN(n4865) );
  NOR2_X1 U4987 ( .A1(n4477), .A2(n4474), .ZN(n4473) );
  INV_X1 U4988 ( .A(n7748), .ZN(n4474) );
  AOI21_X1 U4989 ( .B1(n4479), .B2(n4481), .A(n4478), .ZN(n4477) );
  NOR2_X1 U4990 ( .A1(n4253), .A2(n4484), .ZN(n4478) );
  NAND2_X1 U4991 ( .A1(n4303), .A2(n7748), .ZN(n4476) );
  OR2_X1 U4992 ( .A1(n8350), .A2(n8158), .ZN(n7826) );
  NOR2_X1 U4993 ( .A1(n7821), .A2(n8170), .ZN(n4799) );
  OR2_X1 U4994 ( .A1(n8371), .A2(n7946), .ZN(n8169) );
  OR2_X1 U4995 ( .A1(n8380), .A2(n7872), .ZN(n7814) );
  NAND2_X1 U4996 ( .A1(n8298), .A2(n8308), .ZN(n4414) );
  OR2_X1 U4997 ( .A1(n4414), .A2(n8276), .ZN(n4413) );
  NOR2_X1 U4998 ( .A1(n7787), .A2(n4714), .ZN(n4713) );
  NOR2_X1 U4999 ( .A1(n4424), .A2(n8419), .ZN(n4423) );
  INV_X1 U5000 ( .A(n4425), .ZN(n4424) );
  NOR2_X1 U5001 ( .A1(n7488), .A2(n8424), .ZN(n4425) );
  AOI21_X1 U5002 ( .B1(n4603), .B2(n4601), .A(n4301), .ZN(n4600) );
  INV_X1 U5003 ( .A(n7676), .ZN(n4601) );
  INV_X1 U5004 ( .A(n4603), .ZN(n4602) );
  AND2_X1 U5005 ( .A1(n7778), .A2(n7671), .ZN(n4603) );
  NOR2_X1 U5006 ( .A1(n8434), .A2(n4418), .ZN(n4417) );
  INV_X1 U5007 ( .A(n4419), .ZN(n4418) );
  INV_X1 U5008 ( .A(n7662), .ZN(n4581) );
  OAI21_X1 U5009 ( .B1(n7774), .B2(n4579), .A(n7666), .ZN(n4578) );
  NAND2_X1 U5010 ( .A1(n7773), .A2(n7662), .ZN(n4579) );
  NAND2_X1 U5011 ( .A1(n6758), .A2(n9953), .ZN(n7641) );
  INV_X1 U5012 ( .A(n6363), .ZN(n4389) );
  INV_X1 U5013 ( .A(n8330), .ZN(n6729) );
  INV_X1 U5014 ( .A(n4430), .ZN(n4428) );
  NAND2_X1 U5015 ( .A1(n8332), .A2(n7653), .ZN(n9858) );
  NOR2_X1 U5016 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n4731) );
  AND4_X1 U5017 ( .A1(n4814), .A2(n4813), .A3(n4812), .A4(n4811), .ZN(n4815)
         );
  NOR2_X1 U5018 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n4814) );
  NOR2_X1 U5019 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4813) );
  NAND2_X1 U5020 ( .A1(n8550), .A2(n6086), .ZN(n4629) );
  NOR2_X1 U5021 ( .A1(n7501), .A2(n7500), .ZN(n7544) );
  NAND2_X1 U5022 ( .A1(n4513), .A2(n9075), .ZN(n4512) );
  NAND2_X1 U5023 ( .A1(n4673), .A2(n4670), .ZN(n4664) );
  NAND2_X1 U5024 ( .A1(n4673), .A2(n4663), .ZN(n4662) );
  OR2_X1 U5025 ( .A1(n9161), .A2(n9018), .ZN(n4658) );
  AND2_X1 U5026 ( .A1(n8648), .A2(n8788), .ZN(n8988) );
  AND2_X1 U5027 ( .A1(n9521), .A2(n9266), .ZN(n8986) );
  NAND2_X1 U5028 ( .A1(n6819), .A2(n8842), .ZN(n6327) );
  NAND2_X1 U5029 ( .A1(n9752), .A2(n9738), .ZN(n9737) );
  XNOR2_X1 U5030 ( .A(n7610), .B(n7609), .ZN(n7607) );
  NAND2_X1 U5031 ( .A1(n7602), .A2(n7601), .ZN(n7741) );
  OAI21_X1 U5032 ( .B1(n5373), .B2(n4312), .A(n4570), .ZN(n5450) );
  INV_X1 U5033 ( .A(n4571), .ZN(n4570) );
  OAI21_X1 U5034 ( .B1(n4574), .B2(n4312), .A(n5430), .ZN(n4571) );
  OAI21_X1 U5035 ( .B1(n5339), .B2(n5338), .A(n5337), .ZN(n5362) );
  AOI21_X1 U5036 ( .B1(n4568), .B2(n4566), .A(n4565), .ZN(n4564) );
  INV_X1 U5037 ( .A(n4568), .ZN(n4567) );
  INV_X1 U5038 ( .A(n5322), .ZN(n4565) );
  OAI21_X1 U5039 ( .B1(n5262), .B2(n5261), .A(n5260), .ZN(n5279) );
  AND2_X1 U5040 ( .A1(n5241), .A2(n5219), .ZN(n5239) );
  NAND2_X1 U5041 ( .A1(n4541), .A2(n5186), .ZN(n4540) );
  INV_X1 U5042 ( .A(n5214), .ZN(n4541) );
  INV_X1 U5043 ( .A(n5108), .ZN(n4553) );
  NOR2_X1 U5044 ( .A1(n5109), .A2(n4556), .ZN(n4555) );
  INV_X1 U5045 ( .A(n5087), .ZN(n4556) );
  NAND2_X1 U5046 ( .A1(n4533), .A2(n4290), .ZN(n5086) );
  NAND2_X1 U5047 ( .A1(n4806), .A2(n4532), .ZN(n4531) );
  INV_X1 U5048 ( .A(n5036), .ZN(n4534) );
  INV_X1 U5049 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U5050 ( .A1(n4975), .A2(n4974), .ZN(n4995) );
  NAND2_X1 U5051 ( .A1(n4857), .A2(SI_0_), .ZN(n4891) );
  INV_X1 U5052 ( .A(n4736), .ZN(n4735) );
  OAI21_X1 U5053 ( .B1(n4738), .B2(n4737), .A(n7923), .ZN(n4736) );
  INV_X1 U5054 ( .A(n5256), .ZN(n4737) );
  NAND2_X1 U5055 ( .A1(n5395), .A2(n5394), .ZN(n5396) );
  NOR2_X1 U5056 ( .A1(n4746), .A2(n4264), .ZN(n4745) );
  NAND2_X1 U5057 ( .A1(n5224), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5248) );
  INV_X1 U5058 ( .A(n5225), .ZN(n5224) );
  NAND2_X1 U5059 ( .A1(n5378), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5417) );
  AND2_X1 U5060 ( .A1(n4753), .A2(n5034), .ZN(n4752) );
  NAND2_X1 U5061 ( .A1(n6833), .A2(n4754), .ZN(n4753) );
  INV_X1 U5062 ( .A(n4752), .ZN(n4749) );
  NAND2_X1 U5063 ( .A1(n4747), .A2(n4281), .ZN(n4750) );
  INV_X1 U5064 ( .A(n6771), .ZN(n4755) );
  XNOR2_X1 U5065 ( .A(n9937), .B(n4902), .ZN(n4727) );
  NOR2_X1 U5066 ( .A1(n7887), .A2(n4739), .ZN(n4738) );
  INV_X1 U5067 ( .A(n5238), .ZN(n4739) );
  OR2_X1 U5068 ( .A1(n5255), .A2(n5254), .ZN(n5256) );
  NAND2_X1 U5069 ( .A1(n4947), .A2(n4946), .ZN(n6753) );
  NAND2_X1 U5070 ( .A1(n4740), .A2(n4741), .ZN(n6736) );
  AND2_X1 U5071 ( .A1(n4991), .A2(n4744), .ZN(n4740) );
  INV_X1 U5072 ( .A(n6739), .ZN(n4991) );
  NOR2_X1 U5073 ( .A1(n5542), .A2(n9882), .ZN(n5555) );
  INV_X1 U5074 ( .A(n7827), .ZN(n7799) );
  AOI21_X1 U5075 ( .B1(n7835), .B2(n7834), .A(n7833), .ZN(n7838) );
  NOR2_X1 U5076 ( .A1(n7832), .A2(n7831), .ZN(n7833) );
  INV_X1 U5077 ( .A(n6392), .ZN(n7621) );
  AND4_X1 U5078 ( .A1(n5230), .A2(n5229), .A3(n5228), .A4(n5227), .ZN(n7573)
         );
  AND4_X1 U5079 ( .A1(n5030), .A2(n5029), .A3(n5028), .A4(n5027), .ZN(n7157)
         );
  AND4_X1 U5080 ( .A1(n4988), .A2(n4987), .A3(n4986), .A4(n4985), .ZN(n6949)
         );
  OR2_X1 U5081 ( .A1(n5419), .A2(n9394), .ZN(n4796) );
  AND2_X1 U5082 ( .A1(n5533), .A2(n7799), .ZN(n6532) );
  NAND2_X1 U5083 ( .A1(n8177), .A2(n8111), .ZN(n8149) );
  OR2_X1 U5084 ( .A1(n8366), .A2(n8106), .ZN(n8107) );
  AND2_X1 U5085 ( .A1(n5425), .A2(n5424), .ZN(n8210) );
  NAND2_X1 U5086 ( .A1(n4280), .A2(n4386), .ZN(n4385) );
  INV_X1 U5087 ( .A(n8103), .ZN(n4386) );
  NAND2_X1 U5088 ( .A1(n4384), .A2(n4280), .ZN(n4383) );
  NAND2_X1 U5089 ( .A1(n4387), .A2(n4257), .ZN(n4384) );
  INV_X1 U5090 ( .A(n4595), .ZN(n4594) );
  AND2_X1 U5091 ( .A1(n8276), .A2(n8260), .ZN(n4698) );
  OR2_X1 U5092 ( .A1(n8399), .A2(n8314), .ZN(n8101) );
  NOR2_X1 U5093 ( .A1(n4413), .A2(n8303), .ZN(n8271) );
  NOR2_X1 U5094 ( .A1(n8099), .A2(n8402), .ZN(n8098) );
  OR2_X1 U5095 ( .A1(n7528), .A2(n4379), .ZN(n4374) );
  OR2_X1 U5096 ( .A1(n8419), .A2(n7949), .ZN(n7527) );
  AOI21_X1 U5097 ( .B1(n7786), .B2(n4587), .A(n4586), .ZN(n4585) );
  INV_X1 U5098 ( .A(n7699), .ZN(n4587) );
  NAND2_X1 U5099 ( .A1(n7484), .A2(n7699), .ZN(n7485) );
  NAND2_X1 U5100 ( .A1(n4393), .A2(n4392), .ZN(n7489) );
  AOI21_X1 U5101 ( .B1(n4395), .B2(n4397), .A(n4265), .ZN(n4392) );
  AND2_X1 U5102 ( .A1(n7451), .A2(n4686), .ZN(n4685) );
  OR2_X1 U5103 ( .A1(n7449), .A2(n7952), .ZN(n4686) );
  AND2_X1 U5104 ( .A1(n7688), .A2(n7683), .ZN(n7686) );
  NAND2_X1 U5105 ( .A1(n7200), .A2(n4398), .ZN(n4394) );
  AND2_X1 U5106 ( .A1(n7349), .A2(n4705), .ZN(n7369) );
  OR2_X1 U5107 ( .A1(n9976), .A2(n7203), .ZN(n7675) );
  NAND2_X1 U5108 ( .A1(n7199), .A2(n7676), .ZN(n4604) );
  NAND2_X1 U5109 ( .A1(n4604), .A2(n4603), .ZN(n7366) );
  INV_X1 U5110 ( .A(n9861), .ZN(n8313) );
  INV_X1 U5111 ( .A(n7776), .ZN(n6962) );
  AND2_X1 U5112 ( .A1(n7668), .A2(n7669), .ZN(n7776) );
  AND4_X1 U5113 ( .A1(n5055), .A2(n5054), .A3(n5053), .A4(n5052), .ZN(n7162)
         );
  NAND2_X1 U5114 ( .A1(n4980), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5004) );
  NAND2_X1 U5115 ( .A1(n6900), .A2(n6912), .ZN(n6947) );
  AND4_X1 U5116 ( .A1(n5009), .A2(n5008), .A3(n5007), .A4(n5006), .ZN(n6970)
         );
  NOR2_X1 U5117 ( .A1(n6723), .A2(n9953), .ZN(n6905) );
  NAND2_X1 U5118 ( .A1(n6713), .A2(n6712), .ZN(n6911) );
  NAND2_X1 U5119 ( .A1(n6744), .A2(n6745), .ZN(n6713) );
  AND2_X1 U5120 ( .A1(n7639), .A2(n7634), .ZN(n9857) );
  NAND2_X1 U5121 ( .A1(n6593), .A2(n6917), .ZN(n6918) );
  NOR2_X1 U5122 ( .A1(n6584), .A2(n6917), .ZN(n8326) );
  AND2_X1 U5123 ( .A1(n8346), .A2(n9954), .ZN(n4605) );
  INV_X1 U5124 ( .A(n9954), .ZN(n9983) );
  AND2_X1 U5125 ( .A1(n7065), .A2(n6716), .ZN(n7051) );
  AND2_X1 U5126 ( .A1(n5521), .A2(n5520), .ZN(n9883) );
  INV_X1 U5127 ( .A(n5505), .ZN(n4848) );
  AND2_X1 U5128 ( .A1(n4823), .A2(n4856), .ZN(n4610) );
  NAND2_X1 U5129 ( .A1(n5514), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U5130 ( .A1(n8899), .A2(n5621), .ZN(n5703) );
  NOR2_X1 U5131 ( .A1(n8503), .A2(n4359), .ZN(n4358) );
  INV_X1 U5132 ( .A(n4363), .ZN(n4359) );
  NAND2_X1 U5133 ( .A1(n8513), .A2(n5980), .ZN(n4633) );
  OR2_X1 U5134 ( .A1(n8510), .A2(n8513), .ZN(n8511) );
  OR2_X1 U5135 ( .A1(n6035), .A2(n8541), .ZN(n6055) );
  NAND2_X1 U5136 ( .A1(n5639), .A2(n8875), .ZN(n5600) );
  INV_X1 U5137 ( .A(n8830), .ZN(n4558) );
  NAND2_X1 U5138 ( .A1(n8873), .A2(n8604), .ZN(n8834) );
  INV_X1 U5139 ( .A(n5685), .ZN(n6039) );
  NAND2_X1 U5140 ( .A1(n8903), .A2(n4444), .ZN(n6453) );
  OR2_X1 U5141 ( .A1(n6351), .A2(n6277), .ZN(n4444) );
  NAND2_X1 U5142 ( .A1(n6494), .A2(n6493), .ZN(n6935) );
  OR2_X1 U5143 ( .A1(n8929), .A2(n8930), .ZN(n4441) );
  AND2_X1 U5144 ( .A1(n4441), .A2(n4440), .ZN(n6937) );
  NAND2_X1 U5145 ( .A1(n8934), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4440) );
  OR2_X1 U5146 ( .A1(n6937), .A2(n6938), .ZN(n4439) );
  XNOR2_X1 U5147 ( .A(n7544), .B(n7550), .ZN(n7503) );
  AND2_X1 U5148 ( .A1(n9002), .A2(n9000), .ZN(n4777) );
  OR2_X1 U5149 ( .A1(n9473), .A2(n9144), .ZN(n9136) );
  OR2_X1 U5150 ( .A1(n9473), .A2(n9157), .ZN(n9115) );
  NOR2_X1 U5151 ( .A1(n9163), .A2(n4289), .ZN(n4657) );
  OR2_X1 U5152 ( .A1(n9204), .A2(n4658), .ZN(n4653) );
  AND2_X1 U5153 ( .A1(n4660), .A2(n4659), .ZN(n9166) );
  AOI21_X1 U5154 ( .B1(n4785), .B2(n4787), .A(n4302), .ZN(n4784) );
  OR2_X1 U5155 ( .A1(n9204), .A2(n9018), .ZN(n4660) );
  NAND2_X1 U5156 ( .A1(n6003), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6023) );
  INV_X1 U5157 ( .A(n6005), .ZN(n6003) );
  INV_X1 U5158 ( .A(n9194), .ZN(n8991) );
  AOI21_X1 U5159 ( .B1(n9212), .B2(n9017), .A(n9016), .ZN(n9205) );
  AND2_X1 U5160 ( .A1(n9499), .A2(n9242), .ZN(n8990) );
  NAND2_X1 U5161 ( .A1(n9191), .A2(n8991), .ZN(n9192) );
  OR2_X1 U5162 ( .A1(n9262), .A2(n9012), .ZN(n4679) );
  AND2_X1 U5163 ( .A1(n8640), .A2(n8811), .ZN(n8738) );
  NAND2_X1 U5164 ( .A1(n9603), .A2(n7418), .ZN(n4780) );
  NAND2_X1 U5165 ( .A1(n4768), .A2(n6852), .ZN(n6886) );
  OR2_X1 U5166 ( .A1(n8718), .A2(n6443), .ZN(n9723) );
  INV_X1 U5167 ( .A(n9723), .ZN(n9756) );
  NAND2_X1 U5168 ( .A1(n6165), .A2(n6164), .ZN(n9311) );
  NAND2_X1 U5169 ( .A1(n5880), .A2(n5879), .ZN(n9597) );
  INV_X1 U5170 ( .A(n9817), .ZN(n9598) );
  INV_X1 U5171 ( .A(n9742), .ZN(n9819) );
  OR2_X1 U5172 ( .A1(n6469), .A2(n8875), .ZN(n9817) );
  AND2_X1 U5173 ( .A1(n6465), .A2(n6464), .ZN(n6473) );
  NAND2_X1 U5174 ( .A1(n6272), .A2(n6204), .ZN(n9765) );
  NOR2_X1 U5175 ( .A1(n4791), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4790) );
  NAND2_X1 U5176 ( .A1(n4793), .A2(n4792), .ZN(n4791) );
  INV_X1 U5177 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4792) );
  INV_X1 U5178 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5626) );
  NOR2_X1 U5179 ( .A1(n9544), .A2(n5610), .ZN(n5602) );
  INV_X1 U5180 ( .A(n5625), .ZN(n5607) );
  NAND2_X1 U5181 ( .A1(n5476), .A2(n5475), .ZN(n7598) );
  NAND2_X1 U5182 ( .A1(n5474), .A2(n5473), .ZN(n5476) );
  XNOR2_X1 U5183 ( .A(n5595), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U5184 ( .A1(n4573), .A2(n5406), .ZN(n5429) );
  NAND2_X1 U5185 ( .A1(n5373), .A2(n4574), .ZN(n4573) );
  OAI21_X1 U5186 ( .B1(n5362), .B2(n5361), .A(n5360), .ZN(n5371) );
  AND2_X1 U5187 ( .A1(n5372), .A2(n5367), .ZN(n5370) );
  NOR2_X1 U5188 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5574) );
  NAND2_X1 U5189 ( .A1(n4547), .A2(n5186), .ZN(n5215) );
  XNOR2_X1 U5190 ( .A(n5110), .B(n5105), .ZN(n6389) );
  NAND2_X1 U5191 ( .A1(n5088), .A2(n5087), .ZN(n5110) );
  XNOR2_X1 U5192 ( .A(n4912), .B(n4896), .ZN(n4910) );
  AND2_X1 U5193 ( .A1(n5530), .A2(n5529), .ZN(n6530) );
  INV_X1 U5194 ( .A(n4754), .ZN(n4751) );
  NAND2_X1 U5195 ( .A1(n6753), .A2(n4742), .ZN(n4741) );
  NOR2_X1 U5196 ( .A1(n6637), .A2(n4743), .ZN(n4742) );
  INV_X1 U5197 ( .A(n4948), .ZN(n4743) );
  NAND2_X1 U5198 ( .A1(n4968), .A2(n4969), .ZN(n4744) );
  INV_X1 U5199 ( .A(n7848), .ZN(n4469) );
  AND2_X1 U5200 ( .A1(n4880), .A2(n7844), .ZN(n6557) );
  NAND2_X1 U5201 ( .A1(n7618), .A2(n7617), .ZN(n8340) );
  AOI21_X1 U5202 ( .B1(n4256), .B2(n4691), .A(n4318), .ZN(n4689) );
  OAI21_X1 U5203 ( .B1(n8122), .B2(n8292), .A(n8121), .ZN(n4606) );
  NOR2_X1 U5204 ( .A1(n8118), .A2(n8117), .ZN(n8122) );
  OAI21_X1 U5205 ( .B1(n8138), .B2(n8137), .A(n4372), .ZN(n8349) );
  OAI21_X1 U5206 ( .B1(n8147), .B2(n4691), .A(n4256), .ZN(n4372) );
  NAND2_X1 U5207 ( .A1(n8146), .A2(n8112), .ZN(n8138) );
  NAND2_X1 U5208 ( .A1(n8287), .A2(n7808), .ZN(n8266) );
  NAND2_X1 U5209 ( .A1(n8336), .A2(n6724), .ZN(n8307) );
  NAND2_X1 U5210 ( .A1(n7846), .A2(n5540), .ZN(n8272) );
  NAND2_X1 U5211 ( .A1(n6020), .A2(n6019), .ZN(n9493) );
  NOR2_X1 U5212 ( .A1(n4642), .A2(n4638), .ZN(n4637) );
  OR2_X1 U5213 ( .A1(n6179), .A2(n6178), .ZN(n4642) );
  OAI22_X1 U5214 ( .A1(n6354), .A2(n8594), .B1(n5653), .B2(n7613), .ZN(n4789)
         );
  NAND2_X1 U5215 ( .A1(n4618), .A2(n4615), .ZN(n8496) );
  AND2_X1 U5216 ( .A1(n4616), .A2(n8538), .ZN(n4615) );
  NAND2_X1 U5217 ( .A1(n8537), .A2(n4617), .ZN(n4616) );
  INV_X1 U5218 ( .A(n8891), .ZN(n7418) );
  INV_X1 U5219 ( .A(n8888), .ZN(n9285) );
  NAND2_X1 U5220 ( .A1(n6034), .A2(n6033), .ZN(n9487) );
  AND3_X1 U5221 ( .A1(n6232), .A2(n9817), .A3(n8718), .ZN(n8571) );
  AND2_X1 U5222 ( .A1(n6211), .A2(n6145), .ZN(n9085) );
  AND2_X1 U5223 ( .A1(n9222), .A2(n6233), .ZN(n8578) );
  OAI21_X1 U5224 ( .B1(n8968), .B2(n4322), .A(n4448), .ZN(n4447) );
  AOI21_X1 U5225 ( .B1(n8969), .B2(n9707), .A(n9699), .ZN(n4448) );
  AND2_X1 U5226 ( .A1(n5668), .A2(n4527), .ZN(n4526) );
  NAND2_X1 U5227 ( .A1(n8594), .A2(n4528), .ZN(n4527) );
  NAND2_X1 U5228 ( .A1(n4505), .A2(n9585), .ZN(n4504) );
  OR2_X1 U5229 ( .A1(n9084), .A2(n4509), .ZN(n4508) );
  AOI21_X1 U5230 ( .B1(n9079), .B2(n9727), .A(n4325), .ZN(n9314) );
  NAND2_X1 U5231 ( .A1(n4327), .A2(n4326), .ZN(n4325) );
  NAND2_X1 U5232 ( .A1(n9105), .A2(n9739), .ZN(n4326) );
  INV_X1 U5233 ( .A(n9311), .ZN(n9075) );
  NAND2_X1 U5234 ( .A1(n4330), .A2(n4329), .ZN(n4328) );
  NAND2_X1 U5235 ( .A1(n9120), .A2(n9739), .ZN(n4329) );
  NAND2_X1 U5236 ( .A1(n4778), .A2(n9000), .ZN(n9083) );
  NAND2_X1 U5237 ( .A1(n9762), .A2(n6857), .ZN(n9297) );
  INV_X1 U5238 ( .A(n9042), .ZN(n9718) );
  INV_X1 U5239 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9544) );
  MUX2_X1 U5240 ( .A(n7635), .B(n7631), .S(n7754), .Z(n7648) );
  NAND2_X1 U5241 ( .A1(n8614), .A2(n4337), .ZN(n4336) );
  NOR2_X1 U5242 ( .A1(n4287), .A2(n4338), .ZN(n4337) );
  NAND2_X1 U5243 ( .A1(n8798), .A2(n8805), .ZN(n4338) );
  AND2_X1 U5244 ( .A1(n8652), .A2(n9009), .ZN(n4333) );
  OAI21_X1 U5245 ( .B1(n4457), .B2(n4456), .A(n7674), .ZN(n7687) );
  NAND2_X1 U5246 ( .A1(n7670), .A2(n7671), .ZN(n4456) );
  AOI21_X1 U5247 ( .B1(n7664), .B2(n4458), .A(n4300), .ZN(n4457) );
  NAND2_X1 U5248 ( .A1(n4490), .A2(n7698), .ZN(n7703) );
  OAI211_X1 U5249 ( .C1(n7692), .C2(n7754), .A(n4491), .B(n7784), .ZN(n4490)
         );
  NOR2_X1 U5250 ( .A1(n4454), .A2(n7789), .ZN(n4453) );
  INV_X1 U5251 ( .A(n7709), .ZN(n4454) );
  NAND2_X1 U5252 ( .A1(n7717), .A2(n4463), .ZN(n4462) );
  AND2_X1 U5253 ( .A1(n7809), .A2(n7767), .ZN(n4463) );
  NAND2_X1 U5254 ( .A1(n7720), .A2(n4284), .ZN(n4460) );
  NAND2_X1 U5255 ( .A1(n7725), .A2(n4465), .ZN(n4501) );
  INV_X1 U5256 ( .A(n4498), .ZN(n4497) );
  OAI21_X1 U5257 ( .B1(n7724), .B2(n4499), .A(n7723), .ZN(n4498) );
  NAND2_X1 U5258 ( .A1(n8206), .A2(n4500), .ZN(n4499) );
  NAND2_X1 U5259 ( .A1(n8105), .A2(n7947), .ZN(n4500) );
  NAND2_X1 U5260 ( .A1(n7727), .A2(n4465), .ZN(n4494) );
  INV_X1 U5261 ( .A(n4763), .ZN(n4761) );
  NAND2_X1 U5262 ( .A1(n4486), .A2(n4465), .ZN(n4485) );
  AOI21_X1 U5263 ( .B1(n4480), .B2(n4482), .A(n4254), .ZN(n4479) );
  AOI21_X1 U5264 ( .B1(n4496), .B2(n4495), .A(n4493), .ZN(n7734) );
  NAND2_X1 U5265 ( .A1(n7726), .A2(n4465), .ZN(n4495) );
  NAND2_X1 U5266 ( .A1(n8170), .A2(n4494), .ZN(n4493) );
  NAND2_X1 U5267 ( .A1(n4501), .A2(n4497), .ZN(n4496) );
  INV_X1 U5268 ( .A(n7808), .ZN(n4596) );
  NOR2_X1 U5269 ( .A1(n4260), .A2(n8100), .ZN(n4709) );
  NAND2_X1 U5270 ( .A1(n4486), .A2(n8111), .ZN(n4430) );
  OR2_X1 U5271 ( .A1(n9307), .A2(n9035), .ZN(n8767) );
  INV_X1 U5272 ( .A(n4665), .ZN(n4663) );
  NOR2_X1 U5273 ( .A1(n9029), .A2(n4671), .ZN(n4670) );
  INV_X1 U5274 ( .A(n9027), .ZN(n4671) );
  INV_X1 U5275 ( .A(n5406), .ZN(n4572) );
  INV_X1 U5276 ( .A(n5875), .ZN(n4503) );
  INV_X1 U5277 ( .A(n5305), .ZN(n4566) );
  INV_X1 U5278 ( .A(n4805), .ZN(n4550) );
  INV_X1 U5279 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5112) );
  INV_X1 U5280 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5089) );
  INV_X1 U5281 ( .A(n5035), .ZN(n4532) );
  INV_X1 U5282 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5038) );
  INV_X1 U5283 ( .A(n7830), .ZN(n7832) );
  NAND2_X1 U5284 ( .A1(n5121), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5146) );
  INV_X1 U5285 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5145) );
  NOR2_X1 U5286 ( .A1(n8346), .A2(n4430), .ZN(n4429) );
  NOR2_X1 U5287 ( .A1(n4596), .A2(n4593), .ZN(n4592) );
  OAI21_X1 U5288 ( .B1(n7807), .B2(n4596), .A(n7809), .ZN(n4595) );
  AOI21_X1 U5289 ( .B1(n4377), .B2(n4379), .A(n4376), .ZN(n4375) );
  INV_X1 U5290 ( .A(n4709), .ZN(n4376) );
  NAND2_X1 U5291 ( .A1(n4709), .A2(n8098), .ZN(n4708) );
  AND2_X1 U5292 ( .A1(n8276), .A2(n7871), .ZN(n7765) );
  AND2_X1 U5293 ( .A1(n8392), .A2(n8260), .ZN(n7766) );
  INV_X1 U5294 ( .A(n4276), .ZN(n4379) );
  NOR2_X1 U5295 ( .A1(n7701), .A2(n7783), .ZN(n4584) );
  INV_X1 U5296 ( .A(n7704), .ZN(n4586) );
  AND2_X1 U5297 ( .A1(n7686), .A2(n4686), .ZN(n4684) );
  INV_X1 U5298 ( .A(n7362), .ZN(n4397) );
  NOR2_X1 U5299 ( .A1(n7363), .A2(n4399), .ZN(n4398) );
  INV_X1 U5300 ( .A(n7163), .ZN(n4399) );
  NAND2_X1 U5301 ( .A1(n4705), .A2(n4704), .ZN(n7690) );
  NOR2_X1 U5302 ( .A1(n7056), .A2(n9969), .ZN(n4419) );
  AND2_X1 U5303 ( .A1(n7632), .A2(n6898), .ZN(n7635) );
  AND2_X1 U5304 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n4960) );
  NAND2_X1 U5305 ( .A1(n7654), .A2(n6918), .ZN(n7645) );
  NAND2_X1 U5306 ( .A1(n4248), .A2(n9937), .ZN(n7655) );
  INV_X1 U5307 ( .A(n7061), .ZN(n6717) );
  AND3_X1 U5308 ( .A1(n4843), .A2(n4819), .A3(n4818), .ZN(n4822) );
  OR2_X1 U5309 ( .A1(n5117), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5142) );
  AND2_X1 U5310 ( .A1(n5068), .A2(n5067), .ZN(n5091) );
  NOR2_X1 U5311 ( .A1(n4634), .A2(n4349), .ZN(n4348) );
  NOR3_X1 U5312 ( .A1(n4350), .A2(n4611), .A3(n4635), .ZN(n4349) );
  OR2_X1 U5313 ( .A1(n4628), .A2(n4630), .ZN(n4627) );
  AND2_X1 U5314 ( .A1(n6069), .A2(n8550), .ZN(n4630) );
  AND2_X1 U5315 ( .A1(n4364), .A2(n6104), .ZN(n4363) );
  AND2_X1 U5316 ( .A1(n6086), .A2(n6069), .ZN(n4628) );
  AOI21_X1 U5317 ( .B1(n7230), .B2(n5839), .A(n4612), .ZN(n4611) );
  INV_X1 U5318 ( .A(n7335), .ZN(n4612) );
  NAND2_X1 U5319 ( .A1(n4344), .A2(n4346), .ZN(n6015) );
  AOI21_X1 U5320 ( .B1(n4632), .B2(n4347), .A(n4316), .ZN(n4346) );
  OR2_X1 U5321 ( .A1(n9062), .A2(n8705), .ZN(n4562) );
  AND2_X1 U5322 ( .A1(n4439), .A2(n4438), .ZN(n7499) );
  NAND2_X1 U5323 ( .A1(n7266), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4438) );
  NOR2_X1 U5324 ( .A1(n8771), .A2(n4512), .ZN(n4511) );
  AND2_X1 U5325 ( .A1(n8767), .A2(n9031), .ZN(n9030) );
  NOR2_X1 U5326 ( .A1(n9005), .A2(n4666), .ZN(n4665) );
  INV_X1 U5327 ( .A(n4668), .ZN(n4666) );
  AOI21_X1 U5328 ( .B1(n4672), .B2(n4670), .A(n4669), .ZN(n4668) );
  OR2_X1 U5329 ( .A1(n9311), .A2(n9007), .ZN(n8824) );
  INV_X1 U5330 ( .A(n9026), .ZN(n4672) );
  NOR2_X1 U5331 ( .A1(n9487), .A2(n4516), .ZN(n4515) );
  INV_X1 U5332 ( .A(n4517), .ZN(n4516) );
  NOR2_X1 U5333 ( .A1(n9493), .A2(n9499), .ZN(n4517) );
  OR2_X1 U5334 ( .A1(n9493), .A2(n8668), .ZN(n8779) );
  OR2_X1 U5335 ( .A1(n5946), .A2(n7505), .ZN(n5968) );
  OR2_X1 U5336 ( .A1(n9521), .A2(n4523), .ZN(n4522) );
  OR2_X1 U5337 ( .A1(n7435), .A2(n9597), .ZN(n4523) );
  INV_X1 U5338 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U5339 ( .A1(n9784), .A2(n8899), .ZN(n8843) );
  NAND2_X1 U5340 ( .A1(n4774), .A2(n4776), .ZN(n4770) );
  OR2_X1 U5341 ( .A1(n4771), .A2(n8989), .ZN(n4769) );
  NOR2_X1 U5342 ( .A1(n6476), .A2(n6338), .ZN(n6465) );
  INV_X1 U5343 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4794) );
  AND2_X1 U5344 ( .A1(n5451), .A2(n5433), .ZN(n5449) );
  NOR2_X1 U5345 ( .A1(n5407), .A2(n4575), .ZN(n4574) );
  INV_X1 U5346 ( .A(n5372), .ZN(n4575) );
  NAND2_X1 U5347 ( .A1(n9458), .A2(n4369), .ZN(n4368) );
  AND2_X1 U5348 ( .A1(n5322), .A2(n5309), .ZN(n5320) );
  INV_X1 U5349 ( .A(n5277), .ZN(n5278) );
  NAND2_X1 U5350 ( .A1(n4535), .A2(n4536), .ZN(n5262) );
  AOI21_X1 U5351 ( .B1(n4539), .B2(n5187), .A(n4537), .ZN(n4536) );
  INV_X1 U5352 ( .A(n4542), .ZN(n4537) );
  NOR2_X1 U5353 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5571) );
  INV_X1 U5354 ( .A(SI_10_), .ZN(n5063) );
  XNOR2_X1 U5355 ( .A(n5017), .B(SI_7_), .ZN(n5014) );
  XNOR2_X1 U5356 ( .A(n4996), .B(SI_6_), .ZN(n4993) );
  OAI21_X1 U5357 ( .B1(n7613), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n4331), .ZN(
        n4953) );
  NAND2_X1 U5358 ( .A1(n7613), .A2(n6357), .ZN(n4331) );
  INV_X1 U5359 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4717) );
  OR2_X1 U5360 ( .A1(n5146), .A2(n5145), .ZN(n5168) );
  AND2_X1 U5361 ( .A1(n5470), .A2(n5469), .ZN(n5538) );
  INV_X1 U5362 ( .A(n5302), .ZN(n4762) );
  NAND2_X1 U5363 ( .A1(n4765), .A2(n4764), .ZN(n4763) );
  INV_X1 U5364 ( .A(n5318), .ZN(n4764) );
  INV_X1 U5365 ( .A(n5319), .ZN(n4765) );
  INV_X1 U5366 ( .A(n5313), .ZN(n5312) );
  NAND2_X1 U5367 ( .A1(n4723), .A2(n4722), .ZN(n4725) );
  INV_X1 U5368 ( .A(n4726), .ZN(n4722) );
  INV_X1 U5369 ( .A(n5543), .ZN(n7845) );
  AND2_X1 U5370 ( .A1(n4475), .A2(n4472), .ZN(n7753) );
  NOR2_X1 U5371 ( .A1(n4473), .A2(n7830), .ZN(n4472) );
  AND2_X1 U5372 ( .A1(n5355), .A2(n5354), .ZN(n7872) );
  AND4_X1 U5374 ( .A1(n5207), .A2(n5206), .A3(n5205), .A4(n5204), .ZN(n7525)
         );
  AND4_X1 U5375 ( .A1(n5128), .A2(n5127), .A3(n5126), .A4(n5125), .ZN(n7365)
         );
  AND4_X1 U5376 ( .A1(n5079), .A2(n5078), .A3(n5077), .A4(n5076), .ZN(n7203)
         );
  INV_X1 U5377 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4729) );
  NAND2_X1 U5378 ( .A1(n6558), .A2(n4880), .ZN(n6533) );
  NAND2_X1 U5379 ( .A1(n7620), .A2(n7619), .ZN(n8089) );
  AND2_X1 U5380 ( .A1(n8177), .A2(n4426), .ZN(n8088) );
  NOR2_X1 U5381 ( .A1(n8089), .A2(n4427), .ZN(n4426) );
  INV_X1 U5382 ( .A(n4429), .ZN(n4427) );
  OR2_X1 U5383 ( .A1(n8155), .A2(n4691), .ZN(n4690) );
  INV_X1 U5384 ( .A(n8112), .ZN(n4691) );
  NOR2_X1 U5385 ( .A1(n7822), .A2(n4799), .ZN(n7823) );
  OR2_X1 U5386 ( .A1(n8156), .A2(n8155), .ZN(n8160) );
  NOR2_X1 U5387 ( .A1(n8190), .A2(n8362), .ZN(n8177) );
  NAND2_X1 U5388 ( .A1(n8181), .A2(n8157), .ZN(n8109) );
  NAND2_X1 U5389 ( .A1(n8200), .A2(n8191), .ZN(n8190) );
  NOR2_X1 U5390 ( .A1(n4807), .A2(n7627), .ZN(n8228) );
  AND2_X1 U5391 ( .A1(n8205), .A2(n8228), .ZN(n8200) );
  OR2_X1 U5392 ( .A1(n8216), .A2(n8104), .ZN(n8217) );
  INV_X1 U5393 ( .A(n7947), .ZN(n8244) );
  NAND2_X1 U5394 ( .A1(n8258), .A2(n8259), .ZN(n8257) );
  NOR2_X1 U5395 ( .A1(n4413), .A2(n8385), .ZN(n4412) );
  AND2_X1 U5396 ( .A1(n7764), .A2(n8241), .ZN(n8259) );
  NOR2_X1 U5397 ( .A1(n8303), .A2(n4414), .ZN(n8294) );
  INV_X1 U5398 ( .A(n5268), .ZN(n5266) );
  OR2_X1 U5399 ( .A1(n5290), .A2(n5289), .ZN(n5313) );
  NAND2_X1 U5400 ( .A1(n8285), .A2(n7807), .ZN(n8287) );
  NAND2_X1 U5401 ( .A1(n7805), .A2(n7804), .ZN(n8309) );
  AND2_X1 U5402 ( .A1(n7457), .A2(n4421), .ZN(n7576) );
  NOR2_X1 U5403 ( .A1(n7591), .A2(n4422), .ZN(n4421) );
  INV_X1 U5404 ( .A(n4423), .ZN(n4422) );
  AND2_X1 U5405 ( .A1(n7708), .A2(n7707), .ZN(n7787) );
  NAND2_X1 U5406 ( .A1(n5199), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5225) );
  INV_X1 U5407 ( .A(n5201), .ZN(n5199) );
  NAND2_X1 U5408 ( .A1(n7457), .A2(n4425), .ZN(n7491) );
  AOI21_X1 U5409 ( .B1(n7466), .B2(n7784), .A(n4795), .ZN(n7467) );
  AND2_X1 U5410 ( .A1(n7369), .A2(n9984), .ZN(n7457) );
  AOI21_X1 U5411 ( .B1(n4600), .B2(n4602), .A(n4598), .ZN(n4597) );
  INV_X1 U5412 ( .A(n7684), .ZN(n4598) );
  NAND2_X1 U5413 ( .A1(n5072), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5095) );
  INV_X1 U5414 ( .A(n5073), .ZN(n5072) );
  AND2_X1 U5415 ( .A1(n6952), .A2(n4268), .ZN(n7349) );
  INV_X1 U5416 ( .A(n7777), .ZN(n7160) );
  NAND2_X1 U5417 ( .A1(n6952), .A2(n4417), .ZN(n7208) );
  AND2_X1 U5418 ( .A1(n7676), .A2(n7671), .ZN(n7777) );
  OAI21_X1 U5419 ( .B1(n6900), .B2(n4580), .A(n4577), .ZN(n4582) );
  INV_X1 U5420 ( .A(n4578), .ZN(n4577) );
  OR2_X1 U5421 ( .A1(n7774), .A2(n4581), .ZN(n4580) );
  NAND2_X1 U5422 ( .A1(n6952), .A2(n6956), .ZN(n6976) );
  NAND2_X1 U5423 ( .A1(n5003), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5049) );
  OAI211_X1 U5424 ( .C1(n6910), .C2(n6912), .A(n4408), .B(n4401), .ZN(n4404)
         );
  NAND2_X1 U5425 ( .A1(n7773), .A2(n4402), .ZN(n4401) );
  INV_X1 U5426 ( .A(n4279), .ZN(n4402) );
  OR2_X1 U5427 ( .A1(n9870), .A2(n9945), .ZN(n6723) );
  NAND2_X1 U5428 ( .A1(n7641), .A2(n7632), .ZN(n7772) );
  INV_X1 U5429 ( .A(n9855), .ZN(n4371) );
  NAND2_X1 U5430 ( .A1(n7634), .A2(n4589), .ZN(n4588) );
  INV_X1 U5431 ( .A(n7653), .ZN(n4589) );
  AND3_X1 U5432 ( .A1(n4391), .A2(n4390), .A3(n4388), .ZN(n9872) );
  NAND2_X1 U5433 ( .A1(n6405), .A2(n7978), .ZN(n4391) );
  NAND2_X1 U5434 ( .A1(n7743), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4390) );
  NAND2_X1 U5435 ( .A1(n4251), .A2(n4389), .ZN(n4388) );
  INV_X1 U5436 ( .A(n9872), .ZN(n9873) );
  NAND2_X1 U5437 ( .A1(n9871), .A2(n9872), .ZN(n9870) );
  NAND2_X1 U5438 ( .A1(n6729), .A2(n6728), .ZN(n8332) );
  AND2_X1 U5439 ( .A1(n8326), .A2(n9937), .ZN(n9871) );
  NAND2_X1 U5440 ( .A1(n5345), .A2(n5344), .ZN(n8380) );
  NAND2_X1 U5441 ( .A1(n6947), .A2(n7662), .ZN(n6968) );
  NAND2_X1 U5442 ( .A1(n9858), .A2(n9857), .ZN(n9860) );
  NAND2_X1 U5443 ( .A1(n4825), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4826) );
  NOR2_X1 U5444 ( .A1(n5502), .A2(n5501), .ZN(n5507) );
  INV_X1 U5445 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5512) );
  NOR2_X1 U5446 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n4837) );
  INV_X1 U5447 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4838) );
  INV_X1 U5448 ( .A(n6159), .ZN(n4640) );
  NOR2_X1 U5449 ( .A1(n6159), .A2(n4360), .ZN(n4638) );
  OR2_X1 U5450 ( .A1(n6442), .A2(n6855), .ZN(n5642) );
  INV_X1 U5451 ( .A(n4620), .ZN(n4617) );
  NOR2_X1 U5452 ( .A1(n4619), .A2(n8490), .ZN(n4614) );
  INV_X1 U5453 ( .A(n8537), .ZN(n4619) );
  NAND2_X1 U5454 ( .A1(n5881), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U5455 ( .A1(n5966), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5984) );
  INV_X1 U5456 ( .A(n5968), .ZN(n5966) );
  NAND2_X1 U5457 ( .A1(n6089), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6108) );
  OR2_X1 U5458 ( .A1(n7227), .A2(n7230), .ZN(n7228) );
  NAND2_X1 U5459 ( .A1(n6032), .A2(n6031), .ZN(n4620) );
  NAND2_X1 U5460 ( .A1(n5859), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5882) );
  INV_X1 U5461 ( .A(n5861), .ZN(n5859) );
  NAND2_X1 U5462 ( .A1(n4343), .A2(n5680), .ZN(n6623) );
  INV_X1 U5463 ( .A(n6485), .ZN(n5662) );
  NAND2_X1 U5464 ( .A1(n6336), .A2(n9541), .ZN(n6476) );
  OR2_X1 U5465 ( .A1(n8718), .A2(n8875), .ZN(n6336) );
  AND2_X1 U5466 ( .A1(n6227), .A2(n6443), .ZN(n8585) );
  NAND2_X1 U5467 ( .A1(n6206), .A2(n4246), .ZN(n8718) );
  AND3_X1 U5468 ( .A1(n6429), .A2(n6428), .A3(n6427), .ZN(n8977) );
  NAND2_X1 U5469 ( .A1(n5686), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5645) );
  AND2_X1 U5470 ( .A1(n5618), .A2(n5619), .ZN(n4651) );
  AND2_X1 U5471 ( .A1(n8915), .A2(n4450), .ZN(n9628) );
  NAND2_X1 U5472 ( .A1(n8914), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4450) );
  NAND2_X1 U5473 ( .A1(n9628), .A2(n9629), .ZN(n9627) );
  NAND2_X1 U5474 ( .A1(n9627), .A2(n4449), .ZN(n9646) );
  OR2_X1 U5475 ( .A1(n9631), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4449) );
  AOI21_X1 U5476 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6316), .A(n6309), .ZN(
        n6412) );
  NAND2_X1 U5477 ( .A1(n6412), .A2(n6413), .ZN(n6411) );
  NAND2_X1 U5478 ( .A1(n6411), .A2(n4434), .ZN(n9667) );
  OR2_X1 U5479 ( .A1(n6419), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4434) );
  NOR2_X1 U5480 ( .A1(n6491), .A2(n4443), .ZN(n9682) );
  AND2_X1 U5481 ( .A1(n6498), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4443) );
  NOR2_X1 U5482 ( .A1(n9682), .A2(n9681), .ZN(n9680) );
  NOR2_X1 U5483 ( .A1(n9680), .A2(n4442), .ZN(n6494) );
  AND2_X1 U5484 ( .A1(n9674), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4442) );
  OR2_X1 U5485 ( .A1(n5840), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5855) );
  NOR2_X1 U5486 ( .A1(n7503), .A2(n7502), .ZN(n7545) );
  AOI21_X1 U5487 ( .B1(n8962), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8955), .ZN(
        n9694) );
  AND2_X1 U5488 ( .A1(n4509), .A2(n4511), .ZN(n4507) );
  INV_X1 U5489 ( .A(n9585), .ZN(n4509) );
  INV_X1 U5490 ( .A(n4511), .ZN(n4505) );
  AOI21_X1 U5491 ( .B1(n9006), .B2(n9005), .A(n4296), .ZN(n9051) );
  INV_X1 U5492 ( .A(n4512), .ZN(n4510) );
  AND2_X1 U5493 ( .A1(n8824), .A2(n8769), .ZN(n9076) );
  NAND2_X1 U5494 ( .A1(n9078), .A2(n9756), .ZN(n4327) );
  NAND2_X1 U5495 ( .A1(n9090), .A2(n9756), .ZN(n4330) );
  NAND2_X1 U5496 ( .A1(n9095), .A2(n9104), .ZN(n4778) );
  AND2_X1 U5497 ( .A1(n8783), .A2(n9025), .ZN(n9118) );
  NAND2_X1 U5498 ( .A1(n6073), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6091) );
  INV_X1 U5499 ( .A(n6074), .ZN(n6073) );
  AOI21_X1 U5500 ( .B1(n4657), .B2(n4658), .A(n4655), .ZN(n4654) );
  INV_X1 U5501 ( .A(n9021), .ZN(n4655) );
  AND2_X1 U5502 ( .A1(n9236), .A2(n4514), .ZN(n9170) );
  AND2_X1 U5503 ( .A1(n9174), .A2(n4515), .ZN(n4514) );
  AND2_X1 U5504 ( .A1(n9163), .A2(n4785), .ZN(n4783) );
  OAI21_X1 U5505 ( .B1(n4784), .B2(n9020), .A(n4297), .ZN(n4782) );
  NAND2_X1 U5506 ( .A1(n6021), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U5507 ( .A1(n9236), .A2(n4517), .ZN(n9197) );
  AND2_X1 U5508 ( .A1(n8779), .A2(n8722), .ZN(n9194) );
  NAND2_X1 U5509 ( .A1(n9236), .A2(n9227), .ZN(n9228) );
  NOR2_X1 U5510 ( .A1(n4677), .A2(n4675), .ZN(n4674) );
  INV_X1 U5511 ( .A(n9015), .ZN(n4675) );
  AND2_X1 U5512 ( .A1(n8723), .A2(n8787), .ZN(n9218) );
  OR2_X1 U5513 ( .A1(n9271), .A2(n9511), .ZN(n9253) );
  OAI21_X1 U5514 ( .B1(n9282), .B2(n9281), .A(n9011), .ZN(n9263) );
  OR2_X1 U5515 ( .A1(n9589), .A2(n9284), .ZN(n4802) );
  NOR2_X1 U5516 ( .A1(n7324), .A2(n4523), .ZN(n9286) );
  INV_X1 U5517 ( .A(n9266), .ZN(n8985) );
  INV_X1 U5518 ( .A(n8889), .ZN(n9284) );
  NOR2_X1 U5519 ( .A1(n7320), .A2(n7319), .ZN(n7398) );
  NOR2_X1 U5520 ( .A1(n7324), .A2(n9597), .ZN(n7404) );
  OR2_X1 U5521 ( .A1(n7191), .A2(n7193), .ZN(n7324) );
  AND2_X1 U5522 ( .A1(n8637), .A2(n7397), .ZN(n8737) );
  INV_X1 U5523 ( .A(n7129), .ZN(n7131) );
  INV_X1 U5524 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5825) );
  OR2_X1 U5525 ( .A1(n5826), .A2(n5825), .ZN(n5845) );
  AND2_X1 U5526 ( .A1(n7102), .A2(n9818), .ZN(n7138) );
  INV_X1 U5527 ( .A(n8892), .ZN(n7187) );
  AOI21_X1 U5528 ( .B1(n7001), .B2(n7000), .A(n6999), .ZN(n7185) );
  AOI21_X1 U5529 ( .B1(n4649), .B2(n4647), .A(n4646), .ZN(n4645) );
  INV_X1 U5530 ( .A(n4649), .ZN(n4648) );
  NOR2_X1 U5531 ( .A1(n6840), .A2(n8618), .ZN(n4649) );
  OR2_X1 U5532 ( .A1(n6872), .A2(n6998), .ZN(n7005) );
  NAND2_X1 U5533 ( .A1(n6879), .A2(n8851), .ZN(n4650) );
  OR2_X1 U5534 ( .A1(n9716), .A2(n6830), .ZN(n6882) );
  NOR2_X1 U5535 ( .A1(n6882), .A2(n6892), .ZN(n6884) );
  AND2_X1 U5536 ( .A1(n8851), .A2(n8795), .ZN(n8727) );
  NAND2_X1 U5537 ( .A1(n4519), .A2(n9784), .ZN(n9716) );
  INV_X1 U5538 ( .A(n9714), .ZN(n4519) );
  NAND2_X1 U5539 ( .A1(n4520), .A2(n9778), .ZN(n9714) );
  CLKBUF_X1 U5540 ( .A(n5640), .Z(n6340) );
  NAND2_X1 U5541 ( .A1(n6106), .A2(n6105), .ZN(n9327) );
  OR2_X1 U5542 ( .A1(n8705), .A2(n8837), .ZN(n9587) );
  NAND2_X1 U5543 ( .A1(n5843), .A2(n5842), .ZN(n7121) );
  INV_X1 U5544 ( .A(n9815), .ZN(n9524) );
  CLKBUF_X1 U5545 ( .A(n6886), .Z(n6887) );
  NAND2_X1 U5546 ( .A1(n9737), .A2(n6326), .ZN(n6328) );
  XNOR2_X1 U5547 ( .A(n7741), .B(n7740), .ZN(n8606) );
  NAND2_X1 U5548 ( .A1(n5452), .A2(n5451), .ZN(n5474) );
  NAND2_X1 U5549 ( .A1(n5450), .A2(n5449), .ZN(n5452) );
  AND2_X1 U5550 ( .A1(n5475), .A2(n5456), .ZN(n5473) );
  XNOR2_X1 U5551 ( .A(n5450), .B(n5449), .ZN(n7536) );
  NAND2_X1 U5552 ( .A1(n4546), .A2(n5213), .ZN(n5240) );
  NAND2_X1 U5553 ( .A1(n4547), .A2(n4538), .ZN(n4546) );
  INV_X1 U5554 ( .A(n4540), .ZN(n4538) );
  AND2_X1 U5555 ( .A1(n4351), .A2(n5570), .ZN(n5918) );
  AND2_X1 U5556 ( .A1(n4797), .A2(n4353), .ZN(n4351) );
  OAI21_X1 U5557 ( .B1(n5088), .B2(n4273), .A(n4551), .ZN(n5159) );
  AND2_X1 U5558 ( .A1(n4797), .A2(n4354), .ZN(n4352) );
  NAND2_X1 U5559 ( .A1(n4554), .A2(n5108), .ZN(n5137) );
  XNOR2_X1 U5560 ( .A(n5086), .B(n4271), .ZN(n6398) );
  NAND2_X1 U5561 ( .A1(n4530), .A2(n5035), .ZN(n5061) );
  NAND2_X1 U5562 ( .A1(n4693), .A2(n4692), .ZN(n5037) );
  XNOR2_X1 U5563 ( .A(n4953), .B(SI_4_), .ZN(n4951) );
  AND3_X1 U5564 ( .A1(n5669), .A2(n4788), .A3(n5565), .ZN(n5720) );
  NOR2_X1 U5565 ( .A1(n7309), .A2(n10049), .ZN(n7310) );
  NAND2_X1 U5566 ( .A1(n5166), .A2(n5165), .ZN(n7488) );
  AOI21_X1 U5567 ( .B1(n4735), .B2(n4737), .A(n4317), .ZN(n4732) );
  NAND2_X1 U5568 ( .A1(n7582), .A2(n4735), .ZN(n4733) );
  NAND2_X1 U5569 ( .A1(n4758), .A2(n4763), .ZN(n7868) );
  NAND2_X1 U5570 ( .A1(n4341), .A2(n4278), .ZN(n4758) );
  INV_X1 U5571 ( .A(n7951), .ZN(n7693) );
  NAND2_X1 U5572 ( .A1(n7890), .A2(n8313), .ZN(n7939) );
  NAND2_X1 U5573 ( .A1(n4804), .A2(n5401), .ZN(n5402) );
  NAND2_X1 U5574 ( .A1(n5400), .A2(n7898), .ZN(n5401) );
  AOI21_X1 U5575 ( .B1(n6360), .B2(n7742), .A(n4489), .ZN(n4488) );
  NOR2_X1 U5576 ( .A1(n4880), .A2(n6365), .ZN(n4489) );
  NAND2_X1 U5577 ( .A1(n6754), .A2(n4948), .ZN(n6638) );
  AND2_X1 U5578 ( .A1(n5555), .A2(n7845), .ZN(n7890) );
  NAND2_X1 U5579 ( .A1(n4293), .A2(n7914), .ZN(n7896) );
  NAND2_X1 U5580 ( .A1(n5376), .A2(n5375), .ZN(n8371) );
  CLKBUF_X1 U5581 ( .A(n6753), .Z(n6754) );
  NAND2_X1 U5582 ( .A1(n4341), .A2(n5302), .ZN(n7908) );
  NAND2_X1 U5583 ( .A1(n7215), .A2(n5134), .ZN(n7246) );
  NOR2_X1 U5584 ( .A1(n5080), .A2(n4749), .ZN(n4748) );
  NAND2_X1 U5585 ( .A1(n6389), .A2(n7742), .ZN(n4706) );
  NAND2_X1 U5586 ( .A1(n6585), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7925) );
  NAND2_X1 U5587 ( .A1(n7582), .A2(n4738), .ZN(n4734) );
  AND2_X1 U5588 ( .A1(n5555), .A2(n5534), .ZN(n7933) );
  NAND2_X1 U5589 ( .A1(n5198), .A2(n5197), .ZN(n8419) );
  AND2_X1 U5590 ( .A1(n5554), .A2(n5553), .ZN(n8134) );
  INV_X2 U5591 ( .A(P2_U3966), .ZN(n7961) );
  INV_X1 U5592 ( .A(n8082), .ZN(n9850) );
  INV_X1 U5593 ( .A(n9848), .ZN(n9844) );
  AND2_X1 U5594 ( .A1(n5461), .A2(n5437), .ZN(n8178) );
  XNOR2_X1 U5595 ( .A(n8173), .B(n7817), .ZN(n8175) );
  NAND2_X1 U5596 ( .A1(n5414), .A2(n5413), .ZN(n8366) );
  OAI21_X1 U5597 ( .B1(n8250), .B2(n4385), .A(n4383), .ZN(n8223) );
  OAI21_X1 U5598 ( .B1(n8250), .B2(n8103), .A(n4257), .ZN(n8233) );
  AND2_X1 U5599 ( .A1(n4710), .A2(n4711), .ZN(n8284) );
  OR2_X1 U5600 ( .A1(n8301), .A2(n8098), .ZN(n4710) );
  NAND2_X1 U5601 ( .A1(n4712), .A2(n4276), .ZN(n8096) );
  NAND2_X1 U5602 ( .A1(n7485), .A2(n7786), .ZN(n7524) );
  NAND2_X1 U5603 ( .A1(n4687), .A2(n4685), .ZN(n7465) );
  NAND2_X1 U5604 ( .A1(n4687), .A2(n4686), .ZN(n7452) );
  AND2_X1 U5605 ( .A1(n4604), .A2(n7671), .ZN(n7166) );
  OR2_X1 U5606 ( .A1(n8195), .A2(n9985), .ZN(n8278) );
  INV_X1 U5607 ( .A(n9953), .ZN(n6909) );
  INV_X1 U5608 ( .A(n8278), .ZN(n8319) );
  INV_X1 U5609 ( .A(n9857), .ZN(n9856) );
  OAI211_X1 U5610 ( .C1(n4957), .C2(n6359), .A(n4901), .B(n4900), .ZN(n8323)
         );
  INV_X1 U5611 ( .A(n8307), .ZN(n8324) );
  INV_X1 U5612 ( .A(n8321), .ZN(n8325) );
  NAND2_X1 U5613 ( .A1(n4880), .A2(n8469), .ZN(n4409) );
  AND2_X2 U5614 ( .A1(n7065), .A2(n7064), .ZN(n10008) );
  NOR2_X1 U5615 ( .A1(n4606), .A2(n4292), .ZN(n8347) );
  INV_X1 U5616 ( .A(n8349), .ZN(n8354) );
  OR3_X1 U5617 ( .A1(n8396), .A2(n8395), .A3(n8394), .ZN(n8449) );
  AND2_X2 U5618 ( .A1(n7051), .A2(n7050), .ZN(n9993) );
  INV_X1 U5619 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4609) );
  NAND2_X1 U5620 ( .A1(n4851), .A2(n4850), .ZN(n4853) );
  NAND2_X1 U5621 ( .A1(n4823), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4850) );
  NAND2_X1 U5622 ( .A1(n5506), .A2(n5505), .ZN(n7538) );
  XNOR2_X1 U5623 ( .A(n5517), .B(n5516), .ZN(n7392) );
  INV_X1 U5624 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7595) );
  INV_X1 U5625 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7049) );
  INV_X1 U5626 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7025) );
  INV_X1 U5627 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6863) );
  INV_X1 U5628 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6636) );
  INV_X1 U5629 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6592) );
  INV_X1 U5630 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6439) );
  INV_X1 U5631 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6435) );
  INV_X1 U5632 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6426) );
  INV_X1 U5633 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6399) );
  INV_X1 U5634 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6380) );
  NOR2_X1 U5635 ( .A1(n6272), .A2(n6270), .ZN(n6448) );
  AND2_X1 U5636 ( .A1(n5710), .A2(n5708), .ZN(n6624) );
  INV_X1 U5637 ( .A(n8895), .ZN(n7152) );
  OAI211_X1 U5638 ( .C1(n8530), .C2(n4259), .A(n4357), .B(n4356), .ZN(n8569)
         );
  NAND2_X1 U5639 ( .A1(n4360), .A2(n6126), .ZN(n4356) );
  NAND2_X1 U5640 ( .A1(n6128), .A2(n6127), .ZN(n9321) );
  INV_X1 U5641 ( .A(n8898), .ZN(n9722) );
  NAND2_X1 U5642 ( .A1(n4345), .A2(n4632), .ZN(n8519) );
  NAND2_X1 U5643 ( .A1(n8511), .A2(n5980), .ZN(n8520) );
  NAND2_X1 U5644 ( .A1(n8510), .A2(n5980), .ZN(n4345) );
  AND4_X1 U5645 ( .A1(n5812), .A2(n5811), .A3(n5810), .A4(n5809), .ZN(n7235)
         );
  NAND2_X1 U5646 ( .A1(n7411), .A2(n5899), .ZN(n7428) );
  NAND2_X1 U5647 ( .A1(n6070), .A2(n6069), .ZN(n4631) );
  NAND2_X1 U5648 ( .A1(n6072), .A2(n6071), .ZN(n9479) );
  INV_X1 U5649 ( .A(n8890), .ZN(n7433) );
  INV_X1 U5650 ( .A(n8563), .ZN(n8583) );
  INV_X1 U5651 ( .A(n8571), .ZN(n8592) );
  INV_X1 U5652 ( .A(n9265), .ZN(n8645) );
  NAND2_X1 U5653 ( .A1(n5945), .A2(n5944), .ZN(n9514) );
  NAND2_X1 U5654 ( .A1(n8713), .A2(n4558), .ZN(n4557) );
  NAND2_X1 U5655 ( .A1(n6151), .A2(n6150), .ZN(n9105) );
  NAND2_X1 U5656 ( .A1(n6138), .A2(n6137), .ZN(n9120) );
  OR2_X1 U5657 ( .A1(n9099), .A2(n6247), .ZN(n6138) );
  NAND4_X1 U5658 ( .A1(n5755), .A2(n5754), .A3(n5753), .A4(n5752), .ZN(n8896)
         );
  NAND2_X1 U5659 ( .A1(n8905), .A2(n8904), .ZN(n8903) );
  NAND2_X1 U5660 ( .A1(n4432), .A2(n4431), .ZN(n6283) );
  OR2_X1 U5661 ( .A1(n9661), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4431) );
  NAND2_X1 U5662 ( .A1(n9667), .A2(n4433), .ZN(n4432) );
  INV_X1 U5663 ( .A(n9668), .ZN(n4433) );
  INV_X1 U5664 ( .A(n4441), .ZN(n8928) );
  INV_X1 U5665 ( .A(n4439), .ZN(n7265) );
  NAND2_X1 U5666 ( .A1(n4437), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4436) );
  NAND2_X1 U5667 ( .A1(n7546), .A2(n4437), .ZN(n4435) );
  INV_X1 U5668 ( .A(n7548), .ZN(n4437) );
  INV_X1 U5669 ( .A(n9697), .ZN(n9679) );
  NAND2_X1 U5670 ( .A1(n9064), .A2(n9063), .ZN(n9065) );
  NAND2_X1 U5671 ( .A1(n9061), .A2(n9060), .ZN(n9066) );
  NAND2_X1 U5672 ( .A1(n6088), .A2(n6087), .ZN(n9473) );
  NAND2_X1 U5673 ( .A1(n4653), .A2(n4657), .ZN(n9164) );
  NAND2_X1 U5674 ( .A1(n4781), .A2(n4784), .ZN(n9160) );
  NAND2_X1 U5675 ( .A1(n9191), .A2(n4785), .ZN(n4781) );
  AND2_X1 U5676 ( .A1(n9192), .A2(n8992), .ZN(n9178) );
  AND2_X1 U5677 ( .A1(n4676), .A2(n4678), .ZN(n9240) );
  AOI21_X1 U5678 ( .B1(n9247), .B2(n9249), .A(n4773), .ZN(n9235) );
  AND2_X1 U5679 ( .A1(n4679), .A2(n8646), .ZN(n9248) );
  NAND2_X1 U5680 ( .A1(n4779), .A2(n4780), .ZN(n7329) );
  AND2_X1 U5681 ( .A1(n6886), .A2(n6853), .ZN(n6865) );
  NAND2_X1 U5682 ( .A1(n9742), .A2(n6231), .ZN(n9222) );
  INV_X1 U5683 ( .A(n9733), .ZN(n9226) );
  AOI211_X1 U5684 ( .C1(n9742), .C2(n9564), .A(n9584), .B(n9563), .ZN(n9567)
         );
  AOI211_X1 U5685 ( .C1(n9598), .C2(n9585), .A(n9584), .B(n9583), .ZN(n9610)
         );
  AND2_X2 U5686 ( .A1(n6473), .A2(n6466), .ZN(n9828) );
  AND2_X1 U5687 ( .A1(n6191), .A2(n6190), .ZN(n9542) );
  AND2_X1 U5688 ( .A1(n6189), .A2(n6188), .ZN(n6472) );
  INV_X1 U5689 ( .A(n9765), .ZN(n9541) );
  XNOR2_X1 U5690 ( .A(n4529), .B(n7615), .ZN(n9543) );
  NAND2_X1 U5691 ( .A1(n7612), .A2(n7611), .ZN(n4529) );
  NAND2_X1 U5692 ( .A1(n5607), .A2(n5606), .ZN(n5608) );
  NOR2_X1 U5693 ( .A1(n5605), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5606) );
  XNOR2_X1 U5694 ( .A(n7598), .B(n7597), .ZN(n7568) );
  XNOR2_X1 U5695 ( .A(n5474), .B(n5473), .ZN(n7561) );
  INV_X1 U5696 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7244) );
  INV_X1 U5697 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7240) );
  NAND2_X1 U5698 ( .A1(n5576), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5578) );
  INV_X1 U5699 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7047) );
  INV_X1 U5700 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n9348) );
  INV_X1 U5701 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6861) );
  INV_X1 U5702 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9429) );
  INV_X1 U5703 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6508) );
  INV_X1 U5704 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6437) );
  INV_X1 U5705 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9427) );
  INV_X1 U5706 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6403) );
  INV_X1 U5707 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6387) );
  INV_X1 U5708 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9360) );
  OR2_X1 U5709 ( .A1(n5803), .A2(n5802), .ZN(n6381) );
  NAND2_X1 U5710 ( .A1(n4703), .A2(n4913), .ZN(n4929) );
  NAND2_X1 U5711 ( .A1(n4911), .A2(n4910), .ZN(n4703) );
  OAI21_X1 U5712 ( .B1(n5671), .B2(n5670), .A(n5692), .ZN(n6349) );
  XNOR2_X1 U5713 ( .A(n5649), .B(n5650), .ZN(n6351) );
  OAI21_X1 U5714 ( .B1(n6772), .B2(n6771), .A(n4751), .ZN(n6834) );
  NAND2_X1 U5715 ( .A1(n4741), .A2(n4744), .ZN(n6738) );
  AOI21_X1 U5716 ( .B1(n4262), .B2(n7224), .A(n4469), .ZN(n4468) );
  AOI21_X1 U5717 ( .B1(n4606), .B2(n8336), .A(n4298), .ZN(n8130) );
  NAND2_X1 U5718 ( .A1(n4641), .A2(n4313), .ZN(n6262) );
  OAI21_X1 U5719 ( .B1(n8970), .B2(n9744), .A(n4445), .ZN(P1_U3260) );
  AOI21_X1 U5720 ( .B1(n4447), .B2(n9744), .A(n4446), .ZN(n4445) );
  OAI21_X1 U5721 ( .B1(n9689), .B2(n4720), .A(n8971), .ZN(n4446) );
  NOR2_X1 U5722 ( .A1(n9314), .A2(n9234), .ZN(n9080) );
  NOR2_X1 U5723 ( .A1(n9319), .A2(n9291), .ZN(n9092) );
  AND2_X1 U5724 ( .A1(n7737), .A2(n7826), .ZN(n4253) );
  NOR2_X1 U5725 ( .A1(n7746), .A2(n4465), .ZN(n4254) );
  OR2_X1 U5726 ( .A1(n6746), .A2(n6745), .ZN(n4255) );
  AND2_X1 U5727 ( .A1(n8137), .A2(n4690), .ZN(n4256) );
  INV_X1 U5728 ( .A(n8298), .ZN(n8399) );
  AND2_X1 U5729 ( .A1(n5288), .A2(n5287), .ZN(n8298) );
  AND2_X1 U5730 ( .A1(n5468), .A2(n5467), .ZN(n8176) );
  OR2_X1 U5731 ( .A1(n8256), .A2(n8269), .ZN(n4257) );
  NAND2_X1 U5732 ( .A1(n4252), .A2(n5651), .ZN(n4258) );
  OR2_X1 U5733 ( .A1(n8503), .A2(n8528), .ZN(n4259) );
  AND4_X1 U5734 ( .A1(n5100), .A2(n5099), .A3(n5098), .A4(n5097), .ZN(n7368)
         );
  INV_X1 U5735 ( .A(n7368), .ZN(n4704) );
  NOR2_X1 U5736 ( .A1(n8298), .A2(n8268), .ZN(n4260) );
  AND2_X1 U5737 ( .A1(n4282), .A2(n4731), .ZN(n4261) );
  AND2_X1 U5738 ( .A1(n7843), .A2(n7842), .ZN(n4262) );
  INV_X1 U5739 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4354) );
  INV_X1 U5740 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4816) );
  NAND3_X1 U5741 ( .A1(n7795), .A2(n7751), .A3(n4465), .ZN(n4263) );
  AND2_X1 U5742 ( .A1(n7899), .A2(n5399), .ZN(n4264) );
  NAND2_X1 U5743 ( .A1(n4683), .A2(n4311), .ZN(n4265) );
  AND2_X1 U5744 ( .A1(n7801), .A2(n7224), .ZN(n4266) );
  NAND2_X1 U5745 ( .A1(n7591), .A2(n7948), .ZN(n4267) );
  AND2_X1 U5746 ( .A1(n4417), .A2(n4416), .ZN(n4268) );
  AND2_X1 U5747 ( .A1(n4610), .A2(n4609), .ZN(n4269) );
  NAND2_X1 U5748 ( .A1(n5479), .A2(n5478), .ZN(n8350) );
  INV_X1 U5749 ( .A(n8350), .ZN(n4486) );
  NAND2_X1 U5750 ( .A1(n4613), .A2(n4611), .ZN(n7334) );
  NAND2_X1 U5751 ( .A1(n5245), .A2(n5244), .ZN(n8093) );
  NAND2_X1 U5752 ( .A1(n4817), .A2(n4816), .ZN(n5242) );
  INV_X1 U5753 ( .A(n8851), .ZN(n4647) );
  AND2_X1 U5754 ( .A1(n7699), .A2(n7700), .ZN(n7697) );
  AND2_X1 U5755 ( .A1(n4323), .A2(n4866), .ZN(n4270) );
  NAND2_X1 U5756 ( .A1(n5533), .A2(n8077), .ZN(n7797) );
  AND2_X1 U5757 ( .A1(n5087), .A2(n5066), .ZN(n4271) );
  INV_X2 U5758 ( .A(n5643), .ZN(n5701) );
  AND2_X1 U5759 ( .A1(n4626), .A2(n4629), .ZN(n4272) );
  OR2_X1 U5760 ( .A1(n5136), .A2(n4553), .ZN(n4273) );
  OAI211_X1 U5761 ( .C1(n5668), .C2(n6352), .A(n5697), .B(n5696), .ZN(n9713)
         );
  INV_X1 U5762 ( .A(n7774), .ZN(n4400) );
  AND2_X1 U5763 ( .A1(n4583), .A2(n4585), .ZN(n4274) );
  OR2_X1 U5764 ( .A1(n8569), .A2(n6159), .ZN(n4275) );
  AND2_X1 U5765 ( .A1(n7789), .A2(n4267), .ZN(n4276) );
  NAND2_X1 U5766 ( .A1(n5668), .A2(n4789), .ZN(n4277) );
  NOR2_X1 U5767 ( .A1(n7907), .A2(n4762), .ZN(n4278) );
  NOR2_X1 U5768 ( .A1(n7958), .A2(n9953), .ZN(n4279) );
  OR2_X1 U5769 ( .A1(n8380), .A2(n8261), .ZN(n4280) );
  AND2_X1 U5770 ( .A1(n5640), .A2(n6272), .ZN(n5648) );
  INV_X1 U5771 ( .A(n4525), .ZN(n8973) );
  OAI21_X1 U5772 ( .B1(n9543), .B2(n8594), .A(n4526), .ZN(n4525) );
  NAND2_X1 U5773 ( .A1(n7960), .A2(n9872), .ZN(n7634) );
  XNOR2_X1 U5774 ( .A(n4826), .B(P2_IR_REG_29__SCAN_IN), .ZN(n4829) );
  INV_X1 U5775 ( .A(n8503), .ZN(n4360) );
  XNOR2_X1 U5776 ( .A(n5578), .B(n5577), .ZN(n5639) );
  NAND2_X1 U5777 ( .A1(n7731), .A2(n7819), .ZN(n8174) );
  NAND2_X1 U5778 ( .A1(n8610), .A2(n8609), .ZN(n8771) );
  AND2_X1 U5779 ( .A1(n7814), .A2(n7763), .ZN(n8240) );
  INV_X1 U5780 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4856) );
  AND2_X1 U5781 ( .A1(n6833), .A2(n4755), .ZN(n4281) );
  AND4_X1 U5782 ( .A1(n4822), .A2(n4821), .A3(n5500), .A4(n4820), .ZN(n4282)
         );
  AND2_X1 U5783 ( .A1(n5669), .A2(n4788), .ZN(n5717) );
  NAND2_X1 U5784 ( .A1(n4631), .A2(n6085), .ZN(n8547) );
  OR2_X1 U5785 ( .A1(n8402), .A2(n8097), .ZN(n8286) );
  NAND2_X1 U5786 ( .A1(n5983), .A2(n5982), .ZN(n9504) );
  OR2_X1 U5787 ( .A1(n4730), .A2(n4728), .ZN(n4998) );
  AND2_X1 U5788 ( .A1(n7810), .A2(n7808), .ZN(n4283) );
  NAND2_X1 U5789 ( .A1(n5144), .A2(n5143), .ZN(n8424) );
  INV_X1 U5790 ( .A(n4481), .ZN(n4480) );
  OAI21_X1 U5791 ( .B1(n4253), .B2(n4482), .A(n4487), .ZN(n4481) );
  NAND2_X1 U5792 ( .A1(n5223), .A2(n5222), .ZN(n7591) );
  AND2_X1 U5793 ( .A1(n7810), .A2(n8241), .ZN(n4284) );
  NAND2_X1 U5794 ( .A1(n6002), .A2(n6001), .ZN(n9499) );
  OR2_X1 U5795 ( .A1(n9487), .A2(n9168), .ZN(n4285) );
  AND2_X1 U5796 ( .A1(n4667), .A2(n4665), .ZN(n4286) );
  AND2_X1 U5797 ( .A1(n7675), .A2(n7685), .ZN(n7778) );
  NAND2_X1 U5798 ( .A1(n5324), .A2(n5323), .ZN(n8385) );
  NAND2_X1 U5799 ( .A1(n8806), .A2(n8705), .ZN(n4287) );
  OR2_X1 U5800 ( .A1(n8137), .A2(n8155), .ZN(n4288) );
  INV_X1 U5801 ( .A(n4776), .ZN(n4773) );
  NAND2_X1 U5802 ( .A1(n9511), .A2(n9265), .ZN(n4776) );
  NOR2_X1 U5803 ( .A1(n4659), .A2(n9161), .ZN(n4289) );
  AND2_X1 U5804 ( .A1(n8796), .A2(n8850), .ZN(n8729) );
  AND2_X1 U5805 ( .A1(n8286), .A2(n7768), .ZN(n8310) );
  INV_X1 U5806 ( .A(n8310), .ZN(n4593) );
  INV_X1 U5807 ( .A(n9028), .ZN(n4669) );
  AND2_X1 U5808 ( .A1(n4531), .A2(n5062), .ZN(n4290) );
  INV_X1 U5809 ( .A(n8346), .ZN(n8127) );
  NAND2_X1 U5810 ( .A1(n7745), .A2(n7744), .ZN(n8346) );
  AND2_X1 U5811 ( .A1(n7328), .A2(n4780), .ZN(n4291) );
  OAI21_X1 U5812 ( .B1(n5895), .B2(n4635), .A(n7425), .ZN(n4634) );
  OR2_X1 U5813 ( .A1(n8345), .A2(n4605), .ZN(n4292) );
  AND2_X1 U5814 ( .A1(n5359), .A2(n5398), .ZN(n4293) );
  NOR2_X1 U5815 ( .A1(n5085), .A2(n5084), .ZN(n4294) );
  INV_X1 U5816 ( .A(n8528), .ZN(n4364) );
  AND2_X1 U5817 ( .A1(n5017), .A2(SI_7_), .ZN(n4295) );
  AND2_X1 U5818 ( .A1(n9075), .A2(n9007), .ZN(n4296) );
  NAND2_X1 U5819 ( .A1(n9483), .A2(n9186), .ZN(n4297) );
  OR2_X1 U5820 ( .A1(n8129), .A2(n8128), .ZN(n4298) );
  INV_X1 U5821 ( .A(n4484), .ZN(n4483) );
  NAND2_X1 U5822 ( .A1(n7762), .A2(n4485), .ZN(n4484) );
  INV_X1 U5823 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5587) );
  OR2_X1 U5824 ( .A1(n4635), .A2(n4350), .ZN(n4299) );
  INV_X1 U5825 ( .A(n6945), .ZN(n4408) );
  NAND2_X1 U5826 ( .A1(n7667), .A2(n7776), .ZN(n4300) );
  NAND2_X1 U5827 ( .A1(n7690), .A2(n7675), .ZN(n4301) );
  NOR2_X1 U5828 ( .A1(n9183), .A2(n9208), .ZN(n4302) );
  INV_X1 U5829 ( .A(n8206), .ZN(n8198) );
  AND2_X1 U5830 ( .A1(n8169), .A2(n7723), .ZN(n8206) );
  NAND2_X1 U5831 ( .A1(n8309), .A2(n8310), .ZN(n8285) );
  INV_X1 U5832 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4823) );
  OR2_X1 U5833 ( .A1(n4479), .A2(n4483), .ZN(n4303) );
  XNOR2_X1 U5834 ( .A(n8355), .B(n8176), .ZN(n8155) );
  AND2_X1 U5835 ( .A1(n8633), .A2(n8634), .ZN(n8736) );
  INV_X1 U5836 ( .A(n9521), .ZN(n9294) );
  NAND2_X1 U5837 ( .A1(n5920), .A2(n5919), .ZN(n9521) );
  AND2_X1 U5838 ( .A1(n8160), .A2(n7825), .ZN(n8132) );
  AND2_X1 U5839 ( .A1(n5359), .A2(n4745), .ZN(n4304) );
  AND2_X1 U5840 ( .A1(n5311), .A2(n5310), .ZN(n8392) );
  INV_X1 U5841 ( .A(n8392), .ZN(n8276) );
  INV_X1 U5842 ( .A(n7435), .ZN(n9589) );
  NAND2_X1 U5843 ( .A1(n5902), .A2(n5901), .ZN(n7435) );
  OR2_X1 U5844 ( .A1(n9603), .A2(n7418), .ZN(n4305) );
  AND2_X1 U5845 ( .A1(n4893), .A2(n4913), .ZN(n4306) );
  AND2_X1 U5846 ( .A1(n4362), .A2(n6125), .ZN(n4307) );
  NOR2_X1 U5847 ( .A1(n4545), .A2(n4540), .ZN(n4539) );
  AND2_X1 U5848 ( .A1(n5152), .A2(n5134), .ZN(n4308) );
  AND2_X1 U5849 ( .A1(n4534), .A2(n4806), .ZN(n4309) );
  INV_X1 U5850 ( .A(n8989), .ZN(n4774) );
  AND2_X1 U5851 ( .A1(n4708), .A2(n8101), .ZN(n4310) );
  OR2_X1 U5852 ( .A1(n7464), .A2(n7693), .ZN(n4311) );
  AND2_X1 U5853 ( .A1(n4633), .A2(n8521), .ZN(n4632) );
  NAND2_X1 U5854 ( .A1(n7528), .A2(n4713), .ZN(n4712) );
  INV_X1 U5855 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4369) );
  NAND2_X1 U5856 ( .A1(n4706), .A2(n5093), .ZN(n8429) );
  INV_X1 U5857 ( .A(n8429), .ZN(n4705) );
  NAND2_X1 U5858 ( .A1(n7334), .A2(n5874), .ZN(n7378) );
  NOR2_X1 U5859 ( .A1(n9219), .A2(n9218), .ZN(n9217) );
  INV_X1 U5860 ( .A(n5398), .ZN(n4746) );
  AND4_X1 U5861 ( .A1(n5273), .A2(n5272), .A3(n5271), .A4(n5270), .ZN(n8097)
         );
  OR2_X1 U5862 ( .A1(n5428), .A2(n4572), .ZN(n4312) );
  INV_X1 U5863 ( .A(n9078), .ZN(n9035) );
  NAND2_X1 U5864 ( .A1(n5458), .A2(n5457), .ZN(n8355) );
  NAND2_X1 U5865 ( .A1(n7200), .A2(n7163), .ZN(n7364) );
  NAND2_X1 U5866 ( .A1(n5435), .A2(n5434), .ZN(n8362) );
  INV_X1 U5867 ( .A(n8362), .ZN(n8181) );
  NAND2_X1 U5868 ( .A1(n4374), .A2(n4377), .ZN(n8301) );
  NAND2_X1 U5869 ( .A1(n7582), .A2(n5238), .ZN(n7886) );
  AND2_X1 U5870 ( .A1(n7572), .A2(n7707), .ZN(n7803) );
  NAND2_X1 U5871 ( .A1(n4734), .A2(n5256), .ZN(n7922) );
  AND3_X1 U5872 ( .A1(n6257), .A2(n8571), .A3(n6256), .ZN(n4313) );
  NAND2_X1 U5873 ( .A1(n5961), .A2(n8580), .ZN(n8510) );
  NAND2_X1 U5874 ( .A1(n6237), .A2(n6236), .ZN(n9307) );
  INV_X1 U5875 ( .A(n9307), .ZN(n4513) );
  NAND2_X1 U5876 ( .A1(n7228), .A2(n5839), .ZN(n7333) );
  NAND2_X1 U5877 ( .A1(n7747), .A2(n7828), .ZN(n8115) );
  INV_X1 U5878 ( .A(n8115), .ZN(n4487) );
  NOR2_X1 U5879 ( .A1(n7545), .A2(n7546), .ZN(n4314) );
  AND2_X1 U5880 ( .A1(n5333), .A2(n5332), .ZN(n4315) );
  AND4_X1 U5881 ( .A1(n5253), .A2(n5252), .A3(n5251), .A4(n5250), .ZN(n7926)
         );
  INV_X1 U5882 ( .A(n8308), .ZN(n8402) );
  AND2_X1 U5883 ( .A1(n5265), .A2(n5264), .ZN(n8308) );
  NOR3_X1 U5884 ( .A1(n7324), .A2(n9514), .A3(n4522), .ZN(n4524) );
  NAND2_X1 U5885 ( .A1(n9236), .A2(n4515), .ZN(n4518) );
  NAND2_X1 U5886 ( .A1(n7378), .A2(n5895), .ZN(n7411) );
  INV_X1 U5887 ( .A(n4521), .ZN(n9287) );
  NOR2_X1 U5888 ( .A1(n7324), .A2(n4522), .ZN(n4521) );
  NAND2_X1 U5889 ( .A1(n8171), .A2(n7728), .ZN(n8188) );
  AND2_X1 U5890 ( .A1(n5996), .A2(n5995), .ZN(n4316) );
  NOR2_X1 U5891 ( .A1(n8303), .A2(n8402), .ZN(n4415) );
  AND2_X1 U5892 ( .A1(n5276), .A2(n5275), .ZN(n4317) );
  AND2_X1 U5893 ( .A1(n4486), .A2(n8158), .ZN(n4318) );
  NAND2_X1 U5894 ( .A1(n4352), .A2(n5570), .ZN(n4355) );
  INV_X1 U5895 ( .A(n4678), .ZN(n4677) );
  AOI21_X1 U5896 ( .B1(n8646), .B2(n9012), .A(n9014), .ZN(n4678) );
  AND2_X1 U5897 ( .A1(n4712), .A2(n4267), .ZN(n4319) );
  NAND2_X1 U5898 ( .A1(n6053), .A2(n6052), .ZN(n9483) );
  INV_X1 U5899 ( .A(n7754), .ZN(n4465) );
  AND2_X1 U5900 ( .A1(n7457), .A2(n7464), .ZN(n4320) );
  AND2_X1 U5901 ( .A1(n7457), .A2(n4423), .ZN(n4321) );
  NAND2_X1 U5902 ( .A1(n4779), .A2(n4291), .ZN(n7394) );
  NAND2_X1 U5903 ( .A1(n6952), .A2(n4419), .ZN(n4420) );
  NAND2_X1 U5904 ( .A1(n4750), .A2(n4752), .ZN(n7039) );
  OAI21_X1 U5905 ( .B1(n6911), .B2(n4279), .A(n6910), .ZN(n6946) );
  NAND2_X1 U5906 ( .A1(n4394), .A2(n7362), .ZN(n7450) );
  INV_X1 U5907 ( .A(n5592), .ZN(n6202) );
  AND3_X1 U5908 ( .A1(n5620), .A2(n5617), .A3(n4651), .ZN(n6324) );
  INV_X1 U5909 ( .A(n6324), .ZN(n6323) );
  INV_X1 U5910 ( .A(n9976), .ZN(n4416) );
  OAI21_X1 U5911 ( .B1(n9857), .B2(n4371), .A(n6711), .ZN(n6744) );
  INV_X1 U5912 ( .A(n9741), .ZN(n4520) );
  AND2_X1 U5913 ( .A1(n5631), .A2(n5630), .ZN(n6440) );
  INV_X1 U5914 ( .A(n9922), .ZN(n7761) );
  NAND2_X1 U5915 ( .A1(n7052), .A2(n7827), .ZN(n9922) );
  OR2_X1 U5916 ( .A1(n8967), .A2(n8966), .ZN(n4322) );
  AND2_X1 U5917 ( .A1(n7797), .A2(n9922), .ZN(n4323) );
  INV_X1 U5918 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4843) );
  INV_X1 U5919 ( .A(n8077), .ZN(n7839) );
  INV_X1 U5920 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4410) );
  INV_X1 U5921 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n4528) );
  INV_X1 U5922 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4719) );
  NAND2_X1 U5923 ( .A1(n5301), .A2(n5300), .ZN(n7859) );
  NAND2_X1 U5924 ( .A1(n4324), .A2(n4725), .ZN(n6764) );
  NAND3_X1 U5925 ( .A1(n4724), .A2(n6580), .A3(n4883), .ZN(n4324) );
  INV_X1 U5926 ( .A(n4727), .ZN(n4723) );
  NOR2_X1 U5927 ( .A1(n4855), .A2(n4854), .ZN(n4370) );
  NAND2_X2 U5928 ( .A1(n7916), .A2(n7915), .ZN(n7914) );
  INV_X1 U5929 ( .A(n8850), .ZN(n4646) );
  NAND2_X1 U5930 ( .A1(n4667), .A2(n4668), .ZN(n9077) );
  NOR2_X1 U5931 ( .A1(n9205), .A2(n8991), .ZN(n9204) );
  NAND2_X1 U5932 ( .A1(n4956), .A2(n4955), .ZN(n4972) );
  NAND2_X1 U5933 ( .A1(n4599), .A2(n4597), .ZN(n7447) );
  NAND2_X1 U5934 ( .A1(n4694), .A2(n4997), .ZN(n5016) );
  NAND2_X1 U5935 ( .A1(n6841), .A2(n8732), .ZN(n6995) );
  NAND2_X1 U5936 ( .A1(n4332), .A2(n8654), .ZN(n8656) );
  NAND2_X1 U5937 ( .A1(n8653), .A2(n4333), .ZN(n4332) );
  MUX2_X1 U5938 ( .A(n8659), .B(n8658), .S(n8705), .Z(n8662) );
  AND2_X2 U5939 ( .A1(n5592), .A2(n4790), .ZN(n5611) );
  AND2_X2 U5940 ( .A1(n4503), .A2(n5590), .ZN(n5592) );
  NAND2_X1 U5941 ( .A1(n4650), .A2(n8795), .ZN(n6867) );
  NAND3_X1 U5942 ( .A1(n8700), .A2(n9030), .A3(n8701), .ZN(n8703) );
  NAND2_X1 U5943 ( .A1(n4643), .A2(n8843), .ZN(n8847) );
  NAND2_X1 U5944 ( .A1(n4644), .A2(n8842), .ZN(n9720) );
  OAI21_X1 U5945 ( .B1(n8710), .B2(n4559), .A(n4557), .ZN(n8716) );
  OAI211_X1 U5946 ( .C1(n8705), .C2(n4340), .A(n4339), .B(n8667), .ZN(n8670)
         );
  OR2_X1 U5947 ( .A1(n4342), .A2(n5657), .ZN(n5658) );
  NAND2_X1 U5948 ( .A1(n6441), .A2(n5642), .ZN(n4342) );
  NAND2_X1 U5949 ( .A1(n5657), .A2(n4342), .ZN(n6568) );
  INV_X1 U5950 ( .A(n5681), .ZN(n4343) );
  NAND3_X1 U5951 ( .A1(n5961), .A2(n4632), .A3(n8580), .ZN(n4344) );
  INV_X1 U5952 ( .A(n5937), .ZN(n5932) );
  NAND2_X1 U5953 ( .A1(n5570), .A2(n4797), .ZN(n5875) );
  NAND4_X1 U5954 ( .A1(n5570), .A2(n4353), .A3(n4797), .A4(n5571), .ZN(n5962)
         );
  INV_X1 U5955 ( .A(n4355), .ZN(n5877) );
  NAND3_X1 U5956 ( .A1(n4272), .A2(n4363), .A3(n10060), .ZN(n4362) );
  NAND3_X1 U5957 ( .A1(n4272), .A2(n10060), .A3(n4358), .ZN(n4357) );
  AND2_X2 U5958 ( .A1(n4307), .A2(n4361), .ZN(n8504) );
  NAND2_X1 U5959 ( .A1(n4361), .A2(n4362), .ZN(n8532) );
  NAND3_X1 U5960 ( .A1(n4272), .A2(n10060), .A3(n6104), .ZN(n8529) );
  OAI21_X1 U5961 ( .B1(n5580), .B2(n4368), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5582) );
  INV_X1 U5962 ( .A(n4365), .ZN(n5576) );
  NOR2_X2 U5963 ( .A1(n5505), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4855) );
  NAND2_X1 U5964 ( .A1(n4373), .A2(n4375), .ZN(n4707) );
  NAND2_X1 U5965 ( .A1(n7528), .A2(n4377), .ZN(n4373) );
  INV_X1 U5966 ( .A(n4380), .ZN(n8222) );
  INV_X1 U5967 ( .A(n8240), .ZN(n4387) );
  NAND2_X1 U5968 ( .A1(n7200), .A2(n4395), .ZN(n4393) );
  NAND2_X1 U5969 ( .A1(n4405), .A2(n4404), .ZN(n6960) );
  OAI211_X1 U5970 ( .C1(n4405), .C2(n4400), .A(n4403), .B(n6961), .ZN(n6964)
         );
  OAI21_X2 U5971 ( .B1(n4880), .B2(n4410), .A(n4409), .ZN(n6917) );
  INV_X1 U5972 ( .A(n8303), .ZN(n4411) );
  NAND2_X1 U5973 ( .A1(n4412), .A2(n4411), .ZN(n8251) );
  INV_X1 U5974 ( .A(n4415), .ZN(n8302) );
  AND2_X1 U5975 ( .A1(n8177), .A2(n4428), .ZN(n8139) );
  NAND2_X1 U5976 ( .A1(n8177), .A2(n4429), .ZN(n8123) );
  NAND2_X2 U5977 ( .A1(n4817), .A2(n4261), .ZN(n5505) );
  INV_X2 U5978 ( .A(n5220), .ZN(n4817) );
  OAI21_X1 U5979 ( .B1(n7503), .B2(n4436), .A(n4435), .ZN(n8939) );
  MUX2_X1 U5980 ( .A(n6277), .B(P1_REG2_REG_1__SCAN_IN), .S(n6351), .Z(n8905)
         );
  NAND2_X1 U5981 ( .A1(n7715), .A2(n8286), .ZN(n7716) );
  NAND2_X1 U5982 ( .A1(n4455), .A2(n4453), .ZN(n4452) );
  OR2_X1 U5983 ( .A1(n7711), .A2(n7710), .ZN(n4455) );
  INV_X1 U5984 ( .A(n7760), .ZN(n4467) );
  OAI21_X1 U5985 ( .B1(n4467), .B2(n7798), .A(n4266), .ZN(n4470) );
  NAND3_X1 U5986 ( .A1(n4471), .A2(n4470), .A3(n4468), .ZN(P2_U3244) );
  NAND3_X1 U5987 ( .A1(n7760), .A2(n7224), .A3(n4270), .ZN(n4471) );
  OR2_X1 U5988 ( .A1(n7738), .A2(n4476), .ZN(n4475) );
  INV_X1 U5989 ( .A(n8158), .ZN(n4482) );
  NAND4_X1 U5990 ( .A1(n7689), .A2(n7754), .A3(n7688), .A4(n4492), .ZN(n4491)
         );
  NAND2_X4 U5991 ( .A1(n5668), .A2(n8594), .ZN(n8608) );
  XNOR2_X1 U5992 ( .A(n5627), .B(n5626), .ZN(n6280) );
  XNOR2_X2 U5993 ( .A(n5625), .B(P1_IR_REG_28__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U5994 ( .A1(n4502), .A2(n4503), .ZN(n4680) );
  AND2_X1 U5995 ( .A1(n4681), .A2(n5590), .ZN(n4502) );
  AND2_X1 U5996 ( .A1(n9084), .A2(n4510), .ZN(n9052) );
  NAND2_X1 U5997 ( .A1(n9084), .A2(n4511), .ZN(n9041) );
  NAND2_X1 U5998 ( .A1(n9084), .A2(n4507), .ZN(n4506) );
  NAND2_X1 U5999 ( .A1(n9084), .A2(n9075), .ZN(n9070) );
  NAND3_X1 U6000 ( .A1(n4508), .A2(n4506), .A3(n4504), .ZN(n9582) );
  INV_X1 U6001 ( .A(n4518), .ZN(n9179) );
  INV_X1 U6002 ( .A(n4524), .ZN(n9271) );
  NAND3_X1 U6003 ( .A1(n4693), .A2(n4309), .A3(n4692), .ZN(n4533) );
  NAND3_X1 U6004 ( .A1(n4693), .A2(n4692), .A3(n4534), .ZN(n4530) );
  NAND2_X1 U6005 ( .A1(n5188), .A2(n4539), .ZN(n4535) );
  NAND2_X1 U6006 ( .A1(n5088), .A2(n4551), .ZN(n4548) );
  NAND2_X1 U6007 ( .A1(n4548), .A2(n4549), .ZN(n5161) );
  NAND2_X1 U6008 ( .A1(n5088), .A2(n4555), .ZN(n4554) );
  OAI21_X1 U6009 ( .B1(n5304), .B2(n5303), .A(n5305), .ZN(n5321) );
  NAND2_X1 U6010 ( .A1(n5373), .A2(n5372), .ZN(n5408) );
  NAND2_X1 U6011 ( .A1(n5282), .A2(n5281), .ZN(n5304) );
  OAI21_X1 U6012 ( .B1(n4994), .B2(n4697), .A(n5015), .ZN(n4696) );
  INV_X1 U6013 ( .A(n4696), .ZN(n4695) );
  NAND2_X1 U6014 ( .A1(n5371), .A2(n5370), .ZN(n5373) );
  NAND3_X1 U6015 ( .A1(n4808), .A2(n4810), .A3(n4729), .ZN(n4576) );
  NAND2_X1 U6016 ( .A1(n5021), .A2(n4815), .ZN(n5220) );
  NOR2_X2 U6017 ( .A1(n4576), .A2(n4730), .ZN(n5021) );
  NAND2_X1 U6018 ( .A1(n4809), .A2(n4859), .ZN(n4730) );
  INV_X1 U6019 ( .A(n6593), .ZN(n6594) );
  INV_X1 U6020 ( .A(n4582), .ZN(n6969) );
  NAND2_X1 U6021 ( .A1(n7467), .A2(n7697), .ZN(n7484) );
  NAND2_X1 U6022 ( .A1(n7467), .A2(n4584), .ZN(n4583) );
  NAND3_X1 U6023 ( .A1(n4590), .A2(n4588), .A3(n7639), .ZN(n6746) );
  NAND3_X1 U6024 ( .A1(n7634), .A2(n6729), .A3(n6728), .ZN(n4590) );
  NAND2_X1 U6025 ( .A1(n4591), .A2(n4594), .ZN(n7811) );
  NAND2_X1 U6026 ( .A1(n8309), .A2(n4592), .ZN(n4591) );
  NAND2_X1 U6027 ( .A1(n7199), .A2(n4600), .ZN(n4599) );
  NAND2_X1 U6028 ( .A1(n4848), .A2(n4610), .ZN(n4825) );
  NAND2_X1 U6029 ( .A1(n4848), .A2(n4269), .ZN(n8458) );
  NAND2_X1 U6030 ( .A1(n7227), .A2(n5839), .ZN(n4613) );
  NAND3_X1 U6031 ( .A1(n8557), .A2(n6017), .A3(n4622), .ZN(n4621) );
  NAND3_X1 U6032 ( .A1(n8557), .A2(n6017), .A3(n4614), .ZN(n4618) );
  NAND2_X1 U6033 ( .A1(n4621), .A2(n4620), .ZN(n8540) );
  NAND2_X1 U6034 ( .A1(n8557), .A2(n6017), .ZN(n8489) );
  INV_X1 U6035 ( .A(n8490), .ZN(n4622) );
  OAI21_X1 U6036 ( .B1(n6070), .B2(n4625), .A(n4623), .ZN(n8480) );
  NAND2_X1 U6038 ( .A1(n6070), .A2(n4630), .ZN(n4626) );
  NAND2_X1 U6039 ( .A1(n8504), .A2(n4640), .ZN(n4639) );
  INV_X1 U6040 ( .A(n9720), .ZN(n4643) );
  NAND2_X1 U6041 ( .A1(n6820), .A2(n6819), .ZN(n4644) );
  OAI21_X1 U6042 ( .B1(n6879), .B2(n4648), .A(n4645), .ZN(n6841) );
  NAND2_X1 U6043 ( .A1(n9749), .A2(n6325), .ZN(n8725) );
  INV_X2 U6044 ( .A(n6322), .ZN(n8900) );
  AND3_X2 U6045 ( .A1(n4652), .A2(n5645), .A3(n5647), .ZN(n6322) );
  AND2_X1 U6046 ( .A1(n5646), .A2(n5644), .ZN(n4652) );
  NAND2_X1 U6047 ( .A1(n9204), .A2(n4657), .ZN(n4656) );
  INV_X1 U6048 ( .A(n4660), .ZN(n9185) );
  INV_X1 U6049 ( .A(n9103), .ZN(n4661) );
  OAI21_X1 U6050 ( .B1(n4664), .B2(n4661), .A(n4662), .ZN(n9057) );
  NAND2_X1 U6051 ( .A1(n9103), .A2(n4670), .ZN(n4667) );
  NOR2_X1 U6052 ( .A1(n9058), .A2(n9059), .ZN(n4673) );
  OAI21_X1 U6053 ( .B1(n9103), .B2(n4672), .A(n9027), .ZN(n9088) );
  NAND2_X1 U6054 ( .A1(n9262), .A2(n8646), .ZN(n4676) );
  INV_X1 U6055 ( .A(n4679), .ZN(n9250) );
  NAND2_X1 U6056 ( .A1(n5592), .A2(n5591), .ZN(n5597) );
  NAND2_X1 U6057 ( .A1(n7451), .A2(n4684), .ZN(n4683) );
  NAND2_X1 U6058 ( .A1(n4688), .A2(n4689), .ZN(n8113) );
  NAND2_X1 U6059 ( .A1(n8147), .A2(n4256), .ZN(n4688) );
  NAND2_X1 U6060 ( .A1(n8147), .A2(n8155), .ZN(n8146) );
  NAND2_X1 U6061 ( .A1(n4995), .A2(n4695), .ZN(n4693) );
  NAND2_X1 U6062 ( .A1(n4995), .A2(n4994), .ZN(n4694) );
  INV_X1 U6063 ( .A(n4997), .ZN(n4697) );
  INV_X1 U6064 ( .A(n4699), .ZN(n4701) );
  OAI21_X1 U6065 ( .B1(n4910), .B2(n4700), .A(n4928), .ZN(n4699) );
  INV_X1 U6066 ( .A(n4913), .ZN(n4700) );
  NAND2_X1 U6067 ( .A1(n4894), .A2(n4893), .ZN(n4911) );
  NAND2_X1 U6068 ( .A1(n4702), .A2(n4701), .ZN(n4933) );
  NAND2_X1 U6069 ( .A1(n4894), .A2(n4306), .ZN(n4702) );
  NAND2_X1 U6070 ( .A1(n4707), .A2(n4310), .ZN(n8280) );
  INV_X1 U6071 ( .A(n8100), .ZN(n4711) );
  NAND2_X1 U6072 ( .A1(n7528), .A2(n7527), .ZN(n7529) );
  INV_X1 U6073 ( .A(n4712), .ZN(n7575) );
  INV_X1 U6074 ( .A(n7527), .ZN(n4714) );
  NAND3_X1 U6075 ( .A1(n4717), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4715) );
  NAND3_X1 U6076 ( .A1(n4719), .A2(n4720), .A3(n4718), .ZN(n4716) );
  NAND2_X1 U6077 ( .A1(n4725), .A2(n4721), .ZN(n6616) );
  NAND2_X1 U6078 ( .A1(n4727), .A2(n4726), .ZN(n4721) );
  INV_X1 U6079 ( .A(n6616), .ZN(n4724) );
  NAND2_X2 U6080 ( .A1(n4882), .A2(n4881), .ZN(n6580) );
  NAND2_X1 U6081 ( .A1(n6764), .A2(n6765), .ZN(n4919) );
  NAND2_X1 U6082 ( .A1(n6580), .A2(n4883), .ZN(n6617) );
  NAND2_X1 U6083 ( .A1(n4248), .A2(n4250), .ZN(n4726) );
  NAND2_X1 U6084 ( .A1(n4808), .A2(n4810), .ZN(n4728) );
  NAND3_X1 U6085 ( .A1(n4809), .A2(n4860), .A3(n4808), .ZN(n4976) );
  NAND2_X1 U6086 ( .A1(n7215), .A2(n4308), .ZN(n5158) );
  NAND2_X2 U6087 ( .A1(n7217), .A2(n7216), .ZN(n7215) );
  NAND2_X1 U6088 ( .A1(n7914), .A2(n4304), .ZN(n4804) );
  INV_X1 U6089 ( .A(n6772), .ZN(n4747) );
  INV_X1 U6090 ( .A(n6888), .ZN(n4768) );
  NAND3_X1 U6091 ( .A1(n9737), .A2(n6326), .A3(n6327), .ZN(n6816) );
  NAND2_X1 U6092 ( .A1(n4778), .A2(n4777), .ZN(n9004) );
  NAND2_X1 U6093 ( .A1(n7327), .A2(n4305), .ZN(n4779) );
  AOI21_X2 U6094 ( .B1(n9191), .B2(n4783), .A(n4782), .ZN(n9143) );
  NAND4_X1 U6095 ( .A1(n5669), .A2(n4788), .A3(n5565), .A4(n5566), .ZN(n5756)
         );
  NOR2_X2 U6096 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4788) );
  NOR2_X4 U6097 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5669) );
  INV_X1 U6098 ( .A(n8118), .ZN(n7835) );
  AOI21_X1 U6099 ( .B1(n8763), .B2(n8762), .A(n8761), .ZN(n8886) );
  NAND2_X1 U6100 ( .A1(n5663), .A2(n5662), .ZN(n6484) );
  NAND2_X1 U6101 ( .A1(n5820), .A2(n5819), .ZN(n7145) );
  XNOR2_X1 U6102 ( .A(n7607), .B(SI_30_), .ZN(n8595) );
  OR2_X1 U6103 ( .A1(n9305), .A2(n9524), .ZN(n9310) );
  XNOR2_X1 U6104 ( .A(n5429), .B(n5428), .ZN(n7477) );
  NOR2_X2 U6105 ( .A1(n9253), .A2(n9504), .ZN(n9236) );
  NAND2_X1 U6106 ( .A1(n4839), .A2(n4838), .ZN(n5502) );
  INV_X1 U6107 ( .A(n4840), .ZN(n4839) );
  OR2_X1 U6108 ( .A1(n4903), .A2(n4885), .ZN(n4886) );
  NAND2_X1 U6109 ( .A1(n7159), .A2(n7158), .ZN(n7202) );
  XNOR2_X1 U6110 ( .A(n9929), .B(n4902), .ZN(n4868) );
  INV_X1 U6111 ( .A(n5817), .ZN(n5820) );
  NOR2_X2 U6112 ( .A1(n9263), .A2(n9264), .ZN(n9262) );
  NOR2_X1 U6113 ( .A1(n6015), .A2(n6014), .ZN(n6016) );
  INV_X1 U6114 ( .A(n6705), .ZN(n6704) );
  INV_X1 U6115 ( .A(n4829), .ZN(n8468) );
  INV_X1 U6116 ( .A(n5687), .ZN(n6247) );
  NAND2_X1 U6117 ( .A1(n6594), .A2(n6917), .ZN(n6916) );
  INV_X1 U6118 ( .A(n9192), .ZN(n9193) );
  NOR2_X2 U6119 ( .A1(n5403), .A2(n5402), .ZN(n7877) );
  BUF_X4 U6120 ( .A(n4902), .Z(n5415) );
  NOR2_X1 U6121 ( .A1(n9057), .A2(n9032), .ZN(n9034) );
  XNOR2_X2 U6122 ( .A(n5397), .B(n4746), .ZN(n7853) );
  NAND2_X2 U6123 ( .A1(n4831), .A2(n8468), .ZN(n6392) );
  INV_X1 U6124 ( .A(n4831), .ZN(n7596) );
  INV_X1 U6125 ( .A(n6281), .ZN(n8975) );
  INV_X1 U6126 ( .A(n6280), .ZN(n6281) );
  AND2_X1 U6127 ( .A1(n8424), .A2(n7693), .ZN(n4795) );
  NAND2_X2 U6128 ( .A1(n6844), .A2(n9222), .ZN(n9762) );
  INV_X1 U6129 ( .A(n9762), .ZN(n9234) );
  INV_X1 U6130 ( .A(n5639), .ZN(n6206) );
  AND4_X1 U6131 ( .A1(n5569), .A2(n5568), .A3(n5800), .A4(n5567), .ZN(n4797)
         );
  OR2_X1 U6132 ( .A1(n9075), .A2(n8578), .ZN(n4800) );
  OR2_X1 U6133 ( .A1(n8111), .A2(n7945), .ZN(n4801) );
  AND2_X1 U6134 ( .A1(n5626), .A2(n5610), .ZN(n4803) );
  INV_X1 U6135 ( .A(n4895), .ZN(n5111) );
  INV_X1 U6136 ( .A(n7052), .ZN(n5533) );
  AND2_X1 U6137 ( .A1(n5160), .A2(n5141), .ZN(n4805) );
  INV_X1 U6138 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5094) );
  AND2_X1 U6139 ( .A1(n5062), .A2(n5042), .ZN(n4806) );
  NAND2_X1 U6140 ( .A1(n8217), .A2(n7816), .ZN(n8168) );
  INV_X1 U6141 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5610) );
  NAND2_X1 U6142 ( .A1(n6115), .A2(n6114), .ZN(n9127) );
  OR2_X1 U6143 ( .A1(n8718), .A2(n6209), .ZN(n9724) );
  OR2_X1 U6144 ( .A1(n8251), .A2(n8380), .ZN(n4807) );
  INV_X1 U6145 ( .A(n9030), .ZN(n9058) );
  AND2_X1 U6146 ( .A1(n7697), .A2(n7696), .ZN(n7698) );
  INV_X1 U6147 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5567) );
  INV_X1 U6148 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4810) );
  INV_X1 U6149 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U6150 ( .A1(n7899), .A2(n7946), .ZN(n5395) );
  INV_X1 U6151 ( .A(n6351), .ZN(n5651) );
  INV_X1 U6152 ( .A(n5648), .ZN(n5844) );
  INV_X1 U6153 ( .A(n9127), .ZN(n8996) );
  INV_X1 U6154 ( .A(n8736), .ZN(n7130) );
  INV_X1 U6155 ( .A(n5123), .ZN(n5121) );
  NAND2_X1 U6156 ( .A1(n7797), .A2(n4865), .ZN(n4867) );
  INV_X1 U6157 ( .A(n5385), .ZN(n5377) );
  AND2_X1 U6158 ( .A1(n4960), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n4980) );
  INV_X1 U6159 ( .A(n8329), .ZN(n6728) );
  NAND2_X1 U6160 ( .A1(n6704), .A2(n9929), .ZN(n6727) );
  AOI21_X1 U6161 ( .B1(n8470), .B2(n8473), .A(n5938), .ZN(n5957) );
  INV_X1 U6162 ( .A(n6091), .ZN(n6089) );
  NAND2_X1 U6163 ( .A1(n9114), .A2(n8996), .ZN(n8997) );
  INV_X1 U6164 ( .A(n6023), .ZN(n6021) );
  AND2_X1 U6165 ( .A1(n9479), .A2(n9167), .ZN(n8993) );
  NAND2_X1 U6166 ( .A1(n7131), .A2(n7130), .ZN(n7177) );
  INV_X1 U6167 ( .A(n8727), .ZN(n6852) );
  INV_X1 U6168 ( .A(SI_13_), .ZN(n5138) );
  INV_X1 U6169 ( .A(SI_8_), .ZN(n9346) );
  OR2_X1 U6170 ( .A1(n5168), .A2(n5167), .ZN(n5201) );
  INV_X1 U6171 ( .A(n6756), .ZN(n4946) );
  OR2_X1 U6172 ( .A1(n5348), .A2(n5347), .ZN(n5385) );
  NAND2_X1 U6173 ( .A1(n5266), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U6174 ( .A1(n5377), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U6175 ( .A1(n5312), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5348) );
  NOR2_X1 U6176 ( .A1(n8114), .A2(n8115), .ZN(n8118) );
  OR2_X1 U6177 ( .A1(n5095), .A2(n5094), .ZN(n5123) );
  INV_X1 U6178 ( .A(n8434), .ZN(n7171) );
  OR2_X1 U6179 ( .A1(n7772), .A2(n6909), .ZN(n6910) );
  INV_X1 U6180 ( .A(n5923), .ZN(n5921) );
  INV_X1 U6181 ( .A(n5818), .ZN(n5819) );
  OR2_X1 U6182 ( .A1(n8567), .A2(n8568), .ZN(n6159) );
  NAND2_X1 U6183 ( .A1(n6129), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6144) );
  OR2_X1 U6184 ( .A1(n6055), .A2(n6054), .ZN(n6074) );
  OR2_X1 U6185 ( .A1(n5904), .A2(n5903), .ZN(n5923) );
  NOR2_X1 U6186 ( .A1(n9037), .A2(n9036), .ZN(n9038) );
  AND2_X1 U6187 ( .A1(n7182), .A2(n7181), .ZN(n7183) );
  INV_X1 U6188 ( .A(n6327), .ZN(n8726) );
  NAND2_X1 U6189 ( .A1(n7598), .A2(n7597), .ZN(n7602) );
  NAND2_X1 U6190 ( .A1(n5114), .A2(n5113), .ZN(n5135) );
  NAND2_X1 U6191 ( .A1(n5369), .A2(n5368), .ZN(n7627) );
  INV_X1 U6192 ( .A(n7958), .ZN(n6758) );
  OR2_X1 U6193 ( .A1(n5436), .A2(n7937), .ZN(n5461) );
  OR2_X1 U6194 ( .A1(n7864), .A2(n9863), .ZN(n7938) );
  INV_X1 U6195 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5531) );
  OR2_X1 U6196 ( .A1(n8152), .A2(n5419), .ZN(n5468) );
  INV_X1 U6197 ( .A(n8371), .ZN(n8205) );
  AND2_X1 U6198 ( .A1(n8402), .A2(n8099), .ZN(n8100) );
  AND2_X1 U6199 ( .A1(n7761), .A2(n5543), .ZN(n9954) );
  INV_X1 U6200 ( .A(n5557), .ZN(n6560) );
  AND2_X1 U6201 ( .A1(n6182), .A2(n6183), .ZN(n5599) );
  NAND2_X1 U6202 ( .A1(n5921), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5946) );
  OR2_X1 U6203 ( .A1(n5845), .A2(n7337), .ZN(n5861) );
  AND2_X1 U6204 ( .A1(n6163), .A2(n6162), .ZN(n6178) );
  OR2_X1 U6205 ( .A1(n5984), .A2(n8523), .ZN(n6005) );
  OR2_X1 U6206 ( .A1(n6108), .A2(n6107), .ZN(n6131) );
  INV_X1 U6207 ( .A(n9090), .ZN(n9007) );
  INV_X1 U6208 ( .A(n8552), .ZN(n8588) );
  AND2_X1 U6209 ( .A1(n8877), .A2(n5638), .ZN(n8875) );
  CLKBUF_X3 U6210 ( .A(n5711), .Z(n8599) );
  INV_X1 U6211 ( .A(n6381), .ZN(n9661) );
  INV_X1 U6212 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7337) );
  INV_X1 U6213 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7505) );
  INV_X1 U6214 ( .A(n8771), .ZN(n9299) );
  OR2_X1 U6215 ( .A1(n9473), .A2(n9121), .ZN(n8995) );
  INV_X1 U6216 ( .A(n9168), .ZN(n9208) );
  INV_X1 U6217 ( .A(n9214), .ZN(n9252) );
  INV_X1 U6218 ( .A(n8988), .ZN(n9264) );
  INV_X1 U6219 ( .A(n6469), .ZN(n6467) );
  AND2_X1 U6220 ( .A1(n6321), .A2(n6320), .ZN(n9751) );
  NAND2_X1 U6221 ( .A1(n5639), .A2(n8753), .ZN(n6469) );
  OAI22_X1 U6222 ( .A1(n6916), .A2(n5489), .B1(n6917), .B2(n5415), .ZN(n6582)
         );
  AND2_X1 U6223 ( .A1(n5384), .A2(n5383), .ZN(n7946) );
  AND4_X1 U6224 ( .A1(n5174), .A2(n5173), .A3(n5172), .A4(n5171), .ZN(n7517)
         );
  AND2_X1 U6225 ( .A1(n6558), .A2(n6557), .ZN(n9845) );
  AND2_X1 U6226 ( .A1(n6561), .A2(n6560), .ZN(n9556) );
  AND2_X1 U6227 ( .A1(n6532), .A2(n5557), .ZN(n8312) );
  OR2_X1 U6228 ( .A1(n7364), .A2(n7778), .ZN(n7345) );
  INV_X1 U6229 ( .A(n8292), .ZN(n9865) );
  AND2_X1 U6230 ( .A1(n6714), .A2(n7846), .ZN(n7065) );
  INV_X1 U6231 ( .A(n9946), .ZN(n9985) );
  AND2_X1 U6232 ( .A1(n8316), .A2(n8315), .ZN(n8405) );
  INV_X1 U6233 ( .A(n9989), .ZN(n9957) );
  NAND2_X1 U6234 ( .A1(n9854), .A2(n9967), .ZN(n9989) );
  OR2_X1 U6235 ( .A1(n6530), .A2(n9918), .ZN(n9882) );
  INV_X1 U6236 ( .A(n6271), .ZN(n9918) );
  AND2_X1 U6237 ( .A1(n6227), .A2(n6209), .ZN(n8552) );
  INV_X1 U6238 ( .A(n8578), .ZN(n8590) );
  OR2_X1 U6239 ( .A1(n9054), .A2(n6247), .ZN(n6220) );
  INV_X1 U6240 ( .A(n5686), .ZN(n6217) );
  AND2_X1 U6241 ( .A1(n8965), .A2(n6282), .ZN(n9697) );
  AND2_X1 U6242 ( .A1(n8965), .A2(n6303), .ZN(n9699) );
  INV_X1 U6243 ( .A(n9699), .ZN(n9687) );
  INV_X1 U6244 ( .A(n5638), .ZN(n9744) );
  OAI21_X1 U6245 ( .B1(n9040), .B2(n9751), .A(n9039), .ZN(n9302) );
  AND2_X1 U6246 ( .A1(n9211), .A2(n9015), .ZN(n9241) );
  INV_X1 U6247 ( .A(n9724), .ZN(n9739) );
  AND2_X1 U6248 ( .A1(n6467), .A2(n8877), .ZN(n9742) );
  NAND2_X1 U6249 ( .A1(n9759), .A2(n9587), .ZN(n9815) );
  INV_X1 U6250 ( .A(n9587), .ZN(n9822) );
  INV_X1 U6251 ( .A(n6472), .ZN(n6466) );
  XNOR2_X1 U6252 ( .A(n5598), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6183) );
  AND2_X1 U6253 ( .A1(n5878), .A2(n4355), .ZN(n8934) );
  INV_X1 U6254 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9395) );
  AND2_X1 U6255 ( .A1(n6404), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6271) );
  AND2_X1 U6256 ( .A1(n5561), .A2(n5560), .ZN(n5562) );
  INV_X1 U6257 ( .A(n7929), .ZN(n7945) );
  INV_X1 U6258 ( .A(n7933), .ZN(n7931) );
  INV_X1 U6259 ( .A(n7872), .ZN(n8261) );
  INV_X1 U6260 ( .A(n9556), .ZN(n9847) );
  AND2_X1 U6261 ( .A1(n7487), .A2(n7486), .ZN(n8422) );
  NAND2_X1 U6262 ( .A1(n8336), .A2(n6720), .ZN(n8321) );
  NAND2_X2 U6263 ( .A1(n6721), .A2(n8272), .ZN(n8336) );
  INV_X1 U6264 ( .A(n10008), .ZN(n10006) );
  INV_X1 U6265 ( .A(n9993), .ZN(n9991) );
  NOR2_X1 U6266 ( .A1(n9883), .A2(n9882), .ZN(n9898) );
  CLKBUF_X1 U6267 ( .A(n9898), .Z(n9919) );
  INV_X1 U6268 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9428) );
  INV_X1 U6269 ( .A(n8461), .ZN(n8465) );
  AND2_X1 U6270 ( .A1(n6226), .A2(n6478), .ZN(n8563) );
  INV_X1 U6271 ( .A(n6875), .ZN(n9804) );
  NAND2_X1 U6272 ( .A1(n6220), .A2(n6219), .ZN(n9078) );
  OR2_X1 U6273 ( .A1(P1_U3083), .A2(n6448), .ZN(n9689) );
  NAND2_X1 U6274 ( .A1(n9762), .A2(n6225), .ZN(n9733) );
  AND2_X1 U6275 ( .A1(n7101), .A2(n7100), .ZN(n9825) );
  INV_X1 U6276 ( .A(n9843), .ZN(n9840) );
  AND2_X2 U6277 ( .A1(n6473), .A2(n6472), .ZN(n9843) );
  AND2_X1 U6278 ( .A1(n9601), .A2(n9600), .ZN(n9614) );
  AND2_X1 U6279 ( .A1(n9825), .A2(n9824), .ZN(n9842) );
  INV_X1 U6280 ( .A(n9828), .ZN(n9826) );
  OR2_X1 U6281 ( .A1(n9765), .A2(n9764), .ZN(n9771) );
  INV_X1 U6282 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7483) );
  INV_X1 U6283 ( .A(n4246), .ZN(n8753) );
  INV_X1 U6284 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6590) );
  INV_X1 U6285 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6400) );
  NOR2_X1 U6286 ( .A1(n10051), .A2(n10050), .ZN(n10049) );
  AND2_X1 U6287 ( .A1(n6530), .A2(n6271), .ZN(P2_U3966) );
  NOR2_X2 U6288 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4809) );
  NOR2_X2 U6289 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4808) );
  INV_X1 U6290 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4819) );
  INV_X1 U6291 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4818) );
  NOR2_X1 U6292 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n4821) );
  NOR2_X1 U6293 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5500) );
  NOR2_X1 U6294 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n4820) );
  INV_X1 U6296 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n4827) );
  OR2_X1 U6297 ( .A1(n4904), .A2(n4827), .ZN(n4835) );
  INV_X1 U6298 ( .A(n6392), .ZN(n4828) );
  NAND2_X1 U6299 ( .A1(n4828), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4834) );
  NAND2_X2 U6300 ( .A1(n7596), .A2(n4829), .ZN(n4903) );
  INV_X1 U6301 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n4830) );
  OR2_X1 U6302 ( .A1(n4903), .A2(n4830), .ZN(n4833) );
  NAND2_X1 U6303 ( .A1(n4873), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n4832) );
  AND4_X2 U6304 ( .A1(n4835), .A2(n4834), .A3(n4833), .A4(n4832), .ZN(n6705)
         );
  NOR2_X2 U6305 ( .A1(n4836), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n4842) );
  NAND2_X1 U6306 ( .A1(n4842), .A2(n4837), .ZN(n4840) );
  XNOR2_X2 U6307 ( .A(n5513), .B(n5512), .ZN(n7052) );
  NAND2_X1 U6308 ( .A1(n4840), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4841) );
  NAND2_X1 U6309 ( .A1(n4847), .A2(n4843), .ZN(n4844) );
  INV_X1 U6310 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4845) );
  XNOR2_X2 U6311 ( .A(n4847), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8077) );
  AND2_X4 U6312 ( .A1(n7761), .A2(n7845), .ZN(n5489) );
  OR2_X1 U6313 ( .A1(n6705), .A2(n5489), .ZN(n4869) );
  NAND2_X1 U6314 ( .A1(n5505), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4849) );
  NAND2_X1 U6315 ( .A1(n4849), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4851) );
  INV_X1 U6316 ( .A(n4855), .ZN(n4852) );
  INV_X1 U6317 ( .A(n7613), .ZN(n8594) );
  MUX2_X1 U6318 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(P2_DATAO_REG_0__SCAN_IN), 
        .S(n4895), .Z(n4857) );
  XNOR2_X1 U6319 ( .A(n4891), .B(SI_1_), .ZN(n4889) );
  MUX2_X1 U6320 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4895), .Z(n4890) );
  XNOR2_X1 U6321 ( .A(n4889), .B(n4890), .ZN(n6354) );
  NAND2_X1 U6322 ( .A1(n4958), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4864) );
  INV_X1 U6323 ( .A(n4880), .ZN(n4941) );
  NAND2_X1 U6324 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4858) );
  MUX2_X1 U6325 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4858), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n4862) );
  INV_X1 U6326 ( .A(n4860), .ZN(n4861) );
  NAND2_X1 U6327 ( .A1(n4862), .A2(n4861), .ZN(n6536) );
  INV_X1 U6328 ( .A(n6536), .ZN(n7965) );
  NAND2_X1 U6329 ( .A1(n4941), .A2(n7965), .ZN(n4863) );
  OAI211_X2 U6330 ( .C1(n4957), .C2(n6354), .A(n4864), .B(n4863), .ZN(n6584)
         );
  INV_X2 U6331 ( .A(n6584), .ZN(n9929) );
  NAND2_X1 U6332 ( .A1(n4866), .A2(n7799), .ZN(n6719) );
  NAND2_X1 U6333 ( .A1(n4869), .A2(n4868), .ZN(n4883) );
  INV_X1 U6334 ( .A(n4868), .ZN(n4871) );
  INV_X1 U6335 ( .A(n4869), .ZN(n4870) );
  NAND2_X1 U6336 ( .A1(n4871), .A2(n4870), .ZN(n4872) );
  NAND2_X1 U6337 ( .A1(n4883), .A2(n4872), .ZN(n6583) );
  INV_X1 U6338 ( .A(n6583), .ZN(n4882) );
  INV_X2 U6339 ( .A(n4873), .ZN(n5419) );
  INV_X1 U6340 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6600) );
  OR2_X1 U6341 ( .A1(n5419), .A2(n6600), .ZN(n4878) );
  NAND2_X1 U6342 ( .A1(n5420), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n4877) );
  INV_X1 U6343 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9994) );
  OR2_X1 U6344 ( .A1(n4903), .A2(n9994), .ZN(n4876) );
  INV_X1 U6345 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n4874) );
  OR2_X1 U6346 ( .A1(n6392), .A2(n4874), .ZN(n4875) );
  NAND2_X1 U6347 ( .A1(n8594), .A2(SI_0_), .ZN(n4879) );
  XNOR2_X1 U6348 ( .A(n4879), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8469) );
  INV_X1 U6349 ( .A(n6582), .ZN(n4881) );
  INV_X1 U6350 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9394) );
  INV_X1 U6351 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6513) );
  INV_X1 U6352 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n4884) );
  OR2_X1 U6353 ( .A1(n4904), .A2(n4884), .ZN(n4887) );
  INV_X1 U6354 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n4885) );
  AND4_X2 U6355 ( .A1(n4796), .A2(n4888), .A3(n4887), .A4(n4886), .ZN(n6708)
         );
  NAND2_X1 U6356 ( .A1(n4890), .A2(n4889), .ZN(n4894) );
  INV_X1 U6357 ( .A(n4891), .ZN(n4892) );
  NAND2_X1 U6358 ( .A1(n4892), .A2(SI_1_), .ZN(n4893) );
  MUX2_X1 U6359 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4895), .Z(n4912) );
  INV_X1 U6360 ( .A(SI_2_), .ZN(n4896) );
  XNOR2_X1 U6361 ( .A(n4911), .B(n4910), .ZN(n6359) );
  NAND2_X1 U6362 ( .A1(n4958), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4901) );
  NOR2_X1 U6363 ( .A1(n4860), .A2(n4854), .ZN(n4897) );
  INV_X1 U6364 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4898) );
  MUX2_X1 U6365 ( .A(n4854), .B(n4897), .S(P2_IR_REG_2__SCAN_IN), .Z(n4899) );
  AND2_X1 U6366 ( .A1(n4860), .A2(n4898), .ZN(n4935) );
  NOR2_X1 U6367 ( .A1(n4899), .A2(n4935), .ZN(n9555) );
  NAND2_X1 U6368 ( .A1(n4941), .A2(n9555), .ZN(n4900) );
  INV_X1 U6369 ( .A(n8323), .ZN(n9937) );
  NAND2_X1 U6370 ( .A1(n5548), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4909) );
  INV_X1 U6371 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n4905) );
  OR2_X1 U6372 ( .A1(n7624), .A2(n4905), .ZN(n4908) );
  OR2_X1 U6373 ( .A1(n5419), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n4907) );
  INV_X1 U6374 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6514) );
  OR2_X1 U6375 ( .A1(n6392), .A2(n6514), .ZN(n4906) );
  OR2_X1 U6376 ( .A1(n8333), .A2(n5489), .ZN(n4915) );
  NAND2_X1 U6377 ( .A1(n4912), .A2(SI_2_), .ZN(n4913) );
  INV_X1 U6378 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6364) );
  INV_X1 U6379 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6353) );
  MUX2_X1 U6380 ( .A(n6364), .B(n6353), .S(n4895), .Z(n4930) );
  XNOR2_X1 U6381 ( .A(n4930), .B(SI_3_), .ZN(n4928) );
  XNOR2_X1 U6382 ( .A(n4929), .B(n4928), .ZN(n6363) );
  OR2_X1 U6383 ( .A1(n4935), .A2(n4854), .ZN(n4914) );
  XNOR2_X1 U6384 ( .A(n4914), .B(P2_IR_REG_3__SCAN_IN), .ZN(n7978) );
  XNOR2_X1 U6385 ( .A(n5415), .B(n9873), .ZN(n4916) );
  XNOR2_X1 U6386 ( .A(n4915), .B(n4916), .ZN(n6765) );
  INV_X1 U6387 ( .A(n4915), .ZN(n4917) );
  NAND2_X1 U6388 ( .A1(n4917), .A2(n4916), .ZN(n4918) );
  NAND2_X1 U6389 ( .A1(n4919), .A2(n4918), .ZN(n6752) );
  INV_X1 U6390 ( .A(n6752), .ZN(n4947) );
  NAND2_X1 U6391 ( .A1(n5548), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4927) );
  INV_X1 U6392 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6517) );
  OR2_X1 U6393 ( .A1(n6392), .A2(n6517), .ZN(n4926) );
  INV_X1 U6394 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n4920) );
  OR2_X1 U6395 ( .A1(n7624), .A2(n4920), .ZN(n4925) );
  INV_X1 U6396 ( .A(n4960), .ZN(n4961) );
  INV_X1 U6397 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n4922) );
  INV_X1 U6398 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n4921) );
  NAND2_X1 U6399 ( .A1(n4922), .A2(n4921), .ZN(n4923) );
  NAND2_X1 U6400 ( .A1(n4961), .A2(n4923), .ZN(n6757) );
  OR2_X1 U6401 ( .A1(n9862), .A2(n5489), .ZN(n4945) );
  INV_X1 U6402 ( .A(n4930), .ZN(n4931) );
  NAND2_X1 U6403 ( .A1(n4931), .A2(SI_3_), .ZN(n4932) );
  NAND2_X1 U6404 ( .A1(n4933), .A2(n4932), .ZN(n4952) );
  INV_X1 U6405 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6369) );
  INV_X1 U6406 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6357) );
  XNOR2_X1 U6407 ( .A(n4952), .B(n4951), .ZN(n6368) );
  NAND2_X1 U6408 ( .A1(n7616), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n4943) );
  INV_X1 U6409 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4934) );
  AND2_X1 U6410 ( .A1(n4935), .A2(n4934), .ZN(n4938) );
  NOR2_X1 U6411 ( .A1(n4938), .A2(n4854), .ZN(n4936) );
  MUX2_X1 U6412 ( .A(n4854), .B(n4936), .S(P2_IR_REG_4__SCAN_IN), .Z(n4940) );
  INV_X1 U6413 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4937) );
  NAND2_X1 U6414 ( .A1(n4938), .A2(n4937), .ZN(n4949) );
  INV_X1 U6415 ( .A(n4949), .ZN(n4939) );
  NOR2_X1 U6416 ( .A1(n4940), .A2(n4939), .ZN(n7993) );
  NAND2_X1 U6417 ( .A1(n4941), .A2(n7993), .ZN(n4942) );
  OAI211_X1 U6418 ( .C1(n4957), .C2(n6368), .A(n4943), .B(n4942), .ZN(n9945)
         );
  XNOR2_X1 U6419 ( .A(n6759), .B(n5415), .ZN(n4944) );
  NAND2_X1 U6420 ( .A1(n4945), .A2(n4944), .ZN(n4948) );
  OAI21_X1 U6421 ( .B1(n4945), .B2(n4944), .A(n4948), .ZN(n6756) );
  NAND2_X1 U6422 ( .A1(n4949), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4950) );
  XNOR2_X1 U6423 ( .A(n4950), .B(P2_IR_REG_5__SCAN_IN), .ZN(n8006) );
  INV_X1 U6424 ( .A(n8006), .ZN(n6365) );
  NAND2_X1 U6425 ( .A1(n4952), .A2(n4951), .ZN(n4956) );
  INV_X1 U6426 ( .A(n4953), .ZN(n4954) );
  NAND2_X1 U6427 ( .A1(n4954), .A2(SI_4_), .ZN(n4955) );
  MUX2_X1 U6428 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7613), .Z(n4973) );
  XNOR2_X1 U6429 ( .A(n4973), .B(SI_5_), .ZN(n4970) );
  XNOR2_X1 U6430 ( .A(n4972), .B(n4970), .ZN(n6360) );
  NAND2_X1 U6431 ( .A1(n7616), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n4959) );
  XNOR2_X1 U6432 ( .A(n5415), .B(n9953), .ZN(n4968) );
  NAND2_X1 U6433 ( .A1(n5548), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4967) );
  INV_X1 U6434 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6733) );
  OR2_X1 U6435 ( .A1(n6392), .A2(n6733), .ZN(n4966) );
  INV_X1 U6436 ( .A(n4980), .ZN(n4982) );
  INV_X1 U6437 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8004) );
  NAND2_X1 U6438 ( .A1(n4961), .A2(n8004), .ZN(n4962) );
  NAND2_X1 U6439 ( .A1(n4982), .A2(n4962), .ZN(n6725) );
  OR2_X1 U6440 ( .A1(n5419), .A2(n6725), .ZN(n4965) );
  INV_X1 U6441 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n4963) );
  OR2_X1 U6442 ( .A1(n7624), .A2(n4963), .ZN(n4964) );
  NAND4_X1 U6443 ( .A1(n4967), .A2(n4966), .A3(n4965), .A4(n4964), .ZN(n7958)
         );
  AND2_X1 U6444 ( .A1(n7958), .A2(n4250), .ZN(n4969) );
  XNOR2_X1 U6445 ( .A(n4968), .B(n4969), .ZN(n6637) );
  INV_X1 U6446 ( .A(n4970), .ZN(n4971) );
  NAND2_X1 U6447 ( .A1(n4972), .A2(n4971), .ZN(n4975) );
  NAND2_X1 U6448 ( .A1(n4973), .A2(SI_5_), .ZN(n4974) );
  MUX2_X1 U6449 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7613), .Z(n4996) );
  XNOR2_X1 U6450 ( .A(n4995), .B(n4993), .ZN(n6370) );
  NAND2_X1 U6451 ( .A1(n6370), .A2(n7742), .ZN(n4979) );
  NAND2_X1 U6452 ( .A1(n4976), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4977) );
  XNOR2_X1 U6453 ( .A(n4977), .B(P2_IR_REG_6__SCAN_IN), .ZN(n8019) );
  AOI22_X1 U6454 ( .A1(n7616), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6405), .B2(
        n8019), .ZN(n4978) );
  NAND2_X1 U6455 ( .A1(n4979), .A2(n4978), .ZN(n6944) );
  INV_X2 U6456 ( .A(n5415), .ZN(n5490) );
  XNOR2_X1 U6457 ( .A(n6944), .B(n5490), .ZN(n4990) );
  NAND2_X1 U6458 ( .A1(n5548), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4988) );
  INV_X1 U6459 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6520) );
  OR2_X1 U6460 ( .A1(n6392), .A2(n6520), .ZN(n4987) );
  INV_X1 U6461 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n4981) );
  NAND2_X1 U6462 ( .A1(n4982), .A2(n4981), .ZN(n4983) );
  NAND2_X1 U6463 ( .A1(n5004), .A2(n4983), .ZN(n6904) );
  OR2_X1 U6464 ( .A1(n5419), .A2(n6904), .ZN(n4986) );
  INV_X1 U6465 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n4984) );
  OR2_X1 U6466 ( .A1(n7624), .A2(n4984), .ZN(n4985) );
  OR2_X1 U6467 ( .A1(n6949), .A2(n5489), .ZN(n4989) );
  NAND2_X1 U6468 ( .A1(n4990), .A2(n4989), .ZN(n4992) );
  OAI21_X1 U6469 ( .B1(n4990), .B2(n4989), .A(n4992), .ZN(n6739) );
  NAND2_X1 U6470 ( .A1(n6736), .A2(n4992), .ZN(n6772) );
  INV_X1 U6471 ( .A(n4993), .ZN(n4994) );
  NAND2_X1 U6472 ( .A1(n4996), .A2(SI_6_), .ZN(n4997) );
  MUX2_X1 U6473 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7613), .Z(n5017) );
  XNOR2_X1 U6474 ( .A(n5016), .B(n5014), .ZN(n6375) );
  NAND2_X1 U6475 ( .A1(n6375), .A2(n7742), .ZN(n5001) );
  NAND2_X1 U6476 ( .A1(n4998), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4999) );
  XNOR2_X1 U6477 ( .A(n4999), .B(P2_IR_REG_7__SCAN_IN), .ZN(n8031) );
  AOI22_X1 U6478 ( .A1(n7616), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6405), .B2(
        n8031), .ZN(n5000) );
  NAND2_X1 U6479 ( .A1(n5001), .A2(n5000), .ZN(n7056) );
  XNOR2_X1 U6480 ( .A(n7056), .B(n5415), .ZN(n5010) );
  NAND2_X1 U6481 ( .A1(n5548), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5009) );
  INV_X1 U6482 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6951) );
  OR2_X1 U6483 ( .A1(n6392), .A2(n6951), .ZN(n5008) );
  INV_X1 U6484 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5002) );
  OR2_X1 U6485 ( .A1(n7624), .A2(n5002), .ZN(n5007) );
  INV_X1 U6486 ( .A(n5004), .ZN(n5003) );
  INV_X1 U6487 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9410) );
  NAND2_X1 U6488 ( .A1(n5004), .A2(n9410), .ZN(n5005) );
  NAND2_X1 U6489 ( .A1(n5049), .A2(n5005), .ZN(n6955) );
  OR2_X1 U6490 ( .A1(n5419), .A2(n6955), .ZN(n5006) );
  NOR2_X1 U6491 ( .A1(n6970), .A2(n5489), .ZN(n5011) );
  XNOR2_X1 U6492 ( .A(n5010), .B(n5011), .ZN(n6771) );
  INV_X1 U6493 ( .A(n5010), .ZN(n5013) );
  INV_X1 U6494 ( .A(n5011), .ZN(n5012) );
  INV_X1 U6495 ( .A(n5014), .ZN(n5015) );
  MUX2_X1 U6496 ( .A(n6380), .B(n9360), .S(n7613), .Z(n5018) );
  NAND2_X1 U6497 ( .A1(n5018), .A2(n9346), .ZN(n5035) );
  INV_X1 U6498 ( .A(n5018), .ZN(n5019) );
  NAND2_X1 U6499 ( .A1(n5019), .A2(SI_8_), .ZN(n5020) );
  NAND2_X1 U6500 ( .A1(n5035), .A2(n5020), .ZN(n5036) );
  XNOR2_X1 U6501 ( .A(n5037), .B(n5036), .ZN(n6379) );
  NAND2_X1 U6502 ( .A1(n6379), .A2(n7742), .ZN(n5026) );
  NOR2_X1 U6503 ( .A1(n5021), .A2(n4854), .ZN(n5022) );
  MUX2_X1 U6504 ( .A(n4854), .B(n5022), .S(P2_IR_REG_8__SCAN_IN), .Z(n5024) );
  INV_X1 U6505 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5023) );
  AND2_X1 U6506 ( .A1(n5021), .A2(n5023), .ZN(n5068) );
  NOR2_X1 U6507 ( .A1(n5024), .A2(n5068), .ZN(n8044) );
  AOI22_X1 U6508 ( .A1(n7616), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6405), .B2(
        n8044), .ZN(n5025) );
  NAND2_X1 U6509 ( .A1(n5026), .A2(n5025), .ZN(n9969) );
  XNOR2_X1 U6510 ( .A(n9969), .B(n5490), .ZN(n5031) );
  NAND2_X1 U6511 ( .A1(n5548), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5030) );
  INV_X1 U6512 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6975) );
  OR2_X1 U6513 ( .A1(n6392), .A2(n6975), .ZN(n5029) );
  INV_X1 U6514 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5047) );
  XNOR2_X1 U6515 ( .A(n5049), .B(n5047), .ZN(n6974) );
  OR2_X1 U6516 ( .A1(n5419), .A2(n6974), .ZN(n5028) );
  INV_X1 U6517 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9451) );
  OR2_X1 U6518 ( .A1(n7624), .A2(n9451), .ZN(n5027) );
  NOR2_X1 U6519 ( .A1(n7157), .A2(n5489), .ZN(n5032) );
  XNOR2_X1 U6520 ( .A(n5031), .B(n5032), .ZN(n6833) );
  INV_X1 U6521 ( .A(n5031), .ZN(n5033) );
  NAND2_X1 U6522 ( .A1(n5033), .A2(n5032), .ZN(n5034) );
  MUX2_X1 U6523 ( .A(n5038), .B(n6387), .S(n7613), .Z(n5040) );
  INV_X1 U6524 ( .A(SI_9_), .ZN(n5039) );
  NAND2_X1 U6525 ( .A1(n5040), .A2(n5039), .ZN(n5062) );
  INV_X1 U6526 ( .A(n5040), .ZN(n5041) );
  NAND2_X1 U6527 ( .A1(n5041), .A2(SI_9_), .ZN(n5042) );
  XNOR2_X1 U6528 ( .A(n5061), .B(n4806), .ZN(n6383) );
  NAND2_X1 U6529 ( .A1(n6383), .A2(n7742), .ZN(n5045) );
  OR2_X1 U6530 ( .A1(n5068), .A2(n4854), .ZN(n5043) );
  XNOR2_X1 U6531 ( .A(n5043), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8057) );
  AOI22_X1 U6532 ( .A1(n7616), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6405), .B2(
        n8057), .ZN(n5044) );
  NAND2_X1 U6533 ( .A1(n5045), .A2(n5044), .ZN(n8434) );
  XNOR2_X1 U6534 ( .A(n8434), .B(n5490), .ZN(n5056) );
  NAND2_X1 U6535 ( .A1(n5548), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5055) );
  INV_X1 U6536 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7210) );
  OR2_X1 U6537 ( .A1(n6392), .A2(n7210), .ZN(n5054) );
  INV_X1 U6538 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5046) );
  OAI21_X1 U6539 ( .B1(n5049), .B2(n5047), .A(n5046), .ZN(n5050) );
  NAND2_X1 U6540 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5048) );
  NAND2_X1 U6541 ( .A1(n5050), .A2(n5073), .ZN(n7209) );
  OR2_X1 U6542 ( .A1(n5419), .A2(n7209), .ZN(n5053) );
  INV_X1 U6543 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5051) );
  OR2_X1 U6544 ( .A1(n7624), .A2(n5051), .ZN(n5052) );
  OR2_X1 U6545 ( .A1(n7162), .A2(n5489), .ZN(n5057) );
  NAND2_X1 U6546 ( .A1(n5056), .A2(n5057), .ZN(n7108) );
  INV_X1 U6547 ( .A(n5056), .ZN(n5059) );
  INV_X1 U6548 ( .A(n5057), .ZN(n5058) );
  NAND2_X1 U6549 ( .A1(n5059), .A2(n5058), .ZN(n5060) );
  NAND2_X1 U6550 ( .A1(n7108), .A2(n5060), .ZN(n7041) );
  MUX2_X1 U6551 ( .A(n6399), .B(n6400), .S(n7613), .Z(n5064) );
  NAND2_X1 U6552 ( .A1(n5064), .A2(n5063), .ZN(n5087) );
  INV_X1 U6553 ( .A(n5064), .ZN(n5065) );
  NAND2_X1 U6554 ( .A1(n5065), .A2(SI_10_), .ZN(n5066) );
  NAND2_X1 U6555 ( .A1(n6398), .A2(n7742), .ZN(n5071) );
  INV_X1 U6556 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5067) );
  OR2_X1 U6557 ( .A1(n5091), .A2(n4854), .ZN(n5069) );
  XNOR2_X1 U6558 ( .A(n5069), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6551) );
  AOI22_X1 U6559 ( .A1(n7616), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6405), .B2(
        n6551), .ZN(n5070) );
  NAND2_X1 U6560 ( .A1(n5071), .A2(n5070), .ZN(n9976) );
  XNOR2_X1 U6561 ( .A(n9976), .B(n5415), .ZN(n5082) );
  NAND2_X1 U6562 ( .A1(n5420), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5079) );
  INV_X1 U6563 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7170) );
  OR2_X1 U6564 ( .A1(n6392), .A2(n7170), .ZN(n5078) );
  INV_X1 U6565 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6681) );
  NAND2_X1 U6566 ( .A1(n5073), .A2(n6681), .ZN(n5074) );
  NAND2_X1 U6567 ( .A1(n5095), .A2(n5074), .ZN(n7169) );
  OR2_X1 U6568 ( .A1(n5419), .A2(n7169), .ZN(n5077) );
  INV_X1 U6569 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5075) );
  OR2_X1 U6570 ( .A1(n4903), .A2(n5075), .ZN(n5076) );
  NOR2_X1 U6571 ( .A1(n7203), .A2(n5489), .ZN(n5081) );
  AND2_X1 U6572 ( .A1(n5082), .A2(n5081), .ZN(n5085) );
  OR2_X1 U6573 ( .A1(n7041), .A2(n5085), .ZN(n5080) );
  XNOR2_X1 U6574 ( .A(n5082), .B(n5081), .ZN(n7111) );
  INV_X1 U6575 ( .A(n7111), .ZN(n5083) );
  AND2_X1 U6576 ( .A1(n5083), .A2(n7108), .ZN(n5084) );
  NAND2_X1 U6577 ( .A1(n5086), .A2(n4271), .ZN(n5088) );
  MUX2_X1 U6578 ( .A(n5089), .B(n6403), .S(n7613), .Z(n5106) );
  XNOR2_X1 U6579 ( .A(n5106), .B(SI_11_), .ZN(n5105) );
  INV_X1 U6580 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5090) );
  NAND2_X1 U6581 ( .A1(n5091), .A2(n5090), .ZN(n5117) );
  NAND2_X1 U6582 ( .A1(n5117), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5092) );
  XNOR2_X1 U6583 ( .A(n5092), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6609) );
  AOI22_X1 U6584 ( .A1(n7616), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6405), .B2(
        n6609), .ZN(n5093) );
  XNOR2_X1 U6585 ( .A(n8429), .B(n5490), .ZN(n5101) );
  NAND2_X1 U6586 ( .A1(n5420), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5100) );
  INV_X1 U6587 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7352) );
  OR2_X1 U6588 ( .A1(n6392), .A2(n7352), .ZN(n5099) );
  NAND2_X1 U6589 ( .A1(n5095), .A2(n5094), .ZN(n5096) );
  NAND2_X1 U6590 ( .A1(n5123), .A2(n5096), .ZN(n7351) );
  OR2_X1 U6591 ( .A1(n5419), .A2(n7351), .ZN(n5098) );
  INV_X1 U6592 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6552) );
  OR2_X1 U6593 ( .A1(n4903), .A2(n6552), .ZN(n5097) );
  NOR2_X1 U6594 ( .A1(n7368), .A2(n5489), .ZN(n5102) );
  XNOR2_X1 U6595 ( .A(n5101), .B(n5102), .ZN(n7077) );
  INV_X1 U6596 ( .A(n5101), .ZN(n5103) );
  AND2_X1 U6597 ( .A1(n5103), .A2(n5102), .ZN(n5104) );
  INV_X1 U6598 ( .A(n5105), .ZN(n5109) );
  INV_X1 U6599 ( .A(n5106), .ZN(n5107) );
  NAND2_X1 U6600 ( .A1(n5107), .A2(SI_11_), .ZN(n5108) );
  INV_X8 U6601 ( .A(n5111), .ZN(n7613) );
  MUX2_X1 U6602 ( .A(n6426), .B(n5112), .S(n7613), .Z(n5114) );
  INV_X1 U6603 ( .A(SI_12_), .ZN(n5113) );
  INV_X1 U6604 ( .A(n5114), .ZN(n5115) );
  NAND2_X1 U6605 ( .A1(n5115), .A2(SI_12_), .ZN(n5116) );
  NAND2_X1 U6606 ( .A1(n5135), .A2(n5116), .ZN(n5136) );
  XNOR2_X1 U6607 ( .A(n5137), .B(n5136), .ZN(n6409) );
  NAND2_X1 U6608 ( .A1(n6409), .A2(n7742), .ZN(n5120) );
  NAND2_X1 U6609 ( .A1(n5142), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5118) );
  XNOR2_X1 U6610 ( .A(n5118), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6554) );
  AOI22_X1 U6611 ( .A1(n7743), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6405), .B2(
        n6554), .ZN(n5119) );
  NAND2_X1 U6612 ( .A1(n5120), .A2(n5119), .ZN(n7449) );
  XNOR2_X1 U6613 ( .A(n7449), .B(n5490), .ZN(n5129) );
  NAND2_X1 U6614 ( .A1(n5420), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5128) );
  INV_X1 U6615 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6526) );
  OR2_X1 U6616 ( .A1(n6392), .A2(n6526), .ZN(n5127) );
  INV_X1 U6617 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6553) );
  OR2_X1 U6618 ( .A1(n4903), .A2(n6553), .ZN(n5126) );
  INV_X1 U6619 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U6620 ( .A1(n5123), .A2(n5122), .ZN(n5124) );
  NAND2_X1 U6621 ( .A1(n5146), .A2(n5124), .ZN(n7219) );
  OR2_X1 U6622 ( .A1(n5419), .A2(n7219), .ZN(n5125) );
  OR2_X1 U6623 ( .A1(n7365), .A2(n5489), .ZN(n5130) );
  NAND2_X1 U6624 ( .A1(n5129), .A2(n5130), .ZN(n5134) );
  INV_X1 U6625 ( .A(n5129), .ZN(n5132) );
  INV_X1 U6626 ( .A(n5130), .ZN(n5131) );
  NAND2_X1 U6627 ( .A1(n5132), .A2(n5131), .ZN(n5133) );
  AND2_X1 U6628 ( .A1(n5134), .A2(n5133), .ZN(n7216) );
  MUX2_X1 U6629 ( .A(n6435), .B(n9427), .S(n7613), .Z(n5139) );
  INV_X1 U6630 ( .A(n5139), .ZN(n5140) );
  NAND2_X1 U6631 ( .A1(n5140), .A2(SI_13_), .ZN(n5141) );
  XNOR2_X1 U6632 ( .A(n5159), .B(n4805), .ZN(n6432) );
  NAND2_X1 U6633 ( .A1(n6432), .A2(n7742), .ZN(n5144) );
  OAI21_X1 U6634 ( .B1(n5142), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5163) );
  XNOR2_X1 U6635 ( .A(n5163), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6658) );
  AOI22_X1 U6636 ( .A1(n7616), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6405), .B2(
        n6658), .ZN(n5143) );
  XNOR2_X1 U6637 ( .A(n8424), .B(n5490), .ZN(n5153) );
  NAND2_X1 U6638 ( .A1(n5420), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5151) );
  INV_X1 U6639 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6535) );
  OR2_X1 U6640 ( .A1(n4903), .A2(n6535), .ZN(n5150) );
  INV_X1 U6641 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6527) );
  OR2_X1 U6642 ( .A1(n6392), .A2(n6527), .ZN(n5149) );
  NAND2_X1 U6643 ( .A1(n5146), .A2(n5145), .ZN(n5147) );
  NAND2_X1 U6644 ( .A1(n5168), .A2(n5147), .ZN(n7247) );
  OR2_X1 U6645 ( .A1(n5419), .A2(n7247), .ZN(n5148) );
  NAND4_X1 U6646 ( .A1(n5151), .A2(n5150), .A3(n5149), .A4(n5148), .ZN(n7951)
         );
  NAND2_X1 U6647 ( .A1(n7951), .A2(n4250), .ZN(n5154) );
  XNOR2_X1 U6648 ( .A(n5153), .B(n5154), .ZN(n7245) );
  INV_X1 U6649 ( .A(n7245), .ZN(n5152) );
  INV_X1 U6650 ( .A(n5153), .ZN(n5156) );
  INV_X1 U6651 ( .A(n5154), .ZN(n5155) );
  NAND2_X1 U6652 ( .A1(n5156), .A2(n5155), .ZN(n5157) );
  NAND2_X1 U6653 ( .A1(n5158), .A2(n5157), .ZN(n7440) );
  INV_X1 U6654 ( .A(n7440), .ZN(n5181) );
  MUX2_X1 U6655 ( .A(n6439), .B(n6437), .S(n7613), .Z(n5184) );
  XNOR2_X1 U6656 ( .A(n5184), .B(SI_14_), .ZN(n5183) );
  XNOR2_X1 U6657 ( .A(n5188), .B(n5183), .ZN(n6436) );
  NAND2_X1 U6658 ( .A1(n6436), .A2(n7742), .ZN(n5166) );
  INV_X1 U6659 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5162) );
  NAND2_X1 U6660 ( .A1(n5163), .A2(n5162), .ZN(n5164) );
  NAND2_X1 U6661 ( .A1(n5164), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5194) );
  XNOR2_X1 U6662 ( .A(n5194), .B(P2_IR_REG_14__SCAN_IN), .ZN(n6659) );
  AOI22_X1 U6663 ( .A1(n7616), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6659), .B2(
        n6405), .ZN(n5165) );
  XNOR2_X1 U6664 ( .A(n7488), .B(n5490), .ZN(n5175) );
  NAND2_X1 U6665 ( .A1(n5548), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5174) );
  INV_X1 U6666 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7471) );
  OR2_X1 U6667 ( .A1(n6392), .A2(n7471), .ZN(n5173) );
  INV_X1 U6668 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6669 ( .A1(n5168), .A2(n5167), .ZN(n5169) );
  NAND2_X1 U6670 ( .A1(n5201), .A2(n5169), .ZN(n7470) );
  OR2_X1 U6671 ( .A1(n5419), .A2(n7470), .ZN(n5172) );
  INV_X1 U6672 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n5170) );
  OR2_X1 U6673 ( .A1(n7624), .A2(n5170), .ZN(n5171) );
  OR2_X1 U6674 ( .A1(n7517), .A2(n5489), .ZN(n5176) );
  NAND2_X1 U6675 ( .A1(n5175), .A2(n5176), .ZN(n5182) );
  INV_X1 U6676 ( .A(n5175), .ZN(n5178) );
  INV_X1 U6677 ( .A(n5176), .ZN(n5177) );
  NAND2_X1 U6678 ( .A1(n5178), .A2(n5177), .ZN(n5179) );
  NAND2_X1 U6679 ( .A1(n5182), .A2(n5179), .ZN(n7441) );
  INV_X1 U6680 ( .A(n7441), .ZN(n5180) );
  NAND2_X1 U6681 ( .A1(n5181), .A2(n5180), .ZN(n7438) );
  NAND2_X1 U6682 ( .A1(n7438), .A2(n5182), .ZN(n5208) );
  INV_X1 U6683 ( .A(n5183), .ZN(n5187) );
  INV_X1 U6684 ( .A(n5184), .ZN(n5185) );
  NAND2_X1 U6685 ( .A1(n5185), .A2(SI_14_), .ZN(n5186) );
  MUX2_X1 U6686 ( .A(n9428), .B(n6508), .S(n7613), .Z(n5190) );
  INV_X1 U6687 ( .A(SI_15_), .ZN(n5189) );
  NAND2_X1 U6688 ( .A1(n5190), .A2(n5189), .ZN(n5213) );
  INV_X1 U6689 ( .A(n5190), .ZN(n5191) );
  NAND2_X1 U6690 ( .A1(n5191), .A2(SI_15_), .ZN(n5192) );
  NAND2_X1 U6691 ( .A1(n5213), .A2(n5192), .ZN(n5214) );
  XNOR2_X1 U6692 ( .A(n5215), .B(n5214), .ZN(n6507) );
  NAND2_X1 U6693 ( .A1(n6507), .A2(n7742), .ZN(n5198) );
  INV_X1 U6694 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U6695 ( .A1(n5194), .A2(n5193), .ZN(n5195) );
  NAND2_X1 U6696 ( .A1(n5195), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5196) );
  XNOR2_X1 U6697 ( .A(n5196), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6799) );
  AOI22_X1 U6698 ( .A1(n6799), .A2(n6405), .B1(n7743), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5197) );
  XNOR2_X1 U6699 ( .A(n8419), .B(n5415), .ZN(n5209) );
  XNOR2_X1 U6700 ( .A(n5208), .B(n5209), .ZN(n7514) );
  NAND2_X1 U6701 ( .A1(n7621), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5207) );
  INV_X1 U6702 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6661) );
  OR2_X1 U6703 ( .A1(n4903), .A2(n6661), .ZN(n5206) );
  INV_X1 U6704 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U6705 ( .A1(n5201), .A2(n5200), .ZN(n5202) );
  NAND2_X1 U6706 ( .A1(n5225), .A2(n5202), .ZN(n7516) );
  OR2_X1 U6707 ( .A1(n5419), .A2(n7516), .ZN(n5205) );
  INV_X1 U6708 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n5203) );
  OR2_X1 U6709 ( .A1(n7624), .A2(n5203), .ZN(n5204) );
  NOR2_X1 U6710 ( .A1(n7525), .A2(n5489), .ZN(n7515) );
  NAND2_X1 U6711 ( .A1(n7514), .A2(n7515), .ZN(n5212) );
  INV_X1 U6712 ( .A(n5208), .ZN(n5210) );
  NAND2_X1 U6713 ( .A1(n5210), .A2(n5209), .ZN(n5211) );
  NAND2_X1 U6714 ( .A1(n5212), .A2(n5211), .ZN(n7584) );
  INV_X1 U6715 ( .A(n7584), .ZN(n5237) );
  MUX2_X1 U6716 ( .A(n6592), .B(n6590), .S(n7613), .Z(n5217) );
  INV_X1 U6717 ( .A(SI_16_), .ZN(n5216) );
  NAND2_X1 U6718 ( .A1(n5217), .A2(n5216), .ZN(n5241) );
  INV_X1 U6719 ( .A(n5217), .ZN(n5218) );
  NAND2_X1 U6720 ( .A1(n5218), .A2(SI_16_), .ZN(n5219) );
  XNOR2_X1 U6721 ( .A(n5240), .B(n5239), .ZN(n6589) );
  NAND2_X1 U6722 ( .A1(n6589), .A2(n7742), .ZN(n5223) );
  NAND2_X1 U6723 ( .A1(n5220), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5221) );
  XNOR2_X1 U6724 ( .A(n5221), .B(P2_IR_REG_16__SCAN_IN), .ZN(n7089) );
  AOI22_X1 U6725 ( .A1(n7743), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6405), .B2(
        n7089), .ZN(n5222) );
  XNOR2_X1 U6726 ( .A(n7591), .B(n5490), .ZN(n5231) );
  NAND2_X1 U6727 ( .A1(n5420), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5230) );
  INV_X1 U6728 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n6792) );
  OR2_X1 U6729 ( .A1(n4903), .A2(n6792), .ZN(n5229) );
  INV_X1 U6730 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7531) );
  OR2_X1 U6731 ( .A1(n6392), .A2(n7531), .ZN(n5228) );
  INV_X1 U6732 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9392) );
  NAND2_X1 U6733 ( .A1(n5225), .A2(n9392), .ZN(n5226) );
  NAND2_X1 U6734 ( .A1(n5248), .A2(n5226), .ZN(n7589) );
  OR2_X1 U6735 ( .A1(n5419), .A2(n7589), .ZN(n5227) );
  OR2_X1 U6736 ( .A1(n7573), .A2(n5489), .ZN(n5232) );
  NAND2_X1 U6737 ( .A1(n5231), .A2(n5232), .ZN(n5238) );
  INV_X1 U6738 ( .A(n5231), .ZN(n5234) );
  INV_X1 U6739 ( .A(n5232), .ZN(n5233) );
  NAND2_X1 U6740 ( .A1(n5234), .A2(n5233), .ZN(n5235) );
  NAND2_X1 U6741 ( .A1(n5238), .A2(n5235), .ZN(n7585) );
  INV_X1 U6742 ( .A(n7585), .ZN(n5236) );
  NAND2_X2 U6743 ( .A1(n5237), .A2(n5236), .ZN(n7582) );
  MUX2_X1 U6744 ( .A(n6636), .B(n9429), .S(n7613), .Z(n5258) );
  XNOR2_X1 U6745 ( .A(n5258), .B(SI_17_), .ZN(n5257) );
  XNOR2_X1 U6746 ( .A(n5262), .B(n5257), .ZN(n6634) );
  NAND2_X1 U6747 ( .A1(n6634), .A2(n7742), .ZN(n5245) );
  NAND2_X1 U6748 ( .A1(n5242), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5243) );
  XNOR2_X1 U6749 ( .A(n5243), .B(P2_IR_REG_17__SCAN_IN), .ZN(n7280) );
  AOI22_X1 U6750 ( .A1(n7616), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6405), .B2(
        n7280), .ZN(n5244) );
  XNOR2_X1 U6751 ( .A(n8093), .B(n5490), .ZN(n5255) );
  NAND2_X1 U6752 ( .A1(n5420), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5253) );
  INV_X1 U6753 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7577) );
  OR2_X1 U6754 ( .A1(n6392), .A2(n7577), .ZN(n5252) );
  INV_X1 U6755 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n5246) );
  OR2_X1 U6756 ( .A1(n4903), .A2(n5246), .ZN(n5251) );
  INV_X1 U6757 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U6758 ( .A1(n5248), .A2(n5247), .ZN(n5249) );
  NAND2_X1 U6759 ( .A1(n5268), .A2(n5249), .ZN(n7892) );
  OR2_X1 U6760 ( .A1(n5419), .A2(n7892), .ZN(n5250) );
  INV_X1 U6761 ( .A(n7926), .ZN(n8311) );
  NAND2_X1 U6762 ( .A1(n8311), .A2(n4250), .ZN(n5254) );
  XNOR2_X1 U6763 ( .A(n5255), .B(n5254), .ZN(n7887) );
  INV_X1 U6764 ( .A(n5257), .ZN(n5261) );
  INV_X1 U6765 ( .A(n5258), .ZN(n5259) );
  NAND2_X1 U6766 ( .A1(n5259), .A2(SI_17_), .ZN(n5260) );
  MUX2_X1 U6767 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7613), .Z(n5280) );
  XNOR2_X1 U6768 ( .A(n5280), .B(SI_18_), .ZN(n5277) );
  XNOR2_X1 U6769 ( .A(n5279), .B(n5277), .ZN(n6784) );
  NAND2_X1 U6770 ( .A1(n6784), .A2(n7742), .ZN(n5265) );
  NAND2_X1 U6771 ( .A1(n4836), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5263) );
  XNOR2_X1 U6772 ( .A(n5263), .B(P2_IR_REG_18__SCAN_IN), .ZN(n7285) );
  AOI22_X1 U6773 ( .A1(n7743), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6405), .B2(
        n7285), .ZN(n5264) );
  XNOR2_X1 U6774 ( .A(n8308), .B(n5415), .ZN(n5274) );
  INV_X1 U6775 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U6776 ( .A1(n5268), .A2(n5267), .ZN(n5269) );
  NAND2_X1 U6777 ( .A1(n5290), .A2(n5269), .ZN(n8304) );
  OR2_X1 U6778 ( .A1(n8304), .A2(n5419), .ZN(n5273) );
  NAND2_X1 U6779 ( .A1(n7621), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U6780 ( .A1(n5548), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6781 ( .A1(n5420), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5270) );
  NOR2_X1 U6782 ( .A1(n8097), .A2(n5489), .ZN(n5275) );
  XNOR2_X1 U6783 ( .A(n5274), .B(n5275), .ZN(n7923) );
  INV_X1 U6784 ( .A(n5274), .ZN(n5276) );
  INV_X1 U6785 ( .A(n7862), .ZN(n5301) );
  NAND2_X1 U6786 ( .A1(n5279), .A2(n5278), .ZN(n5282) );
  NAND2_X1 U6787 ( .A1(n5280), .A2(SI_18_), .ZN(n5281) );
  MUX2_X1 U6788 ( .A(n6863), .B(n6861), .S(n7613), .Z(n5284) );
  INV_X1 U6789 ( .A(SI_19_), .ZN(n5283) );
  NAND2_X1 U6790 ( .A1(n5284), .A2(n5283), .ZN(n5305) );
  INV_X1 U6791 ( .A(n5284), .ZN(n5285) );
  NAND2_X1 U6792 ( .A1(n5285), .A2(SI_19_), .ZN(n5286) );
  NAND2_X1 U6793 ( .A1(n5305), .A2(n5286), .ZN(n5303) );
  XNOR2_X1 U6794 ( .A(n5304), .B(n5303), .ZN(n6860) );
  NAND2_X1 U6795 ( .A1(n6860), .A2(n7742), .ZN(n5288) );
  AOI22_X1 U6796 ( .A1(n7743), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6405), .B2(
        n8077), .ZN(n5287) );
  XNOR2_X1 U6797 ( .A(n8298), .B(n5415), .ZN(n5295) );
  INV_X1 U6798 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6799 ( .A1(n5290), .A2(n5289), .ZN(n5291) );
  AND2_X1 U6800 ( .A1(n5313), .A2(n5291), .ZN(n8295) );
  NAND2_X1 U6801 ( .A1(n8295), .A2(n5438), .ZN(n5294) );
  AOI22_X1 U6802 ( .A1(n5548), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n7621), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6803 ( .A1(n5420), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5292) );
  OR2_X1 U6804 ( .A1(n8268), .A2(n5489), .ZN(n5296) );
  NAND2_X1 U6805 ( .A1(n5295), .A2(n5296), .ZN(n5302) );
  INV_X1 U6806 ( .A(n5295), .ZN(n5298) );
  INV_X1 U6807 ( .A(n5296), .ZN(n5297) );
  NAND2_X1 U6808 ( .A1(n5298), .A2(n5297), .ZN(n5299) );
  NAND2_X1 U6809 ( .A1(n5302), .A2(n5299), .ZN(n7861) );
  MUX2_X1 U6810 ( .A(n7025), .B(n9348), .S(n7613), .Z(n5307) );
  INV_X1 U6811 ( .A(SI_20_), .ZN(n5306) );
  NAND2_X1 U6812 ( .A1(n5307), .A2(n5306), .ZN(n5322) );
  INV_X1 U6813 ( .A(n5307), .ZN(n5308) );
  NAND2_X1 U6814 ( .A1(n5308), .A2(SI_20_), .ZN(n5309) );
  XNOR2_X1 U6815 ( .A(n5321), .B(n5320), .ZN(n7023) );
  NAND2_X1 U6816 ( .A1(n7023), .A2(n7742), .ZN(n5311) );
  NAND2_X1 U6817 ( .A1(n7743), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5310) );
  XNOR2_X1 U6818 ( .A(n8392), .B(n5415), .ZN(n5319) );
  INV_X1 U6819 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n5317) );
  INV_X1 U6820 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7909) );
  NAND2_X1 U6821 ( .A1(n5313), .A2(n7909), .ZN(n5314) );
  NAND2_X1 U6822 ( .A1(n5348), .A2(n5314), .ZN(n8273) );
  OR2_X1 U6823 ( .A1(n8273), .A2(n5419), .ZN(n5316) );
  AOI22_X1 U6824 ( .A1(n5420), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n7621), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n5315) );
  OAI211_X1 U6825 ( .C1(n4903), .C2(n5317), .A(n5316), .B(n5315), .ZN(n8260)
         );
  NAND2_X1 U6826 ( .A1(n8260), .A2(n4250), .ZN(n5318) );
  XNOR2_X1 U6827 ( .A(n5319), .B(n5318), .ZN(n7907) );
  MUX2_X1 U6828 ( .A(n7049), .B(n7047), .S(n7613), .Z(n5335) );
  XNOR2_X1 U6829 ( .A(n5335), .B(SI_21_), .ZN(n5334) );
  XNOR2_X1 U6830 ( .A(n5339), .B(n5334), .ZN(n7046) );
  NAND2_X1 U6831 ( .A1(n7046), .A2(n7742), .ZN(n5324) );
  NAND2_X1 U6832 ( .A1(n7743), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5323) );
  XNOR2_X1 U6833 ( .A(n8385), .B(n5415), .ZN(n5333) );
  XNOR2_X1 U6834 ( .A(n5348), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n8254) );
  NAND2_X1 U6835 ( .A1(n8254), .A2(n5438), .ZN(n5330) );
  INV_X1 U6836 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6837 ( .A1(n5548), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6838 ( .A1(n7621), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5325) );
  OAI211_X1 U6839 ( .C1(n5327), .C2(n7624), .A(n5326), .B(n5325), .ZN(n5328)
         );
  INV_X1 U6840 ( .A(n5328), .ZN(n5329) );
  NAND2_X1 U6841 ( .A1(n5330), .A2(n5329), .ZN(n8102) );
  NAND2_X1 U6842 ( .A1(n8102), .A2(n4250), .ZN(n5331) );
  XNOR2_X1 U6843 ( .A(n5333), .B(n5331), .ZN(n7869) );
  INV_X1 U6844 ( .A(n5331), .ZN(n5332) );
  INV_X1 U6845 ( .A(n5334), .ZN(n5338) );
  INV_X1 U6846 ( .A(n5335), .ZN(n5336) );
  NAND2_X1 U6847 ( .A1(n5336), .A2(SI_21_), .ZN(n5337) );
  MUX2_X1 U6848 ( .A(n7595), .B(n7240), .S(n7613), .Z(n5341) );
  INV_X1 U6849 ( .A(SI_22_), .ZN(n5340) );
  NAND2_X1 U6850 ( .A1(n5341), .A2(n5340), .ZN(n5360) );
  INV_X1 U6851 ( .A(n5341), .ZN(n5342) );
  NAND2_X1 U6852 ( .A1(n5342), .A2(SI_22_), .ZN(n5343) );
  NAND2_X1 U6853 ( .A1(n5360), .A2(n5343), .ZN(n5361) );
  XNOR2_X1 U6854 ( .A(n5362), .B(n5361), .ZN(n7239) );
  NAND2_X1 U6855 ( .A1(n7239), .A2(n7742), .ZN(n5345) );
  NAND2_X1 U6856 ( .A1(n7616), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5344) );
  XNOR2_X1 U6857 ( .A(n8380), .B(n5490), .ZN(n5356) );
  INV_X1 U6858 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9424) );
  INV_X1 U6859 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5346) );
  OAI21_X1 U6860 ( .B1(n5348), .B2(n9424), .A(n5346), .ZN(n5349) );
  NAND2_X1 U6861 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n5347) );
  NAND2_X1 U6862 ( .A1(n5349), .A2(n5385), .ZN(n8235) );
  OR2_X1 U6863 ( .A1(n8235), .A2(n5419), .ZN(n5355) );
  INV_X1 U6864 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U6865 ( .A1(n7621), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5351) );
  NAND2_X1 U6866 ( .A1(n5548), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5350) );
  OAI211_X1 U6867 ( .C1(n7624), .C2(n5352), .A(n5351), .B(n5350), .ZN(n5353)
         );
  INV_X1 U6868 ( .A(n5353), .ZN(n5354) );
  NAND2_X1 U6869 ( .A1(n8261), .A2(n4250), .ZN(n7915) );
  INV_X1 U6870 ( .A(n5356), .ZN(n5357) );
  OR2_X1 U6871 ( .A1(n5358), .A2(n5357), .ZN(n5359) );
  INV_X1 U6872 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5363) );
  MUX2_X1 U6873 ( .A(n5363), .B(n7244), .S(n7613), .Z(n5365) );
  INV_X1 U6874 ( .A(SI_23_), .ZN(n5364) );
  NAND2_X1 U6875 ( .A1(n5365), .A2(n5364), .ZN(n5372) );
  INV_X1 U6876 ( .A(n5365), .ZN(n5366) );
  NAND2_X1 U6877 ( .A1(n5366), .A2(SI_23_), .ZN(n5367) );
  XNOR2_X1 U6878 ( .A(n5371), .B(n5370), .ZN(n7241) );
  NAND2_X1 U6879 ( .A1(n7241), .A2(n7742), .ZN(n5369) );
  NAND2_X1 U6880 ( .A1(n7743), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5368) );
  XNOR2_X1 U6881 ( .A(n7627), .B(n5415), .ZN(n5398) );
  MUX2_X1 U6882 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n7613), .Z(n5405) );
  INV_X1 U6883 ( .A(SI_24_), .ZN(n5374) );
  XNOR2_X1 U6884 ( .A(n5405), .B(n5374), .ZN(n5404) );
  XNOR2_X1 U6885 ( .A(n5408), .B(n5404), .ZN(n7387) );
  NAND2_X1 U6886 ( .A1(n7387), .A2(n7742), .ZN(n5376) );
  NAND2_X1 U6887 ( .A1(n7743), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5375) );
  XNOR2_X1 U6888 ( .A(n8205), .B(n5415), .ZN(n7899) );
  INV_X1 U6889 ( .A(n5387), .ZN(n5378) );
  INV_X1 U6890 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n7902) );
  NAND2_X1 U6891 ( .A1(n5387), .A2(n7902), .ZN(n5379) );
  NAND2_X1 U6892 ( .A1(n5417), .A2(n5379), .ZN(n8202) );
  OR2_X1 U6893 ( .A1(n8202), .A2(n5419), .ZN(n5384) );
  INV_X1 U6894 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9434) );
  NAND2_X1 U6895 ( .A1(n7621), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U6896 ( .A1(n5548), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5380) );
  OAI211_X1 U6897 ( .C1(n7624), .C2(n9434), .A(n5381), .B(n5380), .ZN(n5382)
         );
  INV_X1 U6898 ( .A(n5382), .ZN(n5383) );
  INV_X1 U6899 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7854) );
  NAND2_X1 U6900 ( .A1(n5385), .A2(n7854), .ZN(n5386) );
  NAND2_X1 U6901 ( .A1(n5387), .A2(n5386), .ZN(n8224) );
  OR2_X1 U6902 ( .A1(n8224), .A2(n5419), .ZN(n5393) );
  INV_X1 U6903 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6904 ( .A1(n5548), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U6905 ( .A1(n7621), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5388) );
  OAI211_X1 U6906 ( .C1(n5390), .C2(n7624), .A(n5389), .B(n5388), .ZN(n5391)
         );
  INV_X1 U6907 ( .A(n5391), .ZN(n5392) );
  NAND2_X1 U6908 ( .A1(n5393), .A2(n5392), .ZN(n7947) );
  NAND2_X1 U6909 ( .A1(n7947), .A2(n4250), .ZN(n7897) );
  INV_X1 U6910 ( .A(n7897), .ZN(n5394) );
  NOR2_X2 U6911 ( .A1(n7853), .A2(n5396), .ZN(n5403) );
  OR2_X1 U6912 ( .A1(n7946), .A2(n5489), .ZN(n5399) );
  INV_X1 U6913 ( .A(n7899), .ZN(n5400) );
  INV_X1 U6914 ( .A(n5399), .ZN(n7898) );
  INV_X1 U6915 ( .A(n5404), .ZN(n5407) );
  NAND2_X1 U6916 ( .A1(n5405), .A2(SI_24_), .ZN(n5406) );
  INV_X1 U6917 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7480) );
  MUX2_X1 U6918 ( .A(n7480), .B(n7483), .S(n7613), .Z(n5410) );
  INV_X1 U6919 ( .A(SI_25_), .ZN(n5409) );
  NAND2_X1 U6920 ( .A1(n5410), .A2(n5409), .ZN(n5430) );
  INV_X1 U6921 ( .A(n5410), .ZN(n5411) );
  NAND2_X1 U6922 ( .A1(n5411), .A2(SI_25_), .ZN(n5412) );
  NAND2_X1 U6923 ( .A1(n5430), .A2(n5412), .ZN(n5428) );
  NAND2_X1 U6924 ( .A1(n7477), .A2(n7742), .ZN(n5414) );
  NAND2_X1 U6925 ( .A1(n7743), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5413) );
  XNOR2_X1 U6926 ( .A(n8366), .B(n5415), .ZN(n5427) );
  INV_X1 U6927 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U6928 ( .A1(n5417), .A2(n5416), .ZN(n5418) );
  NAND2_X1 U6929 ( .A1(n5436), .A2(n5418), .ZN(n8192) );
  OR2_X1 U6930 ( .A1(n8192), .A2(n5419), .ZN(n5425) );
  INV_X1 U6931 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n9450) );
  NAND2_X1 U6932 ( .A1(n5548), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U6933 ( .A1(n5420), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5421) );
  OAI211_X1 U6934 ( .C1(n6392), .C2(n9450), .A(n5422), .B(n5421), .ZN(n5423)
         );
  INV_X1 U6935 ( .A(n5423), .ZN(n5424) );
  NOR2_X1 U6936 ( .A1(n8210), .A2(n5489), .ZN(n5426) );
  NOR2_X1 U6937 ( .A1(n5427), .A2(n5426), .ZN(n7878) );
  NAND2_X1 U6938 ( .A1(n5427), .A2(n5426), .ZN(n7879) );
  OAI21_X1 U6939 ( .B1(n7877), .B2(n7878), .A(n7879), .ZN(n7936) );
  INV_X1 U6940 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7537) );
  INV_X1 U6941 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7539) );
  MUX2_X1 U6942 ( .A(n7537), .B(n7539), .S(n7613), .Z(n5431) );
  INV_X1 U6943 ( .A(SI_26_), .ZN(n9449) );
  NAND2_X1 U6944 ( .A1(n5431), .A2(n9449), .ZN(n5451) );
  INV_X1 U6945 ( .A(n5431), .ZN(n5432) );
  NAND2_X1 U6946 ( .A1(n5432), .A2(SI_26_), .ZN(n5433) );
  NAND2_X1 U6947 ( .A1(n7536), .A2(n7742), .ZN(n5435) );
  NAND2_X1 U6948 ( .A1(n7743), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5434) );
  XNOR2_X1 U6949 ( .A(n8181), .B(n5415), .ZN(n5446) );
  INV_X1 U6950 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7937) );
  NAND2_X1 U6951 ( .A1(n5436), .A2(n7937), .ZN(n5437) );
  NAND2_X1 U6952 ( .A1(n8178), .A2(n5438), .ZN(n5444) );
  INV_X1 U6953 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U6954 ( .A1(n5548), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U6955 ( .A1(n7621), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5439) );
  OAI211_X1 U6956 ( .C1(n5441), .C2(n7624), .A(n5440), .B(n5439), .ZN(n5442)
         );
  INV_X1 U6957 ( .A(n5442), .ZN(n5443) );
  NAND2_X1 U6958 ( .A1(n5444), .A2(n5443), .ZN(n8108) );
  NAND2_X1 U6959 ( .A1(n8108), .A2(n4250), .ZN(n5445) );
  NOR2_X1 U6960 ( .A1(n5446), .A2(n5445), .ZN(n5447) );
  AOI21_X1 U6961 ( .B1(n5446), .B2(n5445), .A(n5447), .ZN(n7935) );
  NAND2_X1 U6962 ( .A1(n7936), .A2(n7935), .ZN(n7934) );
  INV_X1 U6963 ( .A(n5447), .ZN(n5448) );
  NAND2_X1 U6964 ( .A1(n7934), .A2(n5448), .ZN(n6264) );
  INV_X1 U6965 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7563) );
  INV_X1 U6966 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7543) );
  MUX2_X1 U6967 ( .A(n7563), .B(n7543), .S(n7613), .Z(n5454) );
  INV_X1 U6968 ( .A(SI_27_), .ZN(n5453) );
  NAND2_X1 U6969 ( .A1(n5454), .A2(n5453), .ZN(n5475) );
  INV_X1 U6970 ( .A(n5454), .ZN(n5455) );
  NAND2_X1 U6971 ( .A1(n5455), .A2(SI_27_), .ZN(n5456) );
  NAND2_X1 U6972 ( .A1(n7561), .A2(n7742), .ZN(n5458) );
  NAND2_X1 U6973 ( .A1(n7743), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5457) );
  XNOR2_X1 U6974 ( .A(n8355), .B(n5415), .ZN(n5470) );
  INV_X1 U6975 ( .A(n5470), .ZN(n5472) );
  INV_X1 U6976 ( .A(n5461), .ZN(n5459) );
  NAND2_X1 U6977 ( .A1(n5459), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5481) );
  INV_X1 U6978 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U6979 ( .A1(n5461), .A2(n5460), .ZN(n5462) );
  NAND2_X1 U6980 ( .A1(n5481), .A2(n5462), .ZN(n8152) );
  INV_X1 U6981 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U6982 ( .A1(n5548), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U6983 ( .A1(n7621), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5463) );
  OAI211_X1 U6984 ( .C1(n5465), .C2(n7624), .A(n5464), .B(n5463), .ZN(n5466)
         );
  INV_X1 U6985 ( .A(n5466), .ZN(n5467) );
  NOR2_X1 U6986 ( .A1(n8176), .A2(n5489), .ZN(n5469) );
  INV_X1 U6987 ( .A(n5469), .ZN(n5471) );
  AOI21_X1 U6988 ( .B1(n5472), .B2(n5471), .A(n5538), .ZN(n6265) );
  NAND2_X1 U6989 ( .A1(n6264), .A2(n6265), .ZN(n6263) );
  INV_X1 U6990 ( .A(n6263), .ZN(n5535) );
  INV_X1 U6991 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5477) );
  INV_X1 U6992 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7571) );
  MUX2_X1 U6993 ( .A(n5477), .B(n7571), .S(n7613), .Z(n7600) );
  XNOR2_X1 U6994 ( .A(n7600), .B(SI_28_), .ZN(n7597) );
  NAND2_X1 U6995 ( .A1(n7568), .A2(n7742), .ZN(n5479) );
  NAND2_X1 U6996 ( .A1(n7743), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5478) );
  INV_X1 U6997 ( .A(n5481), .ZN(n5480) );
  NAND2_X1 U6998 ( .A1(n5480), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8124) );
  INV_X1 U6999 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U7000 ( .A1(n5481), .A2(n5547), .ZN(n5482) );
  NAND2_X1 U7001 ( .A1(n8124), .A2(n5482), .ZN(n8140) );
  OR2_X1 U7002 ( .A1(n8140), .A2(n5419), .ZN(n5488) );
  INV_X1 U7003 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U7004 ( .A1(n5548), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U7005 ( .A1(n7621), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5483) );
  OAI211_X1 U7006 ( .C1(n5485), .C2(n7624), .A(n5484), .B(n5483), .ZN(n5486)
         );
  INV_X1 U7007 ( .A(n5486), .ZN(n5487) );
  NOR2_X1 U7008 ( .A1(n8158), .A2(n5489), .ZN(n5491) );
  XNOR2_X1 U7009 ( .A(n5491), .B(n5490), .ZN(n5492) );
  XNOR2_X1 U7010 ( .A(n8350), .B(n5492), .ZN(n5536) );
  INV_X1 U7011 ( .A(n5536), .ZN(n5539) );
  NOR4_X1 U7012 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5496) );
  NOR4_X1 U7013 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5495) );
  NOR4_X1 U7014 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n5494) );
  NOR4_X1 U7015 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5493) );
  NAND4_X1 U7016 ( .A1(n5496), .A2(n5495), .A3(n5494), .A4(n5493), .ZN(n5523)
         );
  NOR4_X1 U7017 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n9467) );
  NOR2_X1 U7018 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .ZN(
        n5499) );
  NOR4_X1 U7019 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5498) );
  NOR4_X1 U7020 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n5497) );
  NAND4_X1 U7021 ( .A1(n9467), .A2(n5499), .A3(n5498), .A4(n5497), .ZN(n5522)
         );
  NAND2_X1 U7022 ( .A1(n5500), .A2(n5531), .ZN(n5501) );
  INV_X1 U7023 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U7024 ( .A1(n5507), .A2(n5503), .ZN(n5510) );
  NAND2_X1 U7025 ( .A1(n5510), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5504) );
  MUX2_X1 U7026 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5504), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5506) );
  INV_X1 U7027 ( .A(n7538), .ZN(n5521) );
  INV_X1 U7028 ( .A(n5507), .ZN(n5508) );
  NAND2_X1 U7029 ( .A1(n5508), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5509) );
  MUX2_X1 U7030 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5509), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5511) );
  NAND2_X1 U7031 ( .A1(n5511), .A2(n5510), .ZN(n7478) );
  NAND2_X1 U7032 ( .A1(n5513), .A2(n5512), .ZN(n5514) );
  NAND2_X1 U7033 ( .A1(n5532), .A2(n5531), .ZN(n5515) );
  NAND2_X1 U7034 ( .A1(n5515), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5517) );
  INV_X1 U7035 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5516) );
  INV_X1 U7036 ( .A(P2_B_REG_SCAN_IN), .ZN(n5518) );
  XOR2_X1 U7037 ( .A(n7392), .B(n5518), .Z(n5519) );
  NAND2_X1 U7038 ( .A1(n7478), .A2(n5519), .ZN(n5520) );
  OAI21_X1 U7039 ( .B1(n5523), .B2(n5522), .A(n9883), .ZN(n6714) );
  INV_X1 U7040 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U7041 ( .A1(n9883), .A2(n5524), .ZN(n5525) );
  NAND2_X1 U7042 ( .A1(n7538), .A2(n7478), .ZN(n9917) );
  INV_X1 U7043 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U7044 ( .A1(n9883), .A2(n5526), .ZN(n5527) );
  NAND2_X1 U7045 ( .A1(n7392), .A2(n7538), .ZN(n9915) );
  AND2_X1 U7046 ( .A1(n6717), .A2(n7063), .ZN(n5528) );
  NAND2_X1 U7047 ( .A1(n6714), .A2(n5528), .ZN(n5542) );
  INV_X1 U7048 ( .A(n7392), .ZN(n5530) );
  NOR2_X1 U7049 ( .A1(n7538), .A2(n7478), .ZN(n5529) );
  XNOR2_X1 U7050 ( .A(n5532), .B(n5531), .ZN(n6404) );
  NOR2_X1 U7051 ( .A1(n9954), .A2(n6532), .ZN(n5534) );
  NAND3_X1 U7052 ( .A1(n5535), .A2(n5539), .A3(n7933), .ZN(n5564) );
  INV_X1 U7053 ( .A(n5538), .ZN(n5537) );
  NAND4_X1 U7054 ( .A1(n6263), .A2(n7933), .A3(n5537), .A4(n5536), .ZN(n5563)
         );
  NAND3_X1 U7055 ( .A1(n5539), .A2(n5538), .A3(n7933), .ZN(n5561) );
  INV_X1 U7056 ( .A(n4866), .ZN(n7798) );
  AND2_X1 U7057 ( .A1(n7761), .A2(n7798), .ZN(n6724) );
  NAND2_X1 U7058 ( .A1(n5555), .A2(n6724), .ZN(n5541) );
  NAND2_X1 U7059 ( .A1(n9946), .A2(n8077), .ZN(n7062) );
  INV_X1 U7060 ( .A(n7062), .ZN(n5540) );
  NAND2_X1 U7061 ( .A1(n5542), .A2(n7062), .ZN(n5546) );
  NAND2_X1 U7062 ( .A1(n6532), .A2(n5543), .ZN(n7060) );
  NAND2_X1 U7063 ( .A1(n7060), .A2(n6404), .ZN(n5544) );
  NOR2_X1 U7064 ( .A1(n6530), .A2(n5544), .ZN(n5545) );
  NAND2_X1 U7065 ( .A1(n5546), .A2(n5545), .ZN(n6585) );
  OAI22_X1 U7066 ( .A1(n8140), .A2(n7925), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5547), .ZN(n5559) );
  OR2_X1 U7067 ( .A1(n8124), .A2(n5419), .ZN(n5554) );
  INV_X1 U7068 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U7069 ( .A1(n5548), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U7070 ( .A1(n7621), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5549) );
  OAI211_X1 U7071 ( .C1(n5551), .C2(n7624), .A(n5550), .B(n5549), .ZN(n5552)
         );
  INV_X1 U7072 ( .A(n5552), .ZN(n5553) );
  INV_X1 U7073 ( .A(n5556), .ZN(n5557) );
  INV_X1 U7074 ( .A(n7890), .ZN(n7864) );
  OAI22_X1 U7075 ( .A1(n8134), .A2(n7939), .B1(n8176), .B2(n7938), .ZN(n5558)
         );
  AOI211_X1 U7076 ( .C1(n8350), .C2(n7929), .A(n5559), .B(n5558), .ZN(n5560)
         );
  NAND3_X1 U7077 ( .A1(n5564), .A2(n5563), .A3(n5562), .ZN(P2_U3222) );
  INV_X2 U7078 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U7079 ( .A(n5962), .ZN(n5573) );
  NAND2_X1 U7080 ( .A1(n5573), .A2(n5572), .ZN(n5981) );
  INV_X1 U7081 ( .A(n5981), .ZN(n5575) );
  NAND2_X1 U7082 ( .A1(n5575), .A2(n5574), .ZN(n5580) );
  INV_X1 U7083 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5577) );
  XNOR2_X2 U7084 ( .A(n5579), .B(n9458), .ZN(n8877) );
  NAND2_X1 U7085 ( .A1(n5580), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5581) );
  NOR2_X1 U7086 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5585) );
  NOR2_X1 U7087 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5584) );
  NOR2_X1 U7088 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5583) );
  NAND4_X1 U7089 ( .A1(n5585), .A2(n5584), .A3(n5583), .A4(n9458), .ZN(n5589)
         );
  NAND4_X1 U7090 ( .A1(n5587), .A2(n5939), .A3(n5997), .A4(n5586), .ZN(n5588)
         );
  NOR2_X1 U7091 ( .A1(n5589), .A2(n5588), .ZN(n5590) );
  INV_X1 U7092 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U7093 ( .A1(n5596), .A2(n5593), .ZN(n5594) );
  NAND2_X1 U7094 ( .A1(n5594), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5595) );
  XNOR2_X1 U7095 ( .A(n5596), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U7096 ( .A1(n5597), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5598) );
  NAND2_X2 U7097 ( .A1(n6187), .A2(n5599), .ZN(n6272) );
  NAND2_X2 U7098 ( .A1(n5600), .A2(n5648), .ZN(n5659) );
  NAND2_X1 U7099 ( .A1(n5611), .A2(n5626), .ZN(n5603) );
  NAND2_X1 U7100 ( .A1(n5603), .A2(n5602), .ZN(n5609) );
  NAND2_X1 U7101 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n5604) );
  AND2_X1 U7102 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n5605) );
  NAND2_X1 U7103 ( .A1(n5611), .A2(n4803), .ZN(n9545) );
  INV_X1 U7104 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5612) );
  XNOR2_X2 U7105 ( .A(n5613), .B(n5612), .ZN(n7850) );
  AND2_X4 U7106 ( .A1(n5615), .A2(n5616), .ZN(n5687) );
  NAND2_X1 U7107 ( .A1(n5687), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U7108 ( .A1(n5711), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5619) );
  AND2_X2 U7109 ( .A1(n7850), .A2(n5615), .ZN(n5685) );
  NAND2_X1 U7110 ( .A1(n5685), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5618) );
  AND2_X4 U7111 ( .A1(n5616), .A2(n5614), .ZN(n5686) );
  NAND2_X1 U7112 ( .A1(n5686), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U7113 ( .A1(n5621), .A2(n6323), .ZN(n5631) );
  INV_X1 U7114 ( .A(n5640), .ZN(n5622) );
  INV_X1 U7115 ( .A(n6272), .ZN(n5632) );
  NAND2_X1 U7116 ( .A1(n5622), .A2(n6272), .ZN(n5643) );
  INV_X1 U7117 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U7118 ( .A1(n7613), .A2(SI_0_), .ZN(n5624) );
  INV_X1 U7119 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5623) );
  XNOR2_X1 U7120 ( .A(n5624), .B(n5623), .ZN(n6348) );
  MUX2_X1 U7121 ( .A(n5628), .B(n6348), .S(n5668), .Z(n9743) );
  OAI22_X1 U7122 ( .A1(n5643), .A2(n9743), .B1(n5628), .B2(n6272), .ZN(n5629)
         );
  INV_X1 U7123 ( .A(n5629), .ZN(n5630) );
  NAND2_X1 U7124 ( .A1(n5632), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5633) );
  OAI21_X1 U7125 ( .B1(n5844), .B2(n9743), .A(n5633), .ZN(n5634) );
  INV_X1 U7126 ( .A(n5634), .ZN(n5637) );
  NAND2_X1 U7127 ( .A1(n6323), .A2(n5635), .ZN(n5636) );
  NAND2_X1 U7128 ( .A1(n5637), .A2(n5636), .ZN(n6442) );
  NAND2_X1 U7129 ( .A1(n6440), .A2(n6442), .ZN(n6441) );
  NAND2_X1 U7130 ( .A1(n5687), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5647) );
  NAND2_X1 U7131 ( .A1(n5685), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U7132 ( .A1(n5711), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U7133 ( .A1(n5701), .A2(n8900), .ZN(n5655) );
  INV_X2 U7134 ( .A(n5844), .ZN(n6242) );
  INV_X1 U7135 ( .A(n5668), .ZN(n5652) );
  INV_X1 U7136 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U7137 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5649) );
  INV_X1 U7138 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U7139 ( .A1(n6242), .A2(n6488), .ZN(n5654) );
  NAND2_X1 U7140 ( .A1(n5655), .A2(n5654), .ZN(n5656) );
  XNOR2_X1 U7141 ( .A(n5656), .B(n6855), .ZN(n5657) );
  NAND2_X1 U7142 ( .A1(n5658), .A2(n6568), .ZN(n6483) );
  INV_X1 U7143 ( .A(n6483), .ZN(n5663) );
  OR2_X1 U7144 ( .A1(n6322), .A2(n5659), .ZN(n5661) );
  NAND2_X1 U7145 ( .A1(n5701), .A2(n6488), .ZN(n5660) );
  NAND2_X1 U7146 ( .A1(n5661), .A2(n5660), .ZN(n6485) );
  NAND2_X1 U7147 ( .A1(n6484), .A2(n6568), .ZN(n5684) );
  NAND2_X1 U7148 ( .A1(n5711), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5667) );
  NAND2_X1 U7149 ( .A1(n5685), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5666) );
  NAND2_X1 U7150 ( .A1(n5686), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U7151 ( .A1(n5687), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U7152 ( .A1(n5701), .A2(n9755), .ZN(n5676) );
  OR2_X1 U7153 ( .A1(n5669), .A2(n9544), .ZN(n5671) );
  INV_X1 U7154 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U7155 ( .A1(n5671), .A2(n5670), .ZN(n5692) );
  INV_X1 U7156 ( .A(n8608), .ZN(n5672) );
  OR2_X1 U7157 ( .A1(n5695), .A2(n6359), .ZN(n5673) );
  OAI211_X2 U7158 ( .C1(n5668), .C2(n6349), .A(n5674), .B(n5673), .ZN(n6575)
         );
  NAND2_X1 U7159 ( .A1(n6242), .A2(n6575), .ZN(n5675) );
  NAND2_X1 U7160 ( .A1(n5676), .A2(n5675), .ZN(n5677) );
  XNOR2_X1 U7161 ( .A(n5677), .B(n6855), .ZN(n5680) );
  OR2_X1 U7162 ( .A1(n9725), .A2(n5659), .ZN(n5679) );
  NAND2_X1 U7163 ( .A1(n5701), .A2(n6575), .ZN(n5678) );
  INV_X1 U7164 ( .A(n5680), .ZN(n5682) );
  NAND2_X1 U7165 ( .A1(n5682), .A2(n5681), .ZN(n5683) );
  AND2_X1 U7166 ( .A1(n6623), .A2(n5683), .ZN(n6569) );
  NAND2_X1 U7167 ( .A1(n5684), .A2(n6569), .ZN(n6572) );
  NAND2_X1 U7168 ( .A1(n6572), .A2(n6623), .ZN(n5709) );
  NAND2_X1 U7169 ( .A1(n5711), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5691) );
  NAND2_X1 U7170 ( .A1(n5685), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5690) );
  NAND2_X1 U7171 ( .A1(n5686), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5689) );
  INV_X1 U7172 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9731) );
  NAND2_X1 U7173 ( .A1(n5687), .A2(n9731), .ZN(n5688) );
  NAND4_X1 U7174 ( .A1(n5691), .A2(n5690), .A3(n5689), .A4(n5688), .ZN(n8899)
         );
  NAND2_X1 U7175 ( .A1(n5701), .A2(n8899), .ZN(n5699) );
  NAND2_X1 U7176 ( .A1(n5692), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5694) );
  INV_X1 U7177 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5693) );
  XNOR2_X1 U7178 ( .A(n5694), .B(n5693), .ZN(n6352) );
  OR2_X1 U7179 ( .A1(n8608), .A2(n6353), .ZN(n5697) );
  OR2_X1 U7180 ( .A1(n5695), .A2(n6363), .ZN(n5696) );
  NAND2_X1 U7181 ( .A1(n6242), .A2(n9713), .ZN(n5698) );
  NAND2_X1 U7182 ( .A1(n5699), .A2(n5698), .ZN(n5700) );
  XNOR2_X1 U7183 ( .A(n5700), .B(n6855), .ZN(n5704) );
  NAND2_X1 U7184 ( .A1(n5701), .A2(n9713), .ZN(n5702) );
  AND2_X1 U7185 ( .A1(n5703), .A2(n5702), .ZN(n5705) );
  NAND2_X1 U7186 ( .A1(n5704), .A2(n5705), .ZN(n5710) );
  INV_X1 U7187 ( .A(n5704), .ZN(n5707) );
  INV_X1 U7188 ( .A(n5705), .ZN(n5706) );
  NAND2_X1 U7189 ( .A1(n5707), .A2(n5706), .ZN(n5708) );
  NAND2_X1 U7190 ( .A1(n5709), .A2(n6624), .ZN(n6627) );
  NAND2_X1 U7191 ( .A1(n6627), .A2(n5710), .ZN(n6645) );
  NAND2_X1 U7192 ( .A1(n8599), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U7193 ( .A1(n8600), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U7194 ( .A1(n5686), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5714) );
  INV_X1 U7195 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5712) );
  XNOR2_X1 U7196 ( .A(n5712), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n6643) );
  NAND2_X1 U7197 ( .A1(n5687), .A2(n6643), .ZN(n5713) );
  NAND4_X1 U7198 ( .A1(n5716), .A2(n5715), .A3(n5714), .A4(n5713), .ZN(n8898)
         );
  NAND2_X1 U7199 ( .A1(n5701), .A2(n8898), .ZN(n5726) );
  NOR2_X1 U7200 ( .A1(n5717), .A2(n9544), .ZN(n5718) );
  MUX2_X1 U7201 ( .A(n9544), .B(n5718), .S(P1_IR_REG_4__SCAN_IN), .Z(n5719) );
  INV_X1 U7202 ( .A(n5719), .ZN(n5722) );
  INV_X1 U7203 ( .A(n5720), .ZN(n5721) );
  NAND2_X1 U7204 ( .A1(n5722), .A2(n5721), .ZN(n6356) );
  OR2_X1 U7205 ( .A1(n8608), .A2(n6357), .ZN(n5724) );
  OR2_X1 U7206 ( .A1(n5695), .A2(n6368), .ZN(n5723) );
  OAI211_X1 U7207 ( .C1(n5668), .C2(n6356), .A(n5724), .B(n5723), .ZN(n6830)
         );
  NAND2_X1 U7208 ( .A1(n6242), .A2(n6830), .ZN(n5725) );
  NAND2_X1 U7209 ( .A1(n5726), .A2(n5725), .ZN(n5727) );
  XNOR2_X1 U7210 ( .A(n5727), .B(n6855), .ZN(n5732) );
  OR2_X1 U7211 ( .A1(n9722), .A2(n5659), .ZN(n5729) );
  NAND2_X1 U7212 ( .A1(n5701), .A2(n6830), .ZN(n5728) );
  NAND2_X1 U7213 ( .A1(n5729), .A2(n5728), .ZN(n5730) );
  XNOR2_X1 U7214 ( .A(n5732), .B(n5730), .ZN(n6646) );
  NAND2_X1 U7215 ( .A1(n6645), .A2(n6646), .ZN(n6644) );
  INV_X1 U7216 ( .A(n5730), .ZN(n5731) );
  NAND2_X1 U7217 ( .A1(n5732), .A2(n5731), .ZN(n5733) );
  NAND2_X1 U7218 ( .A1(n6644), .A2(n5733), .ZN(n7012) );
  NAND2_X1 U7219 ( .A1(n8600), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U7220 ( .A1(n8599), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U7221 ( .A1(n5686), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5738) );
  NAND3_X1 U7222 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5750) );
  INV_X1 U7223 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U7224 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5734) );
  NAND2_X1 U7225 ( .A1(n5735), .A2(n5734), .ZN(n5736) );
  AND2_X1 U7226 ( .A1(n5750), .A2(n5736), .ZN(n7020) );
  NAND2_X1 U7227 ( .A1(n5687), .A2(n7020), .ZN(n5737) );
  NAND4_X1 U7228 ( .A1(n5740), .A2(n5739), .A3(n5738), .A4(n5737), .ZN(n8897)
         );
  NAND2_X1 U7229 ( .A1(n5701), .A2(n8897), .ZN(n5745) );
  OR2_X1 U7230 ( .A1(n5720), .A2(n9544), .ZN(n5741) );
  XNOR2_X1 U7231 ( .A(n5741), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6294) );
  INV_X1 U7232 ( .A(n6294), .ZN(n9655) );
  NAND2_X1 U7233 ( .A1(n8605), .A2(n6360), .ZN(n5743) );
  INV_X1 U7234 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6361) );
  OR2_X1 U7235 ( .A1(n8608), .A2(n6361), .ZN(n5742) );
  NAND2_X1 U7236 ( .A1(n6242), .A2(n6892), .ZN(n5744) );
  NAND2_X1 U7237 ( .A1(n5745), .A2(n5744), .ZN(n5746) );
  XNOR2_X1 U7238 ( .A(n5746), .B(n6855), .ZN(n5770) );
  INV_X1 U7239 ( .A(n8897), .ZN(n7034) );
  OR2_X1 U7240 ( .A1(n7034), .A2(n5659), .ZN(n5748) );
  NAND2_X1 U7241 ( .A1(n5701), .A2(n6892), .ZN(n5747) );
  AND2_X1 U7242 ( .A1(n5748), .A2(n5747), .ZN(n7016) );
  AND2_X1 U7243 ( .A1(n5770), .A2(n7016), .ZN(n5774) );
  NAND2_X1 U7244 ( .A1(n8600), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5755) );
  NAND2_X1 U7245 ( .A1(n5686), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U7246 ( .A1(n8599), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5753) );
  INV_X1 U7247 ( .A(n5750), .ZN(n5749) );
  NAND2_X1 U7248 ( .A1(n5749), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5780) );
  INV_X1 U7249 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9340) );
  NAND2_X1 U7250 ( .A1(n5750), .A2(n9340), .ZN(n5751) );
  AND2_X1 U7251 ( .A1(n5780), .A2(n5751), .ZN(n7036) );
  NAND2_X1 U7252 ( .A1(n5687), .A2(n7036), .ZN(n5752) );
  NAND2_X1 U7253 ( .A1(n5701), .A2(n8896), .ZN(n5761) );
  NAND2_X1 U7254 ( .A1(n5756), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5757) );
  XNOR2_X1 U7255 ( .A(n5757), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6316) );
  AOI22_X1 U7256 ( .A1(n6018), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5652), .B2(
        n6316), .ZN(n5759) );
  NAND2_X1 U7257 ( .A1(n6370), .A2(n8605), .ZN(n5758) );
  NAND2_X1 U7258 ( .A1(n5759), .A2(n5758), .ZN(n6875) );
  NAND2_X1 U7259 ( .A1(n6875), .A2(n6242), .ZN(n5760) );
  NAND2_X1 U7260 ( .A1(n5761), .A2(n5760), .ZN(n5762) );
  XNOR2_X1 U7261 ( .A(n5762), .B(n6855), .ZN(n5765) );
  INV_X1 U7262 ( .A(n8896), .ZN(n6881) );
  OR2_X1 U7263 ( .A1(n6881), .A2(n5659), .ZN(n5764) );
  NAND2_X1 U7264 ( .A1(n5635), .A2(n6875), .ZN(n5763) );
  AND2_X1 U7265 ( .A1(n5764), .A2(n5763), .ZN(n5766) );
  NAND2_X1 U7266 ( .A1(n5765), .A2(n5766), .ZN(n6983) );
  INV_X1 U7267 ( .A(n5765), .ZN(n5768) );
  INV_X1 U7268 ( .A(n5766), .ZN(n5767) );
  NAND2_X1 U7269 ( .A1(n5768), .A2(n5767), .ZN(n5769) );
  NAND2_X1 U7270 ( .A1(n6983), .A2(n5769), .ZN(n7028) );
  INV_X1 U7271 ( .A(n5770), .ZN(n7013) );
  INV_X1 U7272 ( .A(n7016), .ZN(n5771) );
  AND2_X1 U7273 ( .A1(n7013), .A2(n5771), .ZN(n5772) );
  NOR2_X1 U7274 ( .A1(n7028), .A2(n5772), .ZN(n5773) );
  OAI21_X1 U7275 ( .B1(n7012), .B2(n5774), .A(n5773), .ZN(n6982) );
  NAND2_X1 U7276 ( .A1(n6982), .A2(n6983), .ZN(n5796) );
  NAND2_X1 U7277 ( .A1(n6375), .A2(n8605), .ZN(n5777) );
  OR2_X1 U7278 ( .A1(n5756), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U7279 ( .A1(n5798), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5775) );
  XNOR2_X1 U7280 ( .A(n5775), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6419) );
  AOI22_X1 U7281 ( .A1(n6018), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5652), .B2(
        n6419), .ZN(n5776) );
  NAND2_X1 U7282 ( .A1(n5777), .A2(n5776), .ZN(n6998) );
  NAND2_X1 U7283 ( .A1(n6998), .A2(n6242), .ZN(n5787) );
  NAND2_X1 U7284 ( .A1(n8599), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U7285 ( .A1(n8600), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5784) );
  NAND2_X1 U7286 ( .A1(n5686), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5783) );
  INV_X1 U7287 ( .A(n5780), .ZN(n5778) );
  NAND2_X1 U7288 ( .A1(n5778), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5807) );
  INV_X1 U7289 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U7290 ( .A1(n5780), .A2(n5779), .ZN(n5781) );
  AND2_X1 U7291 ( .A1(n5807), .A2(n5781), .ZN(n6992) );
  NAND2_X1 U7292 ( .A1(n5687), .A2(n6992), .ZN(n5782) );
  NAND4_X1 U7293 ( .A1(n5785), .A2(n5784), .A3(n5783), .A4(n5782), .ZN(n8895)
         );
  NAND2_X1 U7294 ( .A1(n5701), .A2(n8895), .ZN(n5786) );
  NAND2_X1 U7295 ( .A1(n5787), .A2(n5786), .ZN(n5788) );
  XNOR2_X1 U7296 ( .A(n5788), .B(n6855), .ZN(n5791) );
  NAND2_X1 U7297 ( .A1(n6998), .A2(n5701), .ZN(n5790) );
  OR2_X1 U7298 ( .A1(n7152), .A2(n5659), .ZN(n5789) );
  AND2_X1 U7299 ( .A1(n5790), .A2(n5789), .ZN(n5792) );
  NAND2_X1 U7300 ( .A1(n5791), .A2(n5792), .ZN(n5797) );
  INV_X1 U7301 ( .A(n5791), .ZN(n5794) );
  INV_X1 U7302 ( .A(n5792), .ZN(n5793) );
  NAND2_X1 U7303 ( .A1(n5794), .A2(n5793), .ZN(n5795) );
  AND2_X1 U7304 ( .A1(n5797), .A2(n5795), .ZN(n6984) );
  NAND2_X1 U7305 ( .A1(n5796), .A2(n6984), .ZN(n6986) );
  NAND2_X1 U7306 ( .A1(n6986), .A2(n5797), .ZN(n5817) );
  NAND2_X1 U7307 ( .A1(n6379), .A2(n8605), .ZN(n5805) );
  NOR2_X1 U7308 ( .A1(n5798), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5801) );
  NOR2_X1 U7309 ( .A1(n5801), .A2(n9544), .ZN(n5799) );
  MUX2_X1 U7310 ( .A(n9544), .B(n5799), .S(P1_IR_REG_8__SCAN_IN), .Z(n5803) );
  NAND2_X1 U7311 ( .A1(n5801), .A2(n5800), .ZN(n5840) );
  INV_X1 U7312 ( .A(n5840), .ZN(n5802) );
  AOI22_X1 U7313 ( .A1(n6018), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5652), .B2(
        n9661), .ZN(n5804) );
  NAND2_X1 U7314 ( .A1(n5805), .A2(n5804), .ZN(n7154) );
  NAND2_X1 U7315 ( .A1(n8599), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U7316 ( .A1(n5686), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U7317 ( .A1(n8600), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5810) );
  INV_X1 U7318 ( .A(n5807), .ZN(n5806) );
  NAND2_X1 U7319 ( .A1(n5806), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5826) );
  INV_X1 U7320 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7149) );
  NAND2_X1 U7321 ( .A1(n5807), .A2(n7149), .ZN(n5808) );
  AND2_X1 U7322 ( .A1(n5826), .A2(n5808), .ZN(n7148) );
  NAND2_X1 U7323 ( .A1(n5687), .A2(n7148), .ZN(n5809) );
  NOR2_X1 U7324 ( .A1(n5659), .A2(n7235), .ZN(n5813) );
  AOI21_X1 U7325 ( .B1(n7154), .B2(n5701), .A(n5813), .ZN(n5818) );
  NAND2_X1 U7326 ( .A1(n5817), .A2(n5818), .ZN(n7144) );
  NAND2_X1 U7327 ( .A1(n7154), .A2(n6242), .ZN(n5815) );
  INV_X1 U7328 ( .A(n7235), .ZN(n8894) );
  NAND2_X1 U7329 ( .A1(n5635), .A2(n8894), .ZN(n5814) );
  NAND2_X1 U7330 ( .A1(n5815), .A2(n5814), .ZN(n5816) );
  XNOR2_X1 U7331 ( .A(n5816), .B(n6240), .ZN(n7147) );
  NAND2_X1 U7332 ( .A1(n7144), .A2(n7147), .ZN(n5821) );
  NAND2_X1 U7333 ( .A1(n5821), .A2(n7145), .ZN(n7227) );
  NAND2_X1 U7334 ( .A1(n6383), .A2(n8605), .ZN(n5824) );
  NAND2_X1 U7335 ( .A1(n5840), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5822) );
  XNOR2_X1 U7336 ( .A(n5822), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6498) );
  AOI22_X1 U7337 ( .A1(n6018), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5652), .B2(
        n6498), .ZN(n5823) );
  NAND2_X1 U7338 ( .A1(n5824), .A2(n5823), .ZN(n8623) );
  NAND2_X1 U7339 ( .A1(n8623), .A2(n6242), .ZN(n5833) );
  NAND2_X1 U7340 ( .A1(n8600), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5831) );
  NAND2_X1 U7341 ( .A1(n5686), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U7342 ( .A1(n8599), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5829) );
  NAND2_X1 U7343 ( .A1(n5826), .A2(n5825), .ZN(n5827) );
  AND2_X1 U7344 ( .A1(n5845), .A2(n5827), .ZN(n7231) );
  NAND2_X1 U7345 ( .A1(n5687), .A2(n7231), .ZN(n5828) );
  NAND4_X1 U7346 ( .A1(n5831), .A2(n5830), .A3(n5829), .A4(n5828), .ZN(n8893)
         );
  NAND2_X1 U7347 ( .A1(n5701), .A2(n8893), .ZN(n5832) );
  NAND2_X1 U7348 ( .A1(n5833), .A2(n5832), .ZN(n5834) );
  XNOR2_X1 U7349 ( .A(n5834), .B(n6855), .ZN(n5837) );
  INV_X1 U7350 ( .A(n8893), .ZN(n7339) );
  NOR2_X1 U7351 ( .A1(n5659), .A2(n7339), .ZN(n5835) );
  AOI21_X1 U7352 ( .B1(n8623), .B2(n5701), .A(n5835), .ZN(n5836) );
  NAND2_X1 U7353 ( .A1(n5837), .A2(n5836), .ZN(n5839) );
  OR2_X1 U7354 ( .A1(n5837), .A2(n5836), .ZN(n5838) );
  NAND2_X1 U7355 ( .A1(n5839), .A2(n5838), .ZN(n7230) );
  NAND2_X1 U7356 ( .A1(n6398), .A2(n8605), .ZN(n5843) );
  NAND2_X1 U7357 ( .A1(n5855), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5841) );
  XNOR2_X1 U7358 ( .A(n5841), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9674) );
  AOI22_X1 U7359 ( .A1(n6018), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5652), .B2(
        n9674), .ZN(n5842) );
  NAND2_X1 U7360 ( .A1(n7121), .A2(n6242), .ZN(n5852) );
  NAND2_X1 U7361 ( .A1(n8600), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U7362 ( .A1(n5686), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U7363 ( .A1(n8599), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5848) );
  NAND2_X1 U7364 ( .A1(n5845), .A2(n7337), .ZN(n5846) );
  AND2_X1 U7365 ( .A1(n5861), .A2(n5846), .ZN(n7341) );
  NAND2_X1 U7366 ( .A1(n5687), .A2(n7341), .ZN(n5847) );
  NAND4_X1 U7367 ( .A1(n5850), .A2(n5849), .A3(n5848), .A4(n5847), .ZN(n8892)
         );
  NAND2_X1 U7368 ( .A1(n5701), .A2(n8892), .ZN(n5851) );
  NAND2_X1 U7369 ( .A1(n5852), .A2(n5851), .ZN(n5853) );
  XNOR2_X1 U7370 ( .A(n5853), .B(n6240), .ZN(n5871) );
  NOR2_X1 U7371 ( .A1(n5659), .A2(n7187), .ZN(n5854) );
  AOI21_X1 U7372 ( .B1(n7121), .B2(n5701), .A(n5854), .ZN(n5872) );
  XNOR2_X1 U7373 ( .A(n5871), .B(n5872), .ZN(n7335) );
  NAND2_X1 U7374 ( .A1(n6389), .A2(n8605), .ZN(n5858) );
  OAI21_X1 U7375 ( .B1(n5855), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5856) );
  XNOR2_X1 U7376 ( .A(n5856), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6934) );
  AOI22_X1 U7377 ( .A1(n6018), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5652), .B2(
        n6934), .ZN(n5857) );
  NAND2_X1 U7378 ( .A1(n5858), .A2(n5857), .ZN(n7193) );
  NAND2_X1 U7379 ( .A1(n7193), .A2(n6242), .ZN(n5868) );
  NAND2_X1 U7380 ( .A1(n8599), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U7381 ( .A1(n8600), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5865) );
  NAND2_X1 U7382 ( .A1(n5686), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5864) );
  INV_X1 U7383 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U7384 ( .A1(n5861), .A2(n5860), .ZN(n5862) );
  AND2_X1 U7385 ( .A1(n5882), .A2(n5862), .ZN(n7384) );
  NAND2_X1 U7386 ( .A1(n5687), .A2(n7384), .ZN(n5863) );
  NAND4_X1 U7387 ( .A1(n5866), .A2(n5865), .A3(n5864), .A4(n5863), .ZN(n8891)
         );
  NAND2_X1 U7388 ( .A1(n5701), .A2(n8891), .ZN(n5867) );
  NAND2_X1 U7389 ( .A1(n5868), .A2(n5867), .ZN(n5869) );
  XNOR2_X1 U7390 ( .A(n5869), .B(n6240), .ZN(n5894) );
  NOR2_X1 U7391 ( .A1(n5659), .A2(n7418), .ZN(n5870) );
  AOI21_X1 U7392 ( .B1(n7193), .B2(n5635), .A(n5870), .ZN(n5892) );
  XNOR2_X1 U7393 ( .A(n5894), .B(n5892), .ZN(n7379) );
  INV_X1 U7394 ( .A(n5871), .ZN(n5873) );
  NAND2_X1 U7395 ( .A1(n5873), .A2(n5872), .ZN(n7377) );
  AND2_X1 U7396 ( .A1(n7379), .A2(n7377), .ZN(n5874) );
  NAND2_X1 U7397 ( .A1(n6409), .A2(n8605), .ZN(n5880) );
  NAND2_X1 U7398 ( .A1(n5875), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5876) );
  MUX2_X1 U7399 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5876), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5878) );
  AOI22_X1 U7400 ( .A1(n6018), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5652), .B2(
        n8934), .ZN(n5879) );
  NAND2_X1 U7401 ( .A1(n9597), .A2(n6242), .ZN(n5889) );
  NAND2_X1 U7402 ( .A1(n8599), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5887) );
  NAND2_X1 U7403 ( .A1(n8600), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U7404 ( .A1(n5686), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5885) );
  INV_X1 U7405 ( .A(n5882), .ZN(n5881) );
  INV_X1 U7406 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7416) );
  NAND2_X1 U7407 ( .A1(n5882), .A2(n7416), .ZN(n5883) );
  AND2_X1 U7408 ( .A1(n5904), .A2(n5883), .ZN(n7420) );
  NAND2_X1 U7409 ( .A1(n5687), .A2(n7420), .ZN(n5884) );
  NAND4_X1 U7410 ( .A1(n5887), .A2(n5886), .A3(n5885), .A4(n5884), .ZN(n8890)
         );
  NAND2_X1 U7411 ( .A1(n5635), .A2(n8890), .ZN(n5888) );
  NAND2_X1 U7412 ( .A1(n5889), .A2(n5888), .ZN(n5890) );
  XNOR2_X1 U7413 ( .A(n5890), .B(n6240), .ZN(n5896) );
  NOR2_X1 U7414 ( .A1(n5659), .A2(n7433), .ZN(n5891) );
  AOI21_X1 U7415 ( .B1(n9597), .B2(n5635), .A(n5891), .ZN(n5897) );
  XNOR2_X1 U7416 ( .A(n5896), .B(n5897), .ZN(n7412) );
  INV_X1 U7417 ( .A(n5892), .ZN(n5893) );
  NAND2_X1 U7418 ( .A1(n5894), .A2(n5893), .ZN(n7413) );
  AND2_X1 U7419 ( .A1(n7412), .A2(n7413), .ZN(n5895) );
  INV_X1 U7420 ( .A(n5896), .ZN(n5898) );
  NAND2_X1 U7421 ( .A1(n5898), .A2(n5897), .ZN(n5899) );
  NAND2_X1 U7422 ( .A1(n6432), .A2(n8605), .ZN(n5902) );
  OR2_X1 U7423 ( .A1(n5877), .A2(n9544), .ZN(n5900) );
  XNOR2_X1 U7424 ( .A(n5900), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7266) );
  AOI22_X1 U7425 ( .A1(n6018), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5652), .B2(
        n7266), .ZN(n5901) );
  NAND2_X1 U7426 ( .A1(n7435), .A2(n6242), .ZN(n5911) );
  NAND2_X1 U7427 ( .A1(n8599), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7428 ( .A1(n8600), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U7429 ( .A1(n5686), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U7430 ( .A1(n5904), .A2(n5903), .ZN(n5905) );
  AND2_X1 U7431 ( .A1(n5923), .A2(n5905), .ZN(n7429) );
  NAND2_X1 U7432 ( .A1(n5687), .A2(n7429), .ZN(n5906) );
  NAND4_X1 U7433 ( .A1(n5909), .A2(n5908), .A3(n5907), .A4(n5906), .ZN(n8889)
         );
  NAND2_X1 U7434 ( .A1(n5701), .A2(n8889), .ZN(n5910) );
  NAND2_X1 U7435 ( .A1(n5911), .A2(n5910), .ZN(n5912) );
  XNOR2_X1 U7436 ( .A(n5912), .B(n6855), .ZN(n5914) );
  NOR2_X1 U7437 ( .A1(n5659), .A2(n9284), .ZN(n5913) );
  AOI21_X1 U7438 ( .B1(n7435), .B2(n5701), .A(n5913), .ZN(n5915) );
  AND2_X1 U7439 ( .A1(n5914), .A2(n5915), .ZN(n7424) );
  INV_X1 U7440 ( .A(n5914), .ZN(n5917) );
  INV_X1 U7441 ( .A(n5915), .ZN(n5916) );
  NAND2_X1 U7442 ( .A1(n5917), .A2(n5916), .ZN(n7425) );
  NAND2_X1 U7443 ( .A1(n6436), .A2(n8605), .ZN(n5920) );
  OR2_X1 U7444 ( .A1(n5918), .A2(n9544), .ZN(n5940) );
  XNOR2_X1 U7445 ( .A(n5940), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7507) );
  AOI22_X1 U7446 ( .A1(n6018), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5652), .B2(
        n7507), .ZN(n5919) );
  NAND2_X1 U7447 ( .A1(n9521), .A2(n6242), .ZN(n5930) );
  NAND2_X1 U7448 ( .A1(n8600), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7449 ( .A1(n5686), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U7450 ( .A1(n8599), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5926) );
  INV_X1 U7451 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U7452 ( .A1(n5923), .A2(n5922), .ZN(n5924) );
  AND2_X1 U7453 ( .A1(n5946), .A2(n5924), .ZN(n9290) );
  NAND2_X1 U7454 ( .A1(n5687), .A2(n9290), .ZN(n5925) );
  NAND4_X1 U7455 ( .A1(n5928), .A2(n5927), .A3(n5926), .A4(n5925), .ZN(n9266)
         );
  NAND2_X1 U7456 ( .A1(n5701), .A2(n9266), .ZN(n5929) );
  NAND2_X1 U7457 ( .A1(n5930), .A2(n5929), .ZN(n5931) );
  XNOR2_X1 U7458 ( .A(n5931), .B(n6855), .ZN(n5935) );
  NAND2_X1 U7459 ( .A1(n5932), .A2(n5935), .ZN(n8470) );
  NAND2_X1 U7460 ( .A1(n9521), .A2(n5635), .ZN(n5934) );
  OR2_X1 U7461 ( .A1(n8985), .A2(n5659), .ZN(n5933) );
  NAND2_X1 U7462 ( .A1(n5934), .A2(n5933), .ZN(n8473) );
  INV_X1 U7463 ( .A(n5935), .ZN(n5936) );
  NAND2_X1 U7464 ( .A1(n5937), .A2(n5936), .ZN(n8471) );
  INV_X1 U7465 ( .A(n8471), .ZN(n5938) );
  NAND2_X1 U7466 ( .A1(n6507), .A2(n8605), .ZN(n5945) );
  NAND2_X1 U7467 ( .A1(n5940), .A2(n5939), .ZN(n5941) );
  NAND2_X1 U7468 ( .A1(n5941), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5943) );
  INV_X1 U7469 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5942) );
  XNOR2_X1 U7470 ( .A(n5943), .B(n5942), .ZN(n7550) );
  INV_X1 U7471 ( .A(n7550), .ZN(n7510) );
  AOI22_X1 U7472 ( .A1(n6018), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5652), .B2(
        n7510), .ZN(n5944) );
  NAND2_X1 U7473 ( .A1(n9514), .A2(n6242), .ZN(n5953) );
  NAND2_X1 U7474 ( .A1(n8600), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U7475 ( .A1(n5686), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5950) );
  NAND2_X1 U7476 ( .A1(n8599), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U7477 ( .A1(n5946), .A2(n7505), .ZN(n5947) );
  AND2_X1 U7478 ( .A1(n5968), .A2(n5947), .ZN(n9272) );
  NAND2_X1 U7479 ( .A1(n5687), .A2(n9272), .ZN(n5948) );
  NAND4_X1 U7480 ( .A1(n5951), .A2(n5950), .A3(n5949), .A4(n5948), .ZN(n8888)
         );
  NAND2_X1 U7481 ( .A1(n5635), .A2(n8888), .ZN(n5952) );
  NAND2_X1 U7482 ( .A1(n5953), .A2(n5952), .ZN(n5954) );
  XNOR2_X1 U7483 ( .A(n5954), .B(n6855), .ZN(n5958) );
  NAND2_X1 U7484 ( .A1(n5957), .A2(n5958), .ZN(n8579) );
  NAND2_X1 U7485 ( .A1(n9514), .A2(n5701), .ZN(n5956) );
  OR2_X1 U7486 ( .A1(n9285), .A2(n5659), .ZN(n5955) );
  NAND2_X1 U7487 ( .A1(n5956), .A2(n5955), .ZN(n8582) );
  NAND2_X1 U7488 ( .A1(n8579), .A2(n8582), .ZN(n5961) );
  INV_X1 U7489 ( .A(n5957), .ZN(n5960) );
  INV_X1 U7490 ( .A(n5958), .ZN(n5959) );
  NAND2_X1 U7491 ( .A1(n5960), .A2(n5959), .ZN(n8580) );
  NAND2_X1 U7492 ( .A1(n6589), .A2(n8605), .ZN(n5965) );
  NAND2_X1 U7493 ( .A1(n5962), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5963) );
  XNOR2_X1 U7494 ( .A(n5963), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8944) );
  AOI22_X1 U7495 ( .A1(n6018), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5652), .B2(
        n8944), .ZN(n5964) );
  NAND2_X1 U7496 ( .A1(n9511), .A2(n6242), .ZN(n5975) );
  NAND2_X1 U7497 ( .A1(n8599), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U7498 ( .A1(n8600), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7499 ( .A1(n5686), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5971) );
  INV_X1 U7500 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U7501 ( .A1(n5968), .A2(n5967), .ZN(n5969) );
  AND2_X1 U7502 ( .A1(n5984), .A2(n5969), .ZN(n9255) );
  NAND2_X1 U7503 ( .A1(n5687), .A2(n9255), .ZN(n5970) );
  NAND4_X1 U7504 ( .A1(n5973), .A2(n5972), .A3(n5971), .A4(n5970), .ZN(n9265)
         );
  NAND2_X1 U7505 ( .A1(n5635), .A2(n9265), .ZN(n5974) );
  NAND2_X1 U7506 ( .A1(n5975), .A2(n5974), .ZN(n5976) );
  XNOR2_X1 U7507 ( .A(n5976), .B(n6855), .ZN(n5979) );
  NOR2_X1 U7508 ( .A1(n5659), .A2(n8645), .ZN(n5977) );
  AOI21_X1 U7509 ( .B1(n9511), .B2(n5701), .A(n5977), .ZN(n5978) );
  XNOR2_X1 U7510 ( .A(n5979), .B(n5978), .ZN(n8513) );
  NAND2_X1 U7511 ( .A1(n5979), .A2(n5978), .ZN(n5980) );
  NAND2_X1 U7512 ( .A1(n6634), .A2(n8605), .ZN(n5983) );
  NAND2_X1 U7513 ( .A1(n5981), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5998) );
  XNOR2_X1 U7514 ( .A(n5998), .B(P1_IR_REG_17__SCAN_IN), .ZN(n8962) );
  AOI22_X1 U7515 ( .A1(n6018), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5652), .B2(
        n8962), .ZN(n5982) );
  NAND2_X1 U7516 ( .A1(n9504), .A2(n6242), .ZN(n5991) );
  INV_X1 U7517 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U7518 ( .A1(n5984), .A2(n8523), .ZN(n5985) );
  AND2_X1 U7519 ( .A1(n6005), .A2(n5985), .ZN(n9237) );
  NAND2_X1 U7520 ( .A1(n9237), .A2(n5687), .ZN(n5989) );
  NAND2_X1 U7521 ( .A1(n8599), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U7522 ( .A1(n5686), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7523 ( .A1(n8600), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5986) );
  NAND4_X1 U7524 ( .A1(n5989), .A2(n5988), .A3(n5987), .A4(n5986), .ZN(n9214)
         );
  NAND2_X1 U7525 ( .A1(n5635), .A2(n9214), .ZN(n5990) );
  NAND2_X1 U7526 ( .A1(n5991), .A2(n5990), .ZN(n5992) );
  XNOR2_X1 U7527 ( .A(n5992), .B(n6240), .ZN(n5994) );
  NOR2_X1 U7528 ( .A1(n5659), .A2(n9252), .ZN(n5993) );
  AOI21_X1 U7529 ( .B1(n9504), .B2(n5701), .A(n5993), .ZN(n5995) );
  XNOR2_X1 U7530 ( .A(n5994), .B(n5995), .ZN(n8521) );
  INV_X1 U7531 ( .A(n5994), .ZN(n5996) );
  NAND2_X1 U7532 ( .A1(n6784), .A2(n8605), .ZN(n6002) );
  NAND2_X1 U7533 ( .A1(n5998), .A2(n5997), .ZN(n5999) );
  NAND2_X1 U7534 ( .A1(n5999), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6000) );
  XNOR2_X1 U7535 ( .A(n6000), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9698) );
  AOI22_X1 U7536 ( .A1(n6018), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5652), .B2(
        n9698), .ZN(n6001) );
  NAND2_X1 U7537 ( .A1(n9499), .A2(n6242), .ZN(n6010) );
  INV_X1 U7538 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9224) );
  INV_X1 U7539 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U7540 ( .A1(n6005), .A2(n6004), .ZN(n6006) );
  NAND2_X1 U7541 ( .A1(n6023), .A2(n6006), .ZN(n9223) );
  OR2_X1 U7542 ( .A1(n9223), .A2(n6247), .ZN(n6008) );
  AOI22_X1 U7543 ( .A1(n8599), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n8600), .B2(
        P1_REG1_REG_18__SCAN_IN), .ZN(n6007) );
  OAI211_X1 U7544 ( .C1(n6217), .C2(n9224), .A(n6008), .B(n6007), .ZN(n9242)
         );
  NAND2_X1 U7545 ( .A1(n9242), .A2(n5635), .ZN(n6009) );
  NAND2_X1 U7546 ( .A1(n6010), .A2(n6009), .ZN(n6011) );
  XNOR2_X1 U7547 ( .A(n6011), .B(n6855), .ZN(n6014) );
  NAND2_X1 U7548 ( .A1(n6015), .A2(n6014), .ZN(n8558) );
  NAND2_X1 U7549 ( .A1(n9499), .A2(n5701), .ZN(n6013) );
  NAND2_X1 U7550 ( .A1(n5621), .A2(n9242), .ZN(n6012) );
  NAND2_X1 U7551 ( .A1(n6013), .A2(n6012), .ZN(n8560) );
  NAND2_X1 U7552 ( .A1(n8558), .A2(n8560), .ZN(n6017) );
  INV_X1 U7553 ( .A(n6016), .ZN(n8557) );
  NAND2_X1 U7554 ( .A1(n6860), .A2(n8605), .ZN(n6020) );
  AOI22_X1 U7555 ( .A1(n6018), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9744), .B2(
        n5652), .ZN(n6019) );
  NAND2_X1 U7556 ( .A1(n9493), .A2(n6242), .ZN(n6028) );
  INV_X1 U7557 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9201) );
  INV_X1 U7558 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U7559 ( .A1(n6023), .A2(n6022), .ZN(n6024) );
  NAND2_X1 U7560 ( .A1(n6035), .A2(n6024), .ZN(n9200) );
  OR2_X1 U7561 ( .A1(n9200), .A2(n6247), .ZN(n6026) );
  AOI22_X1 U7562 ( .A1(n8599), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n8600), .B2(
        P1_REG1_REG_19__SCAN_IN), .ZN(n6025) );
  OAI211_X1 U7563 ( .C1(n6217), .C2(n9201), .A(n6026), .B(n6025), .ZN(n9215)
         );
  NAND2_X1 U7564 ( .A1(n9215), .A2(n5701), .ZN(n6027) );
  NAND2_X1 U7565 ( .A1(n6028), .A2(n6027), .ZN(n6029) );
  XNOR2_X1 U7566 ( .A(n6029), .B(n6855), .ZN(n6032) );
  AND2_X1 U7567 ( .A1(n9215), .A2(n5621), .ZN(n6030) );
  AOI21_X1 U7568 ( .B1(n9493), .B2(n5635), .A(n6030), .ZN(n6031) );
  XNOR2_X1 U7569 ( .A(n6032), .B(n6031), .ZN(n8490) );
  NAND2_X1 U7570 ( .A1(n7023), .A2(n8605), .ZN(n6034) );
  OR2_X1 U7571 ( .A1(n8608), .A2(n9348), .ZN(n6033) );
  NAND2_X1 U7572 ( .A1(n9487), .A2(n6242), .ZN(n6044) );
  INV_X1 U7573 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8541) );
  NAND2_X1 U7574 ( .A1(n6035), .A2(n8541), .ZN(n6036) );
  NAND2_X1 U7575 ( .A1(n6055), .A2(n6036), .ZN(n9180) );
  OR2_X1 U7576 ( .A1(n9180), .A2(n6247), .ZN(n6042) );
  INV_X1 U7577 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9454) );
  NAND2_X1 U7578 ( .A1(n5686), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U7579 ( .A1(n8599), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6037) );
  OAI211_X1 U7580 ( .C1(n6039), .C2(n9454), .A(n6038), .B(n6037), .ZN(n6040)
         );
  INV_X1 U7581 ( .A(n6040), .ZN(n6041) );
  NAND2_X1 U7582 ( .A1(n6042), .A2(n6041), .ZN(n9168) );
  NAND2_X1 U7583 ( .A1(n9168), .A2(n5635), .ZN(n6043) );
  NAND2_X1 U7584 ( .A1(n6044), .A2(n6043), .ZN(n6045) );
  XNOR2_X1 U7585 ( .A(n6045), .B(n6240), .ZN(n6048) );
  NAND2_X1 U7586 ( .A1(n9487), .A2(n5701), .ZN(n6047) );
  NAND2_X1 U7587 ( .A1(n9168), .A2(n5621), .ZN(n6046) );
  NAND2_X1 U7588 ( .A1(n6047), .A2(n6046), .ZN(n6049) );
  NAND2_X1 U7589 ( .A1(n6048), .A2(n6049), .ZN(n8537) );
  INV_X1 U7590 ( .A(n6048), .ZN(n6051) );
  INV_X1 U7591 ( .A(n6049), .ZN(n6050) );
  NAND2_X1 U7592 ( .A1(n6051), .A2(n6050), .ZN(n8538) );
  NAND2_X1 U7593 ( .A1(n7046), .A2(n8605), .ZN(n6053) );
  OR2_X1 U7594 ( .A1(n8608), .A2(n7047), .ZN(n6052) );
  NAND2_X1 U7595 ( .A1(n9483), .A2(n6242), .ZN(n6063) );
  INV_X1 U7596 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U7597 ( .A1(n6055), .A2(n6054), .ZN(n6056) );
  AND2_X1 U7598 ( .A1(n6074), .A2(n6056), .ZN(n9171) );
  NAND2_X1 U7599 ( .A1(n9171), .A2(n5687), .ZN(n6061) );
  INV_X1 U7600 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9173) );
  NAND2_X1 U7601 ( .A1(n8599), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7602 ( .A1(n8600), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6057) );
  OAI211_X1 U7603 ( .C1(n6217), .C2(n9173), .A(n6058), .B(n6057), .ZN(n6059)
         );
  INV_X1 U7604 ( .A(n6059), .ZN(n6060) );
  NAND2_X1 U7605 ( .A1(n6061), .A2(n6060), .ZN(n9186) );
  NAND2_X1 U7606 ( .A1(n9186), .A2(n5635), .ZN(n6062) );
  NAND2_X1 U7607 ( .A1(n6063), .A2(n6062), .ZN(n6064) );
  XNOR2_X1 U7608 ( .A(n6064), .B(n6240), .ZN(n6066) );
  AND2_X1 U7609 ( .A1(n9186), .A2(n5621), .ZN(n6065) );
  AOI21_X1 U7610 ( .B1(n9483), .B2(n5701), .A(n6065), .ZN(n6067) );
  XNOR2_X1 U7611 ( .A(n6066), .B(n6067), .ZN(n8497) );
  NAND2_X1 U7612 ( .A1(n8496), .A2(n8497), .ZN(n6070) );
  INV_X1 U7613 ( .A(n6066), .ZN(n6068) );
  NAND2_X1 U7614 ( .A1(n6068), .A2(n6067), .ZN(n6069) );
  NAND2_X1 U7615 ( .A1(n7239), .A2(n8605), .ZN(n6072) );
  OR2_X1 U7616 ( .A1(n8608), .A2(n7240), .ZN(n6071) );
  INV_X1 U7617 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9457) );
  NAND2_X1 U7618 ( .A1(n6074), .A2(n9457), .ZN(n6075) );
  NAND2_X1 U7619 ( .A1(n6091), .A2(n6075), .ZN(n9148) );
  OR2_X1 U7620 ( .A1(n9148), .A2(n6247), .ZN(n6080) );
  INV_X1 U7621 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9149) );
  NAND2_X1 U7622 ( .A1(n8599), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7623 ( .A1(n8600), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6076) );
  OAI211_X1 U7624 ( .C1(n6217), .C2(n9149), .A(n6077), .B(n6076), .ZN(n6078)
         );
  INV_X1 U7625 ( .A(n6078), .ZN(n6079) );
  NAND2_X1 U7626 ( .A1(n6080), .A2(n6079), .ZN(n9167) );
  AND2_X1 U7627 ( .A1(n9167), .A2(n5621), .ZN(n6081) );
  AOI21_X1 U7628 ( .B1(n9479), .B2(n5701), .A(n6081), .ZN(n6085) );
  NAND2_X1 U7629 ( .A1(n9479), .A2(n6242), .ZN(n6083) );
  NAND2_X1 U7630 ( .A1(n9167), .A2(n5635), .ZN(n6082) );
  NAND2_X1 U7631 ( .A1(n6083), .A2(n6082), .ZN(n6084) );
  XNOR2_X1 U7632 ( .A(n6084), .B(n6240), .ZN(n8550) );
  INV_X1 U7633 ( .A(n6085), .ZN(n6086) );
  NAND2_X1 U7634 ( .A1(n7241), .A2(n8605), .ZN(n6088) );
  OR2_X1 U7635 ( .A1(n8608), .A2(n7244), .ZN(n6087) );
  NAND2_X1 U7636 ( .A1(n9473), .A2(n6242), .ZN(n6099) );
  INV_X1 U7637 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7638 ( .A1(n6091), .A2(n6090), .ZN(n6092) );
  NAND2_X1 U7639 ( .A1(n6108), .A2(n6092), .ZN(n9133) );
  OR2_X1 U7640 ( .A1(n9133), .A2(n6247), .ZN(n6097) );
  INV_X1 U7641 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9134) );
  NAND2_X1 U7642 ( .A1(n8599), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7643 ( .A1(n8600), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6093) );
  OAI211_X1 U7644 ( .C1(n9134), .C2(n6217), .A(n6094), .B(n6093), .ZN(n6095)
         );
  INV_X1 U7645 ( .A(n6095), .ZN(n6096) );
  NAND2_X1 U7646 ( .A1(n6097), .A2(n6096), .ZN(n9121) );
  NAND2_X1 U7647 ( .A1(n9121), .A2(n5701), .ZN(n6098) );
  NAND2_X1 U7648 ( .A1(n6099), .A2(n6098), .ZN(n6100) );
  XNOR2_X1 U7649 ( .A(n6100), .B(n6240), .ZN(n6102) );
  AND2_X1 U7650 ( .A1(n9121), .A2(n5621), .ZN(n6101) );
  AOI21_X1 U7651 ( .B1(n9473), .B2(n5701), .A(n6101), .ZN(n8481) );
  NAND2_X1 U7652 ( .A1(n8480), .A2(n8481), .ZN(n8530) );
  INV_X1 U7653 ( .A(n6102), .ZN(n6104) );
  NAND2_X1 U7655 ( .A1(n7387), .A2(n8605), .ZN(n6106) );
  INV_X1 U7656 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7388) );
  OR2_X1 U7657 ( .A1(n8608), .A2(n7388), .ZN(n6105) );
  NAND2_X1 U7658 ( .A1(n9327), .A2(n6242), .ZN(n6117) );
  INV_X1 U7659 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7660 ( .A1(n6108), .A2(n6107), .ZN(n6109) );
  AND2_X1 U7661 ( .A1(n6131), .A2(n6109), .ZN(n9112) );
  NAND2_X1 U7662 ( .A1(n9112), .A2(n5687), .ZN(n6115) );
  INV_X1 U7663 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7664 ( .A1(n8599), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7665 ( .A1(n8600), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6110) );
  OAI211_X1 U7666 ( .C1(n6112), .C2(n6217), .A(n6111), .B(n6110), .ZN(n6113)
         );
  INV_X1 U7667 ( .A(n6113), .ZN(n6114) );
  NAND2_X1 U7668 ( .A1(n9127), .A2(n5635), .ZN(n6116) );
  NAND2_X1 U7669 ( .A1(n6117), .A2(n6116), .ZN(n6118) );
  XNOR2_X1 U7670 ( .A(n6118), .B(n6855), .ZN(n6120) );
  AND2_X1 U7671 ( .A1(n9127), .A2(n5621), .ZN(n6119) );
  AOI21_X1 U7672 ( .B1(n9327), .B2(n5635), .A(n6119), .ZN(n6121) );
  NAND2_X1 U7673 ( .A1(n6120), .A2(n6121), .ZN(n6125) );
  INV_X1 U7674 ( .A(n6120), .ZN(n6123) );
  INV_X1 U7675 ( .A(n6121), .ZN(n6122) );
  NAND2_X1 U7676 ( .A1(n6123), .A2(n6122), .ZN(n6124) );
  NAND2_X1 U7677 ( .A1(n6125), .A2(n6124), .ZN(n8528) );
  INV_X1 U7678 ( .A(n6125), .ZN(n6126) );
  NAND2_X1 U7679 ( .A1(n7477), .A2(n8605), .ZN(n6128) );
  OR2_X1 U7680 ( .A1(n8608), .A2(n7483), .ZN(n6127) );
  INV_X1 U7681 ( .A(n6131), .ZN(n6129) );
  INV_X1 U7682 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U7683 ( .A1(n6131), .A2(n6130), .ZN(n6132) );
  NAND2_X1 U7684 ( .A1(n6144), .A2(n6132), .ZN(n9099) );
  INV_X1 U7685 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7686 ( .A1(n8599), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U7687 ( .A1(n8600), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6133) );
  OAI211_X1 U7688 ( .C1(n6135), .C2(n6217), .A(n6134), .B(n6133), .ZN(n6136)
         );
  INV_X1 U7689 ( .A(n6136), .ZN(n6137) );
  AOI22_X1 U7690 ( .A1(n9321), .A2(n5701), .B1(n5621), .B2(n9120), .ZN(n6156)
         );
  NAND2_X1 U7691 ( .A1(n9321), .A2(n6242), .ZN(n6140) );
  NAND2_X1 U7692 ( .A1(n9120), .A2(n5635), .ZN(n6139) );
  NAND2_X1 U7693 ( .A1(n6140), .A2(n6139), .ZN(n6141) );
  XNOR2_X1 U7694 ( .A(n6141), .B(n6240), .ZN(n6158) );
  XOR2_X1 U7695 ( .A(n6156), .B(n6158), .Z(n8503) );
  NAND2_X1 U7696 ( .A1(n7536), .A2(n8605), .ZN(n6143) );
  OR2_X1 U7697 ( .A1(n8608), .A2(n7539), .ZN(n6142) );
  NAND2_X1 U7698 ( .A1(n9316), .A2(n6242), .ZN(n6153) );
  INV_X1 U7699 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8572) );
  NAND2_X1 U7700 ( .A1(n6144), .A2(n8572), .ZN(n6145) );
  NAND2_X1 U7701 ( .A1(n9085), .A2(n5687), .ZN(n6151) );
  INV_X1 U7702 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7703 ( .A1(n8599), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7704 ( .A1(n8600), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6146) );
  OAI211_X1 U7705 ( .C1(n6217), .C2(n6148), .A(n6147), .B(n6146), .ZN(n6149)
         );
  INV_X1 U7706 ( .A(n6149), .ZN(n6150) );
  NAND2_X1 U7707 ( .A1(n9105), .A2(n5701), .ZN(n6152) );
  NAND2_X1 U7708 ( .A1(n6153), .A2(n6152), .ZN(n6154) );
  XNOR2_X1 U7709 ( .A(n6154), .B(n6855), .ZN(n6160) );
  AND2_X1 U7710 ( .A1(n9105), .A2(n5621), .ZN(n6155) );
  AOI21_X1 U7711 ( .B1(n9316), .B2(n5701), .A(n6155), .ZN(n6161) );
  XNOR2_X1 U7712 ( .A(n6160), .B(n6161), .ZN(n8567) );
  INV_X1 U7713 ( .A(n6156), .ZN(n6157) );
  NOR2_X1 U7714 ( .A1(n6158), .A2(n6157), .ZN(n8568) );
  INV_X1 U7715 ( .A(n6160), .ZN(n6163) );
  INV_X1 U7716 ( .A(n6161), .ZN(n6162) );
  NAND2_X1 U7717 ( .A1(n7561), .A2(n8605), .ZN(n6165) );
  OR2_X1 U7718 ( .A1(n8608), .A2(n7543), .ZN(n6164) );
  NAND2_X1 U7719 ( .A1(n9311), .A2(n6242), .ZN(n6173) );
  XNOR2_X1 U7720 ( .A(n6211), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9073) );
  NAND2_X1 U7721 ( .A1(n9073), .A2(n5687), .ZN(n6171) );
  INV_X1 U7722 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7723 ( .A1(n8599), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U7724 ( .A1(n8600), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6166) );
  OAI211_X1 U7725 ( .C1(n6168), .C2(n6217), .A(n6167), .B(n6166), .ZN(n6169)
         );
  INV_X1 U7726 ( .A(n6169), .ZN(n6170) );
  NAND2_X1 U7727 ( .A1(n9090), .A2(n5635), .ZN(n6172) );
  NAND2_X1 U7728 ( .A1(n6173), .A2(n6172), .ZN(n6174) );
  XNOR2_X1 U7729 ( .A(n6174), .B(n6855), .ZN(n6177) );
  AND2_X1 U7730 ( .A1(n9090), .A2(n5621), .ZN(n6175) );
  AOI21_X1 U7731 ( .B1(n9311), .B2(n5701), .A(n6175), .ZN(n6176) );
  NAND2_X1 U7732 ( .A1(n6177), .A2(n6176), .ZN(n6256) );
  OAI21_X1 U7733 ( .B1(n6177), .B2(n6176), .A(n6256), .ZN(n6179) );
  INV_X1 U7734 ( .A(n6178), .ZN(n6181) );
  INV_X1 U7735 ( .A(n6179), .ZN(n6180) );
  AOI21_X1 U7736 ( .B1(n4275), .B2(n6181), .A(n6180), .ZN(n6207) );
  INV_X1 U7737 ( .A(n6182), .ZN(n7481) );
  INV_X1 U7738 ( .A(n6183), .ZN(n7389) );
  NAND3_X1 U7739 ( .A1(n7481), .A2(P1_B_REG_SCAN_IN), .A3(n7389), .ZN(n6185)
         );
  INV_X1 U7740 ( .A(P1_B_REG_SCAN_IN), .ZN(n8974) );
  NAND2_X1 U7741 ( .A1(n6183), .A2(n8974), .ZN(n6184) );
  INV_X1 U7742 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6186) );
  NAND2_X1 U7743 ( .A1(n9764), .A2(n6186), .ZN(n6189) );
  INV_X1 U7744 ( .A(n6187), .ZN(n7541) );
  NAND2_X1 U7745 ( .A1(n7541), .A2(n7389), .ZN(n6188) );
  INV_X1 U7746 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9455) );
  NAND2_X1 U7747 ( .A1(n9764), .A2(n9455), .ZN(n6191) );
  NAND2_X1 U7748 ( .A1(n7541), .A2(n7481), .ZN(n6190) );
  NOR2_X1 U7749 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .ZN(
        n9464) );
  NOR4_X1 U7750 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6194) );
  NOR4_X1 U7751 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6193) );
  NOR4_X1 U7752 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6192) );
  AND4_X1 U7753 ( .A1(n9464), .A2(n6194), .A3(n6193), .A4(n6192), .ZN(n6200)
         );
  NOR4_X1 U7754 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6198) );
  NOR4_X1 U7755 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6197) );
  NOR4_X1 U7756 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n6196) );
  NOR4_X1 U7757 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6195) );
  AND4_X1 U7758 ( .A1(n6198), .A2(n6197), .A3(n6196), .A4(n6195), .ZN(n6199)
         );
  NAND2_X1 U7759 ( .A1(n6200), .A2(n6199), .ZN(n6201) );
  NAND2_X1 U7760 ( .A1(n9764), .A2(n6201), .ZN(n6337) );
  NAND3_X1 U7761 ( .A1(n6472), .A2(n9542), .A3(n6337), .ZN(n6223) );
  NAND2_X1 U7762 ( .A1(n6202), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6203) );
  XNOR2_X1 U7763 ( .A(n6203), .B(n5591), .ZN(n7242) );
  AND2_X1 U7764 ( .A1(n7242), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6204) );
  NOR2_X1 U7765 ( .A1(n6223), .A2(n9765), .ZN(n6232) );
  OAI21_X1 U7766 ( .B1(n6246), .B2(n6207), .A(n8571), .ZN(n6235) );
  NAND3_X1 U7767 ( .A1(n5622), .A2(n6206), .A3(n5638), .ZN(n8757) );
  INV_X1 U7768 ( .A(n6232), .ZN(n6208) );
  NOR2_X1 U7769 ( .A1(n8757), .A2(n6208), .ZN(n6227) );
  INV_X1 U7770 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6210) );
  INV_X1 U7771 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6253) );
  OAI21_X1 U7772 ( .B1(n6211), .B2(n6210), .A(n6253), .ZN(n6214) );
  INV_X1 U7773 ( .A(n6211), .ZN(n6213) );
  AND2_X1 U7774 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6212) );
  NAND2_X1 U7775 ( .A1(n6213), .A2(n6212), .ZN(n9043) );
  NAND2_X1 U7776 ( .A1(n6214), .A2(n9043), .ZN(n9054) );
  INV_X1 U7777 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9053) );
  NAND2_X1 U7778 ( .A1(n8599), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7779 ( .A1(n8600), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6215) );
  OAI211_X1 U7780 ( .C1(n9053), .C2(n6217), .A(n6216), .B(n6215), .ZN(n6218)
         );
  INV_X1 U7781 ( .A(n6218), .ZN(n6219) );
  AND3_X1 U7782 ( .A1(n6336), .A2(n6272), .A3(n7242), .ZN(n6221) );
  NAND2_X1 U7783 ( .A1(n9817), .A2(n6223), .ZN(n6477) );
  NAND2_X1 U7784 ( .A1(n6221), .A2(n6477), .ZN(n6222) );
  NAND2_X1 U7785 ( .A1(n6222), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6226) );
  OR2_X1 U7786 ( .A1(n6469), .A2(n8877), .ZN(n9740) );
  INV_X1 U7787 ( .A(n9740), .ZN(n6225) );
  AND2_X1 U7788 ( .A1(n6223), .A2(n9541), .ZN(n6224) );
  NAND2_X1 U7789 ( .A1(n6225), .A2(n6224), .ZN(n6478) );
  INV_X1 U7790 ( .A(n9073), .ZN(n6229) );
  INV_X1 U7791 ( .A(n6209), .ZN(n6443) );
  AOI22_X1 U7792 ( .A1(n9105), .A2(n8585), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n6228) );
  OAI21_X1 U7793 ( .B1(n8563), .B2(n6229), .A(n6228), .ZN(n6230) );
  AOI21_X1 U7794 ( .B1(n8552), .B2(n9078), .A(n6230), .ZN(n6234) );
  NOR2_X1 U7795 ( .A1(n9765), .A2(n5638), .ZN(n6231) );
  NAND2_X1 U7796 ( .A1(n6225), .A2(n6232), .ZN(n6233) );
  NAND3_X1 U7797 ( .A1(n6235), .A2(n6234), .A3(n4800), .ZN(P1_U3212) );
  NAND2_X1 U7798 ( .A1(n7568), .A2(n8605), .ZN(n6237) );
  OR2_X1 U7799 ( .A1(n8608), .A2(n7571), .ZN(n6236) );
  NAND2_X1 U7800 ( .A1(n9307), .A2(n5701), .ZN(n6239) );
  NAND2_X1 U7801 ( .A1(n9078), .A2(n5621), .ZN(n6238) );
  NAND2_X1 U7802 ( .A1(n6239), .A2(n6238), .ZN(n6241) );
  XNOR2_X1 U7803 ( .A(n6241), .B(n6240), .ZN(n6244) );
  AOI22_X1 U7804 ( .A1(n9307), .A2(n6242), .B1(n5635), .B2(n9078), .ZN(n6243)
         );
  XNOR2_X1 U7805 ( .A(n6244), .B(n6243), .ZN(n6245) );
  INV_X1 U7806 ( .A(n6245), .ZN(n6257) );
  NAND3_X1 U7807 ( .A1(n6246), .A2(n6245), .A3(n8571), .ZN(n6261) );
  INV_X1 U7808 ( .A(n8585), .ZN(n8573) );
  OR2_X1 U7809 ( .A1(n9043), .A2(n6247), .ZN(n6252) );
  NAND2_X1 U7810 ( .A1(n5686), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U7811 ( .A1(n8599), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6249) );
  NAND2_X1 U7812 ( .A1(n8600), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6248) );
  AND3_X1 U7813 ( .A1(n6250), .A2(n6249), .A3(n6248), .ZN(n6251) );
  NAND2_X1 U7814 ( .A1(n6252), .A2(n6251), .ZN(n9062) );
  OAI22_X1 U7815 ( .A1(n9054), .A2(n8563), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6253), .ZN(n6254) );
  AOI21_X1 U7816 ( .B1(n8552), .B2(n9062), .A(n6254), .ZN(n6255) );
  OAI21_X1 U7817 ( .B1(n9007), .B2(n8573), .A(n6255), .ZN(n6259) );
  NOR3_X1 U7818 ( .A1(n6257), .A2(n8592), .A3(n6256), .ZN(n6258) );
  AOI211_X1 U7819 ( .C1(n9307), .C2(n8590), .A(n6259), .B(n6258), .ZN(n6260)
         );
  NAND3_X1 U7820 ( .A1(n6262), .A2(n6261), .A3(n6260), .ZN(P1_U3218) );
  OAI211_X1 U7821 ( .C1(n6265), .C2(n6264), .A(n6263), .B(n7933), .ZN(n6269)
         );
  NOR2_X1 U7822 ( .A1(n7925), .A2(n8152), .ZN(n6267) );
  INV_X1 U7823 ( .A(n8108), .ZN(n8157) );
  OAI22_X1 U7824 ( .A1(n8158), .A2(n7939), .B1(n8157), .B2(n7938), .ZN(n6266)
         );
  AOI211_X1 U7825 ( .C1(P2_REG3_REG_27__SCAN_IN), .C2(P2_U3152), .A(n6267), 
        .B(n6266), .ZN(n6268) );
  NAND3_X1 U7826 ( .A1(n6269), .A2(n6268), .A3(n4801), .ZN(P2_U3216) );
  INV_X1 U7827 ( .A(n7242), .ZN(n6270) );
  NAND2_X1 U7828 ( .A1(n8718), .A2(n6272), .ZN(n6273) );
  NAND2_X1 U7829 ( .A1(n6273), .A2(n7242), .ZN(n8965) );
  NAND2_X1 U7830 ( .A1(n8965), .A2(n5668), .ZN(n9618) );
  NAND2_X1 U7831 ( .A1(n9618), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AND2_X1 U7832 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7232) );
  INV_X1 U7833 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6274) );
  MUX2_X1 U7834 ( .A(n6274), .B(P1_REG2_REG_9__SCAN_IN), .S(n6498), .Z(n6284)
         );
  INV_X1 U7835 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7003) );
  XNOR2_X1 U7836 ( .A(n6381), .B(n7003), .ZN(n9668) );
  NOR2_X1 U7837 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6419), .ZN(n6275) );
  AOI21_X1 U7838 ( .B1(n6419), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6275), .ZN(
        n6413) );
  INV_X1 U7839 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9415) );
  MUX2_X1 U7840 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9415), .S(n6316), .Z(n6308)
         );
  NOR2_X1 U7841 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6294), .ZN(n6276) );
  AOI21_X1 U7842 ( .B1(n6294), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6276), .ZN(
        n9645) );
  INV_X1 U7843 ( .A(n6356), .ZN(n9631) );
  INV_X1 U7844 ( .A(n6352), .ZN(n8914) );
  INV_X1 U7845 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6278) );
  INV_X1 U7846 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U7847 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6447) );
  INV_X1 U7848 ( .A(n6447), .ZN(n8904) );
  MUX2_X1 U7849 ( .A(n6278), .B(P1_REG2_REG_2__SCAN_IN), .S(n6349), .Z(n6454)
         );
  NAND2_X1 U7850 ( .A1(n6453), .A2(n6454), .ZN(n6452) );
  OAI21_X1 U7851 ( .B1(n6349), .B2(n6278), .A(n6452), .ZN(n8916) );
  XNOR2_X1 U7852 ( .A(n6352), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n8917) );
  NAND2_X1 U7853 ( .A1(n8916), .A2(n8917), .ZN(n8915) );
  XNOR2_X1 U7854 ( .A(n6356), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9629) );
  NAND2_X1 U7855 ( .A1(n9645), .A2(n9646), .ZN(n9644) );
  OAI21_X1 U7856 ( .B1(n6294), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9644), .ZN(
        n6279) );
  INV_X1 U7857 ( .A(n6279), .ZN(n6307) );
  AND2_X1 U7858 ( .A1(n6308), .A2(n6307), .ZN(n6309) );
  NOR2_X1 U7859 ( .A1(n6283), .A2(n6284), .ZN(n6491) );
  OR2_X1 U7860 ( .A1(n6209), .A2(P1_U3084), .ZN(n7569) );
  NOR2_X1 U7861 ( .A1(n7569), .A2(n8975), .ZN(n6282) );
  AOI211_X1 U7862 ( .C1(n6284), .C2(n6283), .A(n6491), .B(n9679), .ZN(n6306)
         );
  NOR2_X1 U7863 ( .A1(n7569), .A2(n6281), .ZN(n6285) );
  XNOR2_X1 U7864 ( .A(n6381), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n9664) );
  OR2_X1 U7865 ( .A1(n6419), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6297) );
  NOR2_X1 U7866 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6419), .ZN(n6286) );
  AOI21_X1 U7867 ( .B1(n6419), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6286), .ZN(
        n6415) );
  INV_X1 U7868 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9831) );
  MUX2_X1 U7869 ( .A(n9831), .B(P1_REG1_REG_2__SCAN_IN), .S(n6349), .Z(n6457)
         );
  INV_X1 U7870 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9829) );
  MUX2_X1 U7871 ( .A(n9829), .B(P1_REG1_REG_1__SCAN_IN), .S(n6351), .Z(n8908)
         );
  AND2_X1 U7872 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n8907) );
  NAND2_X1 U7873 ( .A1(n8908), .A2(n8907), .ZN(n8906) );
  NAND2_X1 U7874 ( .A1(n5651), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U7875 ( .A1(n8906), .A2(n6287), .ZN(n6456) );
  NAND2_X1 U7876 ( .A1(n6457), .A2(n6456), .ZN(n6455) );
  INV_X1 U7877 ( .A(n6349), .ZN(n6451) );
  NAND2_X1 U7878 ( .A1(n6451), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7879 ( .A1(n6455), .A2(n6288), .ZN(n8919) );
  INV_X1 U7880 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6289) );
  OR2_X1 U7881 ( .A1(n6352), .A2(n6289), .ZN(n9632) );
  NAND2_X1 U7882 ( .A1(n6352), .A2(n6289), .ZN(n6290) );
  AND2_X1 U7883 ( .A1(n9632), .A2(n6290), .ZN(n8920) );
  AND2_X1 U7884 ( .A1(n8919), .A2(n8920), .ZN(n9634) );
  INV_X1 U7885 ( .A(n9634), .ZN(n8918) );
  XNOR2_X1 U7886 ( .A(n6356), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9636) );
  AND2_X1 U7887 ( .A1(n9636), .A2(n9632), .ZN(n6291) );
  NAND2_X1 U7888 ( .A1(n8918), .A2(n6291), .ZN(n9635) );
  INV_X1 U7889 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6292) );
  NAND2_X1 U7890 ( .A1(n6356), .A2(n6292), .ZN(n6293) );
  NAND2_X1 U7891 ( .A1(n9635), .A2(n6293), .ZN(n9651) );
  NAND2_X1 U7892 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6294), .ZN(n6295) );
  OAI21_X1 U7893 ( .B1(n6294), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6295), .ZN(
        n9650) );
  OR2_X1 U7894 ( .A1(n9651), .A2(n9650), .ZN(n9647) );
  AND2_X1 U7895 ( .A1(n9647), .A2(n6295), .ZN(n6313) );
  INV_X1 U7896 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6296) );
  XNOR2_X1 U7897 ( .A(n6316), .B(n6296), .ZN(n6314) );
  NAND2_X1 U7898 ( .A1(n6313), .A2(n6314), .ZN(n6312) );
  OAI21_X1 U7899 ( .B1(n6316), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6312), .ZN(
        n6416) );
  NAND2_X1 U7900 ( .A1(n6415), .A2(n6416), .ZN(n6414) );
  AND2_X1 U7901 ( .A1(n6297), .A2(n6414), .ZN(n9663) );
  NAND2_X1 U7902 ( .A1(n9664), .A2(n9663), .ZN(n9662) );
  NAND2_X1 U7903 ( .A1(n9661), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6298) );
  AND2_X1 U7904 ( .A1(n9662), .A2(n6298), .ZN(n6301) );
  NOR2_X1 U7905 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n6498), .ZN(n6299) );
  AOI21_X1 U7906 ( .B1(n6498), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6299), .ZN(
        n6300) );
  NAND2_X1 U7907 ( .A1(n6301), .A2(n6300), .ZN(n6497) );
  OAI21_X1 U7908 ( .B1(n6301), .B2(n6300), .A(n6497), .ZN(n6302) );
  AND2_X1 U7909 ( .A1(n9707), .A2(n6302), .ZN(n6305) );
  INV_X1 U7910 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10048) );
  OR2_X1 U7911 ( .A1(n8975), .A2(P1_U3084), .ZN(n8966) );
  NOR2_X1 U7912 ( .A1(n6443), .A2(n8966), .ZN(n6303) );
  INV_X1 U7913 ( .A(n6498), .ZN(n6385) );
  OAI22_X1 U7914 ( .A1(n9689), .A2(n10048), .B1(n9687), .B2(n6385), .ZN(n6304)
         );
  OR4_X1 U7915 ( .A1(n7232), .A2(n6306), .A3(n6305), .A4(n6304), .ZN(P1_U3250)
         );
  NOR2_X1 U7916 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9340), .ZN(n7032) );
  NOR2_X1 U7917 ( .A1(n6308), .A2(n6307), .ZN(n6310) );
  NOR2_X1 U7918 ( .A1(n6310), .A2(n6309), .ZN(n6311) );
  AND2_X1 U7919 ( .A1(n9697), .A2(n6311), .ZN(n6319) );
  OAI21_X1 U7920 ( .B1(n6314), .B2(n6313), .A(n6312), .ZN(n6315) );
  AND2_X1 U7921 ( .A1(n9707), .A2(n6315), .ZN(n6318) );
  INV_X1 U7922 ( .A(n6316), .ZN(n6372) );
  OAI22_X1 U7923 ( .A1(n9689), .A2(n9395), .B1(n9687), .B2(n6372), .ZN(n6317)
         );
  OR4_X1 U7924 ( .A1(n7032), .A2(n6319), .A3(n6318), .A4(n6317), .ZN(P1_U3247)
         );
  OR2_X1 U7925 ( .A1(n5639), .A2(n5638), .ZN(n6321) );
  INV_X1 U7926 ( .A(n8877), .ZN(n8837) );
  NAND2_X1 U7927 ( .A1(n4246), .A2(n8837), .ZN(n6320) );
  INV_X1 U7928 ( .A(n9743), .ZN(n6811) );
  NAND2_X2 U7929 ( .A1(n8900), .A2(n6343), .ZN(n8841) );
  NAND2_X1 U7930 ( .A1(n8725), .A2(n8841), .ZN(n6820) );
  NAND2_X1 U7931 ( .A1(n9725), .A2(n6575), .ZN(n6819) );
  INV_X2 U7932 ( .A(n6575), .ZN(n9778) );
  NAND2_X1 U7933 ( .A1(n9778), .A2(n9755), .ZN(n8842) );
  XNOR2_X1 U7934 ( .A(n6820), .B(n8726), .ZN(n6335) );
  NAND2_X1 U7935 ( .A1(n6325), .A2(n8841), .ZN(n9752) );
  NOR2_X1 U7936 ( .A1(n6324), .A2(n9743), .ZN(n9738) );
  NAND2_X1 U7937 ( .A1(n8900), .A2(n6488), .ZN(n6326) );
  NAND2_X1 U7938 ( .A1(n6328), .A2(n8726), .ZN(n6329) );
  NAND2_X1 U7939 ( .A1(n6816), .A2(n6329), .ZN(n9782) );
  NAND2_X1 U7940 ( .A1(n6340), .A2(n5638), .ZN(n6331) );
  NAND2_X1 U7941 ( .A1(n4246), .A2(n8875), .ZN(n6330) );
  MUX2_X1 U7942 ( .A(n6331), .B(n6330), .S(n5639), .Z(n9759) );
  INV_X1 U7943 ( .A(n9759), .ZN(n9270) );
  NAND2_X1 U7944 ( .A1(n9782), .A2(n9270), .ZN(n6334) );
  INV_X1 U7945 ( .A(n8899), .ZN(n6821) );
  OAI22_X1 U7946 ( .A1(n6322), .A2(n9724), .B1(n9723), .B2(n6821), .ZN(n6332)
         );
  INV_X1 U7947 ( .A(n6332), .ZN(n6333) );
  OAI211_X1 U7948 ( .C1(n9751), .C2(n6335), .A(n6334), .B(n6333), .ZN(n9780)
         );
  INV_X1 U7949 ( .A(n6337), .ZN(n6338) );
  AND2_X1 U7950 ( .A1(n6466), .A2(n9542), .ZN(n6339) );
  NAND2_X1 U7951 ( .A1(n6465), .A2(n6339), .ZN(n6844) );
  MUX2_X1 U7952 ( .A(n9780), .B(P1_REG2_REG_2__SCAN_IN), .S(n9234), .Z(n6347)
         );
  INV_X1 U7953 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6578) );
  OAI22_X1 U7954 ( .A1(n9733), .A2(n9778), .B1(n6578), .B2(n9222), .ZN(n6346)
         );
  INV_X1 U7955 ( .A(n9782), .ZN(n6344) );
  NOR2_X1 U7956 ( .A1(n6340), .A2(n5638), .ZN(n9761) );
  NAND2_X1 U7957 ( .A1(n9762), .A2(n9761), .ZN(n9276) );
  INV_X1 U7958 ( .A(n8875), .ZN(n6341) );
  NOR2_X1 U7959 ( .A1(n6469), .A2(n6341), .ZN(n6342) );
  NAND2_X1 U7960 ( .A1(n9762), .A2(n6342), .ZN(n9042) );
  NAND2_X1 U7961 ( .A1(n6343), .A2(n9743), .ZN(n9741) );
  OAI21_X1 U7962 ( .B1(n4520), .B2(n9778), .A(n9714), .ZN(n9779) );
  OAI22_X1 U7963 ( .A1(n6344), .A2(n9276), .B1(n9042), .B2(n9779), .ZN(n6345)
         );
  OR3_X1 U7964 ( .A1(n6347), .A2(n6346), .A3(n6345), .ZN(P1_U3289) );
  NAND2_X1 U7965 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_STATE_REG_SCAN_IN), .ZN(
        n6445) );
  OAI21_X1 U7966 ( .B1(n6348), .B2(P1_STATE_REG_SCAN_IN), .A(n6445), .ZN(
        P1_U3353) );
  NOR2_X1 U7967 ( .A1(n7613), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9547) );
  INV_X2 U7968 ( .A(n9547), .ZN(n7852) );
  INV_X1 U7969 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6350) );
  AND2_X1 U7970 ( .A1(n7613), .A2(P1_U3084), .ZN(n7567) );
  OAI222_X1 U7971 ( .A1(n7852), .A2(n6350), .B1(n4249), .B2(n6359), .C1(
        P1_U3084), .C2(n6349), .ZN(P1_U3351) );
  OAI222_X1 U7972 ( .A1(P1_U3084), .A2(n6351), .B1(n4249), .B2(n6354), .C1(
        n5653), .C2(n7852), .ZN(P1_U3352) );
  OAI222_X1 U7973 ( .A1(n7852), .A2(n6353), .B1(n4249), .B2(n6363), .C1(
        P1_U3084), .C2(n6352), .ZN(P1_U3350) );
  AND2_X1 U7974 ( .A1(n7613), .A2(P2_U3152), .ZN(n8461) );
  INV_X1 U7975 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6355) );
  NOR2_X1 U7976 ( .A1(n7613), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8460) );
  INV_X2 U7977 ( .A(n8460), .ZN(n8467) );
  OAI222_X1 U7978 ( .A1(n8465), .A2(n6355), .B1(n8467), .B2(n6354), .C1(n6536), 
        .C2(P2_U3152), .ZN(P2_U3357) );
  OAI222_X1 U7979 ( .A1(n7852), .A2(n6357), .B1(n4249), .B2(n6368), .C1(
        P1_U3084), .C2(n6356), .ZN(P1_U3349) );
  AOI22_X1 U7980 ( .A1(n9555), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n8461), .ZN(n6358) );
  OAI21_X1 U7981 ( .B1(n6359), .B2(n8467), .A(n6358), .ZN(P2_U3356) );
  INV_X1 U7982 ( .A(n6360), .ZN(n6366) );
  OAI222_X1 U7983 ( .A1(n7852), .A2(n6361), .B1(n4249), .B2(n6366), .C1(
        P1_U3084), .C2(n9655), .ZN(P1_U3348) );
  NAND2_X1 U7984 ( .A1(n6472), .A2(n9541), .ZN(n6362) );
  OAI21_X1 U7985 ( .B1(n9541), .B2(n6186), .A(n6362), .ZN(P1_U3440) );
  INV_X1 U7986 ( .A(n7978), .ZN(n6515) );
  OAI222_X1 U7987 ( .A1(n8465), .A2(n6364), .B1(n8467), .B2(n6363), .C1(
        P2_U3152), .C2(n6515), .ZN(P2_U3355) );
  INV_X1 U7988 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6367) );
  OAI222_X1 U7989 ( .A1(n8465), .A2(n6367), .B1(n8467), .B2(n6366), .C1(
        P2_U3152), .C2(n6365), .ZN(P2_U3353) );
  INV_X1 U7990 ( .A(n7993), .ZN(n6516) );
  OAI222_X1 U7991 ( .A1(n8465), .A2(n6369), .B1(n8467), .B2(n6368), .C1(
        P2_U3152), .C2(n6516), .ZN(P2_U3354) );
  INV_X1 U7992 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6371) );
  INV_X1 U7993 ( .A(n6370), .ZN(n6373) );
  INV_X1 U7994 ( .A(n8019), .ZN(n6519) );
  OAI222_X1 U7995 ( .A1(n8465), .A2(n6371), .B1(n8467), .B2(n6373), .C1(
        P2_U3152), .C2(n6519), .ZN(P2_U3352) );
  INV_X1 U7996 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6374) );
  OAI222_X1 U7997 ( .A1(n7852), .A2(n6374), .B1(n4249), .B2(n6373), .C1(
        P1_U3084), .C2(n6372), .ZN(P1_U3347) );
  INV_X1 U7998 ( .A(n6375), .ZN(n6378) );
  AOI22_X1 U7999 ( .A1(n6419), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9547), .ZN(n6376) );
  OAI21_X1 U8000 ( .B1(n6378), .B2(n4249), .A(n6376), .ZN(P1_U3346) );
  AOI22_X1 U8001 ( .A1(n8031), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n8461), .ZN(n6377) );
  OAI21_X1 U8002 ( .B1(n6378), .B2(n8467), .A(n6377), .ZN(P2_U3351) );
  INV_X1 U8003 ( .A(n6379), .ZN(n6382) );
  INV_X1 U8004 ( .A(n8044), .ZN(n6522) );
  OAI222_X1 U8005 ( .A1(n8465), .A2(n6380), .B1(n8467), .B2(n6382), .C1(
        P2_U3152), .C2(n6522), .ZN(P2_U3350) );
  OAI222_X1 U8006 ( .A1(n7852), .A2(n9360), .B1(n4249), .B2(n6382), .C1(
        P1_U3084), .C2(n6381), .ZN(P1_U3345) );
  INV_X1 U8007 ( .A(n6383), .ZN(n6386) );
  AOI22_X1 U8008 ( .A1(n8057), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n8461), .ZN(n6384) );
  OAI21_X1 U8009 ( .B1(n6386), .B2(n8467), .A(n6384), .ZN(P2_U3349) );
  OAI222_X1 U8010 ( .A1(n7852), .A2(n6387), .B1(n4249), .B2(n6386), .C1(n6385), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  NAND2_X1 U8011 ( .A1(n6594), .A2(P2_U3966), .ZN(n6388) );
  OAI21_X1 U8012 ( .B1(n5623), .B2(P2_U3966), .A(n6388), .ZN(P2_U3552) );
  INV_X1 U8013 ( .A(n6389), .ZN(n6402) );
  AOI22_X1 U8014 ( .A1(n6609), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n8461), .ZN(n6390) );
  OAI21_X1 U8015 ( .B1(n6402), .B2(n8467), .A(n6390), .ZN(P2_U3347) );
  INV_X1 U8016 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6391) );
  NOR2_X1 U8017 ( .A1(n4903), .A2(n6391), .ZN(n6396) );
  INV_X1 U8018 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8083) );
  NOR2_X1 U8019 ( .A1(n6392), .A2(n8083), .ZN(n6395) );
  INV_X1 U8020 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6393) );
  NOR2_X1 U8021 ( .A1(n7624), .A2(n6393), .ZN(n6394) );
  OR3_X1 U8022 ( .A1(n6396), .A2(n6395), .A3(n6394), .ZN(n8085) );
  NAND2_X1 U8023 ( .A1(n8085), .A2(P2_U3966), .ZN(n6397) );
  OAI21_X1 U8024 ( .B1(n4528), .B2(P2_U3966), .A(n6397), .ZN(P2_U3583) );
  INV_X1 U8025 ( .A(n6551), .ZN(n6682) );
  INV_X1 U8026 ( .A(n6398), .ZN(n6401) );
  OAI222_X1 U8027 ( .A1(P2_U3152), .A2(n6682), .B1(n8467), .B2(n6401), .C1(
        n6399), .C2(n8465), .ZN(P2_U3348) );
  INV_X1 U8028 ( .A(n9674), .ZN(n9686) );
  OAI222_X1 U8029 ( .A1(P1_U3084), .A2(n9686), .B1(n4249), .B2(n6401), .C1(
        n6400), .C2(n7852), .ZN(P1_U3343) );
  INV_X1 U8030 ( .A(n6934), .ZN(n6495) );
  OAI222_X1 U8031 ( .A1(n7852), .A2(n6403), .B1(n4249), .B2(n6402), .C1(n6495), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  NAND2_X1 U8032 ( .A1(n7846), .A2(n6532), .ZN(n6408) );
  OR2_X1 U8033 ( .A1(n6404), .A2(P2_U3152), .ZN(n7849) );
  NAND2_X1 U8034 ( .A1(n9882), .A2(n7849), .ZN(n6406) );
  NAND2_X1 U8035 ( .A1(n6406), .A2(n6405), .ZN(n6407) );
  AND2_X1 U8036 ( .A1(n6408), .A2(n6407), .ZN(n8082) );
  NOR2_X1 U8037 ( .A1(n9850), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8038 ( .A(n6409), .ZN(n6425) );
  AOI22_X1 U8039 ( .A1(n8934), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9547), .ZN(n6410) );
  OAI21_X1 U8040 ( .B1(n6425), .B2(n4249), .A(n6410), .ZN(P1_U3341) );
  INV_X1 U8041 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6422) );
  OAI21_X1 U8042 ( .B1(n6413), .B2(n6412), .A(n6411), .ZN(n6418) );
  OAI21_X1 U8043 ( .B1(n6416), .B2(n6415), .A(n6414), .ZN(n6417) );
  AOI22_X1 U8044 ( .A1(n9697), .A2(n6418), .B1(n9707), .B2(n6417), .ZN(n6421)
         );
  AND2_X1 U8045 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6989) );
  AOI21_X1 U8046 ( .B1(n9699), .B2(n6419), .A(n6989), .ZN(n6420) );
  OAI211_X1 U8047 ( .C1(n9689), .C2(n6422), .A(n6421), .B(n6420), .ZN(P1_U3248) );
  INV_X1 U8048 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6424) );
  NAND2_X1 U8049 ( .A1(n6323), .A2(P1_U4006), .ZN(n6423) );
  OAI21_X1 U8050 ( .B1(P1_U4006), .B2(n6424), .A(n6423), .ZN(P1_U3555) );
  INV_X1 U8051 ( .A(n6554), .ZN(n6675) );
  OAI222_X1 U8052 ( .A1(n8465), .A2(n6426), .B1(n8467), .B2(n6425), .C1(
        P2_U3152), .C2(n6675), .ZN(P2_U3346) );
  INV_X1 U8053 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6431) );
  NAND2_X1 U8054 ( .A1(n5686), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6429) );
  NAND2_X1 U8055 ( .A1(n8599), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U8056 ( .A1(n8600), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6427) );
  INV_X1 U8057 ( .A(n8977), .ZN(n8717) );
  NAND2_X1 U8058 ( .A1(n8717), .A2(P1_U4006), .ZN(n6430) );
  OAI21_X1 U8059 ( .B1(P1_U4006), .B2(n6431), .A(n6430), .ZN(P1_U3586) );
  INV_X1 U8060 ( .A(n7266), .ZN(n6433) );
  INV_X1 U8061 ( .A(n6432), .ZN(n6434) );
  OAI222_X1 U8062 ( .A1(P1_U3084), .A2(n6433), .B1(n4249), .B2(n6434), .C1(
        n9427), .C2(n7852), .ZN(P1_U3340) );
  INV_X1 U8063 ( .A(n6658), .ZN(n6653) );
  OAI222_X1 U8064 ( .A1(n8465), .A2(n6435), .B1(n8467), .B2(n6434), .C1(n6653), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8065 ( .A(n6436), .ZN(n6438) );
  INV_X1 U8066 ( .A(n7507), .ZN(n7498) );
  OAI222_X1 U8067 ( .A1(n7852), .A2(n6437), .B1(n4249), .B2(n6438), .C1(n7498), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8068 ( .A(n6659), .ZN(n6699) );
  OAI222_X1 U8069 ( .A1(n8465), .A2(n6439), .B1(n8467), .B2(n6438), .C1(n6699), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8070 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6463) );
  OAI21_X1 U8071 ( .B1(n6440), .B2(n6442), .A(n6441), .ZN(n6480) );
  NAND2_X1 U8072 ( .A1(n6443), .A2(n8975), .ZN(n9619) );
  NOR2_X1 U8073 ( .A1(n6480), .A2(n9619), .ZN(n6450) );
  NOR2_X1 U8074 ( .A1(n8975), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6444) );
  OR2_X1 U8075 ( .A1(n7569), .A2(n6444), .ZN(n6446) );
  AND2_X1 U8076 ( .A1(n6446), .A2(n6445), .ZN(n9617) );
  OR2_X1 U8077 ( .A1(n6209), .A2(n8975), .ZN(n8755) );
  NOR2_X1 U8078 ( .A1(n8755), .A2(n6447), .ZN(n9621) );
  INV_X1 U8079 ( .A(n6448), .ZN(n6449) );
  NOR4_X1 U8080 ( .A1(n6450), .A2(n9617), .A3(n9621), .A4(n6449), .ZN(n9638)
         );
  INV_X1 U8081 ( .A(n9638), .ZN(n6462) );
  AOI22_X1 U8082 ( .A1(n9699), .A2(n6451), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        P1_U3084), .ZN(n6460) );
  OAI211_X1 U8083 ( .C1(n6454), .C2(n6453), .A(n9697), .B(n6452), .ZN(n6459)
         );
  OAI211_X1 U8084 ( .C1(n6457), .C2(n6456), .A(n9707), .B(n6455), .ZN(n6458)
         );
  AND3_X1 U8085 ( .A1(n6460), .A2(n6459), .A3(n6458), .ZN(n6461) );
  OAI211_X1 U8086 ( .C1(n6463), .C2(n9689), .A(n6462), .B(n6461), .ZN(P1_U3243) );
  AOI21_X1 U8087 ( .B1(n9742), .B2(n9744), .A(n9542), .ZN(n6464) );
  INV_X1 U8088 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6471) );
  OR2_X1 U8089 ( .A1(n6324), .A2(n6811), .ZN(n8844) );
  INV_X1 U8090 ( .A(n8757), .ZN(n6856) );
  AOI211_X1 U8091 ( .C1(n9749), .C2(n8844), .A(n6467), .B(n6856), .ZN(n6468)
         );
  AOI21_X1 U8092 ( .B1(n9756), .B2(n8900), .A(n6468), .ZN(n6808) );
  OAI21_X1 U8093 ( .B1(n9743), .B2(n6469), .A(n6808), .ZN(n6474) );
  NAND2_X1 U8094 ( .A1(n6474), .A2(n9828), .ZN(n6470) );
  OAI21_X1 U8095 ( .B1(n9828), .B2(n6471), .A(n6470), .ZN(P1_U3454) );
  INV_X1 U8096 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9624) );
  NAND2_X1 U8097 ( .A1(n6474), .A2(n9843), .ZN(n6475) );
  OAI21_X1 U8098 ( .B1(n9843), .B2(n9624), .A(n6475), .ZN(P1_U3523) );
  INV_X1 U8099 ( .A(n6476), .ZN(n6479) );
  AND3_X1 U8100 ( .A1(n6479), .A2(n6478), .A3(n6477), .ZN(n6579) );
  INV_X1 U8101 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6809) );
  AOI22_X1 U8102 ( .A1(n8590), .A2(n6811), .B1(n8552), .B2(n8900), .ZN(n6482)
         );
  NAND2_X1 U8103 ( .A1(n6480), .A2(n8571), .ZN(n6481) );
  OAI211_X1 U8104 ( .C1(n6579), .C2(n6809), .A(n6482), .B(n6481), .ZN(P1_U3230) );
  INV_X1 U8105 ( .A(n6484), .ZN(n6571) );
  AOI21_X1 U8106 ( .B1(n6485), .B2(n6483), .A(n6571), .ZN(n6490) );
  INV_X1 U8107 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n8901) );
  NOR2_X1 U8108 ( .A1(n6579), .A2(n8901), .ZN(n6487) );
  OAI22_X1 U8109 ( .A1(n6324), .A2(n8573), .B1(n8588), .B2(n9725), .ZN(n6486)
         );
  AOI211_X1 U8110 ( .C1(n6488), .C2(n8590), .A(n6487), .B(n6486), .ZN(n6489)
         );
  OAI21_X1 U8111 ( .B1(n6490), .B2(n8592), .A(n6489), .ZN(P1_U3220) );
  INV_X1 U8112 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6506) );
  XNOR2_X1 U8113 ( .A(n9674), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n9681) );
  NOR2_X1 U8114 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6934), .ZN(n6492) );
  AOI21_X1 U8115 ( .B1(n6934), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6492), .ZN(
        n6493) );
  OAI21_X1 U8116 ( .B1(n6494), .B2(n6493), .A(n6935), .ZN(n6503) );
  INV_X1 U8117 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9608) );
  AOI22_X1 U8118 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n6934), .B1(n6495), .B2(
        n9608), .ZN(n6501) );
  INV_X1 U8119 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6496) );
  MUX2_X1 U8120 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6496), .S(n9674), .Z(n6499)
         );
  OAI21_X1 U8121 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n6498), .A(n6497), .ZN(
        n9677) );
  NAND2_X1 U8122 ( .A1(n6499), .A2(n9677), .ZN(n9676) );
  OAI21_X1 U8123 ( .B1(n9674), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9676), .ZN(
        n6500) );
  NAND2_X1 U8124 ( .A1(n6501), .A2(n6500), .ZN(n6928) );
  OAI21_X1 U8125 ( .B1(n6501), .B2(n6500), .A(n6928), .ZN(n6502) );
  AOI22_X1 U8126 ( .A1(n6503), .A2(n9697), .B1(n9707), .B2(n6502), .ZN(n6505)
         );
  AND2_X1 U8127 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7381) );
  AOI21_X1 U8128 ( .B1(n9699), .B2(n6934), .A(n7381), .ZN(n6504) );
  OAI211_X1 U8129 ( .C1(n9689), .C2(n6506), .A(n6505), .B(n6504), .ZN(P1_U3252) );
  INV_X1 U8130 ( .A(n6507), .ZN(n6509) );
  OAI222_X1 U8131 ( .A1(n7852), .A2(n6508), .B1(n4249), .B2(n6509), .C1(
        P1_U3084), .C2(n7550), .ZN(P1_U3338) );
  INV_X1 U8132 ( .A(n6799), .ZN(n6789) );
  OAI222_X1 U8133 ( .A1(n8465), .A2(n9428), .B1(n8467), .B2(n6509), .C1(
        P2_U3152), .C2(n6789), .ZN(P2_U3343) );
  NOR2_X1 U8134 ( .A1(n6609), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6525) );
  NAND2_X1 U8135 ( .A1(n8057), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6523) );
  MUX2_X1 U8136 ( .A(n7210), .B(P2_REG2_REG_9__SCAN_IN), .S(n8057), .Z(n6510)
         );
  INV_X1 U8137 ( .A(n6510), .ZN(n8054) );
  NAND2_X1 U8138 ( .A1(n8031), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6521) );
  MUX2_X1 U8139 ( .A(n6951), .B(P2_REG2_REG_7__SCAN_IN), .S(n8031), .Z(n6511)
         );
  INV_X1 U8140 ( .A(n6511), .ZN(n8029) );
  NAND2_X1 U8141 ( .A1(n8006), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6518) );
  MUX2_X1 U8142 ( .A(n6733), .B(P2_REG2_REG_5__SCAN_IN), .S(n8006), .Z(n6512)
         );
  INV_X1 U8143 ( .A(n6512), .ZN(n8003) );
  MUX2_X1 U8144 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6513), .S(n9555), .Z(n9558)
         );
  INV_X1 U8145 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6925) );
  XNOR2_X1 U8146 ( .A(n6536), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n7964) );
  NAND3_X1 U8147 ( .A1(n7964), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_REG2_REG_0__SCAN_IN), .ZN(n7962) );
  OAI21_X1 U8148 ( .B1(n6925), .B2(n6536), .A(n7962), .ZN(n9559) );
  NAND2_X1 U8149 ( .A1(n9558), .A2(n9559), .ZN(n9557) );
  NAND2_X1 U8150 ( .A1(n9555), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7974) );
  MUX2_X1 U8151 ( .A(n6514), .B(P2_REG2_REG_3__SCAN_IN), .S(n7978), .Z(n7973)
         );
  AOI21_X1 U8152 ( .B1(n9557), .B2(n7974), .A(n7973), .ZN(n7987) );
  NOR2_X1 U8153 ( .A1(n6515), .A2(n6514), .ZN(n7986) );
  MUX2_X1 U8154 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6517), .S(n7993), .Z(n7988)
         );
  OAI21_X1 U8155 ( .B1(n7987), .B2(n7986), .A(n7988), .ZN(n7990) );
  OAI21_X1 U8156 ( .B1(n6517), .B2(n6516), .A(n7990), .ZN(n8002) );
  NAND2_X1 U8157 ( .A1(n8003), .A2(n8002), .ZN(n8001) );
  NAND2_X1 U8158 ( .A1(n6518), .A2(n8001), .ZN(n8016) );
  MUX2_X1 U8159 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6520), .S(n8019), .Z(n8015)
         );
  NAND2_X1 U8160 ( .A1(n8016), .A2(n8015), .ZN(n8014) );
  OAI21_X1 U8161 ( .B1(n6520), .B2(n6519), .A(n8014), .ZN(n8028) );
  NAND2_X1 U8162 ( .A1(n8029), .A2(n8028), .ZN(n8027) );
  NAND2_X1 U8163 ( .A1(n6521), .A2(n8027), .ZN(n8041) );
  MUX2_X1 U8164 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6975), .S(n8044), .Z(n8040)
         );
  NAND2_X1 U8165 ( .A1(n8041), .A2(n8040), .ZN(n8039) );
  OAI21_X1 U8166 ( .B1(n6975), .B2(n6522), .A(n8039), .ZN(n8053) );
  NAND2_X1 U8167 ( .A1(n8054), .A2(n8053), .ZN(n8052) );
  NAND2_X1 U8168 ( .A1(n6523), .A2(n8052), .ZN(n6687) );
  MUX2_X1 U8169 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7170), .S(n6551), .Z(n6686)
         );
  NAND2_X1 U8170 ( .A1(n6687), .A2(n6686), .ZN(n6685) );
  OAI21_X1 U8171 ( .B1(n7170), .B2(n6682), .A(n6685), .ZN(n6607) );
  MUX2_X1 U8172 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n7352), .S(n6609), .Z(n6524)
         );
  INV_X1 U8173 ( .A(n6524), .ZN(n6606) );
  NOR2_X1 U8174 ( .A1(n6607), .A2(n6606), .ZN(n6605) );
  NOR2_X1 U8175 ( .A1(n6525), .A2(n6605), .ZN(n6672) );
  MUX2_X1 U8176 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n6526), .S(n6554), .Z(n6671)
         );
  NAND2_X1 U8177 ( .A1(n6672), .A2(n6671), .ZN(n6670) );
  OAI21_X1 U8178 ( .B1(n6526), .B2(n6675), .A(n6670), .ZN(n6529) );
  MUX2_X1 U8179 ( .A(n6527), .B(P2_REG2_REG_13__SCAN_IN), .S(n6658), .Z(n6528)
         );
  NOR2_X1 U8180 ( .A1(n6529), .A2(n6528), .ZN(n6652) );
  AOI21_X1 U8181 ( .B1(n6529), .B2(n6528), .A(n6652), .ZN(n6567) );
  NOR2_X1 U8182 ( .A1(n6560), .A2(P2_U3152), .ZN(n7564) );
  INV_X1 U8183 ( .A(n7849), .ZN(n7224) );
  AOI21_X1 U8184 ( .B1(n6530), .B2(n7564), .A(n7224), .ZN(n6531) );
  OAI21_X1 U8185 ( .B1(n9882), .B2(n6532), .A(n6531), .ZN(n6558) );
  NAND2_X1 U8186 ( .A1(n6533), .A2(n7961), .ZN(n6561) );
  NOR2_X1 U8187 ( .A1(n6560), .A2(n7844), .ZN(n6534) );
  NAND2_X1 U8188 ( .A1(n6561), .A2(n6534), .ZN(n9848) );
  MUX2_X1 U8189 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n6535), .S(n6658), .Z(n6556)
         );
  MUX2_X1 U8190 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n4885), .S(n9555), .Z(n9552)
         );
  MUX2_X1 U8191 ( .A(n4830), .B(P2_REG1_REG_1__SCAN_IN), .S(n6536), .Z(n7968)
         );
  AND2_X1 U8192 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n7967) );
  NAND2_X1 U8193 ( .A1(n7968), .A2(n7967), .ZN(n7966) );
  NAND2_X1 U8194 ( .A1(n7965), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U8195 ( .A1(n7966), .A2(n6537), .ZN(n9551) );
  NAND2_X1 U8196 ( .A1(n9552), .A2(n9551), .ZN(n9550) );
  NAND2_X1 U8197 ( .A1(n9555), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6538) );
  NAND2_X1 U8198 ( .A1(n9550), .A2(n6538), .ZN(n7980) );
  INV_X1 U8199 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6539) );
  XNOR2_X1 U8200 ( .A(n7978), .B(n6539), .ZN(n7981) );
  NAND2_X1 U8201 ( .A1(n7980), .A2(n7981), .ZN(n7979) );
  NAND2_X1 U8202 ( .A1(n7978), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6540) );
  NAND2_X1 U8203 ( .A1(n7979), .A2(n6540), .ZN(n7995) );
  INV_X1 U8204 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6541) );
  XNOR2_X1 U8205 ( .A(n7993), .B(n6541), .ZN(n7996) );
  NAND2_X1 U8206 ( .A1(n7995), .A2(n7996), .ZN(n7994) );
  NAND2_X1 U8207 ( .A1(n7993), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U8208 ( .A1(n7994), .A2(n6542), .ZN(n8008) );
  OR2_X1 U8209 ( .A1(n8006), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6543) );
  NAND2_X1 U8210 ( .A1(n8006), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6544) );
  AND2_X1 U8211 ( .A1(n6543), .A2(n6544), .ZN(n8009) );
  NAND2_X1 U8212 ( .A1(n8008), .A2(n8009), .ZN(n8007) );
  NAND2_X1 U8213 ( .A1(n8007), .A2(n6544), .ZN(n8021) );
  INV_X1 U8214 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6545) );
  XNOR2_X1 U8215 ( .A(n8019), .B(n6545), .ZN(n8022) );
  NAND2_X1 U8216 ( .A1(n8021), .A2(n8022), .ZN(n8020) );
  NAND2_X1 U8217 ( .A1(n8019), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U8218 ( .A1(n8020), .A2(n6546), .ZN(n8033) );
  INV_X1 U8219 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9437) );
  MUX2_X1 U8220 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9437), .S(n8031), .Z(n8034)
         );
  NAND2_X1 U8221 ( .A1(n8033), .A2(n8034), .ZN(n8032) );
  NAND2_X1 U8222 ( .A1(n8031), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6547) );
  NAND2_X1 U8223 ( .A1(n8032), .A2(n6547), .ZN(n8046) );
  INV_X1 U8224 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10003) );
  MUX2_X1 U8225 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10003), .S(n8044), .Z(n8047)
         );
  NAND2_X1 U8226 ( .A1(n8046), .A2(n8047), .ZN(n8045) );
  NAND2_X1 U8227 ( .A1(n8044), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6548) );
  NAND2_X1 U8228 ( .A1(n8045), .A2(n6548), .ZN(n8059) );
  INV_X1 U8229 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6549) );
  MUX2_X1 U8230 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6549), .S(n8057), .Z(n8060)
         );
  NAND2_X1 U8231 ( .A1(n8059), .A2(n8060), .ZN(n8058) );
  NAND2_X1 U8232 ( .A1(n8057), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U8233 ( .A1(n8058), .A2(n6550), .ZN(n6679) );
  MUX2_X1 U8234 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n5075), .S(n6551), .Z(n6680)
         );
  AND2_X1 U8235 ( .A1(n6679), .A2(n6680), .ZN(n6691) );
  AOI21_X1 U8236 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n6551), .A(n6691), .ZN(
        n6604) );
  MUX2_X1 U8237 ( .A(n6552), .B(P2_REG1_REG_11__SCAN_IN), .S(n6609), .Z(n6603)
         );
  NOR2_X1 U8238 ( .A1(n6604), .A2(n6603), .ZN(n6602) );
  AOI21_X1 U8239 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n6609), .A(n6602), .ZN(
        n6669) );
  MUX2_X1 U8240 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6553), .S(n6554), .Z(n6668)
         );
  NAND2_X1 U8241 ( .A1(n6669), .A2(n6668), .ZN(n6667) );
  OAI21_X1 U8242 ( .B1(n6554), .B2(P2_REG1_REG_12__SCAN_IN), .A(n6667), .ZN(
        n6555) );
  NAND2_X1 U8243 ( .A1(n6555), .A2(n6556), .ZN(n6657) );
  OAI21_X1 U8244 ( .B1(n6556), .B2(n6555), .A(n6657), .ZN(n6559) );
  NAND2_X1 U8245 ( .A1(n6559), .A2(n9845), .ZN(n6566) );
  INV_X1 U8246 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6563) );
  AND2_X1 U8247 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7249) );
  INV_X1 U8248 ( .A(n7249), .ZN(n6562) );
  OAI21_X1 U8249 ( .B1(n8082), .B2(n6563), .A(n6562), .ZN(n6564) );
  AOI21_X1 U8250 ( .B1(n9556), .B2(n6658), .A(n6564), .ZN(n6565) );
  OAI211_X1 U8251 ( .C1(n6567), .C2(n9848), .A(n6566), .B(n6565), .ZN(P2_U3258) );
  INV_X1 U8252 ( .A(n6568), .ZN(n6570) );
  NOR3_X1 U8253 ( .A1(n6571), .A2(n6570), .A3(n6569), .ZN(n6573) );
  INV_X1 U8254 ( .A(n6572), .ZN(n6626) );
  OAI21_X1 U8255 ( .B1(n6573), .B2(n6626), .A(n8571), .ZN(n6577) );
  OAI22_X1 U8256 ( .A1(n6322), .A2(n8573), .B1(n8588), .B2(n6821), .ZN(n6574)
         );
  AOI21_X1 U8257 ( .B1(n6575), .B2(n8590), .A(n6574), .ZN(n6576) );
  OAI211_X1 U8258 ( .C1(n6579), .C2(n6578), .A(n6577), .B(n6576), .ZN(P1_U3235) );
  INV_X1 U8259 ( .A(n6580), .ZN(n6581) );
  AOI21_X1 U8260 ( .B1(n6583), .B2(n6582), .A(n6581), .ZN(n6588) );
  INV_X1 U8261 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6921) );
  OR2_X1 U8262 ( .A1(n6585), .A2(P2_U3152), .ZN(n6619) );
  AOI22_X1 U8263 ( .A1(n7929), .A2(n6584), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n6619), .ZN(n6587) );
  OAI22_X1 U8264 ( .A1(n6593), .A2(n9863), .B1(n6708), .B2(n9861), .ZN(n6919)
         );
  NAND2_X1 U8265 ( .A1(n7890), .A2(n6919), .ZN(n6586) );
  OAI211_X1 U8266 ( .C1(n6588), .C2(n7931), .A(n6587), .B(n6586), .ZN(P2_U3224) );
  INV_X1 U8267 ( .A(n6589), .ZN(n6591) );
  INV_X1 U8268 ( .A(n8944), .ZN(n7557) );
  OAI222_X1 U8269 ( .A1(n7852), .A2(n6590), .B1(n4249), .B2(n6591), .C1(n7557), 
        .C2(P1_U3084), .ZN(P1_U3337) );
  INV_X1 U8270 ( .A(n7089), .ZN(n6803) );
  OAI222_X1 U8271 ( .A1(n8465), .A2(n6592), .B1(n8467), .B2(n6591), .C1(n6803), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  INV_X1 U8272 ( .A(n6619), .ZN(n6601) );
  INV_X1 U8273 ( .A(n7939), .ZN(n6618) );
  AOI22_X1 U8274 ( .A1(n6618), .A2(n6704), .B1(n6917), .B2(n7929), .ZN(n6599)
         );
  INV_X1 U8275 ( .A(n6918), .ZN(n6597) );
  INV_X1 U8276 ( .A(n6917), .ZN(n9921) );
  NAND2_X1 U8277 ( .A1(n6594), .A2(n9921), .ZN(n7651) );
  INV_X1 U8278 ( .A(n7651), .ZN(n6595) );
  MUX2_X1 U8279 ( .A(n6917), .B(n6595), .S(n4250), .Z(n6596) );
  OAI21_X1 U8280 ( .B1(n6597), .B2(n6596), .A(n7933), .ZN(n6598) );
  OAI211_X1 U8281 ( .C1(n6601), .C2(n6600), .A(n6599), .B(n6598), .ZN(P2_U3234) );
  INV_X1 U8282 ( .A(n9845), .ZN(n7283) );
  AOI211_X1 U8283 ( .C1(n6604), .C2(n6603), .A(n7283), .B(n6602), .ZN(n6614)
         );
  AOI21_X1 U8284 ( .B1(n6607), .B2(n6606), .A(n6605), .ZN(n6612) );
  NOR2_X1 U8285 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5094), .ZN(n6608) );
  AOI21_X1 U8286 ( .B1(n9850), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6608), .ZN(
        n6611) );
  NAND2_X1 U8287 ( .A1(n9556), .A2(n6609), .ZN(n6610) );
  OAI211_X1 U8288 ( .C1(n6612), .C2(n9848), .A(n6611), .B(n6610), .ZN(n6613)
         );
  OR2_X1 U8289 ( .A1(n6614), .A2(n6613), .ZN(P2_U3256) );
  NAND2_X1 U8290 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n7961), .ZN(n6615) );
  OAI21_X1 U8291 ( .B1(n8134), .B2(n7961), .A(n6615), .ZN(P2_U3581) );
  XNOR2_X1 U8292 ( .A(n6616), .B(n6617), .ZN(n6622) );
  INV_X1 U8293 ( .A(n7938), .ZN(n6775) );
  AOI22_X1 U8294 ( .A1(n6618), .A2(n7960), .B1(n6775), .B2(n6704), .ZN(n6621)
         );
  AOI22_X1 U8295 ( .A1(n7929), .A2(n8323), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n6619), .ZN(n6620) );
  OAI211_X1 U8296 ( .C1(n6622), .C2(n7931), .A(n6621), .B(n6620), .ZN(P2_U3239) );
  INV_X1 U8297 ( .A(n6623), .ZN(n6625) );
  NOR3_X1 U8298 ( .A1(n6626), .A2(n6625), .A3(n6624), .ZN(n6629) );
  INV_X1 U8299 ( .A(n6627), .ZN(n6628) );
  OAI21_X1 U8300 ( .B1(n6629), .B2(n6628), .A(n8571), .ZN(n6633) );
  AND2_X1 U8301 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8913) );
  AOI21_X1 U8302 ( .B1(n8585), .B2(n9755), .A(n8913), .ZN(n6630) );
  OAI21_X1 U8303 ( .B1(n8588), .B2(n9722), .A(n6630), .ZN(n6631) );
  AOI21_X1 U8304 ( .B1(n9713), .B2(n8590), .A(n6631), .ZN(n6632) );
  OAI211_X1 U8305 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8563), .A(n6633), .B(
        n6632), .ZN(P1_U3216) );
  INV_X1 U8306 ( .A(n6634), .ZN(n6635) );
  INV_X1 U8307 ( .A(n8962), .ZN(n8952) );
  OAI222_X1 U8308 ( .A1(n7852), .A2(n9429), .B1(n4249), .B2(n6635), .C1(n8952), 
        .C2(P1_U3084), .ZN(P1_U3336) );
  INV_X1 U8309 ( .A(n7280), .ZN(n7095) );
  OAI222_X1 U8310 ( .A1(n8465), .A2(n6636), .B1(n8467), .B2(n6635), .C1(n7095), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  XNOR2_X1 U8311 ( .A(n6638), .B(n6637), .ZN(n6642) );
  OAI22_X1 U8312 ( .A1(n9862), .A2(n9863), .B1(n6949), .B2(n9861), .ZN(n6731)
         );
  AOI22_X1 U8313 ( .A1(n7890), .A2(n6731), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n6641) );
  INV_X1 U8314 ( .A(n7925), .ZN(n7942) );
  INV_X1 U8315 ( .A(n6725), .ZN(n6639) );
  AOI22_X1 U8316 ( .A1(n9953), .A2(n7929), .B1(n7942), .B2(n6639), .ZN(n6640)
         );
  OAI211_X1 U8317 ( .C1(n6642), .C2(n7931), .A(n6641), .B(n6640), .ZN(P2_U3229) );
  INV_X1 U8318 ( .A(n6643), .ZN(n6825) );
  OAI21_X1 U8319 ( .B1(n6646), .B2(n6645), .A(n6644), .ZN(n6647) );
  NAND2_X1 U8320 ( .A1(n6647), .A2(n8571), .ZN(n6651) );
  AND2_X1 U8321 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9639) );
  AOI21_X1 U8322 ( .B1(n8552), .B2(n8897), .A(n9639), .ZN(n6648) );
  OAI21_X1 U8323 ( .B1(n8573), .B2(n6821), .A(n6648), .ZN(n6649) );
  AOI21_X1 U8324 ( .B1(n6830), .B2(n8590), .A(n6649), .ZN(n6650) );
  OAI211_X1 U8325 ( .C1(n8563), .C2(n6825), .A(n6651), .B(n6650), .ZN(P1_U3228) );
  NOR2_X1 U8326 ( .A1(n6659), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6654) );
  AOI22_X1 U8327 ( .A1(n6659), .A2(n7471), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n6699), .ZN(n6693) );
  NOR2_X1 U8328 ( .A1(n6694), .A2(n6693), .ZN(n6692) );
  NOR2_X1 U8329 ( .A1(n6654), .A2(n6692), .ZN(n6798) );
  XNOR2_X1 U8330 ( .A(n6798), .B(n6799), .ZN(n6655) );
  NOR2_X1 U8331 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n6655), .ZN(n6800) );
  AOI21_X1 U8332 ( .B1(n6655), .B2(P2_REG2_REG_15__SCAN_IN), .A(n6800), .ZN(
        n6666) );
  AND2_X1 U8333 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7519) );
  NOR2_X1 U8334 ( .A1(n9847), .A2(n6789), .ZN(n6656) );
  AOI211_X1 U8335 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n9850), .A(n7519), .B(
        n6656), .ZN(n6665) );
  INV_X1 U8336 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9578) );
  AOI22_X1 U8337 ( .A1(n6659), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n9578), .B2(
        n6699), .ZN(n6697) );
  OAI21_X1 U8338 ( .B1(n6658), .B2(P2_REG1_REG_13__SCAN_IN), .A(n6657), .ZN(
        n6696) );
  NAND2_X1 U8339 ( .A1(n6697), .A2(n6696), .ZN(n6695) );
  OAI21_X1 U8340 ( .B1(n6659), .B2(P2_REG1_REG_14__SCAN_IN), .A(n6695), .ZN(
        n6788) );
  XNOR2_X1 U8341 ( .A(n6788), .B(n6789), .ZN(n6660) );
  INV_X1 U8342 ( .A(n6660), .ZN(n6663) );
  NOR2_X1 U8343 ( .A1(n6661), .A2(n6660), .ZN(n6790) );
  INV_X1 U8344 ( .A(n6790), .ZN(n6662) );
  OAI211_X1 U8345 ( .C1(n6663), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9845), .B(
        n6662), .ZN(n6664) );
  OAI211_X1 U8346 ( .C1(n6666), .C2(n9848), .A(n6665), .B(n6664), .ZN(P2_U3260) );
  OAI21_X1 U8347 ( .B1(n6669), .B2(n6668), .A(n6667), .ZN(n6677) );
  OAI211_X1 U8348 ( .C1(n6672), .C2(n6671), .A(n6670), .B(n9844), .ZN(n6674)
         );
  AND2_X1 U8349 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7221) );
  AOI21_X1 U8350 ( .B1(n9850), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7221), .ZN(
        n6673) );
  OAI211_X1 U8351 ( .C1(n9847), .C2(n6675), .A(n6674), .B(n6673), .ZN(n6676)
         );
  AOI21_X1 U8352 ( .B1(n9845), .B2(n6677), .A(n6676), .ZN(n6678) );
  INV_X1 U8353 ( .A(n6678), .ZN(P2_U3257) );
  OAI21_X1 U8354 ( .B1(n6680), .B2(n6679), .A(n9845), .ZN(n6690) );
  NOR2_X1 U8355 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6681), .ZN(n6684) );
  NOR2_X1 U8356 ( .A1(n9847), .A2(n6682), .ZN(n6683) );
  AOI211_X1 U8357 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n9850), .A(n6684), .B(
        n6683), .ZN(n6689) );
  OAI211_X1 U8358 ( .C1(n6687), .C2(n6686), .A(n9844), .B(n6685), .ZN(n6688)
         );
  OAI211_X1 U8359 ( .C1(n6691), .C2(n6690), .A(n6689), .B(n6688), .ZN(P2_U3255) );
  AOI21_X1 U8360 ( .B1(n6694), .B2(n6693), .A(n6692), .ZN(n6703) );
  OAI21_X1 U8361 ( .B1(n6697), .B2(n6696), .A(n6695), .ZN(n6701) );
  NAND2_X1 U8362 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7442) );
  NAND2_X1 U8363 ( .A1(n9850), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n6698) );
  OAI211_X1 U8364 ( .C1(n9847), .C2(n6699), .A(n7442), .B(n6698), .ZN(n6700)
         );
  AOI21_X1 U8365 ( .B1(n6701), .B2(n9845), .A(n6700), .ZN(n6702) );
  OAI21_X1 U8366 ( .B1(n6703), .B2(n9848), .A(n6702), .ZN(P2_U3259) );
  NAND2_X1 U8367 ( .A1(n7958), .A2(n6909), .ZN(n7632) );
  NAND2_X1 U8368 ( .A1(n6705), .A2(n6584), .ZN(n7654) );
  NAND2_X1 U8369 ( .A1(n6727), .A2(n7654), .ZN(n6915) );
  NAND2_X1 U8370 ( .A1(n6915), .A2(n6916), .ZN(n6707) );
  NAND2_X1 U8371 ( .A1(n6705), .A2(n9929), .ZN(n6706) );
  NAND2_X1 U8372 ( .A1(n6707), .A2(n6706), .ZN(n8322) );
  NAND2_X1 U8373 ( .A1(n6708), .A2(n8323), .ZN(n7653) );
  NAND2_X1 U8374 ( .A1(n8322), .A2(n8329), .ZN(n6710) );
  NAND2_X1 U8375 ( .A1(n6708), .A2(n9937), .ZN(n6709) );
  NAND2_X1 U8376 ( .A1(n6710), .A2(n6709), .ZN(n9855) );
  NAND2_X1 U8377 ( .A1(n8333), .A2(n9873), .ZN(n7639) );
  NAND2_X1 U8378 ( .A1(n8333), .A2(n9872), .ZN(n6711) );
  NAND2_X1 U8379 ( .A1(n9862), .A2(n9945), .ZN(n7640) );
  INV_X1 U8380 ( .A(n9862), .ZN(n7959) );
  NAND2_X1 U8381 ( .A1(n7959), .A2(n6759), .ZN(n6898) );
  NAND2_X1 U8382 ( .A1(n7640), .A2(n6898), .ZN(n6745) );
  NAND2_X1 U8383 ( .A1(n9862), .A2(n6759), .ZN(n6712) );
  XOR2_X1 U8384 ( .A(n7772), .B(n6911), .Z(n9958) );
  INV_X1 U8385 ( .A(n7060), .ZN(n6715) );
  NOR2_X1 U8386 ( .A1(n7063), .A2(n6715), .ZN(n6716) );
  NAND2_X1 U8387 ( .A1(n7051), .A2(n6717), .ZN(n6721) );
  XNOR2_X1 U8388 ( .A(n5533), .B(n6719), .ZN(n6718) );
  NAND2_X1 U8389 ( .A1(n6718), .A2(n7839), .ZN(n9854) );
  OR2_X1 U8390 ( .A1(n6719), .A2(n7839), .ZN(n6966) );
  NAND2_X1 U8391 ( .A1(n9854), .A2(n6966), .ZN(n6720) );
  INV_X1 U8392 ( .A(n6721), .ZN(n6722) );
  NAND2_X1 U8393 ( .A1(n6722), .A2(n7839), .ZN(n8195) );
  INV_X1 U8394 ( .A(n8195), .ZN(n8328) );
  AOI211_X1 U8395 ( .C1(n9953), .C2(n6723), .A(n9985), .B(n6905), .ZN(n9952)
         );
  OAI22_X1 U8396 ( .A1(n8307), .A2(n6909), .B1(n8272), .B2(n6725), .ZN(n6726)
         );
  AOI21_X1 U8397 ( .B1(n8328), .B2(n9952), .A(n6726), .ZN(n6735) );
  NAND2_X1 U8398 ( .A1(n7645), .A2(n6727), .ZN(n8330) );
  NAND2_X1 U8399 ( .A1(n4255), .A2(n6898), .ZN(n6730) );
  XNOR2_X1 U8400 ( .A(n6730), .B(n7772), .ZN(n6732) );
  NAND2_X1 U8401 ( .A1(n7798), .A2(n7799), .ZN(n7841) );
  AOI21_X1 U8402 ( .B1(n6732), .B2(n9865), .A(n6731), .ZN(n9956) );
  MUX2_X1 U8403 ( .A(n9956), .B(n6733), .S(n4247), .Z(n6734) );
  OAI211_X1 U8404 ( .C1(n9958), .C2(n8321), .A(n6735), .B(n6734), .ZN(P2_U3291) );
  INV_X1 U8405 ( .A(n6736), .ZN(n6737) );
  AOI21_X1 U8406 ( .B1(n6739), .B2(n6738), .A(n6737), .ZN(n6743) );
  NAND2_X1 U8407 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8017) );
  OAI21_X1 U8408 ( .B1(n7925), .B2(n6904), .A(n8017), .ZN(n6741) );
  INV_X1 U8409 ( .A(n6944), .ZN(n9960) );
  OAI22_X1 U8410 ( .A1(n9960), .A2(n7945), .B1(n7939), .B2(n6970), .ZN(n6740)
         );
  AOI211_X1 U8411 ( .C1(n6775), .C2(n7958), .A(n6741), .B(n6740), .ZN(n6742)
         );
  OAI21_X1 U8412 ( .B1(n6743), .B2(n7931), .A(n6742), .ZN(P2_U3241) );
  INV_X1 U8413 ( .A(n6745), .ZN(n7770) );
  XNOR2_X1 U8414 ( .A(n6744), .B(n7770), .ZN(n9950) );
  AOI21_X1 U8415 ( .B1(n6746), .B2(n6745), .A(n8292), .ZN(n6748) );
  OAI22_X1 U8416 ( .A1(n6758), .A2(n9861), .B1(n8333), .B2(n9863), .ZN(n6747)
         );
  AOI21_X1 U8417 ( .B1(n6748), .B2(n4255), .A(n6747), .ZN(n9949) );
  OAI22_X1 U8418 ( .A1(n4247), .A2(n9949), .B1(n6757), .B2(n8272), .ZN(n6749)
         );
  AOI21_X1 U8419 ( .B1(n4247), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6749), .ZN(
        n6751) );
  XNOR2_X1 U8420 ( .A(n9870), .B(n6759), .ZN(n9947) );
  AOI22_X1 U8421 ( .A1(n8319), .A2(n9947), .B1(n8324), .B2(n9945), .ZN(n6750)
         );
  OAI211_X1 U8422 ( .C1(n9950), .C2(n8321), .A(n6751), .B(n6750), .ZN(P2_U3292) );
  INV_X1 U8423 ( .A(n6754), .ZN(n6755) );
  AOI21_X1 U8424 ( .B1(n6752), .B2(n6756), .A(n6755), .ZN(n6763) );
  NAND2_X1 U8425 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7991) );
  OAI21_X1 U8426 ( .B1(n7925), .B2(n6757), .A(n7991), .ZN(n6761) );
  OAI22_X1 U8427 ( .A1(n6759), .A2(n7945), .B1(n7939), .B2(n6758), .ZN(n6760)
         );
  AOI211_X1 U8428 ( .C1(n6775), .C2(n7960), .A(n6761), .B(n6760), .ZN(n6762)
         );
  OAI21_X1 U8429 ( .B1(n6763), .B2(n7931), .A(n6762), .ZN(P2_U3232) );
  XNOR2_X1 U8430 ( .A(n6764), .B(n6765), .ZN(n6770) );
  NOR2_X1 U8431 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4922), .ZN(n7977) );
  INV_X1 U8432 ( .A(n7977), .ZN(n6766) );
  OAI21_X1 U8433 ( .B1(n7925), .B2(P2_REG3_REG_3__SCAN_IN), .A(n6766), .ZN(
        n6768) );
  OAI22_X1 U8434 ( .A1(n9872), .A2(n7945), .B1(n7939), .B2(n9862), .ZN(n6767)
         );
  AOI211_X1 U8435 ( .C1(n6775), .C2(n4248), .A(n6768), .B(n6767), .ZN(n6769)
         );
  OAI21_X1 U8436 ( .B1(n7931), .B2(n6770), .A(n6769), .ZN(P2_U3220) );
  XNOR2_X1 U8437 ( .A(n6772), .B(n6771), .ZN(n6777) );
  INV_X1 U8438 ( .A(n6949), .ZN(n7957) );
  OAI22_X1 U8439 ( .A1(n7925), .A2(n6955), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9410), .ZN(n6774) );
  INV_X1 U8440 ( .A(n7056), .ZN(n6956) );
  OAI22_X1 U8441 ( .A1(n6956), .A2(n7945), .B1(n7939), .B2(n7157), .ZN(n6773)
         );
  AOI211_X1 U8442 ( .C1(n6775), .C2(n7957), .A(n6774), .B(n6773), .ZN(n6776)
         );
  OAI21_X1 U8443 ( .B1(n6777), .B2(n7931), .A(n6776), .ZN(P2_U3215) );
  NAND2_X1 U8444 ( .A1(n8278), .A2(n8307), .ZN(n9878) );
  NAND2_X1 U8445 ( .A1(n6918), .A2(n7651), .ZN(n7769) );
  INV_X1 U8446 ( .A(n7769), .ZN(n9923) );
  NAND2_X1 U8447 ( .A1(n7769), .A2(n9865), .ZN(n6779) );
  OR2_X1 U8448 ( .A1(n6705), .A2(n9861), .ZN(n6778) );
  NAND2_X1 U8449 ( .A1(n6779), .A2(n6778), .ZN(n9924) );
  INV_X1 U8450 ( .A(n8272), .ZN(n9869) );
  AOI22_X1 U8451 ( .A1(n8336), .A2(n9924), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n9869), .ZN(n6781) );
  OR2_X1 U8452 ( .A1(n8336), .A2(n4874), .ZN(n6780) );
  OAI211_X1 U8453 ( .C1(n8321), .C2(n9923), .A(n6781), .B(n6780), .ZN(n6782)
         );
  AOI21_X1 U8454 ( .B1(n6917), .B2(n9878), .A(n6782), .ZN(n6783) );
  INV_X1 U8455 ( .A(n6783), .ZN(P2_U3296) );
  INV_X1 U8456 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6785) );
  INV_X1 U8457 ( .A(n6784), .ZN(n6786) );
  INV_X1 U8458 ( .A(n9698), .ZN(n8959) );
  OAI222_X1 U8459 ( .A1(n7852), .A2(n6785), .B1(n4249), .B2(n6786), .C1(
        P1_U3084), .C2(n8959), .ZN(P1_U3335) );
  INV_X1 U8460 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6787) );
  INV_X1 U8461 ( .A(n7285), .ZN(n8069) );
  OAI222_X1 U8462 ( .A1(n8465), .A2(n6787), .B1(n8467), .B2(n6786), .C1(
        P2_U3152), .C2(n8069), .ZN(P2_U3340) );
  NOR2_X1 U8463 ( .A1(n6789), .A2(n6788), .ZN(n6791) );
  NOR2_X1 U8464 ( .A1(n6791), .A2(n6790), .ZN(n6794) );
  XNOR2_X1 U8465 ( .A(n7089), .B(n6792), .ZN(n6793) );
  NAND2_X1 U8466 ( .A1(n6793), .A2(n6794), .ZN(n7088) );
  OAI21_X1 U8467 ( .B1(n6794), .B2(n6793), .A(n7088), .ZN(n6797) );
  NAND2_X1 U8468 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7587) );
  NAND2_X1 U8469 ( .A1(n9850), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n6795) );
  OAI211_X1 U8470 ( .C1(n9847), .C2(n6803), .A(n7587), .B(n6795), .ZN(n6796)
         );
  AOI21_X1 U8471 ( .B1(n6797), .B2(n9845), .A(n6796), .ZN(n6807) );
  NOR2_X1 U8472 ( .A1(n6799), .A2(n6798), .ZN(n6801) );
  NOR2_X1 U8473 ( .A1(n6801), .A2(n6800), .ZN(n6805) );
  NAND2_X1 U8474 ( .A1(n7089), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7084) );
  INV_X1 U8475 ( .A(n7084), .ZN(n6802) );
  AOI21_X1 U8476 ( .B1(n7531), .B2(n6803), .A(n6802), .ZN(n6804) );
  NAND2_X1 U8477 ( .A1(n6804), .A2(n6805), .ZN(n7083) );
  OAI211_X1 U8478 ( .C1(n6805), .C2(n6804), .A(n9844), .B(n7083), .ZN(n6806)
         );
  NAND2_X1 U8479 ( .A1(n6807), .A2(n6806), .ZN(P2_U3261) );
  INV_X1 U8480 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6814) );
  OAI21_X1 U8481 ( .B1(n6809), .B2(n9222), .A(n6808), .ZN(n6810) );
  NAND2_X1 U8482 ( .A1(n6810), .A2(n9762), .ZN(n6813) );
  OAI21_X1 U8483 ( .B1(n9718), .B2(n9226), .A(n6811), .ZN(n6812) );
  OAI211_X1 U8484 ( .C1(n6814), .C2(n9762), .A(n6813), .B(n6812), .ZN(P1_U3291) );
  NAND2_X1 U8485 ( .A1(n9725), .A2(n9778), .ZN(n6815) );
  NAND2_X1 U8486 ( .A1(n6816), .A2(n6815), .ZN(n9712) );
  NAND2_X1 U8487 ( .A1(n6821), .A2(n9713), .ZN(n8849) );
  NAND2_X1 U8488 ( .A1(n8849), .A2(n8843), .ZN(n9721) );
  NAND2_X1 U8489 ( .A1(n9712), .A2(n9721), .ZN(n6818) );
  NAND2_X1 U8490 ( .A1(n6821), .A2(n9784), .ZN(n6817) );
  NAND2_X1 U8491 ( .A1(n6818), .A2(n6817), .ZN(n6849) );
  NAND2_X1 U8492 ( .A1(n9722), .A2(n6830), .ZN(n8848) );
  INV_X1 U8493 ( .A(n6830), .ZN(n9791) );
  NAND2_X1 U8494 ( .A1(n9791), .A2(n8898), .ZN(n8852) );
  NAND2_X1 U8495 ( .A1(n8848), .A2(n8852), .ZN(n6848) );
  INV_X1 U8496 ( .A(n6848), .ZN(n8728) );
  XNOR2_X1 U8497 ( .A(n6849), .B(n8728), .ZN(n9790) );
  NAND2_X1 U8498 ( .A1(n8847), .A2(n8849), .ZN(n6839) );
  XNOR2_X1 U8499 ( .A(n6839), .B(n8728), .ZN(n6823) );
  OAI22_X1 U8500 ( .A1(n6821), .A2(n9724), .B1(n9723), .B2(n7034), .ZN(n6822)
         );
  AOI21_X1 U8501 ( .B1(n6823), .B2(n9727), .A(n6822), .ZN(n6824) );
  OAI21_X1 U8502 ( .B1(n9790), .B2(n9759), .A(n6824), .ZN(n9793) );
  NAND2_X1 U8503 ( .A1(n9793), .A2(n9762), .ZN(n6832) );
  INV_X1 U8504 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6826) );
  OAI22_X1 U8505 ( .A1(n9762), .A2(n6826), .B1(n6825), .B2(n9222), .ZN(n6829)
         );
  INV_X1 U8506 ( .A(n9716), .ZN(n6827) );
  OAI21_X1 U8507 ( .B1(n6827), .B2(n9791), .A(n6882), .ZN(n9792) );
  NOR2_X1 U8508 ( .A1(n9042), .A2(n9792), .ZN(n6828) );
  AOI211_X1 U8509 ( .C1(n9226), .C2(n6830), .A(n6829), .B(n6828), .ZN(n6831)
         );
  OAI211_X1 U8510 ( .C1(n9790), .C2(n9276), .A(n6832), .B(n6831), .ZN(P1_U3287) );
  XNOR2_X1 U8511 ( .A(n6834), .B(n6833), .ZN(n6838) );
  NAND2_X1 U8512 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n8042) );
  OAI21_X1 U8513 ( .B1(n7925), .B2(n6974), .A(n8042), .ZN(n6836) );
  OAI22_X1 U8514 ( .A1(n7162), .A2(n7939), .B1(n7938), .B2(n6970), .ZN(n6835)
         );
  AOI211_X1 U8515 ( .C1(n9969), .C2(n7929), .A(n6836), .B(n6835), .ZN(n6837)
         );
  OAI21_X1 U8516 ( .B1(n6838), .B2(n7931), .A(n6837), .ZN(P2_U3223) );
  OR2_X1 U8517 ( .A1(n6998), .A2(n7152), .ZN(n8798) );
  NAND2_X1 U8518 ( .A1(n6998), .A2(n7152), .ZN(n8619) );
  NAND2_X1 U8519 ( .A1(n8798), .A2(n8619), .ZN(n7000) );
  INV_X1 U8520 ( .A(n7000), .ZN(n8732) );
  OAI21_X1 U8521 ( .B1(n6839), .B2(n6848), .A(n8852), .ZN(n6879) );
  NAND2_X1 U8522 ( .A1(n7034), .A2(n6892), .ZN(n8851) );
  INV_X1 U8523 ( .A(n6892), .ZN(n9800) );
  NAND2_X1 U8524 ( .A1(n9800), .A2(n8897), .ZN(n8795) );
  NAND2_X1 U8525 ( .A1(n9804), .A2(n8896), .ZN(n8796) );
  INV_X1 U8526 ( .A(n8796), .ZN(n6840) );
  NAND2_X1 U8527 ( .A1(n6881), .A2(n6875), .ZN(n8850) );
  OAI21_X1 U8528 ( .B1(n8732), .B2(n6841), .A(n6995), .ZN(n6842) );
  AOI222_X1 U8529 ( .A1(n9727), .A2(n6842), .B1(n8894), .B2(n9756), .C1(n8896), 
        .C2(n9739), .ZN(n9811) );
  NAND2_X1 U8530 ( .A1(n6884), .A2(n9804), .ZN(n6872) );
  INV_X1 U8531 ( .A(n6872), .ZN(n6843) );
  INV_X1 U8532 ( .A(n6998), .ZN(n9812) );
  OAI211_X1 U8533 ( .C1(n6843), .C2(n9812), .A(n9742), .B(n7005), .ZN(n9810)
         );
  INV_X1 U8534 ( .A(n9810), .ZN(n6847) );
  NOR2_X1 U8535 ( .A1(n6844), .A2(n9744), .ZN(n9289) );
  INV_X1 U8536 ( .A(n9222), .ZN(n9747) );
  AOI22_X1 U8537 ( .A1(n9234), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n6992), .B2(
        n9747), .ZN(n6845) );
  OAI21_X1 U8538 ( .B1(n9812), .B2(n9733), .A(n6845), .ZN(n6846) );
  AOI21_X1 U8539 ( .B1(n6847), .B2(n9289), .A(n6846), .ZN(n6859) );
  NAND2_X1 U8540 ( .A1(n6849), .A2(n6848), .ZN(n6851) );
  NAND2_X1 U8541 ( .A1(n9722), .A2(n9791), .ZN(n6850) );
  NAND2_X1 U8542 ( .A1(n6851), .A2(n6850), .ZN(n6888) );
  NAND2_X1 U8543 ( .A1(n8897), .A2(n6892), .ZN(n6853) );
  OR2_X1 U8544 ( .A1(n8896), .A2(n6875), .ZN(n6854) );
  XNOR2_X1 U8545 ( .A(n7001), .B(n7000), .ZN(n9814) );
  NOR2_X1 U8546 ( .A1(n6856), .A2(n6855), .ZN(n6857) );
  INV_X1 U8547 ( .A(n9297), .ZN(n9220) );
  NAND2_X1 U8548 ( .A1(n9814), .A2(n9220), .ZN(n6858) );
  OAI211_X1 U8549 ( .C1(n9811), .C2(n9291), .A(n6859), .B(n6858), .ZN(P1_U3284) );
  INV_X1 U8550 ( .A(n6860), .ZN(n6862) );
  OAI222_X1 U8551 ( .A1(n7852), .A2(n6861), .B1(n4249), .B2(n6862), .C1(n5638), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  OAI222_X1 U8552 ( .A1(n8465), .A2(n6863), .B1(n8467), .B2(n6862), .C1(
        P2_U3152), .C2(n7839), .ZN(P2_U3339) );
  INV_X1 U8553 ( .A(n8729), .ZN(n6868) );
  OAI21_X1 U8554 ( .B1(n6865), .B2(n6868), .A(n6864), .ZN(n9808) );
  INV_X1 U8555 ( .A(n9808), .ZN(n6878) );
  OR2_X1 U8556 ( .A1(n6867), .A2(n6868), .ZN(n8613) );
  INV_X1 U8557 ( .A(n8613), .ZN(n6866) );
  AOI21_X1 U8558 ( .B1(n6868), .B2(n6867), .A(n6866), .ZN(n6869) );
  OAI222_X1 U8559 ( .A1(n9723), .A2(n7152), .B1(n9724), .B2(n7034), .C1(n9751), 
        .C2(n6869), .ZN(n9806) );
  NAND2_X1 U8560 ( .A1(n9806), .A2(n9762), .ZN(n6877) );
  INV_X1 U8561 ( .A(n7036), .ZN(n6870) );
  OAI22_X1 U8562 ( .A1(n9762), .A2(n9415), .B1(n6870), .B2(n9222), .ZN(n6874)
         );
  OR2_X1 U8563 ( .A1(n6884), .A2(n9804), .ZN(n6871) );
  NAND2_X1 U8564 ( .A1(n6872), .A2(n6871), .ZN(n9805) );
  NOR2_X1 U8565 ( .A1(n9805), .A2(n9042), .ZN(n6873) );
  AOI211_X1 U8566 ( .C1(n9226), .C2(n6875), .A(n6874), .B(n6873), .ZN(n6876)
         );
  OAI211_X1 U8567 ( .C1(n9297), .C2(n6878), .A(n6877), .B(n6876), .ZN(P1_U3285) );
  XNOR2_X1 U8568 ( .A(n6879), .B(n8727), .ZN(n6880) );
  OAI222_X1 U8569 ( .A1(n9723), .A2(n6881), .B1(n9724), .B2(n9722), .C1(n9751), 
        .C2(n6880), .ZN(n9802) );
  AND2_X1 U8570 ( .A1(n9762), .A2(n5638), .ZN(n9152) );
  INV_X1 U8571 ( .A(n9152), .ZN(n6895) );
  NAND2_X1 U8572 ( .A1(n6882), .A2(n6892), .ZN(n6883) );
  NAND2_X1 U8573 ( .A1(n6883), .A2(n9742), .ZN(n6885) );
  OR2_X1 U8574 ( .A1(n6885), .A2(n6884), .ZN(n9798) );
  NAND2_X1 U8575 ( .A1(n6888), .A2(n8727), .ZN(n9797) );
  NAND3_X1 U8576 ( .A1(n6887), .A2(n9797), .A3(n9220), .ZN(n6894) );
  INV_X1 U8577 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6890) );
  INV_X1 U8578 ( .A(n7020), .ZN(n6889) );
  OAI22_X1 U8579 ( .A1(n9762), .A2(n6890), .B1(n6889), .B2(n9222), .ZN(n6891)
         );
  AOI21_X1 U8580 ( .B1(n9226), .B2(n6892), .A(n6891), .ZN(n6893) );
  OAI211_X1 U8581 ( .C1(n6895), .C2(n9798), .A(n6894), .B(n6893), .ZN(n6896)
         );
  AOI21_X1 U8582 ( .B1(n9802), .B2(n9762), .A(n6896), .ZN(n6897) );
  INV_X1 U8583 ( .A(n6897), .ZN(P1_U3286) );
  NAND2_X1 U8584 ( .A1(n6949), .A2(n6944), .ZN(n7662) );
  NAND2_X1 U8585 ( .A1(n9960), .A2(n7957), .ZN(n7661) );
  NAND2_X1 U8586 ( .A1(n7662), .A2(n7661), .ZN(n7773) );
  INV_X1 U8587 ( .A(n7773), .ZN(n6912) );
  NAND2_X1 U8588 ( .A1(n4255), .A2(n7635), .ZN(n6899) );
  NAND2_X1 U8589 ( .A1(n6899), .A2(n7641), .ZN(n6900) );
  OAI21_X1 U8590 ( .B1(n6912), .B2(n6900), .A(n6947), .ZN(n6903) );
  NAND2_X1 U8591 ( .A1(n7958), .A2(n8312), .ZN(n6901) );
  OAI21_X1 U8592 ( .B1(n6970), .B2(n9861), .A(n6901), .ZN(n6902) );
  AOI21_X1 U8593 ( .B1(n6903), .B2(n9865), .A(n6902), .ZN(n9966) );
  OAI22_X1 U8594 ( .A1(n8272), .A2(n6904), .B1(n6520), .B2(n8336), .ZN(n6908)
         );
  AND2_X1 U8595 ( .A1(n6905), .A2(n9960), .ZN(n6952) );
  NOR2_X1 U8596 ( .A1(n6905), .A2(n9960), .ZN(n6906) );
  OR2_X1 U8597 ( .A1(n6952), .A2(n6906), .ZN(n9961) );
  NOR2_X1 U8598 ( .A1(n8278), .A2(n9961), .ZN(n6907) );
  AOI211_X1 U8599 ( .C1(n8324), .C2(n6944), .A(n6908), .B(n6907), .ZN(n6914)
         );
  XNOR2_X1 U8600 ( .A(n6946), .B(n6912), .ZN(n9963) );
  NAND2_X1 U8601 ( .A1(n9963), .A2(n8325), .ZN(n6913) );
  OAI211_X1 U8602 ( .C1(n4247), .C2(n9966), .A(n6914), .B(n6913), .ZN(P2_U3290) );
  XNOR2_X1 U8603 ( .A(n6916), .B(n6915), .ZN(n9933) );
  AOI22_X1 U8604 ( .A1(n8325), .A2(n9933), .B1(n8324), .B2(n6584), .ZN(n6924)
         );
  AOI211_X1 U8605 ( .C1(n6917), .C2(n6584), .A(n9985), .B(n8326), .ZN(n9927)
         );
  XNOR2_X1 U8606 ( .A(n6915), .B(n6918), .ZN(n6920) );
  AOI21_X1 U8607 ( .B1(n6920), .B2(n9865), .A(n6919), .ZN(n9930) );
  OAI21_X1 U8608 ( .B1(n6921), .B2(n8272), .A(n9930), .ZN(n6922) );
  AOI22_X1 U8609 ( .A1(n8328), .A2(n9927), .B1(n8336), .B2(n6922), .ZN(n6923)
         );
  OAI211_X1 U8610 ( .C1(n6925), .C2(n8336), .A(n6924), .B(n6923), .ZN(P2_U3295) );
  INV_X1 U8611 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6943) );
  OR2_X1 U8612 ( .A1(n7266), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6927) );
  NAND2_X1 U8613 ( .A1(n7266), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6926) );
  AND2_X1 U8614 ( .A1(n6927), .A2(n6926), .ZN(n6931) );
  OAI21_X1 U8615 ( .B1(n6934), .B2(P1_REG1_REG_11__SCAN_IN), .A(n6928), .ZN(
        n8926) );
  INV_X1 U8616 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6929) );
  MUX2_X1 U8617 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6929), .S(n8934), .Z(n8927)
         );
  NAND2_X1 U8618 ( .A1(n8926), .A2(n8927), .ZN(n8925) );
  OAI21_X1 U8619 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n8934), .A(n8925), .ZN(
        n6930) );
  NAND2_X1 U8620 ( .A1(n6930), .A2(n6931), .ZN(n7261) );
  OAI21_X1 U8621 ( .B1(n6931), .B2(n6930), .A(n7261), .ZN(n6940) );
  INV_X1 U8622 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6933) );
  NOR2_X1 U8623 ( .A1(n7266), .A2(n6933), .ZN(n6932) );
  AOI21_X1 U8624 ( .B1(n7266), .B2(n6933), .A(n6932), .ZN(n6938) );
  OR2_X1 U8625 ( .A1(n6934), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6936) );
  NAND2_X1 U8626 ( .A1(n6936), .A2(n6935), .ZN(n8929) );
  XNOR2_X1 U8627 ( .A(n8934), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n8930) );
  AOI211_X1 U8628 ( .C1(n6938), .C2(n6937), .A(n7265), .B(n9679), .ZN(n6939)
         );
  AOI21_X1 U8629 ( .B1(n9707), .B2(n6940), .A(n6939), .ZN(n6942) );
  AND2_X1 U8630 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7430) );
  AOI21_X1 U8631 ( .B1(n9699), .B2(n7266), .A(n7430), .ZN(n6941) );
  OAI211_X1 U8632 ( .C1(n9689), .C2(n6943), .A(n6942), .B(n6941), .ZN(P1_U3254) );
  AND2_X1 U8633 ( .A1(n7957), .A2(n6944), .ZN(n6945) );
  OR2_X1 U8634 ( .A1(n7056), .A2(n6970), .ZN(n7666) );
  NAND2_X1 U8635 ( .A1(n7056), .A2(n6970), .ZN(n7665) );
  NAND2_X1 U8636 ( .A1(n7666), .A2(n7665), .ZN(n7774) );
  XNOR2_X1 U8637 ( .A(n6960), .B(n4400), .ZN(n7058) );
  XNOR2_X1 U8638 ( .A(n6968), .B(n7774), .ZN(n6948) );
  OAI222_X1 U8639 ( .A1(n9861), .A2(n7157), .B1(n9863), .B2(n6949), .C1(n6948), 
        .C2(n8292), .ZN(n7054) );
  INV_X1 U8640 ( .A(n7054), .ZN(n6950) );
  MUX2_X1 U8641 ( .A(n6951), .B(n6950), .S(n8336), .Z(n6959) );
  INV_X1 U8642 ( .A(n6952), .ZN(n6954) );
  INV_X1 U8643 ( .A(n6976), .ZN(n6953) );
  AOI211_X1 U8644 ( .C1(n7056), .C2(n6954), .A(n9985), .B(n6953), .ZN(n7055)
         );
  OAI22_X1 U8645 ( .A1(n8307), .A2(n6956), .B1(n8272), .B2(n6955), .ZN(n6957)
         );
  AOI21_X1 U8646 ( .B1(n8328), .B2(n7055), .A(n6957), .ZN(n6958) );
  OAI211_X1 U8647 ( .C1(n8321), .C2(n7058), .A(n6959), .B(n6958), .ZN(P2_U3289) );
  INV_X1 U8648 ( .A(n6970), .ZN(n7956) );
  OR2_X1 U8649 ( .A1(n7056), .A2(n7956), .ZN(n6961) );
  INV_X1 U8650 ( .A(n6964), .ZN(n6963) );
  OR2_X1 U8651 ( .A1(n9969), .A2(n7157), .ZN(n7668) );
  NAND2_X1 U8652 ( .A1(n9969), .A2(n7157), .ZN(n7669) );
  NAND2_X1 U8653 ( .A1(n6963), .A2(n6962), .ZN(n7159) );
  NAND2_X1 U8654 ( .A1(n6964), .A2(n7776), .ZN(n6965) );
  NAND2_X1 U8655 ( .A1(n7159), .A2(n6965), .ZN(n9968) );
  INV_X1 U8656 ( .A(n6966), .ZN(n6967) );
  NAND2_X1 U8657 ( .A1(n8336), .A2(n6967), .ZN(n9876) );
  NAND2_X1 U8658 ( .A1(n6969), .A2(n7776), .ZN(n7165) );
  OAI21_X1 U8659 ( .B1(n7776), .B2(n6969), .A(n7165), .ZN(n6972) );
  OAI22_X1 U8660 ( .A1(n6970), .A2(n9863), .B1(n7162), .B2(n9861), .ZN(n6971)
         );
  AOI21_X1 U8661 ( .B1(n6972), .B2(n9865), .A(n6971), .ZN(n6973) );
  OAI21_X1 U8662 ( .B1(n9854), .B2(n9968), .A(n6973), .ZN(n9972) );
  NAND2_X1 U8663 ( .A1(n9972), .A2(n8336), .ZN(n6981) );
  OAI22_X1 U8664 ( .A1(n8336), .A2(n6975), .B1(n6974), .B2(n8272), .ZN(n6979)
         );
  NAND2_X1 U8665 ( .A1(n6976), .A2(n9969), .ZN(n6977) );
  NAND2_X1 U8666 ( .A1(n4420), .A2(n6977), .ZN(n9971) );
  NOR2_X1 U8667 ( .A1(n8278), .A2(n9971), .ZN(n6978) );
  AOI211_X1 U8668 ( .C1(n8324), .C2(n9969), .A(n6979), .B(n6978), .ZN(n6980)
         );
  OAI211_X1 U8669 ( .C1(n9968), .C2(n9876), .A(n6981), .B(n6980), .ZN(P2_U3288) );
  INV_X1 U8670 ( .A(n6982), .ZN(n7030) );
  INV_X1 U8671 ( .A(n6983), .ZN(n6985) );
  NOR3_X1 U8672 ( .A1(n7030), .A2(n6985), .A3(n6984), .ZN(n6988) );
  INV_X1 U8673 ( .A(n6986), .ZN(n6987) );
  OAI21_X1 U8674 ( .B1(n6988), .B2(n6987), .A(n8571), .ZN(n6994) );
  AOI21_X1 U8675 ( .B1(n8585), .B2(n8896), .A(n6989), .ZN(n6990) );
  OAI21_X1 U8676 ( .B1(n8588), .B2(n7235), .A(n6990), .ZN(n6991) );
  AOI21_X1 U8677 ( .B1(n6992), .B2(n8583), .A(n6991), .ZN(n6993) );
  OAI211_X1 U8678 ( .C1(n9812), .C2(n8578), .A(n6994), .B(n6993), .ZN(P1_U3211) );
  OR2_X1 U8679 ( .A1(n7154), .A2(n7235), .ZN(n8805) );
  NAND2_X1 U8680 ( .A1(n7154), .A2(n7235), .ZN(n8631) );
  NAND2_X1 U8681 ( .A1(n8805), .A2(n8631), .ZN(n7179) );
  INV_X1 U8682 ( .A(n7179), .ZN(n8733) );
  NAND2_X1 U8683 ( .A1(n6995), .A2(n8619), .ZN(n6996) );
  NAND2_X1 U8684 ( .A1(n6996), .A2(n8733), .ZN(n7097) );
  OAI21_X1 U8685 ( .B1(n8733), .B2(n6996), .A(n7097), .ZN(n6997) );
  AOI222_X1 U8686 ( .A1(n9727), .A2(n6997), .B1(n8893), .B2(n9756), .C1(n8895), 
        .C2(n9739), .ZN(n7070) );
  NOR2_X1 U8687 ( .A1(n6998), .A2(n8895), .ZN(n6999) );
  NAND2_X1 U8688 ( .A1(n7185), .A2(n7179), .ZN(n7128) );
  OAI21_X1 U8689 ( .B1(n7185), .B2(n7179), .A(n7128), .ZN(n7071) );
  INV_X1 U8690 ( .A(n7148), .ZN(n7002) );
  OAI22_X1 U8691 ( .A1(n9762), .A2(n7003), .B1(n7002), .B2(n9222), .ZN(n7004)
         );
  AOI21_X1 U8692 ( .B1(n9226), .B2(n7154), .A(n7004), .ZN(n7009) );
  NOR2_X1 U8693 ( .A1(n7005), .A2(n7154), .ZN(n7102) );
  NAND2_X1 U8694 ( .A1(n7005), .A2(n7154), .ZN(n7006) );
  NAND2_X1 U8695 ( .A1(n7006), .A2(n9742), .ZN(n7007) );
  NOR2_X1 U8696 ( .A1(n7102), .A2(n7007), .ZN(n7068) );
  NAND2_X1 U8697 ( .A1(n7068), .A2(n9152), .ZN(n7008) );
  OAI211_X1 U8698 ( .C1(n7071), .C2(n9297), .A(n7009), .B(n7008), .ZN(n7010)
         );
  INV_X1 U8699 ( .A(n7010), .ZN(n7011) );
  OAI21_X1 U8700 ( .B1(n7070), .B2(n9234), .A(n7011), .ZN(P1_U3283) );
  INV_X1 U8701 ( .A(n7012), .ZN(n7014) );
  NOR2_X1 U8702 ( .A1(n7014), .A2(n7013), .ZN(n7026) );
  AOI21_X1 U8703 ( .B1(n7014), .B2(n7013), .A(n7026), .ZN(n7015) );
  NAND2_X1 U8704 ( .A1(n7015), .A2(n7016), .ZN(n7029) );
  OAI21_X1 U8705 ( .B1(n7016), .B2(n7015), .A(n7029), .ZN(n7017) );
  NAND2_X1 U8706 ( .A1(n7017), .A2(n8571), .ZN(n7022) );
  AND2_X1 U8707 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9653) );
  AOI21_X1 U8708 ( .B1(n8552), .B2(n8896), .A(n9653), .ZN(n7018) );
  OAI21_X1 U8709 ( .B1(n8573), .B2(n9722), .A(n7018), .ZN(n7019) );
  AOI21_X1 U8710 ( .B1(n7020), .B2(n8583), .A(n7019), .ZN(n7021) );
  OAI211_X1 U8711 ( .C1(n9800), .C2(n8578), .A(n7022), .B(n7021), .ZN(P1_U3225) );
  INV_X1 U8712 ( .A(n7023), .ZN(n7024) );
  OAI222_X1 U8713 ( .A1(P1_U3084), .A2(n8877), .B1(n4249), .B2(n7024), .C1(
        n9348), .C2(n7852), .ZN(P1_U3333) );
  OAI222_X1 U8714 ( .A1(n8465), .A2(n7025), .B1(n8467), .B2(n7024), .C1(n4866), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  INV_X1 U8715 ( .A(n7026), .ZN(n7027) );
  AND3_X1 U8716 ( .A1(n7029), .A2(n7028), .A3(n7027), .ZN(n7031) );
  OAI21_X1 U8717 ( .B1(n7031), .B2(n7030), .A(n8571), .ZN(n7038) );
  AOI21_X1 U8718 ( .B1(n8552), .B2(n8895), .A(n7032), .ZN(n7033) );
  OAI21_X1 U8719 ( .B1(n8573), .B2(n7034), .A(n7033), .ZN(n7035) );
  AOI21_X1 U8720 ( .B1(n7036), .B2(n8583), .A(n7035), .ZN(n7037) );
  OAI211_X1 U8721 ( .C1(n9804), .C2(n8578), .A(n7038), .B(n7037), .ZN(P1_U3237) );
  OR2_X1 U8722 ( .A1(n7039), .A2(n7041), .ZN(n7109) );
  INV_X1 U8723 ( .A(n7109), .ZN(n7040) );
  AOI21_X1 U8724 ( .B1(n7039), .B2(n7041), .A(n7040), .ZN(n7045) );
  NAND2_X1 U8725 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8055) );
  OAI21_X1 U8726 ( .B1(n7925), .B2(n7209), .A(n8055), .ZN(n7043) );
  OAI22_X1 U8727 ( .A1(n7203), .A2(n7939), .B1(n7938), .B2(n7157), .ZN(n7042)
         );
  AOI211_X1 U8728 ( .C1(n8434), .C2(n7929), .A(n7043), .B(n7042), .ZN(n7044)
         );
  OAI21_X1 U8729 ( .B1(n7045), .B2(n7931), .A(n7044), .ZN(P2_U3233) );
  INV_X1 U8730 ( .A(n7046), .ZN(n7048) );
  OAI222_X1 U8731 ( .A1(P1_U3084), .A2(n8753), .B1(n4249), .B2(n7048), .C1(
        n7047), .C2(n7852), .ZN(P1_U3332) );
  OAI222_X1 U8732 ( .A1(n8465), .A2(n7049), .B1(n8467), .B2(n7048), .C1(n7827), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  AND2_X1 U8733 ( .A1(n7061), .A2(n7062), .ZN(n7050) );
  AND2_X1 U8734 ( .A1(n4866), .A2(n8077), .ZN(n7053) );
  NAND2_X1 U8735 ( .A1(n7053), .A2(n7052), .ZN(n9967) );
  AOI211_X1 U8736 ( .C1(n9954), .C2(n7056), .A(n7055), .B(n7054), .ZN(n7057)
         );
  OAI21_X1 U8737 ( .B1(n9957), .B2(n7058), .A(n7057), .ZN(n7066) );
  NAND2_X1 U8738 ( .A1(n7066), .A2(n9993), .ZN(n7059) );
  OAI21_X1 U8739 ( .B1(n9993), .B2(n5002), .A(n7059), .ZN(P2_U3472) );
  AND4_X1 U8740 ( .A1(n7063), .A2(n7062), .A3(n7061), .A4(n7060), .ZN(n7064)
         );
  NAND2_X1 U8741 ( .A1(n7066), .A2(n10008), .ZN(n7067) );
  OAI21_X1 U8742 ( .B1(n10008), .B2(n9437), .A(n7067), .ZN(P2_U3527) );
  INV_X1 U8743 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7073) );
  NAND2_X2 U8744 ( .A1(n5639), .A2(n9744), .ZN(n8705) );
  AOI21_X1 U8745 ( .B1(n9598), .B2(n7154), .A(n7068), .ZN(n7069) );
  OAI211_X1 U8746 ( .C1(n9524), .C2(n7071), .A(n7070), .B(n7069), .ZN(n7074)
         );
  NAND2_X1 U8747 ( .A1(n7074), .A2(n9843), .ZN(n7072) );
  OAI21_X1 U8748 ( .B1(n9843), .B2(n7073), .A(n7072), .ZN(P1_U3531) );
  INV_X1 U8749 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7076) );
  NAND2_X1 U8750 ( .A1(n7074), .A2(n9828), .ZN(n7075) );
  OAI21_X1 U8751 ( .B1(n9828), .B2(n7076), .A(n7075), .ZN(P1_U3478) );
  XNOR2_X1 U8752 ( .A(n7078), .B(n7077), .ZN(n7082) );
  OAI22_X1 U8753 ( .A1(n7925), .A2(n7351), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5094), .ZN(n7080) );
  OAI22_X1 U8754 ( .A1(n7365), .A2(n7939), .B1(n7938), .B2(n7203), .ZN(n7079)
         );
  AOI211_X1 U8755 ( .C1(n8429), .C2(n7929), .A(n7080), .B(n7079), .ZN(n7081)
         );
  OAI21_X1 U8756 ( .B1(n7082), .B2(n7931), .A(n7081), .ZN(P2_U3238) );
  NAND2_X1 U8757 ( .A1(n7084), .A2(n7083), .ZN(n7087) );
  NAND2_X1 U8758 ( .A1(n7280), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7275) );
  INV_X1 U8759 ( .A(n7275), .ZN(n7085) );
  AOI21_X1 U8760 ( .B1(n7577), .B2(n7095), .A(n7085), .ZN(n7086) );
  NAND2_X1 U8761 ( .A1(n7086), .A2(n7087), .ZN(n7274) );
  OAI211_X1 U8762 ( .C1(n7087), .C2(n7086), .A(n9844), .B(n7274), .ZN(n7094)
         );
  AND2_X1 U8763 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7888) );
  OAI21_X1 U8764 ( .B1(n7089), .B2(P2_REG1_REG_16__SCAN_IN), .A(n7088), .ZN(
        n7091) );
  XNOR2_X1 U8765 ( .A(n7280), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n7090) );
  NOR2_X1 U8766 ( .A1(n7090), .A2(n7091), .ZN(n7279) );
  AOI211_X1 U8767 ( .C1(n7091), .C2(n7090), .A(n7279), .B(n7283), .ZN(n7092)
         );
  AOI211_X1 U8768 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n9850), .A(n7888), .B(
        n7092), .ZN(n7093) );
  OAI211_X1 U8769 ( .C1(n9847), .C2(n7095), .A(n7094), .B(n7093), .ZN(P2_U3262) );
  NAND2_X1 U8770 ( .A1(n7154), .A2(n8894), .ZN(n7125) );
  NAND2_X1 U8771 ( .A1(n7128), .A2(n7125), .ZN(n7096) );
  OR2_X1 U8772 ( .A1(n8623), .A2(n8893), .ZN(n7129) );
  NAND2_X1 U8773 ( .A1(n8623), .A2(n8893), .ZN(n7124) );
  NAND2_X1 U8774 ( .A1(n7129), .A2(n7124), .ZN(n8731) );
  XNOR2_X1 U8775 ( .A(n7096), .B(n8731), .ZN(n9823) );
  NAND2_X1 U8776 ( .A1(n9823), .A2(n9270), .ZN(n7101) );
  NAND2_X1 U8777 ( .A1(n7097), .A2(n8631), .ZN(n7120) );
  XNOR2_X1 U8778 ( .A(n7120), .B(n8731), .ZN(n7099) );
  OAI22_X1 U8779 ( .A1(n7187), .A2(n9723), .B1(n9724), .B2(n7235), .ZN(n7098)
         );
  AOI21_X1 U8780 ( .B1(n7099), .B2(n9727), .A(n7098), .ZN(n7100) );
  INV_X1 U8781 ( .A(n9276), .ZN(n9719) );
  INV_X1 U8782 ( .A(n8623), .ZN(n9818) );
  NOR2_X1 U8783 ( .A1(n7102), .A2(n9818), .ZN(n7103) );
  OR2_X1 U8784 ( .A1(n7138), .A2(n7103), .ZN(n9820) );
  INV_X1 U8785 ( .A(n9762), .ZN(n9291) );
  AOI22_X1 U8786 ( .A1(n9291), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7231), .B2(
        n9747), .ZN(n7105) );
  NAND2_X1 U8787 ( .A1(n9226), .A2(n8623), .ZN(n7104) );
  OAI211_X1 U8788 ( .C1(n9820), .C2(n9042), .A(n7105), .B(n7104), .ZN(n7106)
         );
  AOI21_X1 U8789 ( .B1(n9823), .B2(n9719), .A(n7106), .ZN(n7107) );
  OAI21_X1 U8790 ( .B1(n9825), .B2(n9234), .A(n7107), .ZN(P1_U3282) );
  NAND2_X1 U8791 ( .A1(n7109), .A2(n7108), .ZN(n7110) );
  XOR2_X1 U8792 ( .A(n7111), .B(n7110), .Z(n7118) );
  OR2_X1 U8793 ( .A1(n7162), .A2(n9863), .ZN(n7113) );
  OR2_X1 U8794 ( .A1(n7368), .A2(n9861), .ZN(n7112) );
  AND2_X1 U8795 ( .A1(n7113), .A2(n7112), .ZN(n7168) );
  INV_X1 U8796 ( .A(n7168), .ZN(n7114) );
  AOI22_X1 U8797 ( .A1(n7890), .A2(n7114), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n7116) );
  NAND2_X1 U8798 ( .A1(n7929), .A2(n9976), .ZN(n7115) );
  OAI211_X1 U8799 ( .C1(n7925), .C2(n7169), .A(n7116), .B(n7115), .ZN(n7117)
         );
  AOI21_X1 U8800 ( .B1(n7118), .B2(n7933), .A(n7117), .ZN(n7119) );
  INV_X1 U8801 ( .A(n7119), .ZN(P2_U3219) );
  OR2_X1 U8802 ( .A1(n8623), .A2(n7339), .ZN(n8806) );
  NAND2_X1 U8803 ( .A1(n7120), .A2(n8806), .ZN(n7186) );
  NAND2_X1 U8804 ( .A1(n8623), .A2(n7339), .ZN(n8621) );
  NAND2_X1 U8805 ( .A1(n7186), .A2(n8621), .ZN(n7122) );
  OR2_X1 U8806 ( .A1(n7121), .A2(n7187), .ZN(n8633) );
  NAND2_X1 U8807 ( .A1(n7121), .A2(n7187), .ZN(n8634) );
  XNOR2_X1 U8808 ( .A(n7122), .B(n8736), .ZN(n7123) );
  AOI222_X1 U8809 ( .A1(n9727), .A2(n7123), .B1(n8891), .B2(n9756), .C1(n8893), 
        .C2(n9739), .ZN(n7255) );
  AND2_X1 U8810 ( .A1(n7125), .A2(n7124), .ZN(n7127) );
  NAND2_X1 U8811 ( .A1(n7128), .A2(n7127), .ZN(n7126) );
  AND2_X1 U8812 ( .A1(n7126), .A2(n7129), .ZN(n7134) );
  AND2_X1 U8813 ( .A1(n7127), .A2(n7130), .ZN(n7180) );
  NAND2_X1 U8814 ( .A1(n7128), .A2(n7180), .ZN(n7132) );
  NAND2_X1 U8815 ( .A1(n7132), .A2(n7177), .ZN(n7133) );
  AOI21_X1 U8816 ( .B1(n8736), .B2(n7134), .A(n7133), .ZN(n7256) );
  INV_X1 U8817 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7136) );
  INV_X1 U8818 ( .A(n7341), .ZN(n7135) );
  OAI22_X1 U8819 ( .A1(n9762), .A2(n7136), .B1(n7135), .B2(n9222), .ZN(n7137)
         );
  AOI21_X1 U8820 ( .B1(n9226), .B2(n7121), .A(n7137), .ZN(n7141) );
  INV_X1 U8821 ( .A(n7121), .ZN(n7344) );
  NAND2_X1 U8822 ( .A1(n7138), .A2(n7344), .ZN(n7191) );
  OR2_X1 U8823 ( .A1(n7138), .A2(n7344), .ZN(n7139) );
  AND3_X1 U8824 ( .A1(n7191), .A2(n7139), .A3(n9742), .ZN(n7253) );
  NAND2_X1 U8825 ( .A1(n7253), .A2(n9289), .ZN(n7140) );
  OAI211_X1 U8826 ( .C1(n7256), .C2(n9297), .A(n7141), .B(n7140), .ZN(n7142)
         );
  INV_X1 U8827 ( .A(n7142), .ZN(n7143) );
  OAI21_X1 U8828 ( .B1(n9291), .B2(n7255), .A(n7143), .ZN(P1_U3281) );
  NAND2_X1 U8829 ( .A1(n7145), .A2(n7144), .ZN(n7146) );
  XOR2_X1 U8830 ( .A(n7147), .B(n7146), .Z(n7156) );
  NAND2_X1 U8831 ( .A1(n8583), .A2(n7148), .ZN(n7151) );
  NOR2_X1 U8832 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7149), .ZN(n9660) );
  AOI21_X1 U8833 ( .B1(n8552), .B2(n8893), .A(n9660), .ZN(n7150) );
  OAI211_X1 U8834 ( .C1(n7152), .C2(n8573), .A(n7151), .B(n7150), .ZN(n7153)
         );
  AOI21_X1 U8835 ( .B1(n7154), .B2(n8590), .A(n7153), .ZN(n7155) );
  OAI21_X1 U8836 ( .B1(n7156), .B2(n8592), .A(n7155), .ZN(P1_U3219) );
  INV_X1 U8837 ( .A(n7157), .ZN(n7955) );
  NAND2_X1 U8838 ( .A1(n9969), .A2(n7955), .ZN(n7158) );
  INV_X1 U8839 ( .A(n7202), .ZN(n7161) );
  OR2_X1 U8840 ( .A1(n8434), .A2(n7162), .ZN(n7676) );
  NAND2_X1 U8841 ( .A1(n8434), .A2(n7162), .ZN(n7671) );
  NAND2_X1 U8842 ( .A1(n7161), .A2(n7160), .ZN(n7200) );
  INV_X1 U8843 ( .A(n7162), .ZN(n7954) );
  OR2_X1 U8844 ( .A1(n8434), .A2(n7954), .ZN(n7163) );
  NAND2_X1 U8845 ( .A1(n9976), .A2(n7203), .ZN(n7685) );
  NAND2_X1 U8846 ( .A1(n7364), .A2(n7778), .ZN(n7164) );
  NAND2_X1 U8847 ( .A1(n7345), .A2(n7164), .ZN(n9975) );
  NAND2_X1 U8848 ( .A1(n7165), .A2(n7669), .ZN(n7199) );
  OAI211_X1 U8849 ( .C1(n7166), .C2(n7778), .A(n9865), .B(n7366), .ZN(n7167)
         );
  OAI211_X1 U8850 ( .C1(n9975), .C2(n9854), .A(n7168), .B(n7167), .ZN(n9978)
         );
  NAND2_X1 U8851 ( .A1(n9978), .A2(n8336), .ZN(n7176) );
  OAI22_X1 U8852 ( .A1(n8336), .A2(n7170), .B1(n7169), .B2(n8272), .ZN(n7174)
         );
  AND2_X1 U8853 ( .A1(n7208), .A2(n9976), .ZN(n7172) );
  OR2_X1 U8854 ( .A1(n7172), .A2(n7349), .ZN(n9977) );
  NOR2_X1 U8855 ( .A1(n9977), .A2(n8278), .ZN(n7173) );
  AOI211_X1 U8856 ( .C1(n8324), .C2(n9976), .A(n7174), .B(n7173), .ZN(n7175)
         );
  OAI211_X1 U8857 ( .C1(n9975), .C2(n9876), .A(n7176), .B(n7175), .ZN(P2_U3286) );
  OR2_X1 U8858 ( .A1(n7121), .A2(n8892), .ZN(n7178) );
  AND2_X1 U8859 ( .A1(n7178), .A2(n7177), .ZN(n7182) );
  AND2_X1 U8860 ( .A1(n7179), .A2(n7182), .ZN(n7184) );
  INV_X1 U8861 ( .A(n7180), .ZN(n7181) );
  AND2_X1 U8862 ( .A1(n7193), .A2(n7418), .ZN(n7319) );
  INV_X1 U8863 ( .A(n7319), .ZN(n8637) );
  OR2_X1 U8864 ( .A1(n7193), .A2(n7418), .ZN(n7397) );
  XNOR2_X1 U8865 ( .A(n7327), .B(n8737), .ZN(n9602) );
  AND2_X1 U8866 ( .A1(n8634), .A2(n8621), .ZN(n8809) );
  INV_X1 U8867 ( .A(n8633), .ZN(n8807) );
  AOI21_X1 U8868 ( .B1(n7186), .B2(n8809), .A(n8807), .ZN(n7320) );
  XNOR2_X1 U8869 ( .A(n7320), .B(n8737), .ZN(n7189) );
  OAI22_X1 U8870 ( .A1(n7187), .A2(n9724), .B1(n9723), .B2(n7433), .ZN(n7188)
         );
  AOI21_X1 U8871 ( .B1(n7189), .B2(n9727), .A(n7188), .ZN(n7190) );
  OAI21_X1 U8872 ( .B1(n9602), .B2(n9759), .A(n7190), .ZN(n9605) );
  NAND2_X1 U8873 ( .A1(n9605), .A2(n9762), .ZN(n7198) );
  NAND2_X1 U8874 ( .A1(n7191), .A2(n7193), .ZN(n7192) );
  NAND2_X1 U8875 ( .A1(n7324), .A2(n7192), .ZN(n9604) );
  INV_X1 U8876 ( .A(n9604), .ZN(n7196) );
  INV_X1 U8877 ( .A(n7193), .ZN(n9603) );
  AOI22_X1 U8878 ( .A1(n9291), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7384), .B2(
        n9747), .ZN(n7194) );
  OAI21_X1 U8879 ( .B1(n9603), .B2(n9733), .A(n7194), .ZN(n7195) );
  AOI21_X1 U8880 ( .B1(n7196), .B2(n9718), .A(n7195), .ZN(n7197) );
  OAI211_X1 U8881 ( .C1(n9602), .C2(n9276), .A(n7198), .B(n7197), .ZN(P1_U3280) );
  XNOR2_X1 U8882 ( .A(n7199), .B(n7777), .ZN(n7206) );
  INV_X1 U8883 ( .A(n7200), .ZN(n7201) );
  AOI21_X1 U8884 ( .B1(n7777), .B2(n7202), .A(n7201), .ZN(n8438) );
  INV_X1 U8885 ( .A(n7203), .ZN(n7953) );
  AOI22_X1 U8886 ( .A1(n8312), .A2(n7955), .B1(n7953), .B2(n8313), .ZN(n7204)
         );
  OAI21_X1 U8887 ( .B1(n8438), .B2(n9854), .A(n7204), .ZN(n7205) );
  AOI21_X1 U8888 ( .B1(n7206), .B2(n9865), .A(n7205), .ZN(n8437) );
  NAND2_X1 U8889 ( .A1(n4420), .A2(n8434), .ZN(n7207) );
  AND2_X1 U8890 ( .A1(n7208), .A2(n7207), .ZN(n8435) );
  OAI22_X1 U8891 ( .A1(n8336), .A2(n7210), .B1(n7209), .B2(n8272), .ZN(n7212)
         );
  NOR2_X1 U8892 ( .A1(n8307), .A2(n7171), .ZN(n7211) );
  AOI211_X1 U8893 ( .C1(n8435), .C2(n8319), .A(n7212), .B(n7211), .ZN(n7214)
         );
  OR2_X1 U8894 ( .A1(n8438), .A2(n9876), .ZN(n7213) );
  OAI211_X1 U8895 ( .C1(n8437), .C2(n4247), .A(n7214), .B(n7213), .ZN(P2_U3287) );
  INV_X1 U8896 ( .A(n7449), .ZN(n9984) );
  OAI21_X1 U8897 ( .B1(n7217), .B2(n7216), .A(n7215), .ZN(n7218) );
  NAND2_X1 U8898 ( .A1(n7218), .A2(n7933), .ZN(n7223) );
  INV_X1 U8899 ( .A(n7219), .ZN(n7371) );
  OAI22_X1 U8900 ( .A1(n7693), .A2(n7939), .B1(n7938), .B2(n7368), .ZN(n7220)
         );
  AOI211_X1 U8901 ( .C1(n7371), .C2(n7942), .A(n7221), .B(n7220), .ZN(n7222)
         );
  OAI211_X1 U8902 ( .C1(n9984), .C2(n7945), .A(n7223), .B(n7222), .ZN(P2_U3226) );
  INV_X1 U8903 ( .A(n7241), .ZN(n7226) );
  AOI21_X1 U8904 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8461), .A(n7224), .ZN(
        n7225) );
  OAI21_X1 U8905 ( .B1(n7226), .B2(n8467), .A(n7225), .ZN(P2_U3335) );
  INV_X1 U8906 ( .A(n7228), .ZN(n7229) );
  AOI21_X1 U8907 ( .B1(n7230), .B2(n7227), .A(n7229), .ZN(n7238) );
  NAND2_X1 U8908 ( .A1(n8583), .A2(n7231), .ZN(n7234) );
  AOI21_X1 U8909 ( .B1(n8552), .B2(n8892), .A(n7232), .ZN(n7233) );
  OAI211_X1 U8910 ( .C1(n7235), .C2(n8573), .A(n7234), .B(n7233), .ZN(n7236)
         );
  AOI21_X1 U8911 ( .B1(n8623), .B2(n8590), .A(n7236), .ZN(n7237) );
  OAI21_X1 U8912 ( .B1(n7238), .B2(n8592), .A(n7237), .ZN(P1_U3229) );
  INV_X1 U8913 ( .A(n7239), .ZN(n7594) );
  OAI222_X1 U8914 ( .A1(n7852), .A2(n7240), .B1(n4249), .B2(n7594), .C1(n5639), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  NAND2_X1 U8915 ( .A1(n7241), .A2(n7567), .ZN(n7243) );
  OR2_X1 U8916 ( .A1(n7242), .A2(P1_U3084), .ZN(n8839) );
  OAI211_X1 U8917 ( .C1(n7244), .C2(n7852), .A(n7243), .B(n8839), .ZN(P1_U3330) );
  XNOR2_X1 U8918 ( .A(n7246), .B(n7245), .ZN(n7252) );
  INV_X1 U8919 ( .A(n7247), .ZN(n7459) );
  OAI22_X1 U8920 ( .A1(n7517), .A2(n7939), .B1(n7938), .B2(n7365), .ZN(n7248)
         );
  AOI211_X1 U8921 ( .C1(n7942), .C2(n7459), .A(n7249), .B(n7248), .ZN(n7251)
         );
  NAND2_X1 U8922 ( .A1(n8424), .A2(n7929), .ZN(n7250) );
  OAI211_X1 U8923 ( .C1(n7252), .C2(n7931), .A(n7251), .B(n7250), .ZN(P2_U3236) );
  INV_X1 U8924 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7258) );
  AOI21_X1 U8925 ( .B1(n9598), .B2(n7121), .A(n7253), .ZN(n7254) );
  OAI211_X1 U8926 ( .C1(n7256), .C2(n9524), .A(n7255), .B(n7254), .ZN(n7259)
         );
  NAND2_X1 U8927 ( .A1(n7259), .A2(n9828), .ZN(n7257) );
  OAI21_X1 U8928 ( .B1(n9828), .B2(n7258), .A(n7257), .ZN(P1_U3484) );
  NAND2_X1 U8929 ( .A1(n7259), .A2(n9843), .ZN(n7260) );
  OAI21_X1 U8930 ( .B1(n9843), .B2(n6496), .A(n7260), .ZN(P1_U3533) );
  INV_X1 U8931 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7273) );
  OAI21_X1 U8932 ( .B1(n7266), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7261), .ZN(
        n7264) );
  NOR2_X1 U8933 ( .A1(n7507), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7262) );
  AOI21_X1 U8934 ( .B1(n7507), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7262), .ZN(
        n7263) );
  NAND2_X1 U8935 ( .A1(n7263), .A2(n7264), .ZN(n7506) );
  OAI21_X1 U8936 ( .B1(n7264), .B2(n7263), .A(n7506), .ZN(n7271) );
  NAND2_X1 U8937 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8474) );
  OAI21_X1 U8938 ( .B1(n9687), .B2(n7498), .A(n8474), .ZN(n7270) );
  XNOR2_X1 U8939 ( .A(n7498), .B(n7499), .ZN(n7268) );
  INV_X1 U8940 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7267) );
  NOR2_X1 U8941 ( .A1(n7267), .A2(n7268), .ZN(n7500) );
  AOI211_X1 U8942 ( .C1(n7268), .C2(n7267), .A(n7500), .B(n9679), .ZN(n7269)
         );
  AOI211_X1 U8943 ( .C1(n9707), .C2(n7271), .A(n7270), .B(n7269), .ZN(n7272)
         );
  OAI21_X1 U8944 ( .B1(n9689), .B2(n7273), .A(n7272), .ZN(P1_U3255) );
  NAND2_X1 U8945 ( .A1(n7275), .A2(n7274), .ZN(n7276) );
  NOR2_X1 U8946 ( .A1(n7276), .A2(n7285), .ZN(n8066) );
  AOI21_X1 U8947 ( .B1(n7276), .B2(n7285), .A(n8066), .ZN(n7277) );
  INV_X1 U8948 ( .A(n7277), .ZN(n7278) );
  NOR2_X1 U8949 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n7278), .ZN(n8065) );
  AOI21_X1 U8950 ( .B1(n7278), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8065), .ZN(
        n7287) );
  AOI21_X1 U8951 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n7280), .A(n7279), .ZN(
        n8070) );
  XOR2_X1 U8952 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n7285), .Z(n8071) );
  XOR2_X1 U8953 ( .A(n8070), .B(n8071), .Z(n7282) );
  NAND2_X1 U8954 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7924) );
  NAND2_X1 U8955 ( .A1(n9850), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n7281) );
  OAI211_X1 U8956 ( .C1(n7283), .C2(n7282), .A(n7924), .B(n7281), .ZN(n7284)
         );
  AOI21_X1 U8957 ( .B1(n7285), .B2(n9556), .A(n7284), .ZN(n7286) );
  OAI21_X1 U8958 ( .B1(n7287), .B2(n9848), .A(n7286), .ZN(P2_U3263) );
  INV_X1 U8959 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10044) );
  NOR2_X1 U8960 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(P2_ADDR_REG_17__SCAN_IN), 
        .ZN(n7288) );
  AOI21_X1 U8961 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n7288), .ZN(n10015) );
  NOR2_X1 U8962 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7289) );
  AOI21_X1 U8963 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7289), .ZN(n10018) );
  NOR2_X1 U8964 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7290) );
  AOI21_X1 U8965 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7290), .ZN(n10021) );
  NOR2_X1 U8966 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7291) );
  AOI21_X1 U8967 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7291), .ZN(n10024) );
  NOR2_X1 U8968 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7292) );
  AOI21_X1 U8969 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7292), .ZN(n10027) );
  NOR2_X1 U8970 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7299) );
  XNOR2_X1 U8971 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10057) );
  NAND2_X1 U8972 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7297) );
  XOR2_X1 U8973 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10055) );
  NAND2_X1 U8974 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7295) );
  XOR2_X1 U8975 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10053) );
  AOI21_X1 U8976 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10009) );
  INV_X1 U8977 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7293) );
  NAND3_X1 U8978 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10011) );
  OAI21_X1 U8979 ( .B1(n10009), .B2(n7293), .A(n10011), .ZN(n10052) );
  NAND2_X1 U8980 ( .A1(n10053), .A2(n10052), .ZN(n7294) );
  NAND2_X1 U8981 ( .A1(n7295), .A2(n7294), .ZN(n10054) );
  NAND2_X1 U8982 ( .A1(n10055), .A2(n10054), .ZN(n7296) );
  NAND2_X1 U8983 ( .A1(n7297), .A2(n7296), .ZN(n10056) );
  NOR2_X1 U8984 ( .A1(n10057), .A2(n10056), .ZN(n7298) );
  NOR2_X1 U8985 ( .A1(n7299), .A2(n7298), .ZN(n7300) );
  NOR2_X1 U8986 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7300), .ZN(n10039) );
  AND2_X1 U8987 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7300), .ZN(n10038) );
  NOR2_X1 U8988 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10038), .ZN(n7301) );
  NOR2_X1 U8989 ( .A1(n10039), .A2(n7301), .ZN(n7302) );
  NAND2_X1 U8990 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n7302), .ZN(n7304) );
  XNOR2_X1 U8991 ( .A(n7302), .B(n9395), .ZN(n10037) );
  NAND2_X1 U8992 ( .A1(n10037), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7303) );
  NAND2_X1 U8993 ( .A1(n7304), .A2(n7303), .ZN(n7305) );
  NAND2_X1 U8994 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7305), .ZN(n7307) );
  XOR2_X1 U8995 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7305), .Z(n10041) );
  NAND2_X1 U8996 ( .A1(n10041), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7306) );
  NAND2_X1 U8997 ( .A1(n7307), .A2(n7306), .ZN(n7308) );
  AND2_X1 U8998 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7308), .ZN(n7309) );
  INV_X1 U8999 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10051) );
  XNOR2_X1 U9000 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7308), .ZN(n10050) );
  INV_X1 U9001 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7311) );
  NOR2_X1 U9002 ( .A1(n7310), .A2(n7311), .ZN(n7312) );
  XNOR2_X1 U9003 ( .A(n7311), .B(n7310), .ZN(n10047) );
  NOR2_X1 U9004 ( .A1(n10048), .A2(n10047), .ZN(n10046) );
  NOR2_X1 U9005 ( .A1(n7312), .A2(n10046), .ZN(n10036) );
  NAND2_X1 U9006 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7313) );
  OAI21_X1 U9007 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7313), .ZN(n10035) );
  NOR2_X1 U9008 ( .A1(n10036), .A2(n10035), .ZN(n10034) );
  AOI21_X1 U9009 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10034), .ZN(n10033) );
  NAND2_X1 U9010 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7314) );
  OAI21_X1 U9011 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7314), .ZN(n10032) );
  NOR2_X1 U9012 ( .A1(n10033), .A2(n10032), .ZN(n10031) );
  AOI21_X1 U9013 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10031), .ZN(n10030) );
  NOR2_X1 U9014 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7315) );
  AOI21_X1 U9015 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7315), .ZN(n10029) );
  NAND2_X1 U9016 ( .A1(n10030), .A2(n10029), .ZN(n10028) );
  OAI21_X1 U9017 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10028), .ZN(n10026) );
  NAND2_X1 U9018 ( .A1(n10027), .A2(n10026), .ZN(n10025) );
  OAI21_X1 U9019 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10025), .ZN(n10023) );
  NAND2_X1 U9020 ( .A1(n10024), .A2(n10023), .ZN(n10022) );
  OAI21_X1 U9021 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10022), .ZN(n10020) );
  NAND2_X1 U9022 ( .A1(n10021), .A2(n10020), .ZN(n10019) );
  OAI21_X1 U9023 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10019), .ZN(n10017) );
  NAND2_X1 U9024 ( .A1(n10018), .A2(n10017), .ZN(n10016) );
  OAI21_X1 U9025 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10016), .ZN(n10014) );
  NAND2_X1 U9026 ( .A1(n10015), .A2(n10014), .ZN(n10013) );
  OAI21_X1 U9027 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10013), .ZN(n10043) );
  NOR2_X1 U9028 ( .A1(n10044), .A2(n10043), .ZN(n7316) );
  NAND2_X1 U9029 ( .A1(n10044), .A2(n10043), .ZN(n10042) );
  OAI21_X1 U9030 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7316), .A(n10042), .ZN(
        n7318) );
  XNOR2_X1 U9031 ( .A(n4720), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7317) );
  XNOR2_X1 U9032 ( .A(n7318), .B(n7317), .ZN(ADD_1071_U4) );
  OR2_X1 U9033 ( .A1(n9597), .A2(n7433), .ZN(n8640) );
  NAND2_X1 U9034 ( .A1(n9597), .A2(n7433), .ZN(n8811) );
  INV_X1 U9035 ( .A(n7397), .ZN(n7321) );
  NOR2_X1 U9036 ( .A1(n7398), .A2(n7321), .ZN(n7322) );
  XOR2_X1 U9037 ( .A(n8738), .B(n7322), .Z(n7323) );
  OAI222_X1 U9038 ( .A1(n9723), .A2(n9284), .B1(n9724), .B2(n7418), .C1(n9751), 
        .C2(n7323), .ZN(n9595) );
  INV_X1 U9039 ( .A(n9595), .ZN(n7332) );
  AOI211_X1 U9040 ( .C1(n9597), .C2(n7324), .A(n9819), .B(n7404), .ZN(n9596)
         );
  INV_X1 U9041 ( .A(n9597), .ZN(n7423) );
  AOI22_X1 U9042 ( .A1(n9291), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7420), .B2(
        n9747), .ZN(n7325) );
  OAI21_X1 U9043 ( .B1(n7423), .B2(n9733), .A(n7325), .ZN(n7326) );
  AOI21_X1 U9044 ( .B1(n9596), .B2(n9289), .A(n7326), .ZN(n7331) );
  INV_X1 U9045 ( .A(n8738), .ZN(n7328) );
  NAND2_X1 U9046 ( .A1(n7329), .A2(n8738), .ZN(n9599) );
  NAND3_X1 U9047 ( .A1(n7394), .A2(n9599), .A3(n9220), .ZN(n7330) );
  OAI211_X1 U9048 ( .C1(n7332), .C2(n9234), .A(n7331), .B(n7330), .ZN(P1_U3279) );
  OAI21_X1 U9049 ( .B1(n7335), .B2(n7333), .A(n7334), .ZN(n7336) );
  NAND2_X1 U9050 ( .A1(n7336), .A2(n8571), .ZN(n7343) );
  NOR2_X1 U9051 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7337), .ZN(n9684) );
  AOI21_X1 U9052 ( .B1(n8552), .B2(n8891), .A(n9684), .ZN(n7338) );
  OAI21_X1 U9053 ( .B1(n8573), .B2(n7339), .A(n7338), .ZN(n7340) );
  AOI21_X1 U9054 ( .B1(n7341), .B2(n8583), .A(n7340), .ZN(n7342) );
  OAI211_X1 U9055 ( .C1(n7344), .C2(n8578), .A(n7343), .B(n7342), .ZN(P1_U3215) );
  NAND2_X1 U9056 ( .A1(n9976), .A2(n7953), .ZN(n7359) );
  NAND2_X1 U9057 ( .A1(n7345), .A2(n7359), .ZN(n7346) );
  NAND2_X1 U9058 ( .A1(n8429), .A2(n7368), .ZN(n7684) );
  NAND2_X1 U9059 ( .A1(n7690), .A2(n7684), .ZN(n7781) );
  XNOR2_X1 U9060 ( .A(n7346), .B(n7781), .ZN(n8433) );
  NAND2_X1 U9061 ( .A1(n7366), .A2(n7675), .ZN(n7347) );
  XNOR2_X1 U9062 ( .A(n7347), .B(n7781), .ZN(n7348) );
  INV_X1 U9063 ( .A(n7365), .ZN(n7952) );
  AOI222_X1 U9064 ( .A1(n9865), .A2(n7348), .B1(n7952), .B2(n8313), .C1(n7953), 
        .C2(n8312), .ZN(n8432) );
  OR2_X1 U9065 ( .A1(n8432), .A2(n4247), .ZN(n7356) );
  INV_X1 U9066 ( .A(n7349), .ZN(n7350) );
  AOI21_X1 U9067 ( .B1(n8429), .B2(n7350), .A(n7369), .ZN(n8430) );
  NOR2_X1 U9068 ( .A1(n8307), .A2(n4705), .ZN(n7354) );
  OAI22_X1 U9069 ( .A1(n8336), .A2(n7352), .B1(n7351), .B2(n8272), .ZN(n7353)
         );
  AOI211_X1 U9070 ( .C1(n8430), .C2(n8319), .A(n7354), .B(n7353), .ZN(n7355)
         );
  OAI211_X1 U9071 ( .C1(n8433), .C2(n8321), .A(n7356), .B(n7355), .ZN(P2_U3285) );
  NAND2_X1 U9072 ( .A1(n8429), .A2(n4704), .ZN(n7358) );
  INV_X1 U9073 ( .A(n7358), .ZN(n7357) );
  NOR2_X1 U9074 ( .A1(n7357), .A2(n7781), .ZN(n7361) );
  OR2_X1 U9075 ( .A1(n7778), .A2(n7361), .ZN(n7363) );
  AND2_X1 U9076 ( .A1(n7359), .A2(n7358), .ZN(n7360) );
  OR2_X1 U9077 ( .A1(n7361), .A2(n7360), .ZN(n7362) );
  OR2_X1 U9078 ( .A1(n7449), .A2(n7365), .ZN(n7688) );
  NAND2_X1 U9079 ( .A1(n7449), .A2(n7365), .ZN(n7683) );
  XNOR2_X1 U9080 ( .A(n7450), .B(n7686), .ZN(n9990) );
  INV_X1 U9081 ( .A(n9990), .ZN(n7376) );
  INV_X1 U9082 ( .A(n7686), .ZN(n7782) );
  XNOR2_X1 U9083 ( .A(n7447), .B(n7782), .ZN(n7367) );
  OAI222_X1 U9084 ( .A1(n9861), .A2(n7693), .B1(n9863), .B2(n7368), .C1(n7367), 
        .C2(n8292), .ZN(n9987) );
  NOR2_X1 U9085 ( .A1(n7369), .A2(n9984), .ZN(n7370) );
  OR2_X1 U9086 ( .A1(n7457), .A2(n7370), .ZN(n9986) );
  AOI22_X1 U9087 ( .A1(n4247), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7371), .B2(
        n9869), .ZN(n7373) );
  NAND2_X1 U9088 ( .A1(n8324), .A2(n7449), .ZN(n7372) );
  OAI211_X1 U9089 ( .C1(n9986), .C2(n8278), .A(n7373), .B(n7372), .ZN(n7374)
         );
  AOI21_X1 U9090 ( .B1(n9987), .B2(n8336), .A(n7374), .ZN(n7375) );
  OAI21_X1 U9091 ( .B1(n8321), .B2(n7376), .A(n7375), .ZN(P2_U3284) );
  AND2_X1 U9092 ( .A1(n7334), .A2(n7377), .ZN(n7380) );
  OAI211_X1 U9093 ( .C1(n7380), .C2(n7379), .A(n8571), .B(n7378), .ZN(n7386)
         );
  AOI21_X1 U9094 ( .B1(n8585), .B2(n8892), .A(n7381), .ZN(n7382) );
  OAI21_X1 U9095 ( .B1(n8588), .B2(n7433), .A(n7382), .ZN(n7383) );
  AOI21_X1 U9096 ( .B1(n7384), .B2(n8583), .A(n7383), .ZN(n7385) );
  OAI211_X1 U9097 ( .C1(n9603), .C2(n8578), .A(n7386), .B(n7385), .ZN(P1_U3234) );
  INV_X1 U9098 ( .A(n7387), .ZN(n7391) );
  OAI222_X1 U9099 ( .A1(P1_U3084), .A2(n7389), .B1(n4249), .B2(n7391), .C1(
        n7388), .C2(n7852), .ZN(P1_U3329) );
  INV_X1 U9100 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7390) );
  OAI222_X1 U9101 ( .A1(P2_U3152), .A2(n7392), .B1(n8467), .B2(n7391), .C1(
        n7390), .C2(n8465), .ZN(P2_U3334) );
  NAND2_X1 U9102 ( .A1(n9597), .A2(n8890), .ZN(n7393) );
  NAND2_X1 U9103 ( .A1(n7394), .A2(n7393), .ZN(n7395) );
  OR2_X1 U9104 ( .A1(n7435), .A2(n9284), .ZN(n8639) );
  NAND2_X1 U9105 ( .A1(n7435), .A2(n9284), .ZN(n9009) );
  NAND2_X1 U9106 ( .A1(n8639), .A2(n9009), .ZN(n8740) );
  NAND2_X1 U9107 ( .A1(n7395), .A2(n8740), .ZN(n8984) );
  OR2_X1 U9108 ( .A1(n7395), .A2(n8740), .ZN(n7396) );
  NAND2_X1 U9109 ( .A1(n8984), .A2(n7396), .ZN(n9588) );
  INV_X1 U9110 ( .A(n8740), .ZN(n7400) );
  NAND2_X1 U9111 ( .A1(n8640), .A2(n7397), .ZN(n8810) );
  OAI21_X1 U9112 ( .B1(n7398), .B2(n8810), .A(n8811), .ZN(n7399) );
  NAND2_X1 U9113 ( .A1(n7399), .A2(n7400), .ZN(n9010) );
  OAI21_X1 U9114 ( .B1(n7400), .B2(n7399), .A(n9010), .ZN(n7402) );
  OAI22_X1 U9115 ( .A1(n7433), .A2(n9724), .B1(n9723), .B2(n8985), .ZN(n7401)
         );
  AOI21_X1 U9116 ( .B1(n7402), .B2(n9727), .A(n7401), .ZN(n7403) );
  OAI21_X1 U9117 ( .B1(n9588), .B2(n9759), .A(n7403), .ZN(n9591) );
  NAND2_X1 U9118 ( .A1(n9591), .A2(n9762), .ZN(n7410) );
  NOR2_X1 U9119 ( .A1(n7404), .A2(n9589), .ZN(n7405) );
  OR2_X1 U9120 ( .A1(n9286), .A2(n7405), .ZN(n9590) );
  INV_X1 U9121 ( .A(n9590), .ZN(n7408) );
  AOI22_X1 U9122 ( .A1(n9291), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7429), .B2(
        n9747), .ZN(n7406) );
  OAI21_X1 U9123 ( .B1(n9589), .B2(n9733), .A(n7406), .ZN(n7407) );
  AOI21_X1 U9124 ( .B1(n7408), .B2(n9718), .A(n7407), .ZN(n7409) );
  OAI211_X1 U9125 ( .C1(n9588), .C2(n9276), .A(n7410), .B(n7409), .ZN(P1_U3278) );
  INV_X1 U9126 ( .A(n7411), .ZN(n7415) );
  AOI21_X1 U9127 ( .B1(n7378), .B2(n7413), .A(n7412), .ZN(n7414) );
  OAI21_X1 U9128 ( .B1(n7415), .B2(n7414), .A(n8571), .ZN(n7422) );
  NOR2_X1 U9129 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7416), .ZN(n8933) );
  AOI21_X1 U9130 ( .B1(n8552), .B2(n8889), .A(n8933), .ZN(n7417) );
  OAI21_X1 U9131 ( .B1(n8573), .B2(n7418), .A(n7417), .ZN(n7419) );
  AOI21_X1 U9132 ( .B1(n7420), .B2(n8583), .A(n7419), .ZN(n7421) );
  OAI211_X1 U9133 ( .C1(n7423), .C2(n8578), .A(n7422), .B(n7421), .ZN(P1_U3222) );
  INV_X1 U9134 ( .A(n7424), .ZN(n7426) );
  NAND2_X1 U9135 ( .A1(n7426), .A2(n7425), .ZN(n7427) );
  XNOR2_X1 U9136 ( .A(n7428), .B(n7427), .ZN(n7437) );
  NAND2_X1 U9137 ( .A1(n8583), .A2(n7429), .ZN(n7432) );
  AOI21_X1 U9138 ( .B1(n8552), .B2(n9266), .A(n7430), .ZN(n7431) );
  OAI211_X1 U9139 ( .C1(n7433), .C2(n8573), .A(n7432), .B(n7431), .ZN(n7434)
         );
  AOI21_X1 U9140 ( .B1(n7435), .B2(n8590), .A(n7434), .ZN(n7436) );
  OAI21_X1 U9141 ( .B1(n7437), .B2(n8592), .A(n7436), .ZN(P1_U3232) );
  INV_X1 U9142 ( .A(n7438), .ZN(n7439) );
  AOI21_X1 U9143 ( .B1(n7441), .B2(n7440), .A(n7439), .ZN(n7446) );
  OAI21_X1 U9144 ( .B1(n7925), .B2(n7470), .A(n7442), .ZN(n7444) );
  OAI22_X1 U9145 ( .A1(n7525), .A2(n7939), .B1(n7938), .B2(n7693), .ZN(n7443)
         );
  AOI211_X1 U9146 ( .C1(n7488), .C2(n7929), .A(n7444), .B(n7443), .ZN(n7445)
         );
  OAI21_X1 U9147 ( .B1(n7446), .B2(n7931), .A(n7445), .ZN(P2_U3217) );
  NAND2_X1 U9148 ( .A1(n7447), .A2(n7688), .ZN(n7448) );
  NAND2_X1 U9149 ( .A1(n7448), .A2(n7683), .ZN(n7466) );
  XNOR2_X1 U9150 ( .A(n8424), .B(n7951), .ZN(n7784) );
  XNOR2_X1 U9151 ( .A(n7466), .B(n7784), .ZN(n7456) );
  INV_X1 U9152 ( .A(n7784), .ZN(n7451) );
  NAND2_X1 U9153 ( .A1(n7452), .A2(n7784), .ZN(n7453) );
  NAND2_X1 U9154 ( .A1(n7465), .A2(n7453), .ZN(n8428) );
  INV_X1 U9155 ( .A(n7517), .ZN(n7950) );
  AOI22_X1 U9156 ( .A1(n8312), .A2(n7952), .B1(n7950), .B2(n8313), .ZN(n7454)
         );
  OAI21_X1 U9157 ( .B1(n8428), .B2(n9854), .A(n7454), .ZN(n7455) );
  AOI21_X1 U9158 ( .B1(n9865), .B2(n7456), .A(n7455), .ZN(n8427) );
  INV_X1 U9159 ( .A(n7457), .ZN(n7458) );
  INV_X1 U9160 ( .A(n8424), .ZN(n7464) );
  AOI21_X1 U9161 ( .B1(n8424), .B2(n7458), .A(n4320), .ZN(n8425) );
  AOI22_X1 U9162 ( .A1(n4247), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7459), .B2(
        n9869), .ZN(n7460) );
  OAI21_X1 U9163 ( .B1(n7464), .B2(n8307), .A(n7460), .ZN(n7462) );
  NOR2_X1 U9164 ( .A1(n8428), .A2(n9876), .ZN(n7461) );
  AOI211_X1 U9165 ( .C1(n8425), .C2(n8319), .A(n7462), .B(n7461), .ZN(n7463)
         );
  OAI21_X1 U9166 ( .B1(n4247), .B2(n8427), .A(n7463), .ZN(P2_U3283) );
  NAND2_X1 U9167 ( .A1(n7488), .A2(n7517), .ZN(n7700) );
  XNOR2_X1 U9168 ( .A(n7489), .B(n7697), .ZN(n9577) );
  INV_X1 U9169 ( .A(n9577), .ZN(n7476) );
  INV_X1 U9170 ( .A(n7697), .ZN(n7783) );
  OAI211_X1 U9171 ( .C1(n7467), .C2(n7697), .A(n9865), .B(n7484), .ZN(n7469)
         );
  INV_X1 U9172 ( .A(n7525), .ZN(n7949) );
  AOI22_X1 U9173 ( .A1(n7949), .A2(n8313), .B1(n8312), .B2(n7951), .ZN(n7468)
         );
  NAND2_X1 U9174 ( .A1(n7469), .A2(n7468), .ZN(n9575) );
  INV_X1 U9175 ( .A(n7488), .ZN(n9573) );
  OAI21_X1 U9176 ( .B1(n4320), .B2(n9573), .A(n7491), .ZN(n9574) );
  OAI22_X1 U9177 ( .A1(n8336), .A2(n7471), .B1(n7470), .B2(n8272), .ZN(n7472)
         );
  AOI21_X1 U9178 ( .B1(n7488), .B2(n8324), .A(n7472), .ZN(n7473) );
  OAI21_X1 U9179 ( .B1(n9574), .B2(n8278), .A(n7473), .ZN(n7474) );
  AOI21_X1 U9180 ( .B1(n9575), .B2(n8336), .A(n7474), .ZN(n7475) );
  OAI21_X1 U9181 ( .B1(n7476), .B2(n8321), .A(n7475), .ZN(P2_U3282) );
  INV_X1 U9182 ( .A(n7477), .ZN(n7482) );
  OAI222_X1 U9183 ( .A1(n8465), .A2(n7480), .B1(n8467), .B2(n7482), .C1(
        P2_U3152), .C2(n7478), .ZN(P2_U3333) );
  OAI222_X1 U9184 ( .A1(n7852), .A2(n7483), .B1(n4249), .B2(n7482), .C1(
        P1_U3084), .C2(n7481), .ZN(P1_U3328) );
  NAND2_X1 U9185 ( .A1(n8419), .A2(n7525), .ZN(n7705) );
  NAND2_X1 U9186 ( .A1(n7704), .A2(n7705), .ZN(n7701) );
  INV_X1 U9187 ( .A(n7701), .ZN(n7786) );
  OAI211_X1 U9188 ( .C1(n7485), .C2(n7786), .A(n7524), .B(n9865), .ZN(n7487)
         );
  INV_X1 U9189 ( .A(n7573), .ZN(n7948) );
  AOI22_X1 U9190 ( .A1(n8312), .A2(n7950), .B1(n7948), .B2(n8313), .ZN(n7486)
         );
  OAI22_X1 U9191 ( .A1(n7489), .A2(n7697), .B1(n7488), .B2(n7950), .ZN(n7490)
         );
  NAND2_X1 U9192 ( .A1(n7490), .A2(n7701), .ZN(n7528) );
  OAI21_X1 U9193 ( .B1(n7490), .B2(n7701), .A(n7528), .ZN(n8418) );
  NAND2_X1 U9194 ( .A1(n8418), .A2(n8325), .ZN(n7497) );
  AOI21_X1 U9195 ( .B1(n8419), .B2(n7491), .A(n4321), .ZN(n8420) );
  INV_X1 U9196 ( .A(n8419), .ZN(n7492) );
  NOR2_X1 U9197 ( .A1(n7492), .A2(n8307), .ZN(n7495) );
  INV_X1 U9198 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7493) );
  OAI22_X1 U9199 ( .A1(n8336), .A2(n7493), .B1(n7516), .B2(n8272), .ZN(n7494)
         );
  AOI211_X1 U9200 ( .C1(n8420), .C2(n8319), .A(n7495), .B(n7494), .ZN(n7496)
         );
  OAI211_X1 U9201 ( .C1(n4247), .C2(n8422), .A(n7497), .B(n7496), .ZN(P2_U3281) );
  INV_X1 U9202 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7513) );
  NOR2_X1 U9203 ( .A1(n7499), .A2(n7498), .ZN(n7501) );
  INV_X1 U9204 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7502) );
  AOI211_X1 U9205 ( .C1(n7503), .C2(n7502), .A(n7545), .B(n9679), .ZN(n7504)
         );
  INV_X1 U9206 ( .A(n7504), .ZN(n7512) );
  NOR2_X1 U9207 ( .A1(n7505), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8584) );
  OAI21_X1 U9208 ( .B1(n7507), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7506), .ZN(
        n7549) );
  XNOR2_X1 U9209 ( .A(n7550), .B(n7549), .ZN(n7508) );
  INV_X1 U9210 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9435) );
  NOR2_X1 U9211 ( .A1(n9435), .A2(n7508), .ZN(n7551) );
  INV_X1 U9212 ( .A(n9707), .ZN(n9648) );
  AOI211_X1 U9213 ( .C1(n7508), .C2(n9435), .A(n7551), .B(n9648), .ZN(n7509)
         );
  AOI211_X1 U9214 ( .C1(n7510), .C2(n9699), .A(n8584), .B(n7509), .ZN(n7511)
         );
  OAI211_X1 U9215 ( .C1(n9689), .C2(n7513), .A(n7512), .B(n7511), .ZN(P1_U3256) );
  XNOR2_X1 U9216 ( .A(n7514), .B(n7515), .ZN(n7523) );
  INV_X1 U9217 ( .A(n7516), .ZN(n7520) );
  OAI22_X1 U9218 ( .A1(n7573), .A2(n7939), .B1(n7938), .B2(n7517), .ZN(n7518)
         );
  AOI211_X1 U9219 ( .C1(n7942), .C2(n7520), .A(n7519), .B(n7518), .ZN(n7522)
         );
  NAND2_X1 U9220 ( .A1(n8419), .A2(n7929), .ZN(n7521) );
  OAI211_X1 U9221 ( .C1(n7523), .C2(n7931), .A(n7522), .B(n7521), .ZN(P2_U3243) );
  OR2_X1 U9222 ( .A1(n7591), .A2(n7573), .ZN(n7708) );
  NAND2_X1 U9223 ( .A1(n7591), .A2(n7573), .ZN(n7707) );
  NAND2_X1 U9224 ( .A1(n4274), .A2(n7787), .ZN(n7572) );
  OAI21_X1 U9225 ( .B1(n4274), .B2(n7787), .A(n7572), .ZN(n7526) );
  OAI22_X1 U9226 ( .A1(n7525), .A2(n9863), .B1(n7926), .B2(n9861), .ZN(n7586)
         );
  AOI21_X1 U9227 ( .B1(n7526), .B2(n9865), .A(n7586), .ZN(n8416) );
  AOI21_X1 U9228 ( .B1(n7787), .B2(n7529), .A(n7575), .ZN(n8415) );
  INV_X1 U9229 ( .A(n7591), .ZN(n8413) );
  OAI21_X1 U9230 ( .B1(n4321), .B2(n8413), .A(n9946), .ZN(n7530) );
  OR2_X1 U9231 ( .A1(n7530), .A2(n7576), .ZN(n8412) );
  OAI22_X1 U9232 ( .A1(n8336), .A2(n7531), .B1(n7589), .B2(n8272), .ZN(n7532)
         );
  AOI21_X1 U9233 ( .B1(n7591), .B2(n8324), .A(n7532), .ZN(n7533) );
  OAI21_X1 U9234 ( .B1(n8412), .B2(n8195), .A(n7533), .ZN(n7534) );
  AOI21_X1 U9235 ( .B1(n8415), .B2(n8325), .A(n7534), .ZN(n7535) );
  OAI21_X1 U9236 ( .B1(n4247), .B2(n8416), .A(n7535), .ZN(P2_U3280) );
  INV_X1 U9237 ( .A(n7536), .ZN(n7540) );
  OAI222_X1 U9238 ( .A1(P2_U3152), .A2(n7538), .B1(n8467), .B2(n7540), .C1(
        n7537), .C2(n8465), .ZN(P2_U3332) );
  OAI222_X1 U9239 ( .A1(P1_U3084), .A2(n7541), .B1(n4249), .B2(n7540), .C1(
        n7539), .C2(n7852), .ZN(P1_U3327) );
  NAND2_X1 U9240 ( .A1(n7561), .A2(n7567), .ZN(n7542) );
  OAI211_X1 U9241 ( .C1(n7852), .C2(n7543), .A(n7542), .B(n8966), .ZN(P1_U3326) );
  NOR2_X1 U9242 ( .A1(n7544), .A2(n7550), .ZN(n7546) );
  NAND2_X1 U9243 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n8944), .ZN(n7547) );
  OAI21_X1 U9244 ( .B1(n8944), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7547), .ZN(
        n7548) );
  AOI211_X1 U9245 ( .C1(n4314), .C2(n7548), .A(n8939), .B(n9679), .ZN(n7560)
         );
  NOR2_X1 U9246 ( .A1(n7550), .A2(n7549), .ZN(n7552) );
  NOR2_X1 U9247 ( .A1(n7552), .A2(n7551), .ZN(n7554) );
  XNOR2_X1 U9248 ( .A(n8944), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7553) );
  NOR2_X1 U9249 ( .A1(n7554), .A2(n7553), .ZN(n8943) );
  AOI211_X1 U9250 ( .C1(n7554), .C2(n7553), .A(n8943), .B(n9648), .ZN(n7559)
         );
  INV_X1 U9251 ( .A(n9689), .ZN(n9706) );
  NAND2_X1 U9252 ( .A1(n9706), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7556) );
  NAND2_X1 U9253 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n7555) );
  OAI211_X1 U9254 ( .C1(n9687), .C2(n7557), .A(n7556), .B(n7555), .ZN(n7558)
         );
  OR3_X1 U9255 ( .A1(n7560), .A2(n7559), .A3(n7558), .ZN(P1_U3257) );
  INV_X1 U9256 ( .A(n7561), .ZN(n7562) );
  OAI222_X1 U9257 ( .A1(n8465), .A2(n7563), .B1(n8467), .B2(n7562), .C1(n7844), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U9258 ( .A(n7568), .ZN(n7566) );
  AOI21_X1 U9259 ( .B1(n8461), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n7564), .ZN(
        n7565) );
  OAI21_X1 U9260 ( .B1(n7566), .B2(n8467), .A(n7565), .ZN(P2_U3330) );
  NAND2_X1 U9261 ( .A1(n7568), .A2(n7567), .ZN(n7570) );
  OAI211_X1 U9262 ( .C1(n7852), .C2(n7571), .A(n7570), .B(n7569), .ZN(P1_U3325) );
  NAND2_X1 U9263 ( .A1(n8093), .A2(n7926), .ZN(n7628) );
  NAND2_X1 U9264 ( .A1(n7804), .A2(n7628), .ZN(n7789) );
  XNOR2_X1 U9265 ( .A(n7803), .B(n7789), .ZN(n7574) );
  OAI22_X1 U9266 ( .A1(n8097), .A2(n9861), .B1(n7573), .B2(n9863), .ZN(n7889)
         );
  AOI21_X1 U9267 ( .B1(n7574), .B2(n9865), .A(n7889), .ZN(n8410) );
  OAI21_X1 U9268 ( .B1(n4319), .B2(n7789), .A(n8096), .ZN(n8409) );
  NAND2_X1 U9269 ( .A1(n7576), .A2(n8094), .ZN(n8303) );
  OAI211_X1 U9270 ( .C1(n7576), .C2(n8094), .A(n9946), .B(n8303), .ZN(n8407)
         );
  OAI22_X1 U9271 ( .A1(n8336), .A2(n7577), .B1(n7892), .B2(n8272), .ZN(n7578)
         );
  AOI21_X1 U9272 ( .B1(n8093), .B2(n8324), .A(n7578), .ZN(n7579) );
  OAI21_X1 U9273 ( .B1(n8407), .B2(n8195), .A(n7579), .ZN(n7580) );
  AOI21_X1 U9274 ( .B1(n8409), .B2(n8325), .A(n7580), .ZN(n7581) );
  OAI21_X1 U9275 ( .B1(n4247), .B2(n8410), .A(n7581), .ZN(P2_U3279) );
  INV_X1 U9276 ( .A(n7582), .ZN(n7583) );
  AOI21_X1 U9277 ( .B1(n7585), .B2(n7584), .A(n7583), .ZN(n7593) );
  NAND2_X1 U9278 ( .A1(n7890), .A2(n7586), .ZN(n7588) );
  OAI211_X1 U9279 ( .C1(n7925), .C2(n7589), .A(n7588), .B(n7587), .ZN(n7590)
         );
  AOI21_X1 U9280 ( .B1(n7591), .B2(n7929), .A(n7590), .ZN(n7592) );
  OAI21_X1 U9281 ( .B1(n7593), .B2(n7931), .A(n7592), .ZN(P2_U3228) );
  OAI222_X1 U9282 ( .A1(n8465), .A2(n7595), .B1(n8467), .B2(n7594), .C1(
        P2_U3152), .C2(n7052), .ZN(P2_U3336) );
  INV_X1 U9283 ( .A(SI_28_), .ZN(n7599) );
  NAND2_X1 U9284 ( .A1(n7600), .A2(n7599), .ZN(n7601) );
  INV_X1 U9285 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9436) );
  INV_X1 U9286 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8607) );
  MUX2_X1 U9287 ( .A(n9436), .B(n8607), .S(n7613), .Z(n7739) );
  INV_X1 U9288 ( .A(SI_29_), .ZN(n7603) );
  AND2_X1 U9289 ( .A1(n7739), .A2(n7603), .ZN(n7604) );
  INV_X1 U9290 ( .A(n7739), .ZN(n7605) );
  NAND2_X1 U9291 ( .A1(n7605), .A2(SI_29_), .ZN(n7606) );
  MUX2_X1 U9292 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7613), .Z(n7609) );
  INV_X1 U9293 ( .A(n8595), .ZN(n7851) );
  INV_X1 U9294 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9356) );
  OAI222_X1 U9295 ( .A1(P2_U3152), .A2(n7596), .B1(n8467), .B2(n7851), .C1(
        n9356), .C2(n8465), .ZN(P2_U3328) );
  INV_X1 U9296 ( .A(n7607), .ZN(n7608) );
  NAND2_X1 U9297 ( .A1(n7608), .A2(SI_30_), .ZN(n7612) );
  NAND2_X1 U9298 ( .A1(n7610), .A2(n7609), .ZN(n7611) );
  MUX2_X1 U9299 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7613), .Z(n7614) );
  XNOR2_X1 U9300 ( .A(n7614), .B(SI_31_), .ZN(n7615) );
  NAND2_X1 U9301 ( .A1(n9543), .A2(n7742), .ZN(n7618) );
  NAND2_X1 U9302 ( .A1(n7743), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7617) );
  INV_X1 U9303 ( .A(n8085), .ZN(n7625) );
  NAND2_X1 U9304 ( .A1(n8340), .A2(n7625), .ZN(n7836) );
  NAND2_X1 U9305 ( .A1(n8595), .A2(n7742), .ZN(n7620) );
  NAND2_X1 U9306 ( .A1(n7743), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7619) );
  INV_X1 U9307 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9579) );
  NAND2_X1 U9308 ( .A1(n7621), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7623) );
  INV_X1 U9309 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9572) );
  OR2_X1 U9310 ( .A1(n4903), .A2(n9572), .ZN(n7622) );
  OAI211_X1 U9311 ( .C1(n7624), .C2(n9579), .A(n7623), .B(n7622), .ZN(n8119)
         );
  INV_X1 U9312 ( .A(n8119), .ZN(n7749) );
  NOR2_X1 U9313 ( .A1(n8089), .A2(n7749), .ZN(n7830) );
  NAND2_X1 U9314 ( .A1(n7836), .A2(n7832), .ZN(n7795) );
  OR2_X1 U9315 ( .A1(n8340), .A2(n7625), .ZN(n7751) );
  NOR2_X1 U9316 ( .A1(n7839), .A2(n7827), .ZN(n7626) );
  AND2_X1 U9317 ( .A1(n7052), .A2(n7626), .ZN(n7754) );
  INV_X1 U9318 ( .A(n8169), .ZN(n7727) );
  NAND2_X1 U9319 ( .A1(n8366), .A2(n8210), .ZN(n7728) );
  NAND2_X1 U9320 ( .A1(n8371), .A2(n7946), .ZN(n7723) );
  AND2_X1 U9321 ( .A1(n7627), .A2(n8244), .ZN(n7815) );
  INV_X1 U9322 ( .A(n7815), .ZN(n8207) );
  NAND2_X1 U9323 ( .A1(n7723), .A2(n8207), .ZN(n7726) );
  XNOR2_X1 U9324 ( .A(n7627), .B(n7947), .ZN(n8218) );
  INV_X1 U9325 ( .A(n8260), .ZN(n7871) );
  INV_X1 U9326 ( .A(n7765), .ZN(n7810) );
  INV_X1 U9327 ( .A(n7804), .ZN(n7630) );
  NAND2_X1 U9328 ( .A1(n8402), .A2(n8097), .ZN(n7768) );
  NAND2_X1 U9329 ( .A1(n7768), .A2(n7628), .ZN(n7629) );
  MUX2_X1 U9330 ( .A(n7630), .B(n7629), .S(n7754), .Z(n7712) );
  AND2_X1 U9331 ( .A1(n7641), .A2(n7640), .ZN(n7631) );
  INV_X1 U9332 ( .A(n7648), .ZN(n7633) );
  NAND2_X1 U9333 ( .A1(n7633), .A2(n7632), .ZN(n7638) );
  NAND2_X1 U9334 ( .A1(n7635), .A2(n7634), .ZN(n7637) );
  INV_X1 U9335 ( .A(n7661), .ZN(n7636) );
  AOI21_X1 U9336 ( .B1(n7638), .B2(n7637), .A(n7636), .ZN(n7660) );
  NAND2_X1 U9337 ( .A1(n7640), .A2(n7639), .ZN(n7643) );
  NAND2_X1 U9338 ( .A1(n7662), .A2(n7641), .ZN(n7642) );
  AOI21_X1 U9339 ( .B1(n7648), .B2(n7643), .A(n7642), .ZN(n7650) );
  AND2_X1 U9340 ( .A1(n7651), .A2(n7799), .ZN(n7644) );
  OAI211_X1 U9341 ( .C1(n7645), .C2(n7644), .A(n6727), .B(n7655), .ZN(n7646)
         );
  NAND3_X1 U9342 ( .A1(n7646), .A2(n7653), .A3(n4465), .ZN(n7647) );
  NAND3_X1 U9343 ( .A1(n7648), .A2(n9857), .A3(n7647), .ZN(n7649) );
  OAI21_X1 U9344 ( .B1(n7650), .B2(n7754), .A(n7649), .ZN(n7658) );
  NAND2_X1 U9345 ( .A1(n6727), .A2(n7651), .ZN(n7652) );
  NAND3_X1 U9346 ( .A1(n7654), .A2(n7653), .A3(n7652), .ZN(n7656) );
  NAND3_X1 U9347 ( .A1(n7656), .A2(n7754), .A3(n7655), .ZN(n7657) );
  NAND2_X1 U9348 ( .A1(n7658), .A2(n7657), .ZN(n7659) );
  OAI21_X1 U9349 ( .B1(n7660), .B2(n4465), .A(n7659), .ZN(n7664) );
  MUX2_X1 U9350 ( .A(n7662), .B(n7661), .S(n4465), .Z(n7663) );
  MUX2_X1 U9351 ( .A(n7666), .B(n7665), .S(n4465), .Z(n7667) );
  MUX2_X1 U9352 ( .A(n7669), .B(n7668), .S(n4465), .Z(n7670) );
  NAND2_X1 U9353 ( .A1(n7778), .A2(n7777), .ZN(n7673) );
  NAND3_X1 U9354 ( .A1(n7675), .A2(n7754), .A3(n7676), .ZN(n7672) );
  NAND2_X1 U9355 ( .A1(n7673), .A2(n7672), .ZN(n7674) );
  INV_X1 U9356 ( .A(n7685), .ZN(n7677) );
  OAI211_X1 U9357 ( .C1(n7677), .C2(n7676), .A(n7690), .B(n7675), .ZN(n7678)
         );
  INV_X1 U9358 ( .A(n7678), .ZN(n7679) );
  NAND3_X1 U9359 ( .A1(n7687), .A2(n7686), .A3(n7679), .ZN(n7682) );
  NAND2_X1 U9360 ( .A1(n7683), .A2(n7684), .ZN(n7680) );
  NAND2_X1 U9361 ( .A1(n7680), .A2(n7688), .ZN(n7681) );
  NAND2_X1 U9362 ( .A1(n7682), .A2(n7681), .ZN(n7692) );
  INV_X1 U9363 ( .A(n7683), .ZN(n7691) );
  NAND4_X1 U9364 ( .A1(n7687), .A2(n7686), .A3(n7685), .A4(n7684), .ZN(n7689)
         );
  NAND2_X1 U9365 ( .A1(n7951), .A2(n7754), .ZN(n7695) );
  NAND2_X1 U9366 ( .A1(n7693), .A2(n4465), .ZN(n7694) );
  MUX2_X1 U9367 ( .A(n7695), .B(n7694), .S(n8424), .Z(n7696) );
  MUX2_X1 U9368 ( .A(n7700), .B(n7699), .S(n4465), .Z(n7702) );
  AOI21_X1 U9369 ( .B1(n7703), .B2(n7702), .A(n7701), .ZN(n7711) );
  MUX2_X1 U9370 ( .A(n7705), .B(n7704), .S(n4465), .Z(n7706) );
  NAND2_X1 U9371 ( .A1(n7787), .A2(n7706), .ZN(n7710) );
  INV_X1 U9372 ( .A(n7789), .ZN(n7802) );
  MUX2_X1 U9373 ( .A(n7708), .B(n7707), .S(n4465), .Z(n7709) );
  NAND2_X1 U9374 ( .A1(n7715), .A2(n7768), .ZN(n7713) );
  OR2_X1 U9375 ( .A1(n8399), .A2(n8268), .ZN(n7767) );
  NAND2_X1 U9376 ( .A1(n7713), .A2(n7767), .ZN(n7714) );
  NAND2_X1 U9377 ( .A1(n8399), .A2(n8268), .ZN(n7808) );
  INV_X1 U9378 ( .A(n7766), .ZN(n7809) );
  NAND2_X1 U9379 ( .A1(n7716), .A2(n7808), .ZN(n7717) );
  NAND2_X1 U9380 ( .A1(n8385), .A2(n8269), .ZN(n8241) );
  OR2_X1 U9381 ( .A1(n8385), .A2(n8269), .ZN(n7764) );
  NAND2_X1 U9382 ( .A1(n8380), .A2(n7872), .ZN(n7763) );
  AOI21_X1 U9383 ( .B1(n7718), .B2(n7763), .A(n4465), .ZN(n7719) );
  NAND3_X1 U9384 ( .A1(n7720), .A2(n7764), .A3(n7809), .ZN(n7721) );
  NAND3_X1 U9385 ( .A1(n7721), .A2(n7763), .A3(n8241), .ZN(n7722) );
  NAND3_X1 U9386 ( .A1(n7724), .A2(n7814), .A3(n7722), .ZN(n7725) );
  INV_X1 U9387 ( .A(n7627), .ZN(n8105) );
  NAND2_X1 U9388 ( .A1(n8181), .A2(n8108), .ZN(n7731) );
  NAND2_X1 U9389 ( .A1(n7731), .A2(n8171), .ZN(n7730) );
  NAND2_X1 U9390 ( .A1(n8362), .A2(n8157), .ZN(n7819) );
  INV_X1 U9391 ( .A(n8174), .ZN(n7817) );
  NAND2_X1 U9392 ( .A1(n7817), .A2(n7728), .ZN(n7729) );
  MUX2_X1 U9393 ( .A(n7730), .B(n7729), .S(n4465), .Z(n7733) );
  INV_X1 U9394 ( .A(n8155), .ZN(n7792) );
  MUX2_X1 U9395 ( .A(n7819), .B(n7731), .S(n4465), .Z(n7732) );
  OAI211_X1 U9396 ( .C1(n7734), .C2(n7733), .A(n7792), .B(n7732), .ZN(n7738)
         );
  OR2_X1 U9397 ( .A1(n8355), .A2(n8176), .ZN(n7825) );
  NAND2_X1 U9398 ( .A1(n8350), .A2(n8158), .ZN(n7762) );
  INV_X1 U9399 ( .A(n7762), .ZN(n7735) );
  AOI21_X1 U9400 ( .B1(n8176), .B2(n8355), .A(n7735), .ZN(n7736) );
  MUX2_X1 U9401 ( .A(n7825), .B(n7736), .S(n4465), .Z(n7737) );
  XNOR2_X1 U9402 ( .A(n7739), .B(SI_29_), .ZN(n7740) );
  NAND2_X1 U9403 ( .A1(n8606), .A2(n7742), .ZN(n7745) );
  NAND2_X1 U9404 ( .A1(n7616), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7744) );
  NAND2_X1 U9405 ( .A1(n8346), .A2(n8134), .ZN(n7828) );
  INV_X1 U9406 ( .A(n7747), .ZN(n7746) );
  MUX2_X1 U9407 ( .A(n7828), .B(n7747), .S(n4465), .Z(n7748) );
  NAND2_X1 U9408 ( .A1(n8089), .A2(n7749), .ZN(n7750) );
  NAND2_X1 U9409 ( .A1(n7751), .A2(n7750), .ZN(n7837) );
  INV_X1 U9410 ( .A(n7837), .ZN(n7752) );
  NAND2_X1 U9411 ( .A1(n7753), .A2(n7752), .ZN(n7756) );
  NAND2_X1 U9412 ( .A1(n7837), .A2(n7754), .ZN(n7755) );
  NAND3_X1 U9413 ( .A1(n4263), .A2(n7756), .A3(n7755), .ZN(n7759) );
  INV_X1 U9414 ( .A(n7836), .ZN(n7757) );
  NAND2_X1 U9415 ( .A1(n7757), .A2(n7754), .ZN(n7758) );
  NAND2_X1 U9416 ( .A1(n7759), .A2(n7758), .ZN(n7760) );
  NAND2_X1 U9417 ( .A1(n7826), .A2(n7762), .ZN(n8137) );
  INV_X1 U9418 ( .A(n8137), .ZN(n8133) );
  NAND2_X1 U9419 ( .A1(n7767), .A2(n7808), .ZN(n8290) );
  NOR4_X1 U9420 ( .A1(n8329), .A2(n7769), .A3(n6915), .A4(n4866), .ZN(n7771)
         );
  NAND3_X1 U9421 ( .A1(n7771), .A2(n7770), .A3(n9857), .ZN(n7775) );
  NOR4_X1 U9422 ( .A1(n7775), .A2(n7774), .A3(n7773), .A4(n7772), .ZN(n7779)
         );
  NAND4_X1 U9423 ( .A1(n7779), .A2(n7778), .A3(n7777), .A4(n7776), .ZN(n7780)
         );
  NOR4_X1 U9424 ( .A1(n7783), .A2(n7782), .A3(n7781), .A4(n7780), .ZN(n7785)
         );
  NAND4_X1 U9425 ( .A1(n7787), .A2(n7786), .A3(n7785), .A4(n7784), .ZN(n7788)
         );
  NOR4_X1 U9426 ( .A1(n8290), .A2(n4593), .A3(n7789), .A4(n7788), .ZN(n7790)
         );
  NAND4_X1 U9427 ( .A1(n8240), .A2(n8259), .A3(n8279), .A4(n7790), .ZN(n7791)
         );
  NOR4_X1 U9428 ( .A1(n8188), .A2(n8198), .A3(n8104), .A4(n7791), .ZN(n7793)
         );
  NAND4_X1 U9429 ( .A1(n8133), .A2(n7817), .A3(n7793), .A4(n7792), .ZN(n7794)
         );
  NOR4_X1 U9430 ( .A1(n7837), .A2(n7795), .A3(n8115), .A4(n7794), .ZN(n7796)
         );
  XNOR2_X1 U9431 ( .A(n7796), .B(n8077), .ZN(n7800) );
  OAI22_X1 U9432 ( .A1(n7800), .A2(n7799), .B1(n7798), .B2(n7797), .ZN(n7801)
         );
  NAND2_X1 U9433 ( .A1(n7803), .A2(n7802), .ZN(n7805) );
  INV_X1 U9434 ( .A(n8286), .ZN(n7806) );
  NOR2_X1 U9435 ( .A1(n8290), .A2(n7806), .ZN(n7807) );
  NAND2_X1 U9436 ( .A1(n7811), .A2(n7810), .ZN(n8258) );
  INV_X1 U9437 ( .A(n8241), .ZN(n7812) );
  NOR2_X1 U9438 ( .A1(n4387), .A2(n7812), .ZN(n7813) );
  NAND2_X1 U9439 ( .A1(n8257), .A2(n7813), .ZN(n8239) );
  NAND2_X1 U9440 ( .A1(n8239), .A2(n7814), .ZN(n8216) );
  NOR2_X1 U9441 ( .A1(n8198), .A2(n7815), .ZN(n7816) );
  AND2_X1 U9442 ( .A1(n8169), .A2(n7820), .ZN(n7818) );
  NAND2_X1 U9443 ( .A1(n8168), .A2(n7818), .ZN(n7824) );
  INV_X1 U9444 ( .A(n7819), .ZN(n7822) );
  INV_X1 U9445 ( .A(n7820), .ZN(n7821) );
  INV_X1 U9446 ( .A(n8188), .ZN(n8170) );
  NAND2_X1 U9447 ( .A1(n7824), .A2(n7823), .ZN(n8156) );
  NOR2_X1 U9448 ( .A1(n8085), .A2(n7827), .ZN(n7831) );
  INV_X1 U9449 ( .A(n7828), .ZN(n7829) );
  AOI21_X1 U9450 ( .B1(n8089), .B2(n7831), .A(n7829), .ZN(n7834) );
  OAI21_X1 U9451 ( .B1(n7838), .B2(n7837), .A(n7836), .ZN(n7840) );
  XNOR2_X1 U9452 ( .A(n7840), .B(n8077), .ZN(n7843) );
  NAND2_X1 U9453 ( .A1(n4250), .A2(n7841), .ZN(n7842) );
  INV_X1 U9454 ( .A(n7844), .ZN(n8084) );
  NAND4_X1 U9455 ( .A1(n7846), .A2(n8084), .A3(n7845), .A4(n8312), .ZN(n7847)
         );
  OAI211_X1 U9456 ( .C1(n5533), .C2(n7849), .A(n7847), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7848) );
  INV_X1 U9457 ( .A(n8606), .ZN(n8466) );
  OAI222_X1 U9458 ( .A1(n7852), .A2(n8607), .B1(P1_U3084), .B2(n5614), .C1(
        n4249), .C2(n8466), .ZN(P1_U3324) );
  INV_X1 U9459 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8596) );
  OAI222_X1 U9460 ( .A1(n7852), .A2(n8596), .B1(n4249), .B2(n7851), .C1(n7850), 
        .C2(P1_U3084), .ZN(P1_U3323) );
  XNOR2_X1 U9461 ( .A(n7853), .B(n7897), .ZN(n7858) );
  OAI22_X1 U9462 ( .A1(n7925), .A2(n8224), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7854), .ZN(n7856) );
  OAI22_X1 U9463 ( .A1(n7946), .A2(n7939), .B1(n7938), .B2(n7872), .ZN(n7855)
         );
  AOI211_X1 U9464 ( .C1(n7627), .C2(n7929), .A(n7856), .B(n7855), .ZN(n7857)
         );
  OAI21_X1 U9465 ( .B1(n7858), .B2(n7931), .A(n7857), .ZN(P2_U3218) );
  INV_X1 U9466 ( .A(n4341), .ZN(n7860) );
  AOI21_X1 U9467 ( .B1(n7862), .B2(n7861), .A(n7860), .ZN(n7867) );
  INV_X1 U9468 ( .A(n8097), .ZN(n8099) );
  AOI22_X1 U9469 ( .A1(n8260), .A2(n8313), .B1(n8099), .B2(n8312), .ZN(n8291)
         );
  NAND2_X1 U9470 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8080) );
  NAND2_X1 U9471 ( .A1(n7942), .A2(n8295), .ZN(n7863) );
  OAI211_X1 U9472 ( .C1(n7864), .C2(n8291), .A(n8080), .B(n7863), .ZN(n7865)
         );
  AOI21_X1 U9473 ( .B1(n8399), .B2(n7929), .A(n7865), .ZN(n7866) );
  OAI21_X1 U9474 ( .B1(n7867), .B2(n7931), .A(n7866), .ZN(P2_U3221) );
  XNOR2_X1 U9475 ( .A(n7868), .B(n7869), .ZN(n7876) );
  INV_X1 U9476 ( .A(n8254), .ZN(n7870) );
  OAI22_X1 U9477 ( .A1(n7925), .A2(n7870), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9424), .ZN(n7874) );
  OAI22_X1 U9478 ( .A1(n7872), .A2(n7939), .B1(n7938), .B2(n7871), .ZN(n7873)
         );
  AOI211_X1 U9479 ( .C1(n8385), .C2(n7929), .A(n7874), .B(n7873), .ZN(n7875)
         );
  OAI21_X1 U9480 ( .B1(n7876), .B2(n7931), .A(n7875), .ZN(P2_U3225) );
  INV_X1 U9481 ( .A(n7878), .ZN(n7880) );
  NAND2_X1 U9482 ( .A1(n7880), .A2(n7879), .ZN(n7881) );
  XNOR2_X1 U9483 ( .A(n7877), .B(n7881), .ZN(n7885) );
  OAI22_X1 U9484 ( .A1(n8157), .A2(n9861), .B1(n7946), .B2(n9863), .ZN(n8185)
         );
  AOI22_X1 U9485 ( .A1(n8185), .A2(n7890), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n7882) );
  OAI21_X1 U9486 ( .B1(n8192), .B2(n7925), .A(n7882), .ZN(n7883) );
  AOI21_X1 U9487 ( .B1(n8366), .B2(n7929), .A(n7883), .ZN(n7884) );
  OAI21_X1 U9488 ( .B1(n7885), .B2(n7931), .A(n7884), .ZN(P2_U3227) );
  XNOR2_X1 U9489 ( .A(n7886), .B(n7887), .ZN(n7895) );
  AOI21_X1 U9490 ( .B1(n7890), .B2(n7889), .A(n7888), .ZN(n7891) );
  OAI21_X1 U9491 ( .B1(n7892), .B2(n7925), .A(n7891), .ZN(n7893) );
  AOI21_X1 U9492 ( .B1(n8093), .B2(n7929), .A(n7893), .ZN(n7894) );
  OAI21_X1 U9493 ( .B1(n7895), .B2(n7931), .A(n7894), .ZN(P2_U3230) );
  OAI21_X1 U9494 ( .B1(n7853), .B2(n7897), .A(n7896), .ZN(n7901) );
  XNOR2_X1 U9495 ( .A(n7899), .B(n7898), .ZN(n7900) );
  XNOR2_X1 U9496 ( .A(n7901), .B(n7900), .ZN(n7906) );
  OAI22_X1 U9497 ( .A1(n7925), .A2(n8202), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7902), .ZN(n7904) );
  OAI22_X1 U9498 ( .A1(n8210), .A2(n7939), .B1(n7938), .B2(n8244), .ZN(n7903)
         );
  AOI211_X1 U9499 ( .C1(n8371), .C2(n7929), .A(n7904), .B(n7903), .ZN(n7905)
         );
  OAI21_X1 U9500 ( .B1(n7906), .B2(n7931), .A(n7905), .ZN(P2_U3231) );
  XNOR2_X1 U9501 ( .A(n7908), .B(n7907), .ZN(n7913) );
  OAI22_X1 U9502 ( .A1(n7925), .A2(n8273), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7909), .ZN(n7911) );
  OAI22_X1 U9503 ( .A1(n8269), .A2(n7939), .B1(n7938), .B2(n8268), .ZN(n7910)
         );
  AOI211_X1 U9504 ( .C1(n8276), .C2(n7929), .A(n7911), .B(n7910), .ZN(n7912)
         );
  OAI21_X1 U9505 ( .B1(n7913), .B2(n7931), .A(n7912), .ZN(P2_U3235) );
  INV_X1 U9506 ( .A(n8380), .ZN(n8238) );
  OAI21_X1 U9507 ( .B1(n7916), .B2(n7915), .A(n7914), .ZN(n7917) );
  NAND2_X1 U9508 ( .A1(n7917), .A2(n7933), .ZN(n7921) );
  NOR2_X1 U9509 ( .A1(n7925), .A2(n8235), .ZN(n7919) );
  OAI22_X1 U9510 ( .A1(n8244), .A2(n7939), .B1(n7938), .B2(n8269), .ZN(n7918)
         );
  AOI211_X1 U9511 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3152), .A(n7919), 
        .B(n7918), .ZN(n7920) );
  OAI211_X1 U9512 ( .C1(n8238), .C2(n7945), .A(n7921), .B(n7920), .ZN(P2_U3237) );
  XNOR2_X1 U9513 ( .A(n7922), .B(n7923), .ZN(n7932) );
  OAI21_X1 U9514 ( .B1(n7925), .B2(n8304), .A(n7924), .ZN(n7928) );
  OAI22_X1 U9515 ( .A1(n8268), .A2(n7939), .B1(n7938), .B2(n7926), .ZN(n7927)
         );
  AOI211_X1 U9516 ( .C1(n8402), .C2(n7929), .A(n7928), .B(n7927), .ZN(n7930)
         );
  OAI21_X1 U9517 ( .B1(n7932), .B2(n7931), .A(n7930), .ZN(P2_U3240) );
  OAI211_X1 U9518 ( .C1(n7936), .C2(n7935), .A(n7934), .B(n7933), .ZN(n7944)
         );
  NOR2_X1 U9519 ( .A1(n7937), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7941) );
  OAI22_X1 U9520 ( .A1(n8176), .A2(n7939), .B1(n7938), .B2(n8210), .ZN(n7940)
         );
  AOI211_X1 U9521 ( .C1(n7942), .C2(n8178), .A(n7941), .B(n7940), .ZN(n7943)
         );
  OAI211_X1 U9522 ( .C1(n8181), .C2(n7945), .A(n7944), .B(n7943), .ZN(P2_U3242) );
  MUX2_X1 U9523 ( .A(n8119), .B(P2_DATAO_REG_30__SCAN_IN), .S(n7961), .Z(
        P2_U3582) );
  MUX2_X1 U9524 ( .A(n4482), .B(P2_DATAO_REG_28__SCAN_IN), .S(n7961), .Z(
        P2_U3580) );
  INV_X1 U9525 ( .A(n8176), .ZN(n8110) );
  MUX2_X1 U9526 ( .A(n8110), .B(P2_DATAO_REG_27__SCAN_IN), .S(n7961), .Z(
        P2_U3579) );
  MUX2_X1 U9527 ( .A(n8108), .B(P2_DATAO_REG_26__SCAN_IN), .S(n7961), .Z(
        P2_U3578) );
  INV_X1 U9528 ( .A(n8210), .ZN(n8106) );
  MUX2_X1 U9529 ( .A(n8106), .B(P2_DATAO_REG_25__SCAN_IN), .S(n7961), .Z(
        P2_U3577) );
  INV_X1 U9530 ( .A(n7946), .ZN(n8220) );
  MUX2_X1 U9531 ( .A(n8220), .B(P2_DATAO_REG_24__SCAN_IN), .S(n7961), .Z(
        P2_U3576) );
  MUX2_X1 U9532 ( .A(n7947), .B(P2_DATAO_REG_23__SCAN_IN), .S(n7961), .Z(
        P2_U3575) );
  MUX2_X1 U9533 ( .A(n8261), .B(P2_DATAO_REG_22__SCAN_IN), .S(n7961), .Z(
        P2_U3574) );
  MUX2_X1 U9534 ( .A(n8102), .B(P2_DATAO_REG_21__SCAN_IN), .S(n7961), .Z(
        P2_U3573) );
  MUX2_X1 U9535 ( .A(n8260), .B(P2_DATAO_REG_20__SCAN_IN), .S(n7961), .Z(
        P2_U3572) );
  INV_X1 U9536 ( .A(n8268), .ZN(n8314) );
  MUX2_X1 U9537 ( .A(n8314), .B(P2_DATAO_REG_19__SCAN_IN), .S(n7961), .Z(
        P2_U3571) );
  MUX2_X1 U9538 ( .A(n8099), .B(P2_DATAO_REG_18__SCAN_IN), .S(n7961), .Z(
        P2_U3570) );
  MUX2_X1 U9539 ( .A(n8311), .B(P2_DATAO_REG_17__SCAN_IN), .S(n7961), .Z(
        P2_U3569) );
  MUX2_X1 U9540 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n7948), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9541 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n7949), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9542 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n7950), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9543 ( .A(n7951), .B(P2_DATAO_REG_13__SCAN_IN), .S(n7961), .Z(
        P2_U3565) );
  MUX2_X1 U9544 ( .A(n7952), .B(P2_DATAO_REG_12__SCAN_IN), .S(n7961), .Z(
        P2_U3564) );
  MUX2_X1 U9545 ( .A(n4704), .B(P2_DATAO_REG_11__SCAN_IN), .S(n7961), .Z(
        P2_U3563) );
  MUX2_X1 U9546 ( .A(n7953), .B(P2_DATAO_REG_10__SCAN_IN), .S(n7961), .Z(
        P2_U3562) );
  MUX2_X1 U9547 ( .A(n7954), .B(P2_DATAO_REG_9__SCAN_IN), .S(n7961), .Z(
        P2_U3561) );
  MUX2_X1 U9548 ( .A(n7955), .B(P2_DATAO_REG_8__SCAN_IN), .S(n7961), .Z(
        P2_U3560) );
  MUX2_X1 U9549 ( .A(n7956), .B(P2_DATAO_REG_7__SCAN_IN), .S(n7961), .Z(
        P2_U3559) );
  MUX2_X1 U9550 ( .A(n7957), .B(P2_DATAO_REG_6__SCAN_IN), .S(n7961), .Z(
        P2_U3558) );
  MUX2_X1 U9551 ( .A(n7958), .B(P2_DATAO_REG_5__SCAN_IN), .S(n7961), .Z(
        P2_U3557) );
  MUX2_X1 U9552 ( .A(n7959), .B(P2_DATAO_REG_4__SCAN_IN), .S(n7961), .Z(
        P2_U3556) );
  MUX2_X1 U9553 ( .A(n7960), .B(P2_DATAO_REG_3__SCAN_IN), .S(n7961), .Z(
        P2_U3555) );
  MUX2_X1 U9554 ( .A(n4248), .B(P2_DATAO_REG_2__SCAN_IN), .S(n7961), .Z(
        P2_U3554) );
  MUX2_X1 U9555 ( .A(n6704), .B(P2_DATAO_REG_1__SCAN_IN), .S(n7961), .Z(
        P2_U3553) );
  NOR2_X1 U9556 ( .A1(n4410), .A2(n4874), .ZN(n7963) );
  OAI211_X1 U9557 ( .C1(n7964), .C2(n7963), .A(n9844), .B(n7962), .ZN(n7972)
         );
  AOI22_X1 U9558 ( .A1(n9850), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n7971) );
  NAND2_X1 U9559 ( .A1(n9556), .A2(n7965), .ZN(n7970) );
  OAI211_X1 U9560 ( .C1(n7968), .C2(n7967), .A(n9845), .B(n7966), .ZN(n7969)
         );
  NAND4_X1 U9561 ( .A1(n7972), .A2(n7971), .A3(n7970), .A4(n7969), .ZN(
        P2_U3246) );
  INV_X1 U9562 ( .A(n7987), .ZN(n7976) );
  NAND3_X1 U9563 ( .A1(n9557), .A2(n7974), .A3(n7973), .ZN(n7975) );
  NAND3_X1 U9564 ( .A1(n9844), .A2(n7976), .A3(n7975), .ZN(n7985) );
  AOI21_X1 U9565 ( .B1(n9850), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n7977), .ZN(
        n7984) );
  NAND2_X1 U9566 ( .A1(n9556), .A2(n7978), .ZN(n7983) );
  OAI211_X1 U9567 ( .C1(n7981), .C2(n7980), .A(n9845), .B(n7979), .ZN(n7982)
         );
  NAND4_X1 U9568 ( .A1(n7985), .A2(n7984), .A3(n7983), .A4(n7982), .ZN(
        P2_U3248) );
  OR3_X1 U9569 ( .A1(n7988), .A2(n7987), .A3(n7986), .ZN(n7989) );
  NAND3_X1 U9570 ( .A1(n9844), .A2(n7990), .A3(n7989), .ZN(n8000) );
  INV_X1 U9571 ( .A(n7991), .ZN(n7992) );
  AOI21_X1 U9572 ( .B1(n9850), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n7992), .ZN(
        n7999) );
  NAND2_X1 U9573 ( .A1(n9556), .A2(n7993), .ZN(n7998) );
  OAI211_X1 U9574 ( .C1(n7996), .C2(n7995), .A(n9845), .B(n7994), .ZN(n7997)
         );
  NAND4_X1 U9575 ( .A1(n8000), .A2(n7999), .A3(n7998), .A4(n7997), .ZN(
        P2_U3249) );
  OAI211_X1 U9576 ( .C1(n8003), .C2(n8002), .A(n9844), .B(n8001), .ZN(n8013)
         );
  NOR2_X1 U9577 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8004), .ZN(n8005) );
  AOI21_X1 U9578 ( .B1(n9850), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8005), .ZN(
        n8012) );
  NAND2_X1 U9579 ( .A1(n9556), .A2(n8006), .ZN(n8011) );
  OAI211_X1 U9580 ( .C1(n8009), .C2(n8008), .A(n9845), .B(n8007), .ZN(n8010)
         );
  NAND4_X1 U9581 ( .A1(n8013), .A2(n8012), .A3(n8011), .A4(n8010), .ZN(
        P2_U3250) );
  OAI211_X1 U9582 ( .C1(n8016), .C2(n8015), .A(n9844), .B(n8014), .ZN(n8026)
         );
  INV_X1 U9583 ( .A(n8017), .ZN(n8018) );
  AOI21_X1 U9584 ( .B1(n9850), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8018), .ZN(
        n8025) );
  NAND2_X1 U9585 ( .A1(n9556), .A2(n8019), .ZN(n8024) );
  OAI211_X1 U9586 ( .C1(n8022), .C2(n8021), .A(n9845), .B(n8020), .ZN(n8023)
         );
  NAND4_X1 U9587 ( .A1(n8026), .A2(n8025), .A3(n8024), .A4(n8023), .ZN(
        P2_U3251) );
  OAI211_X1 U9588 ( .C1(n8029), .C2(n8028), .A(n9844), .B(n8027), .ZN(n8038)
         );
  NOR2_X1 U9589 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9410), .ZN(n8030) );
  AOI21_X1 U9590 ( .B1(n9850), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8030), .ZN(
        n8037) );
  NAND2_X1 U9591 ( .A1(n9556), .A2(n8031), .ZN(n8036) );
  OAI211_X1 U9592 ( .C1(n8034), .C2(n8033), .A(n9845), .B(n8032), .ZN(n8035)
         );
  NAND4_X1 U9593 ( .A1(n8038), .A2(n8037), .A3(n8036), .A4(n8035), .ZN(
        P2_U3252) );
  OAI211_X1 U9594 ( .C1(n8041), .C2(n8040), .A(n9844), .B(n8039), .ZN(n8051)
         );
  INV_X1 U9595 ( .A(n8042), .ZN(n8043) );
  AOI21_X1 U9596 ( .B1(n9850), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8043), .ZN(
        n8050) );
  NAND2_X1 U9597 ( .A1(n9556), .A2(n8044), .ZN(n8049) );
  OAI211_X1 U9598 ( .C1(n8047), .C2(n8046), .A(n9845), .B(n8045), .ZN(n8048)
         );
  NAND4_X1 U9599 ( .A1(n8051), .A2(n8050), .A3(n8049), .A4(n8048), .ZN(
        P2_U3253) );
  OAI211_X1 U9600 ( .C1(n8054), .C2(n8053), .A(n9844), .B(n8052), .ZN(n8064)
         );
  INV_X1 U9601 ( .A(n8055), .ZN(n8056) );
  AOI21_X1 U9602 ( .B1(n9850), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8056), .ZN(
        n8063) );
  NAND2_X1 U9603 ( .A1(n9556), .A2(n8057), .ZN(n8062) );
  OAI211_X1 U9604 ( .C1(n8060), .C2(n8059), .A(n9845), .B(n8058), .ZN(n8061)
         );
  NAND4_X1 U9605 ( .A1(n8064), .A2(n8063), .A3(n8062), .A4(n8061), .ZN(
        P2_U3254) );
  NOR2_X1 U9606 ( .A1(n8066), .A2(n8065), .ZN(n8067) );
  XOR2_X1 U9607 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8067), .Z(n8074) );
  INV_X1 U9608 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8068) );
  AOI22_X1 U9609 ( .A1(n8071), .A2(n8070), .B1(n8069), .B2(n8068), .ZN(n8072)
         );
  XNOR2_X1 U9610 ( .A(n8072), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8076) );
  INV_X1 U9611 ( .A(n8076), .ZN(n8073) );
  AOI22_X1 U9612 ( .A1(n8074), .A2(n9844), .B1(n8073), .B2(n9845), .ZN(n8079)
         );
  NOR2_X1 U9613 ( .A1(n8074), .A2(n9848), .ZN(n8075) );
  AOI211_X1 U9614 ( .C1(n9845), .C2(n8076), .A(n9556), .B(n8075), .ZN(n8078)
         );
  MUX2_X1 U9615 ( .A(n8079), .B(n8078), .S(n8077), .Z(n8081) );
  OAI211_X1 U9616 ( .C1(n8082), .C2(n4719), .A(n8081), .B(n8080), .ZN(P2_U3264) );
  INV_X1 U9617 ( .A(n8385), .ZN(n8256) );
  INV_X1 U9618 ( .A(n8366), .ZN(n8191) );
  XOR2_X1 U9619 ( .A(n8340), .B(n8088), .Z(n8342) );
  NOR2_X1 U9620 ( .A1(n8336), .A2(n8083), .ZN(n8086) );
  AOI21_X1 U9621 ( .B1(n8084), .B2(P2_B_REG_SCAN_IN), .A(n9861), .ZN(n8120) );
  NAND2_X1 U9622 ( .A1(n8120), .A2(n8085), .ZN(n9568) );
  NOR2_X1 U9623 ( .A1(n4247), .A2(n9568), .ZN(n8090) );
  AOI211_X1 U9624 ( .C1(n8340), .C2(n8324), .A(n8086), .B(n8090), .ZN(n8087)
         );
  OAI21_X1 U9625 ( .B1(n8342), .B2(n8278), .A(n8087), .ZN(P2_U3265) );
  INV_X1 U9626 ( .A(n8089), .ZN(n9569) );
  AOI21_X1 U9627 ( .B1(n8089), .B2(n8123), .A(n8088), .ZN(n9571) );
  NAND2_X1 U9628 ( .A1(n9571), .A2(n8319), .ZN(n8092) );
  AOI21_X1 U9629 ( .B1(n4247), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8090), .ZN(
        n8091) );
  OAI211_X1 U9630 ( .C1(n9569), .C2(n8307), .A(n8092), .B(n8091), .ZN(P2_U3266) );
  INV_X1 U9631 ( .A(n8093), .ZN(n8094) );
  NAND2_X1 U9632 ( .A1(n8094), .A2(n7926), .ZN(n8095) );
  NOR2_X1 U9633 ( .A1(n8280), .A2(n8279), .ZN(n8391) );
  NOR2_X1 U9634 ( .A1(n8385), .A2(n8102), .ZN(n8103) );
  INV_X1 U9635 ( .A(n8218), .ZN(n8104) );
  OAI21_X1 U9636 ( .B1(n8105), .B2(n8244), .A(n8222), .ZN(n8199) );
  OAI22_X1 U9637 ( .A1(n8199), .A2(n8206), .B1(n8220), .B2(n8371), .ZN(n8189)
         );
  NAND2_X1 U9638 ( .A1(n8189), .A2(n8188), .ZN(n8187) );
  NAND2_X1 U9639 ( .A1(n8187), .A2(n8107), .ZN(n8166) );
  NAND2_X1 U9640 ( .A1(n8166), .A2(n8174), .ZN(n8165) );
  NAND2_X1 U9641 ( .A1(n8165), .A2(n8109), .ZN(n8147) );
  INV_X1 U9642 ( .A(n8355), .ZN(n8111) );
  XNOR2_X1 U9643 ( .A(n8113), .B(n8115), .ZN(n8343) );
  INV_X1 U9644 ( .A(n8343), .ZN(n8131) );
  INV_X1 U9645 ( .A(n8114), .ZN(n8116) );
  NOR2_X1 U9646 ( .A1(n8116), .A2(n4487), .ZN(n8117) );
  AOI22_X1 U9647 ( .A1(n4482), .A2(n8312), .B1(n8120), .B2(n8119), .ZN(n8121)
         );
  OAI21_X1 U9648 ( .B1(n8139), .B2(n8127), .A(n8123), .ZN(n8344) );
  NOR2_X1 U9649 ( .A1(n8344), .A2(n8278), .ZN(n8129) );
  INV_X1 U9650 ( .A(n8124), .ZN(n8125) );
  AOI22_X1 U9651 ( .A1(n4247), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8125), .B2(
        n9869), .ZN(n8126) );
  OAI21_X1 U9652 ( .B1(n8127), .B2(n8307), .A(n8126), .ZN(n8128) );
  OAI21_X1 U9653 ( .B1(n8131), .B2(n8321), .A(n8130), .ZN(P2_U3267) );
  XNOR2_X1 U9654 ( .A(n8132), .B(n8133), .ZN(n8136) );
  OAI22_X1 U9655 ( .A1(n8134), .A2(n9861), .B1(n8176), .B2(n9863), .ZN(n8135)
         );
  AOI21_X1 U9656 ( .B1(n8136), .B2(n9865), .A(n8135), .ZN(n8353) );
  AOI21_X1 U9657 ( .B1(n8350), .B2(n8149), .A(n8139), .ZN(n8351) );
  NAND2_X1 U9658 ( .A1(n8351), .A2(n8319), .ZN(n8143) );
  INV_X1 U9659 ( .A(n8140), .ZN(n8141) );
  AOI22_X1 U9660 ( .A1(n4247), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8141), .B2(
        n9869), .ZN(n8142) );
  OAI211_X1 U9661 ( .C1(n4486), .C2(n8307), .A(n8143), .B(n8142), .ZN(n8144)
         );
  AOI21_X1 U9662 ( .B1(n8349), .B2(n8325), .A(n8144), .ZN(n8145) );
  OAI21_X1 U9663 ( .B1(n4247), .B2(n8353), .A(n8145), .ZN(P2_U3268) );
  OAI21_X1 U9664 ( .B1(n8147), .B2(n8155), .A(n8146), .ZN(n8148) );
  INV_X1 U9665 ( .A(n8148), .ZN(n8359) );
  INV_X1 U9666 ( .A(n8177), .ZN(n8151) );
  INV_X1 U9667 ( .A(n8149), .ZN(n8150) );
  AOI21_X1 U9668 ( .B1(n8355), .B2(n8151), .A(n8150), .ZN(n8356) );
  INV_X1 U9669 ( .A(n8152), .ZN(n8153) );
  AOI22_X1 U9670 ( .A1(n4247), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8153), .B2(
        n9869), .ZN(n8154) );
  OAI21_X1 U9671 ( .B1(n8111), .B2(n8307), .A(n8154), .ZN(n8163) );
  AOI21_X1 U9672 ( .B1(n8156), .B2(n8155), .A(n8292), .ZN(n8161) );
  OAI22_X1 U9673 ( .A1(n8158), .A2(n9861), .B1(n8157), .B2(n9863), .ZN(n8159)
         );
  AOI21_X1 U9674 ( .B1(n8161), .B2(n8160), .A(n8159), .ZN(n8358) );
  NOR2_X1 U9675 ( .A1(n8358), .A2(n4247), .ZN(n8162) );
  AOI211_X1 U9676 ( .C1(n8356), .C2(n8319), .A(n8163), .B(n8162), .ZN(n8164)
         );
  OAI21_X1 U9677 ( .B1(n8359), .B2(n8321), .A(n8164), .ZN(P2_U3269) );
  OAI21_X1 U9678 ( .B1(n8166), .B2(n8174), .A(n8165), .ZN(n8167) );
  INV_X1 U9679 ( .A(n8167), .ZN(n8364) );
  NAND2_X1 U9680 ( .A1(n8168), .A2(n8169), .ZN(n8184) );
  NAND2_X1 U9681 ( .A1(n8184), .A2(n8170), .ZN(n8172) );
  NAND2_X1 U9682 ( .A1(n8172), .A2(n8171), .ZN(n8173) );
  OAI222_X1 U9683 ( .A1(n9861), .A2(n8176), .B1(n9863), .B2(n8210), .C1(n8292), 
        .C2(n8175), .ZN(n8360) );
  AOI211_X1 U9684 ( .C1(n8362), .C2(n8190), .A(n9985), .B(n8177), .ZN(n8361)
         );
  NAND2_X1 U9685 ( .A1(n8361), .A2(n8328), .ZN(n8180) );
  AOI22_X1 U9686 ( .A1(n4247), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8178), .B2(
        n9869), .ZN(n8179) );
  OAI211_X1 U9687 ( .C1(n8181), .C2(n8307), .A(n8180), .B(n8179), .ZN(n8182)
         );
  AOI21_X1 U9688 ( .B1(n8360), .B2(n8336), .A(n8182), .ZN(n8183) );
  OAI21_X1 U9689 ( .B1(n8364), .B2(n8321), .A(n8183), .ZN(P2_U3270) );
  XNOR2_X1 U9690 ( .A(n8184), .B(n8188), .ZN(n8186) );
  AOI21_X1 U9691 ( .B1(n8186), .B2(n9865), .A(n8185), .ZN(n8369) );
  OAI21_X1 U9692 ( .B1(n8189), .B2(n8188), .A(n8187), .ZN(n8365) );
  OAI211_X1 U9693 ( .C1(n8191), .C2(n8200), .A(n9946), .B(n8190), .ZN(n8368)
         );
  OAI22_X1 U9694 ( .A1(n8336), .A2(n9450), .B1(n8192), .B2(n8272), .ZN(n8193)
         );
  AOI21_X1 U9695 ( .B1(n8366), .B2(n8324), .A(n8193), .ZN(n8194) );
  OAI21_X1 U9696 ( .B1(n8368), .B2(n8195), .A(n8194), .ZN(n8196) );
  AOI21_X1 U9697 ( .B1(n8365), .B2(n8325), .A(n8196), .ZN(n8197) );
  OAI21_X1 U9698 ( .B1(n4247), .B2(n8369), .A(n8197), .ZN(P2_U3271) );
  XNOR2_X1 U9699 ( .A(n8199), .B(n8198), .ZN(n8375) );
  INV_X1 U9700 ( .A(n8228), .ZN(n8201) );
  AOI21_X1 U9701 ( .B1(n8371), .B2(n8201), .A(n8200), .ZN(n8372) );
  INV_X1 U9702 ( .A(n8202), .ZN(n8203) );
  AOI22_X1 U9703 ( .A1(n4247), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8203), .B2(
        n9869), .ZN(n8204) );
  OAI21_X1 U9704 ( .B1(n8205), .B2(n8307), .A(n8204), .ZN(n8214) );
  INV_X1 U9705 ( .A(n8168), .ZN(n8209) );
  AOI21_X1 U9706 ( .B1(n8217), .B2(n8207), .A(n8206), .ZN(n8208) );
  NOR3_X1 U9707 ( .A1(n8209), .A2(n8208), .A3(n8292), .ZN(n8212) );
  OAI22_X1 U9708 ( .A1(n8210), .A2(n9861), .B1(n8244), .B2(n9863), .ZN(n8211)
         );
  NOR2_X1 U9709 ( .A1(n8212), .A2(n8211), .ZN(n8374) );
  NOR2_X1 U9710 ( .A1(n8374), .A2(n4247), .ZN(n8213) );
  AOI211_X1 U9711 ( .C1(n8372), .C2(n8319), .A(n8214), .B(n8213), .ZN(n8215)
         );
  OAI21_X1 U9712 ( .B1(n8375), .B2(n8321), .A(n8215), .ZN(P2_U3272) );
  INV_X1 U9713 ( .A(n8216), .ZN(n8219) );
  OAI21_X1 U9714 ( .B1(n8219), .B2(n8218), .A(n8217), .ZN(n8221) );
  AOI222_X1 U9715 ( .A1(n9865), .A2(n8221), .B1(n8261), .B2(n8312), .C1(n8220), 
        .C2(n8313), .ZN(n8378) );
  OAI21_X1 U9716 ( .B1(n8223), .B2(n8104), .A(n8222), .ZN(n8379) );
  INV_X1 U9717 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8225) );
  OAI22_X1 U9718 ( .A1(n8336), .A2(n8225), .B1(n8224), .B2(n8272), .ZN(n8226)
         );
  AOI21_X1 U9719 ( .B1(n7627), .B2(n8324), .A(n8226), .ZN(n8230) );
  AND2_X1 U9720 ( .A1(n7627), .A2(n4807), .ZN(n8227) );
  NOR2_X1 U9721 ( .A1(n8228), .A2(n8227), .ZN(n8376) );
  NAND2_X1 U9722 ( .A1(n8376), .A2(n8319), .ZN(n8229) );
  OAI211_X1 U9723 ( .C1(n8379), .C2(n8321), .A(n8230), .B(n8229), .ZN(n8231)
         );
  INV_X1 U9724 ( .A(n8231), .ZN(n8232) );
  OAI21_X1 U9725 ( .B1(n4247), .B2(n8378), .A(n8232), .ZN(P2_U3273) );
  XNOR2_X1 U9726 ( .A(n8233), .B(n4387), .ZN(n8384) );
  INV_X1 U9727 ( .A(n4807), .ZN(n8234) );
  AOI21_X1 U9728 ( .B1(n8380), .B2(n8251), .A(n8234), .ZN(n8381) );
  INV_X1 U9729 ( .A(n8235), .ZN(n8236) );
  AOI22_X1 U9730 ( .A1(n4247), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8236), .B2(
        n9869), .ZN(n8237) );
  OAI21_X1 U9731 ( .B1(n8238), .B2(n8307), .A(n8237), .ZN(n8248) );
  INV_X1 U9732 ( .A(n8239), .ZN(n8243) );
  AOI21_X1 U9733 ( .B1(n8257), .B2(n8241), .A(n8240), .ZN(n8242) );
  NOR3_X1 U9734 ( .A1(n8243), .A2(n8242), .A3(n8292), .ZN(n8246) );
  OAI22_X1 U9735 ( .A1(n8244), .A2(n9861), .B1(n8269), .B2(n9863), .ZN(n8245)
         );
  NOR2_X1 U9736 ( .A1(n8246), .A2(n8245), .ZN(n8383) );
  NOR2_X1 U9737 ( .A1(n8383), .A2(n4247), .ZN(n8247) );
  AOI211_X1 U9738 ( .C1(n8381), .C2(n8319), .A(n8248), .B(n8247), .ZN(n8249)
         );
  OAI21_X1 U9739 ( .B1(n8384), .B2(n8321), .A(n8249), .ZN(P2_U3274) );
  XNOR2_X1 U9740 ( .A(n8250), .B(n8259), .ZN(n8389) );
  INV_X1 U9741 ( .A(n8271), .ZN(n8253) );
  INV_X1 U9742 ( .A(n8251), .ZN(n8252) );
  AOI21_X1 U9743 ( .B1(n8385), .B2(n8253), .A(n8252), .ZN(n8386) );
  AOI22_X1 U9744 ( .A1(n4247), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8254), .B2(
        n9869), .ZN(n8255) );
  OAI21_X1 U9745 ( .B1(n8256), .B2(n8307), .A(n8255), .ZN(n8264) );
  OAI21_X1 U9746 ( .B1(n8259), .B2(n8258), .A(n8257), .ZN(n8262) );
  AOI222_X1 U9747 ( .A1(n9865), .A2(n8262), .B1(n8261), .B2(n8313), .C1(n8260), 
        .C2(n8312), .ZN(n8388) );
  NOR2_X1 U9748 ( .A1(n8388), .A2(n4247), .ZN(n8263) );
  AOI211_X1 U9749 ( .C1(n8386), .C2(n8319), .A(n8264), .B(n8263), .ZN(n8265)
         );
  OAI21_X1 U9750 ( .B1(n8389), .B2(n8321), .A(n8265), .ZN(P2_U3275) );
  XOR2_X1 U9751 ( .A(n8266), .B(n8279), .Z(n8267) );
  OAI222_X1 U9752 ( .A1(n9861), .A2(n8269), .B1(n9863), .B2(n8268), .C1(n8267), 
        .C2(n8292), .ZN(n8395) );
  NOR2_X1 U9753 ( .A1(n8294), .A2(n8392), .ZN(n8270) );
  OR2_X1 U9754 ( .A1(n8271), .A2(n8270), .ZN(n8393) );
  INV_X1 U9755 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8274) );
  OAI22_X1 U9756 ( .A1(n8336), .A2(n8274), .B1(n8273), .B2(n8272), .ZN(n8275)
         );
  AOI21_X1 U9757 ( .B1(n8276), .B2(n8324), .A(n8275), .ZN(n8277) );
  OAI21_X1 U9758 ( .B1(n8393), .B2(n8278), .A(n8277), .ZN(n8282) );
  AND2_X1 U9759 ( .A1(n8280), .A2(n8279), .ZN(n8390) );
  NOR3_X1 U9760 ( .A1(n8391), .A2(n8390), .A3(n8321), .ZN(n8281) );
  AOI211_X1 U9761 ( .C1(n8336), .C2(n8395), .A(n8282), .B(n8281), .ZN(n8283)
         );
  INV_X1 U9762 ( .A(n8283), .ZN(P2_U3276) );
  XOR2_X1 U9763 ( .A(n8284), .B(n8290), .Z(n8401) );
  NAND2_X1 U9764 ( .A1(n8285), .A2(n8286), .ZN(n8289) );
  INV_X1 U9765 ( .A(n8287), .ZN(n8288) );
  AOI21_X1 U9766 ( .B1(n8290), .B2(n8289), .A(n8288), .ZN(n8293) );
  OAI21_X1 U9767 ( .B1(n8293), .B2(n8292), .A(n8291), .ZN(n8397) );
  AOI211_X1 U9768 ( .C1(n8399), .C2(n8302), .A(n9985), .B(n8294), .ZN(n8398)
         );
  NAND2_X1 U9769 ( .A1(n8398), .A2(n8328), .ZN(n8297) );
  AOI22_X1 U9770 ( .A1(n4247), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8295), .B2(
        n9869), .ZN(n8296) );
  OAI211_X1 U9771 ( .C1(n8298), .C2(n8307), .A(n8297), .B(n8296), .ZN(n8299)
         );
  AOI21_X1 U9772 ( .B1(n8397), .B2(n8336), .A(n8299), .ZN(n8300) );
  OAI21_X1 U9773 ( .B1(n8401), .B2(n8321), .A(n8300), .ZN(P2_U3277) );
  XNOR2_X1 U9774 ( .A(n8301), .B(n8310), .ZN(n8406) );
  AOI21_X1 U9775 ( .B1(n8402), .B2(n8303), .A(n4415), .ZN(n8403) );
  INV_X1 U9776 ( .A(n8304), .ZN(n8305) );
  AOI22_X1 U9777 ( .A1(n4247), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8305), .B2(
        n9869), .ZN(n8306) );
  OAI21_X1 U9778 ( .B1(n8308), .B2(n8307), .A(n8306), .ZN(n8318) );
  OAI211_X1 U9779 ( .C1(n8310), .C2(n8309), .A(n8285), .B(n9865), .ZN(n8316)
         );
  AOI22_X1 U9780 ( .A1(n8314), .A2(n8313), .B1(n8312), .B2(n8311), .ZN(n8315)
         );
  NOR2_X1 U9781 ( .A1(n8405), .A2(n4247), .ZN(n8317) );
  AOI211_X1 U9782 ( .C1(n8403), .C2(n8319), .A(n8318), .B(n8317), .ZN(n8320)
         );
  OAI21_X1 U9783 ( .B1(n8406), .B2(n8321), .A(n8320), .ZN(P2_U3278) );
  XNOR2_X1 U9784 ( .A(n8329), .B(n8322), .ZN(n9939) );
  AOI22_X1 U9785 ( .A1(n8325), .A2(n9939), .B1(n8324), .B2(n8323), .ZN(n8339)
         );
  OAI21_X1 U9786 ( .B1(n8326), .B2(n9937), .A(n9946), .ZN(n8327) );
  NOR2_X1 U9787 ( .A1(n8327), .A2(n9871), .ZN(n9934) );
  AOI22_X1 U9788 ( .A1(n8328), .A2(n9934), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n9869), .ZN(n8338) );
  NAND2_X1 U9789 ( .A1(n8330), .A2(n8329), .ZN(n8331) );
  NAND2_X1 U9790 ( .A1(n8332), .A2(n8331), .ZN(n8335) );
  OAI22_X1 U9791 ( .A1(n6705), .A2(n9863), .B1(n8333), .B2(n9861), .ZN(n8334)
         );
  AOI21_X1 U9792 ( .B1(n8335), .B2(n9865), .A(n8334), .ZN(n9936) );
  MUX2_X1 U9793 ( .A(n6513), .B(n9936), .S(n8336), .Z(n8337) );
  NAND3_X1 U9794 ( .A1(n8339), .A2(n8338), .A3(n8337), .ZN(P2_U3294) );
  NAND2_X1 U9795 ( .A1(n8340), .A2(n9954), .ZN(n8341) );
  OAI211_X1 U9796 ( .C1(n8342), .C2(n9985), .A(n9568), .B(n8341), .ZN(n8439)
         );
  MUX2_X1 U9797 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8439), .S(n10008), .Z(
        P2_U3551) );
  NAND2_X1 U9798 ( .A1(n8343), .A2(n9989), .ZN(n8348) );
  NOR2_X1 U9799 ( .A1(n8344), .A2(n9985), .ZN(n8345) );
  NAND2_X1 U9800 ( .A1(n8348), .A2(n8347), .ZN(n8440) );
  MUX2_X1 U9801 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8440), .S(n10008), .Z(
        P2_U3549) );
  AOI22_X1 U9802 ( .A1(n8351), .A2(n9946), .B1(n9954), .B2(n8350), .ZN(n8352)
         );
  OAI211_X1 U9803 ( .C1(n8354), .C2(n9957), .A(n8353), .B(n8352), .ZN(n8441)
         );
  MUX2_X1 U9804 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8441), .S(n10008), .Z(
        P2_U3548) );
  AOI22_X1 U9805 ( .A1(n8356), .A2(n9946), .B1(n9954), .B2(n8355), .ZN(n8357)
         );
  OAI211_X1 U9806 ( .C1(n8359), .C2(n9957), .A(n8358), .B(n8357), .ZN(n8442)
         );
  MUX2_X1 U9807 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8442), .S(n10008), .Z(
        P2_U3547) );
  OAI21_X1 U9808 ( .B1(n8364), .B2(n9957), .A(n8363), .ZN(n8443) );
  MUX2_X1 U9809 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8443), .S(n10008), .Z(
        P2_U3546) );
  NAND2_X1 U9810 ( .A1(n8365), .A2(n9989), .ZN(n8370) );
  NAND2_X1 U9811 ( .A1(n8366), .A2(n9954), .ZN(n8367) );
  NAND4_X1 U9812 ( .A1(n8370), .A2(n8369), .A3(n8368), .A4(n8367), .ZN(n8444)
         );
  MUX2_X1 U9813 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8444), .S(n10008), .Z(
        P2_U3545) );
  AOI22_X1 U9814 ( .A1(n8372), .A2(n9946), .B1(n9954), .B2(n8371), .ZN(n8373)
         );
  OAI211_X1 U9815 ( .C1(n8375), .C2(n9957), .A(n8374), .B(n8373), .ZN(n8445)
         );
  MUX2_X1 U9816 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8445), .S(n10008), .Z(
        P2_U3544) );
  AOI22_X1 U9817 ( .A1(n8376), .A2(n9946), .B1(n9954), .B2(n7627), .ZN(n8377)
         );
  OAI211_X1 U9818 ( .C1(n8379), .C2(n9957), .A(n8378), .B(n8377), .ZN(n8446)
         );
  MUX2_X1 U9819 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8446), .S(n10008), .Z(
        P2_U3543) );
  AOI22_X1 U9820 ( .A1(n8381), .A2(n9946), .B1(n9954), .B2(n8380), .ZN(n8382)
         );
  OAI211_X1 U9821 ( .C1(n8384), .C2(n9957), .A(n8383), .B(n8382), .ZN(n8447)
         );
  MUX2_X1 U9822 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8447), .S(n10008), .Z(
        P2_U3542) );
  AOI22_X1 U9823 ( .A1(n8386), .A2(n9946), .B1(n9954), .B2(n8385), .ZN(n8387)
         );
  OAI211_X1 U9824 ( .C1(n8389), .C2(n9957), .A(n8388), .B(n8387), .ZN(n8448)
         );
  MUX2_X1 U9825 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8448), .S(n10008), .Z(
        P2_U3541) );
  NOR3_X1 U9826 ( .A1(n8391), .A2(n8390), .A3(n9957), .ZN(n8396) );
  OAI22_X1 U9827 ( .A1(n8393), .A2(n9985), .B1(n8392), .B2(n9983), .ZN(n8394)
         );
  MUX2_X1 U9828 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8449), .S(n10008), .Z(
        P2_U3540) );
  AOI211_X1 U9829 ( .C1(n9954), .C2(n8399), .A(n8398), .B(n8397), .ZN(n8400)
         );
  OAI21_X1 U9830 ( .B1(n8401), .B2(n9957), .A(n8400), .ZN(n8450) );
  MUX2_X1 U9831 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8450), .S(n10008), .Z(
        P2_U3539) );
  AOI22_X1 U9832 ( .A1(n8403), .A2(n9946), .B1(n9954), .B2(n8402), .ZN(n8404)
         );
  OAI211_X1 U9833 ( .C1(n8406), .C2(n9957), .A(n8405), .B(n8404), .ZN(n8451)
         );
  MUX2_X1 U9834 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8451), .S(n10008), .Z(
        P2_U3538) );
  OAI21_X1 U9835 ( .B1(n8094), .B2(n9983), .A(n8407), .ZN(n8408) );
  AOI21_X1 U9836 ( .B1(n8409), .B2(n9989), .A(n8408), .ZN(n8411) );
  NAND2_X1 U9837 ( .A1(n8411), .A2(n8410), .ZN(n8452) );
  MUX2_X1 U9838 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8452), .S(n10008), .Z(
        P2_U3537) );
  OAI21_X1 U9839 ( .B1(n8413), .B2(n9983), .A(n8412), .ZN(n8414) );
  AOI21_X1 U9840 ( .B1(n8415), .B2(n9989), .A(n8414), .ZN(n8417) );
  NAND2_X1 U9841 ( .A1(n8417), .A2(n8416), .ZN(n8453) );
  MUX2_X1 U9842 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8453), .S(n10008), .Z(
        P2_U3536) );
  INV_X1 U9843 ( .A(n8418), .ZN(n8423) );
  AOI22_X1 U9844 ( .A1(n8420), .A2(n9946), .B1(n9954), .B2(n8419), .ZN(n8421)
         );
  OAI211_X1 U9845 ( .C1(n8423), .C2(n9957), .A(n8422), .B(n8421), .ZN(n8454)
         );
  MUX2_X1 U9846 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8454), .S(n10008), .Z(
        P2_U3535) );
  AOI22_X1 U9847 ( .A1(n8425), .A2(n9946), .B1(n9954), .B2(n8424), .ZN(n8426)
         );
  OAI211_X1 U9848 ( .C1(n9967), .C2(n8428), .A(n8427), .B(n8426), .ZN(n8455)
         );
  MUX2_X1 U9849 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8455), .S(n10008), .Z(
        P2_U3533) );
  AOI22_X1 U9850 ( .A1(n8430), .A2(n9946), .B1(n9954), .B2(n8429), .ZN(n8431)
         );
  OAI211_X1 U9851 ( .C1(n9957), .C2(n8433), .A(n8432), .B(n8431), .ZN(n8456)
         );
  MUX2_X1 U9852 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n8456), .S(n10008), .Z(
        P2_U3531) );
  AOI22_X1 U9853 ( .A1(n8435), .A2(n9946), .B1(n9954), .B2(n8434), .ZN(n8436)
         );
  OAI211_X1 U9854 ( .C1(n8438), .C2(n9967), .A(n8437), .B(n8436), .ZN(n8457)
         );
  MUX2_X1 U9855 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n8457), .S(n10008), .Z(
        P2_U3529) );
  MUX2_X1 U9856 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8439), .S(n9993), .Z(
        P2_U3519) );
  MUX2_X1 U9857 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8440), .S(n9993), .Z(
        P2_U3517) );
  MUX2_X1 U9858 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8441), .S(n9993), .Z(
        P2_U3516) );
  MUX2_X1 U9859 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8442), .S(n9993), .Z(
        P2_U3515) );
  MUX2_X1 U9860 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8443), .S(n9993), .Z(
        P2_U3514) );
  MUX2_X1 U9861 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8444), .S(n9993), .Z(
        P2_U3513) );
  MUX2_X1 U9862 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8445), .S(n9993), .Z(
        P2_U3512) );
  MUX2_X1 U9863 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8446), .S(n9993), .Z(
        P2_U3511) );
  MUX2_X1 U9864 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8447), .S(n9993), .Z(
        P2_U3510) );
  MUX2_X1 U9865 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8448), .S(n9993), .Z(
        P2_U3509) );
  MUX2_X1 U9866 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8449), .S(n9993), .Z(
        P2_U3508) );
  MUX2_X1 U9867 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8450), .S(n9993), .Z(
        P2_U3507) );
  MUX2_X1 U9868 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8451), .S(n9993), .Z(
        P2_U3505) );
  MUX2_X1 U9869 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8452), .S(n9993), .Z(
        P2_U3502) );
  MUX2_X1 U9870 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8453), .S(n9993), .Z(
        P2_U3499) );
  MUX2_X1 U9871 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8454), .S(n9993), .Z(
        P2_U3496) );
  MUX2_X1 U9872 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8455), .S(n9993), .Z(
        P2_U3490) );
  MUX2_X1 U9873 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n8456), .S(n9993), .Z(
        P2_U3484) );
  MUX2_X1 U9874 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n8457), .S(n9993), .Z(
        P2_U3478) );
  INV_X1 U9875 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8459) );
  NAND3_X1 U9876 ( .A1(n8459), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8464) );
  NAND2_X1 U9877 ( .A1(n9543), .A2(n8460), .ZN(n8463) );
  NAND2_X1 U9878 ( .A1(n8461), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8462) );
  OAI211_X1 U9879 ( .C1(n8458), .C2(n8464), .A(n8463), .B(n8462), .ZN(P2_U3327) );
  OAI222_X1 U9880 ( .A1(n8468), .A2(P2_U3152), .B1(n8467), .B2(n8466), .C1(
        n9436), .C2(n8465), .ZN(P2_U3329) );
  MUX2_X1 U9881 ( .A(n8469), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U9882 ( .A1(n8470), .A2(n8471), .ZN(n8472) );
  XOR2_X1 U9883 ( .A(n8473), .B(n8472), .Z(n8479) );
  NAND2_X1 U9884 ( .A1(n8585), .A2(n8889), .ZN(n8475) );
  OAI211_X1 U9885 ( .C1(n8588), .C2(n9285), .A(n8475), .B(n8474), .ZN(n8477)
         );
  NOR2_X1 U9886 ( .A1(n9294), .A2(n8578), .ZN(n8476) );
  AOI211_X1 U9887 ( .C1(n9290), .C2(n8583), .A(n8477), .B(n8476), .ZN(n8478)
         );
  OAI21_X1 U9888 ( .B1(n8479), .B2(n8592), .A(n8478), .ZN(P1_U3213) );
  INV_X1 U9889 ( .A(n8530), .ZN(n8483) );
  AOI21_X1 U9890 ( .B1(n8480), .B2(n8529), .A(n8481), .ZN(n8482) );
  AOI21_X1 U9891 ( .B1(n8483), .B2(n8529), .A(n8482), .ZN(n8488) );
  NAND2_X1 U9892 ( .A1(n9127), .A2(n8552), .ZN(n8485) );
  AOI22_X1 U9893 ( .A1(n9167), .A2(n8585), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8484) );
  OAI211_X1 U9894 ( .C1(n8563), .C2(n9133), .A(n8485), .B(n8484), .ZN(n8486)
         );
  AOI21_X1 U9895 ( .B1(n9473), .B2(n8590), .A(n8486), .ZN(n8487) );
  OAI21_X1 U9896 ( .B1(n8488), .B2(n8592), .A(n8487), .ZN(P1_U3214) );
  XOR2_X1 U9897 ( .A(n8490), .B(n8489), .Z(n8495) );
  AOI22_X1 U9898 ( .A1(n8552), .A2(n9168), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3084), .ZN(n8492) );
  NAND2_X1 U9899 ( .A1(n8585), .A2(n9242), .ZN(n8491) );
  OAI211_X1 U9900 ( .C1(n8563), .C2(n9200), .A(n8492), .B(n8491), .ZN(n8493)
         );
  AOI21_X1 U9901 ( .B1(n9493), .B2(n8590), .A(n8493), .ZN(n8494) );
  OAI21_X1 U9902 ( .B1(n8495), .B2(n8592), .A(n8494), .ZN(P1_U3217) );
  XOR2_X1 U9903 ( .A(n8496), .B(n8497), .Z(n8502) );
  INV_X1 U9904 ( .A(n9167), .ZN(n8680) );
  AOI22_X1 U9905 ( .A1(n8585), .A2(n9168), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8499) );
  NAND2_X1 U9906 ( .A1(n8583), .A2(n9171), .ZN(n8498) );
  OAI211_X1 U9907 ( .C1(n8680), .C2(n8588), .A(n8499), .B(n8498), .ZN(n8500)
         );
  AOI21_X1 U9908 ( .B1(n9483), .B2(n8590), .A(n8500), .ZN(n8501) );
  OAI21_X1 U9909 ( .B1(n8502), .B2(n8592), .A(n8501), .ZN(P1_U3221) );
  AOI21_X1 U9910 ( .B1(n8504), .B2(n8503), .A(n8569), .ZN(n8509) );
  NAND2_X1 U9911 ( .A1(n9105), .A2(n8552), .ZN(n8506) );
  AOI22_X1 U9912 ( .A1(n9127), .A2(n8585), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8505) );
  OAI211_X1 U9913 ( .C1(n8563), .C2(n9099), .A(n8506), .B(n8505), .ZN(n8507)
         );
  AOI21_X1 U9914 ( .B1(n9321), .B2(n8590), .A(n8507), .ZN(n8508) );
  OAI21_X1 U9915 ( .B1(n8509), .B2(n8592), .A(n8508), .ZN(P1_U3223) );
  INV_X1 U9916 ( .A(n8511), .ZN(n8512) );
  AOI21_X1 U9917 ( .B1(n8513), .B2(n8510), .A(n8512), .ZN(n8518) );
  NAND2_X1 U9918 ( .A1(n8583), .A2(n9255), .ZN(n8515) );
  AOI22_X1 U9919 ( .A1(n8552), .A2(n9214), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n8514) );
  OAI211_X1 U9920 ( .C1(n9285), .C2(n8573), .A(n8515), .B(n8514), .ZN(n8516)
         );
  AOI21_X1 U9921 ( .B1(n9511), .B2(n8590), .A(n8516), .ZN(n8517) );
  OAI21_X1 U9922 ( .B1(n8518), .B2(n8592), .A(n8517), .ZN(P1_U3224) );
  INV_X1 U9923 ( .A(n9504), .ZN(n9239) );
  OAI21_X1 U9924 ( .B1(n8521), .B2(n8520), .A(n8519), .ZN(n8522) );
  NAND2_X1 U9925 ( .A1(n8522), .A2(n8571), .ZN(n8527) );
  NOR2_X1 U9926 ( .A1(n8523), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8949) );
  AOI21_X1 U9927 ( .B1(n8552), .B2(n9242), .A(n8949), .ZN(n8524) );
  OAI21_X1 U9928 ( .B1(n8573), .B2(n8645), .A(n8524), .ZN(n8525) );
  AOI21_X1 U9929 ( .B1(n9237), .B2(n8583), .A(n8525), .ZN(n8526) );
  OAI211_X1 U9930 ( .C1(n9239), .C2(n8578), .A(n8527), .B(n8526), .ZN(P1_U3226) );
  INV_X1 U9931 ( .A(n9327), .ZN(n9114) );
  AND3_X1 U9932 ( .A1(n8530), .A2(n8529), .A3(n8528), .ZN(n8531) );
  OAI21_X1 U9933 ( .B1(n8532), .B2(n8531), .A(n8571), .ZN(n8536) );
  AOI22_X1 U9934 ( .A1(n9121), .A2(n8585), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8533) );
  OAI21_X1 U9935 ( .B1(n8999), .B2(n8588), .A(n8533), .ZN(n8534) );
  AOI21_X1 U9936 ( .B1(n9112), .B2(n8583), .A(n8534), .ZN(n8535) );
  OAI211_X1 U9937 ( .C1(n9114), .C2(n8578), .A(n8536), .B(n8535), .ZN(P1_U3227) );
  NAND2_X1 U9938 ( .A1(n8538), .A2(n8537), .ZN(n8539) );
  XNOR2_X1 U9939 ( .A(n8540), .B(n8539), .ZN(n8546) );
  INV_X1 U9940 ( .A(n9186), .ZN(n9156) );
  OAI22_X1 U9941 ( .A1(n9156), .A2(n8588), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8541), .ZN(n8542) );
  AOI21_X1 U9942 ( .B1(n8585), .B2(n9215), .A(n8542), .ZN(n8543) );
  OAI21_X1 U9943 ( .B1(n8563), .B2(n9180), .A(n8543), .ZN(n8544) );
  AOI21_X1 U9944 ( .B1(n9487), .B2(n8590), .A(n8544), .ZN(n8545) );
  OAI21_X1 U9945 ( .B1(n8546), .B2(n8592), .A(n8545), .ZN(P1_U3231) );
  NAND2_X1 U9946 ( .A1(n10060), .A2(n8547), .ZN(n8549) );
  XOR2_X1 U9947 ( .A(n8550), .B(n8549), .Z(n8556) );
  OAI22_X1 U9948 ( .A1(n9156), .A2(n8573), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9457), .ZN(n8551) );
  AOI21_X1 U9949 ( .B1(n8552), .B2(n9121), .A(n8551), .ZN(n8553) );
  OAI21_X1 U9950 ( .B1(n8563), .B2(n9148), .A(n8553), .ZN(n8554) );
  AOI21_X1 U9951 ( .B1(n9479), .B2(n8590), .A(n8554), .ZN(n8555) );
  OAI21_X1 U9952 ( .B1(n8556), .B2(n8592), .A(n8555), .ZN(P1_U3233) );
  NAND2_X1 U9953 ( .A1(n8557), .A2(n8558), .ZN(n8559) );
  XOR2_X1 U9954 ( .A(n8560), .B(n8559), .Z(n8566) );
  INV_X1 U9955 ( .A(n9215), .ZN(n8668) );
  NAND2_X1 U9956 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9700) );
  OAI21_X1 U9957 ( .B1(n8588), .B2(n8668), .A(n9700), .ZN(n8561) );
  AOI21_X1 U9958 ( .B1(n8585), .B2(n9214), .A(n8561), .ZN(n8562) );
  OAI21_X1 U9959 ( .B1(n8563), .B2(n9223), .A(n8562), .ZN(n8564) );
  AOI21_X1 U9960 ( .B1(n9499), .B2(n8590), .A(n8564), .ZN(n8565) );
  OAI21_X1 U9961 ( .B1(n8566), .B2(n8592), .A(n8565), .ZN(P1_U3236) );
  INV_X1 U9962 ( .A(n9316), .ZN(n9087) );
  OAI21_X1 U9963 ( .B1(n8569), .B2(n8568), .A(n8567), .ZN(n8570) );
  NAND3_X1 U9964 ( .A1(n4275), .A2(n8571), .A3(n8570), .ZN(n8577) );
  OAI22_X1 U9965 ( .A1(n8999), .A2(n8573), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8572), .ZN(n8575) );
  NOR2_X1 U9966 ( .A1(n9007), .A2(n8588), .ZN(n8574) );
  AOI211_X1 U9967 ( .C1(n9085), .C2(n8583), .A(n8575), .B(n8574), .ZN(n8576)
         );
  OAI211_X1 U9968 ( .C1(n9087), .C2(n8578), .A(n8577), .B(n8576), .ZN(P1_U3238) );
  NAND2_X1 U9969 ( .A1(n8579), .A2(n8580), .ZN(n8581) );
  XOR2_X1 U9970 ( .A(n8582), .B(n8581), .Z(n8593) );
  NAND2_X1 U9971 ( .A1(n8583), .A2(n9272), .ZN(n8587) );
  AOI21_X1 U9972 ( .B1(n8585), .B2(n9266), .A(n8584), .ZN(n8586) );
  OAI211_X1 U9973 ( .C1(n8645), .C2(n8588), .A(n8587), .B(n8586), .ZN(n8589)
         );
  AOI21_X1 U9974 ( .B1(n9514), .B2(n8590), .A(n8589), .ZN(n8591) );
  OAI21_X1 U9975 ( .B1(n8593), .B2(n8592), .A(n8591), .ZN(P1_U3239) );
  NAND2_X1 U9976 ( .A1(n8873), .A2(n8705), .ZN(n8713) );
  NAND2_X1 U9977 ( .A1(n8595), .A2(n8605), .ZN(n8598) );
  OR2_X1 U9978 ( .A1(n8608), .A2(n8596), .ZN(n8597) );
  NAND2_X1 U9979 ( .A1(n8599), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8603) );
  NAND2_X1 U9980 ( .A1(n5686), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8602) );
  NAND2_X1 U9981 ( .A1(n8600), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8601) );
  AND3_X1 U9982 ( .A1(n8603), .A2(n8602), .A3(n8601), .ZN(n9036) );
  NOR2_X1 U9983 ( .A1(n9585), .A2(n9036), .ZN(n8751) );
  NAND2_X1 U9984 ( .A1(n8973), .A2(n8751), .ZN(n8604) );
  NAND2_X1 U9985 ( .A1(n8606), .A2(n8605), .ZN(n8610) );
  OR2_X1 U9986 ( .A1(n8608), .A2(n8607), .ZN(n8609) );
  NAND2_X1 U9987 ( .A1(n9307), .A2(n9035), .ZN(n9031) );
  NAND2_X1 U9988 ( .A1(n9311), .A2(n9007), .ZN(n8769) );
  MUX2_X1 U9989 ( .A(n8824), .B(n8769), .S(n8705), .Z(n8701) );
  OR2_X1 U9990 ( .A1(n9327), .A2(n8996), .ZN(n8783) );
  NAND2_X1 U9991 ( .A1(n9327), .A2(n8996), .ZN(n9025) );
  INV_X1 U9992 ( .A(n9121), .ZN(n9157) );
  NAND2_X1 U9993 ( .A1(n9473), .A2(n9157), .ZN(n9024) );
  NAND2_X1 U9994 ( .A1(n9115), .A2(n9024), .ZN(n9130) );
  INV_X1 U9995 ( .A(n9130), .ZN(n8747) );
  NAND2_X1 U9996 ( .A1(n9118), .A2(n8747), .ZN(n8612) );
  NAND3_X1 U9997 ( .A1(n9025), .A2(n8705), .A3(n9024), .ZN(n8611) );
  NAND2_X1 U9998 ( .A1(n8612), .A2(n8611), .ZN(n8689) );
  NAND3_X1 U9999 ( .A1(n8613), .A2(n8850), .A3(n8619), .ZN(n8614) );
  INV_X1 U10000 ( .A(n8852), .ZN(n8615) );
  OR2_X1 U10001 ( .A1(n8847), .A2(n8615), .ZN(n8794) );
  INV_X1 U10002 ( .A(n8795), .ZN(n8618) );
  NAND2_X1 U10003 ( .A1(n8849), .A2(n8848), .ZN(n8616) );
  NAND3_X1 U10004 ( .A1(n8616), .A2(n8795), .A3(n8852), .ZN(n8617) );
  AND2_X1 U10005 ( .A1(n8617), .A2(n8851), .ZN(n8802) );
  OAI211_X1 U10006 ( .C1(n8794), .C2(n8618), .A(n8729), .B(n8802), .ZN(n8620)
         );
  AND2_X1 U10007 ( .A1(n8798), .A2(n8796), .ZN(n8800) );
  NAND2_X1 U10008 ( .A1(n8631), .A2(n8619), .ZN(n8792) );
  AOI21_X1 U10009 ( .B1(n8620), .B2(n8800), .A(n8792), .ZN(n8629) );
  INV_X1 U10010 ( .A(n8705), .ZN(n8714) );
  NAND2_X1 U10011 ( .A1(n8621), .A2(n8714), .ZN(n8626) );
  INV_X1 U10012 ( .A(n8626), .ZN(n8628) );
  AND2_X1 U10013 ( .A1(n8714), .A2(n8893), .ZN(n8624) );
  OAI21_X1 U10014 ( .B1(n8714), .B2(n8893), .A(n8623), .ZN(n8622) );
  OAI21_X1 U10015 ( .B1(n8624), .B2(n8623), .A(n8622), .ZN(n8625) );
  OAI21_X1 U10016 ( .B1(n8626), .B2(n8805), .A(n8625), .ZN(n8627) );
  AOI21_X1 U10017 ( .B1(n8629), .B2(n8628), .A(n8627), .ZN(n8630) );
  NAND2_X1 U10018 ( .A1(n8632), .A2(n8736), .ZN(n8636) );
  MUX2_X1 U10019 ( .A(n8634), .B(n8633), .S(n8714), .Z(n8635) );
  NAND3_X1 U10020 ( .A1(n8636), .A2(n8737), .A3(n8635), .ZN(n8650) );
  AND2_X1 U10021 ( .A1(n8811), .A2(n8637), .ZN(n8638) );
  AND2_X1 U10022 ( .A1(n9009), .A2(n8638), .ZN(n8790) );
  OR2_X1 U10023 ( .A1(n9521), .A2(n8985), .ZN(n9011) );
  NAND2_X1 U10024 ( .A1(n9011), .A2(n8639), .ZN(n8816) );
  AOI21_X1 U10025 ( .B1(n8650), .B2(n8790), .A(n8816), .ZN(n8644) );
  INV_X1 U10026 ( .A(n8811), .ZN(n8642) );
  INV_X1 U10027 ( .A(n8640), .ZN(n8641) );
  MUX2_X1 U10028 ( .A(n8642), .B(n8641), .S(n8714), .Z(n8651) );
  NAND2_X1 U10029 ( .A1(n8651), .A2(n9009), .ZN(n8643) );
  AND2_X1 U10030 ( .A1(n9521), .A2(n8985), .ZN(n8789) );
  AOI21_X1 U10031 ( .B1(n8644), .B2(n8643), .A(n8789), .ZN(n8647) );
  OR2_X1 U10032 ( .A1(n9514), .A2(n9285), .ZN(n8648) );
  NAND2_X1 U10033 ( .A1(n9514), .A2(n9285), .ZN(n8788) );
  OR2_X1 U10034 ( .A1(n9511), .A2(n8645), .ZN(n8660) );
  NAND2_X1 U10035 ( .A1(n9511), .A2(n8645), .ZN(n9013) );
  NAND2_X1 U10036 ( .A1(n8660), .A2(n9013), .ZN(n9249) );
  INV_X1 U10037 ( .A(n9249), .ZN(n8646) );
  OAI211_X1 U10038 ( .C1(n8647), .C2(n9264), .A(n8646), .B(n8788), .ZN(n8659)
         );
  AND2_X1 U10039 ( .A1(n8660), .A2(n8648), .ZN(n8818) );
  INV_X1 U10040 ( .A(n8810), .ZN(n8649) );
  NAND2_X1 U10041 ( .A1(n8650), .A2(n8649), .ZN(n8653) );
  INV_X1 U10042 ( .A(n8651), .ZN(n8652) );
  INV_X1 U10043 ( .A(n8816), .ZN(n8654) );
  INV_X1 U10044 ( .A(n8789), .ZN(n8655) );
  NAND3_X1 U10045 ( .A1(n8656), .A2(n8988), .A3(n8655), .ZN(n8657) );
  NAND2_X1 U10046 ( .A1(n8818), .A2(n8657), .ZN(n8658) );
  MUX2_X1 U10047 ( .A(n8660), .B(n9013), .S(n8705), .Z(n8661) );
  NAND2_X1 U10048 ( .A1(n8662), .A2(n8661), .ZN(n8665) );
  INV_X1 U10049 ( .A(n9242), .ZN(n9207) );
  NAND2_X1 U10050 ( .A1(n9499), .A2(n9207), .ZN(n8787) );
  NAND2_X1 U10051 ( .A1(n9504), .A2(n9252), .ZN(n9015) );
  OAI211_X1 U10052 ( .C1(n8665), .C2(n9214), .A(n8787), .B(n9015), .ZN(n8664)
         );
  OR2_X1 U10053 ( .A1(n9499), .A2(n9207), .ZN(n8723) );
  OR2_X1 U10054 ( .A1(n9504), .A2(n9252), .ZN(n9211) );
  AND2_X1 U10055 ( .A1(n8723), .A2(n9211), .ZN(n9017) );
  OAI21_X1 U10056 ( .B1(n8665), .B2(n9504), .A(n9017), .ZN(n8663) );
  INV_X1 U10057 ( .A(n8665), .ZN(n8666) );
  AND2_X1 U10058 ( .A1(n9504), .A2(n9214), .ZN(n8989) );
  NAND2_X1 U10059 ( .A1(n8666), .A2(n8989), .ZN(n8667) );
  NAND3_X1 U10060 ( .A1(n8670), .A2(n8779), .A3(n8723), .ZN(n8669) );
  AND2_X1 U10061 ( .A1(n9487), .A2(n9208), .ZN(n9161) );
  NAND2_X1 U10062 ( .A1(n9493), .A2(n8668), .ZN(n8722) );
  INV_X1 U10063 ( .A(n8722), .ZN(n9018) );
  NOR2_X1 U10064 ( .A1(n9161), .A2(n9018), .ZN(n8777) );
  NAND2_X1 U10065 ( .A1(n8669), .A2(n8777), .ZN(n8673) );
  NAND3_X1 U10066 ( .A1(n8670), .A2(n8787), .A3(n8722), .ZN(n8671) );
  AOI21_X1 U10067 ( .B1(n8671), .B2(n8779), .A(n9161), .ZN(n8672) );
  INV_X1 U10068 ( .A(n8674), .ZN(n8676) );
  NAND2_X1 U10069 ( .A1(n9483), .A2(n9156), .ZN(n9021) );
  OR2_X1 U10070 ( .A1(n9483), .A2(n9156), .ZN(n8675) );
  NAND2_X1 U10071 ( .A1(n9021), .A2(n8675), .ZN(n9163) );
  NOR2_X1 U10072 ( .A1(n9487), .A2(n9208), .ZN(n9019) );
  NOR2_X1 U10073 ( .A1(n9163), .A2(n9019), .ZN(n8677) );
  NAND2_X1 U10074 ( .A1(n8676), .A2(n8677), .ZN(n8686) );
  INV_X1 U10075 ( .A(n8677), .ZN(n8678) );
  NAND2_X1 U10076 ( .A1(n8678), .A2(n9021), .ZN(n8679) );
  OR2_X1 U10077 ( .A1(n9479), .A2(n8680), .ZN(n8721) );
  AND2_X1 U10078 ( .A1(n8679), .A2(n8721), .ZN(n8775) );
  NAND2_X1 U10079 ( .A1(n8686), .A2(n8775), .ZN(n8681) );
  NAND2_X1 U10080 ( .A1(n9479), .A2(n8680), .ZN(n9022) );
  NAND2_X1 U10081 ( .A1(n8681), .A2(n9022), .ZN(n8685) );
  INV_X1 U10082 ( .A(n9024), .ZN(n8682) );
  NAND2_X1 U10083 ( .A1(n8783), .A2(n8682), .ZN(n8683) );
  AND2_X1 U10084 ( .A1(n8683), .A2(n9025), .ZN(n8684) );
  NAND2_X1 U10085 ( .A1(n9321), .A2(n8999), .ZN(n9026) );
  NAND2_X1 U10086 ( .A1(n8684), .A2(n9026), .ZN(n8865) );
  AOI21_X1 U10087 ( .B1(n8689), .B2(n8685), .A(n8865), .ZN(n8692) );
  NAND3_X1 U10088 ( .A1(n8686), .A2(n9021), .A3(n9022), .ZN(n8687) );
  NAND3_X1 U10089 ( .A1(n8687), .A2(n9115), .A3(n8721), .ZN(n8690) );
  NAND2_X1 U10090 ( .A1(n9027), .A2(n8783), .ZN(n8688) );
  AOI21_X1 U10091 ( .B1(n8690), .B2(n8689), .A(n8688), .ZN(n8691) );
  MUX2_X1 U10092 ( .A(n8692), .B(n8691), .S(n8705), .Z(n8699) );
  NOR2_X1 U10093 ( .A1(n9316), .A2(n9105), .ZN(n9001) );
  NAND2_X1 U10094 ( .A1(n9316), .A2(n9105), .ZN(n9003) );
  INV_X1 U10095 ( .A(n9003), .ZN(n8693) );
  MUX2_X1 U10096 ( .A(n9027), .B(n9026), .S(n8705), .Z(n8694) );
  NAND2_X1 U10097 ( .A1(n9089), .A2(n8694), .ZN(n8698) );
  INV_X1 U10098 ( .A(n9105), .ZN(n8695) );
  NAND2_X1 U10099 ( .A1(n9316), .A2(n8695), .ZN(n9028) );
  NOR2_X1 U10100 ( .A1(n9316), .A2(n8695), .ZN(n9029) );
  MUX2_X1 U10101 ( .A(n4669), .B(n9029), .S(n8705), .Z(n8696) );
  INV_X1 U10102 ( .A(n8696), .ZN(n8697) );
  OAI211_X1 U10103 ( .C1(n8699), .C2(n8698), .A(n9076), .B(n8697), .ZN(n8700)
         );
  MUX2_X1 U10104 ( .A(n9031), .B(n8767), .S(n8705), .Z(n8702) );
  NAND2_X1 U10105 ( .A1(n8703), .A2(n8702), .ZN(n8704) );
  INV_X1 U10106 ( .A(n8704), .ZN(n8711) );
  INV_X1 U10107 ( .A(n9062), .ZN(n8770) );
  NAND3_X1 U10108 ( .A1(n8704), .A2(n8770), .A3(n9299), .ZN(n8708) );
  NAND2_X1 U10109 ( .A1(n9062), .A2(n8705), .ZN(n8707) );
  NAND2_X1 U10110 ( .A1(n8771), .A2(n8714), .ZN(n8706) );
  NAND3_X1 U10111 ( .A1(n8708), .A2(n8707), .A3(n8706), .ZN(n8709) );
  NOR2_X1 U10112 ( .A1(n8834), .A2(n8709), .ZN(n8710) );
  INV_X1 U10113 ( .A(n9036), .ZN(n8887) );
  NAND2_X1 U10114 ( .A1(n8887), .A2(n8717), .ZN(n8712) );
  NAND2_X1 U10115 ( .A1(n9585), .A2(n8712), .ZN(n8830) );
  NAND2_X1 U10116 ( .A1(n8834), .A2(n8714), .ZN(n8715) );
  NAND2_X1 U10117 ( .A1(n8716), .A2(n8715), .ZN(n8766) );
  INV_X1 U10118 ( .A(n8766), .ZN(n8763) );
  NAND2_X1 U10119 ( .A1(n4525), .A2(n8717), .ZN(n8764) );
  INV_X1 U10120 ( .A(n8718), .ZN(n8719) );
  AND2_X1 U10121 ( .A1(n8764), .A2(n8719), .ZN(n8762) );
  NAND2_X1 U10122 ( .A1(n9585), .A2(n9036), .ZN(n8720) );
  AND2_X1 U10123 ( .A1(n8764), .A2(n8720), .ZN(n8872) );
  XNOR2_X1 U10124 ( .A(n8771), .B(n9062), .ZN(n9033) );
  NAND2_X1 U10125 ( .A1(n9027), .A2(n9026), .ZN(n9104) );
  NAND2_X1 U10126 ( .A1(n8721), .A2(n9022), .ZN(n9153) );
  INV_X1 U10127 ( .A(n9153), .ZN(n9142) );
  XNOR2_X1 U10128 ( .A(n9487), .B(n9208), .ZN(n9184) );
  INV_X1 U10129 ( .A(n8841), .ZN(n8724) );
  NOR2_X1 U10130 ( .A1(n8725), .A2(n8724), .ZN(n9750) );
  INV_X1 U10131 ( .A(n9721), .ZN(n9711) );
  AND4_X1 U10132 ( .A1(n9750), .A2(n9711), .A3(n8726), .A4(n8844), .ZN(n8730)
         );
  AND4_X1 U10133 ( .A1(n8730), .A2(n8729), .A3(n8728), .A4(n8727), .ZN(n8734)
         );
  AND4_X1 U10134 ( .A1(n8734), .A2(n8733), .A3(n8732), .A4(n8731), .ZN(n8735)
         );
  NAND4_X1 U10135 ( .A1(n8738), .A2(n8737), .A3(n8736), .A4(n8735), .ZN(n8739)
         );
  NOR2_X1 U10136 ( .A1(n8740), .A2(n8739), .ZN(n8742) );
  XNOR2_X1 U10137 ( .A(n9521), .B(n8985), .ZN(n9281) );
  INV_X1 U10138 ( .A(n9281), .ZN(n8741) );
  NAND3_X1 U10139 ( .A1(n8988), .A2(n8742), .A3(n8741), .ZN(n8743) );
  NOR2_X1 U10140 ( .A1(n9249), .A2(n8743), .ZN(n8744) );
  NAND4_X1 U10141 ( .A1(n9194), .A2(n9218), .A3(n9241), .A4(n8744), .ZN(n8745)
         );
  NOR3_X1 U10142 ( .A1(n9163), .A2(n9184), .A3(n8745), .ZN(n8746) );
  NAND4_X1 U10143 ( .A1(n9118), .A2(n8747), .A3(n9142), .A4(n8746), .ZN(n8748)
         );
  NOR2_X1 U10144 ( .A1(n9104), .A2(n8748), .ZN(n8749) );
  AND2_X1 U10145 ( .A1(n9089), .A2(n8749), .ZN(n8750) );
  AND4_X1 U10146 ( .A1(n9033), .A2(n9030), .A3(n9076), .A4(n8750), .ZN(n8752)
         );
  INV_X1 U10147 ( .A(n8751), .ZN(n8869) );
  NAND4_X1 U10148 ( .A1(n8872), .A2(n8752), .A3(n8873), .A4(n8869), .ZN(n8754)
         );
  NAND2_X1 U10149 ( .A1(n8754), .A2(n8753), .ZN(n8836) );
  OR2_X1 U10150 ( .A1(n9765), .A2(n8755), .ZN(n8756) );
  OR2_X1 U10151 ( .A1(n8757), .A2(n8756), .ZN(n8760) );
  INV_X1 U10152 ( .A(n8839), .ZN(n8758) );
  AOI21_X1 U10153 ( .B1(n5639), .B2(n8758), .A(n8974), .ZN(n8759) );
  NAND2_X1 U10154 ( .A1(n8760), .A2(n8759), .ZN(n8878) );
  NAND4_X1 U10155 ( .A1(n8836), .A2(n9744), .A3(n8837), .A4(n8878), .ZN(n8761)
         );
  NAND2_X1 U10156 ( .A1(n8764), .A2(n4246), .ZN(n8831) );
  NOR2_X1 U10157 ( .A1(n8831), .A2(n6206), .ZN(n8765) );
  NAND2_X1 U10158 ( .A1(n8766), .A2(n8765), .ZN(n8885) );
  OR2_X1 U10159 ( .A1(n8771), .A2(n8770), .ZN(n8768) );
  NAND2_X1 U10160 ( .A1(n8768), .A2(n8767), .ZN(n8827) );
  INV_X1 U10161 ( .A(n8827), .ZN(n8774) );
  INV_X1 U10162 ( .A(n8824), .ZN(n9059) );
  OAI211_X1 U10163 ( .C1(n9059), .C2(n9028), .A(n9031), .B(n8769), .ZN(n8773)
         );
  AND2_X1 U10164 ( .A1(n8771), .A2(n8770), .ZN(n8772) );
  AOI21_X1 U10165 ( .B1(n8774), .B2(n8773), .A(n8772), .ZN(n8867) );
  INV_X1 U10166 ( .A(n8775), .ZN(n8776) );
  NAND2_X1 U10167 ( .A1(n8776), .A2(n9022), .ZN(n8782) );
  AND2_X1 U10168 ( .A1(n8777), .A2(n9021), .ZN(n8778) );
  AND2_X1 U10169 ( .A1(n8778), .A2(n9022), .ZN(n8785) );
  INV_X1 U10170 ( .A(n8787), .ZN(n9016) );
  OAI21_X1 U10171 ( .B1(n9017), .B2(n9016), .A(n8779), .ZN(n8780) );
  NAND2_X1 U10172 ( .A1(n8785), .A2(n8780), .ZN(n8781) );
  AND3_X1 U10173 ( .A1(n8782), .A2(n9115), .A3(n8781), .ZN(n8784) );
  NAND2_X1 U10174 ( .A1(n8784), .A2(n8783), .ZN(n8863) );
  INV_X1 U10175 ( .A(n8785), .ZN(n8861) );
  AND2_X1 U10176 ( .A1(n9015), .A2(n9013), .ZN(n8786) );
  NAND2_X1 U10177 ( .A1(n8787), .A2(n8786), .ZN(n8817) );
  INV_X1 U10178 ( .A(n8788), .ZN(n9012) );
  OR3_X1 U10179 ( .A1(n8817), .A2(n9012), .A3(n8789), .ZN(n8820) );
  INV_X1 U10180 ( .A(n8790), .ZN(n8814) );
  INV_X1 U10181 ( .A(n8809), .ZN(n8791) );
  OR3_X1 U10182 ( .A1(n8814), .A2(n8792), .A3(n8791), .ZN(n8793) );
  NOR2_X1 U10183 ( .A1(n8820), .A2(n8793), .ZN(n8855) );
  INV_X1 U10184 ( .A(n8794), .ZN(n8804) );
  NAND2_X1 U10185 ( .A1(n8796), .A2(n8795), .ZN(n8797) );
  NAND2_X1 U10186 ( .A1(n8797), .A2(n8850), .ZN(n8799) );
  AND2_X1 U10187 ( .A1(n8799), .A2(n8798), .ZN(n8854) );
  INV_X1 U10188 ( .A(n8800), .ZN(n8801) );
  AOI21_X1 U10189 ( .B1(n8802), .B2(n8850), .A(n8801), .ZN(n8803) );
  AOI21_X1 U10190 ( .B1(n8804), .B2(n8854), .A(n8803), .ZN(n8821) );
  NAND2_X1 U10191 ( .A1(n8806), .A2(n8805), .ZN(n8808) );
  AOI21_X1 U10192 ( .B1(n8809), .B2(n8808), .A(n8807), .ZN(n8813) );
  NAND3_X1 U10193 ( .A1(n9009), .A2(n8811), .A3(n8810), .ZN(n8812) );
  OAI21_X1 U10194 ( .B1(n8814), .B2(n8813), .A(n8812), .ZN(n8815) );
  NOR2_X1 U10195 ( .A1(n8816), .A2(n8815), .ZN(n8819) );
  OAI22_X1 U10196 ( .A1(n8820), .A2(n8819), .B1(n8818), .B2(n8817), .ZN(n8840)
         );
  AOI21_X1 U10197 ( .B1(n8855), .B2(n8821), .A(n8840), .ZN(n8822) );
  NOR2_X1 U10198 ( .A1(n8861), .A2(n8822), .ZN(n8823) );
  NOR2_X1 U10199 ( .A1(n8863), .A2(n8823), .ZN(n8828) );
  INV_X1 U10200 ( .A(n9029), .ZN(n8825) );
  NAND3_X1 U10201 ( .A1(n8825), .A2(n8824), .A3(n9027), .ZN(n8826) );
  NOR2_X1 U10202 ( .A1(n8827), .A2(n8826), .ZN(n8864) );
  OAI21_X1 U10203 ( .B1(n8828), .B2(n8865), .A(n8864), .ZN(n8829) );
  AND3_X1 U10204 ( .A1(n8830), .A2(n8867), .A3(n8829), .ZN(n8833) );
  INV_X1 U10205 ( .A(n8831), .ZN(n8832) );
  OAI21_X1 U10206 ( .B1(n8834), .B2(n8833), .A(n8832), .ZN(n8835) );
  NAND2_X1 U10207 ( .A1(n8836), .A2(n8835), .ZN(n8838) );
  NAND4_X1 U10208 ( .A1(n8838), .A2(n8837), .A3(n5638), .A4(n8878), .ZN(n8883)
         );
  NAND2_X1 U10209 ( .A1(n8878), .A2(n8839), .ZN(n8882) );
  INV_X1 U10210 ( .A(n8840), .ZN(n8859) );
  AND2_X1 U10211 ( .A1(n8841), .A2(n4246), .ZN(n8845) );
  NAND4_X1 U10212 ( .A1(n8845), .A2(n8844), .A3(n8843), .A4(n8842), .ZN(n8846)
         );
  NAND4_X1 U10213 ( .A1(n8849), .A2(n8848), .A3(n8847), .A4(n8846), .ZN(n8853)
         );
  AOI211_X1 U10214 ( .C1(n8853), .C2(n8852), .A(n4646), .B(n4647), .ZN(n8857)
         );
  INV_X1 U10215 ( .A(n8854), .ZN(n8856) );
  OAI21_X1 U10216 ( .B1(n8857), .B2(n8856), .A(n8855), .ZN(n8858) );
  AND2_X1 U10217 ( .A1(n8859), .A2(n8858), .ZN(n8860) );
  NOR2_X1 U10218 ( .A1(n8861), .A2(n8860), .ZN(n8862) );
  NOR2_X1 U10219 ( .A1(n8863), .A2(n8862), .ZN(n8866) );
  OAI21_X1 U10220 ( .B1(n8866), .B2(n8865), .A(n8864), .ZN(n8868) );
  NAND2_X1 U10221 ( .A1(n8868), .A2(n8867), .ZN(n8870) );
  NAND2_X1 U10222 ( .A1(n8870), .A2(n8869), .ZN(n8871) );
  NAND2_X1 U10223 ( .A1(n8872), .A2(n8871), .ZN(n8874) );
  AND2_X1 U10224 ( .A1(n8874), .A2(n8873), .ZN(n8879) );
  INV_X1 U10225 ( .A(n8879), .ZN(n8876) );
  NAND3_X1 U10226 ( .A1(n8876), .A2(n8875), .A3(n8878), .ZN(n8881) );
  NAND4_X1 U10227 ( .A1(n8879), .A2(n9744), .A3(n8878), .A4(n8877), .ZN(n8880)
         );
  NAND4_X1 U10228 ( .A1(n8883), .A2(n8882), .A3(n8881), .A4(n8880), .ZN(n8884)
         );
  AOI21_X1 U10229 ( .B1(n8886), .B2(n8885), .A(n8884), .ZN(P1_U3240) );
  MUX2_X1 U10230 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n8887), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10231 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9062), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10232 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9078), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10233 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9090), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10234 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9105), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10235 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9120), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10236 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9127), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10237 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9121), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10238 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9167), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10239 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9186), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10240 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9168), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10241 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9215), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10242 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9242), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10243 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9214), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10244 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9265), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10245 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n8888), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10246 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9266), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10247 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8889), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10248 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8890), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10249 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n8891), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10250 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n8892), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10251 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n8893), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10252 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n8894), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10253 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8895), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10254 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8896), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10255 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n8897), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10256 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n8898), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10257 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n8899), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10258 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9755), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10259 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n8900), .S(P1_U4006), .Z(
        P1_U3556) );
  NAND2_X1 U10260 ( .A1(n9706), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n8912) );
  NOR2_X1 U10261 ( .A1(n8901), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8902) );
  AOI21_X1 U10262 ( .B1(n9699), .B2(n5651), .A(n8902), .ZN(n8911) );
  OAI211_X1 U10263 ( .C1(n8905), .C2(n8904), .A(n9697), .B(n8903), .ZN(n8910)
         );
  OAI211_X1 U10264 ( .C1(n8908), .C2(n8907), .A(n9707), .B(n8906), .ZN(n8909)
         );
  NAND4_X1 U10265 ( .A1(n8912), .A2(n8911), .A3(n8910), .A4(n8909), .ZN(
        P1_U3242) );
  NAND2_X1 U10266 ( .A1(n9706), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n8924) );
  AOI21_X1 U10267 ( .B1(n9699), .B2(n8914), .A(n8913), .ZN(n8923) );
  OAI211_X1 U10268 ( .C1(n8917), .C2(n8916), .A(n9697), .B(n8915), .ZN(n8922)
         );
  OAI211_X1 U10269 ( .C1(n8920), .C2(n8919), .A(n9707), .B(n8918), .ZN(n8921)
         );
  NAND4_X1 U10270 ( .A1(n8924), .A2(n8923), .A3(n8922), .A4(n8921), .ZN(
        P1_U3244) );
  OAI21_X1 U10271 ( .B1(n8927), .B2(n8926), .A(n8925), .ZN(n8932) );
  AOI211_X1 U10272 ( .C1(n8930), .C2(n8929), .A(n8928), .B(n9679), .ZN(n8931)
         );
  AOI21_X1 U10273 ( .B1(n9707), .B2(n8932), .A(n8931), .ZN(n8938) );
  INV_X1 U10274 ( .A(n8933), .ZN(n8937) );
  NAND2_X1 U10275 ( .A1(n9706), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n8936) );
  NAND2_X1 U10276 ( .A1(n9699), .A2(n8934), .ZN(n8935) );
  NAND4_X1 U10277 ( .A1(n8938), .A2(n8937), .A3(n8936), .A4(n8935), .ZN(
        P1_U3253) );
  AOI21_X1 U10278 ( .B1(n8944), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8939), .ZN(
        n8942) );
  NAND2_X1 U10279 ( .A1(n8962), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8940) );
  OAI21_X1 U10280 ( .B1(n8962), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8940), .ZN(
        n8941) );
  NOR2_X1 U10281 ( .A1(n8942), .A2(n8941), .ZN(n8955) );
  AOI211_X1 U10282 ( .C1(n8942), .C2(n8941), .A(n8955), .B(n9679), .ZN(n8948)
         );
  AOI21_X1 U10283 ( .B1(n8944), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8943), .ZN(
        n8946) );
  XNOR2_X1 U10284 ( .A(n8962), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n8945) );
  NOR2_X1 U10285 ( .A1(n8946), .A2(n8945), .ZN(n8961) );
  AOI211_X1 U10286 ( .C1(n8946), .C2(n8945), .A(n8961), .B(n9648), .ZN(n8947)
         );
  NOR2_X1 U10287 ( .A1(n8948), .A2(n8947), .ZN(n8951) );
  INV_X1 U10288 ( .A(n8949), .ZN(n8950) );
  OAI211_X1 U10289 ( .C1(n8952), .C2(n9687), .A(n8951), .B(n8950), .ZN(n8953)
         );
  AOI21_X1 U10290 ( .B1(n9706), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n8953), .ZN(
        n8954) );
  INV_X1 U10291 ( .A(n8954), .ZN(P1_U3258) );
  OR2_X1 U10292 ( .A1(n9698), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8957) );
  NAND2_X1 U10293 ( .A1(n9698), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8956) );
  NAND2_X1 U10294 ( .A1(n8957), .A2(n8956), .ZN(n9695) );
  NOR2_X1 U10295 ( .A1(n9694), .A2(n9695), .ZN(n9693) );
  AOI21_X1 U10296 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9698), .A(n9693), .ZN(
        n8958) );
  XNOR2_X1 U10297 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n8958), .ZN(n8968) );
  INV_X1 U10298 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8960) );
  AOI22_X1 U10299 ( .A1(n9698), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n8960), .B2(
        n8959), .ZN(n9705) );
  AOI21_X1 U10300 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n8962), .A(n8961), .ZN(
        n9704) );
  NAND2_X1 U10301 ( .A1(n9705), .A2(n9704), .ZN(n9703) );
  OAI21_X1 U10302 ( .B1(n9698), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9703), .ZN(
        n8963) );
  XNOR2_X1 U10303 ( .A(n8963), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n8964) );
  AOI22_X1 U10304 ( .A1(n8968), .A2(n9697), .B1(n9707), .B2(n8964), .ZN(n8970)
         );
  INV_X1 U10305 ( .A(n8964), .ZN(n8969) );
  INV_X1 U10306 ( .A(n8965), .ZN(n8967) );
  NAND2_X1 U10307 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3084), .ZN(n8971) );
  INV_X1 U10308 ( .A(n9321), .ZN(n9102) );
  INV_X1 U10309 ( .A(n9479), .ZN(n9147) );
  INV_X1 U10310 ( .A(n9483), .ZN(n9174) );
  INV_X1 U10311 ( .A(n9499), .ZN(n9227) );
  NAND2_X1 U10312 ( .A1(n9147), .A2(n9170), .ZN(n9144) );
  NOR2_X2 U10313 ( .A1(n9327), .A2(n9136), .ZN(n9111) );
  NAND2_X1 U10314 ( .A1(n9102), .A2(n9111), .ZN(n9096) );
  NOR2_X2 U10315 ( .A1(n9096), .A2(n9316), .ZN(n9084) );
  NOR2_X1 U10316 ( .A1(n9585), .A2(n9041), .ZN(n8972) );
  XNOR2_X1 U10317 ( .A(n8973), .B(n8972), .ZN(n9564) );
  NAND2_X1 U10318 ( .A1(n9564), .A2(n9718), .ZN(n8980) );
  OR2_X1 U10319 ( .A1(n8975), .A2(n8974), .ZN(n8976) );
  NAND2_X1 U10320 ( .A1(n9756), .A2(n8976), .ZN(n9037) );
  NOR2_X1 U10321 ( .A1(n9037), .A2(n8977), .ZN(n9584) );
  INV_X1 U10322 ( .A(n9584), .ZN(n8978) );
  NOR2_X1 U10323 ( .A1(n9234), .A2(n8978), .ZN(n8981) );
  AOI21_X1 U10324 ( .B1(n9234), .B2(P1_REG2_REG_31__SCAN_IN), .A(n8981), .ZN(
        n8979) );
  OAI211_X1 U10325 ( .C1(n4525), .C2(n9733), .A(n8980), .B(n8979), .ZN(
        P1_U3261) );
  INV_X1 U10326 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9425) );
  NOR2_X1 U10327 ( .A1(n9762), .A2(n9425), .ZN(n8982) );
  AOI211_X1 U10328 ( .C1(n9585), .C2(n9226), .A(n8982), .B(n8981), .ZN(n8983)
         );
  OAI21_X1 U10329 ( .B1(n9582), .B2(n9042), .A(n8983), .ZN(P1_U3262) );
  NAND2_X1 U10330 ( .A1(n8984), .A2(n4802), .ZN(n9280) );
  NAND2_X1 U10331 ( .A1(n9294), .A2(n8985), .ZN(n8987) );
  AOI21_X2 U10332 ( .B1(n9280), .B2(n8987), .A(n8986), .ZN(n9261) );
  INV_X1 U10333 ( .A(n9514), .ZN(n9274) );
  OR2_X2 U10334 ( .A1(n9217), .A2(n8990), .ZN(n9191) );
  NAND2_X1 U10335 ( .A1(n9493), .A2(n9215), .ZN(n8992) );
  INV_X1 U10336 ( .A(n9487), .ZN(n9183) );
  INV_X1 U10337 ( .A(n9143), .ZN(n8994) );
  AOI21_X1 U10338 ( .B1(n8994), .B2(n9153), .A(n8993), .ZN(n9131) );
  NAND2_X1 U10339 ( .A1(n9131), .A2(n9130), .ZN(n9129) );
  NAND2_X1 U10340 ( .A1(n9129), .A2(n8995), .ZN(n9110) );
  NAND2_X1 U10341 ( .A1(n9110), .A2(n4798), .ZN(n8998) );
  NAND2_X1 U10342 ( .A1(n9102), .A2(n8999), .ZN(n9000) );
  INV_X1 U10343 ( .A(n9001), .ZN(n9002) );
  NAND2_X1 U10344 ( .A1(n9004), .A2(n9003), .ZN(n9069) );
  INV_X1 U10345 ( .A(n9069), .ZN(n9006) );
  INV_X1 U10346 ( .A(n9076), .ZN(n9005) );
  OAI21_X1 U10347 ( .B1(n9035), .B2(n4513), .A(n9050), .ZN(n9008) );
  XNOR2_X1 U10348 ( .A(n9008), .B(n9033), .ZN(n9298) );
  INV_X1 U10349 ( .A(n9298), .ZN(n9049) );
  NAND2_X1 U10350 ( .A1(n9010), .A2(n9009), .ZN(n9282) );
  INV_X1 U10351 ( .A(n9013), .ZN(n9014) );
  INV_X1 U10352 ( .A(n9163), .ZN(n9020) );
  INV_X1 U10353 ( .A(n9022), .ZN(n9023) );
  AOI21_X1 U10354 ( .B1(n9154), .B2(n9142), .A(n9023), .ZN(n9126) );
  NAND2_X1 U10355 ( .A1(n9126), .A2(n9024), .ZN(n9116) );
  NAND3_X1 U10356 ( .A1(n9116), .A2(n9118), .A3(n9115), .ZN(n9117) );
  INV_X1 U10357 ( .A(n9031), .ZN(n9032) );
  OAI21_X1 U10358 ( .B1(n9052), .B2(n9299), .A(n9041), .ZN(n9300) );
  NOR2_X1 U10359 ( .A1(n9300), .A2(n9042), .ZN(n9047) );
  INV_X1 U10360 ( .A(n9043), .ZN(n9044) );
  AOI22_X1 U10361 ( .A1(n9044), .A2(n9747), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9234), .ZN(n9045) );
  OAI21_X1 U10362 ( .B1(n9299), .B2(n9733), .A(n9045), .ZN(n9046) );
  AOI211_X1 U10363 ( .C1(n9302), .C2(n9762), .A(n9047), .B(n9046), .ZN(n9048)
         );
  OAI21_X1 U10364 ( .B1(n9049), .B2(n9297), .A(n9048), .ZN(P1_U3355) );
  OAI21_X1 U10365 ( .B1(n9051), .B2(n9058), .A(n9050), .ZN(n9305) );
  AOI211_X1 U10366 ( .C1(n9307), .C2(n9070), .A(n9819), .B(n9052), .ZN(n9306)
         );
  NOR2_X1 U10367 ( .A1(n4513), .A2(n9733), .ZN(n9056) );
  OAI22_X1 U10368 ( .A1(n9054), .A2(n9222), .B1(n9053), .B2(n9762), .ZN(n9055)
         );
  AOI211_X1 U10369 ( .C1(n9306), .C2(n9152), .A(n9056), .B(n9055), .ZN(n9068)
         );
  INV_X1 U10370 ( .A(n9057), .ZN(n9061) );
  OAI21_X1 U10371 ( .B1(n4286), .B2(n9059), .A(n9058), .ZN(n9060) );
  NAND2_X1 U10372 ( .A1(n9090), .A2(n9739), .ZN(n9064) );
  NAND2_X1 U10373 ( .A1(n9062), .A2(n9756), .ZN(n9063) );
  OR2_X1 U10374 ( .A1(n9309), .A2(n9234), .ZN(n9067) );
  OAI211_X1 U10375 ( .C1(n9305), .C2(n9297), .A(n9068), .B(n9067), .ZN(
        P1_U3263) );
  XNOR2_X1 U10376 ( .A(n9069), .B(n9005), .ZN(n9315) );
  INV_X1 U10377 ( .A(n9084), .ZN(n9072) );
  INV_X1 U10378 ( .A(n9070), .ZN(n9071) );
  AOI21_X1 U10379 ( .B1(n9311), .B2(n9072), .A(n9071), .ZN(n9312) );
  AOI22_X1 U10380 ( .A1(n9073), .A2(n9747), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9234), .ZN(n9074) );
  OAI21_X1 U10381 ( .B1(n9075), .B2(n9733), .A(n9074), .ZN(n9081) );
  XNOR2_X1 U10382 ( .A(n9077), .B(n9076), .ZN(n9079) );
  AOI211_X1 U10383 ( .C1(n9312), .C2(n9718), .A(n9081), .B(n9080), .ZN(n9082)
         );
  OAI21_X1 U10384 ( .B1(n9315), .B2(n9297), .A(n9082), .ZN(P1_U3264) );
  XNOR2_X1 U10385 ( .A(n9083), .B(n9089), .ZN(n9320) );
  AOI21_X1 U10386 ( .B1(n9316), .B2(n9096), .A(n9084), .ZN(n9317) );
  AOI22_X1 U10387 ( .A1(n9085), .A2(n9747), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9234), .ZN(n9086) );
  OAI21_X1 U10388 ( .B1(n9087), .B2(n9733), .A(n9086), .ZN(n9093) );
  XOR2_X1 U10389 ( .A(n9089), .B(n9088), .Z(n9091) );
  AOI211_X1 U10390 ( .C1(n9317), .C2(n9718), .A(n9093), .B(n9092), .ZN(n9094)
         );
  OAI21_X1 U10391 ( .B1(n9297), .B2(n9320), .A(n9094), .ZN(P1_U3265) );
  XOR2_X1 U10392 ( .A(n9104), .B(n9095), .Z(n9325) );
  INV_X1 U10393 ( .A(n9111), .ZN(n9098) );
  INV_X1 U10394 ( .A(n9096), .ZN(n9097) );
  AOI21_X1 U10395 ( .B1(n9321), .B2(n9098), .A(n9097), .ZN(n9322) );
  INV_X1 U10396 ( .A(n9099), .ZN(n9100) );
  AOI22_X1 U10397 ( .A1(n9100), .A2(n9747), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9234), .ZN(n9101) );
  OAI21_X1 U10398 ( .B1(n9102), .B2(n9733), .A(n9101), .ZN(n9108) );
  XOR2_X1 U10399 ( .A(n9104), .B(n9103), .Z(n9106) );
  AOI222_X1 U10400 ( .A1(n9727), .A2(n9106), .B1(n9127), .B2(n9739), .C1(n9105), .C2(n9756), .ZN(n9324) );
  NOR2_X1 U10401 ( .A1(n9324), .A2(n9234), .ZN(n9107) );
  AOI211_X1 U10402 ( .C1(n9322), .C2(n9718), .A(n9108), .B(n9107), .ZN(n9109)
         );
  OAI21_X1 U10403 ( .B1(n9325), .B2(n9297), .A(n9109), .ZN(P1_U3266) );
  XNOR2_X1 U10404 ( .A(n9110), .B(n9118), .ZN(n9330) );
  AOI211_X1 U10405 ( .C1(n9327), .C2(n9136), .A(n9819), .B(n9111), .ZN(n9326)
         );
  AOI22_X1 U10406 ( .A1(n9112), .A2(n9747), .B1(n9291), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n9113) );
  OAI21_X1 U10407 ( .B1(n9114), .B2(n9733), .A(n9113), .ZN(n9124) );
  AND2_X1 U10408 ( .A1(n9116), .A2(n9115), .ZN(n9119) );
  OAI21_X1 U10409 ( .B1(n9119), .B2(n9118), .A(n9117), .ZN(n9122) );
  AOI222_X1 U10410 ( .A1(n9727), .A2(n9122), .B1(n9121), .B2(n9739), .C1(n9120), .C2(n9756), .ZN(n9329) );
  NOR2_X1 U10411 ( .A1(n9329), .A2(n9234), .ZN(n9123) );
  AOI211_X1 U10412 ( .C1(n9152), .C2(n9326), .A(n9124), .B(n9123), .ZN(n9125)
         );
  OAI21_X1 U10413 ( .B1(n9330), .B2(n9297), .A(n9125), .ZN(P1_U3267) );
  XNOR2_X1 U10414 ( .A(n9126), .B(n9130), .ZN(n9128) );
  AOI222_X1 U10415 ( .A1(n9727), .A2(n9128), .B1(n9127), .B2(n9756), .C1(n9167), .C2(n9739), .ZN(n9475) );
  OAI21_X1 U10416 ( .B1(n9131), .B2(n9130), .A(n9129), .ZN(n9132) );
  INV_X1 U10417 ( .A(n9132), .ZN(n9476) );
  OAI22_X1 U10418 ( .A1(n9762), .A2(n9134), .B1(n9133), .B2(n9222), .ZN(n9135)
         );
  AOI21_X1 U10419 ( .B1(n9473), .B2(n9226), .A(n9135), .ZN(n9139) );
  AOI21_X1 U10420 ( .B1(n9473), .B2(n9144), .A(n9819), .ZN(n9137) );
  AND2_X1 U10421 ( .A1(n9137), .A2(n9136), .ZN(n9472) );
  NAND2_X1 U10422 ( .A1(n9472), .A2(n9152), .ZN(n9138) );
  OAI211_X1 U10423 ( .C1(n9476), .C2(n9297), .A(n9139), .B(n9138), .ZN(n9140)
         );
  INV_X1 U10424 ( .A(n9140), .ZN(n9141) );
  OAI21_X1 U10425 ( .B1(n9234), .B2(n9475), .A(n9141), .ZN(P1_U3268) );
  XNOR2_X1 U10426 ( .A(n9143), .B(n9142), .ZN(n9481) );
  INV_X1 U10427 ( .A(n9170), .ZN(n9146) );
  INV_X1 U10428 ( .A(n9144), .ZN(n9145) );
  AOI211_X1 U10429 ( .C1(n9479), .C2(n9146), .A(n9819), .B(n9145), .ZN(n9478)
         );
  NOR2_X1 U10430 ( .A1(n9147), .A2(n9733), .ZN(n9151) );
  OAI22_X1 U10431 ( .A1(n9762), .A2(n9149), .B1(n9148), .B2(n9222), .ZN(n9150)
         );
  AOI211_X1 U10432 ( .C1(n9478), .C2(n9152), .A(n9151), .B(n9150), .ZN(n9159)
         );
  XNOR2_X1 U10433 ( .A(n9154), .B(n9153), .ZN(n9155) );
  OAI222_X1 U10434 ( .A1(n9723), .A2(n9157), .B1(n9724), .B2(n9156), .C1(n9155), .C2(n9751), .ZN(n9477) );
  NAND2_X1 U10435 ( .A1(n9477), .A2(n9762), .ZN(n9158) );
  OAI211_X1 U10436 ( .C1(n9481), .C2(n9297), .A(n9159), .B(n9158), .ZN(
        P1_U3269) );
  XNOR2_X1 U10437 ( .A(n9160), .B(n9163), .ZN(n9486) );
  INV_X1 U10438 ( .A(n9161), .ZN(n9162) );
  NAND2_X1 U10439 ( .A1(n9163), .A2(n9162), .ZN(n9165) );
  OAI21_X1 U10440 ( .B1(n9166), .B2(n9165), .A(n9164), .ZN(n9169) );
  AOI222_X1 U10441 ( .A1(n9727), .A2(n9169), .B1(n9168), .B2(n9739), .C1(n9167), .C2(n9756), .ZN(n9485) );
  AOI211_X1 U10442 ( .C1(n9483), .C2(n4518), .A(n9819), .B(n9170), .ZN(n9482)
         );
  AOI22_X1 U10443 ( .A1(n9482), .A2(n5638), .B1(n9747), .B2(n9171), .ZN(n9172)
         );
  AOI21_X1 U10444 ( .B1(n9485), .B2(n9172), .A(n9291), .ZN(n9176) );
  OAI22_X1 U10445 ( .A1(n9174), .A2(n9733), .B1(n9173), .B2(n9762), .ZN(n9175)
         );
  NOR2_X1 U10446 ( .A1(n9176), .A2(n9175), .ZN(n9177) );
  OAI21_X1 U10447 ( .B1(n9297), .B2(n9486), .A(n9177), .ZN(P1_U3270) );
  XOR2_X1 U10448 ( .A(n9184), .B(n9178), .Z(n9491) );
  AOI21_X1 U10449 ( .B1(n9487), .B2(n9197), .A(n9179), .ZN(n9488) );
  INV_X1 U10450 ( .A(n9180), .ZN(n9181) );
  AOI22_X1 U10451 ( .A1(n9291), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9181), .B2(
        n9747), .ZN(n9182) );
  OAI21_X1 U10452 ( .B1(n9183), .B2(n9733), .A(n9182), .ZN(n9189) );
  XNOR2_X1 U10453 ( .A(n9185), .B(n9184), .ZN(n9187) );
  AOI222_X1 U10454 ( .A1(n9727), .A2(n9187), .B1(n9186), .B2(n9756), .C1(n9215), .C2(n9739), .ZN(n9490) );
  NOR2_X1 U10455 ( .A1(n9490), .A2(n9234), .ZN(n9188) );
  AOI211_X1 U10456 ( .C1(n9488), .C2(n9718), .A(n9189), .B(n9188), .ZN(n9190)
         );
  OAI21_X1 U10457 ( .B1(n9491), .B2(n9297), .A(n9190), .ZN(P1_U3271) );
  INV_X1 U10458 ( .A(n9191), .ZN(n9195) );
  AOI21_X1 U10459 ( .B1(n9195), .B2(n9194), .A(n9193), .ZN(n9196) );
  INV_X1 U10460 ( .A(n9196), .ZN(n9497) );
  INV_X1 U10461 ( .A(n9197), .ZN(n9198) );
  AOI21_X1 U10462 ( .B1(n9493), .B2(n9228), .A(n9198), .ZN(n9494) );
  INV_X1 U10463 ( .A(n9493), .ZN(n9199) );
  NOR2_X1 U10464 ( .A1(n9199), .A2(n9733), .ZN(n9203) );
  OAI22_X1 U10465 ( .A1(n9762), .A2(n9201), .B1(n9200), .B2(n9222), .ZN(n9202)
         );
  AOI211_X1 U10466 ( .C1(n9494), .C2(n9718), .A(n9203), .B(n9202), .ZN(n9210)
         );
  AOI21_X1 U10467 ( .B1(n9205), .B2(n8991), .A(n9204), .ZN(n9206) );
  OAI222_X1 U10468 ( .A1(n9723), .A2(n9208), .B1(n9724), .B2(n9207), .C1(n9751), .C2(n9206), .ZN(n9492) );
  NAND2_X1 U10469 ( .A1(n9492), .A2(n9762), .ZN(n9209) );
  OAI211_X1 U10470 ( .C1(n9497), .C2(n9297), .A(n9210), .B(n9209), .ZN(
        P1_U3272) );
  NAND2_X1 U10471 ( .A1(n9212), .A2(n9211), .ZN(n9213) );
  XOR2_X1 U10472 ( .A(n9218), .B(n9213), .Z(n9216) );
  AOI222_X1 U10473 ( .A1(n9727), .A2(n9216), .B1(n9215), .B2(n9756), .C1(n9214), .C2(n9739), .ZN(n9502) );
  INV_X1 U10474 ( .A(n9217), .ZN(n9221) );
  NAND2_X1 U10475 ( .A1(n9219), .A2(n9218), .ZN(n9498) );
  NAND3_X1 U10476 ( .A1(n9221), .A2(n9220), .A3(n9498), .ZN(n9232) );
  OAI22_X1 U10477 ( .A1(n9762), .A2(n9224), .B1(n9223), .B2(n9222), .ZN(n9225)
         );
  AOI21_X1 U10478 ( .B1(n9499), .B2(n9226), .A(n9225), .ZN(n9231) );
  OR2_X1 U10479 ( .A1(n9236), .A2(n9227), .ZN(n9229) );
  AND2_X1 U10480 ( .A1(n9229), .A2(n9228), .ZN(n9500) );
  NAND2_X1 U10481 ( .A1(n9500), .A2(n9718), .ZN(n9230) );
  AND3_X1 U10482 ( .A1(n9232), .A2(n9231), .A3(n9230), .ZN(n9233) );
  OAI21_X1 U10483 ( .B1(n9502), .B2(n9234), .A(n9233), .ZN(P1_U3273) );
  XNOR2_X1 U10484 ( .A(n9235), .B(n9241), .ZN(n9508) );
  AOI21_X1 U10485 ( .B1(n9504), .B2(n9253), .A(n9236), .ZN(n9505) );
  AOI22_X1 U10486 ( .A1(n9291), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9237), .B2(
        n9747), .ZN(n9238) );
  OAI21_X1 U10487 ( .B1(n9239), .B2(n9733), .A(n9238), .ZN(n9245) );
  XOR2_X1 U10488 ( .A(n9241), .B(n9240), .Z(n9243) );
  AOI222_X1 U10489 ( .A1(n9727), .A2(n9243), .B1(n9242), .B2(n9756), .C1(n9265), .C2(n9739), .ZN(n9507) );
  NOR2_X1 U10490 ( .A1(n9507), .A2(n9234), .ZN(n9244) );
  AOI211_X1 U10491 ( .C1(n9505), .C2(n9718), .A(n9245), .B(n9244), .ZN(n9246)
         );
  OAI21_X1 U10492 ( .B1(n9297), .B2(n9508), .A(n9246), .ZN(P1_U3274) );
  XNOR2_X1 U10493 ( .A(n9247), .B(n9249), .ZN(n9513) );
  AOI21_X1 U10494 ( .B1(n9250), .B2(n9249), .A(n9248), .ZN(n9251) );
  OAI222_X1 U10495 ( .A1(n9723), .A2(n9252), .B1(n9724), .B2(n9285), .C1(n9751), .C2(n9251), .ZN(n9509) );
  INV_X1 U10496 ( .A(n9511), .ZN(n9258) );
  INV_X1 U10497 ( .A(n9253), .ZN(n9254) );
  AOI211_X1 U10498 ( .C1(n9511), .C2(n9271), .A(n9819), .B(n9254), .ZN(n9510)
         );
  NAND2_X1 U10499 ( .A1(n9510), .A2(n9289), .ZN(n9257) );
  AOI22_X1 U10500 ( .A1(n9291), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9255), .B2(
        n9747), .ZN(n9256) );
  OAI211_X1 U10501 ( .C1(n9258), .C2(n9733), .A(n9257), .B(n9256), .ZN(n9259)
         );
  AOI21_X1 U10502 ( .B1(n9509), .B2(n9762), .A(n9259), .ZN(n9260) );
  OAI21_X1 U10503 ( .B1(n9297), .B2(n9513), .A(n9260), .ZN(P1_U3275) );
  XNOR2_X1 U10504 ( .A(n9261), .B(n9264), .ZN(n9275) );
  AOI21_X1 U10505 ( .B1(n9264), .B2(n9263), .A(n9262), .ZN(n9268) );
  AOI22_X1 U10506 ( .A1(n9739), .A2(n9266), .B1(n9756), .B2(n9265), .ZN(n9267)
         );
  OAI21_X1 U10507 ( .B1(n9268), .B2(n9751), .A(n9267), .ZN(n9269) );
  AOI21_X1 U10508 ( .B1(n9270), .B2(n9275), .A(n9269), .ZN(n9517) );
  AOI21_X1 U10509 ( .B1(n9514), .B2(n9287), .A(n4524), .ZN(n9515) );
  AOI22_X1 U10510 ( .A1(n9291), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9272), .B2(
        n9747), .ZN(n9273) );
  OAI21_X1 U10511 ( .B1(n9274), .B2(n9733), .A(n9273), .ZN(n9278) );
  INV_X1 U10512 ( .A(n9275), .ZN(n9518) );
  NOR2_X1 U10513 ( .A1(n9518), .A2(n9276), .ZN(n9277) );
  AOI211_X1 U10514 ( .C1(n9515), .C2(n9718), .A(n9278), .B(n9277), .ZN(n9279)
         );
  OAI21_X1 U10515 ( .B1(n9291), .B2(n9517), .A(n9279), .ZN(P1_U3276) );
  XNOR2_X1 U10516 ( .A(n9280), .B(n9281), .ZN(n9523) );
  XNOR2_X1 U10517 ( .A(n9282), .B(n9281), .ZN(n9283) );
  OAI222_X1 U10518 ( .A1(n9723), .A2(n9285), .B1(n9724), .B2(n9284), .C1(n9751), .C2(n9283), .ZN(n9519) );
  INV_X1 U10519 ( .A(n9286), .ZN(n9288) );
  AOI211_X1 U10520 ( .C1(n9521), .C2(n9288), .A(n9819), .B(n4521), .ZN(n9520)
         );
  NAND2_X1 U10521 ( .A1(n9520), .A2(n9289), .ZN(n9293) );
  AOI22_X1 U10522 ( .A1(n9291), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9290), .B2(
        n9747), .ZN(n9292) );
  OAI211_X1 U10523 ( .C1(n9294), .C2(n9733), .A(n9293), .B(n9292), .ZN(n9295)
         );
  AOI21_X1 U10524 ( .B1(n9519), .B2(n9762), .A(n9295), .ZN(n9296) );
  OAI21_X1 U10525 ( .B1(n9523), .B2(n9297), .A(n9296), .ZN(P1_U3277) );
  NAND2_X1 U10526 ( .A1(n9298), .A2(n9815), .ZN(n9304) );
  OAI22_X1 U10527 ( .A1(n9300), .A2(n9819), .B1(n9299), .B2(n9817), .ZN(n9301)
         );
  NOR2_X1 U10528 ( .A1(n9302), .A2(n9301), .ZN(n9303) );
  NAND2_X1 U10529 ( .A1(n9304), .A2(n9303), .ZN(n9525) );
  MUX2_X1 U10530 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9525), .S(n9843), .Z(
        P1_U3552) );
  AOI21_X1 U10531 ( .B1(n9598), .B2(n9307), .A(n9306), .ZN(n9308) );
  NAND3_X1 U10532 ( .A1(n9310), .A2(n9309), .A3(n9308), .ZN(n9526) );
  MUX2_X1 U10533 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9526), .S(n9843), .Z(
        P1_U3551) );
  AOI22_X1 U10534 ( .A1(n9312), .A2(n9742), .B1(n9598), .B2(n9311), .ZN(n9313)
         );
  OAI211_X1 U10535 ( .C1(n9315), .C2(n9524), .A(n9314), .B(n9313), .ZN(n9527)
         );
  MUX2_X1 U10536 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9527), .S(n9843), .Z(
        P1_U3550) );
  AOI22_X1 U10537 ( .A1(n9317), .A2(n9742), .B1(n9598), .B2(n9316), .ZN(n9318)
         );
  OAI211_X1 U10538 ( .C1(n9320), .C2(n9524), .A(n9319), .B(n9318), .ZN(n9528)
         );
  MUX2_X1 U10539 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9528), .S(n9843), .Z(
        P1_U3549) );
  AOI22_X1 U10540 ( .A1(n9322), .A2(n9742), .B1(n9598), .B2(n9321), .ZN(n9323)
         );
  OAI211_X1 U10541 ( .C1(n9325), .C2(n9524), .A(n9324), .B(n9323), .ZN(n9529)
         );
  MUX2_X1 U10542 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9529), .S(n9843), .Z(
        P1_U3548) );
  AOI21_X1 U10543 ( .B1(n9598), .B2(n9327), .A(n9326), .ZN(n9328) );
  OAI211_X1 U10544 ( .C1(n9330), .C2(n9524), .A(n9329), .B(n9328), .ZN(n9530)
         );
  MUX2_X1 U10545 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9530), .S(n9843), .Z(n9471) );
  INV_X1 U10546 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n9332) );
  AOI22_X1 U10547 ( .A1(n9332), .A2(keyinput17), .B1(n6274), .B2(keyinput59), 
        .ZN(n9331) );
  OAI221_X1 U10548 ( .B1(n9332), .B2(keyinput17), .C1(n6274), .C2(keyinput59), 
        .A(n9331), .ZN(n9336) );
  INV_X1 U10549 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n9905) );
  INV_X1 U10550 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9767) );
  AOI22_X1 U10551 ( .A1(n9905), .A2(keyinput16), .B1(n9767), .B2(keyinput49), 
        .ZN(n9333) );
  OAI221_X1 U10552 ( .B1(n9905), .B2(keyinput16), .C1(n9767), .C2(keyinput49), 
        .A(n9333), .ZN(n9335) );
  INV_X1 U10553 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9769) );
  XNOR2_X1 U10554 ( .A(n9769), .B(keyinput25), .ZN(n9334) );
  NOR3_X1 U10555 ( .A1(n9336), .A2(n9335), .A3(n9334), .ZN(n9354) );
  INV_X1 U10556 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9426) );
  AOI22_X1 U10557 ( .A1(n9425), .A2(keyinput27), .B1(n9426), .B2(keyinput38), 
        .ZN(n9337) );
  OAI221_X1 U10558 ( .B1(n9425), .B2(keyinput27), .C1(n9426), .C2(keyinput38), 
        .A(n9337), .ZN(n9343) );
  INV_X1 U10559 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9456) );
  AOI22_X1 U10560 ( .A1(n9457), .A2(keyinput8), .B1(keyinput11), .B2(n9456), 
        .ZN(n9338) );
  OAI221_X1 U10561 ( .B1(n9457), .B2(keyinput8), .C1(n9456), .C2(keyinput11), 
        .A(n9338), .ZN(n9342) );
  AOI22_X1 U10562 ( .A1(n10051), .A2(keyinput28), .B1(n9340), .B2(keyinput48), 
        .ZN(n9339) );
  OAI221_X1 U10563 ( .B1(n10051), .B2(keyinput28), .C1(n9340), .C2(keyinput48), 
        .A(n9339), .ZN(n9341) );
  NOR3_X1 U10564 ( .A1(n9343), .A2(n9342), .A3(n9341), .ZN(n9353) );
  INV_X1 U10565 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9615) );
  AOI22_X1 U10566 ( .A1(n9615), .A2(keyinput13), .B1(keyinput51), .B2(n9578), 
        .ZN(n9344) );
  OAI221_X1 U10567 ( .B1(n9615), .B2(keyinput13), .C1(n9578), .C2(keyinput51), 
        .A(n9344), .ZN(n9351) );
  AOI22_X1 U10568 ( .A1(n9450), .A2(keyinput57), .B1(n9346), .B2(keyinput22), 
        .ZN(n9345) );
  OAI221_X1 U10569 ( .B1(n9450), .B2(keyinput57), .C1(n9346), .C2(keyinput22), 
        .A(n9345), .ZN(n9350) );
  AOI22_X1 U10570 ( .A1(n9458), .A2(keyinput3), .B1(keyinput4), .B2(n9348), 
        .ZN(n9347) );
  OAI221_X1 U10571 ( .B1(n9458), .B2(keyinput3), .C1(n9348), .C2(keyinput4), 
        .A(n9347), .ZN(n9349) );
  NOR3_X1 U10572 ( .A1(n9351), .A2(n9350), .A3(n9349), .ZN(n9352) );
  AND3_X1 U10573 ( .A1(n9354), .A2(n9353), .A3(n9352), .ZN(n9389) );
  AOI22_X1 U10574 ( .A1(n9436), .A2(keyinput45), .B1(keyinput33), .B2(n9356), 
        .ZN(n9355) );
  OAI221_X1 U10575 ( .B1(n9436), .B2(keyinput45), .C1(n9356), .C2(keyinput33), 
        .A(n9355), .ZN(n9364) );
  AOI22_X1 U10576 ( .A1(n5002), .A2(keyinput10), .B1(n9429), .B2(keyinput6), 
        .ZN(n9357) );
  OAI221_X1 U10577 ( .B1(n5002), .B2(keyinput10), .C1(n9429), .C2(keyinput6), 
        .A(n9357), .ZN(n9363) );
  AOI22_X1 U10578 ( .A1(n4884), .A2(keyinput46), .B1(n9449), .B2(keyinput58), 
        .ZN(n9358) );
  OAI221_X1 U10579 ( .B1(n4884), .B2(keyinput46), .C1(n9449), .C2(keyinput58), 
        .A(n9358), .ZN(n9362) );
  INV_X1 U10580 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n9907) );
  AOI22_X1 U10581 ( .A1(n9907), .A2(keyinput54), .B1(n9360), .B2(keyinput18), 
        .ZN(n9359) );
  OAI221_X1 U10582 ( .B1(n9907), .B2(keyinput54), .C1(n9360), .C2(keyinput18), 
        .A(n9359), .ZN(n9361) );
  NOR4_X1 U10583 ( .A1(n9364), .A2(n9363), .A3(n9362), .A4(n9361), .ZN(n9388)
         );
  INV_X1 U10584 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n9893) );
  AOI22_X1 U10585 ( .A1(n9893), .A2(keyinput0), .B1(keyinput21), .B2(n4922), 
        .ZN(n9365) );
  OAI221_X1 U10586 ( .B1(n9893), .B2(keyinput0), .C1(n4922), .C2(keyinput21), 
        .A(n9365), .ZN(n9368) );
  AOI22_X1 U10587 ( .A1(n9428), .A2(keyinput5), .B1(keyinput39), .B2(n9437), 
        .ZN(n9366) );
  OAI221_X1 U10588 ( .B1(n9428), .B2(keyinput5), .C1(n9437), .C2(keyinput39), 
        .A(n9366), .ZN(n9367) );
  NOR2_X1 U10589 ( .A1(n9368), .A2(n9367), .ZN(n9387) );
  INV_X1 U10590 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9914) );
  INV_X1 U10591 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9370) );
  AOI22_X1 U10592 ( .A1(n9914), .A2(keyinput42), .B1(n9370), .B2(keyinput12), 
        .ZN(n9369) );
  OAI221_X1 U10593 ( .B1(n9914), .B2(keyinput42), .C1(n9370), .C2(keyinput12), 
        .A(n9369), .ZN(n9385) );
  INV_X1 U10594 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n9372) );
  AOI22_X1 U10595 ( .A1(n9372), .A2(keyinput24), .B1(n9435), .B2(keyinput55), 
        .ZN(n9371) );
  OAI221_X1 U10596 ( .B1(n9372), .B2(keyinput24), .C1(n9435), .C2(keyinput55), 
        .A(n9371), .ZN(n9384) );
  XNOR2_X1 U10597 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput52), .ZN(n9375) );
  XNOR2_X1 U10598 ( .A(SI_2_), .B(keyinput9), .ZN(n9374) );
  XNOR2_X1 U10599 ( .A(keyinput32), .B(P2_REG3_REG_1__SCAN_IN), .ZN(n9373) );
  AND3_X1 U10600 ( .A1(n9375), .A2(n9374), .A3(n9373), .ZN(n9382) );
  XNOR2_X1 U10601 ( .A(keyinput1), .B(n4934), .ZN(n9378) );
  INV_X1 U10602 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n9376) );
  XNOR2_X1 U10603 ( .A(keyinput50), .B(n9376), .ZN(n9377) );
  NOR2_X1 U10604 ( .A1(n9378), .A2(n9377), .ZN(n9381) );
  XNOR2_X1 U10605 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput36), .ZN(n9380) );
  XNOR2_X1 U10606 ( .A(P2_REG2_REG_1__SCAN_IN), .B(keyinput63), .ZN(n9379) );
  NAND4_X1 U10607 ( .A1(n9382), .A2(n9381), .A3(n9380), .A4(n9379), .ZN(n9383)
         );
  NOR3_X1 U10608 ( .A1(n9385), .A2(n9384), .A3(n9383), .ZN(n9386) );
  AND4_X1 U10609 ( .A1(n9389), .A2(n9388), .A3(n9387), .A4(n9386), .ZN(n9423)
         );
  AOI22_X1 U10610 ( .A1(n9424), .A2(keyinput56), .B1(n9455), .B2(keyinput15), 
        .ZN(n9390) );
  OAI221_X1 U10611 ( .B1(n9424), .B2(keyinput56), .C1(n9455), .C2(keyinput15), 
        .A(n9390), .ZN(n9400) );
  INV_X1 U10612 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n9911) );
  AOI22_X1 U10613 ( .A1(n9911), .A2(keyinput19), .B1(keyinput60), .B2(n9392), 
        .ZN(n9391) );
  OAI221_X1 U10614 ( .B1(n9911), .B2(keyinput19), .C1(n9392), .C2(keyinput60), 
        .A(n9391), .ZN(n9399) );
  AOI22_X1 U10615 ( .A1(n9395), .A2(keyinput29), .B1(n9394), .B2(keyinput37), 
        .ZN(n9393) );
  OAI221_X1 U10616 ( .B1(n9395), .B2(keyinput29), .C1(n9394), .C2(keyinput37), 
        .A(n9393), .ZN(n9398) );
  INV_X1 U10617 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n9901) );
  AOI22_X1 U10618 ( .A1(n9901), .A2(keyinput44), .B1(n6186), .B2(keyinput2), 
        .ZN(n9396) );
  OAI221_X1 U10619 ( .B1(n9901), .B2(keyinput44), .C1(n6186), .C2(keyinput2), 
        .A(n9396), .ZN(n9397) );
  NOR4_X1 U10620 ( .A1(n9400), .A2(n9399), .A3(n9398), .A4(n9397), .ZN(n9422)
         );
  INV_X1 U10621 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n9886) );
  INV_X1 U10622 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9766) );
  AOI22_X1 U10623 ( .A1(n9886), .A2(keyinput43), .B1(n9766), .B2(keyinput23), 
        .ZN(n9401) );
  OAI221_X1 U10624 ( .B1(n9886), .B2(keyinput43), .C1(n9766), .C2(keyinput23), 
        .A(n9401), .ZN(n9408) );
  AOI22_X1 U10625 ( .A1(n6148), .A2(keyinput7), .B1(keyinput47), .B2(n4920), 
        .ZN(n9402) );
  OAI221_X1 U10626 ( .B1(n6148), .B2(keyinput7), .C1(n4920), .C2(keyinput47), 
        .A(n9402), .ZN(n9407) );
  AOI22_X1 U10627 ( .A1(n9624), .A2(keyinput62), .B1(keyinput14), .B2(n9451), 
        .ZN(n9403) );
  OAI221_X1 U10628 ( .B1(n9624), .B2(keyinput62), .C1(n9451), .C2(keyinput14), 
        .A(n9403), .ZN(n9406) );
  INV_X1 U10629 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9768) );
  AOI22_X1 U10630 ( .A1(n9454), .A2(keyinput41), .B1(n9768), .B2(keyinput34), 
        .ZN(n9404) );
  OAI221_X1 U10631 ( .B1(n9454), .B2(keyinput41), .C1(n9768), .C2(keyinput34), 
        .A(n9404), .ZN(n9405) );
  NOR4_X1 U10632 ( .A1(n9408), .A2(n9407), .A3(n9406), .A4(n9405), .ZN(n9421)
         );
  AOI22_X1 U10633 ( .A1(n9410), .A2(keyinput53), .B1(n9427), .B2(keyinput31), 
        .ZN(n9409) );
  OAI221_X1 U10634 ( .B1(n9410), .B2(keyinput53), .C1(n9427), .C2(keyinput31), 
        .A(n9409), .ZN(n9419) );
  INV_X1 U10635 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9446) );
  AOI22_X1 U10636 ( .A1(n4843), .A2(keyinput35), .B1(keyinput20), .B2(n9446), 
        .ZN(n9411) );
  OAI221_X1 U10637 ( .B1(n4843), .B2(keyinput35), .C1(n9446), .C2(keyinput20), 
        .A(n9411), .ZN(n9418) );
  INV_X1 U10638 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9413) );
  AOI22_X1 U10639 ( .A1(n9413), .A2(keyinput61), .B1(keyinput30), .B2(n9434), 
        .ZN(n9412) );
  OAI221_X1 U10640 ( .B1(n9413), .B2(keyinput61), .C1(n9434), .C2(keyinput30), 
        .A(n9412), .ZN(n9417) );
  AOI22_X1 U10641 ( .A1(n5374), .A2(keyinput26), .B1(keyinput40), .B2(n9415), 
        .ZN(n9414) );
  OAI221_X1 U10642 ( .B1(n5374), .B2(keyinput26), .C1(n9415), .C2(keyinput40), 
        .A(n9414), .ZN(n9416) );
  NOR4_X1 U10643 ( .A1(n9419), .A2(n9418), .A3(n9417), .A4(n9416), .ZN(n9420)
         );
  NAND4_X1 U10644 ( .A1(n9423), .A2(n9422), .A3(n9421), .A4(n9420), .ZN(n9469)
         );
  NOR4_X1 U10645 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .A3(n9911), .A4(n9424), .ZN(n9466) );
  AND4_X1 U10646 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_REG2_REG_30__SCAN_IN), 
        .A3(n9426), .A4(n9425), .ZN(n9433) );
  AND4_X1 U10647 ( .A1(SI_8_), .A2(P2_DATAO_REG_8__SCAN_IN), .A3(n9428), .A4(
        n9427), .ZN(n9432) );
  AND3_X1 U10648 ( .A1(P1_REG2_REG_26__SCAN_IN), .A2(P2_REG0_REG_4__SCAN_IN), 
        .A3(P2_REG0_REG_2__SCAN_IN), .ZN(n9431) );
  NOR3_X1 U10649 ( .A1(SI_24_), .A2(P2_DATAO_REG_20__SCAN_IN), .A3(n9429), 
        .ZN(n9430) );
  NAND4_X1 U10650 ( .A1(n9433), .A2(n9432), .A3(n9431), .A4(n9430), .ZN(n9443)
         );
  NOR4_X1 U10651 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .A3(P2_REG3_REG_2__SCAN_IN), .A4(n9434), .ZN(n9441) );
  NOR4_X1 U10652 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(P1_REG2_REG_6__SCAN_IN), 
        .A3(P1_REG1_REG_0__SCAN_IN), .A4(P2_REG3_REG_1__SCAN_IN), .ZN(n9440)
         );
  NOR4_X1 U10653 ( .A1(P1_REG0_REG_15__SCAN_IN), .A2(P1_REG1_REG_14__SCAN_IN), 
        .A3(P1_REG0_REG_11__SCAN_IN), .A4(n9435), .ZN(n9439) );
  NOR4_X1 U10654 ( .A1(P2_REG0_REG_7__SCAN_IN), .A2(P1_DATAO_REG_30__SCAN_IN), 
        .A3(n9437), .A4(n9436), .ZN(n9438) );
  NAND4_X1 U10655 ( .A1(n9441), .A2(n9440), .A3(n9439), .A4(n9438), .ZN(n9442)
         );
  NOR2_X1 U10656 ( .A1(n9443), .A2(n9442), .ZN(n9444) );
  AND2_X1 U10657 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(n9444), .ZN(n9445) );
  NAND4_X1 U10658 ( .A1(n9445), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P1_ADDR_REG_6__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n9448) );
  NAND4_X1 U10659 ( .A1(n9446), .A2(n9768), .A3(n10051), .A4(
        P2_ADDR_REG_12__SCAN_IN), .ZN(n9447) );
  NOR2_X1 U10660 ( .A1(n9448), .A2(n9447), .ZN(n9463) );
  NAND4_X1 U10661 ( .A1(n9450), .A2(n9449), .A3(n4854), .A4(SI_2_), .ZN(n9453)
         );
  NAND4_X1 U10662 ( .A1(n9372), .A2(n9451), .A3(P2_REG1_REG_14__SCAN_IN), .A4(
        P2_REG2_REG_1__SCAN_IN), .ZN(n9452) );
  NOR2_X1 U10663 ( .A1(n9453), .A2(n9452), .ZN(n9462) );
  NAND4_X1 U10664 ( .A1(n9456), .A2(n9455), .A3(n9454), .A4(
        P1_D_REG_0__SCAN_IN), .ZN(n9460) );
  NAND4_X1 U10665 ( .A1(n9458), .A2(n9457), .A3(P1_IR_REG_24__SCAN_IN), .A4(
        P1_REG3_REG_6__SCAN_IN), .ZN(n9459) );
  NOR2_X1 U10666 ( .A1(n9460), .A2(n9459), .ZN(n9461) );
  AND4_X1 U10667 ( .A1(n9464), .A2(n9463), .A3(n9462), .A4(n9461), .ZN(n9465)
         );
  NAND3_X1 U10668 ( .A1(n9467), .A2(n9466), .A3(n9465), .ZN(n9468) );
  XNOR2_X1 U10669 ( .A(n9469), .B(n9468), .ZN(n9470) );
  XNOR2_X1 U10670 ( .A(n9471), .B(n9470), .ZN(P1_U3547) );
  AOI21_X1 U10671 ( .B1(n9598), .B2(n9473), .A(n9472), .ZN(n9474) );
  OAI211_X1 U10672 ( .C1(n9476), .C2(n9524), .A(n9475), .B(n9474), .ZN(n9531)
         );
  MUX2_X1 U10673 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9531), .S(n9843), .Z(
        P1_U3546) );
  AOI211_X1 U10674 ( .C1(n9598), .C2(n9479), .A(n9478), .B(n9477), .ZN(n9480)
         );
  OAI21_X1 U10675 ( .B1(n9481), .B2(n9524), .A(n9480), .ZN(n9532) );
  MUX2_X1 U10676 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9532), .S(n9843), .Z(
        P1_U3545) );
  AOI21_X1 U10677 ( .B1(n9598), .B2(n9483), .A(n9482), .ZN(n9484) );
  OAI211_X1 U10678 ( .C1(n9486), .C2(n9524), .A(n9485), .B(n9484), .ZN(n9533)
         );
  MUX2_X1 U10679 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9533), .S(n9843), .Z(
        P1_U3544) );
  AOI22_X1 U10680 ( .A1(n9488), .A2(n9742), .B1(n9598), .B2(n9487), .ZN(n9489)
         );
  OAI211_X1 U10681 ( .C1(n9491), .C2(n9524), .A(n9490), .B(n9489), .ZN(n9534)
         );
  MUX2_X1 U10682 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9534), .S(n9843), .Z(
        P1_U3543) );
  INV_X1 U10683 ( .A(n9492), .ZN(n9496) );
  AOI22_X1 U10684 ( .A1(n9494), .A2(n9742), .B1(n9598), .B2(n9493), .ZN(n9495)
         );
  OAI211_X1 U10685 ( .C1(n9497), .C2(n9524), .A(n9496), .B(n9495), .ZN(n9535)
         );
  MUX2_X1 U10686 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9535), .S(n9843), .Z(
        P1_U3542) );
  NAND2_X1 U10687 ( .A1(n9498), .A2(n9815), .ZN(n9503) );
  AOI22_X1 U10688 ( .A1(n9500), .A2(n9742), .B1(n9598), .B2(n9499), .ZN(n9501)
         );
  OAI211_X1 U10689 ( .C1(n9217), .C2(n9503), .A(n9502), .B(n9501), .ZN(n9536)
         );
  MUX2_X1 U10690 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9536), .S(n9843), .Z(
        P1_U3541) );
  AOI22_X1 U10691 ( .A1(n9505), .A2(n9742), .B1(n9598), .B2(n9504), .ZN(n9506)
         );
  OAI211_X1 U10692 ( .C1(n9524), .C2(n9508), .A(n9507), .B(n9506), .ZN(n9537)
         );
  MUX2_X1 U10693 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9537), .S(n9843), .Z(
        P1_U3540) );
  AOI211_X1 U10694 ( .C1(n9598), .C2(n9511), .A(n9510), .B(n9509), .ZN(n9512)
         );
  OAI21_X1 U10695 ( .B1(n9524), .B2(n9513), .A(n9512), .ZN(n9538) );
  MUX2_X1 U10696 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9538), .S(n9843), .Z(
        P1_U3539) );
  AOI22_X1 U10697 ( .A1(n9515), .A2(n9742), .B1(n9598), .B2(n9514), .ZN(n9516)
         );
  OAI211_X1 U10698 ( .C1(n9587), .C2(n9518), .A(n9517), .B(n9516), .ZN(n9539)
         );
  MUX2_X1 U10699 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9539), .S(n9843), .Z(
        P1_U3538) );
  AOI211_X1 U10700 ( .C1(n9598), .C2(n9521), .A(n9520), .B(n9519), .ZN(n9522)
         );
  OAI21_X1 U10701 ( .B1(n9524), .B2(n9523), .A(n9522), .ZN(n9540) );
  MUX2_X1 U10702 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9540), .S(n9843), .Z(
        P1_U3537) );
  MUX2_X1 U10703 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9525), .S(n9828), .Z(
        P1_U3520) );
  MUX2_X1 U10704 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9526), .S(n9828), .Z(
        P1_U3519) );
  MUX2_X1 U10705 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9527), .S(n9828), .Z(
        P1_U3518) );
  MUX2_X1 U10706 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9528), .S(n9828), .Z(
        P1_U3517) );
  MUX2_X1 U10707 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9529), .S(n9828), .Z(
        P1_U3516) );
  MUX2_X1 U10708 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9530), .S(n9828), .Z(
        P1_U3515) );
  MUX2_X1 U10709 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9531), .S(n9828), .Z(
        P1_U3514) );
  MUX2_X1 U10710 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9532), .S(n9828), .Z(
        P1_U3513) );
  MUX2_X1 U10711 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9533), .S(n9828), .Z(
        P1_U3512) );
  MUX2_X1 U10712 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9534), .S(n9828), .Z(
        P1_U3511) );
  MUX2_X1 U10713 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9535), .S(n9828), .Z(
        P1_U3510) );
  MUX2_X1 U10714 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9536), .S(n9828), .Z(
        P1_U3508) );
  MUX2_X1 U10715 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9537), .S(n9828), .Z(
        P1_U3505) );
  MUX2_X1 U10716 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9538), .S(n9828), .Z(
        P1_U3502) );
  MUX2_X1 U10717 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9539), .S(n9828), .Z(
        P1_U3499) );
  MUX2_X1 U10718 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9540), .S(n9828), .Z(
        P1_U3496) );
  MUX2_X1 U10719 ( .A(P1_D_REG_1__SCAN_IN), .B(n9542), .S(n9541), .Z(P1_U3441)
         );
  INV_X1 U10720 ( .A(n9543), .ZN(n9549) );
  NOR4_X1 U10721 ( .A1(n9545), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9544), .A4(
        P1_U3084), .ZN(n9546) );
  AOI21_X1 U10722 ( .B1(n9547), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9546), .ZN(
        n9548) );
  OAI21_X1 U10723 ( .B1(n9549), .B2(n4249), .A(n9548), .ZN(P1_U3322) );
  AOI22_X1 U10724 ( .A1(n9850), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9562) );
  OAI21_X1 U10725 ( .B1(n9552), .B2(n9551), .A(n9550), .ZN(n9553) );
  INV_X1 U10726 ( .A(n9553), .ZN(n9554) );
  AOI22_X1 U10727 ( .A1(n9556), .A2(n9555), .B1(n9845), .B2(n9554), .ZN(n9561)
         );
  OAI211_X1 U10728 ( .C1(n9559), .C2(n9558), .A(n9844), .B(n9557), .ZN(n9560)
         );
  NAND3_X1 U10729 ( .A1(n9562), .A2(n9561), .A3(n9560), .ZN(P2_U3247) );
  NOR2_X1 U10730 ( .A1(n4525), .A2(n9817), .ZN(n9563) );
  INV_X1 U10731 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9565) );
  AOI22_X1 U10732 ( .A1(n9843), .A2(n9567), .B1(n9565), .B2(n9840), .ZN(
        P1_U3554) );
  INV_X1 U10733 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9566) );
  AOI22_X1 U10734 ( .A1(n9828), .A2(n9567), .B1(n9566), .B2(n9826), .ZN(
        P1_U3522) );
  OAI21_X1 U10735 ( .B1(n9569), .B2(n9983), .A(n9568), .ZN(n9570) );
  AOI21_X1 U10736 ( .B1(n9571), .B2(n9946), .A(n9570), .ZN(n9580) );
  AOI22_X1 U10737 ( .A1(n10008), .A2(n9580), .B1(n9572), .B2(n10006), .ZN(
        P2_U3550) );
  OAI22_X1 U10738 ( .A1(n9574), .A2(n9985), .B1(n9573), .B2(n9983), .ZN(n9576)
         );
  AOI211_X1 U10739 ( .C1(n9577), .C2(n9989), .A(n9576), .B(n9575), .ZN(n9581)
         );
  AOI22_X1 U10740 ( .A1(n10008), .A2(n9581), .B1(n9578), .B2(n10006), .ZN(
        P2_U3534) );
  AOI22_X1 U10741 ( .A1(n9993), .A2(n9580), .B1(n9579), .B2(n9991), .ZN(
        P2_U3518) );
  AOI22_X1 U10742 ( .A1(n9993), .A2(n9581), .B1(n5170), .B2(n9991), .ZN(
        P2_U3493) );
  NOR2_X1 U10743 ( .A1(n9582), .A2(n9819), .ZN(n9583) );
  INV_X1 U10744 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9586) );
  AOI22_X1 U10745 ( .A1(n9843), .A2(n9610), .B1(n9586), .B2(n9840), .ZN(
        P1_U3553) );
  INV_X1 U10746 ( .A(n9588), .ZN(n9593) );
  OAI22_X1 U10747 ( .A1(n9590), .A2(n9819), .B1(n9589), .B2(n9817), .ZN(n9592)
         );
  AOI211_X1 U10748 ( .C1(n9822), .C2(n9593), .A(n9592), .B(n9591), .ZN(n9612)
         );
  INV_X1 U10749 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9594) );
  AOI22_X1 U10750 ( .A1(n9843), .A2(n9612), .B1(n9594), .B2(n9840), .ZN(
        P1_U3536) );
  AOI211_X1 U10751 ( .C1(n9598), .C2(n9597), .A(n9596), .B(n9595), .ZN(n9601)
         );
  NAND3_X1 U10752 ( .A1(n7394), .A2(n9599), .A3(n9815), .ZN(n9600) );
  AOI22_X1 U10753 ( .A1(n9843), .A2(n9614), .B1(n6929), .B2(n9840), .ZN(
        P1_U3535) );
  INV_X1 U10754 ( .A(n9602), .ZN(n9607) );
  OAI22_X1 U10755 ( .A1(n9604), .A2(n9819), .B1(n9603), .B2(n9817), .ZN(n9606)
         );
  AOI211_X1 U10756 ( .C1(n9822), .C2(n9607), .A(n9606), .B(n9605), .ZN(n9616)
         );
  AOI22_X1 U10757 ( .A1(n9843), .A2(n9616), .B1(n9608), .B2(n9840), .ZN(
        P1_U3534) );
  INV_X1 U10758 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9609) );
  AOI22_X1 U10759 ( .A1(n9828), .A2(n9610), .B1(n9609), .B2(n9826), .ZN(
        P1_U3521) );
  INV_X1 U10760 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9611) );
  AOI22_X1 U10761 ( .A1(n9828), .A2(n9612), .B1(n9611), .B2(n9826), .ZN(
        P1_U3493) );
  INV_X1 U10762 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9613) );
  AOI22_X1 U10763 ( .A1(n9828), .A2(n9614), .B1(n9613), .B2(n9826), .ZN(
        P1_U3490) );
  AOI22_X1 U10764 ( .A1(n9828), .A2(n9616), .B1(n9615), .B2(n9826), .ZN(
        P1_U3487) );
  XNOR2_X1 U10765 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10766 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NOR2_X1 U10767 ( .A1(n9618), .A2(n9617), .ZN(n9623) );
  INV_X1 U10768 ( .A(n9619), .ZN(n9620) );
  OAI22_X1 U10769 ( .A1(n9621), .A2(n9620), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n9624), .ZN(n9622) );
  AOI22_X1 U10770 ( .A1(n9706), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(n9623), .B2(
        n9622), .ZN(n9626) );
  NAND3_X1 U10771 ( .A1(n9707), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9624), .ZN(
        n9625) );
  OAI211_X1 U10772 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n6809), .A(n9626), .B(
        n9625), .ZN(P1_U3241) );
  INV_X1 U10773 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9643) );
  OAI21_X1 U10774 ( .B1(n9629), .B2(n9628), .A(n9627), .ZN(n9630) );
  AOI22_X1 U10775 ( .A1(n9631), .A2(n9699), .B1(n9697), .B2(n9630), .ZN(n9642)
         );
  INV_X1 U10776 ( .A(n9632), .ZN(n9633) );
  NOR2_X1 U10777 ( .A1(n9634), .A2(n9633), .ZN(n9637) );
  OAI21_X1 U10778 ( .B1(n9637), .B2(n9636), .A(n9635), .ZN(n9640) );
  AOI211_X1 U10779 ( .C1(n9707), .C2(n9640), .A(n9639), .B(n9638), .ZN(n9641)
         );
  OAI211_X1 U10780 ( .C1(n9689), .C2(n9643), .A(n9642), .B(n9641), .ZN(
        P1_U3245) );
  OAI21_X1 U10781 ( .B1(n9646), .B2(n9645), .A(n9644), .ZN(n9654) );
  INV_X1 U10782 ( .A(n9647), .ZN(n9649) );
  AOI211_X1 U10783 ( .C1(n9651), .C2(n9650), .A(n9649), .B(n9648), .ZN(n9652)
         );
  AOI211_X1 U10784 ( .C1(n9697), .C2(n9654), .A(n9653), .B(n9652), .ZN(n9659)
         );
  INV_X1 U10785 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9656) );
  OAI22_X1 U10786 ( .A1(n9689), .A2(n9656), .B1(n9687), .B2(n9655), .ZN(n9657)
         );
  INV_X1 U10787 ( .A(n9657), .ZN(n9658) );
  NAND2_X1 U10788 ( .A1(n9659), .A2(n9658), .ZN(P1_U3246) );
  AOI21_X1 U10789 ( .B1(n9699), .B2(n9661), .A(n9660), .ZN(n9666) );
  OAI211_X1 U10790 ( .C1(n9664), .C2(n9663), .A(n9707), .B(n9662), .ZN(n9665)
         );
  AND2_X1 U10791 ( .A1(n9666), .A2(n9665), .ZN(n9673) );
  INV_X1 U10792 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9670) );
  XNOR2_X1 U10793 ( .A(n9668), .B(n9667), .ZN(n9669) );
  OAI22_X1 U10794 ( .A1(n9689), .A2(n9670), .B1(n9679), .B2(n9669), .ZN(n9671)
         );
  INV_X1 U10795 ( .A(n9671), .ZN(n9672) );
  NAND2_X1 U10796 ( .A1(n9673), .A2(n9672), .ZN(P1_U3249) );
  MUX2_X1 U10797 ( .A(n6496), .B(P1_REG1_REG_10__SCAN_IN), .S(n9674), .Z(n9675) );
  INV_X1 U10798 ( .A(n9675), .ZN(n9678) );
  OAI21_X1 U10799 ( .B1(n9678), .B2(n9677), .A(n9676), .ZN(n9685) );
  AOI211_X1 U10800 ( .C1(n9682), .C2(n9681), .A(n9680), .B(n9679), .ZN(n9683)
         );
  AOI211_X1 U10801 ( .C1(n9707), .C2(n9685), .A(n9684), .B(n9683), .ZN(n9692)
         );
  INV_X1 U10802 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9688) );
  OAI22_X1 U10803 ( .A1(n9689), .A2(n9688), .B1(n9687), .B2(n9686), .ZN(n9690)
         );
  INV_X1 U10804 ( .A(n9690), .ZN(n9691) );
  NAND2_X1 U10805 ( .A1(n9692), .A2(n9691), .ZN(P1_U3251) );
  AOI21_X1 U10806 ( .B1(n9695), .B2(n9694), .A(n9693), .ZN(n9696) );
  NAND2_X1 U10807 ( .A1(n9697), .A2(n9696), .ZN(n9702) );
  NAND2_X1 U10808 ( .A1(n9699), .A2(n9698), .ZN(n9701) );
  AND3_X1 U10809 ( .A1(n9702), .A2(n9701), .A3(n9700), .ZN(n9710) );
  OAI21_X1 U10810 ( .B1(n9705), .B2(n9704), .A(n9703), .ZN(n9708) );
  AOI22_X1 U10811 ( .A1(n9708), .A2(n9707), .B1(n9706), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n9709) );
  NAND2_X1 U10812 ( .A1(n9710), .A2(n9709), .ZN(P1_U3259) );
  XNOR2_X1 U10813 ( .A(n9712), .B(n9711), .ZN(n9730) );
  INV_X1 U10814 ( .A(n9730), .ZN(n9788) );
  NAND2_X1 U10815 ( .A1(n9714), .A2(n9713), .ZN(n9715) );
  NAND2_X1 U10816 ( .A1(n9716), .A2(n9715), .ZN(n9785) );
  INV_X1 U10817 ( .A(n9785), .ZN(n9717) );
  AOI22_X1 U10818 ( .A1(n9788), .A2(n9719), .B1(n9718), .B2(n9717), .ZN(n9736)
         );
  XNOR2_X1 U10819 ( .A(n9720), .B(n9721), .ZN(n9728) );
  OAI22_X1 U10820 ( .A1(n9725), .A2(n9724), .B1(n9723), .B2(n9722), .ZN(n9726)
         );
  AOI21_X1 U10821 ( .B1(n9728), .B2(n9727), .A(n9726), .ZN(n9729) );
  OAI21_X1 U10822 ( .B1(n9730), .B2(n9759), .A(n9729), .ZN(n9786) );
  AOI22_X1 U10823 ( .A1(n9234), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9747), .B2(
        n9731), .ZN(n9732) );
  OAI21_X1 U10824 ( .B1(n9784), .B2(n9733), .A(n9732), .ZN(n9734) );
  AOI21_X1 U10825 ( .B1(n9786), .B2(n9762), .A(n9734), .ZN(n9735) );
  NAND2_X1 U10826 ( .A1(n9736), .A2(n9735), .ZN(P1_U3288) );
  OAI21_X1 U10827 ( .B1(n9738), .B2(n9752), .A(n9737), .ZN(n9758) );
  INV_X1 U10828 ( .A(n9758), .ZN(n9776) );
  NAND2_X1 U10829 ( .A1(n9739), .A2(n6323), .ZN(n9772) );
  OAI21_X1 U10830 ( .B1(n6343), .B2(n9740), .A(n9772), .ZN(n9746) );
  OAI211_X1 U10831 ( .C1(n6343), .C2(n9743), .A(n9742), .B(n9741), .ZN(n9773)
         );
  NOR2_X1 U10832 ( .A1(n9773), .A2(n9744), .ZN(n9745) );
  AOI211_X1 U10833 ( .C1(n9747), .C2(P1_REG3_REG_1__SCAN_IN), .A(n9746), .B(
        n9745), .ZN(n9748) );
  INV_X1 U10834 ( .A(n9748), .ZN(n9760) );
  INV_X1 U10835 ( .A(n9749), .ZN(n9753) );
  AOI211_X1 U10836 ( .C1(n9753), .C2(n9752), .A(n9751), .B(n9750), .ZN(n9754)
         );
  AOI21_X1 U10837 ( .B1(n9756), .B2(n9755), .A(n9754), .ZN(n9757) );
  OAI21_X1 U10838 ( .B1(n9759), .B2(n9758), .A(n9757), .ZN(n9774) );
  AOI211_X1 U10839 ( .C1(n9761), .C2(n9776), .A(n9760), .B(n9774), .ZN(n9763)
         );
  AOI22_X1 U10840 ( .A1(n9234), .A2(n6277), .B1(n9763), .B2(n9762), .ZN(
        P1_U3290) );
  AND2_X1 U10841 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9771), .ZN(P1_U3292) );
  AND2_X1 U10842 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9771), .ZN(P1_U3293) );
  AND2_X1 U10843 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9771), .ZN(P1_U3294) );
  AND2_X1 U10844 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9771), .ZN(P1_U3295) );
  AND2_X1 U10845 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9771), .ZN(P1_U3296) );
  AND2_X1 U10846 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9771), .ZN(P1_U3297) );
  AND2_X1 U10847 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9771), .ZN(P1_U3298) );
  AND2_X1 U10848 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9771), .ZN(P1_U3299) );
  INV_X1 U10849 ( .A(n9771), .ZN(n9770) );
  NOR2_X1 U10850 ( .A1(n9770), .A2(n9766), .ZN(P1_U3300) );
  AND2_X1 U10851 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9771), .ZN(P1_U3301) );
  AND2_X1 U10852 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9771), .ZN(P1_U3302) );
  AND2_X1 U10853 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9771), .ZN(P1_U3303) );
  NOR2_X1 U10854 ( .A1(n9770), .A2(n9767), .ZN(P1_U3304) );
  AND2_X1 U10855 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9771), .ZN(P1_U3305) );
  AND2_X1 U10856 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9771), .ZN(P1_U3306) );
  NOR2_X1 U10857 ( .A1(n9770), .A2(n9768), .ZN(P1_U3307) );
  AND2_X1 U10858 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9771), .ZN(P1_U3308) );
  AND2_X1 U10859 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9771), .ZN(P1_U3309) );
  AND2_X1 U10860 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9771), .ZN(P1_U3310) );
  NOR2_X1 U10861 ( .A1(n9770), .A2(n9769), .ZN(P1_U3311) );
  AND2_X1 U10862 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9771), .ZN(P1_U3312) );
  AND2_X1 U10863 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9771), .ZN(P1_U3313) );
  AND2_X1 U10864 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9771), .ZN(P1_U3314) );
  AND2_X1 U10865 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9771), .ZN(P1_U3315) );
  AND2_X1 U10866 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9771), .ZN(P1_U3316) );
  AND2_X1 U10867 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9771), .ZN(P1_U3317) );
  AND2_X1 U10868 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9771), .ZN(P1_U3318) );
  AND2_X1 U10869 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9771), .ZN(P1_U3319) );
  AND2_X1 U10870 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9771), .ZN(P1_U3320) );
  AND2_X1 U10871 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9771), .ZN(P1_U3321) );
  OAI211_X1 U10872 ( .C1(n6343), .C2(n9817), .A(n9773), .B(n9772), .ZN(n9775)
         );
  AOI211_X1 U10873 ( .C1(n9822), .C2(n9776), .A(n9775), .B(n9774), .ZN(n9830)
         );
  INV_X1 U10874 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9777) );
  AOI22_X1 U10875 ( .A1(n9828), .A2(n9830), .B1(n9777), .B2(n9826), .ZN(
        P1_U3457) );
  OAI22_X1 U10876 ( .A1(n9779), .A2(n9819), .B1(n9778), .B2(n9817), .ZN(n9781)
         );
  AOI211_X1 U10877 ( .C1(n9822), .C2(n9782), .A(n9781), .B(n9780), .ZN(n9832)
         );
  INV_X1 U10878 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9783) );
  AOI22_X1 U10879 ( .A1(n9828), .A2(n9832), .B1(n9783), .B2(n9826), .ZN(
        P1_U3460) );
  OAI22_X1 U10880 ( .A1(n9785), .A2(n9819), .B1(n9784), .B2(n9817), .ZN(n9787)
         );
  AOI211_X1 U10881 ( .C1(n9822), .C2(n9788), .A(n9787), .B(n9786), .ZN(n9833)
         );
  INV_X1 U10882 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9789) );
  AOI22_X1 U10883 ( .A1(n9828), .A2(n9833), .B1(n9789), .B2(n9826), .ZN(
        P1_U3463) );
  INV_X1 U10884 ( .A(n9790), .ZN(n9795) );
  OAI22_X1 U10885 ( .A1(n9792), .A2(n9819), .B1(n9791), .B2(n9817), .ZN(n9794)
         );
  AOI211_X1 U10886 ( .C1(n9822), .C2(n9795), .A(n9794), .B(n9793), .ZN(n9834)
         );
  INV_X1 U10887 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9796) );
  AOI22_X1 U10888 ( .A1(n9828), .A2(n9834), .B1(n9796), .B2(n9826), .ZN(
        P1_U3466) );
  NAND3_X1 U10889 ( .A1(n6887), .A2(n9797), .A3(n9815), .ZN(n9799) );
  OAI211_X1 U10890 ( .C1(n9800), .C2(n9817), .A(n9799), .B(n9798), .ZN(n9801)
         );
  NOR2_X1 U10891 ( .A1(n9802), .A2(n9801), .ZN(n9836) );
  INV_X1 U10892 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9803) );
  AOI22_X1 U10893 ( .A1(n9828), .A2(n9836), .B1(n9803), .B2(n9826), .ZN(
        P1_U3469) );
  OAI22_X1 U10894 ( .A1(n9805), .A2(n9819), .B1(n9804), .B2(n9817), .ZN(n9807)
         );
  AOI211_X1 U10895 ( .C1(n9815), .C2(n9808), .A(n9807), .B(n9806), .ZN(n9837)
         );
  INV_X1 U10896 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9809) );
  AOI22_X1 U10897 ( .A1(n9828), .A2(n9837), .B1(n9809), .B2(n9826), .ZN(
        P1_U3472) );
  OAI211_X1 U10898 ( .C1(n9812), .C2(n9817), .A(n9811), .B(n9810), .ZN(n9813)
         );
  AOI21_X1 U10899 ( .B1(n9815), .B2(n9814), .A(n9813), .ZN(n9839) );
  INV_X1 U10900 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9816) );
  AOI22_X1 U10901 ( .A1(n9828), .A2(n9839), .B1(n9816), .B2(n9826), .ZN(
        P1_U3475) );
  OAI22_X1 U10902 ( .A1(n9820), .A2(n9819), .B1(n9818), .B2(n9817), .ZN(n9821)
         );
  AOI21_X1 U10903 ( .B1(n9823), .B2(n9822), .A(n9821), .ZN(n9824) );
  INV_X1 U10904 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9827) );
  AOI22_X1 U10905 ( .A1(n9828), .A2(n9842), .B1(n9827), .B2(n9826), .ZN(
        P1_U3481) );
  AOI22_X1 U10906 ( .A1(n9843), .A2(n9830), .B1(n9829), .B2(n9840), .ZN(
        P1_U3524) );
  AOI22_X1 U10907 ( .A1(n9843), .A2(n9832), .B1(n9831), .B2(n9840), .ZN(
        P1_U3525) );
  AOI22_X1 U10908 ( .A1(n9843), .A2(n9833), .B1(n6289), .B2(n9840), .ZN(
        P1_U3526) );
  AOI22_X1 U10909 ( .A1(n9843), .A2(n9834), .B1(n6292), .B2(n9840), .ZN(
        P1_U3527) );
  INV_X1 U10910 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9835) );
  AOI22_X1 U10911 ( .A1(n9843), .A2(n9836), .B1(n9835), .B2(n9840), .ZN(
        P1_U3528) );
  AOI22_X1 U10912 ( .A1(n9843), .A2(n9837), .B1(n6296), .B2(n9840), .ZN(
        P1_U3529) );
  INV_X1 U10913 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9838) );
  AOI22_X1 U10914 ( .A1(n9843), .A2(n9839), .B1(n9838), .B2(n9840), .ZN(
        P1_U3530) );
  INV_X1 U10915 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9841) );
  AOI22_X1 U10916 ( .A1(n9843), .A2(n9842), .B1(n9841), .B2(n9840), .ZN(
        P1_U3532) );
  AOI22_X1 U10917 ( .A1(n9844), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9845), .ZN(n9853) );
  NAND2_X1 U10918 ( .A1(n9845), .A2(n9994), .ZN(n9846) );
  OAI211_X1 U10919 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n9848), .A(n9847), .B(
        n9846), .ZN(n9849) );
  INV_X1 U10920 ( .A(n9849), .ZN(n9852) );
  AOI22_X1 U10921 ( .A1(n9850), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9851) );
  OAI221_X1 U10922 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9853), .C1(n4410), .C2(
        n9852), .A(n9851), .ZN(P2_U3245) );
  INV_X1 U10923 ( .A(n9854), .ZN(n9868) );
  XNOR2_X1 U10924 ( .A(n9856), .B(n9855), .ZN(n9941) );
  OR2_X1 U10925 ( .A1(n9858), .A2(n9857), .ZN(n9859) );
  NAND2_X1 U10926 ( .A1(n9860), .A2(n9859), .ZN(n9866) );
  OAI22_X1 U10927 ( .A1(n6708), .A2(n9863), .B1(n9862), .B2(n9861), .ZN(n9864)
         );
  AOI21_X1 U10928 ( .B1(n9866), .B2(n9865), .A(n9864), .ZN(n9944) );
  INV_X1 U10929 ( .A(n9944), .ZN(n9867) );
  AOI21_X1 U10930 ( .B1(n9868), .B2(n9941), .A(n9867), .ZN(n9881) );
  AOI22_X1 U10931 ( .A1(n9869), .A2(n4922), .B1(P2_REG2_REG_3__SCAN_IN), .B2(
        n4247), .ZN(n9880) );
  OAI211_X1 U10932 ( .C1(n9872), .C2(n9871), .A(n9870), .B(n9946), .ZN(n9875)
         );
  NAND2_X1 U10933 ( .A1(n9873), .A2(n9954), .ZN(n9874) );
  NAND2_X1 U10934 ( .A1(n9875), .A2(n9874), .ZN(n9940) );
  INV_X1 U10935 ( .A(n9876), .ZN(n9877) );
  AOI22_X1 U10936 ( .A1(n9878), .A2(n9940), .B1(n9877), .B2(n9941), .ZN(n9879)
         );
  OAI211_X1 U10937 ( .C1(n4247), .C2(n9881), .A(n9880), .B(n9879), .ZN(
        P2_U3293) );
  INV_X1 U10938 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n9884) );
  NOR2_X1 U10939 ( .A1(n9919), .A2(n9884), .ZN(P2_U3297) );
  INV_X1 U10940 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n9885) );
  NOR2_X1 U10941 ( .A1(n9919), .A2(n9885), .ZN(P2_U3298) );
  NOR2_X1 U10942 ( .A1(n9919), .A2(n9886), .ZN(P2_U3299) );
  INV_X1 U10943 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n9887) );
  NOR2_X1 U10944 ( .A1(n9919), .A2(n9887), .ZN(P2_U3300) );
  INV_X1 U10945 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n9888) );
  NOR2_X1 U10946 ( .A1(n9898), .A2(n9888), .ZN(P2_U3301) );
  INV_X1 U10947 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n9889) );
  NOR2_X1 U10948 ( .A1(n9898), .A2(n9889), .ZN(P2_U3302) );
  INV_X1 U10949 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9890) );
  NOR2_X1 U10950 ( .A1(n9898), .A2(n9890), .ZN(P2_U3303) );
  INV_X1 U10951 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n9891) );
  NOR2_X1 U10952 ( .A1(n9898), .A2(n9891), .ZN(P2_U3304) );
  INV_X1 U10953 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n9892) );
  NOR2_X1 U10954 ( .A1(n9898), .A2(n9892), .ZN(P2_U3305) );
  NOR2_X1 U10955 ( .A1(n9898), .A2(n9893), .ZN(P2_U3306) );
  INV_X1 U10956 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n9894) );
  NOR2_X1 U10957 ( .A1(n9898), .A2(n9894), .ZN(P2_U3307) );
  INV_X1 U10958 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n9895) );
  NOR2_X1 U10959 ( .A1(n9898), .A2(n9895), .ZN(P2_U3308) );
  INV_X1 U10960 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n9896) );
  NOR2_X1 U10961 ( .A1(n9898), .A2(n9896), .ZN(P2_U3309) );
  INV_X1 U10962 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n9897) );
  NOR2_X1 U10963 ( .A1(n9898), .A2(n9897), .ZN(P2_U3310) );
  INV_X1 U10964 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n9899) );
  NOR2_X1 U10965 ( .A1(n9919), .A2(n9899), .ZN(P2_U3311) );
  INV_X1 U10966 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9900) );
  NOR2_X1 U10967 ( .A1(n9919), .A2(n9900), .ZN(P2_U3312) );
  NOR2_X1 U10968 ( .A1(n9919), .A2(n9901), .ZN(P2_U3313) );
  INV_X1 U10969 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n9902) );
  NOR2_X1 U10970 ( .A1(n9919), .A2(n9902), .ZN(P2_U3314) );
  INV_X1 U10971 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n9903) );
  NOR2_X1 U10972 ( .A1(n9919), .A2(n9903), .ZN(P2_U3315) );
  INV_X1 U10973 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n9904) );
  NOR2_X1 U10974 ( .A1(n9919), .A2(n9904), .ZN(P2_U3316) );
  NOR2_X1 U10975 ( .A1(n9919), .A2(n9905), .ZN(P2_U3317) );
  INV_X1 U10976 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n9906) );
  NOR2_X1 U10977 ( .A1(n9919), .A2(n9906), .ZN(P2_U3318) );
  NOR2_X1 U10978 ( .A1(n9919), .A2(n9907), .ZN(P2_U3319) );
  INV_X1 U10979 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n9908) );
  NOR2_X1 U10980 ( .A1(n9919), .A2(n9908), .ZN(P2_U3320) );
  INV_X1 U10981 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n9909) );
  NOR2_X1 U10982 ( .A1(n9919), .A2(n9909), .ZN(P2_U3321) );
  INV_X1 U10983 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n9910) );
  NOR2_X1 U10984 ( .A1(n9919), .A2(n9910), .ZN(P2_U3322) );
  NOR2_X1 U10985 ( .A1(n9919), .A2(n9911), .ZN(P2_U3323) );
  INV_X1 U10986 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n9912) );
  NOR2_X1 U10987 ( .A1(n9919), .A2(n9912), .ZN(P2_U3324) );
  INV_X1 U10988 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n9913) );
  NOR2_X1 U10989 ( .A1(n9919), .A2(n9913), .ZN(P2_U3325) );
  NOR2_X1 U10990 ( .A1(n9919), .A2(n9914), .ZN(P2_U3326) );
  OAI22_X1 U10991 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n9919), .B1(n9918), .B2(
        n9915), .ZN(n9916) );
  INV_X1 U10992 ( .A(n9916), .ZN(P2_U3437) );
  OAI22_X1 U10993 ( .A1(P2_D_REG_1__SCAN_IN), .A2(n9919), .B1(n9918), .B2(
        n9917), .ZN(n9920) );
  INV_X1 U10994 ( .A(n9920), .ZN(P2_U3438) );
  OAI22_X1 U10995 ( .A1(n9923), .A2(n9957), .B1(n9922), .B2(n9921), .ZN(n9925)
         );
  NOR2_X1 U10996 ( .A1(n9925), .A2(n9924), .ZN(n9995) );
  INV_X1 U10997 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9926) );
  AOI22_X1 U10998 ( .A1(n9993), .A2(n9995), .B1(n9926), .B2(n9991), .ZN(
        P2_U3451) );
  INV_X1 U10999 ( .A(n9927), .ZN(n9928) );
  OAI21_X1 U11000 ( .B1(n9929), .B2(n9983), .A(n9928), .ZN(n9932) );
  INV_X1 U11001 ( .A(n9930), .ZN(n9931) );
  AOI211_X1 U11002 ( .C1(n9989), .C2(n9933), .A(n9932), .B(n9931), .ZN(n9996)
         );
  AOI22_X1 U11003 ( .A1(n9993), .A2(n9996), .B1(n4827), .B2(n9991), .ZN(
        P2_U3454) );
  INV_X1 U11004 ( .A(n9934), .ZN(n9935) );
  OAI211_X1 U11005 ( .C1(n9937), .C2(n9983), .A(n9936), .B(n9935), .ZN(n9938)
         );
  AOI21_X1 U11006 ( .B1(n9989), .B2(n9939), .A(n9938), .ZN(n9997) );
  AOI22_X1 U11007 ( .A1(n9993), .A2(n9997), .B1(n4884), .B2(n9991), .ZN(
        P2_U3457) );
  INV_X1 U11008 ( .A(n9940), .ZN(n9943) );
  NAND2_X1 U11009 ( .A1(n9941), .A2(n9989), .ZN(n9942) );
  AND3_X1 U11010 ( .A1(n9944), .A2(n9943), .A3(n9942), .ZN(n9998) );
  AOI22_X1 U11011 ( .A1(n9993), .A2(n9998), .B1(n4905), .B2(n9991), .ZN(
        P2_U3460) );
  AOI22_X1 U11012 ( .A1(n9947), .A2(n9946), .B1(n9954), .B2(n9945), .ZN(n9948)
         );
  OAI211_X1 U11013 ( .C1(n9950), .C2(n9957), .A(n9949), .B(n9948), .ZN(n9951)
         );
  INV_X1 U11014 ( .A(n9951), .ZN(n9999) );
  AOI22_X1 U11015 ( .A1(n9993), .A2(n9999), .B1(n4920), .B2(n9991), .ZN(
        P2_U3463) );
  AOI21_X1 U11016 ( .B1(n9954), .B2(n9953), .A(n9952), .ZN(n9955) );
  OAI211_X1 U11017 ( .C1(n9958), .C2(n9957), .A(n9956), .B(n9955), .ZN(n9959)
         );
  INV_X1 U11018 ( .A(n9959), .ZN(n10001) );
  AOI22_X1 U11019 ( .A1(n9993), .A2(n10001), .B1(n4963), .B2(n9991), .ZN(
        P2_U3466) );
  OAI22_X1 U11020 ( .A1(n9961), .A2(n9985), .B1(n9960), .B2(n9983), .ZN(n9962)
         );
  INV_X1 U11021 ( .A(n9962), .ZN(n9965) );
  NAND2_X1 U11022 ( .A1(n9963), .A2(n9989), .ZN(n9964) );
  AND3_X1 U11023 ( .A1(n9966), .A2(n9965), .A3(n9964), .ZN(n10002) );
  AOI22_X1 U11024 ( .A1(n9993), .A2(n10002), .B1(n4984), .B2(n9991), .ZN(
        P2_U3469) );
  INV_X1 U11025 ( .A(n9967), .ZN(n9981) );
  INV_X1 U11026 ( .A(n9968), .ZN(n9974) );
  INV_X1 U11027 ( .A(n9969), .ZN(n9970) );
  OAI22_X1 U11028 ( .A1(n9971), .A2(n9985), .B1(n9970), .B2(n9983), .ZN(n9973)
         );
  AOI211_X1 U11029 ( .C1(n9981), .C2(n9974), .A(n9973), .B(n9972), .ZN(n10004)
         );
  AOI22_X1 U11030 ( .A1(n9993), .A2(n10004), .B1(n9451), .B2(n9991), .ZN(
        P2_U3475) );
  INV_X1 U11031 ( .A(n9975), .ZN(n9980) );
  OAI22_X1 U11032 ( .A1(n9977), .A2(n9985), .B1(n4416), .B2(n9983), .ZN(n9979)
         );
  AOI211_X1 U11033 ( .C1(n9981), .C2(n9980), .A(n9979), .B(n9978), .ZN(n10005)
         );
  INV_X1 U11034 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9982) );
  AOI22_X1 U11035 ( .A1(n9993), .A2(n10005), .B1(n9982), .B2(n9991), .ZN(
        P2_U3481) );
  OAI22_X1 U11036 ( .A1(n9986), .A2(n9985), .B1(n9984), .B2(n9983), .ZN(n9988)
         );
  AOI211_X1 U11037 ( .C1(n9990), .C2(n9989), .A(n9988), .B(n9987), .ZN(n10007)
         );
  INV_X1 U11038 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9992) );
  AOI22_X1 U11039 ( .A1(n9993), .A2(n10007), .B1(n9992), .B2(n9991), .ZN(
        P2_U3487) );
  AOI22_X1 U11040 ( .A1(n10008), .A2(n9995), .B1(n9994), .B2(n10006), .ZN(
        P2_U3520) );
  AOI22_X1 U11041 ( .A1(n10008), .A2(n9996), .B1(n4830), .B2(n10006), .ZN(
        P2_U3521) );
  AOI22_X1 U11042 ( .A1(n10008), .A2(n9997), .B1(n4885), .B2(n10006), .ZN(
        P2_U3522) );
  AOI22_X1 U11043 ( .A1(n10008), .A2(n9998), .B1(n6539), .B2(n10006), .ZN(
        P2_U3523) );
  AOI22_X1 U11044 ( .A1(n10008), .A2(n9999), .B1(n6541), .B2(n10006), .ZN(
        P2_U3524) );
  INV_X1 U11045 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10000) );
  AOI22_X1 U11046 ( .A1(n10008), .A2(n10001), .B1(n10000), .B2(n10006), .ZN(
        P2_U3525) );
  AOI22_X1 U11047 ( .A1(n10008), .A2(n10002), .B1(n6545), .B2(n10006), .ZN(
        P2_U3526) );
  AOI22_X1 U11048 ( .A1(n10008), .A2(n10004), .B1(n10003), .B2(n10006), .ZN(
        P2_U3528) );
  AOI22_X1 U11049 ( .A1(n10008), .A2(n10005), .B1(n5075), .B2(n10006), .ZN(
        P2_U3530) );
  AOI22_X1 U11050 ( .A1(n10008), .A2(n10007), .B1(n6553), .B2(n10006), .ZN(
        P2_U3532) );
  INV_X1 U11051 ( .A(n10009), .ZN(n10010) );
  NAND2_X1 U11052 ( .A1(n10011), .A2(n10010), .ZN(n10012) );
  XNOR2_X1 U11053 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10012), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11054 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11055 ( .B1(n10015), .B2(n10014), .A(n10013), .ZN(ADD_1071_U56) );
  OAI21_X1 U11056 ( .B1(n10018), .B2(n10017), .A(n10016), .ZN(ADD_1071_U57) );
  OAI21_X1 U11057 ( .B1(n10021), .B2(n10020), .A(n10019), .ZN(ADD_1071_U58) );
  OAI21_X1 U11058 ( .B1(n10024), .B2(n10023), .A(n10022), .ZN(ADD_1071_U59) );
  OAI21_X1 U11059 ( .B1(n10027), .B2(n10026), .A(n10025), .ZN(ADD_1071_U60) );
  OAI21_X1 U11060 ( .B1(n10030), .B2(n10029), .A(n10028), .ZN(ADD_1071_U61) );
  AOI21_X1 U11061 ( .B1(n10033), .B2(n10032), .A(n10031), .ZN(ADD_1071_U62) );
  AOI21_X1 U11062 ( .B1(n10036), .B2(n10035), .A(n10034), .ZN(ADD_1071_U63) );
  XOR2_X1 U11063 ( .A(n10037), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11064 ( .A1(n10039), .A2(n10038), .ZN(n10040) );
  XOR2_X1 U11065 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10040), .Z(ADD_1071_U51) );
  XOR2_X1 U11066 ( .A(n10041), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  OAI21_X1 U11067 ( .B1(n10044), .B2(n10043), .A(n10042), .ZN(n10045) );
  XNOR2_X1 U11068 ( .A(n10045), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11069 ( .B1(n10048), .B2(n10047), .A(n10046), .ZN(ADD_1071_U47) );
  AOI21_X1 U11070 ( .B1(n10051), .B2(n10050), .A(n10049), .ZN(ADD_1071_U48) );
  XOR2_X1 U11071 ( .A(n10053), .B(n10052), .Z(ADD_1071_U54) );
  XOR2_X1 U11072 ( .A(n10055), .B(n10054), .Z(ADD_1071_U53) );
  XNOR2_X1 U11073 ( .A(n10057), .B(n10056), .ZN(ADD_1071_U52) );
  CLKBUF_X3 U4754 ( .A(n4958), .Z(n7743) );
  CLKBUF_X1 U4772 ( .A(n4873), .Z(n5438) );
  XNOR2_X1 U5373 ( .A(n4824), .B(P2_IR_REG_30__SCAN_IN), .ZN(n4831) );
  CLKBUF_X1 U6037 ( .A(n6205), .Z(n4246) );
  NAND2_X1 U6295 ( .A1(n6070), .A2(n4628), .ZN(n10060) );
endmodule

