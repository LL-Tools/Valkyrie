

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10744;

  AND2_X1 U4993 ( .A1(n9895), .A2(n9898), .ZN(n9992) );
  AND2_X1 U4994 ( .A1(n8362), .A2(n8358), .ZN(n8356) );
  INV_X1 U4995 ( .A(n5633), .ZN(n5662) );
  CLKBUF_X1 U4996 ( .A(n5753), .Z(n6446) );
  CLKBUF_X2 U4997 ( .A(n6864), .Z(n8291) );
  CLKBUF_X2 U4998 ( .A(n6990), .Z(n7587) );
  NAND4_X1 U4999 ( .A1(n5659), .A2(n5658), .A3(n5657), .A4(n5656), .ZN(n5664)
         );
  NAND4_X1 U5000 ( .A1(n5676), .A2(n5675), .A3(n5674), .A4(n5673), .ZN(n5692)
         );
  INV_X1 U5001 ( .A(n6644), .ZN(n6725) );
  CLKBUF_X1 U5002 ( .A(n6746), .Z(n4931) );
  INV_X1 U5004 ( .A(n10744), .ZN(n4930) );
  INV_X1 U5005 ( .A(n7674), .ZN(n8344) );
  NAND2_X1 U5006 ( .A1(n7233), .A2(n7232), .ZN(n7274) );
  NAND2_X1 U5007 ( .A1(n5648), .A2(n8278), .ZN(n5735) );
  INV_X1 U5008 ( .A(n8859), .ZN(n8879) );
  INV_X1 U5009 ( .A(n8491), .ZN(n8492) );
  INV_X1 U5010 ( .A(n6291), .ZN(n6247) );
  NAND2_X2 U5012 ( .A1(n6478), .A2(n6482), .ZN(n8249) );
  AND2_X1 U5014 ( .A1(n5499), .A2(n9644), .ZN(n9645) );
  XNOR2_X1 U5015 ( .A(n5593), .B(n5592), .ZN(n5609) );
  INV_X2 U5016 ( .A(n6572), .ZN(n8825) );
  OR2_X1 U5017 ( .A1(n9616), .A2(n9826), .ZN(n9895) );
  OAI21_X2 U5018 ( .B1(n5815), .B2(n5478), .A(n5476), .ZN(n5475) );
  AOI21_X2 U5019 ( .B1(n5298), .B2(n8989), .A(n8257), .ZN(n9013) );
  NOR4_X2 U5020 ( .A1(n8876), .A2(n8867), .A3(n8459), .A4(n8330), .ZN(n8331)
         );
  OAI22_X2 U5021 ( .A1(n8511), .A2(n5364), .B1(n5366), .B2(n8516), .ZN(n8688)
         );
  AOI211_X2 U5022 ( .C1(n9891), .C2(n9688), .A(n9687), .B(n9686), .ZN(n9689)
         );
  OAI22_X2 U5023 ( .A1(n9873), .A2(n9872), .B1(n9975), .B2(n9889), .ZN(n9854)
         );
  AOI21_X2 U5024 ( .B1(n9634), .B2(n9633), .A(n5237), .ZN(n9873) );
  AOI21_X2 U5025 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6705), .A(n6704), .ZN(
        n6790) );
  XNOR2_X2 U5026 ( .A(n6372), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6428) );
  XNOR2_X2 U5027 ( .A(n6397), .B(n6396), .ZN(n7064) );
  AOI22_X2 U5028 ( .A1(P1_REG2_REG_1__SCAN_IN), .A2(n6725), .B1(n6644), .B2(
        n5655), .ZN(n6717) );
  XNOR2_X1 U5029 ( .A(n6391), .B(n6390), .ZN(n6746) );
  XNOR2_X2 U5030 ( .A(n5649), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6644) );
  NAND2_X1 U5031 ( .A1(n8080), .A2(n8053), .ZN(n8052) );
  NAND2_X1 U5032 ( .A1(n7514), .A2(n7442), .ZN(n9403) );
  INV_X1 U5033 ( .A(n7214), .ZN(n7507) );
  INV_X1 U5034 ( .A(n8713), .ZN(n7315) );
  CLKBUF_X2 U5035 ( .A(n5653), .Z(n5083) );
  NAND2_X2 U5036 ( .A1(n7081), .A2(n7072), .ZN(n8349) );
  INV_X1 U5037 ( .A(n8716), .ZN(n7081) );
  INV_X1 U5038 ( .A(n5692), .ZN(n7203) );
  INV_X1 U5039 ( .A(n6997), .ZN(n7078) );
  CLKBUF_X2 U5040 ( .A(n6743), .Z(n8208) );
  CLKBUF_X2 U5041 ( .A(n5671), .Z(n6283) );
  NAND2_X1 U5042 ( .A1(n6638), .A2(n5567), .ZN(n5571) );
  NAND2_X1 U5043 ( .A1(n5323), .A2(n6934), .ZN(n5322) );
  CLKBUF_X1 U5044 ( .A(n6373), .Z(n6374) );
  AND2_X1 U5045 ( .A1(n5547), .A2(n4964), .ZN(n5546) );
  INV_X1 U5046 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6414) );
  OAI21_X1 U5047 ( .B1(n8535), .B2(n5375), .A(n4971), .ZN(n8596) );
  AND2_X1 U5048 ( .A1(n8245), .A2(n8244), .ZN(n8246) );
  NAND2_X1 U5049 ( .A1(n5324), .A2(n8819), .ZN(n8778) );
  NAND2_X1 U5050 ( .A1(n5147), .A2(n5146), .ZN(n9805) );
  AND2_X1 U5051 ( .A1(n9653), .A2(n9492), .ZN(n9793) );
  OR2_X1 U5052 ( .A1(n7609), .A2(n5345), .ZN(n5342) );
  NAND2_X1 U5053 ( .A1(n8199), .A2(n8198), .ZN(n8700) );
  AND2_X1 U5054 ( .A1(n7748), .A2(n7747), .ZN(n7861) );
  OR2_X1 U5055 ( .A1(n7628), .A2(n7627), .ZN(n7748) );
  AOI21_X1 U5056 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n7623), .A(n7622), .ZN(
        n7628) );
  NOR2_X1 U5057 ( .A1(n8767), .A2(n8766), .ZN(n8768) );
  AND2_X1 U5058 ( .A1(n5307), .A2(n5306), .ZN(n8733) );
  NAND2_X1 U5059 ( .A1(n5835), .A2(n5834), .ZN(n7676) );
  INV_X1 U5060 ( .A(n7483), .ZN(n7277) );
  AND2_X1 U5061 ( .A1(n7128), .A2(n5090), .ZN(n7483) );
  OAI211_X1 U5062 ( .C1(n5086), .C2(n6665), .A(n5772), .B(n5771), .ZN(n7432)
         );
  INV_X1 U5063 ( .A(n6861), .ZN(n6592) );
  NAND2_X1 U5064 ( .A1(n5810), .A2(n5036), .ZN(n7235) );
  NAND2_X2 U5065 ( .A1(n6591), .A2(n6590), .ZN(n6861) );
  OR2_X1 U5066 ( .A1(n7059), .A2(n7058), .ZN(n7186) );
  NAND2_X1 U5067 ( .A1(n5765), .A2(n5764), .ZN(n5769) );
  INV_X1 U5069 ( .A(n6879), .ZN(n10548) );
  NAND2_X1 U5070 ( .A1(n5734), .A2(n5733), .ZN(n5765) );
  BUF_X2 U5071 ( .A(n6865), .Z(n8159) );
  AND2_X1 U5072 ( .A1(n6525), .A2(n9153), .ZN(n6864) );
  NAND2_X2 U5073 ( .A1(n8344), .A2(n8505), .ZN(n8491) );
  OAI21_X1 U5074 ( .B1(n5480), .B2(n5479), .A(n4987), .ZN(n5477) );
  NAND4_X1 U5075 ( .A1(n5625), .A2(n5624), .A3(n5623), .A4(n5622), .ZN(n6474)
         );
  XNOR2_X1 U5076 ( .A(n6415), .B(n6414), .ZN(n7674) );
  AND2_X1 U5077 ( .A1(n5792), .A2(n5109), .ZN(n5289) );
  NAND2_X1 U5078 ( .A1(n6379), .A2(n6374), .ZN(n7957) );
  NAND2_X1 U5079 ( .A1(n9148), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6521) );
  NAND2_X2 U5080 ( .A1(n5571), .A2(n5570), .ZN(n5648) );
  OR2_X1 U5081 ( .A1(n5482), .A2(n5479), .ZN(n5478) );
  INV_X1 U5082 ( .A(n5753), .ZN(n4932) );
  AND2_X1 U5083 ( .A1(n5809), .A2(n5791), .ZN(n5792) );
  INV_X1 U5084 ( .A(n6377), .ZN(n6387) );
  XNOR2_X1 U5085 ( .A(n5618), .B(n5617), .ZN(n10279) );
  NAND2_X1 U5086 ( .A1(n5358), .A2(n5360), .ZN(n6373) );
  AND3_X1 U5087 ( .A1(n5356), .A2(n6367), .A3(n6368), .ZN(n5360) );
  NAND3_X1 U5088 ( .A1(n5957), .A2(n5548), .A3(n5612), .ZN(n5569) );
  INV_X2 U5089 ( .A(n9150), .ZN(n9156) );
  OR2_X1 U5090 ( .A1(n7134), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7241) );
  INV_X8 U5091 ( .A(n8278), .ZN(n6594) );
  AND2_X1 U5092 ( .A1(n5566), .A2(n5549), .ZN(n5548) );
  AND3_X1 U5093 ( .A1(n5440), .A2(n5359), .A3(n6395), .ZN(n5358) );
  AND2_X2 U5094 ( .A1(n6389), .A2(n6390), .ZN(n6395) );
  NOR2_X1 U5095 ( .A1(n6370), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U5096 ( .A1(n5573), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5485) );
  AND4_X1 U5097 ( .A1(n5244), .A2(n5245), .A3(n5246), .A4(n5557), .ZN(n5817)
         );
  INV_X1 U5098 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6026) );
  INV_X1 U5099 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7042) );
  INV_X1 U5100 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5592) );
  NOR2_X1 U5101 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5583) );
  INV_X1 U5102 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5594) );
  INV_X4 U5103 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5104 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6316) );
  INV_X1 U5105 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6583) );
  NOR2_X1 U5106 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5245) );
  NOR2_X1 U5107 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5246) );
  INV_X1 U5108 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7084) );
  INV_X1 U5109 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6455) );
  NOR2_X1 U5110 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5547) );
  NOR2_X1 U5111 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n6365) );
  NOR2_X1 U5112 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n6366) );
  INV_X1 U5113 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6390) );
  INV_X1 U5114 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7285) );
  INV_X1 U5115 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6548) );
  INV_X1 U5116 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6970) );
  INV_X1 U5117 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n6520) );
  NOR2_X1 U5118 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5244) );
  OAI21_X2 U5119 ( .B1(n8875), .B2(n8468), .A(n8307), .ZN(n8865) );
  OAI21_X4 U5120 ( .B1(n9342), .B2(n5250), .A(n5248), .ZN(n9835) );
  NAND2_X2 U5121 ( .A1(n9341), .A2(n9378), .ZN(n9342) );
  INV_X4 U5122 ( .A(n6592), .ZN(n8552) );
  OAI22_X2 U5123 ( .A1(n8016), .A2(n9451), .B1(n9987), .B2(n7969), .ZN(n9634)
         );
  CLKBUF_X3 U5124 ( .A(n6741), .Z(n8187) );
  OR2_X1 U5125 ( .A1(n8259), .A2(n8846), .ZN(n8494) );
  INV_X1 U5126 ( .A(n9501), .ZN(n5116) );
  NAND2_X1 U5127 ( .A1(n8554), .A2(n5101), .ZN(n8475) );
  INV_X1 U5128 ( .A(n9080), .ZN(n5101) );
  OR2_X1 U5129 ( .A1(n9123), .A2(n8945), .ZN(n8434) );
  NOR2_X1 U5130 ( .A1(n5361), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n5359) );
  INV_X1 U5131 ( .A(n9245), .ZN(n5406) );
  AND2_X1 U5132 ( .A1(n5626), .A2(n6363), .ZN(n5082) );
  NAND2_X1 U5133 ( .A1(n5569), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6332) );
  AOI21_X1 U5134 ( .B1(n5465), .B2(n5463), .A(n5018), .ZN(n5462) );
  INV_X1 U5135 ( .A(n6157), .ZN(n5463) );
  NAND2_X1 U5136 ( .A1(n5489), .A2(n5488), .ZN(n6127) );
  AOI21_X1 U5137 ( .B1(n4939), .B2(n5492), .A(n5019), .ZN(n5488) );
  NAND2_X1 U5138 ( .A1(n8501), .A2(n5427), .ZN(n5426) );
  NAND2_X1 U5139 ( .A1(n5429), .A2(n7674), .ZN(n5427) );
  AND2_X1 U5140 ( .A1(n6525), .A2(n6526), .ZN(n6865) );
  AND2_X1 U5141 ( .A1(n8508), .A2(n6526), .ZN(n6990) );
  NAND2_X1 U5142 ( .A1(n8299), .A2(n8242), .ZN(n8842) );
  INV_X1 U5143 ( .A(n8187), .ZN(n8288) );
  NAND2_X1 U5144 ( .A1(n5113), .A2(n5115), .ZN(n5112) );
  INV_X1 U5145 ( .A(n9504), .ZN(n5126) );
  INV_X1 U5146 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6410) );
  INV_X1 U5147 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6371) );
  NOR2_X1 U5148 ( .A1(n8543), .A2(n5377), .ZN(n5376) );
  INV_X1 U5149 ( .A(n8538), .ZN(n5377) );
  NAND2_X1 U5150 ( .A1(n7891), .A2(n7893), .ZN(n5335) );
  AND2_X1 U5151 ( .A1(n8522), .A2(n5021), .ZN(n5354) );
  INV_X1 U5152 ( .A(n5316), .ZN(n5313) );
  INV_X1 U5153 ( .A(n5315), .ZN(n5314) );
  OAI21_X1 U5154 ( .B1(n7183), .B2(n4934), .A(n7393), .ZN(n5315) );
  NAND2_X1 U5155 ( .A1(n7186), .A2(n7184), .ZN(n7182) );
  OR2_X1 U5156 ( .A1(n10467), .A2(n5325), .ZN(n5324) );
  NOR2_X1 U5157 ( .A1(n10457), .A2(n8776), .ZN(n5325) );
  INV_X1 U5158 ( .A(n8233), .ZN(n5434) );
  OR2_X1 U5159 ( .A1(n9074), .A2(n8237), .ZN(n8299) );
  OR2_X1 U5160 ( .A1(n8632), .A2(n8898), .ZN(n8464) );
  OR2_X1 U5161 ( .A1(n9142), .A2(n8610), .ZN(n8421) );
  XNOR2_X1 U5162 ( .A(n6411), .B(n6410), .ZN(n6478) );
  OAI21_X1 U5163 ( .B1(n6373), .B2(n5453), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6411) );
  NAND2_X1 U5164 ( .A1(n6408), .A2(n6375), .ZN(n5453) );
  AND2_X2 U5165 ( .A1(n5194), .A2(n5193), .ZN(n6389) );
  INV_X1 U5166 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5193) );
  INV_X1 U5167 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5194) );
  XNOR2_X1 U5168 ( .A(n5663), .B(n5633), .ZN(n5667) );
  INV_X1 U5169 ( .A(n8003), .ZN(n5415) );
  NAND2_X1 U5170 ( .A1(n9786), .A2(n9638), .ZN(n5235) );
  NOR2_X1 U5171 ( .A1(n9944), .A2(n5208), .ZN(n5207) );
  INV_X1 U5172 ( .A(n5209), .ZN(n5208) );
  OR2_X1 U5173 ( .A1(n7958), .A2(n9167), .ZN(n9454) );
  INV_X1 U5174 ( .A(n10279), .ZN(n5621) );
  XNOR2_X1 U5175 ( .A(n10539), .B(n5664), .ZN(n7494) );
  NAND2_X1 U5176 ( .A1(n5499), .A2(n5498), .ZN(n9516) );
  NAND2_X1 U5177 ( .A1(n8225), .A2(n8224), .ZN(n8271) );
  NOR2_X1 U5178 ( .A1(n5099), .A2(n5565), .ZN(n5566) );
  INV_X1 U5179 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5563) );
  XNOR2_X1 U5180 ( .A(n6060), .B(n10188), .ZN(n6061) );
  NAND2_X1 U5181 ( .A1(n6046), .A2(n6045), .ZN(n6062) );
  NAND2_X1 U5182 ( .A1(n5500), .A2(n4945), .ZN(n6046) );
  NAND2_X1 U5183 ( .A1(n5980), .A2(n5979), .ZN(n6001) );
  INV_X1 U5184 ( .A(n5481), .ZN(n5480) );
  OAI21_X1 U5185 ( .B1(n5482), .B2(n5814), .A(n5854), .ZN(n5481) );
  OAI21_X1 U5186 ( .B1(n8553), .B2(n5387), .A(n5386), .ZN(n5385) );
  NAND2_X1 U5187 ( .A1(n8553), .A2(n5390), .ZN(n5386) );
  NOR2_X1 U5188 ( .A1(n5388), .A2(n8559), .ZN(n5387) );
  NAND2_X1 U5189 ( .A1(n5372), .A2(n8706), .ZN(n5371) );
  NAND2_X2 U5190 ( .A1(n7888), .A2(n7887), .ZN(n7989) );
  BUF_X1 U5191 ( .A(n8160), .Z(n8183) );
  AND2_X2 U5192 ( .A1(n8508), .A2(n9153), .ZN(n8160) );
  NAND2_X1 U5193 ( .A1(n6492), .A2(n6491), .ZN(n6685) );
  NOR2_X1 U5194 ( .A1(n7393), .A2(n4934), .ZN(n5316) );
  XNOR2_X1 U5195 ( .A(n8768), .B(n10371), .ZN(n10382) );
  NOR2_X1 U5196 ( .A1(n10381), .A2(n10382), .ZN(n10380) );
  OR2_X1 U5197 ( .A1(n8128), .A2(n5295), .ZN(n5293) );
  AND2_X1 U5198 ( .A1(n8129), .A2(n5296), .ZN(n5295) );
  NAND2_X1 U5199 ( .A1(n8963), .A2(n5554), .ZN(n5296) );
  NAND2_X1 U5200 ( .A1(n5297), .A2(n5554), .ZN(n5294) );
  NAND2_X1 U5201 ( .A1(n8954), .A2(n8955), .ZN(n8232) );
  AOI21_X1 U5202 ( .B1(n4933), .B2(n5269), .A(n4944), .ZN(n5267) );
  INV_X1 U5203 ( .A(n8208), .ZN(n8132) );
  NAND2_X1 U5204 ( .A1(n7674), .A2(n7758), .ZN(n10715) );
  NAND2_X1 U5205 ( .A1(n8249), .A2(n8278), .ZN(n6741) );
  XNOR2_X1 U5206 ( .A(n6524), .B(P2_IR_REG_29__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U5207 ( .A1(n6523), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6524) );
  XNOR2_X1 U5208 ( .A(n6552), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8833) );
  XNOR2_X1 U5209 ( .A(n5742), .B(n5633), .ZN(n5749) );
  NAND3_X1 U5210 ( .A1(n5569), .A2(P1_IR_REG_31__SCAN_IN), .A3(n5568), .ZN(
        n5570) );
  NAND3_X1 U5211 ( .A1(n5041), .A2(n5610), .A3(n6363), .ZN(n6291) );
  AOI21_X1 U5212 ( .B1(n6185), .B2(n5051), .A(n5049), .ZN(n5048) );
  NAND2_X1 U5213 ( .A1(n5050), .A2(n6210), .ZN(n5049) );
  NAND2_X1 U5214 ( .A1(n5051), .A2(n5053), .ZN(n5050) );
  NAND2_X1 U5215 ( .A1(n5620), .A2(n5621), .ZN(n5753) );
  NAND2_X1 U5216 ( .A1(n5257), .A2(n5260), .ZN(n9701) );
  INV_X1 U5217 ( .A(n9698), .ZN(n5260) );
  AOI22_X1 U5218 ( .A1(n9744), .A2(n9641), .B1(n9729), .B2(n9746), .ZN(n9732)
         );
  OAI21_X1 U5219 ( .B1(n9654), .B2(n5134), .A(n5132), .ZN(n9756) );
  INV_X1 U5220 ( .A(n5133), .ZN(n5132) );
  OAI21_X1 U5221 ( .B1(n5135), .B2(n5134), .A(n9760), .ZN(n5133) );
  INV_X1 U5222 ( .A(n9655), .ZN(n5134) );
  INV_X1 U5223 ( .A(n5249), .ZN(n5248) );
  OAI21_X1 U5224 ( .B1(n5252), .B2(n5250), .A(n9475), .ZN(n5249) );
  NAND2_X1 U5225 ( .A1(n5251), .A2(n9466), .ZN(n5250) );
  NAND2_X1 U5226 ( .A1(n7805), .A2(n7803), .ZN(n5534) );
  INV_X1 U5227 ( .A(n5726), .ZN(n9335) );
  NAND2_X1 U5228 ( .A1(n10052), .A2(n10279), .ZN(n5755) );
  AND2_X1 U5229 ( .A1(n5620), .A2(n10279), .ZN(n5671) );
  AND2_X1 U5230 ( .A1(n9701), .A2(n5258), .ZN(n9681) );
  NOR2_X1 U5231 ( .A1(n9679), .A2(n5259), .ZN(n5258) );
  INV_X1 U5232 ( .A(n9661), .ZN(n5259) );
  NAND2_X1 U5233 ( .A1(n7212), .A2(n7211), .ZN(n9852) );
  OR2_X1 U5234 ( .A1(n8285), .A2(n8284), .ZN(n8287) );
  XNOR2_X1 U5235 ( .A(n5606), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6302) );
  OR2_X1 U5236 ( .A1(n5605), .A2(n5604), .ZN(n5606) );
  OAI21_X1 U5237 ( .B1(n6158), .B2(n5464), .A(n5462), .ZN(n6213) );
  NAND2_X1 U5238 ( .A1(n5506), .A2(n5502), .ZN(n6025) );
  NAND2_X1 U5239 ( .A1(n5683), .A2(n5682), .ZN(n5687) );
  AOI21_X1 U5240 ( .B1(n5447), .B2(n4942), .A(n4992), .ZN(n5446) );
  AND2_X1 U5241 ( .A1(n8334), .A2(n8336), .ZN(n5429) );
  OR2_X1 U5242 ( .A1(n8333), .A2(n8344), .ZN(n8334) );
  XNOR2_X1 U5243 ( .A(n5091), .B(n8247), .ZN(n5298) );
  OAI21_X1 U5244 ( .B1(n8845), .B2(n8219), .A(n5016), .ZN(n5091) );
  AND2_X1 U5245 ( .A1(n5213), .A2(n5212), .ZN(n9903) );
  AOI21_X1 U5246 ( .B1(n9673), .B2(n9904), .A(n9826), .ZN(n5212) );
  INV_X1 U5247 ( .A(n9645), .ZN(n5213) );
  INV_X1 U5248 ( .A(n9630), .ZN(n10003) );
  OAI21_X1 U5249 ( .B1(n8397), .B2(n8396), .A(n8395), .ZN(n5196) );
  AOI21_X1 U5250 ( .B1(n8419), .B2(n5167), .A(n5166), .ZN(n5165) );
  OAI21_X1 U5251 ( .B1(n9467), .B2(n9465), .A(n9469), .ZN(n5120) );
  NOR2_X1 U5252 ( .A1(n5119), .A2(n9511), .ZN(n5118) );
  INV_X1 U5253 ( .A(n8474), .ZN(n5176) );
  AND2_X1 U5254 ( .A1(n5177), .A2(n5175), .ZN(n5174) );
  NOR2_X1 U5255 ( .A1(n4957), .A2(n5172), .ZN(n5171) );
  NAND2_X1 U5256 ( .A1(n8462), .A2(n8890), .ZN(n5172) );
  OR2_X1 U5257 ( .A1(n5116), .A2(n9499), .ZN(n5115) );
  INV_X1 U5258 ( .A(n8548), .ZN(n5392) );
  INV_X1 U5259 ( .A(n5098), .ZN(n9366) );
  NOR2_X1 U5260 ( .A1(n9800), .A2(n9813), .ZN(n5209) );
  INV_X1 U5261 ( .A(n5471), .ZN(n5470) );
  OAI21_X1 U5262 ( .B1(n5473), .B2(n5472), .A(n6275), .ZN(n5471) );
  INV_X1 U5263 ( .A(n6255), .ZN(n5472) );
  NAND2_X1 U5264 ( .A1(n5493), .A2(n5491), .ZN(n5490) );
  INV_X1 U5265 ( .A(n6102), .ZN(n5495) );
  INV_X1 U5266 ( .A(n5493), .ZN(n5492) );
  INV_X1 U5267 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U5268 ( .A1(n5374), .A2(n5376), .ZN(n5373) );
  INV_X1 U5269 ( .A(n5378), .ZN(n5374) );
  NOR2_X1 U5270 ( .A1(n8147), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5103) );
  AOI21_X1 U5271 ( .B1(n5346), .B2(n5344), .A(n4979), .ZN(n5343) );
  NAND2_X1 U5272 ( .A1(n8490), .A2(n8492), .ZN(n8493) );
  NAND2_X1 U5273 ( .A1(n6389), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6503) );
  NOR2_X1 U5274 ( .A1(n10398), .A2(n5015), .ZN(n8771) );
  NAND2_X1 U5275 ( .A1(n10389), .A2(n5189), .ZN(n8757) );
  OR2_X1 U5276 ( .A1(n10388), .A2(n10700), .ZN(n5189) );
  NAND2_X1 U5277 ( .A1(n10424), .A2(n5188), .ZN(n8760) );
  OR2_X1 U5278 ( .A1(n10423), .A2(n8759), .ZN(n5188) );
  NOR2_X1 U5279 ( .A1(n10432), .A2(n5095), .ZN(n8773) );
  NOR2_X1 U5280 ( .A1(n10423), .A2(n5096), .ZN(n5095) );
  OR2_X1 U5281 ( .A1(n8922), .A2(n8703), .ZN(n8451) );
  NOR2_X1 U5282 ( .A1(n8096), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6986) );
  NAND2_X1 U5283 ( .A1(n7483), .A2(n8713), .ZN(n8361) );
  OR2_X1 U5284 ( .A1(n9086), .A2(n8879), .ZN(n8471) );
  AND2_X1 U5285 ( .A1(n5276), .A2(n4963), .ZN(n5275) );
  AND2_X1 U5286 ( .A1(n5277), .A2(n4963), .ZN(n5273) );
  AND2_X1 U5287 ( .A1(n8460), .A2(n8461), .ZN(n8458) );
  INV_X1 U5288 ( .A(n8421), .ZN(n5418) );
  NAND2_X1 U5289 ( .A1(n7760), .A2(n8320), .ZN(n5439) );
  OR2_X1 U5290 ( .A1(n7883), .A2(n10672), .ZN(n8392) );
  AOI21_X1 U5291 ( .B1(n5413), .B2(n7901), .A(n5057), .ZN(n5056) );
  INV_X1 U5292 ( .A(n5978), .ZN(n5057) );
  NAND2_X1 U5293 ( .A1(n5056), .A2(n5414), .ZN(n5055) );
  AND2_X1 U5294 ( .A1(n5628), .A2(n5627), .ZN(n5634) );
  NAND2_X1 U5295 ( .A1(n5653), .A2(n10533), .ZN(n5628) );
  AND2_X1 U5296 ( .A1(n5896), .A2(n5402), .ZN(n5401) );
  NAND2_X1 U5297 ( .A1(n5123), .A2(n9510), .ZN(n5122) );
  OR2_X1 U5298 ( .A1(n9349), .A2(n9620), .ZN(n9523) );
  INV_X1 U5299 ( .A(n9640), .ZN(n5225) );
  NOR2_X1 U5300 ( .A1(n9776), .A2(n5136), .ZN(n5135) );
  INV_X1 U5301 ( .A(n9653), .ZN(n5136) );
  NAND2_X1 U5302 ( .A1(n5089), .A2(n4952), .ZN(n5107) );
  OR2_X1 U5303 ( .A1(n9868), .A2(n9968), .ZN(n9475) );
  AND2_X1 U5304 ( .A1(n9872), .A2(n9468), .ZN(n5252) );
  NOR2_X1 U5305 ( .A1(n5204), .A2(n9171), .ZN(n5203) );
  INV_X1 U5306 ( .A(n5205), .ZN(n5204) );
  NAND2_X1 U5307 ( .A1(n9375), .A2(n4959), .ZN(n5529) );
  NOR2_X1 U5308 ( .A1(n7719), .A2(n10680), .ZN(n7787) );
  INV_X1 U5309 ( .A(n7661), .ZN(n5526) );
  OR2_X1 U5310 ( .A1(n7676), .A2(n7698), .ZN(n7708) );
  AOI21_X1 U5311 ( .B1(n7428), .B2(n7427), .A(n9310), .ZN(n9398) );
  NOR2_X2 U5312 ( .A1(n6319), .A2(n5608), .ZN(n9511) );
  OR2_X1 U5313 ( .A1(n9693), .A2(n9911), .ZN(n9661) );
  INV_X1 U5314 ( .A(n9681), .ZN(n5256) );
  INV_X1 U5315 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5612) );
  INV_X1 U5316 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6331) );
  INV_X1 U5317 ( .A(n6212), .ZN(n5460) );
  INV_X1 U5318 ( .A(n6167), .ZN(n5466) );
  NAND2_X1 U5319 ( .A1(n5595), .A2(n5585), .ZN(n5593) );
  NAND2_X1 U5320 ( .A1(n6002), .A2(SI_15_), .ZN(n6024) );
  NOR2_X1 U5321 ( .A1(n5922), .A2(n5517), .ZN(n5516) );
  INV_X1 U5322 ( .A(n5898), .ZN(n5517) );
  INV_X1 U5323 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5560) );
  NOR2_X1 U5324 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5556) );
  NOR2_X1 U5325 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5555) );
  OAI211_X1 U5326 ( .C1(n5487), .C2(P1_DATAO_REG_3__SCAN_IN), .A(n5218), .B(
        n5217), .ZN(n5711) );
  NAND2_X1 U5327 ( .A1(n5129), .A2(n5220), .ZN(n5218) );
  NAND3_X1 U5328 ( .A1(n5301), .A2(n5303), .A3(n5302), .ZN(n5684) );
  NAND2_X1 U5329 ( .A1(n5304), .A2(n5485), .ZN(n5303) );
  NAND2_X1 U5330 ( .A1(n8278), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5104) );
  INV_X1 U5331 ( .A(n5354), .ZN(n5349) );
  NAND2_X1 U5332 ( .A1(n7609), .A2(n7608), .ZN(n7733) );
  INV_X1 U5333 ( .A(n5335), .ZN(n5334) );
  NOR2_X1 U5334 ( .A1(n8663), .A2(n5352), .ZN(n5351) );
  INV_X1 U5335 ( .A(n8524), .ZN(n5352) );
  NAND2_X1 U5336 ( .A1(n8523), .A2(n5354), .ZN(n5353) );
  AND2_X1 U5337 ( .A1(n8249), .A2(n6573), .ZN(n6948) );
  OAI21_X1 U5338 ( .B1(n4936), .B2(n5368), .A(n8566), .ZN(n5367) );
  NAND2_X1 U5339 ( .A1(n6428), .A2(n6382), .ZN(n6494) );
  AND2_X1 U5340 ( .A1(n6381), .A2(n6380), .ZN(n6382) );
  NAND2_X1 U5341 ( .A1(n6685), .A2(n6684), .ZN(n5323) );
  NOR2_X1 U5342 ( .A1(n5321), .A2(n6934), .ZN(n5320) );
  INV_X1 U5343 ( .A(n6684), .ZN(n5321) );
  OAI211_X1 U5344 ( .C1(n7182), .C2(n5313), .A(n5312), .B(n5310), .ZN(n7410)
         );
  AOI21_X1 U5345 ( .B1(n5314), .B2(n4934), .A(n5311), .ZN(n5310) );
  OAI21_X1 U5346 ( .B1(n5313), .B2(n7183), .A(P2_REG2_REG_7__SCAN_IN), .ZN(
        n5311) );
  OR2_X1 U5347 ( .A1(n7541), .A2(n8742), .ZN(n5308) );
  AND2_X1 U5348 ( .A1(n7541), .A2(n8742), .ZN(n8730) );
  NAND2_X1 U5349 ( .A1(n5308), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5306) );
  OR2_X1 U5350 ( .A1(n6581), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n6582) );
  NOR2_X1 U5351 ( .A1(n10380), .A2(n8769), .ZN(n10400) );
  NAND2_X1 U5352 ( .A1(n10390), .A2(n10391), .ZN(n10389) );
  XNOR2_X1 U5353 ( .A(n8771), .B(n10406), .ZN(n10417) );
  NOR2_X1 U5354 ( .A1(n10417), .A2(n10416), .ZN(n10415) );
  XNOR2_X1 U5355 ( .A(n8757), .B(n10406), .ZN(n10408) );
  NAND2_X1 U5356 ( .A1(n10425), .A2(n10426), .ZN(n10424) );
  XNOR2_X1 U5357 ( .A(n8760), .B(n10440), .ZN(n10442) );
  NAND2_X1 U5358 ( .A1(n10477), .A2(n8763), .ZN(n10495) );
  NAND2_X1 U5359 ( .A1(n7047), .A2(n7046), .ZN(n8194) );
  INV_X1 U5360 ( .A(n8192), .ZN(n7047) );
  NOR2_X1 U5361 ( .A1(n5285), .A2(n8309), .ZN(n5284) );
  NOR2_X1 U5362 ( .A1(n4954), .A2(n8934), .ZN(n5285) );
  AOI21_X1 U5363 ( .B1(n5284), .B2(n4954), .A(n5283), .ZN(n5282) );
  INV_X1 U5364 ( .A(n8451), .ZN(n5283) );
  NAND2_X1 U5365 ( .A1(n5039), .A2(n8400), .ZN(n8035) );
  AND4_X1 U5366 ( .A1(n7593), .A2(n7592), .A3(n7591), .A4(n7590), .ZN(n7893)
         );
  NAND2_X1 U5367 ( .A1(n7272), .A2(n8365), .ZN(n7250) );
  AND2_X1 U5368 ( .A1(n8369), .A2(n8370), .ZN(n8312) );
  NAND2_X1 U5369 ( .A1(n7250), .A2(n8312), .ZN(n7461) );
  AND2_X1 U5370 ( .A1(n8350), .A2(n8357), .ZN(n8314) );
  INV_X1 U5371 ( .A(n8842), .ZN(n8844) );
  NAND2_X1 U5372 ( .A1(n8290), .A2(n8289), .ZN(n8303) );
  OR2_X1 U5373 ( .A1(n8865), .A2(n8240), .ZN(n5450) );
  INV_X1 U5374 ( .A(n8297), .ZN(n5449) );
  NAND2_X1 U5375 ( .A1(n5035), .A2(n8464), .ZN(n8875) );
  NAND2_X1 U5376 ( .A1(n5437), .A2(n5435), .ZN(n5035) );
  NOR2_X1 U5377 ( .A1(n8459), .A2(n5436), .ZN(n5435) );
  INV_X1 U5378 ( .A(n8461), .ZN(n5436) );
  AND3_X1 U5379 ( .A1(n8186), .A2(n8185), .A3(n8184), .ZN(n8898) );
  OR2_X1 U5380 ( .A1(n5281), .A2(n8308), .ZN(n5277) );
  INV_X1 U5381 ( .A(n5282), .ZN(n5281) );
  OR2_X1 U5382 ( .A1(n5279), .A2(n8308), .ZN(n5276) );
  AOI21_X1 U5383 ( .B1(n5280), .B2(n5282), .A(n4988), .ZN(n5279) );
  INV_X1 U5384 ( .A(n5284), .ZN(n5280) );
  OR2_X1 U5385 ( .A1(n8947), .A2(n8957), .ZN(n8141) );
  AOI21_X1 U5386 ( .B1(n5293), .B2(n5294), .A(n4985), .ZN(n5292) );
  OR2_X1 U5387 ( .A1(n6948), .A2(n8491), .ZN(n10566) );
  INV_X1 U5388 ( .A(n8458), .ZN(n8895) );
  OR2_X1 U5389 ( .A1(n5430), .A2(n8921), .ZN(n5030) );
  NAND2_X1 U5390 ( .A1(n5032), .A2(n8948), .ZN(n5031) );
  AND2_X1 U5391 ( .A1(n8434), .A2(n8429), .ZN(n8955) );
  NAND2_X1 U5392 ( .A1(n8966), .A2(n8965), .ZN(n8964) );
  INV_X1 U5393 ( .A(n8976), .ZN(n8973) );
  NAND2_X1 U5394 ( .A1(n8231), .A2(n8421), .ZN(n8974) );
  OR2_X1 U5395 ( .A1(n8326), .A2(n5269), .ZN(n5268) );
  NAND2_X1 U5396 ( .A1(n8105), .A2(n8418), .ZN(n8992) );
  NAND2_X1 U5397 ( .A1(n6800), .A2(n6799), .ZN(n8989) );
  INV_X1 U5398 ( .A(n10566), .ZN(n8995) );
  NAND2_X1 U5399 ( .A1(n8035), .A2(n5443), .ZN(n8086) );
  NOR2_X1 U5400 ( .A1(n8081), .A2(n5444), .ZN(n5443) );
  INV_X1 U5401 ( .A(n8034), .ZN(n5444) );
  NAND2_X1 U5402 ( .A1(n8086), .A2(n5441), .ZN(n8230) );
  NOR2_X1 U5403 ( .A1(n8326), .A2(n5442), .ZN(n5441) );
  INV_X1 U5404 ( .A(n8407), .ZN(n5442) );
  INV_X1 U5405 ( .A(n8989), .ZN(n10562) );
  OR2_X1 U5406 ( .A1(n8491), .A2(n6801), .ZN(n6840) );
  XNOR2_X1 U5407 ( .A(n5197), .B(n6409), .ZN(n6482) );
  OAI21_X1 U5408 ( .B1(n6373), .B2(n4990), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5197) );
  INV_X1 U5409 ( .A(n6478), .ZN(n6572) );
  INV_X1 U5410 ( .A(n5361), .ZN(n5357) );
  NAND2_X1 U5411 ( .A1(n6413), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U5412 ( .A1(n6549), .A2(n6548), .ZN(n6551) );
  INV_X1 U5413 ( .A(n6389), .ZN(n5309) );
  NAND2_X1 U5414 ( .A1(n5412), .A2(n5411), .ZN(n9162) );
  AOI21_X1 U5415 ( .B1(n7901), .B2(n5413), .A(n4993), .ZN(n5411) );
  OAI21_X1 U5416 ( .B1(n7696), .B2(n7692), .A(n7693), .ZN(n5403) );
  INV_X1 U5417 ( .A(n5403), .ZN(n5400) );
  INV_X1 U5418 ( .A(n9183), .ZN(n5061) );
  NAND2_X1 U5419 ( .A1(n9254), .A2(n6080), .ZN(n5070) );
  NAND2_X1 U5420 ( .A1(n5062), .A2(n9252), .ZN(n5069) );
  OR2_X1 U5421 ( .A1(n9254), .A2(n6080), .ZN(n5062) );
  AND2_X1 U5422 ( .A1(n6032), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U5423 ( .A1(n6050), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6090) );
  AND2_X1 U5424 ( .A1(n5004), .A2(n4937), .ZN(n5053) );
  NOR2_X1 U5425 ( .A1(n5052), .A2(n5405), .ZN(n5051) );
  NOR2_X1 U5426 ( .A1(n4937), .A2(n6184), .ZN(n5052) );
  XNOR2_X1 U5427 ( .A(n5720), .B(n5633), .ZN(n5744) );
  AND2_X1 U5428 ( .A1(n7089), .A2(n7090), .ZN(n5100) );
  NAND2_X1 U5429 ( .A1(n5067), .A2(n5058), .ZN(n9231) );
  AOI21_X1 U5430 ( .B1(n9254), .B2(n5065), .A(n5063), .ZN(n5067) );
  AOI21_X1 U5431 ( .B1(n9254), .B2(n5060), .A(n5059), .ZN(n5058) );
  NOR2_X1 U5432 ( .A1(n9233), .A2(n5066), .ZN(n5065) );
  NAND2_X1 U5433 ( .A1(n5085), .A2(n5084), .ZN(n5416) );
  NOR2_X1 U5434 ( .A1(n5401), .A2(n5399), .ZN(n5398) );
  INV_X1 U5435 ( .A(n7693), .ZN(n5399) );
  AND2_X1 U5436 ( .A1(n5396), .A2(n5395), .ZN(n5394) );
  OR2_X1 U5437 ( .A1(n5896), .A2(n5402), .ZN(n5395) );
  OR2_X1 U5438 ( .A1(n5401), .A2(n5397), .ZN(n5396) );
  NAND2_X1 U5439 ( .A1(n7692), .A2(n7693), .ZN(n5397) );
  NAND2_X1 U5440 ( .A1(n4932), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5656) );
  OR2_X1 U5441 ( .A1(n5753), .A2(n10534), .ZN(n5622) );
  NAND2_X1 U5442 ( .A1(n5106), .A2(n5012), .ZN(n9715) );
  INV_X1 U5443 ( .A(n9702), .ZN(n9730) );
  NAND2_X1 U5444 ( .A1(n9756), .A2(n9656), .ZN(n9752) );
  NAND2_X1 U5445 ( .A1(n5232), .A2(n5235), .ZN(n5228) );
  NAND2_X1 U5446 ( .A1(n4997), .A2(n5235), .ZN(n5227) );
  NAND2_X1 U5447 ( .A1(n5232), .A2(n5231), .ZN(n5230) );
  INV_X1 U5448 ( .A(n5233), .ZN(n5231) );
  AND2_X1 U5449 ( .A1(n9497), .A2(n9656), .ZN(n9760) );
  NAND2_X1 U5450 ( .A1(n9654), .A2(n5135), .ZN(n9773) );
  OR2_X1 U5451 ( .A1(n9800), .A2(n9778), .ZN(n9653) );
  NOR2_X1 U5452 ( .A1(n9793), .A2(n5234), .ZN(n5233) );
  NOR2_X1 U5453 ( .A1(n4935), .A2(n9803), .ZN(n5234) );
  AOI21_X1 U5454 ( .B1(n5148), .B2(n9473), .A(n9803), .ZN(n5146) );
  NAND2_X1 U5455 ( .A1(n9835), .A2(n5148), .ZN(n5147) );
  INV_X1 U5456 ( .A(n5107), .ZN(n9804) );
  AND2_X1 U5457 ( .A1(n9485), .A2(n9484), .ZN(n9823) );
  NAND2_X1 U5458 ( .A1(n9342), .A2(n5252), .ZN(n9874) );
  OR2_X1 U5459 ( .A1(n9632), .A2(n9879), .ZN(n9468) );
  AND2_X1 U5460 ( .A1(n9632), .A2(n9631), .ZN(n5237) );
  AND2_X1 U5461 ( .A1(n7917), .A2(n5533), .ZN(n5532) );
  NAND2_X1 U5462 ( .A1(n7804), .A2(n7803), .ZN(n5533) );
  NAND2_X1 U5463 ( .A1(n9454), .A2(n9456), .ZN(n9375) );
  OAI21_X1 U5464 ( .B1(n7235), .B2(n5726), .A(n5242), .ZN(n7456) );
  NOR2_X1 U5465 ( .A1(n4967), .A2(n5243), .ZN(n5242) );
  NOR2_X1 U5466 ( .A1(n5086), .A2(n6784), .ZN(n5243) );
  NAND2_X1 U5467 ( .A1(n10052), .A2(n5621), .ZN(n5751) );
  NAND2_X1 U5468 ( .A1(n4932), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5673) );
  OR2_X1 U5469 ( .A1(n9522), .A2(n10347), .ZN(n9880) );
  NAND2_X1 U5470 ( .A1(n7494), .A2(n7493), .ZN(n7492) );
  NOR2_X1 U5471 ( .A1(n6474), .A2(n5611), .ZN(n9363) );
  AND4_X1 U5472 ( .A1(n6290), .A2(n6289), .A3(n6288), .A4(n6287), .ZN(n9902)
         );
  NAND2_X1 U5473 ( .A1(n9337), .A2(n9336), .ZN(n9621) );
  NAND2_X1 U5474 ( .A1(n5963), .A2(n5962), .ZN(n7958) );
  NAND2_X1 U5475 ( .A1(n5905), .A2(n5904), .ZN(n7802) );
  INV_X1 U5476 ( .A(n10729), .ZN(n10705) );
  NAND3_X1 U5477 ( .A1(n6302), .A2(n6300), .A3(n6301), .ZN(n10042) );
  XNOR2_X1 U5478 ( .A(n5615), .B(n10046), .ZN(n5620) );
  NAND2_X1 U5479 ( .A1(n5265), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5615) );
  OR2_X1 U5480 ( .A1(n8271), .A2(n8270), .ZN(n8272) );
  INV_X1 U5481 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U5482 ( .A1(n5469), .A2(n6255), .ZN(n6276) );
  NAND2_X1 U5483 ( .A1(n6233), .A2(n5473), .ZN(n5469) );
  OAI21_X1 U5484 ( .B1(n5593), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5586) );
  AND2_X1 U5485 ( .A1(n6167), .A2(n6156), .ZN(n6157) );
  NAND2_X1 U5486 ( .A1(n6082), .A2(n6081), .ZN(n6103) );
  NAND2_X1 U5487 ( .A1(n5494), .A2(n5493), .ZN(n6082) );
  OAI21_X1 U5488 ( .B1(n5078), .B2(n5581), .A(n5077), .ZN(n5076) );
  NAND2_X1 U5489 ( .A1(n5582), .A2(n5589), .ZN(n5078) );
  NAND2_X1 U5490 ( .A1(n5604), .A2(n5589), .ZN(n5077) );
  NAND2_X1 U5491 ( .A1(n5508), .A2(n5507), .ZN(n5506) );
  NOR2_X1 U5492 ( .A1(n5925), .A2(n5515), .ZN(n5512) );
  INV_X1 U5493 ( .A(n5477), .ZN(n5476) );
  XNOR2_X1 U5494 ( .A(n5131), .B(n5874), .ZN(n7580) );
  OAI21_X1 U5495 ( .B1(n5815), .B2(n5482), .A(n5480), .ZN(n5131) );
  NAND2_X1 U5496 ( .A1(n5769), .A2(n4962), .ZN(n5788) );
  OAI21_X1 U5497 ( .B1(n5684), .B2(SI_2_), .A(n5707), .ZN(n5685) );
  NOR2_X1 U5498 ( .A1(n5643), .A2(n10105), .ZN(n5644) );
  INV_X1 U5499 ( .A(n7478), .ZN(n10638) );
  INV_X1 U5500 ( .A(n8967), .ZN(n8945) );
  NOR2_X1 U5501 ( .A1(n5383), .A2(n8683), .ZN(n5381) );
  AND2_X1 U5502 ( .A1(n5385), .A2(n4966), .ZN(n5383) );
  NAND2_X1 U5503 ( .A1(n5385), .A2(n5389), .ZN(n5384) );
  NAND2_X1 U5504 ( .A1(n8553), .A2(n8559), .ZN(n5389) );
  NAND2_X1 U5505 ( .A1(n8547), .A2(n5007), .ZN(n8549) );
  INV_X1 U5506 ( .A(n8704), .ZN(n8944) );
  XNOR2_X1 U5507 ( .A(n8533), .B(n8703), .ZN(n8590) );
  NAND2_X1 U5508 ( .A1(n8073), .A2(n8072), .ZN(n8511) );
  AND4_X1 U5509 ( .A1(n8101), .A2(n8100), .A3(n8099), .A4(n8098), .ZN(n8619)
         );
  INV_X1 U5510 ( .A(n8679), .ZN(n8689) );
  NAND2_X1 U5511 ( .A1(n8146), .A2(n8145), .ZN(n8642) );
  INV_X1 U5512 ( .A(n8993), .ZN(n8692) );
  NAND2_X1 U5513 ( .A1(n8038), .A2(n8037), .ZN(n8652) );
  AND3_X1 U5514 ( .A1(n6993), .A2(n6992), .A3(n6991), .ZN(n8907) );
  AND4_X1 U5515 ( .A1(n8118), .A2(n8117), .A3(n8116), .A4(n8115), .ZN(n8668)
         );
  NAND2_X1 U5516 ( .A1(n6578), .A2(n10570), .ZN(n8681) );
  INV_X1 U5517 ( .A(n5426), .ZN(n5425) );
  AND2_X1 U5518 ( .A1(n5184), .A2(n8506), .ZN(n5423) );
  OAI211_X1 U5519 ( .C1(n5426), .C2(n4947), .A(n5185), .B(n5428), .ZN(n5184)
         );
  NAND2_X1 U5520 ( .A1(n7153), .A2(n7152), .ZN(n8554) );
  OAI211_X1 U5521 ( .C1(n8215), .C2(n9105), .A(n8173), .B(n8172), .ZN(n8702)
         );
  NAND4_X1 U5522 ( .A1(n6603), .A2(n6602), .A3(n6601), .A4(n6600), .ZN(n8716)
         );
  XNOR2_X1 U5523 ( .A(n10495), .B(n10494), .ZN(n5201) );
  NAND2_X1 U5524 ( .A1(n5200), .A2(n5199), .ZN(n5198) );
  INV_X1 U5525 ( .A(n10497), .ZN(n5199) );
  NAND2_X1 U5526 ( .A1(n10498), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n5200) );
  NOR2_X1 U5527 ( .A1(n8832), .A2(n5329), .ZN(n5328) );
  NAND2_X1 U5528 ( .A1(n8784), .A2(n5330), .ZN(n5329) );
  OAI211_X1 U5529 ( .C1(n8778), .C2(n8777), .A(n5093), .B(n5092), .ZN(n8781)
         );
  OR2_X1 U5530 ( .A1(n8779), .A2(n10510), .ZN(n5092) );
  NAND2_X1 U5531 ( .A1(n10504), .A2(n5094), .ZN(n5093) );
  NAND2_X1 U5532 ( .A1(n8176), .A2(n8175), .ZN(n8902) );
  NAND2_X1 U5533 ( .A1(n7929), .A2(n7928), .ZN(n8401) );
  AOI21_X1 U5534 ( .B1(n10050), .B2(n8288), .A(n8283), .ZN(n9067) );
  AND2_X1 U5535 ( .A1(n9011), .A2(n5553), .ZN(n9012) );
  OR2_X1 U5536 ( .A1(n9010), .A2(n10715), .ZN(n5553) );
  NAND2_X1 U5537 ( .A1(n8210), .A2(n8209), .ZN(n9074) );
  OR2_X1 U5538 ( .A1(n8208), .A2(n8207), .ZN(n8209) );
  NAND2_X1 U5539 ( .A1(n8112), .A2(n8111), .ZN(n9129) );
  NAND2_X1 U5540 ( .A1(n8104), .A2(n8103), .ZN(n9135) );
  NAND2_X1 U5541 ( .A1(n8108), .A2(n8107), .ZN(n9142) );
  NAND2_X1 U5542 ( .A1(n5607), .A2(n6302), .ZN(n6363) );
  XNOR2_X1 U5543 ( .A(n6317), .B(n6316), .ZN(n7814) );
  NAND2_X1 U5544 ( .A1(n6315), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6317) );
  AND2_X1 U5545 ( .A1(n5551), .A2(n9259), .ZN(n5043) );
  NAND2_X1 U5546 ( .A1(n6281), .A2(n6280), .ZN(n9630) );
  NAND2_X2 U5547 ( .A1(n5652), .A2(n5651), .ZN(n7496) );
  OR2_X1 U5548 ( .A1(n5735), .A2(n6399), .ZN(n5652) );
  NAND2_X1 U5549 ( .A1(n6031), .A2(n6030), .ZN(n9982) );
  NAND2_X1 U5550 ( .A1(n6192), .A2(n6191), .ZN(n9933) );
  NAND2_X1 U5551 ( .A1(n6161), .A2(n6160), .ZN(n9944) );
  OR2_X1 U5552 ( .A1(n6335), .A2(n10347), .ZN(n9276) );
  NAND2_X1 U5553 ( .A1(n9196), .A2(n6252), .ZN(n9260) );
  AND2_X1 U5554 ( .A1(n6442), .A2(n6637), .ZN(n10350) );
  NAND2_X1 U5555 ( .A1(n9298), .A2(n9297), .ZN(n9628) );
  INV_X1 U5556 ( .A(n9907), .ZN(n5155) );
  NAND2_X1 U5557 ( .A1(n6236), .A2(n6235), .ZN(n9724) );
  INV_X1 U5558 ( .A(n9635), .ZN(n9968) );
  NAND2_X1 U5559 ( .A1(n6083), .A2(n6630), .ZN(n5518) );
  NAND2_X1 U5560 ( .A1(n10525), .A2(n7350), .ZN(n9888) );
  OAI211_X1 U5561 ( .C1(n9670), .C2(n5497), .A(n5543), .B(n5537), .ZN(n9907)
         );
  NAND2_X1 U5562 ( .A1(n9664), .A2(n5006), .ZN(n5543) );
  NAND2_X1 U5563 ( .A1(n9670), .A2(n5542), .ZN(n5537) );
  NOR2_X1 U5564 ( .A1(n9664), .A2(n5006), .ZN(n5542) );
  INV_X1 U5565 ( .A(n5541), .ZN(n5540) );
  OAI21_X1 U5566 ( .B1(n9905), .B2(n10737), .A(n5022), .ZN(n5541) );
  INV_X1 U5567 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5545) );
  AND2_X1 U5568 ( .A1(n9667), .A2(n9666), .ZN(n5157) );
  AND2_X1 U5569 ( .A1(n5241), .A2(n5240), .ZN(n10001) );
  AND2_X1 U5570 ( .A1(n4998), .A2(n9910), .ZN(n5240) );
  OAI211_X1 U5571 ( .C1(n8399), .C2(n8491), .A(n8400), .B(n5195), .ZN(n8406)
         );
  NAND2_X1 U5572 ( .A1(n8973), .A2(n8422), .ZN(n5166) );
  NAND2_X1 U5573 ( .A1(n5163), .A2(n8425), .ZN(n8432) );
  NAND2_X1 U5574 ( .A1(n5163), .A2(n4969), .ZN(n8431) );
  INV_X1 U5575 ( .A(n8426), .ZN(n5164) );
  AND2_X1 U5576 ( .A1(n8874), .A2(n8466), .ZN(n5177) );
  NAND3_X1 U5577 ( .A1(n8462), .A2(n8890), .A3(n8895), .ZN(n5175) );
  OAI21_X1 U5578 ( .B1(n9472), .B2(n9515), .A(n5117), .ZN(n9481) );
  AOI21_X1 U5579 ( .B1(n5120), .B2(n5118), .A(n9636), .ZN(n5117) );
  NAND2_X1 U5580 ( .A1(n5173), .A2(n8856), .ZN(n5170) );
  INV_X1 U5581 ( .A(n6061), .ZN(n5491) );
  INV_X1 U5582 ( .A(n5346), .ZN(n5345) );
  INV_X1 U5583 ( .A(n7608), .ZN(n5344) );
  INV_X1 U5584 ( .A(n8338), .ZN(n8310) );
  NAND2_X1 U5585 ( .A1(n10572), .A2(n8716), .ZN(n8351) );
  OR2_X1 U5586 ( .A1(n9505), .A2(n5126), .ZN(n5125) );
  OAI21_X1 U5587 ( .B1(n9500), .B2(n5115), .A(n5113), .ZN(n9506) );
  NAND2_X1 U5588 ( .A1(n5126), .A2(n9511), .ZN(n5124) );
  AOI21_X1 U5589 ( .B1(n9751), .B2(n9657), .A(n5145), .ZN(n5144) );
  INV_X1 U5590 ( .A(SI_20_), .ZN(n10186) );
  INV_X1 U5591 ( .A(SI_17_), .ZN(n10188) );
  NAND2_X1 U5592 ( .A1(n6000), .A2(n5502), .ZN(n5501) );
  INV_X1 U5593 ( .A(n6041), .ZN(n5503) );
  INV_X1 U5594 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5881) );
  INV_X1 U5595 ( .A(SI_9_), .ZN(n10203) );
  INV_X1 U5596 ( .A(SI_8_), .ZN(n10210) );
  NAND2_X1 U5597 ( .A1(n5129), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5128) );
  NOR2_X1 U5598 ( .A1(n5305), .A2(n5486), .ZN(n5304) );
  NAND2_X1 U5599 ( .A1(n7042), .A2(n5572), .ZN(n5484) );
  INV_X1 U5600 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5572) );
  AND2_X1 U5601 ( .A1(n5391), .A2(n5393), .ZN(n5390) );
  NAND2_X1 U5602 ( .A1(n8551), .A2(n8554), .ZN(n5393) );
  NAND2_X1 U5603 ( .A1(n8559), .A2(n5392), .ZN(n5391) );
  NAND2_X1 U5604 ( .A1(n5190), .A2(n8489), .ZN(n8499) );
  NAND2_X1 U5605 ( .A1(n8495), .A2(n8487), .ZN(n5190) );
  NAND2_X1 U5606 ( .A1(n6389), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U5607 ( .A1(n5309), .A2(n4970), .ZN(n6501) );
  OR2_X1 U5608 ( .A1(n8745), .A2(n8722), .ZN(n8765) );
  OR2_X1 U5609 ( .A1(n7536), .A2(n5186), .ZN(n8741) );
  NOR2_X1 U5610 ( .A1(n7571), .A2(n10658), .ZN(n5186) );
  NAND2_X1 U5611 ( .A1(n10458), .A2(n5187), .ZN(n8762) );
  OR2_X1 U5612 ( .A1(n10457), .A2(n9057), .ZN(n5187) );
  NAND2_X1 U5613 ( .A1(n8247), .A2(n4956), .ZN(n8244) );
  INV_X1 U5614 ( .A(n5103), .ZN(n8157) );
  INV_X1 U5615 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10239) );
  NOR2_X1 U5616 ( .A1(n7767), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5102) );
  NAND2_X1 U5617 ( .A1(n10614), .A2(n8712), .ZN(n8369) );
  INV_X1 U5618 ( .A(n10572), .ZN(n7072) );
  NAND2_X1 U5619 ( .A1(n8342), .A2(n8346), .ZN(n6946) );
  OR2_X1 U5620 ( .A1(n8491), .A2(n6563), .ZN(n6813) );
  NOR2_X1 U5621 ( .A1(n5433), .A2(n8921), .ZN(n5032) );
  OR2_X1 U5622 ( .A1(n6547), .A2(n6546), .ZN(n6806) );
  NAND2_X1 U5623 ( .A1(n6371), .A2(n5362), .ZN(n5361) );
  INV_X1 U5624 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5362) );
  NAND4_X1 U5625 ( .A1(n7282), .A2(n7098), .A3(n6970), .A4(n7285), .ZN(n6370)
         );
  INV_X1 U5626 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5363) );
  INV_X1 U5627 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7098) );
  INV_X1 U5628 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6454) );
  INV_X1 U5629 ( .A(n9252), .ZN(n5066) );
  NOR2_X1 U5630 ( .A1(n9233), .A2(n5061), .ZN(n5059) );
  NOR2_X1 U5631 ( .A1(n9233), .A2(n9251), .ZN(n5060) );
  NAND2_X1 U5632 ( .A1(n9252), .A2(n6080), .ZN(n5064) );
  INV_X1 U5633 ( .A(n7821), .ZN(n5402) );
  NOR2_X1 U5634 ( .A1(n9672), .A2(n9630), .ZN(n9644) );
  NAND2_X1 U5635 ( .A1(n9691), .A2(n9615), .ZN(n9672) );
  NOR2_X1 U5636 ( .A1(n9720), .A2(n9724), .ZN(n9691) );
  AOI21_X1 U5637 ( .B1(n5144), .B2(n9391), .A(n5141), .ZN(n5140) );
  INV_X1 U5638 ( .A(n9659), .ZN(n5141) );
  OR2_X1 U5639 ( .A1(n9752), .A2(n5142), .ZN(n5139) );
  INV_X1 U5640 ( .A(n5144), .ZN(n5142) );
  NAND2_X1 U5641 ( .A1(n9724), .A2(n9730), .ZN(n9660) );
  OR2_X1 U5642 ( .A1(n9724), .A2(n9730), .ZN(n9504) );
  NAND2_X1 U5643 ( .A1(n9745), .A2(n10014), .ZN(n9720) );
  AOI21_X1 U5644 ( .B1(n5151), .B2(n5150), .A(n5149), .ZN(n5148) );
  INV_X1 U5645 ( .A(n9484), .ZN(n5149) );
  OR2_X1 U5646 ( .A1(n9171), .A2(n9987), .ZN(n9460) );
  NOR2_X1 U5647 ( .A1(n6012), .A2(n6011), .ZN(n6032) );
  OR2_X1 U5648 ( .A1(n5985), .A2(n5984), .ZN(n6012) );
  AND2_X1 U5649 ( .A1(n9460), .A2(n9300), .ZN(n9451) );
  NOR2_X1 U5650 ( .A1(n10706), .A2(n7958), .ZN(n5205) );
  OR2_X1 U5651 ( .A1(n10706), .A2(n8008), .ZN(n9453) );
  OR2_X1 U5652 ( .A1(n7712), .A2(n9367), .ZN(n7713) );
  NOR2_X1 U5653 ( .A1(n7210), .A2(n5254), .ZN(n5253) );
  INV_X1 U5654 ( .A(n7207), .ZN(n5254) );
  AND2_X1 U5655 ( .A1(n7562), .A2(n7659), .ZN(n7668) );
  XNOR2_X1 U5656 ( .A(n8271), .B(n8269), .ZN(n8268) );
  NAND2_X1 U5657 ( .A1(n5468), .A2(n5467), .ZN(n8221) );
  AOI21_X1 U5658 ( .B1(n5470), .B2(n5472), .A(n5026), .ZN(n5467) );
  NOR2_X1 U5659 ( .A1(n6256), .A2(n5474), .ZN(n5473) );
  INV_X1 U5660 ( .A(n6232), .ZN(n5474) );
  AND2_X1 U5661 ( .A1(n5010), .A2(n6067), .ZN(n5493) );
  INV_X1 U5662 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5900) );
  INV_X1 U5663 ( .A(n5874), .ZN(n5479) );
  INV_X1 U5664 ( .A(SI_10_), .ZN(n10199) );
  NAND2_X1 U5665 ( .A1(n5483), .A2(n5830), .ZN(n5482) );
  INV_X1 U5666 ( .A(n5855), .ZN(n5483) );
  INV_X1 U5667 ( .A(n5711), .ZN(n5709) );
  INV_X1 U5668 ( .A(n5040), .ZN(n5129) );
  INV_X1 U5669 ( .A(n5390), .ZN(n5388) );
  NAND2_X1 U5670 ( .A1(n7369), .A2(n7368), .ZN(n7607) );
  NAND2_X1 U5671 ( .A1(n6978), .A2(n6977), .ZN(n7371) );
  INV_X1 U5672 ( .A(n7241), .ZN(n6978) );
  XNOR2_X1 U5673 ( .A(n6861), .B(n6997), .ZN(n6597) );
  INV_X1 U5674 ( .A(n5376), .ZN(n5375) );
  OAI21_X1 U5675 ( .B1(n7131), .B2(n7130), .A(n7129), .ZN(n7310) );
  INV_X1 U5676 ( .A(n8539), .ZN(n8623) );
  NAND2_X1 U5677 ( .A1(n8657), .A2(n8538), .ZN(n8576) );
  NOR2_X1 U5678 ( .A1(n7734), .A2(n5347), .ZN(n5346) );
  INV_X1 U5679 ( .A(n7732), .ZN(n5347) );
  OR2_X1 U5680 ( .A1(n7371), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7574) );
  NAND2_X1 U5681 ( .A1(n6980), .A2(n6979), .ZN(n7588) );
  INV_X1 U5682 ( .A(n7574), .ZN(n6980) );
  NAND2_X1 U5683 ( .A1(n8530), .A2(n8529), .ZN(n8635) );
  INV_X1 U5684 ( .A(n8638), .ZN(n8529) );
  NOR2_X1 U5685 ( .A1(n8655), .A2(n5379), .ZN(n5378) );
  INV_X1 U5686 ( .A(n8534), .ZN(n5379) );
  NAND2_X1 U5687 ( .A1(n5103), .A2(n6988), .ZN(n8169) );
  NAND2_X1 U5688 ( .A1(n5333), .A2(n7991), .ZN(n8069) );
  INV_X1 U5689 ( .A(n5102), .ZN(n7830) );
  NOR2_X1 U5690 ( .A1(n7312), .A2(n7313), .ZN(n7363) );
  NOR2_X1 U5691 ( .A1(n5448), .A2(n4986), .ZN(n5447) );
  NOR2_X1 U5692 ( .A1(n5449), .A2(n8300), .ZN(n5448) );
  NAND2_X1 U5693 ( .A1(n8303), .A2(n8301), .ZN(n8490) );
  NAND2_X1 U5694 ( .A1(n5426), .A2(n8833), .ZN(n5185) );
  AND4_X1 U5695 ( .A1(n6570), .A2(n6569), .A3(n6568), .A4(n6567), .ZN(n6943)
         );
  OAI21_X1 U5696 ( .B1(n7173), .B2(n5180), .A(n5178), .ZN(n5182) );
  AOI21_X1 U5697 ( .B1(n5183), .B2(n5179), .A(n7175), .ZN(n5178) );
  INV_X1 U5698 ( .A(n5183), .ZN(n5180) );
  AND2_X1 U5699 ( .A1(n5182), .A2(n5181), .ZN(n7391) );
  NAND2_X1 U5700 ( .A1(n7326), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5181) );
  XNOR2_X1 U5701 ( .A(n8741), .B(n7581), .ZN(n7538) );
  INV_X1 U5702 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10242) );
  NAND2_X1 U5703 ( .A1(n10372), .A2(n8756), .ZN(n10390) );
  NOR2_X1 U5704 ( .A1(n10415), .A2(n8772), .ZN(n10434) );
  NAND2_X1 U5705 ( .A1(n10407), .A2(n8758), .ZN(n10425) );
  NAND2_X1 U5706 ( .A1(n10441), .A2(n8761), .ZN(n10459) );
  NAND2_X1 U5707 ( .A1(n10459), .A2(n10460), .ZN(n10458) );
  NOR2_X1 U5708 ( .A1(n8774), .A2(n10449), .ZN(n10469) );
  NOR2_X1 U5709 ( .A1(n10469), .A2(n10468), .ZN(n10467) );
  XNOR2_X1 U5710 ( .A(n8762), .B(n10475), .ZN(n10478) );
  OAI21_X1 U5711 ( .B1(n5324), .B2(n8819), .A(n8778), .ZN(n10487) );
  INV_X1 U5712 ( .A(n8778), .ZN(n10505) );
  NAND2_X1 U5713 ( .A1(n10476), .A2(n8833), .ZN(n5330) );
  INV_X1 U5714 ( .A(n10507), .ZN(n5094) );
  OR2_X1 U5715 ( .A1(n8211), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8260) );
  AND2_X1 U5716 ( .A1(n7144), .A2(n10265), .ZN(n7146) );
  OR2_X1 U5717 ( .A1(n8468), .A2(n8467), .ZN(n8876) );
  AOI21_X1 U5718 ( .B1(n5432), .B2(n5434), .A(n4981), .ZN(n5430) );
  NAND2_X1 U5719 ( .A1(n6987), .A2(n10239), .ZN(n8147) );
  INV_X1 U5720 ( .A(n8135), .ZN(n6987) );
  INV_X1 U5721 ( .A(n8055), .ZN(n6984) );
  INV_X1 U5722 ( .A(n6986), .ZN(n8113) );
  OR2_X1 U5723 ( .A1(n8042), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8055) );
  NAND2_X1 U5724 ( .A1(n5102), .A2(n10242), .ZN(n7933) );
  NAND2_X1 U5725 ( .A1(n6982), .A2(n6981), .ZN(n8042) );
  INV_X1 U5726 ( .A(n7933), .ZN(n6982) );
  INV_X1 U5727 ( .A(n8405), .ZN(n8081) );
  AND2_X1 U5728 ( .A1(n8408), .A2(n8407), .ZN(n8405) );
  NAND2_X1 U5729 ( .A1(n7842), .A2(n7841), .ZN(n7939) );
  AND2_X1 U5730 ( .A1(n7845), .A2(n8392), .ZN(n5438) );
  NAND2_X1 U5731 ( .A1(n7601), .A2(n8379), .ZN(n5038) );
  NAND2_X1 U5732 ( .A1(n5270), .A2(n7644), .ZN(n7636) );
  NAND2_X1 U5733 ( .A1(n7634), .A2(n7633), .ZN(n5270) );
  NAND2_X1 U5734 ( .A1(n7470), .A2(n8315), .ZN(n7634) );
  OR2_X1 U5735 ( .A1(n7229), .A2(n7231), .ZN(n7233) );
  NAND2_X1 U5736 ( .A1(n6803), .A2(n6840), .ZN(n8256) );
  CLKBUF_X1 U5737 ( .A(n6946), .Z(n8338) );
  CLKBUF_X1 U5738 ( .A(n6943), .Z(n10563) );
  INV_X1 U5739 ( .A(n8876), .ZN(n8874) );
  INV_X1 U5740 ( .A(n8700), .ZN(n8887) );
  AOI21_X1 U5741 ( .B1(n5273), .B2(n5276), .A(n4980), .ZN(n5272) );
  NAND2_X1 U5742 ( .A1(n8168), .A2(n8167), .ZN(n9035) );
  OR2_X1 U5743 ( .A1(n8165), .A2(n8187), .ZN(n8168) );
  AOI21_X1 U5744 ( .B1(n5420), .B2(n4941), .A(n4978), .ZN(n5034) );
  INV_X1 U5745 ( .A(n8991), .ZN(n8986) );
  NAND2_X1 U5746 ( .A1(n8041), .A2(n8040), .ZN(n8514) );
  NAND2_X1 U5747 ( .A1(n5439), .A2(n8392), .ZN(n7844) );
  NAND2_X1 U5748 ( .A1(n6852), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6560) );
  NAND2_X1 U5749 ( .A1(n5454), .A2(n5452), .ZN(n5451) );
  NOR2_X1 U5750 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n5452) );
  NAND2_X1 U5751 ( .A1(n4960), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6372) );
  XNOR2_X1 U5752 ( .A(n6418), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8505) );
  INV_X1 U5753 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7282) );
  INV_X1 U5754 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6462) );
  OR2_X1 U5755 ( .A1(n6402), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n6406) );
  INV_X1 U5756 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6396) );
  NAND2_X1 U5757 ( .A1(n5054), .A2(n4977), .ZN(n9163) );
  NAND2_X1 U5758 ( .A1(n5085), .A2(n5056), .ZN(n5054) );
  NAND2_X1 U5759 ( .A1(n9243), .A2(n9245), .ZN(n9176) );
  NAND2_X1 U5760 ( .A1(n5669), .A2(n5668), .ZN(n6832) );
  INV_X1 U5761 ( .A(n5667), .ZN(n5668) );
  OR2_X1 U5762 ( .A1(n9205), .A2(n9206), .ZN(n5410) );
  AND2_X1 U5763 ( .A1(n6210), .A2(n6209), .ZN(n9221) );
  XNOR2_X1 U5764 ( .A(n5744), .B(n5745), .ZN(n7104) );
  OR2_X1 U5765 ( .A1(n6090), .A2(n6089), .ZN(n6106) );
  NOR2_X1 U5766 ( .A1(n5934), .A2(n5933), .ZN(n5964) );
  AND2_X1 U5767 ( .A1(n5698), .A2(n5699), .ZN(n6878) );
  NOR2_X1 U5768 ( .A1(n5779), .A2(n7259), .ZN(n5047) );
  NAND2_X1 U5769 ( .A1(n7291), .A2(n7292), .ZN(n7290) );
  NAND2_X1 U5770 ( .A1(n5122), .A2(n5121), .ZN(n9519) );
  NOR2_X1 U5771 ( .A1(n9664), .A2(n9514), .ZN(n5121) );
  NOR4_X1 U5772 ( .A1(n9520), .A2(n9386), .A3(n9385), .A4(n9384), .ZN(n9532)
         );
  NAND2_X1 U5773 ( .A1(n5497), .A2(n5496), .ZN(n9384) );
  NOR3_X1 U5774 ( .A1(n9383), .A2(n9698), .A3(n9679), .ZN(n5496) );
  AND3_X1 U5775 ( .A1(n6451), .A2(n6450), .A3(n6449), .ZN(n9620) );
  INV_X1 U5776 ( .A(n6283), .ZN(n6223) );
  AOI21_X1 U5777 ( .B1(n6771), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6766), .ZN(
        n6914) );
  OR2_X1 U5778 ( .A1(n6914), .A2(n6913), .ZN(n6911) );
  OR2_X1 U5779 ( .A1(n6780), .A2(n6779), .ZN(n6777) );
  NOR2_X1 U5780 ( .A1(n7863), .A2(n7862), .ZN(n7866) );
  AOI21_X1 U5781 ( .B1(n9564), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9563), .ZN(
        n9567) );
  NAND2_X1 U5782 ( .A1(n9711), .A2(n9660), .ZN(n9699) );
  NAND2_X1 U5783 ( .A1(n9661), .A2(n9354), .ZN(n9698) );
  NAND2_X1 U5784 ( .A1(n5139), .A2(n5140), .ZN(n9709) );
  NAND2_X1 U5785 ( .A1(n5139), .A2(n5137), .ZN(n9711) );
  NOR2_X1 U5786 ( .A1(n5138), .A2(n9716), .ZN(n5137) );
  INV_X1 U5787 ( .A(n5140), .ZN(n5138) );
  INV_X1 U5788 ( .A(n5228), .ZN(n5226) );
  NAND2_X1 U5789 ( .A1(n9812), .A2(n4968), .ZN(n9762) );
  NAND2_X1 U5790 ( .A1(n9812), .A2(n5207), .ZN(n9780) );
  OAI21_X1 U5791 ( .B1(n9835), .B2(n9473), .A(n5148), .ZN(n9806) );
  NAND2_X1 U5792 ( .A1(n10031), .A2(n9822), .ZN(n5536) );
  AND2_X1 U5793 ( .A1(n7809), .A2(n4949), .ZN(n9883) );
  NAND2_X1 U5794 ( .A1(n7809), .A2(n5203), .ZN(n8019) );
  NAND2_X1 U5795 ( .A1(n5529), .A2(n4972), .ZN(n5528) );
  AND2_X1 U5796 ( .A1(n9375), .A2(n5532), .ZN(n5530) );
  OR2_X1 U5797 ( .A1(n7962), .A2(n7961), .ZN(n8014) );
  NAND2_X1 U5798 ( .A1(n7809), .A2(n7808), .ZN(n7919) );
  OR2_X1 U5799 ( .A1(n5907), .A2(n5906), .ZN(n5934) );
  OR2_X1 U5800 ( .A1(n5886), .A2(n5885), .ZN(n5907) );
  NAND2_X1 U5801 ( .A1(n7668), .A2(n10648), .ZN(n7718) );
  NAND2_X1 U5802 ( .A1(n7658), .A2(n5524), .ZN(n5521) );
  NAND2_X1 U5803 ( .A1(n7553), .A2(n9409), .ZN(n7710) );
  AOI21_X1 U5804 ( .B1(n9403), .B2(n9398), .A(n5247), .ZN(n7553) );
  INV_X1 U5805 ( .A(n9306), .ZN(n5247) );
  NAND2_X1 U5806 ( .A1(n9410), .A2(n9409), .ZN(n9400) );
  INV_X1 U5807 ( .A(n7344), .ZN(n5041) );
  INV_X1 U5808 ( .A(n9398), .ZN(n7446) );
  NAND2_X1 U5809 ( .A1(n10532), .A2(n7744), .ZN(n9826) );
  NAND2_X1 U5810 ( .A1(n7208), .A2(n7207), .ZN(n5255) );
  CLKBUF_X1 U5811 ( .A(n7494), .Z(n5098) );
  OR2_X1 U5812 ( .A1(n7946), .A2(n5609), .ZN(n7342) );
  NAND2_X1 U5813 ( .A1(n6319), .A2(n5608), .ZN(n7198) );
  AND2_X1 U5814 ( .A1(n6304), .A2(n10044), .ZN(n7340) );
  NAND2_X1 U5815 ( .A1(n9511), .A2(n7744), .ZN(n7946) );
  NAND2_X1 U5816 ( .A1(n9712), .A2(n10704), .ZN(n5263) );
  AOI21_X1 U5817 ( .B1(n9684), .B2(n9852), .A(n9683), .ZN(n9910) );
  OAI211_X1 U5818 ( .C1(n5086), .C2(n6401), .A(n5717), .B(n5716), .ZN(n7214)
         );
  NOR2_X1 U5819 ( .A1(n7220), .A2(n10041), .ZN(n7341) );
  NAND2_X1 U5820 ( .A1(n7814), .A2(n6318), .ZN(n10041) );
  AND2_X1 U5821 ( .A1(n6363), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6318) );
  XNOR2_X1 U5822 ( .A(n8221), .B(n8220), .ZN(n8206) );
  NAND2_X1 U5823 ( .A1(n5465), .A2(n6212), .ZN(n5461) );
  INV_X1 U5824 ( .A(n5459), .ZN(n5458) );
  OAI21_X1 U5825 ( .B1(n5462), .B2(n5460), .A(n5017), .ZN(n5459) );
  AND2_X1 U5826 ( .A1(n5548), .A2(n5957), .ZN(n5605) );
  AOI21_X1 U5827 ( .B1(n6127), .B2(n6126), .A(n6125), .ZN(n6132) );
  NAND2_X1 U5828 ( .A1(n5602), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U5829 ( .A1(n5080), .A2(n5079), .ZN(n5588) );
  NOR2_X1 U5830 ( .A1(n5581), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U5831 ( .A1(n6025), .A2(n6024), .ZN(n6042) );
  OAI21_X1 U5832 ( .B1(n5899), .B2(n5511), .A(n5509), .ZN(n5955) );
  INV_X1 U5833 ( .A(n5510), .ZN(n5509) );
  OAI21_X1 U5834 ( .B1(n5516), .B2(n5511), .A(n5948), .ZN(n5510) );
  INV_X1 U5835 ( .A(n5512), .ZN(n5511) );
  AND2_X1 U5836 ( .A1(n5979), .A2(n5953), .ZN(n5954) );
  NAND2_X1 U5837 ( .A1(n5955), .A2(n5954), .ZN(n5980) );
  AND2_X1 U5838 ( .A1(n5961), .A2(n6006), .ZN(n7623) );
  INV_X1 U5839 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U5840 ( .A1(n5288), .A2(n5286), .ZN(n5815) );
  AOI21_X1 U5841 ( .B1(n5289), .B2(n5290), .A(n5287), .ZN(n5286) );
  INV_X1 U5842 ( .A(n5809), .ZN(n5287) );
  AND2_X1 U5843 ( .A1(n5830), .A2(n5813), .ZN(n5814) );
  INV_X1 U5844 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5558) );
  AND2_X1 U5845 ( .A1(n5556), .A2(n5555), .ZN(n5535) );
  NOR2_X1 U5846 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5679) );
  NAND2_X1 U5847 ( .A1(n5365), .A2(n5370), .ZN(n8567) );
  NAND2_X1 U5848 ( .A1(n8511), .A2(n4936), .ZN(n5365) );
  AND2_X1 U5849 ( .A1(n7989), .A2(n7891), .ZN(n7892) );
  NOR2_X1 U5850 ( .A1(n6857), .A2(n6748), .ZN(n5338) );
  OAI21_X1 U5851 ( .B1(n8523), .B2(n5350), .A(n5348), .ZN(n8584) );
  INV_X1 U5852 ( .A(n5351), .ZN(n5350) );
  AOI21_X1 U5853 ( .B1(n5351), .B2(n5349), .A(n4975), .ZN(n5348) );
  INV_X1 U5854 ( .A(n8709), .ZN(n7883) );
  NAND2_X1 U5855 ( .A1(n8156), .A2(n8155), .ZN(n8922) );
  NAND2_X1 U5856 ( .A1(n8191), .A2(n8190), .ZN(n9026) );
  OR2_X1 U5857 ( .A1(n8188), .A2(n8187), .ZN(n8191) );
  NAND2_X1 U5858 ( .A1(n8180), .A2(n8179), .ZN(n8632) );
  NAND2_X1 U5859 ( .A1(n7733), .A2(n7732), .ZN(n7735) );
  NAND2_X1 U5860 ( .A1(n7733), .A2(n5346), .ZN(n7885) );
  NAND2_X1 U5861 ( .A1(n8511), .A2(n5371), .ZN(n8647) );
  NAND2_X1 U5862 ( .A1(n8535), .A2(n8534), .ZN(n8656) );
  INV_X1 U5863 ( .A(n8676), .ZN(n8691) );
  NAND2_X1 U5864 ( .A1(n5353), .A2(n8524), .ZN(n8664) );
  NAND2_X1 U5865 ( .A1(n5353), .A2(n5351), .ZN(n8665) );
  INV_X1 U5866 ( .A(n8554), .ZN(n8869) );
  OR2_X1 U5867 ( .A1(n6574), .A2(n6948), .ZN(n8679) );
  NAND2_X1 U5868 ( .A1(n5370), .A2(n5369), .ZN(n5364) );
  INV_X1 U5869 ( .A(n5367), .ZN(n5366) );
  NAND2_X1 U5870 ( .A1(n6854), .A2(n8507), .ZN(n8694) );
  INV_X1 U5871 ( .A(n8507), .ZN(n5428) );
  NAND2_X1 U5872 ( .A1(n7052), .A2(n7051), .ZN(n8859) );
  INV_X1 U5873 ( .A(n8907), .ZN(n8624) );
  INV_X1 U5874 ( .A(n7893), .ZN(n8708) );
  NAND4_X1 U5875 ( .A1(n6530), .A2(n6529), .A3(n6528), .A4(n6527), .ZN(n8717)
         );
  NAND2_X1 U5876 ( .A1(n5319), .A2(n5322), .ZN(n6687) );
  AOI21_X1 U5877 ( .B1(n7173), .B2(P2_REG1_REG_5__SCAN_IN), .A(n5180), .ZN(
        n7174) );
  XNOR2_X1 U5878 ( .A(n7391), .B(n7393), .ZN(n7394) );
  NAND2_X1 U5879 ( .A1(n5317), .A2(n7408), .ZN(n7328) );
  NOR2_X1 U5880 ( .A1(n7395), .A2(n7396), .ZN(n7536) );
  NAND2_X1 U5881 ( .A1(n5307), .A2(n5308), .ZN(n7542) );
  NOR2_X1 U5882 ( .A1(n5306), .A2(n8730), .ZN(n8729) );
  AND2_X1 U5883 ( .A1(n6585), .A2(n6609), .ZN(n10371) );
  AND2_X1 U5884 ( .A1(n6496), .A2(n6495), .ZN(n10498) );
  NAND2_X1 U5885 ( .A1(n5437), .A2(n8461), .ZN(n8891) );
  NAND2_X1 U5886 ( .A1(n5278), .A2(n5282), .ZN(n8905) );
  NAND2_X1 U5887 ( .A1(n8929), .A2(n5284), .ZN(n5278) );
  AOI21_X1 U5888 ( .B1(n8929), .B2(n8934), .A(n4954), .ZN(n8917) );
  NAND2_X1 U5889 ( .A1(n5431), .A2(n8233), .ZN(n8933) );
  NAND2_X1 U5890 ( .A1(n8948), .A2(n8941), .ZN(n5431) );
  OAI21_X1 U5891 ( .B1(n8966), .B2(n5294), .A(n5293), .ZN(n8942) );
  NAND2_X1 U5892 ( .A1(n8134), .A2(n8133), .ZN(n8947) );
  NAND2_X1 U5893 ( .A1(n7461), .A2(n8370), .ZN(n7462) );
  OAI21_X1 U5894 ( .B1(n7364), .B2(n8187), .A(n5299), .ZN(n7478) );
  AND2_X1 U5895 ( .A1(n7366), .A2(n5300), .ZN(n5299) );
  NAND2_X1 U5896 ( .A1(n8131), .A2(n5318), .ZN(n5300) );
  OR2_X1 U5897 ( .A1(n6824), .A2(n10571), .ZN(n8937) );
  INV_X1 U5898 ( .A(n9004), .ZN(n8950) );
  INV_X1 U5899 ( .A(n10715), .ZN(n10671) );
  INV_X1 U5900 ( .A(n10570), .ZN(n8983) );
  AOI21_X1 U5901 ( .B1(n8554), .B2(n8994), .A(n8847), .ZN(n8848) );
  NOR2_X1 U5902 ( .A1(n8846), .A2(n10566), .ZN(n8847) );
  AND2_X1 U5903 ( .A1(n7127), .A2(n4961), .ZN(n5090) );
  OR2_X1 U5904 ( .A1(n8187), .A2(n7126), .ZN(n7128) );
  NAND2_X1 U5905 ( .A1(n10723), .A2(n10671), .ZN(n9050) );
  INV_X1 U5906 ( .A(n10723), .ZN(n10721) );
  AND2_X1 U5907 ( .A1(n5450), .A2(n5449), .ZN(n8843) );
  NAND2_X1 U5908 ( .A1(n8205), .A2(n8204), .ZN(n9080) );
  OR2_X1 U5909 ( .A1(n8208), .A2(n8266), .ZN(n8204) );
  NAND2_X1 U5910 ( .A1(n8202), .A2(n8201), .ZN(n9086) );
  OR2_X1 U5911 ( .A1(n8208), .A2(n9160), .ZN(n8201) );
  NAND2_X1 U5912 ( .A1(n5271), .A2(n5276), .ZN(n8896) );
  OR2_X1 U5913 ( .A1(n8929), .A2(n5277), .ZN(n5271) );
  INV_X1 U5914 ( .A(n8947), .ZN(n9120) );
  NAND2_X1 U5915 ( .A1(n8121), .A2(n8120), .ZN(n9123) );
  NAND2_X1 U5916 ( .A1(n8964), .A2(n5554), .ZN(n8956) );
  AND2_X1 U5917 ( .A1(n8969), .A2(n8968), .ZN(n9128) );
  INV_X1 U5918 ( .A(n5419), .ZN(n8962) );
  AOI21_X1 U5919 ( .B1(n8974), .B2(n8973), .A(n4955), .ZN(n5419) );
  AND2_X1 U5920 ( .A1(n8981), .A2(n8980), .ZN(n9134) );
  AND2_X1 U5921 ( .A1(n8998), .A2(n8997), .ZN(n9140) );
  OAI21_X1 U5922 ( .B1(n8052), .B2(n5269), .A(n4933), .ZN(n8990) );
  INV_X1 U5923 ( .A(n8514), .ZN(n8575) );
  AND2_X1 U5924 ( .A1(n8086), .A2(n8407), .ZN(n8048) );
  AND2_X1 U5925 ( .A1(n10727), .A2(n10671), .ZN(n9141) );
  AND2_X2 U5926 ( .A1(n6848), .A2(n6847), .ZN(n10727) );
  CLKBUF_X1 U5927 ( .A(n6482), .Z(n6483) );
  XNOR2_X1 U5928 ( .A(n6376), .B(n6375), .ZN(n7956) );
  NAND2_X1 U5929 ( .A1(n6374), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6376) );
  MUX2_X1 U5930 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6378), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n6379) );
  NAND2_X1 U5931 ( .A1(n6551), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6415) );
  INV_X1 U5932 ( .A(n10388), .ZN(n8804) );
  NAND2_X1 U5933 ( .A1(n5309), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6391) );
  AND3_X1 U5934 ( .A1(n9176), .A2(n9174), .A3(n9175), .ZN(n9223) );
  NAND2_X1 U5935 ( .A1(n5403), .A2(n5896), .ZN(n7819) );
  NAND2_X1 U5936 ( .A1(n5400), .A2(n5897), .ZN(n7820) );
  OAI21_X1 U5937 ( .B1(n7761), .B2(n5726), .A(n5884), .ZN(n10680) );
  AND2_X1 U5938 ( .A1(n5070), .A2(n5061), .ZN(n5068) );
  NAND2_X1 U5939 ( .A1(n6085), .A2(n6084), .ZN(n9962) );
  INV_X1 U5940 ( .A(n6323), .ZN(n6358) );
  NAND2_X1 U5941 ( .A1(n5072), .A2(n5071), .ZN(n7900) );
  AOI21_X1 U5942 ( .B1(n5394), .B2(n5073), .A(n5023), .ZN(n5072) );
  NOR2_X1 U5943 ( .A1(n5398), .A2(n7873), .ZN(n5073) );
  AND2_X1 U5944 ( .A1(n5410), .A2(n4953), .ZN(n9215) );
  OAI21_X1 U5945 ( .B1(n6185), .B2(n5053), .A(n5051), .ZN(n9220) );
  XNOR2_X1 U5946 ( .A(n5749), .B(n5747), .ZN(n7089) );
  OAI21_X1 U5947 ( .B1(n7006), .B2(n5726), .A(n5214), .ZN(n10597) );
  NOR2_X1 U5948 ( .A1(n4958), .A2(n5215), .ZN(n5214) );
  NOR2_X1 U5949 ( .A1(n5648), .A2(n6918), .ZN(n5215) );
  NAND2_X1 U5950 ( .A1(n5130), .A2(n5858), .ZN(n10662) );
  NAND2_X1 U5951 ( .A1(n7580), .A2(n9335), .ZN(n5130) );
  NAND2_X1 U5952 ( .A1(n5416), .A2(n5947), .ZN(n8004) );
  NAND2_X1 U5953 ( .A1(n5416), .A2(n5413), .ZN(n8005) );
  NAND2_X1 U5954 ( .A1(n6694), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9275) );
  NAND2_X1 U5955 ( .A1(n5075), .A2(n5394), .ZN(n7875) );
  NAND2_X1 U5956 ( .A1(n7696), .A2(n5398), .ZN(n5075) );
  AOI21_X1 U5957 ( .B1(n4938), .B2(n9206), .A(n5009), .ZN(n5408) );
  INV_X1 U5958 ( .A(n7456), .ZN(n10622) );
  OR2_X1 U5959 ( .A1(n5751), .A2(n5654), .ZN(n5658) );
  OR2_X1 U5960 ( .A1(n5755), .A2(n5655), .ZN(n5657) );
  OR2_X1 U5961 ( .A1(n5755), .A2(n5619), .ZN(n5625) );
  OR2_X1 U5962 ( .A1(n5751), .A2(n10521), .ZN(n5624) );
  XNOR2_X1 U5963 ( .A(n6333), .B(P1_IR_REG_28__SCAN_IN), .ZN(n10347) );
  AOI21_X1 U5964 ( .B1(n6630), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6953), .ZN(
        n6768) );
  NOR2_X1 U5965 ( .A1(n6768), .A2(n6767), .ZN(n6766) );
  AND2_X1 U5966 ( .A1(n6911), .A2(n6635), .ZN(n6642) );
  AOI21_X1 U5967 ( .B1(n6656), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6655), .ZN(
        n6780) );
  NAND2_X1 U5968 ( .A1(n6727), .A2(n5097), .ZN(n6729) );
  OR2_X1 U5969 ( .A1(n6728), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5097) );
  AOI21_X1 U5970 ( .B1(n6886), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6885), .ZN(
        n6888) );
  AOI21_X1 U5971 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9602), .A(n9601), .ZN(
        n9604) );
  NAND2_X1 U5972 ( .A1(n5143), .A2(n9657), .ZN(n9727) );
  OR2_X1 U5973 ( .A1(n9752), .A2(n9751), .ZN(n5143) );
  NAND2_X1 U5974 ( .A1(n9773), .A2(n9655), .ZN(n9757) );
  NAND2_X1 U5975 ( .A1(n5223), .A2(n5227), .ZN(n9761) );
  OR2_X1 U5976 ( .A1(n9804), .A2(n5228), .ZN(n5223) );
  NAND2_X1 U5977 ( .A1(n9654), .A2(n9653), .ZN(n9775) );
  NAND2_X1 U5978 ( .A1(n5229), .A2(n5232), .ZN(n9772) );
  NAND2_X1 U5979 ( .A1(n9804), .A2(n5233), .ZN(n5229) );
  AOI21_X1 U5980 ( .B1(n9804), .B2(n9803), .A(n4935), .ZN(n9794) );
  OR2_X1 U5981 ( .A1(n8153), .A2(n5726), .ZN(n6137) );
  AND2_X1 U5982 ( .A1(n5152), .A2(n5153), .ZN(n9820) );
  NAND2_X1 U5983 ( .A1(n9835), .A2(n9840), .ZN(n5152) );
  NAND2_X1 U5984 ( .A1(n9874), .A2(n9466), .ZN(n9850) );
  INV_X1 U5985 ( .A(n9554), .ZN(n9975) );
  NAND2_X1 U5986 ( .A1(n6049), .A2(n6048), .ZN(n9868) );
  NAND2_X1 U5987 ( .A1(n9342), .A2(n9468), .ZN(n9876) );
  INV_X1 U5988 ( .A(n9555), .ZN(n9987) );
  INV_X1 U5989 ( .A(n5527), .ZN(n7959) );
  AOI21_X1 U5990 ( .B1(n5534), .B2(n5532), .A(n4959), .ZN(n5527) );
  OR2_X1 U5991 ( .A1(n7805), .A2(n7804), .ZN(n5531) );
  NAND2_X1 U5992 ( .A1(n5523), .A2(n7661), .ZN(n7675) );
  NAND2_X1 U5993 ( .A1(n7658), .A2(n7657), .ZN(n5523) );
  INV_X1 U5994 ( .A(n9559), .ZN(n10632) );
  NAND2_X1 U5995 ( .A1(n5820), .A2(n5819), .ZN(n7566) );
  INV_X1 U5996 ( .A(n10597), .ZN(n7522) );
  OR2_X1 U5997 ( .A1(n5751), .A2(n7351), .ZN(n5676) );
  OR2_X1 U5998 ( .A1(n5755), .A2(n5672), .ZN(n5674) );
  INV_X1 U5999 ( .A(n9888), .ZN(n9869) );
  INV_X1 U6000 ( .A(n9891), .ZN(n9865) );
  OR2_X1 U6001 ( .A1(n7342), .A2(n10041), .ZN(n10522) );
  NOR2_X1 U6002 ( .A1(n9903), .A2(n5210), .ZN(n9905) );
  NAND2_X1 U6003 ( .A1(n5211), .A2(n5008), .ZN(n5210) );
  NAND2_X1 U6004 ( .A1(n9904), .A2(n10705), .ZN(n5211) );
  INV_X1 U6005 ( .A(n9621), .ZN(n9995) );
  INV_X1 U6006 ( .A(n7958), .ZN(n8033) );
  INV_X1 U6007 ( .A(n7802), .ZN(n7955) );
  AND2_X1 U6008 ( .A1(n5614), .A2(n5617), .ZN(n5264) );
  XNOR2_X1 U6009 ( .A(n8282), .B(n8281), .ZN(n10050) );
  NAND2_X1 U6010 ( .A1(n8287), .A2(n8286), .ZN(n10055) );
  OAI21_X1 U6011 ( .B1(n5602), .B2(n5601), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5417) );
  NAND2_X1 U6012 ( .A1(n6168), .A2(n6167), .ZN(n6190) );
  OR2_X1 U6013 ( .A1(n5586), .A2(n5600), .ZN(n5587) );
  NAND2_X1 U6014 ( .A1(n5506), .A2(n5504), .ZN(n6004) );
  NAND2_X1 U6015 ( .A1(n5513), .A2(n5512), .ZN(n5949) );
  NAND2_X1 U6016 ( .A1(n5513), .A2(n5514), .ZN(n5926) );
  NAND2_X1 U6017 ( .A1(n5108), .A2(n5899), .ZN(n7761) );
  NAND2_X1 U6018 ( .A1(n5475), .A2(n5880), .ZN(n5108) );
  NAND2_X1 U6019 ( .A1(n5831), .A2(n5816), .ZN(n7364) );
  OR2_X1 U6020 ( .A1(n5815), .A2(n5814), .ZN(n5816) );
  OAI21_X1 U6021 ( .B1(n5769), .B2(n5290), .A(n5289), .ZN(n5810) );
  NAND2_X1 U6022 ( .A1(n5788), .A2(n5037), .ZN(n5036) );
  NOR2_X1 U6023 ( .A1(n5792), .A2(n5290), .ZN(n5037) );
  NAND2_X1 U6024 ( .A1(n5456), .A2(n5685), .ZN(n5688) );
  NAND2_X1 U6025 ( .A1(n5105), .A2(n5682), .ZN(n5646) );
  NAND2_X1 U6026 ( .A1(n5384), .A2(n8685), .ZN(n5382) );
  NAND2_X1 U6027 ( .A1(n4995), .A2(n5428), .ZN(n5424) );
  AOI21_X1 U6028 ( .B1(n5201), .B2(n10483), .A(n5198), .ZN(n10517) );
  NAND2_X1 U6029 ( .A1(n5331), .A2(n5326), .ZN(P2_U3201) );
  INV_X1 U6030 ( .A(n5327), .ZN(n5326) );
  OAI21_X1 U6031 ( .B1(n8834), .B2(n10496), .A(n5328), .ZN(n5327) );
  AND2_X1 U6032 ( .A1(n7814), .A2(n6364), .ZN(P1_U3973) );
  AOI21_X1 U6033 ( .B1(n9260), .B2(n5043), .A(n5020), .ZN(n5044) );
  AOI211_X1 U6034 ( .C1(n9724), .C2(n9281), .A(n9265), .B(n9264), .ZN(n9266)
         );
  OR2_X1 U6035 ( .A1(n9593), .A2(n5087), .ZN(P1_U3261) );
  AOI21_X1 U6036 ( .B1(n10350), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n9594), .ZN(
        n5088) );
  OAI211_X1 U6037 ( .C1(n9906), .C2(n9685), .A(n5156), .B(n5154), .ZN(P1_U3356) );
  AOI21_X1 U6038 ( .B1(n9903), .B2(n9891), .A(n9669), .ZN(n5156) );
  NAND2_X1 U6039 ( .A1(n5155), .A2(n9855), .ZN(n5154) );
  OAI21_X1 U6040 ( .B1(n10001), .B2(n10735), .A(n5238), .ZN(P1_U3550) );
  INV_X1 U6041 ( .A(n5239), .ZN(n5238) );
  OAI22_X1 U6042 ( .A1(n10003), .A2(n9991), .B1(n10736), .B2(n9913), .ZN(n5239) );
  NAND2_X1 U6043 ( .A1(n10740), .A2(n10711), .ZN(n5544) );
  INV_X1 U6044 ( .A(n5539), .ZN(n5538) );
  OAI21_X1 U6045 ( .B1(n9906), .B2(n10737), .A(n5540), .ZN(n5539) );
  OAI21_X1 U6046 ( .B1(n10001), .B2(n10737), .A(n5261), .ZN(P1_U3518) );
  INV_X1 U6047 ( .A(n5262), .ZN(n5261) );
  OAI22_X1 U6048 ( .A1(n10003), .A2(n10040), .B1(n10740), .B2(n10002), .ZN(
        n5262) );
  XNOR2_X2 U6049 ( .A(n5591), .B(n5590), .ZN(n5608) );
  AND2_X1 U6050 ( .A1(n8991), .A2(n5268), .ZN(n4933) );
  AND2_X1 U6051 ( .A1(n7326), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4934) );
  AND2_X1 U6052 ( .A1(n9823), .A2(n5153), .ZN(n5151) );
  NAND2_X1 U6053 ( .A1(n6137), .A2(n6136), .ZN(n9800) );
  INV_X1 U6054 ( .A(n9800), .ZN(n5236) );
  AND2_X1 U6055 ( .A1(n8475), .A2(n8476), .ZN(n8856) );
  NOR2_X1 U6056 ( .A1(n9813), .A2(n9553), .ZN(n4935) );
  AND2_X1 U6057 ( .A1(n4973), .A2(n5371), .ZN(n4936) );
  OR2_X1 U6058 ( .A1(n9222), .A2(n5406), .ZN(n4937) );
  AND2_X1 U6059 ( .A1(n5550), .A2(n4953), .ZN(n4938) );
  AND2_X1 U6060 ( .A1(n5490), .A2(n5013), .ZN(n4939) );
  NAND2_X1 U6061 ( .A1(n7465), .A2(n7471), .ZN(n8370) );
  NAND2_X1 U6062 ( .A1(n6073), .A2(n6072), .ZN(n9847) );
  INV_X1 U6063 ( .A(n9847), .ZN(n10031) );
  AND2_X1 U6064 ( .A1(n5068), .A2(n5069), .ZN(n4940) );
  OR2_X1 U6065 ( .A1(n4955), .A2(n5418), .ZN(n4941) );
  OR2_X1 U6066 ( .A1(n8240), .A2(n8300), .ZN(n4942) );
  AND2_X1 U6067 ( .A1(n5226), .A2(n9640), .ZN(n4943) );
  AND2_X1 U6068 ( .A1(n9142), .A2(n8978), .ZN(n4944) );
  AND2_X1 U6069 ( .A1(n5501), .A2(n5014), .ZN(n4945) );
  NAND2_X1 U6070 ( .A1(n9291), .A2(n9290), .ZN(n9904) );
  INV_X1 U6071 ( .A(n9904), .ZN(n5499) );
  AOI21_X1 U6072 ( .B1(n5233), .B2(n4935), .A(n4991), .ZN(n5232) );
  NAND2_X1 U6073 ( .A1(n5494), .A2(n5010), .ZN(n4946) );
  NOR2_X1 U6074 ( .A1(n5429), .A2(n7418), .ZN(n4947) );
  AND4_X1 U6075 ( .A1(n5960), .A2(n6026), .A3(n5564), .A4(n5582), .ZN(n4948)
         );
  AND2_X1 U6076 ( .A1(n5203), .A2(n5202), .ZN(n4949) );
  INV_X1 U6077 ( .A(n5114), .ZN(n5113) );
  OAI21_X1 U6078 ( .B1(n5116), .B2(n4982), .A(n9502), .ZN(n5114) );
  AND2_X1 U6079 ( .A1(n5848), .A2(n5829), .ZN(n4950) );
  INV_X1 U6080 ( .A(n9636), .ZN(n5251) );
  INV_X1 U6081 ( .A(n9642), .ZN(n9921) );
  NAND2_X1 U6082 ( .A1(n9812), .A2(n5209), .ZN(n4951) );
  NAND2_X1 U6083 ( .A1(n9962), .A2(n9836), .ZN(n4952) );
  INV_X1 U6084 ( .A(n9712), .ZN(n9911) );
  NAND2_X1 U6085 ( .A1(n7809), .A2(n5205), .ZN(n5206) );
  NAND2_X1 U6086 ( .A1(n5599), .A2(n5598), .ZN(n6299) );
  NAND2_X1 U6087 ( .A1(n6551), .A2(n6550), .ZN(n7691) );
  AND2_X2 U6088 ( .A1(n5928), .A2(n5561), .ZN(n5957) );
  NAND2_X1 U6089 ( .A1(n6040), .A2(n6039), .ZN(n4953) );
  AND2_X1 U6090 ( .A1(n9115), .A2(n8944), .ZN(n4954) );
  NOR2_X1 U6091 ( .A1(n9135), .A2(n8619), .ZN(n4955) );
  NAND2_X1 U6092 ( .A1(n7268), .A2(n6371), .ZN(n6383) );
  NAND2_X1 U6093 ( .A1(n5404), .A2(n5407), .ZN(n9174) );
  NAND2_X1 U6094 ( .A1(n8243), .A2(n8299), .ZN(n4956) );
  OR2_X1 U6095 ( .A1(n8867), .A2(n8469), .ZN(n4957) );
  INV_X1 U6096 ( .A(n5433), .ZN(n5432) );
  OAI21_X1 U6097 ( .B1(n8941), .B2(n5434), .A(n8928), .ZN(n5433) );
  NOR2_X1 U6098 ( .A1(n9296), .A2(n6398), .ZN(n4958) );
  AND2_X1 U6099 ( .A1(n10706), .A2(n9556), .ZN(n4959) );
  INV_X1 U6100 ( .A(n5778), .ZN(n5779) );
  INV_X1 U6101 ( .A(n5475), .ZN(n5879) );
  OR2_X1 U6102 ( .A1(n6374), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4960) );
  INV_X1 U6103 ( .A(n9466), .ZN(n5119) );
  NAND2_X1 U6104 ( .A1(n8523), .A2(n8522), .ZN(n8614) );
  OR2_X1 U6105 ( .A1(n8249), .A2(n7177), .ZN(n4961) );
  INV_X1 U6106 ( .A(n9809), .ZN(n9778) );
  OAI21_X1 U6107 ( .B1(n5648), .B2(n5576), .A(n5575), .ZN(n10533) );
  AND2_X1 U6108 ( .A1(n5768), .A2(n5787), .ZN(n4962) );
  NAND2_X1 U6109 ( .A1(n8494), .A2(n8478), .ZN(n8480) );
  INV_X1 U6110 ( .A(n8480), .ZN(n8247) );
  INV_X1 U6111 ( .A(n8715), .ZN(n10565) );
  INV_X1 U6112 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6394) );
  INV_X1 U6113 ( .A(n7901), .ZN(n5084) );
  INV_X1 U6114 ( .A(n6184), .ZN(n5407) );
  NAND2_X1 U6115 ( .A1(n9517), .A2(n9516), .ZN(n9664) );
  INV_X1 U6116 ( .A(n9664), .ZN(n5497) );
  NAND2_X1 U6117 ( .A1(n6170), .A2(n6169), .ZN(n9764) );
  INV_X1 U6118 ( .A(n9764), .ZN(n10019) );
  OR2_X1 U6119 ( .A1(n9100), .A2(n8907), .ZN(n4963) );
  NAND2_X1 U6120 ( .A1(n5069), .A2(n5070), .ZN(n9182) );
  AND3_X1 U6121 ( .A1(n5900), .A2(n5881), .A3(n5560), .ZN(n4964) );
  INV_X1 U6122 ( .A(n8418), .ZN(n5269) );
  AND2_X1 U6123 ( .A1(n10557), .A2(n5162), .ZN(n4965) );
  NAND2_X1 U6124 ( .A1(n5931), .A2(n5930), .ZN(n10706) );
  OR2_X1 U6125 ( .A1(n8553), .A2(n5388), .ZN(n4966) );
  NOR2_X1 U6126 ( .A1(n9296), .A2(n6407), .ZN(n4967) );
  AND2_X1 U6127 ( .A1(n5207), .A2(n10019), .ZN(n4968) );
  NAND2_X1 U6128 ( .A1(n5681), .A2(n5705), .ZN(n6961) );
  NAND2_X1 U6129 ( .A1(n5983), .A2(n5982), .ZN(n9171) );
  INV_X1 U6130 ( .A(n9944), .ZN(n9786) );
  AND2_X1 U6131 ( .A1(n8425), .A2(n5164), .ZN(n4969) );
  AND2_X1 U6132 ( .A1(n6518), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4970) );
  INV_X1 U6133 ( .A(n9813), .ZN(n9614) );
  NAND2_X1 U6134 ( .A1(n6105), .A2(n6104), .ZN(n9813) );
  AND2_X1 U6135 ( .A1(n8542), .A2(n5373), .ZN(n4971) );
  NAND2_X1 U6136 ( .A1(n7958), .A2(n7964), .ZN(n4972) );
  OR2_X1 U6137 ( .A1(n8645), .A2(n8569), .ZN(n4973) );
  NOR2_X1 U6138 ( .A1(n7986), .A2(n8707), .ZN(n4974) );
  AND2_X1 U6139 ( .A1(n8526), .A2(n8967), .ZN(n4975) );
  INV_X1 U6140 ( .A(n5414), .ZN(n5413) );
  NAND2_X1 U6141 ( .A1(n5415), .A2(n5947), .ZN(n5414) );
  AND2_X1 U6142 ( .A1(n8347), .A2(n8346), .ZN(n4976) );
  AND2_X1 U6143 ( .A1(n5055), .A2(n5997), .ZN(n4977) );
  INV_X1 U6144 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6375) );
  OR2_X1 U6145 ( .A1(n8430), .A2(n8668), .ZN(n5554) );
  NOR2_X1 U6146 ( .A1(n9129), .A2(n8668), .ZN(n4978) );
  NOR2_X1 U6147 ( .A1(n7884), .A2(n7883), .ZN(n4979) );
  NOR2_X1 U6148 ( .A1(n8902), .A2(n8624), .ZN(n4980) );
  NOR2_X1 U6149 ( .A1(n8642), .A2(n8944), .ZN(n4981) );
  AND2_X1 U6150 ( .A1(n9743), .A2(n9498), .ZN(n4982) );
  INV_X1 U6151 ( .A(n5455), .ZN(n5454) );
  NAND2_X1 U6152 ( .A1(n6408), .A2(n6410), .ZN(n5455) );
  INV_X1 U6153 ( .A(n5505), .ZN(n5504) );
  NOR2_X1 U6154 ( .A1(n5999), .A2(SI_14_), .ZN(n5505) );
  INV_X1 U6155 ( .A(n5515), .ZN(n5514) );
  NOR2_X1 U6156 ( .A1(n5921), .A2(SI_11_), .ZN(n5515) );
  INV_X1 U6157 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5638) );
  OAI21_X1 U6158 ( .B1(n9175), .B2(n9222), .A(n9221), .ZN(n5405) );
  INV_X1 U6159 ( .A(n5457), .ZN(n6218) );
  OAI21_X1 U6160 ( .B1(n6158), .B2(n5461), .A(n5458), .ZN(n5457) );
  INV_X1 U6161 ( .A(n7873), .ZN(n5074) );
  OR2_X1 U6162 ( .A1(n8249), .A2(n4931), .ZN(n4983) );
  NAND2_X1 U6163 ( .A1(n9680), .A2(n9679), .ZN(n4984) );
  INV_X1 U6164 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5486) );
  NOR2_X1 U6165 ( .A1(n9120), .A2(n8931), .ZN(n4985) );
  INV_X1 U6166 ( .A(n5421), .ZN(n5420) );
  OAI21_X1 U6167 ( .B1(n8973), .B2(n4955), .A(n8963), .ZN(n5421) );
  INV_X1 U6168 ( .A(n6856), .ZN(n6857) );
  NAND2_X1 U6169 ( .A1(n8494), .A2(n8299), .ZN(n4986) );
  OR2_X1 U6170 ( .A1(n5873), .A2(SI_9_), .ZN(n4987) );
  AND2_X1 U6171 ( .A1(n9035), .A2(n8702), .ZN(n4988) );
  NAND2_X1 U6172 ( .A1(n9764), .A2(n9639), .ZN(n4989) );
  INV_X1 U6173 ( .A(n6000), .ZN(n5507) );
  XNOR2_X1 U6174 ( .A(n5999), .B(SI_14_), .ZN(n6000) );
  OR2_X1 U6175 ( .A1(n5455), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4990) );
  OAI21_X1 U6176 ( .B1(n9233), .B2(n5064), .A(n9232), .ZN(n5063) );
  OAI21_X1 U6177 ( .B1(n5227), .B2(n5225), .A(n4989), .ZN(n5224) );
  AND2_X1 U6178 ( .A1(n5236), .A2(n9778), .ZN(n4991) );
  OAI21_X1 U6179 ( .B1(n5174), .B2(n4957), .A(n5176), .ZN(n5173) );
  INV_X1 U6180 ( .A(n8371), .ZN(n8315) );
  AND2_X1 U6181 ( .A1(n8378), .A2(n7643), .ZN(n8371) );
  NAND2_X1 U6182 ( .A1(n8490), .A2(n8478), .ZN(n4992) );
  NAND2_X1 U6183 ( .A1(n5978), .A2(n5996), .ZN(n4993) );
  AND2_X1 U6184 ( .A1(n8371), .A2(n8370), .ZN(n4994) );
  AND2_X1 U6185 ( .A1(n5425), .A2(n8833), .ZN(n4995) );
  INV_X1 U6186 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5582) );
  AND3_X1 U6187 ( .A1(n5594), .A2(n5592), .A3(n6316), .ZN(n4996) );
  NAND2_X1 U6188 ( .A1(n5230), .A2(n9776), .ZN(n4997) );
  AND2_X1 U6189 ( .A1(n9909), .A2(n5263), .ZN(n4998) );
  AND2_X1 U6190 ( .A1(n9868), .A2(n9635), .ZN(n4999) );
  NOR2_X1 U6191 ( .A1(n7676), .A2(n10661), .ZN(n5000) );
  NOR2_X1 U6192 ( .A1(n6003), .A2(n5505), .ZN(n5502) );
  AND3_X1 U6193 ( .A1(n5440), .A2(n5357), .A3(n6395), .ZN(n5001) );
  OR2_X1 U6194 ( .A1(n10031), .A2(n9822), .ZN(n5002) );
  AND2_X1 U6195 ( .A1(n9469), .A2(n9466), .ZN(n9872) );
  AND2_X1 U6196 ( .A1(n5112), .A2(n9660), .ZN(n5003) );
  NAND2_X1 U6197 ( .A1(n5633), .A2(n6291), .ZN(n5653) );
  INV_X1 U6198 ( .A(n8128), .ZN(n5297) );
  AND2_X1 U6199 ( .A1(n9123), .A2(n8967), .ZN(n8128) );
  INV_X1 U6200 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5617) );
  OR2_X1 U6201 ( .A1(n9222), .A2(n6184), .ZN(n5004) );
  INV_X1 U6202 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5305) );
  INV_X1 U6203 ( .A(n6074), .ZN(n5844) );
  AND2_X1 U6204 ( .A1(n6363), .A2(n6328), .ZN(n6074) );
  INV_X1 U6205 ( .A(n9840), .ZN(n5150) );
  INV_X1 U6206 ( .A(n9851), .ZN(n9822) );
  NAND2_X1 U6207 ( .A1(n5334), .A2(n7989), .ZN(n7990) );
  AND2_X1 U6208 ( .A1(n9812), .A2(n9614), .ZN(n5005) );
  NOR2_X1 U6209 ( .A1(n10003), .A2(n9902), .ZN(n5006) );
  OR2_X1 U6211 ( .A1(n8674), .A2(n8859), .ZN(n5007) );
  INV_X1 U6212 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5219) );
  INV_X1 U6213 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5220) );
  OR2_X1 U6214 ( .A1(n9902), .A2(n10631), .ZN(n5008) );
  OAI21_X1 U6215 ( .B1(n8231), .B2(n5421), .A(n5034), .ZN(n8954) );
  NAND2_X1 U6216 ( .A1(n5531), .A2(n7803), .ZN(n7918) );
  INV_X1 U6217 ( .A(n9658), .ZN(n5145) );
  XNOR2_X1 U6218 ( .A(n6436), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7571) );
  AND2_X1 U6219 ( .A1(n9213), .A2(n6059), .ZN(n5009) );
  INV_X1 U6220 ( .A(n5857), .ZN(n5080) );
  NOR2_X1 U6221 ( .A1(n9844), .A2(n9962), .ZN(n9812) );
  OR2_X1 U6222 ( .A1(n6060), .A2(SI_17_), .ZN(n5010) );
  NAND2_X1 U6223 ( .A1(n5817), .A2(n5559), .ZN(n5832) );
  NAND2_X1 U6224 ( .A1(n6222), .A2(n6221), .ZN(n9735) );
  INV_X1 U6225 ( .A(n9735), .ZN(n10014) );
  INV_X1 U6226 ( .A(n8569), .ZN(n8705) );
  AND4_X1 U6227 ( .A1(n7938), .A2(n7937), .A3(n7936), .A4(n7935), .ZN(n8569)
         );
  NAND2_X1 U6228 ( .A1(n8052), .A2(n8326), .ZN(n8105) );
  AND2_X1 U6229 ( .A1(n8035), .A2(n8034), .ZN(n5011) );
  OR2_X1 U6230 ( .A1(n10014), .A2(n9921), .ZN(n5012) );
  AND2_X1 U6231 ( .A1(n5495), .A2(n6081), .ZN(n5013) );
  AND2_X1 U6232 ( .A1(n5503), .A2(n6024), .ZN(n5014) );
  NAND2_X1 U6233 ( .A1(n6260), .A2(n6259), .ZN(n9693) );
  NOR2_X1 U6234 ( .A1(n9824), .A2(n9823), .ZN(n9965) );
  INV_X1 U6235 ( .A(n9965), .ZN(n5089) );
  AND2_X1 U6236 ( .A1(n8804), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5015) );
  OR2_X1 U6237 ( .A1(n8237), .A2(n9015), .ZN(n5016) );
  INV_X1 U6238 ( .A(n8516), .ZN(n5369) );
  OR2_X1 U6239 ( .A1(n6211), .A2(SI_24_), .ZN(n5017) );
  AND2_X1 U6240 ( .A1(n6188), .A2(n10162), .ZN(n5018) );
  AND2_X1 U6241 ( .A1(n6101), .A2(n10192), .ZN(n5019) );
  INV_X1 U6242 ( .A(n5465), .ZN(n5464) );
  NOR2_X1 U6243 ( .A1(n6189), .A2(n5466), .ZN(n5465) );
  NAND2_X1 U6244 ( .A1(n6362), .A2(n6361), .ZN(n5020) );
  INV_X1 U6245 ( .A(n5370), .ZN(n5368) );
  NAND2_X1 U6246 ( .A1(n8645), .A2(n8569), .ZN(n5370) );
  OR2_X1 U6247 ( .A1(n8615), .A2(n8668), .ZN(n5021) );
  INV_X1 U6248 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5562) );
  INV_X1 U6249 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6369) );
  INV_X1 U6250 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5600) );
  XNOR2_X1 U6251 ( .A(n5595), .B(n5594), .ZN(n7744) );
  NAND2_X1 U6252 ( .A1(n6009), .A2(n6008), .ZN(n9632) );
  INV_X1 U6253 ( .A(n9632), .ZN(n5202) );
  INV_X1 U6254 ( .A(n9894), .ZN(n9855) );
  INV_X1 U6255 ( .A(n8683), .ZN(n8685) );
  NAND2_X1 U6256 ( .A1(n4994), .A2(n7461), .ZN(n7600) );
  INV_X1 U6257 ( .A(n5332), .ZN(n6810) );
  OAI21_X1 U6258 ( .B1(n6547), .B2(P2_D_REG_0__SCAN_IN), .A(n6534), .ZN(n5332)
         );
  NAND2_X1 U6259 ( .A1(n5081), .A2(n7649), .ZN(n7696) );
  NAND2_X1 U6260 ( .A1(n6427), .A2(n6428), .ZN(n6547) );
  OR2_X1 U6261 ( .A1(n10740), .A2(n5545), .ZN(n5022) );
  OR2_X1 U6262 ( .A1(n6562), .A2(n6561), .ZN(n8683) );
  AND2_X1 U6263 ( .A1(n5920), .A2(n5919), .ZN(n5023) );
  AND4_X1 U6264 ( .A1(n6341), .A2(n6340), .A3(n6339), .A4(n6338), .ZN(n9682)
         );
  INV_X1 U6265 ( .A(n9682), .ZN(n5498) );
  OR2_X1 U6266 ( .A1(n5857), .A2(n5581), .ZN(n5024) );
  AND2_X1 U6267 ( .A1(n5588), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5025) );
  AND2_X1 U6268 ( .A1(n6279), .A2(n6278), .ZN(n5026) );
  INV_X1 U6269 ( .A(n8730), .ZN(n5307) );
  AND3_X2 U6270 ( .A1(n7225), .A2(n7341), .A3(n7339), .ZN(n10740) );
  AND3_X2 U6271 ( .A1(n7225), .A2(n7341), .A3(n7224), .ZN(n10736) );
  INV_X1 U6272 ( .A(n10457), .ZN(n8787) );
  INV_X1 U6273 ( .A(n10423), .ZN(n8795) );
  INV_X1 U6274 ( .A(n10496), .ZN(n10483) );
  OR2_X1 U6275 ( .A1(n10360), .A2(n9596), .ZN(n5027) );
  OR2_X1 U6276 ( .A1(n6332), .A2(n6331), .ZN(n6638) );
  AND2_X1 U6277 ( .A1(n7786), .A2(n7946), .ZN(n10528) );
  AND2_X1 U6278 ( .A1(n5340), .A2(n5341), .ZN(n5028) );
  NAND3_X1 U6279 ( .A1(n5548), .A2(n5957), .A3(n5264), .ZN(n5265) );
  INV_X1 U6280 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5096) );
  AND2_X1 U6281 ( .A1(n5428), .A2(n7418), .ZN(n5029) );
  INV_X1 U6282 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5179) );
  NAND2_X1 U6283 ( .A1(n7057), .A2(n7177), .ZN(n7184) );
  NAND3_X1 U6284 ( .A1(n5031), .A2(n8234), .A3(n5030), .ZN(n8909) );
  NAND2_X1 U6285 ( .A1(n5033), .A2(n5430), .ZN(n8920) );
  NAND2_X1 U6286 ( .A1(n8948), .A2(n5432), .ZN(n5033) );
  NAND2_X1 U6287 ( .A1(n7273), .A2(n8313), .ZN(n7272) );
  NAND2_X1 U6288 ( .A1(n8865), .A2(n8471), .ZN(n8235) );
  NAND3_X1 U6289 ( .A1(n5105), .A2(n5682), .A3(n5644), .ZN(n5683) );
  INV_X1 U6290 ( .A(n5038), .ZN(n7760) );
  XNOR2_X1 U6291 ( .A(n5038), .B(n8320), .ZN(n10670) );
  NAND2_X1 U6292 ( .A1(n7931), .A2(n8398), .ZN(n5039) );
  NAND2_X4 U6293 ( .A1(n5487), .A2(n5040), .ZN(n8278) );
  NAND2_X2 U6294 ( .A1(n5484), .A2(n5486), .ZN(n5040) );
  NAND3_X1 U6295 ( .A1(n5040), .A2(n5487), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n5637) );
  NAND3_X1 U6296 ( .A1(n5040), .A2(n5487), .A3(n5641), .ZN(n5158) );
  NAND3_X1 U6297 ( .A1(n5040), .A2(n5487), .A3(P2_DATAO_REG_2__SCAN_IN), .ZN(
        n5301) );
  NAND3_X1 U6298 ( .A1(n5040), .A2(n5487), .A3(n5219), .ZN(n5217) );
  NAND3_X1 U6299 ( .A1(n5040), .A2(n5487), .A3(P2_DATAO_REG_5__SCAN_IN), .ZN(
        n5127) );
  NAND2_X1 U6300 ( .A1(n7786), .A2(n5041), .ZN(n7425) );
  NOR2_X1 U6301 ( .A1(n9288), .A2(n9521), .ZN(n7344) );
  NAND2_X1 U6302 ( .A1(n9260), .A2(n5551), .ZN(n6323) );
  NAND2_X1 U6303 ( .A1(n5042), .A2(n5044), .ZN(P1_U3214) );
  NAND2_X1 U6304 ( .A1(n6357), .A2(n9259), .ZN(n5042) );
  NAND2_X1 U6305 ( .A1(n5777), .A2(n5778), .ZN(n7257) );
  NAND2_X1 U6306 ( .A1(n5045), .A2(n5779), .ZN(n7258) );
  INV_X1 U6307 ( .A(n5777), .ZN(n5045) );
  OAI21_X1 U6308 ( .B1(n5777), .B2(n5047), .A(n5046), .ZN(n7291) );
  NAND2_X1 U6309 ( .A1(n5779), .A2(n7259), .ZN(n5046) );
  NAND2_X1 U6310 ( .A1(n6185), .A2(n6184), .ZN(n9243) );
  INV_X1 U6311 ( .A(n5048), .ZN(n9197) );
  INV_X1 U6312 ( .A(n6185), .ZN(n5404) );
  NAND4_X1 U6313 ( .A1(n5394), .A2(n5081), .A3(n5074), .A4(n7649), .ZN(n5071)
         );
  OAI21_X1 U6314 ( .B1(n5080), .B2(n5604), .A(n5076), .ZN(n6070) );
  NAND2_X1 U6315 ( .A1(n7383), .A2(n7384), .ZN(n7382) );
  OAI21_X1 U6316 ( .B1(n9269), .B2(n9272), .A(n9270), .ZN(n9205) );
  NOR2_X1 U6317 ( .A1(n6023), .A2(n6022), .ZN(n9269) );
  NAND2_X1 U6318 ( .A1(n6877), .A2(n6878), .ZN(n6876) );
  NAND2_X1 U6319 ( .A1(n7382), .A2(n4950), .ZN(n7648) );
  NAND2_X1 U6320 ( .A1(n7290), .A2(n5802), .ZN(n7383) );
  NAND2_X1 U6321 ( .A1(n5670), .A2(n6832), .ZN(n6877) );
  NAND2_X1 U6322 ( .A1(n7648), .A2(n7650), .ZN(n5081) );
  NAND2_X2 U6323 ( .A1(n7198), .A2(n5082), .ZN(n5633) );
  NAND2_X1 U6324 ( .A1(n7088), .A2(n5100), .ZN(n7087) );
  NAND2_X1 U6325 ( .A1(n5587), .A2(n6315), .ZN(n9533) );
  NAND2_X1 U6326 ( .A1(n9197), .A2(n9198), .ZN(n9196) );
  INV_X1 U6327 ( .A(n9533), .ZN(n6319) );
  NAND2_X1 U6328 ( .A1(n5409), .A2(n5408), .ZN(n9254) );
  NAND2_X1 U6329 ( .A1(n5851), .A2(n5850), .ZN(n7649) );
  NAND2_X1 U6330 ( .A1(n6831), .A2(n6833), .ZN(n5670) );
  NAND2_X1 U6331 ( .A1(n5666), .A2(n5667), .ZN(n6831) );
  NAND2_X1 U6332 ( .A1(n9231), .A2(n6123), .ZN(n9189) );
  INV_X1 U6333 ( .A(n7900), .ZN(n5085) );
  INV_X1 U6334 ( .A(n5609), .ZN(n9521) );
  NAND2_X1 U6335 ( .A1(n9188), .A2(n6151), .ZN(n6185) );
  NAND3_X1 U6337 ( .A1(n9595), .A2(n5088), .A3(n5027), .ZN(n5087) );
  NOR2_X1 U6338 ( .A1(n9592), .A2(n9591), .ZN(n9601) );
  NOR2_X1 U6339 ( .A1(n6730), .A2(n6729), .ZN(n6885) );
  NAND2_X1 U6340 ( .A1(n6708), .A2(n6707), .ZN(n6727) );
  NOR2_X1 U6341 ( .A1(n6662), .A2(n6661), .ZN(n6704) );
  NOR2_X1 U6342 ( .A1(n6888), .A2(n6887), .ZN(n7156) );
  NOR2_X1 U6343 ( .A1(n6790), .A2(n6789), .ZN(n6788) );
  NOR2_X1 U6344 ( .A1(n6955), .A2(n6954), .ZN(n6953) );
  NOR2_X1 U6345 ( .A1(n6642), .A2(n6641), .ZN(n6655) );
  NAND2_X1 U6346 ( .A1(n5634), .A2(n5629), .ZN(n6696) );
  NAND2_X1 U6347 ( .A1(n8688), .A2(n8687), .ZN(n8686) );
  NAND2_X2 U6348 ( .A1(n8589), .A2(n8590), .ZN(n8535) );
  NOR2_X1 U6349 ( .A1(n7011), .A2(n7010), .ZN(n7131) );
  NAND2_X1 U6350 ( .A1(n5221), .A2(n7781), .ZN(n7805) );
  NAND2_X1 U6351 ( .A1(n7422), .A2(n7421), .ZN(n7517) );
  NAND2_X1 U6352 ( .A1(n5222), .A2(n7552), .ZN(n7658) );
  NAND2_X1 U6353 ( .A1(n9732), .A2(n9643), .ZN(n5106) );
  NAND2_X1 U6354 ( .A1(n9671), .A2(n9679), .ZN(n9670) );
  NAND2_X1 U6355 ( .A1(n4948), .A2(n4996), .ZN(n5099) );
  NAND2_X1 U6356 ( .A1(n9637), .A2(n5536), .ZN(n9824) );
  NAND2_X1 U6357 ( .A1(n5788), .A2(n5770), .ZN(n7126) );
  OAI21_X2 U6358 ( .B1(n8909), .B2(n8455), .A(n8453), .ZN(n8894) );
  NAND2_X1 U6359 ( .A1(n5714), .A2(n5713), .ZN(n5728) );
  NAND2_X1 U6360 ( .A1(n8987), .A2(n8986), .ZN(n8231) );
  NAND2_X1 U6361 ( .A1(n8082), .A2(n8081), .ZN(n8080) );
  AOI22_X2 U6362 ( .A1(n8885), .A2(n8459), .B1(n8898), .B2(n9095), .ZN(n8877)
         );
  NAND2_X1 U6363 ( .A1(n7765), .A2(n7764), .ZN(n7840) );
  OAI22_X1 U6364 ( .A1(n8050), .A2(n8049), .B1(n8706), .B2(n8401), .ZN(n8051)
         );
  NAND2_X2 U6365 ( .A1(n8142), .A2(n8141), .ZN(n8929) );
  AND3_X2 U6366 ( .A1(n6744), .A2(n6745), .A3(n4983), .ZN(n10572) );
  AOI22_X1 U6367 ( .A1(n8866), .A2(n8203), .B1(n9022), .B2(n8879), .ZN(n8857)
         );
  OAI21_X1 U6368 ( .B1(n7468), .B2(n7467), .A(n7466), .ZN(n7469) );
  NOR2_X2 U6369 ( .A1(n10487), .A2(n10486), .ZN(n10504) );
  NAND2_X1 U6370 ( .A1(n7056), .A2(n7055), .ZN(n7057) );
  NAND2_X1 U6371 ( .A1(n7540), .A2(n7539), .ZN(n7541) );
  NAND2_X1 U6372 ( .A1(n8782), .A2(n10509), .ZN(n5331) );
  NAND2_X1 U6373 ( .A1(n7338), .A2(n9356), .ZN(n7337) );
  NAND2_X1 U6374 ( .A1(n9839), .A2(n5002), .ZN(n9637) );
  AOI22_X1 U6375 ( .A1(n9690), .A2(n9698), .B1(n9615), .B2(n9911), .ZN(n9671)
         );
  AOI21_X1 U6376 ( .B1(n9854), .B2(n9636), .A(n4999), .ZN(n9839) );
  NAND2_X1 U6377 ( .A1(n9189), .A2(n9190), .ZN(n9188) );
  NAND2_X1 U6378 ( .A1(n5817), .A2(n5547), .ZN(n5857) );
  NAND2_X1 U6379 ( .A1(n7103), .A2(n7104), .ZN(n7088) );
  NAND2_X1 U6380 ( .A1(n5636), .A2(n5635), .ZN(n5666) );
  AOI21_X1 U6381 ( .B1(n5524), .B2(n5526), .A(n5000), .ZN(n5522) );
  OAI21_X1 U6382 ( .B1(n7657), .B2(n5526), .A(n9418), .ZN(n5525) );
  AOI21_X1 U6383 ( .B1(n8495), .B2(n8494), .A(n8493), .ZN(n8498) );
  INV_X1 U6384 ( .A(n8486), .ZN(n5191) );
  NAND2_X1 U6385 ( .A1(n7045), .A2(n10158), .ZN(n8192) );
  NAND3_X1 U6386 ( .A1(n5170), .A2(n5169), .A3(n8477), .ZN(n8481) );
  NAND2_X1 U6387 ( .A1(n5104), .A2(n5637), .ZN(n5639) );
  NAND2_X1 U6388 ( .A1(n5640), .A2(n10221), .ZN(n5105) );
  INV_X1 U6389 ( .A(n5525), .ZN(n5524) );
  AOI21_X2 U6390 ( .B1(n5107), .B2(n4943), .A(n5224), .ZN(n9744) );
  NAND2_X1 U6391 ( .A1(n5274), .A2(n5272), .ZN(n8885) );
  OAI22_X1 U6392 ( .A1(n7274), .A2(n7234), .B1(n7277), .B2(n8713), .ZN(n7468)
         );
  INV_X1 U6393 ( .A(n7469), .ZN(n7470) );
  OAI21_X2 U6394 ( .B1(n8619), .B2(n8109), .A(n8975), .ZN(n8966) );
  NAND2_X1 U6395 ( .A1(n8894), .A2(n8460), .ZN(n5437) );
  NAND2_X1 U6396 ( .A1(n7780), .A2(n9370), .ZN(n5221) );
  NAND2_X1 U6397 ( .A1(n7551), .A2(n9400), .ZN(n5222) );
  NAND2_X1 U6398 ( .A1(n9912), .A2(n10711), .ZN(n5241) );
  NAND2_X1 U6399 ( .A1(n7445), .A2(n7444), .ZN(n7551) );
  NAND2_X1 U6400 ( .A1(n7707), .A2(n7706), .ZN(n7780) );
  OAI211_X1 U6401 ( .C1(n9907), .C2(n10528), .A(n9905), .B(n9906), .ZN(n10000)
         );
  NAND2_X1 U6402 ( .A1(n9163), .A2(n5998), .ZN(n6023) );
  NAND2_X2 U6403 ( .A1(n5879), .A2(n5878), .ZN(n5899) );
  INV_X1 U6404 ( .A(n5768), .ZN(n5110) );
  NAND2_X1 U6405 ( .A1(n5110), .A2(n5787), .ZN(n5109) );
  INV_X1 U6406 ( .A(n5787), .ZN(n5290) );
  INV_X1 U6407 ( .A(n9500), .ZN(n5111) );
  OAI21_X1 U6408 ( .B1(n5111), .B2(n5114), .A(n5003), .ZN(n9503) );
  NAND3_X1 U6409 ( .A1(n5125), .A2(n9509), .A3(n5124), .ZN(n5123) );
  OAI211_X1 U6410 ( .C1(n5487), .C2(n6473), .A(n5128), .B(n5127), .ZN(n5766)
         );
  NAND2_X2 U6411 ( .A1(n5485), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5487) );
  INV_X1 U6412 ( .A(n9477), .ZN(n5153) );
  AOI21_X2 U6413 ( .B1(n9668), .B2(n9852), .A(n5157), .ZN(n9906) );
  OAI211_X1 U6414 ( .C1(n5487), .C2(P1_DATAO_REG_0__SCAN_IN), .A(n5159), .B(
        n5158), .ZN(n5643) );
  NAND2_X1 U6415 ( .A1(n5129), .A2(n5642), .ZN(n5159) );
  NAND2_X1 U6416 ( .A1(n5160), .A2(n8356), .ZN(n8364) );
  NAND2_X1 U6417 ( .A1(n8355), .A2(n5161), .ZN(n5160) );
  OAI21_X1 U6418 ( .B1(n8348), .B2(n8491), .A(n4965), .ZN(n5161) );
  NAND2_X1 U6419 ( .A1(n4976), .A2(n8491), .ZN(n5162) );
  NAND2_X1 U6420 ( .A1(n5165), .A2(n5168), .ZN(n5163) );
  AND2_X1 U6421 ( .A1(n8986), .A2(n5269), .ZN(n5167) );
  NAND2_X1 U6422 ( .A1(n8416), .A2(n8415), .ZN(n5168) );
  NAND3_X1 U6423 ( .A1(n8463), .A2(n8856), .A3(n5171), .ZN(n5169) );
  INV_X1 U6424 ( .A(n5182), .ZN(n7325) );
  NAND2_X1 U6425 ( .A1(n7172), .A2(n7177), .ZN(n5183) );
  NAND3_X1 U6426 ( .A1(n5191), .A2(n8485), .A3(n8247), .ZN(n8495) );
  XNOR2_X2 U6427 ( .A(n5192), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6934) );
  NOR2_X1 U6428 ( .A1(n6395), .A2(n9147), .ZN(n5192) );
  NAND3_X1 U6429 ( .A1(n5196), .A2(n8491), .A3(n8398), .ZN(n5195) );
  NAND2_X1 U6430 ( .A1(n6997), .A2(n6943), .ZN(n8346) );
  NAND2_X1 U6431 ( .A1(n7078), .A2(n6942), .ZN(n8342) );
  NAND3_X1 U6432 ( .A1(n8342), .A2(n8345), .A3(n8346), .ZN(n7074) );
  OR2_X2 U6433 ( .A1(n7718), .A2(n10662), .ZN(n7719) );
  NOR2_X2 U6434 ( .A1(n7450), .A2(n7456), .ZN(n7562) );
  INV_X1 U6435 ( .A(n5206), .ZN(n7970) );
  NAND2_X1 U6436 ( .A1(n5765), .A2(n5216), .ZN(n7006) );
  OR2_X1 U6437 ( .A1(n5734), .A2(n5733), .ZN(n5216) );
  INV_X2 U6438 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5573) );
  NAND2_X1 U6439 ( .A1(n7208), .A2(n5253), .ZN(n9304) );
  XNOR2_X1 U6440 ( .A(n5255), .B(n9356), .ZN(n7348) );
  INV_X1 U6441 ( .A(n9699), .ZN(n5257) );
  NAND2_X1 U6442 ( .A1(n4984), .A2(n5256), .ZN(n9684) );
  NAND2_X1 U6443 ( .A1(n9701), .A2(n9661), .ZN(n9680) );
  NAND3_X1 U6444 ( .A1(n5548), .A2(n5957), .A3(n5614), .ZN(n5616) );
  NAND2_X1 U6445 ( .A1(n8052), .A2(n4933), .ZN(n5266) );
  NAND2_X1 U6446 ( .A1(n5266), .A2(n5267), .ZN(n8977) );
  NAND2_X1 U6447 ( .A1(n8929), .A2(n5275), .ZN(n5274) );
  NAND2_X1 U6448 ( .A1(n5769), .A2(n5289), .ZN(n5288) );
  NAND2_X1 U6449 ( .A1(n8966), .A2(n5293), .ZN(n5291) );
  NAND2_X1 U6450 ( .A1(n5291), .A2(n5292), .ZN(n8142) );
  NAND2_X1 U6451 ( .A1(n9013), .A2(n9012), .ZN(n9071) );
  OAI21_X2 U6452 ( .B1(n7939), .B2(n4974), .A(n7940), .ZN(n8050) );
  NAND3_X1 U6453 ( .A1(n5484), .A2(n5486), .A3(P1_DATAO_REG_2__SCAN_IN), .ZN(
        n5302) );
  NAND2_X1 U6454 ( .A1(n7182), .A2(n5314), .ZN(n5312) );
  OAI21_X1 U6455 ( .B1(n7182), .B2(n4934), .A(n5314), .ZN(n7408) );
  NAND2_X1 U6456 ( .A1(n7327), .A2(n5316), .ZN(n5317) );
  NAND2_X1 U6457 ( .A1(n7182), .A2(n7183), .ZN(n7327) );
  INV_X1 U6458 ( .A(n7393), .ZN(n5318) );
  NAND3_X1 U6459 ( .A1(n5322), .A2(n5319), .A3(P2_REG2_REG_3__SCAN_IN), .ZN(
        n6926) );
  NAND2_X1 U6460 ( .A1(n6685), .A2(n5320), .ZN(n5319) );
  NAND2_X1 U6461 ( .A1(n6926), .A2(n5322), .ZN(n6927) );
  NOR2_X1 U6462 ( .A1(n10450), .A2(n10451), .ZN(n10449) );
  NOR2_X1 U6463 ( .A1(n10400), .A2(n10399), .ZN(n10398) );
  NOR2_X1 U6464 ( .A1(n10434), .A2(n10433), .ZN(n10432) );
  OAI22_X1 U6465 ( .A1(n8857), .A2(n8856), .B1(n9080), .B2(n8554), .ZN(n8845)
         );
  OAI21_X1 U6466 ( .B1(n8849), .B2(n10562), .A(n8848), .ZN(n9014) );
  NAND2_X1 U6467 ( .A1(n7715), .A2(n7716), .ZN(n7798) );
  NAND2_X1 U6468 ( .A1(n7912), .A2(n7911), .ZN(n7960) );
  NAND2_X2 U6469 ( .A1(n8014), .A2(n9460), .ZN(n9341) );
  NOR2_X1 U6470 ( .A1(n8732), .A2(n8733), .ZN(n8767) );
  XNOR2_X2 U6471 ( .A(n6393), .B(n6392), .ZN(n6612) );
  NAND2_X1 U6472 ( .A1(n5831), .A2(n5830), .ZN(n5856) );
  NAND2_X1 U6473 ( .A1(n5335), .A2(n7989), .ZN(n5333) );
  INV_X1 U6474 ( .A(n6751), .ZN(n5340) );
  NAND2_X1 U6475 ( .A1(n5339), .A2(n6747), .ZN(n5341) );
  NAND2_X1 U6476 ( .A1(n5337), .A2(n5336), .ZN(n6863) );
  NAND2_X1 U6477 ( .A1(n6856), .A2(n6751), .ZN(n5336) );
  NAND2_X1 U6478 ( .A1(n5339), .A2(n5338), .ZN(n5337) );
  INV_X1 U6479 ( .A(n6749), .ZN(n5339) );
  INV_X1 U6480 ( .A(n5341), .ZN(n6750) );
  NOR2_X1 U6481 ( .A1(n6598), .A2(n6599), .ZN(n6749) );
  NAND2_X1 U6482 ( .A1(n5342), .A2(n5343), .ZN(n7890) );
  INV_X1 U6483 ( .A(n6416), .ZN(n5355) );
  NAND2_X1 U6484 ( .A1(n5355), .A2(n5363), .ZN(n6384) );
  INV_X1 U6485 ( .A(n6384), .ZN(n5356) );
  AND2_X1 U6486 ( .A1(n5360), .A2(n5001), .ZN(n6377) );
  AND4_X1 U6487 ( .A1(n5440), .A2(n6367), .A3(n6368), .A4(n6395), .ZN(n7268)
         );
  INV_X1 U6488 ( .A(n8512), .ZN(n5372) );
  NAND2_X1 U6489 ( .A1(n8535), .A2(n5378), .ZN(n8657) );
  NAND2_X1 U6490 ( .A1(n8549), .A2(n5381), .ZN(n5380) );
  OAI211_X1 U6491 ( .C1(n8549), .C2(n5382), .A(n5380), .B(n8558), .ZN(P2_U3160) );
  NAND2_X1 U6492 ( .A1(n8549), .A2(n8548), .ZN(n8560) );
  NAND2_X1 U6493 ( .A1(n9205), .A2(n4938), .ZN(n5409) );
  INV_X1 U6494 ( .A(n5410), .ZN(n9204) );
  NAND2_X1 U6495 ( .A1(n7382), .A2(n5829), .ZN(n5851) );
  NAND2_X1 U6496 ( .A1(n7900), .A2(n5413), .ZN(n5412) );
  NAND4_X1 U6497 ( .A1(n5555), .A2(n5556), .A3(n5557), .A4(n5558), .ZN(n5762)
         );
  NAND3_X1 U6498 ( .A1(n5555), .A2(n5556), .A3(n5557), .ZN(n5724) );
  INV_X1 U6499 ( .A(n5603), .ZN(n6298) );
  XNOR2_X1 U6500 ( .A(n5417), .B(n5562), .ZN(n5603) );
  NAND2_X1 U6501 ( .A1(n5584), .A2(n5583), .ZN(n5602) );
  OAI211_X1 U6502 ( .C1(n8335), .C2(n5424), .A(n5423), .B(n5422), .ZN(P2_U3296) );
  NAND3_X1 U6503 ( .A1(n8335), .A2(n5029), .A3(n5429), .ZN(n5422) );
  NAND2_X1 U6504 ( .A1(n5439), .A2(n5438), .ZN(n7926) );
  NAND4_X1 U6505 ( .A1(n6368), .A2(n6367), .A3(n6395), .A4(n6369), .ZN(n6900)
         );
  NAND3_X1 U6506 ( .A1(n6368), .A2(n6395), .A3(n6367), .ZN(n6795) );
  NAND2_X1 U6507 ( .A1(n8865), .A2(n5447), .ZN(n5445) );
  NAND2_X1 U6508 ( .A1(n5445), .A2(n5446), .ZN(n8302) );
  INV_X1 U6509 ( .A(n5450), .ZN(n8298) );
  NOR2_X2 U6510 ( .A1(n6373), .A2(n5451), .ZN(n6522) );
  INV_X1 U6511 ( .A(n5687), .ZN(n5456) );
  NAND2_X1 U6512 ( .A1(n6158), .A2(n6157), .ZN(n6168) );
  NAND2_X1 U6513 ( .A1(n6233), .A2(n5470), .ZN(n5468) );
  NAND2_X1 U6514 ( .A1(n6233), .A2(n6232), .ZN(n6257) );
  NAND2_X1 U6515 ( .A1(n5815), .A2(n5814), .ZN(n5831) );
  NAND2_X1 U6516 ( .A1(n6062), .A2(n4939), .ZN(n5489) );
  NAND2_X1 U6517 ( .A1(n6062), .A2(n6061), .ZN(n5494) );
  INV_X1 U6518 ( .A(n6001), .ZN(n5508) );
  NAND2_X1 U6519 ( .A1(n6001), .A2(n5502), .ZN(n5500) );
  NAND2_X1 U6520 ( .A1(n5899), .A2(n5516), .ZN(n5513) );
  NAND2_X1 U6521 ( .A1(n5899), .A2(n5898), .ZN(n5923) );
  OAI211_X1 U6522 ( .C1(n6742), .C2(n5726), .A(n5519), .B(n5518), .ZN(n6879)
         );
  NAND2_X1 U6523 ( .A1(n5520), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5519) );
  INV_X2 U6524 ( .A(n5735), .ZN(n5520) );
  NAND2_X2 U6525 ( .A1(n5648), .A2(n6594), .ZN(n5726) );
  NAND2_X1 U6526 ( .A1(n5521), .A2(n5522), .ZN(n7705) );
  AOI21_X2 U6527 ( .B1(n5534), .B2(n5530), .A(n5528), .ZN(n8016) );
  NOR2_X1 U6528 ( .A1(n5535), .A2(n5604), .ZN(n5722) );
  OAI21_X1 U6529 ( .B1(n9907), .B2(n5544), .A(n5538), .ZN(P1_U3519) );
  AND2_X2 U6530 ( .A1(n5817), .A2(n5546), .ZN(n5928) );
  NAND2_X1 U6531 ( .A1(n5957), .A2(n5566), .ZN(n5596) );
  XNOR2_X1 U6532 ( .A(n6855), .B(n7081), .ZN(n6751) );
  NAND2_X1 U6533 ( .A1(n6855), .A2(n7081), .ZN(n6856) );
  XNOR2_X1 U6534 ( .A(n6610), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10388) );
  INV_X1 U6535 ( .A(n8303), .ZN(n9070) );
  INV_X1 U6536 ( .A(n6526), .ZN(n9153) );
  XNOR2_X1 U6537 ( .A(n8845), .B(n8844), .ZN(n8849) );
  CLKBUF_X1 U6538 ( .A(n8596), .Z(n8597) );
  NAND2_X1 U6539 ( .A1(n8287), .A2(n8277), .ZN(n8282) );
  XNOR2_X1 U6540 ( .A(n7072), .B(n6861), .ZN(n6855) );
  NAND2_X1 U6541 ( .A1(n6946), .A2(n6947), .ZN(n10558) );
  NAND2_X1 U6542 ( .A1(n6153), .A2(n6152), .ZN(n6158) );
  INV_X1 U6543 ( .A(n9628), .ZN(n9999) );
  INV_X1 U6544 ( .A(n5666), .ZN(n5669) );
  INV_X1 U6545 ( .A(n5639), .ZN(n5640) );
  NAND2_X1 U6546 ( .A1(n8500), .A2(n7691), .ZN(n8501) );
  XNOR2_X1 U6547 ( .A(n8268), .B(n8226), .ZN(n9289) );
  NAND2_X1 U6548 ( .A1(n5648), .A2(n10288), .ZN(n5575) );
  XNOR2_X1 U6549 ( .A(n6276), .B(n6275), .ZN(n8265) );
  INV_X1 U6550 ( .A(n5620), .ZN(n10052) );
  OR2_X1 U6551 ( .A1(n9213), .A2(n6059), .ZN(n5550) );
  NAND2_X2 U6552 ( .A1(n7343), .A2(n10522), .ZN(n10525) );
  AND2_X1 U6553 ( .A1(n6330), .A2(n6343), .ZN(n9259) );
  AND2_X1 U6554 ( .A1(n6355), .A2(n6356), .ZN(n5551) );
  INV_X1 U6555 ( .A(n8994), .ZN(n10564) );
  INV_X1 U6556 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6981) );
  AND2_X1 U6557 ( .A1(n6321), .A2(n9259), .ZN(n5552) );
  INV_X1 U6558 ( .A(n9242), .ZN(n9281) );
  INV_X1 U6559 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6979) );
  INV_X1 U6560 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6866) );
  INV_X1 U6561 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6985) );
  INV_X1 U6562 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6975) );
  INV_X1 U6563 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6977) );
  INV_X1 U6564 ( .A(n9171), .ZN(n7969) );
  NAND2_X2 U6565 ( .A1(n6824), .A2(n10570), .ZN(n10577) );
  NAND2_X1 U6566 ( .A1(n8484), .A2(n8483), .ZN(n8485) );
  INV_X1 U6567 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5564) );
  INV_X1 U6568 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6408) );
  INV_X1 U6569 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5561) );
  OR2_X1 U6570 ( .A1(n6150), .A2(n6149), .ZN(n6151) );
  INV_X1 U6571 ( .A(n8707), .ZN(n8067) );
  INV_X1 U6572 ( .A(n8710), .ZN(n7731) );
  AOI211_X1 U6573 ( .C1(n9067), .C2(n8303), .A(n8496), .B(n8302), .ZN(n8305)
         );
  INV_X1 U6574 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6412) );
  INV_X1 U6575 ( .A(n5850), .ZN(n5848) );
  INV_X1 U6576 ( .A(n9693), .ZN(n9615) );
  INV_X1 U6577 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5568) );
  INV_X1 U6578 ( .A(SI_26_), .ZN(n10170) );
  INV_X1 U6579 ( .A(SI_22_), .ZN(n10180) );
  INV_X1 U6580 ( .A(SI_16_), .ZN(n10195) );
  INV_X1 U6581 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5557) );
  AND2_X1 U6582 ( .A1(n7361), .A2(n8712), .ZN(n7362) );
  INV_X1 U6583 ( .A(n7001), .ZN(n7002) );
  NAND2_X1 U6584 ( .A1(n8533), .A2(n8932), .ZN(n8534) );
  INV_X1 U6585 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6983) );
  NOR2_X1 U6586 ( .A1(n8171), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n7045) );
  OR2_X1 U6587 ( .A1(n6547), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6533) );
  INV_X1 U6588 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6519) );
  NAND2_X1 U6589 ( .A1(n5695), .A2(n5694), .ZN(n5698) );
  AND2_X1 U6590 ( .A1(n6139), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6162) );
  NOR2_X1 U6591 ( .A1(n6194), .A2(n9226), .ZN(n6224) );
  INV_X1 U6592 ( .A(n9522), .ZN(n9526) );
  INV_X1 U6593 ( .A(n9340), .ZN(n7197) );
  INV_X1 U6594 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10046) );
  INV_X1 U6595 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5589) );
  OR2_X1 U6596 ( .A1(n6006), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6007) );
  NOR2_X1 U6597 ( .A1(n7363), .A2(n7362), .ZN(n7369) );
  OR2_X1 U6598 ( .A1(n7588), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7767) );
  OR2_X1 U6599 ( .A1(n8208), .A2(n8189), .ZN(n8190) );
  NAND2_X1 U6600 ( .A1(n7002), .A2(n8715), .ZN(n7003) );
  OR2_X1 U6601 ( .A1(n8169), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8171) );
  OAI21_X1 U6602 ( .B1(n7311), .B2(n8713), .A(n7310), .ZN(n7312) );
  NAND2_X1 U6603 ( .A1(n6984), .A2(n6983), .ZN(n8096) );
  AND2_X1 U6604 ( .A1(n8296), .A2(n7305), .ZN(n8846) );
  NAND2_X1 U6605 ( .A1(n7146), .A2(n7145), .ZN(n8211) );
  NAND2_X1 U6606 ( .A1(n6986), .A2(n6985), .ZN(n8122) );
  NAND2_X1 U6607 ( .A1(n6533), .A2(n6532), .ZN(n6819) );
  AND2_X1 U6608 ( .A1(n6535), .A2(n6810), .ZN(n6808) );
  NAND2_X1 U6609 ( .A1(n6494), .A2(n6566), .ZN(n6577) );
  INV_X1 U6610 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6456) );
  INV_X1 U6611 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9147) );
  AND3_X1 U6612 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5780) );
  NOR2_X1 U6613 ( .A1(n6106), .A2(n9236), .ZN(n6139) );
  AND2_X1 U6614 ( .A1(n9261), .A2(n9262), .ZN(n6252) );
  AND2_X1 U6615 ( .A1(n5608), .A2(n7744), .ZN(n9340) );
  AND2_X1 U6616 ( .A1(n6162), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6171) );
  INV_X1 U6617 ( .A(n9691), .ZN(n9721) );
  INV_X1 U6618 ( .A(n9758), .ZN(n9729) );
  INV_X1 U6619 ( .A(n9553), .ZN(n9949) );
  INV_X1 U6620 ( .A(n9631), .ZN(n9879) );
  INV_X1 U6621 ( .A(n9451), .ZN(n7961) );
  INV_X1 U6622 ( .A(n9677), .ZN(n9861) );
  OR2_X1 U6623 ( .A1(n10042), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6303) );
  OR2_X1 U6624 ( .A1(n9620), .A2(n9619), .ZN(n9898) );
  OR2_X1 U6625 ( .A1(n9296), .A2(n7985), .ZN(n6221) );
  OR2_X1 U6626 ( .A1(n9296), .A2(n7746), .ZN(n6104) );
  OR2_X1 U6627 ( .A1(n10518), .A2(n7201), .ZN(n7786) );
  NAND2_X1 U6628 ( .A1(n9526), .A2(n10347), .ZN(n10631) );
  NAND2_X1 U6629 ( .A1(n10532), .A2(n7197), .ZN(n10729) );
  INV_X1 U6630 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5576) );
  INV_X1 U6631 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5590) );
  AND2_X1 U6632 ( .A1(n6604), .A2(n6948), .ZN(n8676) );
  AND2_X1 U6633 ( .A1(n8218), .A2(n8217), .ZN(n8237) );
  INV_X1 U6634 ( .A(n8183), .ZN(n8215) );
  OR2_X1 U6635 ( .A1(n6513), .A2(n8825), .ZN(n10489) );
  INV_X1 U6636 ( .A(n8830), .ZN(n10513) );
  OR2_X1 U6637 ( .A1(n10715), .A2(n6554), .ZN(n10571) );
  AND2_X1 U6638 ( .A1(n6948), .A2(n8492), .ZN(n8994) );
  INV_X1 U6639 ( .A(n8937), .ZN(n9001) );
  OR2_X1 U6640 ( .A1(n6577), .A2(n6809), .ZN(n10570) );
  INV_X1 U6641 ( .A(n9050), .ZN(n9061) );
  NOR2_X1 U6642 ( .A1(n6808), .A2(n6807), .ZN(n6822) );
  INV_X1 U6643 ( .A(n8856), .ZN(n8854) );
  OR2_X1 U6644 ( .A1(n8308), .A2(n4988), .ZN(n8908) );
  NAND2_X1 U6645 ( .A1(n8256), .A2(n10689), .ZN(n10720) );
  INV_X1 U6646 ( .A(n8267), .ZN(n7817) );
  AND2_X1 U6647 ( .A1(n6324), .A2(n9259), .ZN(n6320) );
  INV_X1 U6648 ( .A(n9276), .ZN(n8011) );
  INV_X1 U6649 ( .A(n10366), .ZN(n9590) );
  INV_X1 U6650 ( .A(n10362), .ZN(n9582) );
  NOR2_X1 U6651 ( .A1(n10353), .A2(n10347), .ZN(n9609) );
  INV_X1 U6652 ( .A(n9826), .ZN(n9884) );
  INV_X1 U6653 ( .A(n10631), .ZN(n10704) );
  AND2_X1 U6654 ( .A1(n10525), .A2(n5608), .ZN(n9891) );
  INV_X1 U6655 ( .A(n9880), .ZN(n10519) );
  AND2_X1 U6656 ( .A1(n6303), .A2(n10045), .ZN(n7224) );
  INV_X1 U6657 ( .A(n10528), .ZN(n10711) );
  AND2_X1 U6658 ( .A1(n9533), .A2(n9521), .ZN(n10532) );
  NAND2_X1 U6659 ( .A1(n6132), .A2(n6131), .ZN(n6153) );
  INV_X1 U6660 ( .A(n8249), .ZN(n8131) );
  INV_X1 U6661 ( .A(n8694), .ZN(n7381) );
  INV_X1 U6662 ( .A(n8237), .ZN(n8858) );
  INV_X1 U6663 ( .A(n8619), .ZN(n8996) );
  OR2_X1 U6664 ( .A1(n6494), .A2(n6560), .ZN(n10503) );
  OR2_X1 U6665 ( .A1(n6513), .A2(n6572), .ZN(n10496) );
  NAND2_X1 U6666 ( .A1(n10577), .A2(n10576), .ZN(n9004) );
  NAND2_X1 U6667 ( .A1(n10723), .A2(n10720), .ZN(n9064) );
  AND2_X2 U6668 ( .A1(n6822), .A2(n6815), .ZN(n10723) );
  INV_X1 U6669 ( .A(n8642), .ZN(n9115) );
  NAND2_X1 U6670 ( .A1(n10727), .A2(n10720), .ZN(n9145) );
  AND3_X1 U6671 ( .A1(n10675), .A2(n10674), .A3(n10673), .ZN(n10678) );
  INV_X1 U6672 ( .A(n10727), .ZN(n10724) );
  INV_X1 U6673 ( .A(n6560), .ZN(n6566) );
  NAND2_X1 U6674 ( .A1(n6847), .A2(n6547), .ZN(n6433) );
  INV_X1 U6675 ( .A(n8505), .ZN(n7758) );
  NAND2_X1 U6676 ( .A1(n6358), .A2(n6320), .ZN(n6354) );
  NAND2_X1 U6677 ( .A1(n7261), .A2(n10705), .ZN(n9242) );
  INV_X1 U6678 ( .A(n9259), .ZN(n9284) );
  OR2_X1 U6679 ( .A1(n6144), .A2(n6143), .ZN(n9809) );
  INV_X2 U6680 ( .A(P1_U3973), .ZN(n9561) );
  OR2_X1 U6681 ( .A1(n6637), .A2(n6636), .ZN(n10353) );
  INV_X1 U6682 ( .A(n9609), .ZN(n10360) );
  NAND2_X1 U6683 ( .A1(n10525), .A2(n7425), .ZN(n9894) );
  INV_X1 U6684 ( .A(n10525), .ZN(n9685) );
  NAND2_X1 U6685 ( .A1(n10736), .A2(n10705), .ZN(n9991) );
  INV_X1 U6686 ( .A(n10736), .ZN(n10735) );
  NAND2_X1 U6687 ( .A1(n10740), .A2(n10705), .ZN(n10040) );
  INV_X1 U6688 ( .A(n10740), .ZN(n10737) );
  INV_X1 U6689 ( .A(n10053), .ZN(n10284) );
  INV_X1 U6690 ( .A(n10503), .ZN(P2_U3893) );
  NAND4_X1 U6691 ( .A1(n5583), .A2(n5563), .A3(n5600), .A4(n5562), .ZN(n5565)
         );
  NOR2_X1 U6692 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n5613) );
  INV_X1 U6693 ( .A(n5613), .ZN(n5567) );
  NOR2_X1 U6694 ( .A1(n8278), .A2(n10105), .ZN(n5574) );
  INV_X1 U6695 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5641) );
  XNOR2_X1 U6696 ( .A(n5574), .B(n5641), .ZN(n10288) );
  INV_X1 U6697 ( .A(n10533), .ZN(n5611) );
  NOR2_X1 U6698 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5580) );
  NOR2_X1 U6699 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5579) );
  NOR2_X1 U6700 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5578) );
  NOR2_X1 U6701 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5577) );
  NAND4_X1 U6702 ( .A1(n5580), .A2(n5579), .A3(n5578), .A4(n5577), .ZN(n5581)
         );
  INV_X1 U6703 ( .A(n5588), .ZN(n5584) );
  NAND2_X1 U6704 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n5585) );
  NAND2_X1 U6705 ( .A1(n5586), .A2(n5600), .ZN(n6315) );
  NAND2_X1 U6706 ( .A1(n6070), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U6707 ( .A1(n5609), .A2(n7744), .ZN(n5626) );
  NAND2_X1 U6708 ( .A1(n5596), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5597) );
  MUX2_X1 U6709 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5597), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5599) );
  INV_X1 U6710 ( .A(n5605), .ZN(n5598) );
  NAND2_X1 U6711 ( .A1(n4996), .A2(n5600), .ZN(n5601) );
  NOR2_X1 U6712 ( .A1(n6299), .A2(n5603), .ZN(n5607) );
  INV_X1 U6713 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U6714 ( .A1(n9533), .A2(n9340), .ZN(n5610) );
  INV_X1 U6715 ( .A(n5608), .ZN(n9610) );
  NAND2_X1 U6716 ( .A1(n9610), .A2(n7744), .ZN(n9288) );
  AND2_X1 U6717 ( .A1(n5613), .A2(n5612), .ZN(n5614) );
  NAND2_X1 U6718 ( .A1(n5616), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5618) );
  INV_X1 U6719 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5619) );
  INV_X1 U6720 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10521) );
  NAND2_X1 U6721 ( .A1(n5671), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5623) );
  INV_X1 U6722 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10534) );
  INV_X1 U6723 ( .A(n5626), .ZN(n6328) );
  NAND2_X1 U6724 ( .A1(n6474), .A2(n6074), .ZN(n5627) );
  INV_X1 U6725 ( .A(n6363), .ZN(n6439) );
  NAND2_X1 U6726 ( .A1(n6439), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U6727 ( .A1(n6474), .A2(n6247), .ZN(n5632) );
  NOR2_X1 U6728 ( .A1(n6363), .A2(n5576), .ZN(n5630) );
  AOI21_X1 U6729 ( .B1(n10533), .B2(n6074), .A(n5630), .ZN(n5631) );
  NAND2_X1 U6730 ( .A1(n5632), .A2(n5631), .ZN(n6695) );
  NAND2_X1 U6731 ( .A1(n6696), .A2(n6695), .ZN(n5636) );
  NAND2_X1 U6732 ( .A1(n5634), .A2(n5662), .ZN(n5635) );
  INV_X1 U6733 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U6734 ( .A1(n5639), .A2(SI_1_), .ZN(n5682) );
  INV_X1 U6735 ( .A(SI_1_), .ZN(n10221) );
  INV_X1 U6736 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5642) );
  INV_X1 U6737 ( .A(n5644), .ZN(n5645) );
  NAND2_X1 U6738 ( .A1(n5646), .A2(n5645), .ZN(n5647) );
  NAND2_X1 U6739 ( .A1(n5683), .A2(n5647), .ZN(n6593) );
  NAND2_X1 U6740 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5649) );
  OAI22_X1 U6741 ( .A1(n5726), .A2(n6593), .B1(n5648), .B2(n6725), .ZN(n5650)
         );
  INV_X1 U6742 ( .A(n5650), .ZN(n5651) );
  NAND2_X1 U6743 ( .A1(n7496), .A2(n5653), .ZN(n5661) );
  NAND2_X1 U6744 ( .A1(n5671), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5659) );
  INV_X1 U6745 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n5654) );
  INV_X1 U6746 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U6747 ( .A1(n5664), .A2(n6074), .ZN(n5660) );
  NAND2_X1 U6748 ( .A1(n5661), .A2(n5660), .ZN(n5663) );
  AND2_X1 U6749 ( .A1(n7496), .A2(n6074), .ZN(n5665) );
  AOI21_X1 U6750 ( .B1(n5664), .B2(n6247), .A(n5665), .ZN(n6833) );
  INV_X1 U6751 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7351) );
  NAND2_X1 U6752 ( .A1(n5671), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5675) );
  INV_X1 U6753 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5672) );
  NAND2_X1 U6754 ( .A1(n5692), .A2(n6074), .ZN(n5690) );
  INV_X1 U6755 ( .A(n5679), .ZN(n5677) );
  NAND2_X1 U6756 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5677), .ZN(n5678) );
  INV_X1 U6757 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5680) );
  MUX2_X1 U6758 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5678), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n5681) );
  NAND2_X1 U6759 ( .A1(n5680), .A2(n5679), .ZN(n5705) );
  INV_X1 U6760 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6400) );
  NAND2_X1 U6761 ( .A1(n5684), .A2(SI_2_), .ZN(n5707) );
  INV_X1 U6762 ( .A(n5685), .ZN(n5686) );
  NAND2_X1 U6763 ( .A1(n5687), .A2(n5686), .ZN(n5708) );
  NAND2_X1 U6764 ( .A1(n5688), .A2(n5708), .ZN(n6742) );
  NAND2_X1 U6765 ( .A1(n6879), .A2(n5653), .ZN(n5689) );
  NAND2_X1 U6766 ( .A1(n5690), .A2(n5689), .ZN(n5691) );
  XNOR2_X1 U6767 ( .A(n5691), .B(n5662), .ZN(n5697) );
  INV_X1 U6768 ( .A(n5697), .ZN(n5695) );
  AND2_X1 U6769 ( .A1(n6879), .A2(n6074), .ZN(n5693) );
  AOI21_X1 U6770 ( .B1(n5692), .B2(n6247), .A(n5693), .ZN(n5696) );
  INV_X1 U6771 ( .A(n5696), .ZN(n5694) );
  NAND2_X1 U6772 ( .A1(n5697), .A2(n5696), .ZN(n5699) );
  NAND2_X1 U6773 ( .A1(n6876), .A2(n5699), .ZN(n7103) );
  NAND2_X1 U6774 ( .A1(n5671), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5704) );
  OR2_X1 U6775 ( .A1(n5751), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5703) );
  INV_X1 U6776 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5700) );
  OR2_X1 U6777 ( .A1(n5755), .A2(n5700), .ZN(n5702) );
  INV_X1 U6778 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6643) );
  OR2_X1 U6779 ( .A1(n5753), .A2(n6643), .ZN(n5701) );
  NAND4_X1 U6780 ( .A1(n5704), .A2(n5703), .A3(n5702), .A4(n5701), .ZN(n10598)
         );
  NAND2_X1 U6781 ( .A1(n10598), .A2(n6074), .ZN(n5719) );
  NAND2_X1 U6782 ( .A1(n5705), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5706) );
  XNOR2_X1 U6783 ( .A(n5706), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6771) );
  INV_X1 U6784 ( .A(n6771), .ZN(n6401) );
  OR2_X1 U6785 ( .A1(n5735), .A2(n5219), .ZN(n5717) );
  NAND2_X1 U6786 ( .A1(n5708), .A2(n5707), .ZN(n5714) );
  NAND2_X1 U6787 ( .A1(n5709), .A2(SI_3_), .ZN(n5727) );
  INV_X1 U6788 ( .A(SI_3_), .ZN(n5710) );
  NAND2_X1 U6789 ( .A1(n5711), .A2(n5710), .ZN(n5712) );
  AND2_X1 U6790 ( .A1(n5727), .A2(n5712), .ZN(n5713) );
  OR2_X1 U6791 ( .A1(n5714), .A2(n5713), .ZN(n5715) );
  NAND2_X1 U6792 ( .A1(n5728), .A2(n5715), .ZN(n6858) );
  OR2_X1 U6793 ( .A1(n5726), .A2(n6858), .ZN(n5716) );
  NAND2_X1 U6794 ( .A1(n7214), .A2(n5653), .ZN(n5718) );
  NAND2_X1 U6795 ( .A1(n5719), .A2(n5718), .ZN(n5720) );
  AND2_X1 U6796 ( .A1(n7214), .A2(n6074), .ZN(n5721) );
  AOI21_X1 U6797 ( .B1(n10598), .B2(n6247), .A(n5721), .ZN(n5745) );
  MUX2_X1 U6798 ( .A(n5604), .B(n5722), .S(P1_IR_REG_4__SCAN_IN), .Z(n5723) );
  INV_X1 U6799 ( .A(n5723), .ZN(n5725) );
  NAND2_X1 U6800 ( .A1(n5725), .A2(n5724), .ZN(n6918) );
  NAND2_X1 U6801 ( .A1(n5728), .A2(n5727), .ZN(n5734) );
  MUX2_X1 U6802 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n6594), .Z(n5729) );
  NAND2_X1 U6803 ( .A1(n5729), .A2(SI_4_), .ZN(n5764) );
  INV_X1 U6804 ( .A(n5729), .ZN(n5731) );
  INV_X1 U6805 ( .A(SI_4_), .ZN(n5730) );
  NAND2_X1 U6806 ( .A1(n5731), .A2(n5730), .ZN(n5732) );
  AND2_X1 U6807 ( .A1(n5764), .A2(n5732), .ZN(n5733) );
  INV_X1 U6808 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6398) );
  NAND2_X1 U6809 ( .A1(n10597), .A2(n5653), .ZN(n5741) );
  NAND2_X1 U6810 ( .A1(n6283), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5739) );
  INV_X1 U6811 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6633) );
  OR2_X1 U6812 ( .A1(n5755), .A2(n6633), .ZN(n5738) );
  XNOR2_X1 U6813 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7518) );
  OR2_X1 U6814 ( .A1(n5751), .A2(n7518), .ZN(n5737) );
  INV_X1 U6815 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6646) );
  OR2_X1 U6816 ( .A1(n5753), .A2(n6646), .ZN(n5736) );
  NAND4_X1 U6817 ( .A1(n5739), .A2(n5738), .A3(n5737), .A4(n5736), .ZN(n9560)
         );
  NAND2_X1 U6818 ( .A1(n9560), .A2(n6074), .ZN(n5740) );
  NAND2_X1 U6819 ( .A1(n5741), .A2(n5740), .ZN(n5742) );
  AND2_X1 U6820 ( .A1(n10597), .A2(n6074), .ZN(n5743) );
  AOI21_X1 U6821 ( .B1(n9560), .B2(n6247), .A(n5743), .ZN(n5747) );
  INV_X1 U6822 ( .A(n5744), .ZN(n5746) );
  NAND2_X1 U6823 ( .A1(n5746), .A2(n5745), .ZN(n7090) );
  INV_X1 U6824 ( .A(n5747), .ZN(n5748) );
  NAND2_X1 U6825 ( .A1(n5749), .A2(n5748), .ZN(n5750) );
  NAND2_X1 U6826 ( .A1(n7087), .A2(n5750), .ZN(n5777) );
  INV_X1 U6827 ( .A(n6337), .ZN(n6108) );
  AOI21_X1 U6828 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5752) );
  NOR2_X1 U6829 ( .A1(n5752), .A2(n5780), .ZN(n7434) );
  NAND2_X1 U6830 ( .A1(n6108), .A2(n7434), .ZN(n5760) );
  INV_X1 U6831 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6647) );
  OR2_X1 U6832 ( .A1(n6446), .A2(n6647), .ZN(n5759) );
  INV_X1 U6833 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5754) );
  OR2_X1 U6834 ( .A1(n6223), .A2(n5754), .ZN(n5758) );
  INV_X1 U6835 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5756) );
  OR2_X1 U6836 ( .A1(n6448), .A2(n5756), .ZN(n5757) );
  NAND4_X1 U6837 ( .A1(n5760), .A2(n5759), .A3(n5758), .A4(n5757), .ZN(n7514)
         );
  NAND2_X1 U6838 ( .A1(n7514), .A2(n6074), .ZN(n5774) );
  NAND2_X1 U6839 ( .A1(n5724), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5761) );
  MUX2_X1 U6840 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5761), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5763) );
  AND2_X1 U6841 ( .A1(n5763), .A2(n5762), .ZN(n6656) );
  INV_X1 U6842 ( .A(n6656), .ZN(n6665) );
  NAND2_X1 U6843 ( .A1(n5766), .A2(SI_5_), .ZN(n5787) );
  INV_X1 U6844 ( .A(n5766), .ZN(n5767) );
  INV_X1 U6845 ( .A(SI_5_), .ZN(n10098) );
  NAND2_X1 U6846 ( .A1(n5767), .A2(n10098), .ZN(n5768) );
  OR2_X1 U6847 ( .A1(n5769), .A2(n4962), .ZN(n5770) );
  OR2_X1 U6848 ( .A1(n5726), .A2(n7126), .ZN(n5772) );
  INV_X1 U6849 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6405) );
  OR2_X1 U6850 ( .A1(n9296), .A2(n6405), .ZN(n5771) );
  NAND2_X1 U6851 ( .A1(n7432), .A2(n5083), .ZN(n5773) );
  NAND2_X1 U6852 ( .A1(n5774), .A2(n5773), .ZN(n5775) );
  XNOR2_X1 U6853 ( .A(n5775), .B(n5633), .ZN(n5778) );
  AND2_X1 U6854 ( .A1(n7432), .A2(n6282), .ZN(n5776) );
  AOI21_X1 U6855 ( .B1(n7514), .B2(n6247), .A(n5776), .ZN(n7259) );
  NAND2_X1 U6856 ( .A1(n6283), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5784) );
  INV_X1 U6857 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6666) );
  OR2_X1 U6858 ( .A1(n6446), .A2(n6666), .ZN(n5783) );
  NAND2_X1 U6859 ( .A1(n5780), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5838) );
  OAI21_X1 U6860 ( .B1(n5780), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5838), .ZN(
        n7453) );
  OR2_X1 U6861 ( .A1(n6337), .A2(n7453), .ZN(n5782) );
  INV_X1 U6862 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7454) );
  OR2_X1 U6863 ( .A1(n6448), .A2(n7454), .ZN(n5781) );
  NAND4_X1 U6864 ( .A1(n5784), .A2(n5783), .A3(n5782), .A4(n5781), .ZN(n9559)
         );
  NAND2_X1 U6865 ( .A1(n9559), .A2(n6074), .ZN(n5794) );
  NAND2_X1 U6866 ( .A1(n5762), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5786) );
  INV_X1 U6867 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5785) );
  XNOR2_X1 U6868 ( .A(n5786), .B(n5785), .ZN(n6784) );
  MUX2_X1 U6869 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6594), .Z(n5789) );
  NAND2_X1 U6870 ( .A1(n5789), .A2(SI_6_), .ZN(n5809) );
  INV_X1 U6871 ( .A(n5789), .ZN(n5790) );
  INV_X1 U6872 ( .A(SI_6_), .ZN(n10097) );
  NAND2_X1 U6873 ( .A1(n5790), .A2(n10097), .ZN(n5791) );
  INV_X1 U6874 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U6875 ( .A1(n7456), .A2(n5083), .ZN(n5793) );
  NAND2_X1 U6876 ( .A1(n5794), .A2(n5793), .ZN(n5795) );
  XNOR2_X1 U6877 ( .A(n5795), .B(n5662), .ZN(n5797) );
  AND2_X1 U6878 ( .A1(n7456), .A2(n6282), .ZN(n5796) );
  AOI21_X1 U6879 ( .B1(n9559), .B2(n6247), .A(n5796), .ZN(n5798) );
  NAND2_X1 U6880 ( .A1(n5797), .A2(n5798), .ZN(n5802) );
  INV_X1 U6881 ( .A(n5797), .ZN(n5800) );
  INV_X1 U6882 ( .A(n5798), .ZN(n5799) );
  NAND2_X1 U6883 ( .A1(n5800), .A2(n5799), .ZN(n5801) );
  AND2_X1 U6884 ( .A1(n5802), .A2(n5801), .ZN(n7292) );
  NAND2_X1 U6885 ( .A1(n6283), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5808) );
  INV_X1 U6886 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5803) );
  OR2_X1 U6887 ( .A1(n6448), .A2(n5803), .ZN(n5807) );
  INV_X1 U6888 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5804) );
  XNOR2_X1 U6889 ( .A(n5838), .B(n5804), .ZN(n7559) );
  OR2_X1 U6890 ( .A1(n6337), .A2(n7559), .ZN(n5806) );
  INV_X1 U6891 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6663) );
  OR2_X1 U6892 ( .A1(n6446), .A2(n6663), .ZN(n5805) );
  NAND4_X1 U6893 ( .A1(n5808), .A2(n5807), .A3(n5806), .A4(n5805), .ZN(n9558)
         );
  NAND2_X1 U6894 ( .A1(n9558), .A2(n6282), .ZN(n5822) );
  MUX2_X1 U6895 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6594), .Z(n5811) );
  NAND2_X1 U6896 ( .A1(n5811), .A2(SI_7_), .ZN(n5830) );
  INV_X1 U6897 ( .A(n5811), .ZN(n5812) );
  INV_X1 U6898 ( .A(SI_7_), .ZN(n10208) );
  NAND2_X1 U6899 ( .A1(n5812), .A2(n10208), .ZN(n5813) );
  OR2_X1 U6900 ( .A1(n7364), .A2(n5726), .ZN(n5820) );
  INV_X2 U6901 ( .A(n5086), .ZN(n6083) );
  OR2_X1 U6902 ( .A1(n5817), .A2(n5604), .ZN(n5818) );
  XNOR2_X1 U6903 ( .A(n5818), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6705) );
  AOI22_X1 U6904 ( .A1(n5520), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6083), .B2(
        n6705), .ZN(n5819) );
  NAND2_X1 U6905 ( .A1(n7566), .A2(n5083), .ZN(n5821) );
  NAND2_X1 U6906 ( .A1(n5822), .A2(n5821), .ZN(n5823) );
  XNOR2_X1 U6907 ( .A(n5823), .B(n5662), .ZN(n5828) );
  NAND2_X1 U6908 ( .A1(n9558), .A2(n6247), .ZN(n5825) );
  NAND2_X1 U6909 ( .A1(n7566), .A2(n6074), .ZN(n5824) );
  NAND2_X1 U6910 ( .A1(n5825), .A2(n5824), .ZN(n5826) );
  XNOR2_X1 U6911 ( .A(n5828), .B(n5826), .ZN(n7384) );
  INV_X1 U6912 ( .A(n5826), .ZN(n5827) );
  NAND2_X1 U6913 ( .A1(n5828), .A2(n5827), .ZN(n5829) );
  MUX2_X1 U6914 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n6594), .Z(n5852) );
  XNOR2_X1 U6915 ( .A(n5852), .B(SI_8_), .ZN(n5855) );
  XNOR2_X1 U6916 ( .A(n5856), .B(n5855), .ZN(n7570) );
  NAND2_X1 U6917 ( .A1(n7570), .A2(n9335), .ZN(n5835) );
  NAND2_X1 U6918 ( .A1(n5832), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5833) );
  XNOR2_X1 U6919 ( .A(n5833), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6706) );
  AOI22_X1 U6920 ( .A1(n5520), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6083), .B2(
        n6706), .ZN(n5834) );
  NAND2_X1 U6921 ( .A1(n7676), .A2(n5083), .ZN(n5846) );
  NAND2_X1 U6922 ( .A1(n4932), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5843) );
  OR2_X1 U6923 ( .A1(n6223), .A2(n10652), .ZN(n5842) );
  INV_X1 U6924 ( .A(n5838), .ZN(n5836) );
  AOI21_X1 U6925 ( .B1(n5836), .B2(P1_REG3_REG_7__SCAN_IN), .A(
        P1_REG3_REG_8__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U6926 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n5837) );
  NOR2_X1 U6927 ( .A1(n5838), .A2(n5837), .ZN(n5859) );
  OR2_X1 U6928 ( .A1(n5839), .A2(n5859), .ZN(n7666) );
  OR2_X1 U6929 ( .A1(n6337), .A2(n7666), .ZN(n5841) );
  INV_X1 U6930 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7667) );
  OR2_X1 U6931 ( .A1(n6448), .A2(n7667), .ZN(n5840) );
  NAND4_X1 U6932 ( .A1(n5843), .A2(n5842), .A3(n5841), .A4(n5840), .ZN(n10661)
         );
  INV_X2 U6933 ( .A(n5844), .ZN(n6282) );
  NAND2_X1 U6934 ( .A1(n10661), .A2(n6282), .ZN(n5845) );
  NAND2_X1 U6935 ( .A1(n5846), .A2(n5845), .ZN(n5847) );
  XNOR2_X1 U6936 ( .A(n5847), .B(n5662), .ZN(n5850) );
  AND2_X1 U6937 ( .A1(n10661), .A2(n6247), .ZN(n5849) );
  AOI21_X1 U6938 ( .B1(n7676), .B2(n6282), .A(n5849), .ZN(n7650) );
  INV_X1 U6939 ( .A(n5852), .ZN(n5853) );
  NAND2_X1 U6940 ( .A1(n5853), .A2(n10210), .ZN(n5854) );
  MUX2_X1 U6941 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n6594), .Z(n5873) );
  XNOR2_X1 U6942 ( .A(n5873), .B(n10203), .ZN(n5874) );
  NAND2_X1 U6943 ( .A1(n5857), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5882) );
  XNOR2_X1 U6944 ( .A(n5882), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6728) );
  AOI22_X1 U6945 ( .A1(n5520), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6083), .B2(
        n6728), .ZN(n5858) );
  NAND2_X1 U6946 ( .A1(n10662), .A2(n5083), .ZN(n5866) );
  NAND2_X1 U6947 ( .A1(n6283), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5864) );
  INV_X1 U6948 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6699) );
  OR2_X1 U6949 ( .A1(n6446), .A2(n6699), .ZN(n5863) );
  NAND2_X1 U6950 ( .A1(n5859), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5886) );
  OR2_X1 U6951 ( .A1(n5859), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U6952 ( .A1(n5886), .A2(n5860), .ZN(n7697) );
  OR2_X1 U6953 ( .A1(n6337), .A2(n7697), .ZN(n5862) );
  INV_X1 U6954 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7680) );
  OR2_X1 U6955 ( .A1(n6448), .A2(n7680), .ZN(n5861) );
  NAND4_X1 U6956 ( .A1(n5864), .A2(n5863), .A3(n5862), .A4(n5861), .ZN(n10679)
         );
  NAND2_X1 U6957 ( .A1(n10679), .A2(n6282), .ZN(n5865) );
  NAND2_X1 U6958 ( .A1(n5866), .A2(n5865), .ZN(n5867) );
  XNOR2_X1 U6959 ( .A(n5867), .B(n5662), .ZN(n5869) );
  AND2_X1 U6960 ( .A1(n10679), .A2(n6247), .ZN(n5868) );
  AOI21_X1 U6961 ( .B1(n10662), .B2(n6282), .A(n5868), .ZN(n5870) );
  AND2_X1 U6962 ( .A1(n5869), .A2(n5870), .ZN(n7692) );
  INV_X1 U6963 ( .A(n5869), .ZN(n5872) );
  INV_X1 U6964 ( .A(n5870), .ZN(n5871) );
  NAND2_X1 U6965 ( .A1(n5872), .A2(n5871), .ZN(n7693) );
  MUX2_X1 U6966 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6594), .Z(n5875) );
  NAND2_X1 U6967 ( .A1(n5875), .A2(SI_10_), .ZN(n5898) );
  INV_X1 U6968 ( .A(n5875), .ZN(n5876) );
  NAND2_X1 U6969 ( .A1(n5876), .A2(n10199), .ZN(n5877) );
  NAND2_X1 U6970 ( .A1(n5898), .A2(n5877), .ZN(n5880) );
  INV_X1 U6971 ( .A(n5880), .ZN(n5878) );
  NAND2_X1 U6972 ( .A1(n5882), .A2(n5881), .ZN(n5883) );
  NAND2_X1 U6973 ( .A1(n5883), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5901) );
  XNOR2_X1 U6974 ( .A(n5901), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6886) );
  AOI22_X1 U6975 ( .A1(n5520), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6083), .B2(
        n6886), .ZN(n5884) );
  NAND2_X1 U6976 ( .A1(n10680), .A2(n5083), .ZN(n5893) );
  NAND2_X1 U6977 ( .A1(n6283), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5891) );
  INV_X1 U6978 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6733) );
  OR2_X1 U6979 ( .A1(n6446), .A2(n6733), .ZN(n5890) );
  INV_X1 U6980 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U6981 ( .A1(n5886), .A2(n5885), .ZN(n5887) );
  NAND2_X1 U6982 ( .A1(n5907), .A2(n5887), .ZN(n7824) );
  OR2_X1 U6983 ( .A1(n6337), .A2(n7824), .ZN(n5889) );
  INV_X1 U6984 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7722) );
  OR2_X1 U6985 ( .A1(n6448), .A2(n7722), .ZN(n5888) );
  NAND4_X1 U6986 ( .A1(n5891), .A2(n5890), .A3(n5889), .A4(n5888), .ZN(n9557)
         );
  NAND2_X1 U6987 ( .A1(n9557), .A2(n6282), .ZN(n5892) );
  NAND2_X1 U6988 ( .A1(n5893), .A2(n5892), .ZN(n5894) );
  XNOR2_X1 U6989 ( .A(n5894), .B(n5633), .ZN(n5896) );
  AND2_X1 U6990 ( .A1(n9557), .A2(n6247), .ZN(n5895) );
  AOI21_X1 U6991 ( .B1(n10680), .B2(n6282), .A(n5895), .ZN(n7821) );
  INV_X1 U6992 ( .A(n5896), .ZN(n5897) );
  MUX2_X1 U6993 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6594), .Z(n5921) );
  XNOR2_X1 U6994 ( .A(n5921), .B(SI_11_), .ZN(n5922) );
  XNOR2_X1 U6995 ( .A(n5923), .B(n5922), .ZN(n7836) );
  NAND2_X1 U6996 ( .A1(n7836), .A2(n9335), .ZN(n5905) );
  NAND2_X1 U6997 ( .A1(n5901), .A2(n5900), .ZN(n5902) );
  NAND2_X1 U6998 ( .A1(n5902), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5903) );
  XNOR2_X1 U6999 ( .A(n5903), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7157) );
  AOI22_X1 U7000 ( .A1(n5520), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6083), .B2(
        n7157), .ZN(n5904) );
  NAND2_X1 U7001 ( .A1(n7802), .A2(n5083), .ZN(n5914) );
  NAND2_X1 U7002 ( .A1(n6283), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5912) );
  INV_X1 U7003 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6889) );
  OR2_X1 U7004 ( .A1(n6446), .A2(n6889), .ZN(n5911) );
  INV_X1 U7005 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7006 ( .A1(n5907), .A2(n5906), .ZN(n5908) );
  NAND2_X1 U7007 ( .A1(n5934), .A2(n5908), .ZN(n7877) );
  OR2_X1 U7008 ( .A1(n6337), .A2(n7877), .ZN(n5910) );
  INV_X1 U7009 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7789) );
  OR2_X1 U7010 ( .A1(n6448), .A2(n7789), .ZN(n5909) );
  NAND4_X1 U7011 ( .A1(n5912), .A2(n5911), .A3(n5910), .A4(n5909), .ZN(n10703)
         );
  NAND2_X1 U7012 ( .A1(n10703), .A2(n6282), .ZN(n5913) );
  NAND2_X1 U7013 ( .A1(n5914), .A2(n5913), .ZN(n5915) );
  XNOR2_X1 U7014 ( .A(n5915), .B(n5662), .ZN(n5917) );
  AND2_X1 U7015 ( .A1(n10703), .A2(n6247), .ZN(n5916) );
  AOI21_X1 U7016 ( .B1(n7802), .B2(n6282), .A(n5916), .ZN(n5918) );
  AND2_X1 U7017 ( .A1(n5917), .A2(n5918), .ZN(n7873) );
  INV_X1 U7018 ( .A(n5917), .ZN(n5920) );
  INV_X1 U7019 ( .A(n5918), .ZN(n5919) );
  MUX2_X1 U7020 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6594), .Z(n5924) );
  NAND2_X1 U7021 ( .A1(n5924), .A2(SI_12_), .ZN(n5948) );
  OAI21_X1 U7022 ( .B1(n5924), .B2(SI_12_), .A(n5948), .ZN(n5925) );
  NAND2_X1 U7023 ( .A1(n5926), .A2(n5925), .ZN(n5927) );
  NAND2_X1 U7024 ( .A1(n5927), .A2(n5949), .ZN(n7927) );
  OR2_X1 U7025 ( .A1(n7927), .A2(n5726), .ZN(n5931) );
  OR2_X1 U7026 ( .A1(n5928), .A2(n5604), .ZN(n5929) );
  XNOR2_X1 U7027 ( .A(n5929), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7162) );
  AOI22_X1 U7028 ( .A1(n5520), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6083), .B2(
        n7162), .ZN(n5930) );
  NAND2_X1 U7029 ( .A1(n10706), .A2(n5083), .ZN(n5942) );
  NAND2_X1 U7030 ( .A1(n6283), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5940) );
  INV_X1 U7031 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5932) );
  OR2_X1 U7032 ( .A1(n6446), .A2(n5932), .ZN(n5939) );
  INV_X1 U7033 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5933) );
  AND2_X1 U7034 ( .A1(n5934), .A2(n5933), .ZN(n5935) );
  OR2_X1 U7035 ( .A1(n5935), .A2(n5964), .ZN(n7902) );
  OR2_X1 U7036 ( .A1(n6337), .A2(n7902), .ZN(n5938) );
  INV_X1 U7037 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n5936) );
  OR2_X1 U7038 ( .A1(n6448), .A2(n5936), .ZN(n5937) );
  NAND4_X1 U7039 ( .A1(n5940), .A2(n5939), .A3(n5938), .A4(n5937), .ZN(n9556)
         );
  NAND2_X1 U7040 ( .A1(n9556), .A2(n6282), .ZN(n5941) );
  NAND2_X1 U7041 ( .A1(n5942), .A2(n5941), .ZN(n5943) );
  XNOR2_X1 U7042 ( .A(n5943), .B(n5662), .ZN(n5946) );
  AND2_X1 U7043 ( .A1(n9556), .A2(n6247), .ZN(n5944) );
  AOI21_X1 U7044 ( .B1(n10706), .B2(n6282), .A(n5944), .ZN(n5945) );
  XNOR2_X1 U7045 ( .A(n5946), .B(n5945), .ZN(n7901) );
  NAND2_X1 U7046 ( .A1(n5946), .A2(n5945), .ZN(n5947) );
  MUX2_X1 U7047 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6594), .Z(n5950) );
  NAND2_X1 U7048 ( .A1(n5950), .A2(SI_13_), .ZN(n5979) );
  INV_X1 U7049 ( .A(n5950), .ZN(n5952) );
  INV_X1 U7050 ( .A(SI_13_), .ZN(n5951) );
  NAND2_X1 U7051 ( .A1(n5952), .A2(n5951), .ZN(n5953) );
  OR2_X1 U7052 ( .A1(n5955), .A2(n5954), .ZN(n5956) );
  NAND2_X1 U7053 ( .A1(n5980), .A2(n5956), .ZN(n8036) );
  OR2_X1 U7054 ( .A1(n8036), .A2(n5726), .ZN(n5963) );
  NOR2_X1 U7055 ( .A1(n5957), .A2(n5604), .ZN(n5958) );
  MUX2_X1 U7056 ( .A(n5604), .B(n5958), .S(P1_IR_REG_13__SCAN_IN), .Z(n5959)
         );
  INV_X1 U7057 ( .A(n5959), .ZN(n5961) );
  NAND2_X1 U7058 ( .A1(n5957), .A2(n5960), .ZN(n6006) );
  AOI22_X1 U7059 ( .A1(n5520), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6083), .B2(
        n7623), .ZN(n5962) );
  NAND2_X1 U7060 ( .A1(n7958), .A2(n5083), .ZN(n5971) );
  NAND2_X1 U7061 ( .A1(n6283), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5969) );
  INV_X1 U7062 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7164) );
  OR2_X1 U7063 ( .A1(n6446), .A2(n7164), .ZN(n5968) );
  NAND2_X1 U7064 ( .A1(n5964), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5985) );
  OR2_X1 U7065 ( .A1(n5964), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7066 ( .A1(n5985), .A2(n5965), .ZN(n8007) );
  OR2_X1 U7067 ( .A1(n6337), .A2(n8007), .ZN(n5967) );
  INV_X1 U7068 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7920) );
  OR2_X1 U7069 ( .A1(n6448), .A2(n7920), .ZN(n5966) );
  NAND4_X1 U7070 ( .A1(n5969), .A2(n5968), .A3(n5967), .A4(n5966), .ZN(n7964)
         );
  NAND2_X1 U7071 ( .A1(n7964), .A2(n6282), .ZN(n5970) );
  NAND2_X1 U7072 ( .A1(n5971), .A2(n5970), .ZN(n5972) );
  XNOR2_X1 U7073 ( .A(n5972), .B(n5662), .ZN(n5974) );
  AND2_X1 U7074 ( .A1(n7964), .A2(n6247), .ZN(n5973) );
  AOI21_X1 U7075 ( .B1(n7958), .B2(n6282), .A(n5973), .ZN(n5975) );
  XNOR2_X1 U7076 ( .A(n5974), .B(n5975), .ZN(n8003) );
  INV_X1 U7077 ( .A(n5974), .ZN(n5977) );
  INV_X1 U7078 ( .A(n5975), .ZN(n5976) );
  NAND2_X1 U7079 ( .A1(n5977), .A2(n5976), .ZN(n5978) );
  MUX2_X1 U7080 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6594), .Z(n5999) );
  XNOR2_X1 U7081 ( .A(n6001), .B(n6000), .ZN(n8039) );
  NAND2_X1 U7082 ( .A1(n8039), .A2(n9335), .ZN(n5983) );
  NAND2_X1 U7083 ( .A1(n6006), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5981) );
  XNOR2_X1 U7084 ( .A(n5981), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7624) );
  AOI22_X1 U7085 ( .A1(n5520), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6083), .B2(
        n7624), .ZN(n5982) );
  NAND2_X1 U7086 ( .A1(n9171), .A2(n5083), .ZN(n5992) );
  NAND2_X1 U7087 ( .A1(n6283), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5990) );
  INV_X1 U7088 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7617) );
  OR2_X1 U7089 ( .A1(n6446), .A2(n7617), .ZN(n5989) );
  INV_X1 U7090 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7091 ( .A1(n5985), .A2(n5984), .ZN(n5986) );
  NAND2_X1 U7092 ( .A1(n6012), .A2(n5986), .ZN(n9168) );
  OR2_X1 U7093 ( .A1(n6337), .A2(n9168), .ZN(n5988) );
  INV_X1 U7094 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7972) );
  OR2_X1 U7095 ( .A1(n6448), .A2(n7972), .ZN(n5987) );
  NAND4_X1 U7096 ( .A1(n5990), .A2(n5989), .A3(n5988), .A4(n5987), .ZN(n9555)
         );
  NAND2_X1 U7097 ( .A1(n9555), .A2(n6282), .ZN(n5991) );
  NAND2_X1 U7098 ( .A1(n5992), .A2(n5991), .ZN(n5993) );
  XNOR2_X1 U7099 ( .A(n5993), .B(n5662), .ZN(n5996) );
  NAND2_X1 U7100 ( .A1(n9171), .A2(n6282), .ZN(n5995) );
  NAND2_X1 U7101 ( .A1(n9555), .A2(n6247), .ZN(n5994) );
  NAND2_X1 U7102 ( .A1(n5995), .A2(n5994), .ZN(n9165) );
  NAND2_X1 U7103 ( .A1(n9162), .A2(n9165), .ZN(n5998) );
  INV_X1 U7104 ( .A(n5996), .ZN(n5997) );
  MUX2_X1 U7105 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6594), .Z(n6002) );
  OAI21_X1 U7106 ( .B1(n6002), .B2(SI_15_), .A(n6024), .ZN(n6003) );
  NAND2_X1 U7107 ( .A1(n6004), .A2(n6003), .ZN(n6005) );
  NAND2_X1 U7108 ( .A1(n6005), .A2(n6025), .ZN(n8106) );
  OR2_X1 U7109 ( .A1(n8106), .A2(n5726), .ZN(n6009) );
  NAND2_X1 U7110 ( .A1(n6007), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6027) );
  XNOR2_X1 U7111 ( .A(n6027), .B(P1_IR_REG_15__SCAN_IN), .ZN(n7853) );
  AOI22_X1 U7112 ( .A1(n5520), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6083), .B2(
        n7853), .ZN(n6008) );
  NAND2_X1 U7113 ( .A1(n9632), .A2(n5083), .ZN(n6020) );
  NAND2_X1 U7114 ( .A1(n6283), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6018) );
  INV_X1 U7115 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6010) );
  OR2_X1 U7116 ( .A1(n6446), .A2(n6010), .ZN(n6017) );
  INV_X1 U7117 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6011) );
  AND2_X1 U7118 ( .A1(n6012), .A2(n6011), .ZN(n6013) );
  OR2_X1 U7119 ( .A1(n6013), .A2(n6032), .ZN(n9274) );
  OR2_X1 U7120 ( .A1(n6337), .A2(n9274), .ZN(n6016) );
  INV_X1 U7121 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6014) );
  OR2_X1 U7122 ( .A1(n6448), .A2(n6014), .ZN(n6015) );
  NAND4_X1 U7123 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .ZN(n9631)
         );
  NAND2_X1 U7124 ( .A1(n9631), .A2(n6282), .ZN(n6019) );
  NAND2_X1 U7125 ( .A1(n6020), .A2(n6019), .ZN(n6021) );
  XNOR2_X1 U7126 ( .A(n6021), .B(n5633), .ZN(n6022) );
  AOI22_X1 U7127 ( .A1(n9632), .A2(n6282), .B1(n6247), .B2(n9631), .ZN(n9272)
         );
  NAND2_X1 U7128 ( .A1(n6023), .A2(n6022), .ZN(n9270) );
  MUX2_X1 U7129 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6594), .Z(n6043) );
  XNOR2_X1 U7130 ( .A(n6043), .B(SI_16_), .ZN(n6041) );
  XNOR2_X1 U7131 ( .A(n6042), .B(n6041), .ZN(n8102) );
  NAND2_X1 U7132 ( .A1(n8102), .A2(n9335), .ZN(n6031) );
  NAND2_X1 U7133 ( .A1(n6027), .A2(n6026), .ZN(n6028) );
  NAND2_X1 U7134 ( .A1(n6028), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6029) );
  XNOR2_X1 U7135 ( .A(n6029), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9564) );
  AOI22_X1 U7136 ( .A1(n5520), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6083), .B2(
        n9564), .ZN(n6030) );
  NAND2_X1 U7137 ( .A1(n6283), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6037) );
  INV_X1 U7138 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9887) );
  OR2_X1 U7139 ( .A1(n6448), .A2(n9887), .ZN(n6036) );
  NOR2_X1 U7140 ( .A1(n6032), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6033) );
  OR2_X1 U7141 ( .A1(n6050), .A2(n6033), .ZN(n9881) );
  OR2_X1 U7142 ( .A1(n6337), .A2(n9881), .ZN(n6035) );
  INV_X1 U7143 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7856) );
  OR2_X1 U7144 ( .A1(n6446), .A2(n7856), .ZN(n6034) );
  NAND4_X1 U7145 ( .A1(n6037), .A2(n6036), .A3(n6035), .A4(n6034), .ZN(n9554)
         );
  AOI22_X1 U7146 ( .A1(n9982), .A2(n5083), .B1(n6282), .B2(n9554), .ZN(n6038)
         );
  XNOR2_X1 U7147 ( .A(n6038), .B(n5633), .ZN(n6040) );
  AOI22_X1 U7148 ( .A1(n9982), .A2(n6074), .B1(n6247), .B2(n9554), .ZN(n6039)
         );
  XNOR2_X1 U7149 ( .A(n6040), .B(n6039), .ZN(n9206) );
  INV_X1 U7150 ( .A(n6043), .ZN(n6044) );
  NAND2_X1 U7151 ( .A1(n6044), .A2(n10195), .ZN(n6045) );
  MUX2_X1 U7152 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n6594), .Z(n6060) );
  XNOR2_X1 U7153 ( .A(n6062), .B(n6061), .ZN(n8110) );
  NAND2_X1 U7154 ( .A1(n8110), .A2(n9335), .ZN(n6049) );
  NAND2_X1 U7155 ( .A1(n5024), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6047) );
  XNOR2_X1 U7156 ( .A(n6047), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9587) );
  AOI22_X1 U7157 ( .A1(n5520), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6083), .B2(
        n9587), .ZN(n6048) );
  NAND2_X1 U7158 ( .A1(n6283), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6055) );
  INV_X1 U7159 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9978) );
  OR2_X1 U7160 ( .A1(n6446), .A2(n9978), .ZN(n6054) );
  OR2_X1 U7161 ( .A1(n6050), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7162 ( .A1(n6090), .A2(n6051), .ZN(n9856) );
  OR2_X1 U7163 ( .A1(n6337), .A2(n9856), .ZN(n6053) );
  INV_X1 U7164 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9565) );
  OR2_X1 U7165 ( .A1(n6448), .A2(n9565), .ZN(n6052) );
  NAND4_X1 U7166 ( .A1(n6055), .A2(n6054), .A3(n6053), .A4(n6052), .ZN(n9635)
         );
  AOI22_X1 U7167 ( .A1(n9868), .A2(n5083), .B1(n6282), .B2(n9635), .ZN(n6056)
         );
  XOR2_X1 U7168 ( .A(n5633), .B(n6056), .Z(n9213) );
  NAND2_X1 U7169 ( .A1(n9868), .A2(n6282), .ZN(n6058) );
  NAND2_X1 U7170 ( .A1(n9635), .A2(n6247), .ZN(n6057) );
  NAND2_X1 U7171 ( .A1(n6058), .A2(n6057), .ZN(n6059) );
  INV_X1 U7172 ( .A(n6059), .ZN(n9212) );
  MUX2_X1 U7173 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6594), .Z(n6063) );
  NAND2_X1 U7174 ( .A1(n6063), .A2(SI_18_), .ZN(n6081) );
  INV_X1 U7175 ( .A(n6063), .ZN(n6065) );
  INV_X1 U7176 ( .A(SI_18_), .ZN(n6064) );
  NAND2_X1 U7177 ( .A1(n6065), .A2(n6064), .ZN(n6066) );
  NAND2_X1 U7178 ( .A1(n6081), .A2(n6066), .ZN(n6068) );
  INV_X1 U7179 ( .A(n6068), .ZN(n6067) );
  NAND2_X1 U7180 ( .A1(n4946), .A2(n6068), .ZN(n6069) );
  NAND2_X1 U7181 ( .A1(n6082), .A2(n6069), .ZN(n8119) );
  OR2_X1 U7182 ( .A1(n8119), .A2(n5726), .ZN(n6073) );
  NAND2_X1 U7183 ( .A1(n5025), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n6071) );
  AND2_X1 U7184 ( .A1(n6071), .A2(n6070), .ZN(n9602) );
  AOI22_X1 U7185 ( .A1(n5520), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6083), .B2(
        n9602), .ZN(n6072) );
  NAND2_X1 U7186 ( .A1(n4932), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6078) );
  INV_X1 U7187 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10029) );
  OR2_X1 U7188 ( .A1(n6223), .A2(n10029), .ZN(n6077) );
  INV_X1 U7189 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6088) );
  XNOR2_X1 U7190 ( .A(n6090), .B(n6088), .ZN(n9841) );
  OR2_X1 U7191 ( .A1(n6337), .A2(n9841), .ZN(n6076) );
  INV_X1 U7192 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9588) );
  OR2_X1 U7193 ( .A1(n6448), .A2(n9588), .ZN(n6075) );
  NAND4_X1 U7194 ( .A1(n6078), .A2(n6077), .A3(n6076), .A4(n6075), .ZN(n9851)
         );
  OAI22_X1 U7195 ( .A1(n10031), .A2(n5844), .B1(n9822), .B2(n6291), .ZN(n6080)
         );
  AOI22_X1 U7196 ( .A1(n9847), .A2(n5083), .B1(n6282), .B2(n9851), .ZN(n6079)
         );
  XOR2_X1 U7197 ( .A(n5633), .B(n6079), .Z(n9252) );
  INV_X1 U7198 ( .A(n6080), .ZN(n9251) );
  MUX2_X1 U7199 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n6594), .Z(n6100) );
  XNOR2_X1 U7200 ( .A(n6100), .B(SI_19_), .ZN(n6102) );
  XNOR2_X1 U7201 ( .A(n6103), .B(n6102), .ZN(n8130) );
  NAND2_X1 U7202 ( .A1(n8130), .A2(n9335), .ZN(n6085) );
  AOI22_X1 U7203 ( .A1(n5520), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9610), .B2(
        n6083), .ZN(n6084) );
  NAND2_X1 U7204 ( .A1(n6283), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6095) );
  INV_X1 U7205 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n6086) );
  OR2_X1 U7206 ( .A1(n6446), .A2(n6086), .ZN(n6094) );
  INV_X1 U7207 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6087) );
  OAI21_X1 U7208 ( .B1(n6090), .B2(n6088), .A(n6087), .ZN(n6091) );
  NAND2_X1 U7209 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n6089) );
  NAND2_X1 U7210 ( .A1(n6091), .A2(n6106), .ZN(n9828) );
  OR2_X1 U7211 ( .A1(n6337), .A2(n9828), .ZN(n6093) );
  INV_X1 U7212 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9829) );
  OR2_X1 U7213 ( .A1(n6448), .A2(n9829), .ZN(n6092) );
  NAND4_X1 U7214 ( .A1(n6095), .A2(n6094), .A3(n6093), .A4(n6092), .ZN(n9836)
         );
  AOI22_X1 U7215 ( .A1(n9962), .A2(n5083), .B1(n6282), .B2(n9836), .ZN(n6096)
         );
  XNOR2_X1 U7216 ( .A(n6096), .B(n5633), .ZN(n6098) );
  AOI22_X1 U7217 ( .A1(n9962), .A2(n6282), .B1(n6247), .B2(n9836), .ZN(n6097)
         );
  NAND2_X1 U7218 ( .A1(n6098), .A2(n6097), .ZN(n6099) );
  OAI21_X1 U7219 ( .B1(n6098), .B2(n6097), .A(n6099), .ZN(n9183) );
  INV_X1 U7220 ( .A(n6099), .ZN(n9233) );
  INV_X1 U7221 ( .A(n6100), .ZN(n6101) );
  INV_X1 U7222 ( .A(SI_19_), .ZN(n10192) );
  MUX2_X1 U7223 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6594), .Z(n6124) );
  XNOR2_X1 U7224 ( .A(n6124), .B(n10186), .ZN(n6126) );
  XNOR2_X1 U7225 ( .A(n6127), .B(n6126), .ZN(n8143) );
  NAND2_X1 U7226 ( .A1(n8143), .A2(n9335), .ZN(n6105) );
  INV_X1 U7227 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7746) );
  NAND2_X1 U7228 ( .A1(n9813), .A2(n5083), .ZN(n6115) );
  INV_X1 U7229 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9236) );
  AND2_X1 U7230 ( .A1(n6106), .A2(n9236), .ZN(n6107) );
  NOR2_X1 U7231 ( .A1(n6139), .A2(n6107), .ZN(n9814) );
  NAND2_X1 U7232 ( .A1(n6108), .A2(n9814), .ZN(n6113) );
  INV_X1 U7233 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10025) );
  OR2_X1 U7234 ( .A1(n6223), .A2(n10025), .ZN(n6112) );
  INV_X1 U7235 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9957) );
  OR2_X1 U7236 ( .A1(n6446), .A2(n9957), .ZN(n6111) );
  INV_X1 U7237 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n6109) );
  OR2_X1 U7238 ( .A1(n6448), .A2(n6109), .ZN(n6110) );
  NAND4_X1 U7239 ( .A1(n6113), .A2(n6112), .A3(n6111), .A4(n6110), .ZN(n9553)
         );
  NAND2_X1 U7240 ( .A1(n9553), .A2(n6282), .ZN(n6114) );
  NAND2_X1 U7241 ( .A1(n6115), .A2(n6114), .ZN(n6116) );
  XNOR2_X1 U7242 ( .A(n6116), .B(n5662), .ZN(n6118) );
  AND2_X1 U7243 ( .A1(n9553), .A2(n6247), .ZN(n6117) );
  AOI21_X1 U7244 ( .B1(n9813), .B2(n6282), .A(n6117), .ZN(n6119) );
  NAND2_X1 U7245 ( .A1(n6118), .A2(n6119), .ZN(n6123) );
  INV_X1 U7246 ( .A(n6118), .ZN(n6121) );
  INV_X1 U7247 ( .A(n6119), .ZN(n6120) );
  NAND2_X1 U7248 ( .A1(n6121), .A2(n6120), .ZN(n6122) );
  AND2_X1 U7249 ( .A1(n6123), .A2(n6122), .ZN(n9232) );
  NOR2_X1 U7250 ( .A1(n6124), .A2(SI_20_), .ZN(n6125) );
  MUX2_X1 U7251 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n6594), .Z(n6128) );
  NAND2_X1 U7252 ( .A1(n6128), .A2(SI_21_), .ZN(n6152) );
  INV_X1 U7253 ( .A(n6128), .ZN(n6129) );
  INV_X1 U7254 ( .A(SI_21_), .ZN(n10183) );
  NAND2_X1 U7255 ( .A1(n6129), .A2(n10183), .ZN(n6130) );
  NAND2_X1 U7256 ( .A1(n6152), .A2(n6130), .ZN(n6133) );
  INV_X1 U7257 ( .A(n6133), .ZN(n6131) );
  INV_X1 U7258 ( .A(n6132), .ZN(n6134) );
  NAND2_X1 U7259 ( .A1(n6134), .A2(n6133), .ZN(n6135) );
  NAND2_X1 U7260 ( .A1(n6153), .A2(n6135), .ZN(n8153) );
  INV_X1 U7261 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7729) );
  OR2_X1 U7262 ( .A1(n9296), .A2(n7729), .ZN(n6136) );
  NAND2_X1 U7263 ( .A1(n9800), .A2(n5083), .ZN(n6146) );
  INV_X1 U7264 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U7265 ( .A1(n6283), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6138) );
  OAI21_X1 U7266 ( .B1(n6446), .B2(n9952), .A(n6138), .ZN(n6144) );
  NOR2_X1 U7267 ( .A1(n6139), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6140) );
  OR2_X1 U7268 ( .A1(n6162), .A2(n6140), .ZN(n9795) );
  INV_X1 U7269 ( .A(n6448), .ZN(n6141) );
  NAND2_X1 U7270 ( .A1(n6141), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6142) );
  OAI21_X1 U7271 ( .B1(n9795), .B2(n6337), .A(n6142), .ZN(n6143) );
  NAND2_X1 U7272 ( .A1(n9809), .A2(n6282), .ZN(n6145) );
  NAND2_X1 U7273 ( .A1(n6146), .A2(n6145), .ZN(n6147) );
  XNOR2_X1 U7274 ( .A(n6147), .B(n5633), .ZN(n6150) );
  AOI22_X1 U7275 ( .A1(n9800), .A2(n6074), .B1(n6247), .B2(n9809), .ZN(n6148)
         );
  XNOR2_X1 U7276 ( .A(n6150), .B(n6148), .ZN(n9190) );
  INV_X1 U7277 ( .A(n6148), .ZN(n6149) );
  MUX2_X1 U7278 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n6594), .Z(n6154) );
  NAND2_X1 U7279 ( .A1(n6154), .A2(SI_22_), .ZN(n6167) );
  INV_X1 U7280 ( .A(n6154), .ZN(n6155) );
  NAND2_X1 U7281 ( .A1(n6155), .A2(n10180), .ZN(n6156) );
  OR2_X1 U7282 ( .A1(n6158), .A2(n6157), .ZN(n6159) );
  NAND2_X1 U7283 ( .A1(n6168), .A2(n6159), .ZN(n8165) );
  OR2_X1 U7284 ( .A1(n8165), .A2(n5726), .ZN(n6161) );
  INV_X1 U7285 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8095) );
  OR2_X1 U7286 ( .A1(n9296), .A2(n8095), .ZN(n6160) );
  NOR2_X1 U7287 ( .A1(n6162), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6163) );
  OR2_X1 U7288 ( .A1(n6171), .A2(n6163), .ZN(n9782) );
  AOI22_X1 U7289 ( .A1(n4932), .A2(P1_REG1_REG_22__SCAN_IN), .B1(n6283), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7290 ( .A1(n6141), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6164) );
  OAI211_X1 U7291 ( .C1(n9782), .C2(n6337), .A(n6165), .B(n6164), .ZN(n9791)
         );
  AOI22_X1 U7292 ( .A1(n9944), .A2(n5083), .B1(n6282), .B2(n9791), .ZN(n6166)
         );
  XNOR2_X1 U7293 ( .A(n6166), .B(n5633), .ZN(n6184) );
  INV_X1 U7294 ( .A(n9791), .ZN(n9638) );
  OAI22_X1 U7295 ( .A1(n9786), .A2(n5844), .B1(n9638), .B2(n6291), .ZN(n9245)
         );
  MUX2_X1 U7296 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n6594), .Z(n6187) );
  XNOR2_X1 U7297 ( .A(n6187), .B(SI_23_), .ZN(n6189) );
  XNOR2_X1 U7298 ( .A(n6190), .B(n6189), .ZN(n8174) );
  NAND2_X1 U7299 ( .A1(n8174), .A2(n9335), .ZN(n6170) );
  INV_X1 U7300 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7816) );
  OR2_X1 U7301 ( .A1(n9296), .A2(n7816), .ZN(n6169) );
  NAND2_X1 U7302 ( .A1(n9764), .A2(n5083), .ZN(n6176) );
  OR2_X1 U7303 ( .A1(n6171), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7304 ( .A1(n6171), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7305 ( .A1(n6172), .A2(n6194), .ZN(n9765) );
  AOI22_X1 U7306 ( .A1(n4932), .A2(P1_REG1_REG_23__SCAN_IN), .B1(n6283), .B2(
        P1_REG0_REG_23__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7307 ( .A1(n6141), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6173) );
  OAI211_X1 U7308 ( .C1(n9765), .C2(n6337), .A(n6174), .B(n6173), .ZN(n9639)
         );
  NAND2_X1 U7309 ( .A1(n9639), .A2(n6282), .ZN(n6175) );
  NAND2_X1 U7310 ( .A1(n6176), .A2(n6175), .ZN(n6177) );
  XNOR2_X1 U7311 ( .A(n6177), .B(n5662), .ZN(n6179) );
  AND2_X1 U7312 ( .A1(n9639), .A2(n6247), .ZN(n6178) );
  AOI21_X1 U7313 ( .B1(n9764), .B2(n6282), .A(n6178), .ZN(n6180) );
  NAND2_X1 U7314 ( .A1(n6179), .A2(n6180), .ZN(n6186) );
  INV_X1 U7315 ( .A(n6179), .ZN(n6182) );
  INV_X1 U7316 ( .A(n6180), .ZN(n6181) );
  NAND2_X1 U7317 ( .A1(n6182), .A2(n6181), .ZN(n6183) );
  AND2_X1 U7318 ( .A1(n6186), .A2(n6183), .ZN(n9175) );
  INV_X1 U7319 ( .A(n6186), .ZN(n9222) );
  INV_X1 U7320 ( .A(n6187), .ZN(n6188) );
  INV_X1 U7321 ( .A(SI_23_), .ZN(n10162) );
  MUX2_X1 U7322 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n6594), .Z(n6211) );
  INV_X1 U7323 ( .A(SI_24_), .ZN(n10177) );
  XNOR2_X1 U7324 ( .A(n6211), .B(n10177), .ZN(n6212) );
  XNOR2_X1 U7325 ( .A(n6213), .B(n6212), .ZN(n8177) );
  NAND2_X1 U7326 ( .A1(n8177), .A2(n9335), .ZN(n6192) );
  INV_X1 U7327 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8000) );
  OR2_X1 U7328 ( .A1(n9296), .A2(n8000), .ZN(n6191) );
  NAND2_X1 U7329 ( .A1(n9933), .A2(n5083), .ZN(n6202) );
  NAND2_X1 U7330 ( .A1(n6283), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6200) );
  INV_X1 U7331 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6193) );
  OR2_X1 U7332 ( .A1(n6446), .A2(n6193), .ZN(n6199) );
  INV_X1 U7333 ( .A(n6194), .ZN(n6196) );
  INV_X1 U7334 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9226) );
  INV_X1 U7335 ( .A(n6224), .ZN(n6195) );
  OAI21_X1 U7336 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n6196), .A(n6195), .ZN(
        n9747) );
  OR2_X1 U7337 ( .A1(n6337), .A2(n9747), .ZN(n6198) );
  INV_X1 U7338 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9748) );
  OR2_X1 U7339 ( .A1(n6448), .A2(n9748), .ZN(n6197) );
  NAND4_X1 U7340 ( .A1(n6200), .A2(n6199), .A3(n6198), .A4(n6197), .ZN(n9758)
         );
  NAND2_X1 U7341 ( .A1(n9758), .A2(n6282), .ZN(n6201) );
  NAND2_X1 U7342 ( .A1(n6202), .A2(n6201), .ZN(n6203) );
  XNOR2_X1 U7343 ( .A(n6203), .B(n5662), .ZN(n6205) );
  AND2_X1 U7344 ( .A1(n9758), .A2(n6247), .ZN(n6204) );
  AOI21_X1 U7345 ( .B1(n9933), .B2(n6282), .A(n6204), .ZN(n6206) );
  NAND2_X1 U7346 ( .A1(n6205), .A2(n6206), .ZN(n6210) );
  INV_X1 U7347 ( .A(n6205), .ZN(n6208) );
  INV_X1 U7348 ( .A(n6206), .ZN(n6207) );
  NAND2_X1 U7349 ( .A1(n6208), .A2(n6207), .ZN(n6209) );
  MUX2_X1 U7350 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n6594), .Z(n6214) );
  NAND2_X1 U7351 ( .A1(n6214), .A2(SI_25_), .ZN(n6232) );
  INV_X1 U7352 ( .A(n6214), .ZN(n6215) );
  INV_X1 U7353 ( .A(SI_25_), .ZN(n10163) );
  NAND2_X1 U7354 ( .A1(n6215), .A2(n10163), .ZN(n6216) );
  NAND2_X1 U7355 ( .A1(n6232), .A2(n6216), .ZN(n6219) );
  INV_X1 U7356 ( .A(n6219), .ZN(n6217) );
  NAND2_X1 U7357 ( .A1(n6218), .A2(n6217), .ZN(n6233) );
  NAND2_X1 U7358 ( .A1(n5457), .A2(n6219), .ZN(n6220) );
  NAND2_X1 U7359 ( .A1(n6233), .A2(n6220), .ZN(n8188) );
  OR2_X1 U7360 ( .A1(n8188), .A2(n5726), .ZN(n6222) );
  INV_X1 U7361 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7985) );
  NAND2_X1 U7362 ( .A1(n9735), .A2(n5083), .ZN(n6230) );
  NAND2_X1 U7363 ( .A1(n4932), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6228) );
  INV_X1 U7364 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10012) );
  OR2_X1 U7365 ( .A1(n6223), .A2(n10012), .ZN(n6227) );
  NAND2_X1 U7366 ( .A1(n6224), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6237) );
  OAI21_X1 U7367 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n6224), .A(n6237), .ZN(
        n9736) );
  OR2_X1 U7368 ( .A1(n6337), .A2(n9736), .ZN(n6226) );
  INV_X1 U7369 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9737) );
  OR2_X1 U7370 ( .A1(n6448), .A2(n9737), .ZN(n6225) );
  NAND4_X1 U7371 ( .A1(n6228), .A2(n6227), .A3(n6226), .A4(n6225), .ZN(n9642)
         );
  NAND2_X1 U7372 ( .A1(n9642), .A2(n6282), .ZN(n6229) );
  NAND2_X1 U7373 ( .A1(n6230), .A2(n6229), .ZN(n6231) );
  XNOR2_X1 U7374 ( .A(n6231), .B(n5633), .ZN(n6249) );
  AOI22_X1 U7375 ( .A1(n9735), .A2(n6282), .B1(n6247), .B2(n9642), .ZN(n6250)
         );
  XNOR2_X1 U7376 ( .A(n6249), .B(n6250), .ZN(n9198) );
  MUX2_X1 U7377 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n6594), .Z(n6253) );
  XNOR2_X1 U7378 ( .A(n6253), .B(SI_26_), .ZN(n6256) );
  XNOR2_X1 U7379 ( .A(n6257), .B(n6256), .ZN(n9157) );
  NAND2_X1 U7380 ( .A1(n9157), .A2(n9335), .ZN(n6236) );
  INV_X1 U7381 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n6234) );
  OR2_X1 U7382 ( .A1(n9296), .A2(n6234), .ZN(n6235) );
  NAND2_X1 U7383 ( .A1(n9724), .A2(n5083), .ZN(n6245) );
  NAND2_X1 U7384 ( .A1(n6283), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6243) );
  INV_X1 U7385 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9924) );
  OR2_X1 U7386 ( .A1(n6446), .A2(n9924), .ZN(n6242) );
  INV_X1 U7387 ( .A(n6237), .ZN(n6238) );
  NAND2_X1 U7388 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n6238), .ZN(n6263) );
  OAI21_X1 U7389 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n6238), .A(n6263), .ZN(
        n9717) );
  OR2_X1 U7390 ( .A1(n6337), .A2(n9717), .ZN(n6241) );
  INV_X1 U7391 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6239) );
  OR2_X1 U7392 ( .A1(n6448), .A2(n6239), .ZN(n6240) );
  NAND4_X1 U7393 ( .A1(n6243), .A2(n6242), .A3(n6241), .A4(n6240), .ZN(n9702)
         );
  NAND2_X1 U7394 ( .A1(n9702), .A2(n6282), .ZN(n6244) );
  NAND2_X1 U7395 ( .A1(n6245), .A2(n6244), .ZN(n6246) );
  XNOR2_X1 U7396 ( .A(n6246), .B(n5633), .ZN(n6274) );
  AND2_X1 U7397 ( .A1(n9702), .A2(n6247), .ZN(n6248) );
  AOI21_X1 U7398 ( .B1(n9724), .B2(n6282), .A(n6248), .ZN(n6272) );
  XNOR2_X1 U7399 ( .A(n6274), .B(n6272), .ZN(n9261) );
  INV_X1 U7400 ( .A(n6249), .ZN(n6251) );
  NAND2_X1 U7401 ( .A1(n6251), .A2(n6250), .ZN(n9262) );
  INV_X1 U7402 ( .A(n6253), .ZN(n6254) );
  NAND2_X1 U7403 ( .A1(n6254), .A2(n10170), .ZN(n6255) );
  MUX2_X1 U7404 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n6594), .Z(n6277) );
  INV_X1 U7405 ( .A(SI_27_), .ZN(n6278) );
  XNOR2_X1 U7406 ( .A(n6277), .B(n6278), .ZN(n6275) );
  NAND2_X1 U7407 ( .A1(n8265), .A2(n9335), .ZN(n6260) );
  INV_X1 U7408 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n6258) );
  OR2_X1 U7409 ( .A1(n9296), .A2(n6258), .ZN(n6259) );
  NAND2_X1 U7410 ( .A1(n6283), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6268) );
  INV_X1 U7411 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9917) );
  OR2_X1 U7412 ( .A1(n6446), .A2(n9917), .ZN(n6267) );
  INV_X1 U7413 ( .A(n6263), .ZN(n6261) );
  NAND2_X1 U7414 ( .A1(n6261), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6285) );
  INV_X1 U7415 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6262) );
  NAND2_X1 U7416 ( .A1(n6263), .A2(n6262), .ZN(n6264) );
  NAND2_X1 U7417 ( .A1(n6285), .A2(n6264), .ZN(n9694) );
  OR2_X1 U7418 ( .A1(n6337), .A2(n9694), .ZN(n6266) );
  INV_X1 U7419 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9695) );
  OR2_X1 U7420 ( .A1(n6448), .A2(n9695), .ZN(n6265) );
  NAND4_X1 U7421 ( .A1(n6268), .A2(n6267), .A3(n6266), .A4(n6265), .ZN(n9712)
         );
  AOI22_X1 U7422 ( .A1(n9693), .A2(n5083), .B1(n6282), .B2(n9712), .ZN(n6269)
         );
  XOR2_X1 U7423 ( .A(n5633), .B(n6269), .Z(n6271) );
  OAI22_X1 U7424 ( .A1(n9615), .A2(n5844), .B1(n9911), .B2(n6291), .ZN(n6270)
         );
  NOR2_X1 U7425 ( .A1(n6271), .A2(n6270), .ZN(n6325) );
  AOI21_X1 U7426 ( .B1(n6271), .B2(n6270), .A(n6325), .ZN(n6355) );
  INV_X1 U7427 ( .A(n6272), .ZN(n6273) );
  NAND2_X1 U7428 ( .A1(n6274), .A2(n6273), .ZN(n6356) );
  INV_X1 U7429 ( .A(n6277), .ZN(n6279) );
  MUX2_X1 U7430 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6594), .Z(n8222) );
  INV_X1 U7431 ( .A(SI_28_), .ZN(n10062) );
  XNOR2_X1 U7432 ( .A(n8222), .B(n10062), .ZN(n8220) );
  NAND2_X1 U7433 ( .A1(n8206), .A2(n9335), .ZN(n6281) );
  INV_X1 U7434 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10280) );
  OR2_X1 U7435 ( .A1(n9296), .A2(n10280), .ZN(n6280) );
  NAND2_X1 U7436 ( .A1(n9630), .A2(n6282), .ZN(n6293) );
  NAND2_X1 U7437 ( .A1(n6283), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6290) );
  INV_X1 U7438 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9913) );
  OR2_X1 U7439 ( .A1(n6446), .A2(n9913), .ZN(n6289) );
  INV_X1 U7440 ( .A(n6285), .ZN(n6284) );
  NAND2_X1 U7441 ( .A1(n6284), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9646) );
  INV_X1 U7442 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U7443 ( .A1(n6285), .A2(n6334), .ZN(n6286) );
  NAND2_X1 U7444 ( .A1(n9646), .A2(n6286), .ZN(n9674) );
  OR2_X1 U7445 ( .A1(n6337), .A2(n9674), .ZN(n6288) );
  INV_X1 U7446 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9675) );
  OR2_X1 U7447 ( .A1(n6448), .A2(n9675), .ZN(n6287) );
  OR2_X1 U7448 ( .A1(n9902), .A2(n6291), .ZN(n6292) );
  NAND2_X1 U7449 ( .A1(n6293), .A2(n6292), .ZN(n6294) );
  XNOR2_X1 U7450 ( .A(n6294), .B(n5662), .ZN(n6297) );
  NAND2_X1 U7451 ( .A1(n9630), .A2(n5083), .ZN(n6295) );
  OAI21_X1 U7452 ( .B1(n9902), .B2(n5844), .A(n6295), .ZN(n6296) );
  XNOR2_X1 U7453 ( .A(n6297), .B(n6296), .ZN(n6324) );
  INV_X1 U7454 ( .A(P1_B_REG_SCAN_IN), .ZN(n9617) );
  NAND2_X1 U7455 ( .A1(n6298), .A2(n9617), .ZN(n6301) );
  NAND3_X1 U7456 ( .A1(n5603), .A2(P1_B_REG_SCAN_IN), .A3(n6299), .ZN(n6300)
         );
  INV_X1 U7457 ( .A(n6302), .ZN(n10287) );
  NAND2_X1 U7458 ( .A1(n10287), .A2(n5603), .ZN(n10045) );
  OR2_X1 U7459 ( .A1(n10042), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6304) );
  NAND2_X1 U7460 ( .A1(n10287), .A2(n6299), .ZN(n10044) );
  NOR4_X1 U7461 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6313) );
  NOR4_X1 U7462 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6312) );
  OR4_X1 U7463 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6310) );
  NOR4_X1 U7464 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6308) );
  NOR4_X1 U7465 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6307) );
  NOR4_X1 U7466 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6306) );
  NOR4_X1 U7467 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6305) );
  NAND4_X1 U7468 ( .A1(n6308), .A2(n6307), .A3(n6306), .A4(n6305), .ZN(n6309)
         );
  NOR4_X1 U7469 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n6310), .A4(n6309), .ZN(n6311) );
  AND3_X1 U7470 ( .A1(n6313), .A2(n6312), .A3(n6311), .ZN(n6314) );
  OR2_X1 U7471 ( .A1(n10042), .A2(n6314), .ZN(n7218) );
  NAND3_X1 U7472 ( .A1(n7224), .A2(n7340), .A3(n7218), .ZN(n6345) );
  NOR2_X1 U7473 ( .A1(n6345), .A2(n10041), .ZN(n6330) );
  NAND2_X1 U7474 ( .A1(n6319), .A2(n5609), .ZN(n9522) );
  AND2_X1 U7475 ( .A1(n10729), .A2(n9522), .ZN(n6343) );
  INV_X1 U7476 ( .A(n6324), .ZN(n6322) );
  INV_X1 U7477 ( .A(n6325), .ZN(n6321) );
  NAND3_X1 U7478 ( .A1(n6323), .A2(n6322), .A3(n5552), .ZN(n6353) );
  NAND3_X1 U7479 ( .A1(n6325), .A2(n6324), .A3(n9259), .ZN(n6352) );
  INV_X1 U7480 ( .A(n6330), .ZN(n6327) );
  INV_X1 U7481 ( .A(n7744), .ZN(n9544) );
  OR2_X1 U7482 ( .A1(n10041), .A2(n9544), .ZN(n6326) );
  NAND2_X1 U7483 ( .A1(n6327), .A2(n6326), .ZN(n7261) );
  INV_X1 U7484 ( .A(n7198), .ZN(n6329) );
  AND2_X1 U7485 ( .A1(n6329), .A2(n6328), .ZN(n10518) );
  NAND2_X1 U7486 ( .A1(n6330), .A2(n10518), .ZN(n6335) );
  NAND2_X1 U7487 ( .A1(n6332), .A2(n6331), .ZN(n6639) );
  NAND2_X1 U7488 ( .A1(n6639), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6333) );
  INV_X1 U7489 ( .A(n10347), .ZN(n10282) );
  OR2_X2 U7490 ( .A1(n6335), .A2(n10282), .ZN(n9278) );
  OAI22_X1 U7491 ( .A1(n9278), .A2(n9911), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6334), .ZN(n6350) );
  NAND2_X1 U7492 ( .A1(n5671), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6341) );
  INV_X1 U7493 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6336) );
  OR2_X1 U7494 ( .A1(n6446), .A2(n6336), .ZN(n6340) );
  OR2_X1 U7495 ( .A1(n6337), .A2(n9646), .ZN(n6339) );
  INV_X1 U7496 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9647) );
  OR2_X1 U7497 ( .A1(n6448), .A2(n9647), .ZN(n6338) );
  INV_X1 U7498 ( .A(n10518), .ZN(n6342) );
  OR2_X1 U7499 ( .A1(n6342), .A2(n10041), .ZN(n9287) );
  INV_X1 U7500 ( .A(n6343), .ZN(n6344) );
  NAND2_X1 U7501 ( .A1(n10532), .A2(n9544), .ZN(n7349) );
  NAND3_X1 U7502 ( .A1(n9287), .A2(n6344), .A3(n7349), .ZN(n6346) );
  NAND2_X1 U7503 ( .A1(n6346), .A2(n6345), .ZN(n6348) );
  NAND2_X1 U7504 ( .A1(n9526), .A2(n7197), .ZN(n7219) );
  AND3_X1 U7505 ( .A1(n7219), .A2(n7814), .A3(n6363), .ZN(n6347) );
  NAND2_X1 U7506 ( .A1(n6348), .A2(n6347), .ZN(n6694) );
  OAI22_X1 U7507 ( .A1(n9276), .A2(n9682), .B1(n9275), .B2(n9674), .ZN(n6349)
         );
  AOI211_X1 U7508 ( .C1(n9630), .C2(n9281), .A(n6350), .B(n6349), .ZN(n6351)
         );
  NAND4_X1 U7509 ( .A1(n6354), .A2(n6353), .A3(n6352), .A4(n6351), .ZN(
        P1_U3220) );
  AOI21_X1 U7510 ( .B1(n9260), .B2(n6356), .A(n6355), .ZN(n6357) );
  NOR2_X1 U7511 ( .A1(n9278), .A2(n9730), .ZN(n6360) );
  OAI22_X1 U7512 ( .A1(n9276), .A2(n9902), .B1(n9275), .B2(n9694), .ZN(n6359)
         );
  AOI211_X1 U7513 ( .C1(P1_REG3_REG_27__SCAN_IN), .C2(P1_U3086), .A(n6360), 
        .B(n6359), .ZN(n6362) );
  NAND2_X1 U7514 ( .A1(n9693), .A2(n9281), .ZN(n6361) );
  NOR2_X1 U7515 ( .A1(n6363), .A2(P1_U3086), .ZN(n6364) );
  AND4_X2 U7516 ( .A1(n6366), .A2(n6365), .A3(n6583), .A4(n6456), .ZN(n6368)
         );
  AND4_X2 U7517 ( .A1(n6454), .A2(n6396), .A3(n6455), .A4(n6394), .ZN(n6367)
         );
  NAND3_X1 U7518 ( .A1(n6548), .A2(n6412), .A3(n6414), .ZN(n6416) );
  INV_X1 U7519 ( .A(n7956), .ZN(n6381) );
  NAND2_X1 U7520 ( .A1(n6387), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6378) );
  INV_X1 U7521 ( .A(n7957), .ZN(n6380) );
  OR2_X1 U7522 ( .A1(n6383), .A2(n6384), .ZN(n6385) );
  NAND2_X1 U7523 ( .A1(n6385), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6386) );
  MUX2_X1 U7524 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6386), .S(
        P2_IR_REG_23__SCAN_IN), .Z(n6388) );
  NAND2_X1 U7525 ( .A1(n6388), .A2(n6387), .ZN(n6852) );
  INV_X2 U7526 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NAND2_X1 U7527 ( .A1(n8278), .A2(P2_U3151), .ZN(n8267) );
  INV_X1 U7528 ( .A(n7817), .ZN(n9159) );
  NOR2_X1 U7529 ( .A1(n8278), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9150) );
  OAI222_X1 U7530 ( .A1(n9159), .A2(n6742), .B1(n9156), .B2(n5305), .C1(
        P2_U3151), .C2(n4931), .ZN(P2_U3293) );
  INV_X1 U7531 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U7532 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6392) );
  OAI222_X1 U7533 ( .A1(n9159), .A2(n6593), .B1(n9156), .B2(n5638), .C1(
        P2_U3151), .C2(n6612), .ZN(P2_U3294) );
  OAI222_X1 U7534 ( .A1(n9156), .A2(n5220), .B1(n6934), .B2(P2_U3151), .C1(
        n9159), .C2(n6858), .ZN(P2_U3292) );
  INV_X1 U7535 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7005) );
  NAND2_X1 U7536 ( .A1(n6395), .A2(n6394), .ZN(n6402) );
  NAND2_X1 U7537 ( .A1(n6402), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6397) );
  OAI222_X1 U7538 ( .A1(n9156), .A2(n7005), .B1(n7064), .B2(P2_U3151), .C1(
        n9159), .C2(n7006), .ZN(P2_U3291) );
  NAND2_X1 U7539 ( .A1(n8278), .A2(P1_U3086), .ZN(n10285) );
  INV_X1 U7540 ( .A(n10285), .ZN(n10053) );
  NOR2_X1 U7541 ( .A1(n8278), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10054) );
  INV_X2 U7542 ( .A(n10054), .ZN(n8002) );
  OAI222_X1 U7543 ( .A1(n10284), .A2(n6398), .B1(n8002), .B2(n7006), .C1(n6918), .C2(P1_U3086), .ZN(P1_U3351) );
  OAI222_X1 U7544 ( .A1(P1_U3086), .A2(n6725), .B1(n8002), .B2(n6593), .C1(
        n6399), .C2(n10284), .ZN(P1_U3354) );
  OAI222_X1 U7545 ( .A1(P1_U3086), .A2(n6961), .B1(n8002), .B2(n6742), .C1(
        n6400), .C2(n10284), .ZN(P1_U3353) );
  OAI222_X1 U7546 ( .A1(P1_U3086), .A2(n6401), .B1(n8002), .B2(n6858), .C1(
        n5219), .C2(n10284), .ZN(P1_U3352) );
  INV_X1 U7547 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U7548 ( .A1(n6406), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6404) );
  INV_X1 U7549 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6403) );
  XNOR2_X1 U7550 ( .A(n6404), .B(n6403), .ZN(n7177) );
  OAI222_X1 U7551 ( .A1(n9159), .A2(n7126), .B1(n9156), .B2(n6473), .C1(
        P2_U3151), .C2(n7177), .ZN(P2_U3290) );
  OAI222_X1 U7552 ( .A1(n10284), .A2(n6405), .B1(n8002), .B2(n7126), .C1(n6665), .C2(P1_U3086), .ZN(P1_U3350) );
  NOR2_X1 U7553 ( .A1(n6406), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n6458) );
  OR2_X1 U7554 ( .A1(n6458), .A2(n9147), .ZN(n6421) );
  XNOR2_X1 U7555 ( .A(n6421), .B(n6455), .ZN(n7326) );
  INV_X1 U7556 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7236) );
  OAI222_X1 U7557 ( .A1(n9159), .A2(n7235), .B1(n7326), .B2(P2_U3151), .C1(
        n7236), .C2(n9156), .ZN(P2_U3289) );
  OAI222_X1 U7558 ( .A1(n10284), .A2(n6407), .B1(n8002), .B2(n7235), .C1(n6784), .C2(P1_U3086), .ZN(P1_U3349) );
  INV_X1 U7559 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6409) );
  NAND2_X1 U7560 ( .A1(n6383), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U7561 ( .A1(n6552), .A2(n6412), .ZN(n6413) );
  OR2_X1 U7562 ( .A1(n6383), .A2(n6416), .ZN(n6417) );
  NAND2_X1 U7563 ( .A1(n6417), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6418) );
  NAND2_X1 U7564 ( .A1(n6494), .A2(n8491), .ZN(n6419) );
  NAND2_X1 U7565 ( .A1(n6419), .A2(n6852), .ZN(n6486) );
  INV_X1 U7566 ( .A(n6486), .ZN(n6420) );
  OAI21_X1 U7567 ( .B1(n8131), .B2(n6420), .A(P2_STATE_REG_SCAN_IN), .ZN(
        P2_U3150) );
  AOI21_X1 U7568 ( .B1(n6421), .B2(n6455), .A(n9147), .ZN(n6422) );
  NAND2_X1 U7569 ( .A1(n6422), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n6424) );
  INV_X1 U7570 ( .A(n6422), .ZN(n6423) );
  NAND2_X1 U7571 ( .A1(n6423), .A2(n6456), .ZN(n6435) );
  NAND2_X1 U7572 ( .A1(n6424), .A2(n6435), .ZN(n7393) );
  INV_X1 U7573 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7365) );
  OAI222_X1 U7574 ( .A1(n9159), .A2(n7364), .B1(n7393), .B2(P2_U3151), .C1(
        n7365), .C2(n9156), .ZN(P2_U3288) );
  INV_X1 U7575 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6425) );
  INV_X1 U7576 ( .A(n6705), .ZN(n6671) );
  OAI222_X1 U7577 ( .A1(n10285), .A2(n6425), .B1(n8002), .B2(n7364), .C1(n6671), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U7578 ( .A(n6577), .ZN(n6847) );
  XNOR2_X1 U7579 ( .A(n7957), .B(P2_B_REG_SCAN_IN), .ZN(n6426) );
  NAND2_X1 U7580 ( .A1(n6426), .A2(n7956), .ZN(n6427) );
  INV_X1 U7581 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6430) );
  INV_X1 U7582 ( .A(n6428), .ZN(n9158) );
  NAND2_X1 U7583 ( .A1(n9158), .A2(n7957), .ZN(n6534) );
  INV_X1 U7584 ( .A(n6534), .ZN(n6429) );
  AOI22_X1 U7585 ( .A1(n6433), .A2(n6430), .B1(n6566), .B2(n6429), .ZN(
        P2_U3376) );
  INV_X1 U7586 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6432) );
  NAND2_X1 U7587 ( .A1(n9158), .A2(n7956), .ZN(n6532) );
  INV_X1 U7588 ( .A(n6532), .ZN(n6431) );
  AOI22_X1 U7589 ( .A1(n6433), .A2(n6432), .B1(n6566), .B2(n6431), .ZN(
        P2_U3377) );
  AND2_X1 U7590 ( .A1(n6433), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U7591 ( .A1(n6433), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U7592 ( .A1(n6433), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U7593 ( .A1(n6433), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U7594 ( .A1(n6433), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U7595 ( .A1(n6433), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U7596 ( .A1(n6433), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U7597 ( .A1(n6433), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U7598 ( .A1(n6433), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U7599 ( .A1(n6433), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U7600 ( .A1(n6433), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U7601 ( .A1(n6433), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U7602 ( .A1(n6433), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U7603 ( .A1(n6433), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U7604 ( .A1(n6433), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U7605 ( .A1(n6433), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U7606 ( .A1(n6433), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U7607 ( .A1(n6433), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U7608 ( .A1(n6433), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U7609 ( .A1(n6433), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U7610 ( .A1(n6433), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U7611 ( .A1(n6433), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U7612 ( .A1(n6433), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U7613 ( .A1(n6433), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U7614 ( .A1(n6433), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U7615 ( .A1(n6433), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U7616 ( .A1(n6433), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U7617 ( .A1(n6433), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U7618 ( .A1(n6433), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U7619 ( .A1(n6433), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U7620 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6434) );
  INV_X1 U7621 ( .A(n7570), .ZN(n6437) );
  INV_X1 U7622 ( .A(n6706), .ZN(n6794) );
  OAI222_X1 U7623 ( .A1(n10284), .A2(n6434), .B1(n8002), .B2(n6437), .C1(
        P1_U3086), .C2(n6794), .ZN(P1_U3347) );
  INV_X1 U7624 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6438) );
  NAND2_X1 U7625 ( .A1(n6435), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6436) );
  INV_X1 U7626 ( .A(n7571), .ZN(n7537) );
  OAI222_X1 U7627 ( .A1(n9156), .A2(n6438), .B1(n9159), .B2(n6437), .C1(
        P2_U3151), .C2(n7537), .ZN(P2_U3287) );
  NAND2_X1 U7628 ( .A1(n7814), .A2(n6439), .ZN(n6440) );
  NAND2_X1 U7629 ( .A1(n6440), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6636) );
  INV_X1 U7630 ( .A(n6636), .ZN(n6442) );
  NAND2_X1 U7631 ( .A1(n9526), .A2(n7814), .ZN(n6441) );
  NAND2_X1 U7632 ( .A1(n6441), .A2(n5086), .ZN(n6637) );
  NOR2_X1 U7633 ( .A1(n10350), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U7634 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8509) );
  INV_X1 U7635 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9900) );
  INV_X1 U7636 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9625) );
  OR2_X1 U7637 ( .A1(n6448), .A2(n9625), .ZN(n6444) );
  NAND2_X1 U7638 ( .A1(n5671), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6443) );
  OAI211_X1 U7639 ( .C1(n6446), .C2(n9900), .A(n6444), .B(n6443), .ZN(n9666)
         );
  NAND2_X1 U7640 ( .A1(n9666), .A2(P1_U3973), .ZN(n6445) );
  OAI21_X1 U7641 ( .B1(n8509), .B2(P1_U3973), .A(n6445), .ZN(P1_U3584) );
  INV_X1 U7642 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6453) );
  NAND2_X1 U7643 ( .A1(n5671), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6451) );
  INV_X1 U7644 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9896) );
  OR2_X1 U7645 ( .A1(n6446), .A2(n9896), .ZN(n6450) );
  INV_X1 U7646 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6447) );
  OR2_X1 U7647 ( .A1(n6448), .A2(n6447), .ZN(n6449) );
  INV_X1 U7648 ( .A(n9620), .ZN(n9525) );
  NAND2_X1 U7649 ( .A1(n9525), .A2(P1_U3973), .ZN(n6452) );
  OAI21_X1 U7650 ( .B1(P1_U3973), .B2(n6453), .A(n6452), .ZN(P1_U3585) );
  AND3_X1 U7651 ( .A1(n6456), .A2(n6455), .A3(n6454), .ZN(n6457) );
  AND2_X1 U7652 ( .A1(n6458), .A2(n6457), .ZN(n6461) );
  NAND2_X1 U7653 ( .A1(n6461), .A2(n6462), .ZN(n6581) );
  NAND2_X1 U7654 ( .A1(n6581), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6459) );
  XNOR2_X1 U7655 ( .A(n6459), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8745) );
  INV_X1 U7656 ( .A(n8745), .ZN(n8731) );
  INV_X1 U7657 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6460) );
  OAI222_X1 U7658 ( .A1(n7761), .A2(n9159), .B1(n8731), .B2(P2_U3151), .C1(
        n6460), .C2(n9156), .ZN(P2_U3285) );
  INV_X1 U7659 ( .A(n7580), .ZN(n6470) );
  OR2_X1 U7660 ( .A1(n6461), .A2(n9147), .ZN(n6463) );
  XNOR2_X1 U7661 ( .A(n6463), .B(n6462), .ZN(n8742) );
  INV_X1 U7662 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6464) );
  OAI222_X1 U7663 ( .A1(n8267), .A2(n6470), .B1(n8742), .B2(P2_U3151), .C1(
        n6464), .C2(n9156), .ZN(P2_U3286) );
  INV_X1 U7664 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6465) );
  INV_X1 U7665 ( .A(n6886), .ZN(n6891) );
  OAI222_X1 U7666 ( .A1(n10285), .A2(n6465), .B1(n8002), .B2(n7761), .C1(n6891), .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U7667 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6797) );
  NAND2_X1 U7668 ( .A1(n7964), .A2(P1_U3973), .ZN(n6466) );
  OAI21_X1 U7669 ( .B1(n6797), .B2(P1_U3973), .A(n6466), .ZN(P1_U3567) );
  INV_X1 U7670 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7271) );
  NAND2_X1 U7671 ( .A1(n9851), .A2(P1_U3973), .ZN(n6467) );
  OAI21_X1 U7672 ( .B1(n7271), .B2(P1_U3973), .A(n6467), .ZN(P1_U3572) );
  NAND2_X1 U7673 ( .A1(n5664), .A2(P1_U3973), .ZN(n6468) );
  OAI21_X1 U7674 ( .B1(P1_U3973), .B2(n5638), .A(n6468), .ZN(P1_U3555) );
  NAND2_X1 U7675 ( .A1(n5692), .A2(P1_U3973), .ZN(n6469) );
  OAI21_X1 U7676 ( .B1(P1_U3973), .B2(n5305), .A(n6469), .ZN(P1_U3556) );
  INV_X1 U7677 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6471) );
  INV_X1 U7678 ( .A(n6728), .ZN(n6732) );
  OAI222_X1 U7679 ( .A1(n10285), .A2(n6471), .B1(n8002), .B2(n6470), .C1(n6732), .C2(P1_U3086), .ZN(P1_U3346) );
  NAND2_X1 U7680 ( .A1(n7514), .A2(P1_U3973), .ZN(n6472) );
  OAI21_X1 U7681 ( .B1(P1_U3973), .B2(n6473), .A(n6472), .ZN(P1_U3559) );
  NAND2_X1 U7682 ( .A1(n6474), .A2(P1_U3973), .ZN(n6475) );
  OAI21_X1 U7683 ( .B1(P1_U3973), .B2(n5642), .A(n6475), .ZN(P1_U3554) );
  INV_X1 U7684 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U7685 ( .A1(n9639), .A2(P1_U3973), .ZN(n6476) );
  OAI21_X1 U7686 ( .B1(P1_U3973), .B2(n6477), .A(n6476), .ZN(P1_U3577) );
  MUX2_X1 U7687 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8825), .Z(n6675) );
  XNOR2_X1 U7688 ( .A(n6675), .B(n4931), .ZN(n6485) );
  INV_X1 U7689 ( .A(n6572), .ZN(n6479) );
  MUX2_X1 U7690 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n6479), .Z(n6481) );
  XNOR2_X1 U7691 ( .A(n6481), .B(n6612), .ZN(n6624) );
  INV_X1 U7692 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6480) );
  INV_X1 U7693 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6816) );
  MUX2_X1 U7694 ( .A(n6480), .B(n6816), .S(n6479), .Z(n6512) );
  AND2_X1 U7695 ( .A1(n6512), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6623) );
  NOR2_X1 U7696 ( .A1(n6624), .A2(n6623), .ZN(n6622) );
  AOI21_X1 U7697 ( .B1(n6481), .B2(n6612), .A(n6622), .ZN(n6484) );
  NAND2_X1 U7698 ( .A1(P2_U3893), .A2(n6483), .ZN(n8830) );
  NOR2_X1 U7699 ( .A1(n6484), .A2(n6485), .ZN(n6674) );
  AOI211_X1 U7700 ( .C1(n6485), .C2(n6484), .A(n8830), .B(n6674), .ZN(n6511)
         );
  NAND2_X1 U7701 ( .A1(n6486), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6488) );
  MUX2_X1 U7702 ( .A(n10503), .B(n6488), .S(n6483), .Z(n6487) );
  NOR2_X2 U7703 ( .A1(n6487), .A2(n8131), .ZN(n10476) );
  INV_X1 U7704 ( .A(n10476), .ZN(n10502) );
  OR2_X1 U7705 ( .A1(n6488), .A2(n6483), .ZN(n6513) );
  INV_X1 U7706 ( .A(n10489), .ZN(n10509) );
  INV_X1 U7707 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10579) );
  MUX2_X1 U7708 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10579), .S(n6746), .Z(n6492)
         );
  INV_X1 U7709 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6518) );
  AND2_X1 U7710 ( .A1(n6518), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6489) );
  OAI21_X1 U7711 ( .B1(n6612), .B2(n6489), .A(n6490), .ZN(n6615) );
  INV_X1 U7712 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6616) );
  OR2_X1 U7713 ( .A1(n6615), .A2(n6616), .ZN(n6613) );
  NAND2_X1 U7714 ( .A1(n6613), .A2(n6490), .ZN(n6491) );
  OAI21_X1 U7715 ( .B1(n6492), .B2(n6491), .A(n6685), .ZN(n6499) );
  NAND2_X1 U7716 ( .A1(n8492), .A2(n6852), .ZN(n6493) );
  NAND2_X1 U7717 ( .A1(n8249), .A2(n6493), .ZN(n6496) );
  INV_X1 U7718 ( .A(n6494), .ZN(n6556) );
  AOI21_X1 U7719 ( .B1(n6556), .B2(n6852), .A(P2_U3151), .ZN(n6495) );
  INV_X1 U7720 ( .A(n10498), .ZN(n8738) );
  INV_X1 U7721 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6497) );
  OAI22_X1 U7722 ( .A1(n8738), .A2(n6497), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10263), .ZN(n6498) );
  AOI21_X1 U7723 ( .B1(n10509), .B2(n6499), .A(n6498), .ZN(n6509) );
  INV_X1 U7724 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6500) );
  MUX2_X1 U7725 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6500), .S(n4931), .Z(n6506)
         );
  NAND2_X1 U7726 ( .A1(n6612), .A2(n6503), .ZN(n6502) );
  NAND2_X1 U7727 ( .A1(n6502), .A2(n6501), .ZN(n6617) );
  NAND2_X1 U7728 ( .A1(n6617), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U7729 ( .A1(n6504), .A2(n6503), .ZN(n6505) );
  NAND2_X1 U7730 ( .A1(n6506), .A2(n6505), .ZN(n6680) );
  OAI21_X1 U7731 ( .B1(n6506), .B2(n6505), .A(n6680), .ZN(n6507) );
  NAND2_X1 U7732 ( .A1(n10483), .A2(n6507), .ZN(n6508) );
  OAI211_X1 U7733 ( .C1(n10502), .C2(n4931), .A(n6509), .B(n6508), .ZN(n6510)
         );
  OR2_X1 U7734 ( .A1(n6511), .A2(n6510), .ZN(P2_U3184) );
  AOI22_X1 U7735 ( .A1(n10498), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n6517) );
  NOR2_X1 U7736 ( .A1(n6512), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6515) );
  INV_X1 U7737 ( .A(n6513), .ZN(n6514) );
  OAI22_X1 U7738 ( .A1(n6623), .A2(n6515), .B1(n6514), .B2(n10513), .ZN(n6516)
         );
  OAI211_X1 U7739 ( .C1(n10502), .C2(n6518), .A(n6517), .B(n6516), .ZN(
        P2_U3182) );
  NAND2_X1 U7740 ( .A1(n6522), .A2(n6519), .ZN(n9148) );
  XNOR2_X2 U7741 ( .A(n6521), .B(n6520), .ZN(n8508) );
  INV_X1 U7742 ( .A(n8508), .ZN(n6525) );
  INV_X1 U7743 ( .A(n6522), .ZN(n6523) );
  NAND2_X1 U7744 ( .A1(n6865), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6530) );
  NAND2_X1 U7745 ( .A1(n8160), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U7746 ( .A1(n6864), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U7747 ( .A1(n6990), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6527) );
  NAND2_X1 U7748 ( .A1(n8278), .A2(SI_0_), .ZN(n6531) );
  XNOR2_X1 U7749 ( .A(n6531), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9161) );
  MUX2_X1 U7750 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9161), .S(n8249), .Z(n6805) );
  INV_X1 U7751 ( .A(n6805), .ZN(n6823) );
  AND2_X1 U7752 ( .A1(n8717), .A2(n6823), .ZN(n8341) );
  NOR2_X1 U7753 ( .A1(n8717), .A2(n6823), .ZN(n8345) );
  OR2_X1 U7754 ( .A1(n8341), .A2(n8345), .ZN(n8339) );
  INV_X1 U7755 ( .A(n8339), .ZN(n8311) );
  INV_X1 U7756 ( .A(n6819), .ZN(n6535) );
  NOR2_X1 U7757 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6539) );
  NOR4_X1 U7758 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6538) );
  NOR4_X1 U7759 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6537) );
  NOR4_X1 U7760 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6536) );
  NAND4_X1 U7761 ( .A1(n6539), .A2(n6538), .A3(n6537), .A4(n6536), .ZN(n6545)
         );
  NOR4_X1 U7762 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6543) );
  NOR4_X1 U7763 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6542) );
  NOR4_X1 U7764 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6541) );
  NOR4_X1 U7765 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6540) );
  NAND4_X1 U7766 ( .A1(n6543), .A2(n6542), .A3(n6541), .A4(n6540), .ZN(n6544)
         );
  NOR2_X1 U7767 ( .A1(n6545), .A2(n6544), .ZN(n6546) );
  NAND2_X1 U7768 ( .A1(n6808), .A2(n6806), .ZN(n6846) );
  NAND2_X1 U7769 ( .A1(n8491), .A2(n10715), .ZN(n6559) );
  OR2_X1 U7770 ( .A1(n6549), .A2(n6548), .ZN(n6550) );
  INV_X1 U7771 ( .A(n7691), .ZN(n8336) );
  AND3_X1 U7772 ( .A1(n8336), .A2(n8505), .A3(n8833), .ZN(n6553) );
  AND2_X1 U7773 ( .A1(n6553), .A2(n7674), .ZN(n6839) );
  OR2_X1 U7774 ( .A1(n6559), .A2(n6839), .ZN(n6555) );
  NAND2_X1 U7775 ( .A1(n7691), .A2(n8833), .ZN(n6995) );
  INV_X1 U7776 ( .A(n6995), .ZN(n6554) );
  NAND2_X1 U7777 ( .A1(n6555), .A2(n10571), .ZN(n6842) );
  NAND2_X1 U7778 ( .A1(n6846), .A2(n6842), .ZN(n6558) );
  NAND3_X1 U7779 ( .A1(n6819), .A2(n5332), .A3(n6806), .ZN(n6843) );
  AOI21_X1 U7780 ( .B1(n6843), .B2(n6839), .A(n6556), .ZN(n6557) );
  AND2_X1 U7781 ( .A1(n6558), .A2(n6557), .ZN(n6564) );
  INV_X1 U7782 ( .A(n6564), .ZN(n6562) );
  OR2_X1 U7783 ( .A1(n6560), .A2(n6559), .ZN(n6561) );
  INV_X1 U7784 ( .A(n8833), .ZN(n7418) );
  NAND2_X1 U7785 ( .A1(n7691), .A2(n7418), .ZN(n6801) );
  OR2_X1 U7786 ( .A1(n6577), .A2(n6840), .ZN(n6571) );
  INV_X1 U7787 ( .A(n6571), .ZN(n8503) );
  INV_X1 U7788 ( .A(n6801), .ZN(n6563) );
  AOI21_X1 U7789 ( .B1(n6564), .B2(n6813), .A(P2_U3151), .ZN(n6565) );
  AOI21_X1 U7790 ( .B1(n8503), .B2(n6843), .A(n6565), .ZN(n6854) );
  NAND2_X1 U7791 ( .A1(n6854), .A2(n6566), .ZN(n6758) );
  NAND2_X1 U7792 ( .A1(n6758), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6580) );
  NAND2_X1 U7793 ( .A1(n6865), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6570) );
  NAND2_X1 U7794 ( .A1(n6864), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6569) );
  NAND2_X1 U7795 ( .A1(n6990), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6568) );
  NAND2_X1 U7796 ( .A1(n8160), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6567) );
  NOR2_X1 U7797 ( .A1(n6843), .A2(n6571), .ZN(n6604) );
  INV_X1 U7798 ( .A(n6604), .ZN(n6574) );
  INV_X1 U7799 ( .A(n6483), .ZN(n8502) );
  NAND2_X1 U7800 ( .A1(n8502), .A2(n6572), .ZN(n6573) );
  INV_X1 U7801 ( .A(n6846), .ZN(n6576) );
  NOR2_X1 U7802 ( .A1(n6577), .A2(n10715), .ZN(n6575) );
  NAND2_X1 U7803 ( .A1(n6576), .A2(n6575), .ZN(n6578) );
  OR2_X1 U7804 ( .A1(n10715), .A2(n6995), .ZN(n6809) );
  AOI22_X1 U7805 ( .A1(n6942), .A2(n8689), .B1(n6805), .B2(n8681), .ZN(n6579)
         );
  OAI211_X1 U7806 ( .C1(n8311), .C2(n8683), .A(n6580), .B(n6579), .ZN(P2_U3172) );
  INV_X1 U7807 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6586) );
  INV_X1 U7808 ( .A(n7836), .ZN(n6587) );
  NAND2_X1 U7809 ( .A1(n6582), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6584) );
  OR2_X1 U7810 ( .A1(n6584), .A2(n6583), .ZN(n6585) );
  NAND2_X1 U7811 ( .A1(n6584), .A2(n6583), .ZN(n6609) );
  INV_X1 U7812 ( .A(n10371), .ZN(n8808) );
  OAI222_X1 U7813 ( .A1(n9156), .A2(n6586), .B1(n9159), .B2(n6587), .C1(
        P2_U3151), .C2(n8808), .ZN(P2_U3284) );
  INV_X1 U7814 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6588) );
  INV_X1 U7815 ( .A(n7157), .ZN(n7161) );
  OAI222_X1 U7816 ( .A1(n10285), .A2(n6588), .B1(n8002), .B2(n6587), .C1(
        P1_U3086), .C2(n7161), .ZN(P1_U3344) );
  AND2_X1 U7817 ( .A1(n7674), .A2(n6995), .ZN(n6589) );
  NAND2_X1 U7818 ( .A1(n6810), .A2(n6589), .ZN(n6591) );
  NAND2_X1 U7819 ( .A1(n8344), .A2(n7691), .ZN(n6590) );
  NAND2_X1 U7820 ( .A1(n8717), .A2(n6805), .ZN(n6947) );
  OAI21_X1 U7821 ( .B1(n6805), .B2(n6592), .A(n6947), .ZN(n6599) );
  OR2_X1 U7822 ( .A1(n6741), .A2(n6593), .ZN(n6596) );
  NAND2_X1 U7823 ( .A1(n8249), .A2(n6594), .ZN(n6743) );
  OR2_X1 U7824 ( .A1(n6743), .A2(n5638), .ZN(n6595) );
  OAI211_X2 U7825 ( .C1(n8249), .C2(n6612), .A(n6596), .B(n6595), .ZN(n6997)
         );
  NAND2_X1 U7826 ( .A1(n6597), .A2(n10563), .ZN(n6747) );
  OAI21_X1 U7827 ( .B1(n10563), .B2(n6597), .A(n6747), .ZN(n6598) );
  AOI21_X1 U7828 ( .B1(n6599), .B2(n6598), .A(n6749), .ZN(n6608) );
  NAND2_X1 U7829 ( .A1(n6990), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U7830 ( .A1(n6865), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6602) );
  NAND2_X1 U7831 ( .A1(n8160), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6601) );
  NAND2_X1 U7832 ( .A1(n6864), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6600) );
  AOI22_X1 U7833 ( .A1(n8717), .A2(n8676), .B1(n8681), .B2(n6997), .ZN(n6605)
         );
  OAI21_X1 U7834 ( .B1(n7081), .B2(n8679), .A(n6605), .ZN(n6606) );
  AOI21_X1 U7835 ( .B1(n6758), .B2(P2_REG3_REG_1__SCAN_IN), .A(n6606), .ZN(
        n6607) );
  OAI21_X1 U7836 ( .B1(n6608), .B2(n8683), .A(n6607), .ZN(P2_U3162) );
  NAND2_X1 U7837 ( .A1(n6609), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6610) );
  INV_X1 U7838 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6611) );
  OAI222_X1 U7839 ( .A1(n8267), .A2(n7927), .B1(n8804), .B2(P2_U3151), .C1(
        n6611), .C2(n9156), .ZN(P2_U3283) );
  INV_X1 U7840 ( .A(n6612), .ZN(n6627) );
  INV_X1 U7841 ( .A(n6613), .ZN(n6614) );
  AOI21_X1 U7842 ( .B1(n6616), .B2(n6615), .A(n6614), .ZN(n6621) );
  AOI22_X1 U7843 ( .A1(n10498), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3151), .ZN(n6620) );
  XNOR2_X1 U7844 ( .A(n6617), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n6618) );
  NAND2_X1 U7845 ( .A1(n10483), .A2(n6618), .ZN(n6619) );
  OAI211_X1 U7846 ( .C1(n6621), .C2(n10489), .A(n6620), .B(n6619), .ZN(n6626)
         );
  AOI211_X1 U7847 ( .C1(n6624), .C2(n6623), .A(n8830), .B(n6622), .ZN(n6625)
         );
  AOI211_X1 U7848 ( .C1(n10476), .C2(n6627), .A(n6626), .B(n6625), .ZN(n6628)
         );
  INV_X1 U7849 ( .A(n6628), .ZN(P2_U3183) );
  INV_X1 U7850 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6629) );
  INV_X1 U7851 ( .A(n7162), .ZN(n10361) );
  OAI222_X1 U7852 ( .A1(n10285), .A2(n6629), .B1(n8002), .B2(n7927), .C1(
        n10361), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U7853 ( .A(n6961), .ZN(n6630) );
  NAND2_X1 U7854 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6716) );
  NOR2_X1 U7855 ( .A1(n6717), .A2(n6716), .ZN(n6715) );
  AOI21_X1 U7856 ( .B1(n6644), .B2(P1_REG2_REG_1__SCAN_IN), .A(n6715), .ZN(
        n6955) );
  AOI22_X1 U7857 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n6961), .B1(n6630), .B2(
        n5672), .ZN(n6954) );
  NAND2_X1 U7858 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(n6771), .ZN(n6631) );
  OAI21_X1 U7859 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n6771), .A(n6631), .ZN(
        n6767) );
  INV_X1 U7860 ( .A(n6918), .ZN(n6632) );
  NAND2_X1 U7861 ( .A1(n6632), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6635) );
  NAND2_X1 U7862 ( .A1(n6918), .A2(n6633), .ZN(n6634) );
  NAND2_X1 U7863 ( .A1(n6635), .A2(n6634), .ZN(n6913) );
  AOI22_X1 U7864 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6665), .B1(n6656), .B2(
        n5756), .ZN(n6641) );
  NAND2_X1 U7865 ( .A1(n6638), .A2(n6639), .ZN(n10348) );
  INV_X1 U7866 ( .A(n10348), .ZN(n6640) );
  NAND2_X1 U7867 ( .A1(n10347), .A2(n6640), .ZN(n9286) );
  NOR2_X1 U7868 ( .A1(n10353), .A2(n9286), .ZN(n10366) );
  AOI211_X1 U7869 ( .C1(n6642), .C2(n6641), .A(n6655), .B(n9590), .ZN(n6654)
         );
  NAND2_X1 U7870 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(n6771), .ZN(n6645) );
  MUX2_X1 U7871 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6643), .S(n6771), .Z(n6763)
         );
  INV_X1 U7872 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10552) );
  MUX2_X1 U7873 ( .A(n10552), .B(P1_REG1_REG_2__SCAN_IN), .S(n6961), .Z(n6957)
         );
  INV_X1 U7874 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10544) );
  MUX2_X1 U7875 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10544), .S(n6644), .Z(n6721)
         );
  NAND3_X1 U7876 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .A3(n6721), .ZN(n6720) );
  OAI21_X1 U7877 ( .B1(n6725), .B2(n10544), .A(n6720), .ZN(n6958) );
  NAND2_X1 U7878 ( .A1(n6957), .A2(n6958), .ZN(n6956) );
  OAI21_X1 U7879 ( .B1(n6961), .B2(n10552), .A(n6956), .ZN(n6762) );
  NAND2_X1 U7880 ( .A1(n6763), .A2(n6762), .ZN(n6761) );
  NAND2_X1 U7881 ( .A1(n6645), .A2(n6761), .ZN(n6910) );
  MUX2_X1 U7882 ( .A(n6646), .B(P1_REG1_REG_4__SCAN_IN), .S(n6918), .Z(n6909)
         );
  NAND2_X1 U7883 ( .A1(n6910), .A2(n6909), .ZN(n6908) );
  OAI21_X1 U7884 ( .B1(n6918), .B2(n6646), .A(n6908), .ZN(n6650) );
  MUX2_X1 U7885 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6647), .S(n6656), .Z(n6649)
         );
  INV_X1 U7886 ( .A(n10353), .ZN(n6648) );
  NAND2_X1 U7887 ( .A1(n6648), .A2(n10348), .ZN(n10362) );
  NAND2_X1 U7888 ( .A1(n6649), .A2(n6650), .ZN(n6664) );
  OAI211_X1 U7889 ( .C1(n6650), .C2(n6649), .A(n9582), .B(n6664), .ZN(n6652)
         );
  AND2_X1 U7890 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7263) );
  AOI21_X1 U7891 ( .B1(n10350), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n7263), .ZN(
        n6651) );
  OAI211_X1 U7892 ( .C1(n10360), .C2(n6665), .A(n6652), .B(n6651), .ZN(n6653)
         );
  OR2_X1 U7893 ( .A1(n6654), .A2(n6653), .ZN(P1_U3248) );
  INV_X1 U7894 ( .A(n6784), .ZN(n6657) );
  NAND2_X1 U7895 ( .A1(n6657), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6659) );
  NAND2_X1 U7896 ( .A1(n6784), .A2(n7454), .ZN(n6658) );
  NAND2_X1 U7897 ( .A1(n6659), .A2(n6658), .ZN(n6779) );
  AND2_X1 U7898 ( .A1(n6777), .A2(n6659), .ZN(n6662) );
  NAND2_X1 U7899 ( .A1(n6705), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6660) );
  OAI21_X1 U7900 ( .B1(n6705), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6660), .ZN(
        n6661) );
  AOI211_X1 U7901 ( .C1(n6662), .C2(n6661), .A(n6704), .B(n9590), .ZN(n6673)
         );
  MUX2_X1 U7902 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6663), .S(n6705), .Z(n6668)
         );
  OAI21_X1 U7903 ( .B1(n6665), .B2(n6647), .A(n6664), .ZN(n6774) );
  MUX2_X1 U7904 ( .A(n6666), .B(P1_REG1_REG_6__SCAN_IN), .S(n6784), .Z(n6775)
         );
  NAND2_X1 U7905 ( .A1(n6774), .A2(n6775), .ZN(n6773) );
  OAI21_X1 U7906 ( .B1(n6784), .B2(n6666), .A(n6773), .ZN(n6667) );
  NAND2_X1 U7907 ( .A1(n6668), .A2(n6667), .ZN(n6700) );
  OAI211_X1 U7908 ( .C1(n6668), .C2(n6667), .A(n9582), .B(n6700), .ZN(n6670)
         );
  AND2_X1 U7909 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7387) );
  AOI21_X1 U7910 ( .B1(n10350), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n7387), .ZN(
        n6669) );
  OAI211_X1 U7911 ( .C1(n10360), .C2(n6671), .A(n6670), .B(n6669), .ZN(n6672)
         );
  OR2_X1 U7912 ( .A1(n6673), .A2(n6672), .ZN(P1_U3250) );
  AOI21_X1 U7913 ( .B1(n6675), .B2(n4931), .A(n6674), .ZN(n6677) );
  MUX2_X1 U7914 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8825), .Z(n6935) );
  XOR2_X1 U7915 ( .A(n6934), .B(n6935), .Z(n6676) );
  NAND2_X1 U7916 ( .A1(n6677), .A2(n6676), .ZN(n6933) );
  OAI21_X1 U7917 ( .B1(n6677), .B2(n6676), .A(n6933), .ZN(n6678) );
  NAND2_X1 U7918 ( .A1(n6678), .A2(n10513), .ZN(n6693) );
  NAND2_X1 U7919 ( .A1(n4931), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6679) );
  NAND2_X1 U7920 ( .A1(n6680), .A2(n6679), .ZN(n6921) );
  INV_X1 U7921 ( .A(n6934), .ZN(n6681) );
  XNOR2_X1 U7922 ( .A(n6921), .B(n6681), .ZN(n6922) );
  XNOR2_X1 U7923 ( .A(n6922), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n6691) );
  NAND2_X1 U7924 ( .A1(n10498), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n6683) );
  NOR2_X1 U7925 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7084), .ZN(n6873) );
  INV_X1 U7926 ( .A(n6873), .ZN(n6682) );
  NAND2_X1 U7927 ( .A1(n6683), .A2(n6682), .ZN(n6690) );
  NAND2_X1 U7928 ( .A1(n4931), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6684) );
  INV_X1 U7929 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6686) );
  NAND2_X1 U7930 ( .A1(n6687), .A2(n6686), .ZN(n6688) );
  AOI21_X1 U7931 ( .B1(n6926), .B2(n6688), .A(n10489), .ZN(n6689) );
  AOI211_X1 U7932 ( .C1(n10483), .C2(n6691), .A(n6690), .B(n6689), .ZN(n6692)
         );
  OAI211_X1 U7933 ( .C1(n10502), .C2(n6934), .A(n6693), .B(n6692), .ZN(
        P2_U3185) );
  NOR2_X1 U7934 ( .A1(n6694), .A2(P1_U3086), .ZN(n6880) );
  XOR2_X1 U7935 ( .A(n6695), .B(n6696), .Z(n6904) );
  NAND2_X1 U7936 ( .A1(n6904), .A2(n9259), .ZN(n6698) );
  AOI22_X1 U7937 ( .A1(n8011), .A2(n5664), .B1(n9281), .B2(n10533), .ZN(n6697)
         );
  OAI211_X1 U7938 ( .C1(n6880), .C2(n10521), .A(n6698), .B(n6697), .ZN(
        P1_U3232) );
  MUX2_X1 U7939 ( .A(n6699), .B(P1_REG1_REG_9__SCAN_IN), .S(n6728), .Z(n6703)
         );
  INV_X1 U7940 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10651) );
  NAND2_X1 U7941 ( .A1(n6705), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6701) );
  NAND2_X1 U7942 ( .A1(n6701), .A2(n6700), .ZN(n6787) );
  MUX2_X1 U7943 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10651), .S(n6706), .Z(n6786)
         );
  NAND2_X1 U7944 ( .A1(n6787), .A2(n6786), .ZN(n6785) );
  OAI21_X1 U7945 ( .B1(n10651), .B2(n6794), .A(n6785), .ZN(n6702) );
  NOR2_X1 U7946 ( .A1(n6702), .A2(n6703), .ZN(n6731) );
  AOI21_X1 U7947 ( .B1(n6703), .B2(n6702), .A(n6731), .ZN(n6714) );
  MUX2_X1 U7948 ( .A(n7667), .B(P1_REG2_REG_8__SCAN_IN), .S(n6706), .Z(n6789)
         );
  AOI21_X1 U7949 ( .B1(n6706), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6788), .ZN(
        n6708) );
  AOI22_X1 U7950 ( .A1(n6728), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7680), .B2(
        n6732), .ZN(n6707) );
  AOI221_X1 U7951 ( .B1(n6708), .B2(n6727), .C1(n6707), .C2(n6727), .A(n9590), 
        .ZN(n6709) );
  INV_X1 U7952 ( .A(n6709), .ZN(n6713) );
  INV_X1 U7953 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6710) );
  NOR2_X1 U7954 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6710), .ZN(n7700) );
  NOR2_X1 U7955 ( .A1(n10360), .A2(n6732), .ZN(n6711) );
  AOI211_X1 U7956 ( .C1(n10350), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n7700), .B(
        n6711), .ZN(n6712) );
  OAI211_X1 U7957 ( .C1(n6714), .C2(n10362), .A(n6713), .B(n6712), .ZN(
        P1_U3252) );
  INV_X1 U7958 ( .A(n10350), .ZN(n10370) );
  INV_X1 U7959 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7038) );
  NOR2_X1 U7960 ( .A1(n10370), .A2(n7038), .ZN(n6719) );
  AOI211_X1 U7961 ( .C1(n6717), .C2(n6716), .A(n6715), .B(n9590), .ZN(n6718)
         );
  AOI211_X1 U7962 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(P1_U3086), .A(n6719), .B(
        n6718), .ZN(n6724) );
  NOR2_X1 U7963 ( .A1(n5576), .A2(n10534), .ZN(n6722) );
  OAI211_X1 U7964 ( .C1(n6722), .C2(n6721), .A(n9582), .B(n6720), .ZN(n6723)
         );
  OAI211_X1 U7965 ( .C1(n10360), .C2(n6725), .A(n6724), .B(n6723), .ZN(
        P1_U3244) );
  NAND2_X1 U7966 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n6886), .ZN(n6726) );
  OAI21_X1 U7967 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n6886), .A(n6726), .ZN(
        n6730) );
  AOI211_X1 U7968 ( .C1(n6730), .C2(n6729), .A(n6885), .B(n9590), .ZN(n6740)
         );
  AOI21_X1 U7969 ( .B1(n6699), .B2(n6732), .A(n6731), .ZN(n6735) );
  MUX2_X1 U7970 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6733), .S(n6886), .Z(n6734)
         );
  NAND2_X1 U7971 ( .A1(n6735), .A2(n6734), .ZN(n6890) );
  OAI211_X1 U7972 ( .C1(n6735), .C2(n6734), .A(n6890), .B(n9582), .ZN(n6738)
         );
  NAND2_X1 U7973 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n7823) );
  INV_X1 U7974 ( .A(n7823), .ZN(n6736) );
  AOI21_X1 U7975 ( .B1(n10350), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n6736), .ZN(
        n6737) );
  OAI211_X1 U7976 ( .C1(n10360), .C2(n6891), .A(n6738), .B(n6737), .ZN(n6739)
         );
  OR2_X1 U7977 ( .A1(n6740), .A2(n6739), .ZN(P1_U3253) );
  OR2_X1 U7978 ( .A1(n8187), .A2(n6742), .ZN(n6745) );
  OR2_X1 U7979 ( .A1(n6743), .A2(n5305), .ZN(n6744) );
  INV_X1 U7980 ( .A(n6747), .ZN(n6748) );
  AOI21_X1 U7981 ( .B1(n6751), .B2(n6750), .A(n5028), .ZN(n6760) );
  NAND2_X1 U7982 ( .A1(n6990), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6755) );
  NAND2_X1 U7983 ( .A1(n6865), .A2(n7084), .ZN(n6754) );
  NAND2_X1 U7984 ( .A1(n8160), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6753) );
  NAND2_X1 U7985 ( .A1(n6864), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6752) );
  NAND4_X1 U7986 ( .A1(n6755), .A2(n6754), .A3(n6753), .A4(n6752), .ZN(n8715)
         );
  NOR2_X1 U7987 ( .A1(n10565), .A2(n8679), .ZN(n6757) );
  INV_X1 U7988 ( .A(n8681), .ZN(n8697) );
  OAI22_X1 U7989 ( .A1(n10563), .A2(n8691), .B1(n8697), .B2(n10572), .ZN(n6756) );
  AOI211_X1 U7990 ( .C1(n6758), .C2(P2_REG3_REG_2__SCAN_IN), .A(n6757), .B(
        n6756), .ZN(n6759) );
  OAI21_X1 U7991 ( .B1(n6760), .B2(n8683), .A(n6759), .ZN(P2_U3177) );
  INV_X1 U7992 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6765) );
  OAI211_X1 U7993 ( .C1(n6763), .C2(n6762), .A(n9582), .B(n6761), .ZN(n6764)
         );
  NAND2_X1 U7994 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7106) );
  OAI211_X1 U7995 ( .C1(n10370), .C2(n6765), .A(n6764), .B(n7106), .ZN(n6770)
         );
  AOI211_X1 U7996 ( .C1(n6768), .C2(n6767), .A(n6766), .B(n9590), .ZN(n6769)
         );
  AOI211_X1 U7997 ( .C1(n9609), .C2(n6771), .A(n6770), .B(n6769), .ZN(n6772)
         );
  INV_X1 U7998 ( .A(n6772), .ZN(P1_U3246) );
  OAI211_X1 U7999 ( .C1(n6775), .C2(n6774), .A(n9582), .B(n6773), .ZN(n6783)
         );
  INV_X1 U8000 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6776) );
  NOR2_X1 U8001 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6776), .ZN(n7293) );
  INV_X1 U8002 ( .A(n6777), .ZN(n6778) );
  AOI211_X1 U8003 ( .C1(n6780), .C2(n6779), .A(n6778), .B(n9590), .ZN(n6781)
         );
  AOI211_X1 U8004 ( .C1(n10350), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n7293), .B(
        n6781), .ZN(n6782) );
  OAI211_X1 U8005 ( .C1(n10360), .C2(n6784), .A(n6783), .B(n6782), .ZN(
        P1_U3249) );
  OAI211_X1 U8006 ( .C1(n6787), .C2(n6786), .A(n9582), .B(n6785), .ZN(n6793)
         );
  AND2_X1 U8007 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7653) );
  AOI211_X1 U8008 ( .C1(n6790), .C2(n6789), .A(n6788), .B(n9590), .ZN(n6791)
         );
  AOI211_X1 U8009 ( .C1(n10350), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n7653), .B(
        n6791), .ZN(n6792) );
  OAI211_X1 U8010 ( .C1(n10360), .C2(n6794), .A(n6793), .B(n6792), .ZN(
        P1_U3251) );
  NAND2_X1 U8011 ( .A1(n6795), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6796) );
  XNOR2_X1 U8012 ( .A(n6796), .B(P2_IR_REG_13__SCAN_IN), .ZN(n10406) );
  INV_X1 U8013 ( .A(n10406), .ZN(n8799) );
  OAI222_X1 U8014 ( .A1(n9159), .A2(n8036), .B1(n9156), .B2(n6797), .C1(
        P2_U3151), .C2(n8799), .ZN(P2_U3282) );
  INV_X1 U8015 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6798) );
  INV_X1 U8016 ( .A(n7623), .ZN(n7619) );
  OAI222_X1 U8017 ( .A1(n10285), .A2(n6798), .B1(n8002), .B2(n8036), .C1(n7619), .C2(P1_U3086), .ZN(P1_U3342) );
  NOR2_X1 U8018 ( .A1(n10563), .A2(n10566), .ZN(n6828) );
  OR2_X1 U8019 ( .A1(n7674), .A2(n7691), .ZN(n6800) );
  NAND2_X1 U8020 ( .A1(n8505), .A2(n8833), .ZN(n6799) );
  NAND2_X1 U8021 ( .A1(n8505), .A2(n7418), .ZN(n6811) );
  NAND2_X1 U8022 ( .A1(n6801), .A2(n6811), .ZN(n6802) );
  AND2_X1 U8023 ( .A1(n10715), .A2(n6802), .ZN(n6803) );
  NOR2_X1 U8024 ( .A1(n6995), .A2(n8505), .ZN(n9008) );
  INV_X1 U8025 ( .A(n9008), .ZN(n10689) );
  INV_X1 U8026 ( .A(n10720), .ZN(n10696) );
  AOI21_X1 U8027 ( .B1(n10562), .B2(n10696), .A(n8311), .ZN(n6804) );
  AOI211_X1 U8028 ( .C1(n10671), .C2(n6805), .A(n6828), .B(n6804), .ZN(n6849)
         );
  NAND2_X1 U8029 ( .A1(n6847), .A2(n6806), .ZN(n6807) );
  NAND2_X1 U8030 ( .A1(n6810), .A2(n6809), .ZN(n6814) );
  OR2_X1 U8031 ( .A1(n6811), .A2(n7691), .ZN(n6812) );
  NAND2_X1 U8032 ( .A1(n8491), .A2(n6812), .ZN(n6820) );
  NAND2_X1 U8033 ( .A1(n6813), .A2(n6820), .ZN(n6818) );
  AOI22_X1 U8034 ( .A1(n6814), .A2(n6818), .B1(n6819), .B2(n6820), .ZN(n6815)
         );
  NAND2_X1 U8035 ( .A1(n10721), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6817) );
  OAI21_X1 U8036 ( .B1(n6849), .B2(n10721), .A(n6817), .ZN(P2_U3459) );
  AOI22_X1 U8037 ( .A1(n5332), .A2(n6820), .B1(n6819), .B2(n6818), .ZN(n6821)
         );
  NAND2_X1 U8038 ( .A1(n6822), .A2(n6821), .ZN(n6824) );
  NOR2_X1 U8039 ( .A1(n8937), .A2(n6823), .ZN(n6827) );
  INV_X1 U8040 ( .A(n6840), .ZN(n6825) );
  NOR4_X1 U8041 ( .A1(n8311), .A2(n6825), .A3(n10671), .A4(n6824), .ZN(n6826)
         );
  AOI211_X1 U8042 ( .C1(n8983), .C2(P2_REG3_REG_0__SCAN_IN), .A(n6827), .B(
        n6826), .ZN(n6830) );
  NAND2_X1 U8043 ( .A1(n6828), .A2(n10577), .ZN(n6829) );
  OAI211_X1 U8044 ( .C1(n10577), .C2(n6480), .A(n6830), .B(n6829), .ZN(
        P2_U3233) );
  NAND2_X1 U8045 ( .A1(n6832), .A2(n6831), .ZN(n6834) );
  XNOR2_X1 U8046 ( .A(n6834), .B(n6833), .ZN(n6838) );
  INV_X1 U8047 ( .A(n9278), .ZN(n7264) );
  AOI22_X1 U8048 ( .A1(n7264), .A2(n6474), .B1(n8011), .B2(n5692), .ZN(n6837)
         );
  INV_X1 U8049 ( .A(n6880), .ZN(n6835) );
  AOI22_X1 U8050 ( .A1(n6835), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n9281), .B2(
        n7496), .ZN(n6836) );
  OAI211_X1 U8051 ( .C1(n6838), .C2(n9284), .A(n6837), .B(n6836), .ZN(P1_U3222) );
  INV_X1 U8052 ( .A(n6839), .ZN(n6841) );
  AND2_X1 U8053 ( .A1(n6841), .A2(n6840), .ZN(n6845) );
  INV_X1 U8054 ( .A(n6842), .ZN(n6844) );
  OAI22_X1 U8055 ( .A1(n6846), .A2(n6845), .B1(n6844), .B2(n6843), .ZN(n6848)
         );
  INV_X1 U8056 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6851) );
  OR2_X1 U8057 ( .A1(n6849), .A2(n10724), .ZN(n6850) );
  OAI21_X1 U8058 ( .B1(n10727), .B2(n6851), .A(n6850), .ZN(P2_U3390) );
  INV_X1 U8059 ( .A(n6852), .ZN(n6853) );
  NAND2_X1 U8060 ( .A1(n6853), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8507) );
  OR2_X1 U8061 ( .A1(n8208), .A2(n5220), .ZN(n6860) );
  OR2_X1 U8062 ( .A1(n8187), .A2(n6858), .ZN(n6859) );
  OAI211_X1 U8063 ( .C1(n8249), .C2(n6934), .A(n6860), .B(n6859), .ZN(n7115)
         );
  XNOR2_X1 U8064 ( .A(n7115), .B(n6861), .ZN(n7001) );
  XNOR2_X1 U8065 ( .A(n7001), .B(n8715), .ZN(n6862) );
  NAND2_X1 U8066 ( .A1(n6863), .A2(n6862), .ZN(n7004) );
  OAI211_X1 U8067 ( .C1(n6863), .C2(n6862), .A(n7004), .B(n8685), .ZN(n6875)
         );
  NAND2_X1 U8068 ( .A1(n8291), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6871) );
  NAND2_X1 U8069 ( .A1(n7587), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6870) );
  NAND2_X1 U8070 ( .A1(n6866), .A2(n7084), .ZN(n7012) );
  NAND2_X1 U8071 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6867) );
  NAND2_X1 U8072 ( .A1(n7012), .A2(n6867), .ZN(n7121) );
  NAND2_X1 U8073 ( .A1(n8159), .A2(n7121), .ZN(n6869) );
  NAND2_X1 U8074 ( .A1(n8183), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6868) );
  AND4_X2 U8075 ( .A1(n6871), .A2(n6870), .A3(n6869), .A4(n6868), .ZN(n7276)
         );
  OAI22_X1 U8076 ( .A1(n7081), .A2(n8691), .B1(n7276), .B2(n8679), .ZN(n6872)
         );
  AOI211_X1 U8077 ( .C1(n7115), .C2(n8681), .A(n6873), .B(n6872), .ZN(n6874)
         );
  OAI211_X1 U8078 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n7381), .A(n6875), .B(
        n6874), .ZN(P2_U3158) );
  OAI21_X1 U8079 ( .B1(n6878), .B2(n6877), .A(n6876), .ZN(n6883) );
  INV_X1 U8080 ( .A(n5664), .ZN(n7345) );
  INV_X1 U8081 ( .A(n10598), .ZN(n7524) );
  OAI22_X1 U8082 ( .A1(n7345), .A2(n9278), .B1(n9276), .B2(n7524), .ZN(n6882)
         );
  OAI22_X1 U8083 ( .A1(n6880), .A2(n7351), .B1(n9242), .B2(n10548), .ZN(n6881)
         );
  AOI211_X1 U8084 ( .C1(n6883), .C2(n9259), .A(n6882), .B(n6881), .ZN(n6884)
         );
  INV_X1 U8085 ( .A(n6884), .ZN(P1_U3237) );
  AOI22_X1 U8086 ( .A1(n7157), .A2(n7789), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n7161), .ZN(n6887) );
  AOI211_X1 U8087 ( .C1(n6888), .C2(n6887), .A(n7156), .B(n9590), .ZN(n6897)
         );
  MUX2_X1 U8088 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6889), .S(n7157), .Z(n6893)
         );
  OAI21_X1 U8089 ( .B1(n6891), .B2(n6733), .A(n6890), .ZN(n6892) );
  NAND2_X1 U8090 ( .A1(n6893), .A2(n6892), .ZN(n7160) );
  OAI211_X1 U8091 ( .C1(n6893), .C2(n6892), .A(n9582), .B(n7160), .ZN(n6895)
         );
  AND2_X1 U8092 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7880) );
  AOI21_X1 U8093 ( .B1(n10350), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n7880), .ZN(
        n6894) );
  OAI211_X1 U8094 ( .C1(n10360), .C2(n7161), .A(n6895), .B(n6894), .ZN(n6896)
         );
  OR2_X1 U8095 ( .A1(n6897), .A2(n6896), .ZN(P1_U3254) );
  INV_X1 U8096 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9155) );
  NAND2_X1 U8097 ( .A1(n5498), .A2(P1_U3973), .ZN(n6898) );
  OAI21_X1 U8098 ( .B1(n9155), .B2(P1_U3973), .A(n6898), .ZN(P1_U3583) );
  INV_X1 U8099 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6899) );
  INV_X1 U8100 ( .A(n8039), .ZN(n6901) );
  INV_X1 U8101 ( .A(n7624), .ZN(n7751) );
  OAI222_X1 U8102 ( .A1(n10285), .A2(n6899), .B1(n8002), .B2(n6901), .C1(
        P1_U3086), .C2(n7751), .ZN(P1_U3341) );
  INV_X1 U8103 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6902) );
  NAND2_X1 U8104 ( .A1(n6900), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6971) );
  XNOR2_X1 U8105 ( .A(n6971), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10423) );
  OAI222_X1 U8106 ( .A1(n9156), .A2(n6902), .B1(n9159), .B2(n6901), .C1(
        P2_U3151), .C2(n8795), .ZN(P2_U3281) );
  NAND2_X1 U8107 ( .A1(n10347), .A2(n10348), .ZN(n6907) );
  NAND2_X1 U8108 ( .A1(n10347), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6903) );
  XOR2_X1 U8109 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6903), .Z(n6906) );
  NOR2_X1 U8110 ( .A1(n6904), .A2(n6907), .ZN(n6905) );
  AOI211_X1 U8111 ( .C1(n6907), .C2(n6906), .A(n9561), .B(n6905), .ZN(n6965)
         );
  AND2_X1 U8112 ( .A1(n10350), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n6920) );
  OAI211_X1 U8113 ( .C1(n6910), .C2(n6909), .A(n9582), .B(n6908), .ZN(n6917)
         );
  AND2_X1 U8114 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7092) );
  INV_X1 U8115 ( .A(n6911), .ZN(n6912) );
  AOI211_X1 U8116 ( .C1(n6914), .C2(n6913), .A(n6912), .B(n9590), .ZN(n6915)
         );
  NOR2_X1 U8117 ( .A1(n7092), .A2(n6915), .ZN(n6916) );
  OAI211_X1 U8118 ( .C1(n10360), .C2(n6918), .A(n6917), .B(n6916), .ZN(n6919)
         );
  OR3_X1 U8119 ( .A1(n6965), .A2(n6920), .A3(n6919), .ZN(P1_U3247) );
  INV_X1 U8120 ( .A(n7064), .ZN(n6940) );
  INV_X1 U8121 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10594) );
  MUX2_X1 U8122 ( .A(n10594), .B(P2_REG1_REG_4__SCAN_IN), .S(n7064), .Z(n6924)
         );
  AOI22_X1 U8123 ( .A1(n6922), .A2(P2_REG1_REG_3__SCAN_IN), .B1(n6934), .B2(
        n6921), .ZN(n6923) );
  NOR2_X1 U8124 ( .A1(n6923), .A2(n6924), .ZN(n7054) );
  AOI21_X1 U8125 ( .B1(n6924), .B2(n6923), .A(n7054), .ZN(n6932) );
  NOR2_X1 U8126 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6866), .ZN(n7019) );
  AOI21_X1 U8127 ( .B1(n10498), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n7019), .ZN(
        n6931) );
  INV_X1 U8128 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6925) );
  MUX2_X1 U8129 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6925), .S(n7064), .Z(n6928)
         );
  NAND2_X1 U8130 ( .A1(n6927), .A2(n6928), .ZN(n7056) );
  OAI21_X1 U8131 ( .B1(n6928), .B2(n6927), .A(n7056), .ZN(n6929) );
  NAND2_X1 U8132 ( .A1(n10509), .A2(n6929), .ZN(n6930) );
  OAI211_X1 U8133 ( .C1(n6932), .C2(n10496), .A(n6931), .B(n6930), .ZN(n6939)
         );
  MUX2_X1 U8134 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8825), .Z(n7065) );
  XNOR2_X1 U8135 ( .A(n7065), .B(n7064), .ZN(n6937) );
  OAI21_X1 U8136 ( .B1(n6935), .B2(n6934), .A(n6933), .ZN(n6936) );
  NOR2_X1 U8137 ( .A1(n6936), .A2(n6937), .ZN(n7063) );
  AOI211_X1 U8138 ( .C1(n6937), .C2(n6936), .A(n8830), .B(n7063), .ZN(n6938)
         );
  AOI211_X1 U8139 ( .C1(n10476), .C2(n6940), .A(n6939), .B(n6938), .ZN(n6941)
         );
  INV_X1 U8140 ( .A(n6941), .ZN(P2_U3186) );
  INV_X1 U8141 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6952) );
  INV_X1 U8142 ( .A(n8345), .ZN(n6945) );
  INV_X1 U8143 ( .A(n6943), .ZN(n6942) );
  INV_X1 U8144 ( .A(n7074), .ZN(n6944) );
  AOI21_X1 U8145 ( .B1(n6945), .B2(n8338), .A(n6944), .ZN(n7000) );
  OAI21_X1 U8146 ( .B1(n6947), .B2(n8338), .A(n10558), .ZN(n6949) );
  AOI222_X1 U8147 ( .A1(n8989), .A2(n6949), .B1(n8716), .B2(n8995), .C1(n8717), 
        .C2(n8994), .ZN(n6996) );
  OAI21_X1 U8148 ( .B1(n10696), .B2(n7000), .A(n6996), .ZN(n6968) );
  NAND2_X1 U8149 ( .A1(n6968), .A2(n10727), .ZN(n6951) );
  NAND2_X1 U8150 ( .A1(n9141), .A2(n6997), .ZN(n6950) );
  OAI211_X1 U8151 ( .C1(n10727), .C2(n6952), .A(n6951), .B(n6950), .ZN(
        P2_U3393) );
  AOI211_X1 U8152 ( .C1(n6955), .C2(n6954), .A(n6953), .B(n9590), .ZN(n6964)
         );
  AOI22_X1 U8153 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(n10350), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6960) );
  OAI211_X1 U8154 ( .C1(n6958), .C2(n6957), .A(n9582), .B(n6956), .ZN(n6959)
         );
  NAND2_X1 U8155 ( .A1(n6960), .A2(n6959), .ZN(n6963) );
  NOR2_X1 U8156 ( .A1(n10360), .A2(n6961), .ZN(n6962) );
  OR4_X1 U8157 ( .A1(n6965), .A2(n6964), .A3(n6963), .A4(n6962), .ZN(P1_U3245)
         );
  INV_X1 U8158 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6966) );
  OAI22_X1 U8159 ( .A1(n9050), .A2(n7078), .B1(n10723), .B2(n6966), .ZN(n6967)
         );
  AOI21_X1 U8160 ( .B1(n6968), .B2(n10723), .A(n6967), .ZN(n6969) );
  INV_X1 U8161 ( .A(n6969), .ZN(P2_U3460) );
  NAND2_X1 U8162 ( .A1(n6971), .A2(n6970), .ZN(n6972) );
  NAND2_X1 U8163 ( .A1(n6972), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7099) );
  XNOR2_X1 U8164 ( .A(n7099), .B(P2_IR_REG_15__SCAN_IN), .ZN(n10440) );
  INV_X1 U8165 ( .A(n10440), .ZN(n8791) );
  INV_X1 U8166 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6973) );
  OAI222_X1 U8167 ( .A1(n9159), .A2(n8106), .B1(n8791), .B2(P2_U3151), .C1(
        n6973), .C2(n9156), .ZN(P2_U3280) );
  INV_X1 U8168 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6974) );
  INV_X1 U8169 ( .A(n7853), .ZN(n7860) );
  OAI222_X1 U8170 ( .A1(n10285), .A2(n6974), .B1(n8002), .B2(n8106), .C1(n7860), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U8171 ( .A(n7012), .ZN(n6976) );
  NAND2_X1 U8172 ( .A1(n6976), .A2(n6975), .ZN(n7134) );
  OR2_X2 U8173 ( .A1(n8122), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8135) );
  INV_X1 U8174 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6988) );
  INV_X1 U8175 ( .A(n7045), .ZN(n8181) );
  NAND2_X1 U8176 ( .A1(n8171), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6989) );
  NAND2_X1 U8177 ( .A1(n8181), .A2(n6989), .ZN(n8901) );
  NAND2_X1 U8178 ( .A1(n8901), .A2(n8159), .ZN(n6993) );
  AOI22_X1 U8179 ( .A1(n8291), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n7587), .B2(
        P2_REG1_REG_23__SCAN_IN), .ZN(n6992) );
  NAND2_X1 U8180 ( .A1(n8160), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6991) );
  NAND2_X1 U8181 ( .A1(n8624), .A2(P2_U3893), .ZN(n6994) );
  OAI21_X1 U8182 ( .B1(P2_U3893), .B2(n7816), .A(n6994), .ZN(P2_U3514) );
  OR2_X1 U8183 ( .A1(n7674), .A2(n6995), .ZN(n7464) );
  NAND2_X1 U8184 ( .A1(n8256), .A2(n7464), .ZN(n10576) );
  MUX2_X1 U8185 ( .A(n6616), .B(n6996), .S(n10577), .Z(n6999) );
  AOI22_X1 U8186 ( .A1(n9001), .A2(n6997), .B1(n8983), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n6998) );
  OAI211_X1 U8187 ( .C1(n9004), .C2(n7000), .A(n6999), .B(n6998), .ZN(P2_U3232) );
  NAND2_X1 U8188 ( .A1(n7004), .A2(n7003), .ZN(n7011) );
  OR2_X1 U8189 ( .A1(n8208), .A2(n7005), .ZN(n7008) );
  OR2_X1 U8190 ( .A1(n8187), .A2(n7006), .ZN(n7007) );
  OAI211_X1 U8191 ( .C1(n8249), .C2(n7064), .A(n7008), .B(n7007), .ZN(n7230)
         );
  XNOR2_X1 U8192 ( .A(n7230), .B(n8552), .ZN(n7009) );
  NAND2_X1 U8193 ( .A1(n7276), .A2(n7009), .ZN(n7125) );
  OAI21_X1 U8194 ( .B1(n7276), .B2(n7009), .A(n7125), .ZN(n7010) );
  AOI21_X1 U8195 ( .B1(n7011), .B2(n7010), .A(n7131), .ZN(n7022) );
  NAND2_X1 U8196 ( .A1(n8291), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7017) );
  NAND2_X1 U8197 ( .A1(n7587), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7016) );
  NAND2_X1 U8198 ( .A1(n7012), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7013) );
  NAND2_X1 U8199 ( .A1(n7134), .A2(n7013), .ZN(n7124) );
  NAND2_X1 U8200 ( .A1(n8159), .A2(n7124), .ZN(n7015) );
  NAND2_X1 U8201 ( .A1(n8183), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7014) );
  NAND4_X1 U8202 ( .A1(n7017), .A2(n7016), .A3(n7015), .A4(n7014), .ZN(n8713)
         );
  OAI22_X1 U8203 ( .A1(n7315), .A2(n8679), .B1(n10565), .B2(n8691), .ZN(n7018)
         );
  AOI211_X1 U8204 ( .C1(n7230), .C2(n8681), .A(n7019), .B(n7018), .ZN(n7021)
         );
  NAND2_X1 U8205 ( .A1(n8694), .A2(n7121), .ZN(n7020) );
  OAI211_X1 U8206 ( .C1(n7022), .C2(n8683), .A(n7021), .B(n7020), .ZN(P2_U3170) );
  NOR2_X1 U8207 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n7023) );
  AOI21_X1 U8208 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n7023), .ZN(n10345) );
  NOR2_X1 U8209 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7024) );
  AOI21_X1 U8210 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7024), .ZN(n10342) );
  NOR2_X1 U8211 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7025) );
  AOI21_X1 U8212 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7025), .ZN(n10339) );
  NOR2_X1 U8213 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7026) );
  AOI21_X1 U8214 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7026), .ZN(n10336) );
  NOR2_X1 U8215 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7027) );
  AOI21_X1 U8216 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7027), .ZN(n10333) );
  NOR2_X1 U8217 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7028) );
  AOI21_X1 U8218 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7028), .ZN(n10330) );
  NOR2_X1 U8219 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7029) );
  AOI21_X1 U8220 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7029), .ZN(n10327) );
  NOR2_X1 U8221 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7030) );
  AOI21_X1 U8222 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7030), .ZN(n10324) );
  NOR2_X1 U8223 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7031) );
  AOI21_X1 U8224 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7031), .ZN(n10321) );
  NOR2_X1 U8225 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7032) );
  AOI21_X1 U8226 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7032), .ZN(n10318) );
  NOR2_X1 U8227 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7033) );
  AOI21_X1 U8228 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7033), .ZN(n10315) );
  NOR2_X1 U8229 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7034) );
  AOI21_X1 U8230 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7034), .ZN(n10312) );
  NOR2_X1 U8231 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7035) );
  AOI21_X1 U8232 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7035), .ZN(n10309) );
  NOR2_X1 U8233 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7036) );
  AOI21_X1 U8234 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7036), .ZN(n10306) );
  NAND2_X1 U8235 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n7037) );
  NAND2_X1 U8236 ( .A1(n7038), .A2(n7037), .ZN(n10292) );
  INV_X1 U8237 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10294) );
  NAND3_X1 U8238 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10293) );
  NAND2_X1 U8239 ( .A1(n10294), .A2(n10293), .ZN(n10290) );
  NAND2_X1 U8240 ( .A1(n10292), .A2(n10290), .ZN(n10297) );
  NAND2_X1 U8241 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7039) );
  OAI21_X1 U8242 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7039), .ZN(n10296) );
  NOR2_X1 U8243 ( .A1(n10297), .A2(n10296), .ZN(n10295) );
  AOI21_X1 U8244 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10295), .ZN(n10300) );
  NAND2_X1 U8245 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7040) );
  OAI21_X1 U8246 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n7040), .ZN(n10299) );
  NOR2_X1 U8247 ( .A1(n10300), .A2(n10299), .ZN(n10298) );
  AOI21_X1 U8248 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10298), .ZN(n10303) );
  NOR2_X1 U8249 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7041) );
  AOI21_X1 U8250 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7041), .ZN(n10302) );
  NAND2_X1 U8251 ( .A1(n10303), .A2(n10302), .ZN(n10301) );
  OAI21_X1 U8252 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10301), .ZN(n10305) );
  NAND2_X1 U8253 ( .A1(n10306), .A2(n10305), .ZN(n10304) );
  OAI21_X1 U8254 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10304), .ZN(n10308) );
  NAND2_X1 U8255 ( .A1(n10309), .A2(n10308), .ZN(n10307) );
  OAI21_X1 U8256 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10307), .ZN(n10311) );
  NAND2_X1 U8257 ( .A1(n10312), .A2(n10311), .ZN(n10310) );
  OAI21_X1 U8258 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10310), .ZN(n10314) );
  NAND2_X1 U8259 ( .A1(n10315), .A2(n10314), .ZN(n10313) );
  OAI21_X1 U8260 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10313), .ZN(n10317) );
  NAND2_X1 U8261 ( .A1(n10318), .A2(n10317), .ZN(n10316) );
  OAI21_X1 U8262 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10316), .ZN(n10320) );
  NAND2_X1 U8263 ( .A1(n10321), .A2(n10320), .ZN(n10319) );
  OAI21_X1 U8264 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10319), .ZN(n10323) );
  NAND2_X1 U8265 ( .A1(n10324), .A2(n10323), .ZN(n10322) );
  OAI21_X1 U8266 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10322), .ZN(n10326) );
  NAND2_X1 U8267 ( .A1(n10327), .A2(n10326), .ZN(n10325) );
  OAI21_X1 U8268 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10325), .ZN(n10329) );
  NAND2_X1 U8269 ( .A1(n10330), .A2(n10329), .ZN(n10328) );
  OAI21_X1 U8270 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10328), .ZN(n10332) );
  NAND2_X1 U8271 ( .A1(n10333), .A2(n10332), .ZN(n10331) );
  OAI21_X1 U8272 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10331), .ZN(n10335) );
  NAND2_X1 U8273 ( .A1(n10336), .A2(n10335), .ZN(n10334) );
  OAI21_X1 U8274 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10334), .ZN(n10338) );
  NAND2_X1 U8275 ( .A1(n10339), .A2(n10338), .ZN(n10337) );
  OAI21_X1 U8276 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10337), .ZN(n10341) );
  NAND2_X1 U8277 ( .A1(n10342), .A2(n10341), .ZN(n10340) );
  OAI21_X1 U8278 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10340), .ZN(n10344) );
  NAND2_X1 U8279 ( .A1(n10345), .A2(n10344), .ZN(n10343) );
  OAI21_X1 U8280 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10343), .ZN(n7044) );
  XNOR2_X1 U8281 ( .A(n7042), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7043) );
  XNOR2_X1 U8282 ( .A(n7044), .B(n7043), .ZN(ADD_1068_U4) );
  INV_X1 U8283 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10158) );
  INV_X1 U8284 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n7046) );
  XNOR2_X1 U8285 ( .A(n8194), .B(P2_REG3_REG_26__SCAN_IN), .ZN(n8871) );
  NAND2_X1 U8286 ( .A1(n8871), .A2(n8159), .ZN(n7052) );
  INV_X1 U8287 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9085) );
  NAND2_X1 U8288 ( .A1(n8291), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n7049) );
  NAND2_X1 U8289 ( .A1(n7587), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n7048) );
  OAI211_X1 U8290 ( .C1(n9085), .C2(n8215), .A(n7049), .B(n7048), .ZN(n7050)
         );
  INV_X1 U8291 ( .A(n7050), .ZN(n7051) );
  NAND2_X1 U8292 ( .A1(n8859), .A2(P2_U3893), .ZN(n7053) );
  OAI21_X1 U8293 ( .B1(P2_U3893), .B2(n6234), .A(n7053), .ZN(P2_U3517) );
  AOI21_X1 U8294 ( .B1(n7064), .B2(P2_REG1_REG_4__SCAN_IN), .A(n7054), .ZN(
        n7171) );
  XNOR2_X1 U8295 ( .A(n7171), .B(n7177), .ZN(n7173) );
  XNOR2_X1 U8296 ( .A(n7173), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n7070) );
  NOR2_X1 U8297 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6975), .ZN(n7141) );
  NAND2_X1 U8298 ( .A1(n7064), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7055) );
  OAI21_X1 U8299 ( .B1(n7057), .B2(n7177), .A(n7184), .ZN(n7059) );
  INV_X1 U8300 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7058) );
  NAND2_X1 U8301 ( .A1(n7059), .A2(n7058), .ZN(n7060) );
  AOI21_X1 U8302 ( .B1(n7186), .B2(n7060), .A(n10489), .ZN(n7061) );
  AOI211_X1 U8303 ( .C1(n10498), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n7141), .B(
        n7061), .ZN(n7062) );
  OAI21_X1 U8304 ( .B1(n7177), .B2(n10502), .A(n7062), .ZN(n7069) );
  MUX2_X1 U8305 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8825), .Z(n7178) );
  XNOR2_X1 U8306 ( .A(n7178), .B(n7177), .ZN(n7067) );
  AOI21_X1 U8307 ( .B1(n7065), .B2(n7064), .A(n7063), .ZN(n7066) );
  NOR2_X1 U8308 ( .A1(n7066), .A2(n7067), .ZN(n7176) );
  AOI211_X1 U8309 ( .C1(n7067), .C2(n7066), .A(n8830), .B(n7176), .ZN(n7068)
         );
  AOI211_X1 U8310 ( .C1(n10483), .C2(n7070), .A(n7069), .B(n7068), .ZN(n7071)
         );
  INV_X1 U8311 ( .A(n7071), .ZN(P2_U3187) );
  NAND2_X1 U8312 ( .A1(n10565), .A2(n7115), .ZN(n8350) );
  INV_X1 U8313 ( .A(n7115), .ZN(n10582) );
  NAND2_X1 U8314 ( .A1(n8715), .A2(n10582), .ZN(n8357) );
  INV_X1 U8315 ( .A(n8349), .ZN(n7073) );
  NOR2_X1 U8316 ( .A1(n8314), .A2(n7073), .ZN(n7077) );
  NAND2_X1 U8317 ( .A1(n8349), .A2(n8351), .ZN(n7079) );
  INV_X1 U8318 ( .A(n7079), .ZN(n10557) );
  NAND2_X1 U8319 ( .A1(n7074), .A2(n8346), .ZN(n8337) );
  NAND2_X1 U8320 ( .A1(n10557), .A2(n8337), .ZN(n10555) );
  NAND2_X1 U8321 ( .A1(n10555), .A2(n8349), .ZN(n7075) );
  NAND2_X1 U8322 ( .A1(n7075), .A2(n8314), .ZN(n7111) );
  INV_X1 U8323 ( .A(n7111), .ZN(n7076) );
  AOI21_X1 U8324 ( .B1(n7077), .B2(n10555), .A(n7076), .ZN(n10583) );
  NAND2_X1 U8325 ( .A1(n10563), .A2(n7078), .ZN(n10556) );
  NAND2_X1 U8326 ( .A1(n10558), .A2(n10556), .ZN(n7080) );
  NAND2_X1 U8327 ( .A1(n7080), .A2(n7079), .ZN(n10560) );
  NAND2_X1 U8328 ( .A1(n7081), .A2(n10572), .ZN(n7082) );
  NAND2_X1 U8329 ( .A1(n10560), .A2(n7082), .ZN(n7117) );
  XOR2_X1 U8330 ( .A(n8314), .B(n7117), .Z(n7083) );
  INV_X1 U8331 ( .A(n7276), .ZN(n8714) );
  AOI222_X1 U8332 ( .A1(n8989), .A2(n7083), .B1(n8714), .B2(n8995), .C1(n8716), 
        .C2(n8994), .ZN(n10581) );
  MUX2_X1 U8333 ( .A(n6686), .B(n10581), .S(n10577), .Z(n7086) );
  AOI22_X1 U8334 ( .A1(n9001), .A2(n7115), .B1(n8983), .B2(n7084), .ZN(n7085)
         );
  OAI211_X1 U8335 ( .C1(n10583), .C2(n9004), .A(n7086), .B(n7085), .ZN(
        P2_U3230) );
  NAND2_X1 U8336 ( .A1(n7087), .A2(n9259), .ZN(n7096) );
  AOI21_X1 U8337 ( .B1(n7088), .B2(n7090), .A(n7089), .ZN(n7095) );
  AOI22_X1 U8338 ( .A1(n7264), .A2(n10598), .B1(n9281), .B2(n10597), .ZN(n7094) );
  NOR2_X1 U8339 ( .A1(n9275), .A2(n7518), .ZN(n7091) );
  AOI211_X1 U8340 ( .C1(n8011), .C2(n7514), .A(n7092), .B(n7091), .ZN(n7093)
         );
  OAI211_X1 U8341 ( .C1(n7096), .C2(n7095), .A(n7094), .B(n7093), .ZN(P1_U3230) );
  INV_X1 U8342 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7097) );
  INV_X1 U8343 ( .A(n8102), .ZN(n7101) );
  INV_X1 U8344 ( .A(n9564), .ZN(n7857) );
  OAI222_X1 U8345 ( .A1(n10285), .A2(n7097), .B1(n8002), .B2(n7101), .C1(
        P1_U3086), .C2(n7857), .ZN(P1_U3339) );
  INV_X1 U8346 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7102) );
  NAND2_X1 U8347 ( .A1(n7099), .A2(n7098), .ZN(n7100) );
  NAND2_X1 U8348 ( .A1(n7100), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7283) );
  XNOR2_X1 U8349 ( .A(n7283), .B(P2_IR_REG_16__SCAN_IN), .ZN(n10457) );
  OAI222_X1 U8350 ( .A1(n9156), .A2(n7102), .B1(n9159), .B2(n7101), .C1(
        P2_U3151), .C2(n8787), .ZN(P2_U3279) );
  OAI21_X1 U8351 ( .B1(n7104), .B2(n7103), .A(n7088), .ZN(n7109) );
  OAI22_X1 U8352 ( .A1(n9278), .A2(n7203), .B1(n9242), .B2(n7507), .ZN(n7108)
         );
  INV_X1 U8353 ( .A(n9560), .ZN(n10609) );
  OR2_X1 U8354 ( .A1(n9275), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7105) );
  OAI211_X1 U8355 ( .C1(n9276), .C2(n10609), .A(n7106), .B(n7105), .ZN(n7107)
         );
  AOI211_X1 U8356 ( .C1(n7109), .C2(n9259), .A(n7108), .B(n7107), .ZN(n7110)
         );
  INV_X1 U8357 ( .A(n7110), .ZN(P1_U3218) );
  OR2_X1 U8358 ( .A1(n7276), .A2(n7230), .ZN(n8362) );
  NAND2_X1 U8359 ( .A1(n7276), .A2(n7230), .ZN(n8358) );
  INV_X1 U8360 ( .A(n8350), .ZN(n8363) );
  NOR2_X1 U8361 ( .A1(n8356), .A2(n8363), .ZN(n7114) );
  NAND2_X1 U8362 ( .A1(n7111), .A2(n8350), .ZN(n7112) );
  NAND2_X1 U8363 ( .A1(n7112), .A2(n8356), .ZN(n7249) );
  INV_X1 U8364 ( .A(n7249), .ZN(n7113) );
  AOI21_X1 U8365 ( .B1(n7114), .B2(n7111), .A(n7113), .ZN(n10591) );
  NAND2_X1 U8366 ( .A1(n8715), .A2(n7115), .ZN(n7116) );
  NAND2_X1 U8367 ( .A1(n7117), .A2(n7116), .ZN(n7119) );
  NAND2_X1 U8368 ( .A1(n10565), .A2(n10582), .ZN(n7118) );
  NAND2_X1 U8369 ( .A1(n7119), .A2(n7118), .ZN(n7229) );
  XOR2_X1 U8370 ( .A(n7229), .B(n8356), .Z(n7120) );
  AOI222_X1 U8371 ( .A1(n8989), .A2(n7120), .B1(n8715), .B2(n8994), .C1(n8713), 
        .C2(n8995), .ZN(n10589) );
  MUX2_X1 U8372 ( .A(n6925), .B(n10589), .S(n10577), .Z(n7123) );
  AOI22_X1 U8373 ( .A1(n9001), .A2(n7230), .B1(n8983), .B2(n7121), .ZN(n7122)
         );
  OAI211_X1 U8374 ( .C1(n10591), .C2(n9004), .A(n7123), .B(n7122), .ZN(
        P2_U3229) );
  INV_X1 U8375 ( .A(n7124), .ZN(n7482) );
  INV_X1 U8376 ( .A(n7125), .ZN(n7130) );
  OR2_X1 U8377 ( .A1(n8208), .A2(n6473), .ZN(n7127) );
  XNOR2_X1 U8378 ( .A(n7277), .B(n8552), .ZN(n7309) );
  XNOR2_X1 U8379 ( .A(n7309), .B(n8713), .ZN(n7129) );
  INV_X1 U8380 ( .A(n7310), .ZN(n7133) );
  NOR3_X1 U8381 ( .A1(n7131), .A2(n7130), .A3(n7129), .ZN(n7132) );
  OAI21_X1 U8382 ( .B1(n7133), .B2(n7132), .A(n8685), .ZN(n7143) );
  NAND2_X1 U8383 ( .A1(n8291), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7139) );
  NAND2_X1 U8384 ( .A1(n7587), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7138) );
  NAND2_X1 U8385 ( .A1(n7134), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7135) );
  NAND2_X1 U8386 ( .A1(n7241), .A2(n7135), .ZN(n7308) );
  NAND2_X1 U8387 ( .A1(n8159), .A2(n7308), .ZN(n7137) );
  NAND2_X1 U8388 ( .A1(n8183), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7136) );
  NAND4_X1 U8389 ( .A1(n7139), .A2(n7138), .A3(n7137), .A4(n7136), .ZN(n8712)
         );
  INV_X1 U8390 ( .A(n8712), .ZN(n7471) );
  OAI22_X1 U8391 ( .A1(n7471), .A2(n8679), .B1(n7276), .B2(n8691), .ZN(n7140)
         );
  AOI211_X1 U8392 ( .C1(n7277), .C2(n8681), .A(n7141), .B(n7140), .ZN(n7142)
         );
  OAI211_X1 U8393 ( .C1(n7482), .C2(n7381), .A(n7143), .B(n7142), .ZN(P2_U3167) );
  INV_X1 U8394 ( .A(n8194), .ZN(n7144) );
  INV_X1 U8395 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10265) );
  INV_X1 U8396 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7145) );
  INV_X1 U8397 ( .A(n7146), .ZN(n7147) );
  NAND2_X1 U8398 ( .A1(n7147), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n7148) );
  NAND2_X1 U8399 ( .A1(n8211), .A2(n7148), .ZN(n8862) );
  NAND2_X1 U8400 ( .A1(n8862), .A2(n8159), .ZN(n7153) );
  INV_X1 U8401 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9079) );
  NAND2_X1 U8402 ( .A1(n8291), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n7150) );
  NAND2_X1 U8403 ( .A1(n7587), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n7149) );
  OAI211_X1 U8404 ( .C1(n9079), .C2(n8215), .A(n7150), .B(n7149), .ZN(n7151)
         );
  INV_X1 U8405 ( .A(n7151), .ZN(n7152) );
  NAND2_X1 U8406 ( .A1(n8554), .A2(P2_U3893), .ZN(n7154) );
  OAI21_X1 U8407 ( .B1(n6258), .B2(P2_U3893), .A(n7154), .ZN(P2_U3518) );
  AOI22_X1 U8408 ( .A1(n7623), .A2(n7920), .B1(P1_REG2_REG_13__SCAN_IN), .B2(
        n7619), .ZN(n7159) );
  NOR2_X1 U8409 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7162), .ZN(n7155) );
  AOI21_X1 U8410 ( .B1(n7162), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7155), .ZN(
        n10356) );
  AOI21_X1 U8411 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7157), .A(n7156), .ZN(
        n10355) );
  NAND2_X1 U8412 ( .A1(n10356), .A2(n10355), .ZN(n10354) );
  OAI21_X1 U8413 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7162), .A(n10354), .ZN(
        n7158) );
  NOR2_X1 U8414 ( .A1(n7159), .A2(n7158), .ZN(n7622) );
  AOI211_X1 U8415 ( .C1(n7159), .C2(n7158), .A(n7622), .B(n9590), .ZN(n7170)
         );
  AOI22_X1 U8416 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n10361), .B1(n7162), .B2(
        n5932), .ZN(n10359) );
  OAI21_X1 U8417 ( .B1(n6889), .B2(n7161), .A(n7160), .ZN(n10358) );
  NOR2_X1 U8418 ( .A1(n10359), .A2(n10358), .ZN(n10357) );
  NOR2_X1 U8419 ( .A1(n7162), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7163) );
  NOR2_X1 U8420 ( .A1(n10357), .A2(n7163), .ZN(n7166) );
  MUX2_X1 U8421 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7164), .S(n7623), .Z(n7165)
         );
  NAND2_X1 U8422 ( .A1(n7166), .A2(n7165), .ZN(n7618) );
  OAI211_X1 U8423 ( .C1(n7166), .C2(n7165), .A(n7618), .B(n9582), .ZN(n7168)
         );
  AND2_X1 U8424 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n8010) );
  AOI21_X1 U8425 ( .B1(n10350), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n8010), .ZN(
        n7167) );
  OAI211_X1 U8426 ( .C1(n10360), .C2(n7619), .A(n7168), .B(n7167), .ZN(n7169)
         );
  OR2_X1 U8427 ( .A1(n7170), .A2(n7169), .ZN(P1_U3256) );
  INV_X1 U8428 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10618) );
  MUX2_X1 U8429 ( .A(n10618), .B(P2_REG1_REG_6__SCAN_IN), .S(n7326), .Z(n7175)
         );
  INV_X1 U8430 ( .A(n7171), .ZN(n7172) );
  AOI21_X1 U8431 ( .B1(n7175), .B2(n7174), .A(n7325), .ZN(n7196) );
  AOI21_X1 U8432 ( .B1(n7178), .B2(n7177), .A(n7176), .ZN(n7180) );
  MUX2_X1 U8433 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8825), .Z(n7324) );
  XOR2_X1 U8434 ( .A(n7326), .B(n7324), .Z(n7179) );
  NAND2_X1 U8435 ( .A1(n7180), .A2(n7179), .ZN(n7323) );
  OAI21_X1 U8436 ( .B1(n7180), .B2(n7179), .A(n7323), .ZN(n7181) );
  NAND2_X1 U8437 ( .A1(n7181), .A2(n10513), .ZN(n7195) );
  INV_X1 U8438 ( .A(n7326), .ZN(n7193) );
  INV_X1 U8439 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7252) );
  MUX2_X1 U8440 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7252), .S(n7326), .Z(n7183)
         );
  INV_X1 U8441 ( .A(n7183), .ZN(n7185) );
  NAND3_X1 U8442 ( .A1(n7186), .A2(n7185), .A3(n7184), .ZN(n7187) );
  AND2_X1 U8443 ( .A1(n7327), .A2(n7187), .ZN(n7191) );
  NAND2_X1 U8444 ( .A1(n10498), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7190) );
  INV_X1 U8445 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7188) );
  NOR2_X1 U8446 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7188), .ZN(n7317) );
  INV_X1 U8447 ( .A(n7317), .ZN(n7189) );
  OAI211_X1 U8448 ( .C1(n10489), .C2(n7191), .A(n7190), .B(n7189), .ZN(n7192)
         );
  AOI21_X1 U8449 ( .B1(n7193), .B2(n10476), .A(n7192), .ZN(n7194) );
  OAI211_X1 U8450 ( .C1(n7196), .C2(n10496), .A(n7195), .B(n7194), .ZN(
        P2_U3188) );
  INV_X1 U8451 ( .A(n10532), .ZN(n7200) );
  NAND2_X1 U8452 ( .A1(n7198), .A2(n7197), .ZN(n7199) );
  NAND2_X1 U8453 ( .A1(n7200), .A2(n7199), .ZN(n7201) );
  INV_X1 U8454 ( .A(n7496), .ZN(n10539) );
  NAND2_X1 U8455 ( .A1(n6474), .A2(n10533), .ZN(n7493) );
  NAND2_X1 U8456 ( .A1(n7345), .A2(n10539), .ZN(n7202) );
  NAND2_X1 U8457 ( .A1(n7492), .A2(n7202), .ZN(n7338) );
  NAND2_X1 U8458 ( .A1(n7203), .A2(n6879), .ZN(n7209) );
  NAND2_X1 U8459 ( .A1(n5692), .A2(n10548), .ZN(n7426) );
  NAND2_X1 U8460 ( .A1(n7209), .A2(n7426), .ZN(n9356) );
  NAND2_X1 U8461 ( .A1(n7203), .A2(n10548), .ZN(n7204) );
  NAND2_X1 U8462 ( .A1(n7337), .A2(n7204), .ZN(n7205) );
  NAND2_X1 U8463 ( .A1(n7524), .A2(n7214), .ZN(n9309) );
  NAND2_X1 U8464 ( .A1(n10598), .A2(n7507), .ZN(n9394) );
  NAND2_X1 U8465 ( .A1(n9309), .A2(n9394), .ZN(n7206) );
  NAND2_X1 U8466 ( .A1(n7205), .A2(n7206), .ZN(n7422) );
  OAI21_X1 U8467 ( .B1(n7205), .B2(n7206), .A(n7422), .ZN(n7509) );
  INV_X1 U8468 ( .A(n7509), .ZN(n7216) );
  INV_X1 U8469 ( .A(n7206), .ZN(n9358) );
  NAND2_X1 U8470 ( .A1(n9366), .A2(n9363), .ZN(n7208) );
  NAND2_X1 U8471 ( .A1(n7345), .A2(n7496), .ZN(n7207) );
  INV_X1 U8472 ( .A(n7209), .ZN(n7210) );
  AND2_X1 U8473 ( .A1(n9304), .A2(n7426), .ZN(n9397) );
  NAND2_X1 U8474 ( .A1(n9397), .A2(n9358), .ZN(n7512) );
  OAI21_X1 U8475 ( .B1(n9358), .B2(n9397), .A(n7512), .ZN(n7213) );
  NAND2_X1 U8476 ( .A1(n6319), .A2(n9610), .ZN(n7212) );
  NAND2_X1 U8477 ( .A1(n5609), .A2(n9544), .ZN(n7211) );
  AOI22_X1 U8478 ( .A1(n7213), .A2(n9852), .B1(n10519), .B2(n9560), .ZN(n7511)
         );
  OR2_X1 U8479 ( .A1(n7496), .A2(n10533), .ZN(n7498) );
  OR2_X1 U8480 ( .A1(n7498), .A2(n6879), .ZN(n7352) );
  NOR2_X2 U8481 ( .A1(n7352), .A2(n7214), .ZN(n7523) );
  AOI211_X1 U8482 ( .C1(n7214), .C2(n7352), .A(n9826), .B(n7523), .ZN(n7503)
         );
  AOI21_X1 U8483 ( .B1(n10704), .B2(n5692), .A(n7503), .ZN(n7215) );
  OAI211_X1 U8484 ( .C1(n10528), .C2(n7216), .A(n7511), .B(n7215), .ZN(n7227)
         );
  INV_X1 U8485 ( .A(n7340), .ZN(n7217) );
  AND2_X1 U8486 ( .A1(n7342), .A2(n7217), .ZN(n7225) );
  NAND2_X1 U8487 ( .A1(n7219), .A2(n7218), .ZN(n7220) );
  INV_X1 U8488 ( .A(n7224), .ZN(n7339) );
  INV_X1 U8489 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7221) );
  OAI22_X1 U8490 ( .A1(n10040), .A2(n7507), .B1(n10740), .B2(n7221), .ZN(n7222) );
  AOI21_X1 U8491 ( .B1(n7227), .B2(n10740), .A(n7222), .ZN(n7223) );
  INV_X1 U8492 ( .A(n7223), .ZN(P1_U3462) );
  OAI22_X1 U8493 ( .A1(n9991), .A2(n7507), .B1(n10736), .B2(n6643), .ZN(n7226)
         );
  AOI21_X1 U8494 ( .B1(n7227), .B2(n10736), .A(n7226), .ZN(n7228) );
  INV_X1 U8495 ( .A(n7228), .ZN(P1_U3525) );
  INV_X1 U8496 ( .A(n7230), .ZN(n10590) );
  AND2_X1 U8497 ( .A1(n7276), .A2(n10590), .ZN(n7231) );
  OR2_X1 U8498 ( .A1(n7276), .A2(n10590), .ZN(n7232) );
  AND2_X1 U8499 ( .A1(n8713), .A2(n7277), .ZN(n7234) );
  OR2_X1 U8500 ( .A1(n8187), .A2(n7235), .ZN(n7238) );
  OR2_X1 U8501 ( .A1(n8208), .A2(n7236), .ZN(n7237) );
  OAI211_X1 U8502 ( .C1(n8249), .C2(n7326), .A(n7238), .B(n7237), .ZN(n7465)
         );
  INV_X1 U8503 ( .A(n7465), .ZN(n10614) );
  INV_X1 U8504 ( .A(n8312), .ZN(n7239) );
  XNOR2_X1 U8505 ( .A(n7468), .B(n7239), .ZN(n7240) );
  NAND2_X1 U8506 ( .A1(n7240), .A2(n8989), .ZN(n7248) );
  NAND2_X1 U8507 ( .A1(n7587), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7246) );
  NAND2_X1 U8508 ( .A1(n8183), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7245) );
  NAND2_X1 U8509 ( .A1(n7241), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7242) );
  NAND2_X1 U8510 ( .A1(n7371), .A2(n7242), .ZN(n7359) );
  NAND2_X1 U8511 ( .A1(n8159), .A2(n7359), .ZN(n7244) );
  NAND2_X1 U8512 ( .A1(n8291), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7243) );
  NAND4_X1 U8513 ( .A1(n7246), .A2(n7245), .A3(n7244), .A4(n7243), .ZN(n8711)
         );
  AOI22_X1 U8514 ( .A1(n8994), .A2(n8713), .B1(n8711), .B2(n8995), .ZN(n7247)
         );
  NAND2_X1 U8515 ( .A1(n7248), .A2(n7247), .ZN(n10615) );
  INV_X1 U8516 ( .A(n10615), .ZN(n7255) );
  INV_X2 U8517 ( .A(n10577), .ZN(n10580) );
  NAND2_X1 U8518 ( .A1(n7249), .A2(n8358), .ZN(n7273) );
  NAND2_X1 U8519 ( .A1(n7315), .A2(n7277), .ZN(n8365) );
  AND2_X1 U8520 ( .A1(n8365), .A2(n8361), .ZN(n8313) );
  OAI21_X1 U8521 ( .B1(n7250), .B2(n8312), .A(n7461), .ZN(n10617) );
  AOI22_X1 U8522 ( .A1(n9001), .A2(n7465), .B1(n8983), .B2(n7308), .ZN(n7251)
         );
  OAI21_X1 U8523 ( .B1(n7252), .B2(n10577), .A(n7251), .ZN(n7253) );
  AOI21_X1 U8524 ( .B1(n10617), .B2(n8950), .A(n7253), .ZN(n7254) );
  OAI21_X1 U8525 ( .B1(n7255), .B2(n10580), .A(n7254), .ZN(P2_U3227) );
  AOI22_X1 U8526 ( .A1(n9602), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10053), .ZN(n7256) );
  OAI21_X1 U8527 ( .B1(n8119), .B2(n8002), .A(n7256), .ZN(P1_U3337) );
  NAND2_X1 U8528 ( .A1(n7258), .A2(n7257), .ZN(n7260) );
  XNOR2_X1 U8529 ( .A(n7260), .B(n7259), .ZN(n7267) );
  INV_X1 U8530 ( .A(n7261), .ZN(n7390) );
  NAND2_X1 U8531 ( .A1(n7432), .A2(n10705), .ZN(n10607) );
  NOR2_X1 U8532 ( .A1(n7390), .A2(n10607), .ZN(n7262) );
  AOI211_X1 U8533 ( .C1(n8011), .C2(n9559), .A(n7263), .B(n7262), .ZN(n7266)
         );
  INV_X1 U8534 ( .A(n9275), .ZN(n9239) );
  AOI22_X1 U8535 ( .A1(n7264), .A2(n9560), .B1(n9239), .B2(n7434), .ZN(n7265)
         );
  OAI211_X1 U8536 ( .C1(n7267), .C2(n9284), .A(n7266), .B(n7265), .ZN(P1_U3227) );
  INV_X1 U8537 ( .A(n7268), .ZN(n7269) );
  NAND2_X1 U8538 ( .A1(n7269), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7270) );
  XNOR2_X1 U8539 ( .A(n7270), .B(P2_IR_REG_18__SCAN_IN), .ZN(n10510) );
  INV_X1 U8540 ( .A(n10510), .ZN(n10512) );
  OAI222_X1 U8541 ( .A1(n9159), .A2(n8119), .B1(n9156), .B2(n7271), .C1(
        P2_U3151), .C2(n10512), .ZN(P2_U3277) );
  OAI21_X1 U8542 ( .B1(n7273), .B2(n8313), .A(n7272), .ZN(n7487) );
  XOR2_X1 U8543 ( .A(n8313), .B(n7274), .Z(n7275) );
  OAI222_X1 U8544 ( .A1(n10564), .A2(n7276), .B1(n10566), .B2(n7471), .C1(
        n7275), .C2(n10562), .ZN(n7484) );
  AOI21_X1 U8545 ( .B1(n10720), .B2(n7487), .A(n7484), .ZN(n7281) );
  AOI22_X1 U8546 ( .A1(n9141), .A2(n7277), .B1(n10724), .B2(
        P2_REG0_REG_5__SCAN_IN), .ZN(n7278) );
  OAI21_X1 U8547 ( .B1(n7281), .B2(n10724), .A(n7278), .ZN(P2_U3405) );
  OAI22_X1 U8548 ( .A1(n9050), .A2(n7483), .B1(n10723), .B2(n5179), .ZN(n7279)
         );
  INV_X1 U8549 ( .A(n7279), .ZN(n7280) );
  OAI21_X1 U8550 ( .B1(n7281), .B2(n10721), .A(n7280), .ZN(P2_U3464) );
  INV_X1 U8551 ( .A(n8110), .ZN(n7288) );
  NAND2_X1 U8552 ( .A1(n7283), .A2(n7282), .ZN(n7284) );
  NAND2_X1 U8553 ( .A1(n7284), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7286) );
  XNOR2_X1 U8554 ( .A(n7286), .B(n7285), .ZN(n8819) );
  INV_X1 U8555 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7287) );
  OAI222_X1 U8556 ( .A1(n9159), .A2(n7288), .B1(n8819), .B2(P2_U3151), .C1(
        n7287), .C2(n9156), .ZN(P2_U3278) );
  INV_X1 U8557 ( .A(n9587), .ZN(n9578) );
  INV_X1 U8558 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7289) );
  OAI222_X1 U8559 ( .A1(P1_U3086), .A2(n9578), .B1(n10284), .B2(n7289), .C1(
        n7288), .C2(n8002), .ZN(P1_U3338) );
  OAI21_X1 U8560 ( .B1(n7292), .B2(n7291), .A(n7290), .ZN(n7298) );
  INV_X1 U8561 ( .A(n7514), .ZN(n7443) );
  OAI22_X1 U8562 ( .A1(n9278), .A2(n7443), .B1(n9242), .B2(n10622), .ZN(n7297)
         );
  INV_X1 U8563 ( .A(n9558), .ZN(n7660) );
  INV_X1 U8564 ( .A(n7293), .ZN(n7295) );
  OR2_X1 U8565 ( .A1(n9275), .A2(n7453), .ZN(n7294) );
  OAI211_X1 U8566 ( .C1(n9276), .C2(n7660), .A(n7295), .B(n7294), .ZN(n7296)
         );
  AOI211_X1 U8567 ( .C1(n7298), .C2(n9259), .A(n7297), .B(n7296), .ZN(n7299)
         );
  INV_X1 U8568 ( .A(n7299), .ZN(P1_U3239) );
  INV_X1 U8569 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10278) );
  INV_X1 U8570 ( .A(n8260), .ZN(n7300) );
  NAND2_X1 U8571 ( .A1(n7300), .A2(n8159), .ZN(n8296) );
  INV_X1 U8572 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n7303) );
  NAND2_X1 U8573 ( .A1(n7587), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7302) );
  NAND2_X1 U8574 ( .A1(n8291), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n7301) );
  OAI211_X1 U8575 ( .C1(n8215), .C2(n7303), .A(n7302), .B(n7301), .ZN(n7304)
         );
  INV_X1 U8576 ( .A(n7304), .ZN(n7305) );
  INV_X1 U8577 ( .A(n8846), .ZN(n7306) );
  NAND2_X1 U8578 ( .A1(n7306), .A2(P2_U3893), .ZN(n7307) );
  OAI21_X1 U8579 ( .B1(n10278), .B2(P2_U3893), .A(n7307), .ZN(P2_U3520) );
  INV_X1 U8580 ( .A(n7308), .ZN(n7320) );
  XNOR2_X1 U8581 ( .A(n7465), .B(n8552), .ZN(n7360) );
  XOR2_X1 U8582 ( .A(n8712), .B(n7360), .Z(n7313) );
  INV_X1 U8583 ( .A(n7309), .ZN(n7311) );
  AOI211_X1 U8584 ( .C1(n7313), .C2(n7312), .A(n8683), .B(n7363), .ZN(n7314)
         );
  INV_X1 U8585 ( .A(n7314), .ZN(n7319) );
  INV_X1 U8586 ( .A(n8711), .ZN(n7569) );
  OAI22_X1 U8587 ( .A1(n7315), .A2(n8691), .B1(n7569), .B2(n8679), .ZN(n7316)
         );
  AOI211_X1 U8588 ( .C1(n7465), .C2(n8681), .A(n7317), .B(n7316), .ZN(n7318)
         );
  OAI211_X1 U8589 ( .C1(n7320), .C2(n7381), .A(n7319), .B(n7318), .ZN(P2_U3179) );
  INV_X1 U8590 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7476) );
  OR2_X1 U8591 ( .A1(n8825), .A2(n7476), .ZN(n7322) );
  NAND2_X1 U8592 ( .A1(n8825), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7321) );
  NAND2_X1 U8593 ( .A1(n7322), .A2(n7321), .ZN(n7397) );
  XOR2_X1 U8594 ( .A(n7393), .B(n7397), .Z(n7399) );
  OAI21_X1 U8595 ( .B1(n7324), .B2(n7326), .A(n7323), .ZN(n7400) );
  XOR2_X1 U8596 ( .A(n7399), .B(n7400), .Z(n7336) );
  XNOR2_X1 U8597 ( .A(n7394), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n7334) );
  NAND2_X1 U8598 ( .A1(n7328), .A2(n7476), .ZN(n7329) );
  AOI21_X1 U8599 ( .B1(n7410), .B2(n7329), .A(n10489), .ZN(n7333) );
  NAND2_X1 U8600 ( .A1(n10476), .A2(n5318), .ZN(n7331) );
  NOR2_X1 U8601 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6977), .ZN(n7378) );
  AOI21_X1 U8602 ( .B1(n10498), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7378), .ZN(
        n7330) );
  NAND2_X1 U8603 ( .A1(n7331), .A2(n7330), .ZN(n7332) );
  AOI211_X1 U8604 ( .C1(n7334), .C2(n10483), .A(n7333), .B(n7332), .ZN(n7335)
         );
  OAI21_X1 U8605 ( .B1(n7336), .B2(n8830), .A(n7335), .ZN(P2_U3189) );
  OAI21_X1 U8606 ( .B1(n7338), .B2(n9356), .A(n7337), .ZN(n10551) );
  INV_X1 U8607 ( .A(n10551), .ZN(n7358) );
  NAND3_X1 U8608 ( .A1(n7341), .A2(n7340), .A3(n7339), .ZN(n7343) );
  AND2_X1 U8609 ( .A1(n10525), .A2(n7344), .ZN(n7976) );
  INV_X1 U8610 ( .A(n7976), .ZN(n7794) );
  INV_X1 U8611 ( .A(n9852), .ZN(n10529) );
  INV_X1 U8612 ( .A(n7786), .ZN(n7968) );
  OAI22_X1 U8613 ( .A1(n7345), .A2(n10631), .B1(n7524), .B2(n9880), .ZN(n7346)
         );
  AOI21_X1 U8614 ( .B1(n10551), .B2(n7968), .A(n7346), .ZN(n7347) );
  OAI21_X1 U8615 ( .B1(n10529), .B2(n7348), .A(n7347), .ZN(n10549) );
  NAND2_X1 U8616 ( .A1(n10549), .A2(n10525), .ZN(n7357) );
  INV_X1 U8617 ( .A(n7349), .ZN(n7350) );
  OAI22_X1 U8618 ( .A1(n10525), .A2(n5672), .B1(n7351), .B2(n10522), .ZN(n7355) );
  INV_X1 U8619 ( .A(n7498), .ZN(n7353) );
  OAI211_X1 U8620 ( .C1(n7353), .C2(n10548), .A(n9884), .B(n7352), .ZN(n10547)
         );
  NOR2_X1 U8621 ( .A1(n9865), .A2(n10547), .ZN(n7354) );
  AOI211_X1 U8622 ( .C1(n9869), .C2(n6879), .A(n7355), .B(n7354), .ZN(n7356)
         );
  OAI211_X1 U8623 ( .C1(n7358), .C2(n7794), .A(n7357), .B(n7356), .ZN(P1_U3291) );
  INV_X1 U8624 ( .A(n7359), .ZN(n7475) );
  INV_X1 U8625 ( .A(n7360), .ZN(n7361) );
  OR2_X1 U8626 ( .A1(n8208), .A2(n7365), .ZN(n7366) );
  XOR2_X1 U8627 ( .A(n8552), .B(n7478), .Z(n7367) );
  NOR2_X1 U8628 ( .A1(n7367), .A2(n8711), .ZN(n7605) );
  AOI21_X1 U8629 ( .B1(n7367), .B2(n8711), .A(n7605), .ZN(n7368) );
  OAI21_X1 U8630 ( .B1(n7369), .B2(n7368), .A(n7607), .ZN(n7370) );
  NAND2_X1 U8631 ( .A1(n7370), .A2(n8685), .ZN(n7380) );
  NAND2_X1 U8632 ( .A1(n7587), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7376) );
  NAND2_X1 U8633 ( .A1(n8183), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7375) );
  NAND2_X1 U8634 ( .A1(n7371), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7372) );
  NAND2_X1 U8635 ( .A1(n7574), .A2(n7372), .ZN(n7638) );
  NAND2_X1 U8636 ( .A1(n8159), .A2(n7638), .ZN(n7374) );
  NAND2_X1 U8637 ( .A1(n8291), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7373) );
  NAND4_X1 U8638 ( .A1(n7376), .A2(n7375), .A3(n7374), .A4(n7373), .ZN(n8710)
         );
  OAI22_X1 U8639 ( .A1(n7731), .A2(n8679), .B1(n8697), .B2(n10638), .ZN(n7377)
         );
  AOI211_X1 U8640 ( .C1(n8676), .C2(n8712), .A(n7378), .B(n7377), .ZN(n7379)
         );
  OAI211_X1 U8641 ( .C1(n7475), .C2(n7381), .A(n7380), .B(n7379), .ZN(P2_U3153) );
  NAND2_X1 U8642 ( .A1(n7566), .A2(n10705), .ZN(n10629) );
  OAI21_X1 U8643 ( .B1(n7384), .B2(n7383), .A(n7382), .ZN(n7385) );
  NAND2_X1 U8644 ( .A1(n7385), .A2(n9259), .ZN(n7389) );
  OAI22_X1 U8645 ( .A1(n9278), .A2(n10632), .B1(n9275), .B2(n7559), .ZN(n7386)
         );
  AOI211_X1 U8646 ( .C1(n8011), .C2(n10661), .A(n7387), .B(n7386), .ZN(n7388)
         );
  OAI211_X1 U8647 ( .C1(n7390), .C2(n10629), .A(n7389), .B(n7388), .ZN(
        P1_U3213) );
  INV_X1 U8648 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10658) );
  MUX2_X1 U8649 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10658), .S(n7571), .Z(n7396)
         );
  INV_X1 U8650 ( .A(n7391), .ZN(n7392) );
  AOI22_X1 U8651 ( .A1(n7394), .A2(P2_REG1_REG_7__SCAN_IN), .B1(n7393), .B2(
        n7392), .ZN(n7395) );
  AOI21_X1 U8652 ( .B1(n7396), .B2(n7395), .A(n7536), .ZN(n7416) );
  INV_X1 U8653 ( .A(n7397), .ZN(n7398) );
  AOI22_X1 U8654 ( .A1(n7400), .A2(n7399), .B1(n5318), .B2(n7398), .ZN(n7530)
         );
  INV_X1 U8655 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7640) );
  OR2_X1 U8656 ( .A1(n8825), .A2(n7640), .ZN(n7402) );
  NAND2_X1 U8657 ( .A1(n8825), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7401) );
  NAND2_X1 U8658 ( .A1(n7402), .A2(n7401), .ZN(n7528) );
  XOR2_X1 U8659 ( .A(n7571), .B(n7528), .Z(n7529) );
  XNOR2_X1 U8660 ( .A(n7530), .B(n7529), .ZN(n7403) );
  NAND2_X1 U8661 ( .A1(n7403), .A2(n10513), .ZN(n7415) );
  INV_X1 U8662 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7405) );
  INV_X1 U8663 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10128) );
  NOR2_X1 U8664 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10128), .ZN(n7612) );
  INV_X1 U8665 ( .A(n7612), .ZN(n7404) );
  OAI21_X1 U8666 ( .B1(n8738), .B2(n7405), .A(n7404), .ZN(n7413) );
  NAND2_X1 U8667 ( .A1(n7410), .A2(n7408), .ZN(n7406) );
  XNOR2_X1 U8668 ( .A(n7571), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7407) );
  NAND2_X1 U8669 ( .A1(n7406), .A2(n7407), .ZN(n7540) );
  INV_X1 U8670 ( .A(n7407), .ZN(n7409) );
  NAND3_X1 U8671 ( .A1(n7410), .A2(n7409), .A3(n7408), .ZN(n7411) );
  AOI21_X1 U8672 ( .B1(n7540), .B2(n7411), .A(n10489), .ZN(n7412) );
  AOI211_X1 U8673 ( .C1(n10476), .C2(n7571), .A(n7413), .B(n7412), .ZN(n7414)
         );
  OAI211_X1 U8674 ( .C1(n7416), .C2(n10496), .A(n7415), .B(n7414), .ZN(
        P2_U3190) );
  INV_X1 U8675 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7417) );
  INV_X1 U8676 ( .A(n8130), .ZN(n7419) );
  OAI222_X1 U8677 ( .A1(n10285), .A2(n7417), .B1(n8002), .B2(n7419), .C1(
        P1_U3086), .C2(n5608), .ZN(P1_U3336) );
  INV_X1 U8678 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7420) );
  OAI222_X1 U8679 ( .A1(n9156), .A2(n7420), .B1(n9159), .B2(n7419), .C1(n7418), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  NAND2_X1 U8680 ( .A1(n7524), .A2(n7507), .ZN(n7421) );
  OAI21_X1 U8681 ( .B1(n7517), .B2(n7522), .A(n10609), .ZN(n7424) );
  NAND2_X1 U8682 ( .A1(n7517), .A2(n7522), .ZN(n7423) );
  NAND2_X1 U8683 ( .A1(n7424), .A2(n7423), .ZN(n7441) );
  NAND2_X1 U8684 ( .A1(n7443), .A2(n7432), .ZN(n9306) );
  INV_X1 U8685 ( .A(n7432), .ZN(n7442) );
  NAND2_X1 U8686 ( .A1(n9306), .A2(n9403), .ZN(n9407) );
  XNOR2_X1 U8687 ( .A(n7441), .B(n9407), .ZN(n10606) );
  INV_X1 U8688 ( .A(n10606), .ZN(n7440) );
  AND2_X1 U8689 ( .A1(n9394), .A2(n7426), .ZN(n9302) );
  NAND2_X1 U8690 ( .A1(n9304), .A2(n9302), .ZN(n7428) );
  INV_X1 U8691 ( .A(n9309), .ZN(n9396) );
  NOR2_X1 U8692 ( .A1(n9560), .A2(n7522), .ZN(n9305) );
  NOR2_X1 U8693 ( .A1(n9396), .A2(n9305), .ZN(n7427) );
  NAND2_X1 U8694 ( .A1(n9560), .A2(n7522), .ZN(n9395) );
  INV_X1 U8695 ( .A(n9395), .ZN(n9310) );
  XNOR2_X1 U8696 ( .A(n7446), .B(n9407), .ZN(n7429) );
  NAND2_X1 U8697 ( .A1(n7429), .A2(n9852), .ZN(n7431) );
  NAND2_X1 U8698 ( .A1(n9559), .A2(n10519), .ZN(n7430) );
  NAND2_X1 U8699 ( .A1(n7431), .A2(n7430), .ZN(n10612) );
  NAND2_X1 U8700 ( .A1(n7523), .A2(n7522), .ZN(n7521) );
  AOI21_X1 U8701 ( .B1(n7521), .B2(n7432), .A(n9826), .ZN(n7433) );
  OR2_X1 U8702 ( .A1(n7521), .A2(n7432), .ZN(n7450) );
  NAND2_X1 U8703 ( .A1(n7433), .A2(n7450), .ZN(n10608) );
  AND2_X1 U8704 ( .A1(n10525), .A2(n10704), .ZN(n9677) );
  INV_X1 U8705 ( .A(n10525), .ZN(n9859) );
  INV_X1 U8706 ( .A(n10522), .ZN(n9857) );
  AOI22_X1 U8707 ( .A1(n9859), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7434), .B2(
        n9857), .ZN(n7435) );
  OAI21_X1 U8708 ( .B1(n7442), .B2(n9888), .A(n7435), .ZN(n7436) );
  AOI21_X1 U8709 ( .B1(n9677), .B2(n9560), .A(n7436), .ZN(n7437) );
  OAI21_X1 U8710 ( .B1(n9865), .B2(n10608), .A(n7437), .ZN(n7438) );
  AOI21_X1 U8711 ( .B1(n10612), .B2(n10525), .A(n7438), .ZN(n7439) );
  OAI21_X1 U8712 ( .B1(n7440), .B2(n9894), .A(n7439), .ZN(P1_U3288) );
  NAND2_X1 U8713 ( .A1(n7441), .A2(n9407), .ZN(n7445) );
  NAND2_X1 U8714 ( .A1(n7443), .A2(n7442), .ZN(n7444) );
  NAND2_X1 U8715 ( .A1(n10632), .A2(n7456), .ZN(n9409) );
  NAND2_X1 U8716 ( .A1(n9559), .A2(n10622), .ZN(n9410) );
  XNOR2_X1 U8717 ( .A(n7551), .B(n9400), .ZN(n10625) );
  INV_X1 U8718 ( .A(n10625), .ZN(n7460) );
  XNOR2_X1 U8719 ( .A(n7553), .B(n9400), .ZN(n7447) );
  NAND2_X1 U8720 ( .A1(n7447), .A2(n9852), .ZN(n7449) );
  AOI22_X1 U8721 ( .A1(n10704), .A2(n7514), .B1(n9558), .B2(n10519), .ZN(n7448) );
  NAND2_X1 U8722 ( .A1(n7449), .A2(n7448), .ZN(n10623) );
  INV_X1 U8723 ( .A(n7450), .ZN(n7452) );
  INV_X1 U8724 ( .A(n7562), .ZN(n7451) );
  OAI211_X1 U8725 ( .C1(n10622), .C2(n7452), .A(n7451), .B(n9884), .ZN(n10621)
         );
  OAI22_X1 U8726 ( .A1(n10525), .A2(n7454), .B1(n7453), .B2(n10522), .ZN(n7455) );
  AOI21_X1 U8727 ( .B1(n9869), .B2(n7456), .A(n7455), .ZN(n7457) );
  OAI21_X1 U8728 ( .B1(n10621), .B2(n9865), .A(n7457), .ZN(n7458) );
  AOI21_X1 U8729 ( .B1(n10623), .B2(n10525), .A(n7458), .ZN(n7459) );
  OAI21_X1 U8730 ( .B1(n7460), .B2(n9894), .A(n7459), .ZN(P1_U3287) );
  NAND2_X1 U8731 ( .A1(n7569), .A2(n7478), .ZN(n8378) );
  NAND2_X1 U8732 ( .A1(n8711), .A2(n10638), .ZN(n7643) );
  NAND2_X1 U8733 ( .A1(n7462), .A2(n8315), .ZN(n7463) );
  NAND2_X1 U8734 ( .A1(n7600), .A2(n7463), .ZN(n10639) );
  NOR2_X1 U8735 ( .A1(n10580), .A2(n7464), .ZN(n8263) );
  INV_X1 U8736 ( .A(n8263), .ZN(n7481) );
  NOR2_X1 U8737 ( .A1(n8712), .A2(n7465), .ZN(n7467) );
  NAND2_X1 U8738 ( .A1(n8712), .A2(n7465), .ZN(n7466) );
  OAI21_X1 U8739 ( .B1(n7470), .B2(n8315), .A(n7634), .ZN(n7473) );
  OAI22_X1 U8740 ( .A1(n7471), .A2(n10564), .B1(n7731), .B2(n10566), .ZN(n7472) );
  AOI21_X1 U8741 ( .B1(n7473), .B2(n8989), .A(n7472), .ZN(n7474) );
  OAI21_X1 U8742 ( .B1(n8256), .B2(n10639), .A(n7474), .ZN(n10641) );
  NAND2_X1 U8743 ( .A1(n10641), .A2(n10577), .ZN(n7480) );
  OAI22_X1 U8744 ( .A1(n10577), .A2(n7476), .B1(n7475), .B2(n10570), .ZN(n7477) );
  AOI21_X1 U8745 ( .B1(n9001), .B2(n7478), .A(n7477), .ZN(n7479) );
  OAI211_X1 U8746 ( .C1(n10639), .C2(n7481), .A(n7480), .B(n7479), .ZN(
        P2_U3226) );
  OAI22_X1 U8747 ( .A1(n8937), .A2(n7483), .B1(n7482), .B2(n10570), .ZN(n7486)
         );
  MUX2_X1 U8748 ( .A(n7484), .B(P2_REG2_REG_5__SCAN_IN), .S(n10580), .Z(n7485)
         );
  AOI211_X1 U8749 ( .C1(n8950), .C2(n7487), .A(n7486), .B(n7485), .ZN(n7488)
         );
  INV_X1 U8750 ( .A(n7488), .ZN(P2_U3228) );
  INV_X1 U8751 ( .A(n9363), .ZN(n7489) );
  XNOR2_X1 U8752 ( .A(n5098), .B(n7489), .ZN(n7491) );
  AND2_X1 U8753 ( .A1(n5692), .A2(n10519), .ZN(n7490) );
  AOI21_X1 U8754 ( .B1(n7491), .B2(n9852), .A(n7490), .ZN(n10543) );
  OAI21_X1 U8755 ( .B1(n5098), .B2(n7493), .A(n7492), .ZN(n10541) );
  AOI22_X1 U8756 ( .A1(n9685), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9857), .ZN(n7495) );
  OAI21_X1 U8757 ( .B1(n10539), .B2(n9888), .A(n7495), .ZN(n7501) );
  INV_X1 U8758 ( .A(n6474), .ZN(n7499) );
  NAND2_X1 U8759 ( .A1(n7496), .A2(n10533), .ZN(n7497) );
  NAND3_X1 U8760 ( .A1(n7498), .A2(n9884), .A3(n7497), .ZN(n10537) );
  OAI22_X1 U8761 ( .A1(n7499), .A2(n9861), .B1(n9865), .B2(n10537), .ZN(n7500)
         );
  AOI211_X1 U8762 ( .C1(n9855), .C2(n10541), .A(n7501), .B(n7500), .ZN(n7502)
         );
  OAI21_X1 U8763 ( .B1(n9685), .B2(n10543), .A(n7502), .ZN(P1_U3292) );
  AOI22_X1 U8764 ( .A1(n7503), .A2(n9891), .B1(n9677), .B2(n5692), .ZN(n7506)
         );
  INV_X1 U8765 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7504) );
  AOI22_X1 U8766 ( .A1(n9685), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9857), .B2(
        n7504), .ZN(n7505) );
  OAI211_X1 U8767 ( .C1(n7507), .C2(n9888), .A(n7506), .B(n7505), .ZN(n7508)
         );
  AOI21_X1 U8768 ( .B1(n7509), .B2(n9855), .A(n7508), .ZN(n7510) );
  OAI21_X1 U8769 ( .B1(n9685), .B2(n7511), .A(n7510), .ZN(P1_U3290) );
  NAND2_X1 U8770 ( .A1(n7512), .A2(n9309), .ZN(n7513) );
  OR2_X1 U8771 ( .A1(n9310), .A2(n9305), .ZN(n7516) );
  INV_X1 U8772 ( .A(n7516), .ZN(n9360) );
  XNOR2_X1 U8773 ( .A(n7513), .B(n9360), .ZN(n7515) );
  AOI22_X1 U8774 ( .A1(n7515), .A2(n9852), .B1(n10519), .B2(n7514), .ZN(n10601) );
  XNOR2_X1 U8775 ( .A(n7517), .B(n7516), .ZN(n10603) );
  INV_X1 U8776 ( .A(n7518), .ZN(n7519) );
  AOI22_X1 U8777 ( .A1(n9685), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7519), .B2(
        n9857), .ZN(n7520) );
  OAI21_X1 U8778 ( .B1(n7522), .B2(n9888), .A(n7520), .ZN(n7526) );
  OAI211_X1 U8779 ( .C1(n7523), .C2(n7522), .A(n7521), .B(n9884), .ZN(n10599)
         );
  OAI22_X1 U8780 ( .A1(n10599), .A2(n9865), .B1(n7524), .B2(n9861), .ZN(n7525)
         );
  AOI211_X1 U8781 ( .C1(n10603), .C2(n9855), .A(n7526), .B(n7525), .ZN(n7527)
         );
  OAI21_X1 U8782 ( .B1(n10601), .B2(n9685), .A(n7527), .ZN(P1_U3289) );
  OAI22_X1 U8783 ( .A1(n7530), .A2(n7529), .B1(n7537), .B2(n7528), .ZN(n8720)
         );
  OR2_X1 U8784 ( .A1(n8825), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7532) );
  INV_X1 U8785 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10676) );
  NAND2_X1 U8786 ( .A1(n8825), .A2(n10676), .ZN(n7531) );
  AND2_X1 U8787 ( .A1(n7532), .A2(n7531), .ZN(n7533) );
  NOR2_X1 U8788 ( .A1(n7533), .A2(n8742), .ZN(n8718) );
  INV_X1 U8789 ( .A(n8718), .ZN(n7534) );
  NAND2_X1 U8790 ( .A1(n7533), .A2(n8742), .ZN(n8719) );
  NAND2_X1 U8791 ( .A1(n7534), .A2(n8719), .ZN(n7535) );
  XNOR2_X1 U8792 ( .A(n8720), .B(n7535), .ZN(n7550) );
  NAND2_X1 U8793 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n7538), .ZN(n8743) );
  OAI21_X1 U8794 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n7538), .A(n8743), .ZN(
        n7548) );
  OR2_X1 U8795 ( .A1(n7571), .A2(n7640), .ZN(n7539) );
  INV_X1 U8796 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7598) );
  AOI21_X1 U8797 ( .B1(n7542), .B2(n7598), .A(n8729), .ZN(n7546) );
  INV_X1 U8798 ( .A(n8742), .ZN(n7581) );
  NOR2_X1 U8799 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6979), .ZN(n7737) );
  INV_X1 U8800 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7543) );
  NOR2_X1 U8801 ( .A1(n8738), .A2(n7543), .ZN(n7544) );
  AOI211_X1 U8802 ( .C1(n10476), .C2(n7581), .A(n7737), .B(n7544), .ZN(n7545)
         );
  OAI21_X1 U8803 ( .B1(n7546), .B2(n10489), .A(n7545), .ZN(n7547) );
  AOI21_X1 U8804 ( .B1(n7548), .B2(n10483), .A(n7547), .ZN(n7549) );
  OAI21_X1 U8805 ( .B1(n7550), .B2(n8830), .A(n7549), .ZN(P2_U3191) );
  NAND2_X1 U8806 ( .A1(n10632), .A2(n10622), .ZN(n7552) );
  NAND2_X1 U8807 ( .A1(n7660), .A2(n7566), .ZN(n7711) );
  INV_X1 U8808 ( .A(n7566), .ZN(n7659) );
  NAND2_X1 U8809 ( .A1(n7659), .A2(n9558), .ZN(n9416) );
  NAND2_X1 U8810 ( .A1(n7711), .A2(n9416), .ZN(n7657) );
  INV_X1 U8811 ( .A(n7657), .ZN(n9412) );
  XNOR2_X1 U8812 ( .A(n7658), .B(n9412), .ZN(n10628) );
  INV_X1 U8813 ( .A(n10661), .ZN(n7698) );
  INV_X1 U8814 ( .A(n9410), .ZN(n7554) );
  NOR2_X1 U8815 ( .A1(n7657), .A2(n7554), .ZN(n7555) );
  NAND2_X1 U8816 ( .A1(n7710), .A2(n7555), .ZN(n7685) );
  INV_X1 U8817 ( .A(n7685), .ZN(n7557) );
  AOI21_X1 U8818 ( .B1(n7710), .B2(n9410), .A(n9412), .ZN(n7556) );
  NOR2_X1 U8819 ( .A1(n7557), .A2(n7556), .ZN(n7558) );
  OAI222_X1 U8820 ( .A1(n9880), .A2(n7698), .B1(n7786), .B2(n10628), .C1(
        n10529), .C2(n7558), .ZN(n10633) );
  NAND2_X1 U8821 ( .A1(n10633), .A2(n10525), .ZN(n7568) );
  INV_X1 U8822 ( .A(n7559), .ZN(n7560) );
  AOI22_X1 U8823 ( .A1(n9859), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7560), .B2(
        n9857), .ZN(n7561) );
  OAI21_X1 U8824 ( .B1(n9861), .B2(n10632), .A(n7561), .ZN(n7565) );
  OAI21_X1 U8825 ( .B1(n7562), .B2(n7659), .A(n9884), .ZN(n7563) );
  OR2_X1 U8826 ( .A1(n7563), .A2(n7668), .ZN(n10630) );
  NOR2_X1 U8827 ( .A1(n10630), .A2(n9865), .ZN(n7564) );
  AOI211_X1 U8828 ( .C1(n9869), .C2(n7566), .A(n7565), .B(n7564), .ZN(n7567)
         );
  OAI211_X1 U8829 ( .C1(n10628), .C2(n7794), .A(n7568), .B(n7567), .ZN(
        P1_U3286) );
  NAND2_X1 U8830 ( .A1(n7569), .A2(n10638), .ZN(n7633) );
  NAND2_X1 U8831 ( .A1(n7570), .A2(n8288), .ZN(n7573) );
  AOI22_X1 U8832 ( .A1(n8132), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8131), .B2(
        n7571), .ZN(n7572) );
  NAND2_X1 U8833 ( .A1(n7573), .A2(n7572), .ZN(n7642) );
  NAND2_X1 U8834 ( .A1(n7731), .A2(n7642), .ZN(n8379) );
  INV_X1 U8835 ( .A(n7642), .ZN(n10655) );
  NAND2_X1 U8836 ( .A1(n10655), .A2(n8710), .ZN(n8375) );
  NAND2_X1 U8837 ( .A1(n8379), .A2(n8375), .ZN(n7644) );
  NAND2_X1 U8838 ( .A1(n7731), .A2(n10655), .ZN(n7585) );
  NAND2_X1 U8839 ( .A1(n7636), .A2(n7585), .ZN(n7584) );
  NAND2_X1 U8840 ( .A1(n8291), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7579) );
  NAND2_X1 U8841 ( .A1(n7587), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7578) );
  NAND2_X1 U8842 ( .A1(n7574), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7575) );
  NAND2_X1 U8843 ( .A1(n7588), .A2(n7575), .ZN(n7740) );
  NAND2_X1 U8844 ( .A1(n8159), .A2(n7740), .ZN(n7577) );
  NAND2_X1 U8845 ( .A1(n8183), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7576) );
  NAND4_X1 U8846 ( .A1(n7579), .A2(n7578), .A3(n7577), .A4(n7576), .ZN(n8709)
         );
  NAND2_X1 U8847 ( .A1(n7580), .A2(n8288), .ZN(n7583) );
  AOI22_X1 U8848 ( .A1(n8132), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8131), .B2(
        n7581), .ZN(n7582) );
  NAND2_X1 U8849 ( .A1(n7583), .A2(n7582), .ZN(n10672) );
  NAND2_X1 U8850 ( .A1(n10672), .A2(n7883), .ZN(n8380) );
  NAND2_X1 U8851 ( .A1(n8392), .A2(n8380), .ZN(n7759) );
  NAND2_X1 U8852 ( .A1(n7584), .A2(n7759), .ZN(n7765) );
  INV_X1 U8853 ( .A(n7759), .ZN(n8320) );
  NAND3_X1 U8854 ( .A1(n7636), .A2(n8320), .A3(n7585), .ZN(n7586) );
  NAND2_X1 U8855 ( .A1(n7765), .A2(n7586), .ZN(n7596) );
  NAND2_X1 U8856 ( .A1(n7587), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7593) );
  NAND2_X1 U8857 ( .A1(n8291), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7592) );
  NAND2_X1 U8858 ( .A1(n7588), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7589) );
  NAND2_X1 U8859 ( .A1(n7767), .A2(n7589), .ZN(n7897) );
  NAND2_X1 U8860 ( .A1(n8159), .A2(n7897), .ZN(n7591) );
  NAND2_X1 U8861 ( .A1(n8183), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7590) );
  NAND2_X1 U8862 ( .A1(n8710), .A2(n8994), .ZN(n7594) );
  OAI21_X1 U8863 ( .B1(n7893), .B2(n10566), .A(n7594), .ZN(n7595) );
  AOI21_X1 U8864 ( .B1(n7596), .B2(n8989), .A(n7595), .ZN(n10675) );
  INV_X1 U8865 ( .A(n7740), .ZN(n7597) );
  OAI22_X1 U8866 ( .A1(n10577), .A2(n7598), .B1(n7597), .B2(n10570), .ZN(n7599) );
  AOI21_X1 U8867 ( .B1(n9001), .B2(n10672), .A(n7599), .ZN(n7603) );
  AND2_X1 U8868 ( .A1(n8375), .A2(n7643), .ZN(n8390) );
  NAND2_X1 U8869 ( .A1(n7600), .A2(n8390), .ZN(n7601) );
  NAND2_X1 U8870 ( .A1(n10670), .A2(n8950), .ZN(n7602) );
  OAI211_X1 U8871 ( .C1(n10675), .C2(n10580), .A(n7603), .B(n7602), .ZN(
        P2_U3224) );
  INV_X1 U8872 ( .A(n7607), .ZN(n7604) );
  XNOR2_X1 U8873 ( .A(n7642), .B(n8552), .ZN(n7730) );
  XNOR2_X1 U8874 ( .A(n7730), .B(n8710), .ZN(n7608) );
  NOR3_X1 U8875 ( .A1(n7604), .A2(n7605), .A3(n7608), .ZN(n7611) );
  INV_X1 U8876 ( .A(n7605), .ZN(n7606) );
  NAND2_X1 U8877 ( .A1(n7607), .A2(n7606), .ZN(n7609) );
  INV_X1 U8878 ( .A(n7733), .ZN(n7610) );
  OAI21_X1 U8879 ( .B1(n7611), .B2(n7610), .A(n8685), .ZN(n7616) );
  AOI21_X1 U8880 ( .B1(n8711), .B2(n8676), .A(n7612), .ZN(n7613) );
  OAI21_X1 U8881 ( .B1(n7883), .B2(n8679), .A(n7613), .ZN(n7614) );
  AOI21_X1 U8882 ( .B1(n8694), .B2(n7638), .A(n7614), .ZN(n7615) );
  OAI211_X1 U8883 ( .C1(n10655), .C2(n8697), .A(n7616), .B(n7615), .ZN(
        P2_U3161) );
  MUX2_X1 U8884 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7617), .S(n7624), .Z(n7621)
         );
  OAI21_X1 U8885 ( .B1(n7619), .B2(n7164), .A(n7618), .ZN(n7620) );
  NAND2_X1 U8886 ( .A1(n7620), .A2(n7621), .ZN(n7750) );
  OAI211_X1 U8887 ( .C1(n7621), .C2(n7620), .A(n9582), .B(n7750), .ZN(n7632)
         );
  NAND2_X1 U8888 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9166) );
  INV_X1 U8889 ( .A(n9166), .ZN(n7630) );
  NAND2_X1 U8890 ( .A1(n7624), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7747) );
  OR2_X1 U8891 ( .A1(n7624), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7625) );
  NAND2_X1 U8892 ( .A1(n7747), .A2(n7625), .ZN(n7627) );
  INV_X1 U8893 ( .A(n7748), .ZN(n7626) );
  AOI211_X1 U8894 ( .C1(n7628), .C2(n7627), .A(n7626), .B(n9590), .ZN(n7629)
         );
  AOI211_X1 U8895 ( .C1(n10350), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n7630), .B(
        n7629), .ZN(n7631) );
  OAI211_X1 U8896 ( .C1(n10360), .C2(n7751), .A(n7632), .B(n7631), .ZN(
        P1_U3257) );
  INV_X1 U8897 ( .A(n7644), .ZN(n8319) );
  NAND3_X1 U8898 ( .A1(n7634), .A2(n8319), .A3(n7633), .ZN(n7635) );
  NAND2_X1 U8899 ( .A1(n7636), .A2(n7635), .ZN(n7637) );
  AOI222_X1 U8900 ( .A1(n8989), .A2(n7637), .B1(n8709), .B2(n8995), .C1(n8711), 
        .C2(n8994), .ZN(n10654) );
  INV_X1 U8901 ( .A(n7638), .ZN(n7639) );
  OAI22_X1 U8902 ( .A1(n10577), .A2(n7640), .B1(n7639), .B2(n10570), .ZN(n7641) );
  AOI21_X1 U8903 ( .B1(n9001), .B2(n7642), .A(n7641), .ZN(n7647) );
  NAND2_X1 U8904 ( .A1(n7600), .A2(n7643), .ZN(n7645) );
  XNOR2_X1 U8905 ( .A(n7645), .B(n7644), .ZN(n10657) );
  NAND2_X1 U8906 ( .A1(n10657), .A2(n8950), .ZN(n7646) );
  OAI211_X1 U8907 ( .C1(n10654), .C2(n10580), .A(n7647), .B(n7646), .ZN(
        P2_U3225) );
  NAND2_X1 U8908 ( .A1(n7648), .A2(n7649), .ZN(n7651) );
  XNOR2_X1 U8909 ( .A(n7651), .B(n7650), .ZN(n7656) );
  OAI22_X1 U8910 ( .A1(n9278), .A2(n7660), .B1(n9275), .B2(n7666), .ZN(n7652)
         );
  AOI211_X1 U8911 ( .C1(n8011), .C2(n10679), .A(n7653), .B(n7652), .ZN(n7655)
         );
  NAND2_X1 U8912 ( .A1(n9281), .A2(n7676), .ZN(n7654) );
  OAI211_X1 U8913 ( .C1(n7656), .C2(n9284), .A(n7655), .B(n7654), .ZN(P1_U3221) );
  NAND2_X1 U8914 ( .A1(n7660), .A2(n7659), .ZN(n7661) );
  NAND2_X1 U8915 ( .A1(n7676), .A2(n7698), .ZN(n9419) );
  NAND2_X1 U8916 ( .A1(n7708), .A2(n9419), .ZN(n9418) );
  XNOR2_X1 U8917 ( .A(n7675), .B(n9418), .ZN(n10645) );
  INV_X1 U8918 ( .A(n10645), .ZN(n7673) );
  NAND2_X1 U8919 ( .A1(n7685), .A2(n7711), .ZN(n7662) );
  XNOR2_X1 U8920 ( .A(n7662), .B(n9418), .ZN(n7665) );
  NAND2_X1 U8921 ( .A1(n10645), .A2(n7968), .ZN(n7664) );
  AOI22_X1 U8922 ( .A1(n10704), .A2(n9558), .B1(n10679), .B2(n10519), .ZN(
        n7663) );
  OAI211_X1 U8923 ( .C1(n7665), .C2(n10529), .A(n7664), .B(n7663), .ZN(n10650)
         );
  NAND2_X1 U8924 ( .A1(n10650), .A2(n10525), .ZN(n7672) );
  OAI22_X1 U8925 ( .A1(n10525), .A2(n7667), .B1(n7666), .B2(n10522), .ZN(n7670) );
  INV_X1 U8926 ( .A(n7676), .ZN(n10648) );
  OAI211_X1 U8927 ( .C1(n7668), .C2(n10648), .A(n9884), .B(n7718), .ZN(n10646)
         );
  NOR2_X1 U8928 ( .A1(n10646), .A2(n9865), .ZN(n7669) );
  AOI211_X1 U8929 ( .C1(n9869), .C2(n7676), .A(n7670), .B(n7669), .ZN(n7671)
         );
  OAI211_X1 U8930 ( .C1(n7673), .C2(n7794), .A(n7672), .B(n7671), .ZN(P1_U3285) );
  INV_X1 U8931 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8154) );
  OAI222_X1 U8932 ( .A1(n9159), .A2(n8153), .B1(P2_U3151), .B2(n7674), .C1(
        n8154), .C2(n9156), .ZN(P2_U3274) );
  INV_X1 U8933 ( .A(n10679), .ZN(n7825) );
  OR2_X1 U8934 ( .A1(n10662), .A2(n7825), .ZN(n9426) );
  NAND2_X1 U8935 ( .A1(n10662), .A2(n7825), .ZN(n9429) );
  NAND2_X1 U8936 ( .A1(n9426), .A2(n9429), .ZN(n7704) );
  XNOR2_X1 U8937 ( .A(n7705), .B(n7704), .ZN(n10667) );
  INV_X1 U8938 ( .A(n10662), .ZN(n7677) );
  XNOR2_X1 U8939 ( .A(n7718), .B(n7677), .ZN(n7679) );
  AND2_X1 U8940 ( .A1(n9557), .A2(n10519), .ZN(n7678) );
  AOI21_X1 U8941 ( .B1(n7679), .B2(n9884), .A(n7678), .ZN(n10664) );
  OAI22_X1 U8942 ( .A1(n10525), .A2(n7680), .B1(n7697), .B2(n10522), .ZN(n7681) );
  AOI21_X1 U8943 ( .B1(n9677), .B2(n10661), .A(n7681), .ZN(n7683) );
  NAND2_X1 U8944 ( .A1(n10662), .A2(n9869), .ZN(n7682) );
  OAI211_X1 U8945 ( .C1(n10664), .C2(n9865), .A(n7683), .B(n7682), .ZN(n7689)
         );
  INV_X1 U8946 ( .A(n7711), .ZN(n7684) );
  NOR2_X1 U8947 ( .A1(n9418), .A2(n7684), .ZN(n9415) );
  INV_X1 U8948 ( .A(n7708), .ZN(n9442) );
  AOI21_X1 U8949 ( .B1(n7685), .B2(n9415), .A(n9442), .ZN(n7686) );
  XOR2_X1 U8950 ( .A(n7704), .B(n7686), .Z(n7687) );
  NAND2_X1 U8951 ( .A1(n7687), .A2(n9852), .ZN(n10665) );
  NOR2_X1 U8952 ( .A1(n10665), .A2(n9685), .ZN(n7688) );
  AOI211_X1 U8953 ( .C1(n9855), .C2(n10667), .A(n7689), .B(n7688), .ZN(n7690)
         );
  INV_X1 U8954 ( .A(n7690), .ZN(P1_U3284) );
  INV_X1 U8955 ( .A(n8143), .ZN(n7745) );
  INV_X1 U8956 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8144) );
  OAI222_X1 U8957 ( .A1(n9159), .A2(n7745), .B1(P2_U3151), .B2(n7691), .C1(
        n8144), .C2(n9156), .ZN(P2_U3275) );
  INV_X1 U8958 ( .A(n7692), .ZN(n7694) );
  NAND2_X1 U8959 ( .A1(n7694), .A2(n7693), .ZN(n7695) );
  XNOR2_X1 U8960 ( .A(n7696), .B(n7695), .ZN(n7703) );
  OAI22_X1 U8961 ( .A1(n9278), .A2(n7698), .B1(n9275), .B2(n7697), .ZN(n7699)
         );
  AOI211_X1 U8962 ( .C1(n8011), .C2(n9557), .A(n7700), .B(n7699), .ZN(n7702)
         );
  NAND2_X1 U8963 ( .A1(n10662), .A2(n9281), .ZN(n7701) );
  OAI211_X1 U8964 ( .C1(n7703), .C2(n9284), .A(n7702), .B(n7701), .ZN(P1_U3231) );
  NAND2_X1 U8965 ( .A1(n7705), .A2(n7704), .ZN(n7707) );
  OR2_X1 U8966 ( .A1(n10662), .A2(n10679), .ZN(n7706) );
  INV_X1 U8967 ( .A(n9557), .ZN(n7878) );
  OR2_X1 U8968 ( .A1(n10680), .A2(n7878), .ZN(n9431) );
  NAND2_X1 U8969 ( .A1(n10680), .A2(n7878), .ZN(n9427) );
  NAND2_X1 U8970 ( .A1(n9431), .A2(n9427), .ZN(n9370) );
  XNOR2_X1 U8971 ( .A(n7780), .B(n9370), .ZN(n10685) );
  INV_X1 U8972 ( .A(n10685), .ZN(n7728) );
  INV_X1 U8973 ( .A(n9370), .ZN(n7716) );
  NAND2_X1 U8974 ( .A1(n9426), .A2(n7708), .ZN(n7712) );
  NAND2_X1 U8975 ( .A1(n9416), .A2(n9410), .ZN(n7709) );
  NOR2_X1 U8976 ( .A1(n7712), .A2(n7709), .ZN(n9373) );
  NAND2_X1 U8977 ( .A1(n7710), .A2(n9373), .ZN(n7714) );
  AND2_X1 U8978 ( .A1(n9419), .A2(n7711), .ZN(n9367) );
  AND2_X1 U8979 ( .A1(n7713), .A2(n9429), .ZN(n9313) );
  NAND2_X1 U8980 ( .A1(n7714), .A2(n9313), .ZN(n7715) );
  OAI21_X1 U8981 ( .B1(n7716), .B2(n7715), .A(n7798), .ZN(n7717) );
  AOI22_X1 U8982 ( .A1(n7717), .A2(n9852), .B1(n10519), .B2(n10703), .ZN(
        n10683) );
  OAI21_X1 U8983 ( .B1(n7824), .B2(n10522), .A(n10683), .ZN(n7726) );
  INV_X1 U8984 ( .A(n10680), .ZN(n7721) );
  INV_X1 U8985 ( .A(n7719), .ZN(n7720) );
  INV_X1 U8986 ( .A(n7787), .ZN(n7788) );
  OAI211_X1 U8987 ( .C1(n7721), .C2(n7720), .A(n7788), .B(n9884), .ZN(n10681)
         );
  OAI22_X1 U8988 ( .A1(n9861), .A2(n7825), .B1(n7722), .B2(n10525), .ZN(n7723)
         );
  AOI21_X1 U8989 ( .B1(n9869), .B2(n10680), .A(n7723), .ZN(n7724) );
  OAI21_X1 U8990 ( .B1(n10681), .B2(n9865), .A(n7724), .ZN(n7725) );
  AOI21_X1 U8991 ( .B1(n7726), .B2(n10525), .A(n7725), .ZN(n7727) );
  OAI21_X1 U8992 ( .B1(n7728), .B2(n9894), .A(n7727), .ZN(P1_U3283) );
  OAI222_X1 U8993 ( .A1(n10285), .A2(n7729), .B1(P1_U3086), .B2(n9521), .C1(
        n8153), .C2(n8002), .ZN(P1_U3334) );
  INV_X1 U8994 ( .A(n10672), .ZN(n7743) );
  NAND2_X1 U8995 ( .A1(n7730), .A2(n7731), .ZN(n7732) );
  XNOR2_X1 U8996 ( .A(n10672), .B(n8552), .ZN(n7884) );
  XOR2_X1 U8997 ( .A(n8709), .B(n7884), .Z(n7734) );
  AOI21_X1 U8998 ( .B1(n7735), .B2(n7734), .A(n8683), .ZN(n7736) );
  NAND2_X1 U8999 ( .A1(n7736), .A2(n7885), .ZN(n7742) );
  AOI21_X1 U9000 ( .B1(n8710), .B2(n8676), .A(n7737), .ZN(n7738) );
  OAI21_X1 U9001 ( .B1(n7893), .B2(n8679), .A(n7738), .ZN(n7739) );
  AOI21_X1 U9002 ( .B1(n8694), .B2(n7740), .A(n7739), .ZN(n7741) );
  OAI211_X1 U9003 ( .C1(n7743), .C2(n8697), .A(n7742), .B(n7741), .ZN(P2_U3171) );
  OAI222_X1 U9004 ( .A1(n10285), .A2(n7746), .B1(n8002), .B2(n7745), .C1(n7744), .C2(P1_U3086), .ZN(P1_U3335) );
  XOR2_X1 U9005 ( .A(n7853), .B(n7861), .Z(n7749) );
  NOR2_X1 U9006 ( .A1(n6014), .A2(n7749), .ZN(n7862) );
  AOI211_X1 U9007 ( .C1(n6014), .C2(n7749), .A(n7862), .B(n9590), .ZN(n7757)
         );
  OAI21_X1 U9008 ( .B1(n7617), .B2(n7751), .A(n7750), .ZN(n7852) );
  XNOR2_X1 U9009 ( .A(n7852), .B(n7860), .ZN(n7752) );
  NAND2_X1 U9010 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n7752), .ZN(n7854) );
  OAI211_X1 U9011 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n7752), .A(n9582), .B(
        n7854), .ZN(n7755) );
  NAND2_X1 U9012 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9277) );
  INV_X1 U9013 ( .A(n9277), .ZN(n7753) );
  AOI21_X1 U9014 ( .B1(n10350), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n7753), .ZN(
        n7754) );
  OAI211_X1 U9015 ( .C1(n10360), .C2(n7860), .A(n7755), .B(n7754), .ZN(n7756)
         );
  OR2_X1 U9016 ( .A1(n7757), .A2(n7756), .ZN(P1_U3258) );
  INV_X1 U9017 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8166) );
  OAI222_X1 U9018 ( .A1(n9159), .A2(n8165), .B1(P2_U3151), .B2(n7758), .C1(
        n8166), .C2(n9156), .ZN(P2_U3273) );
  OR2_X1 U9019 ( .A1(n7761), .A2(n8187), .ZN(n7763) );
  AOI22_X1 U9020 ( .A1(n8132), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8131), .B2(
        n8745), .ZN(n7762) );
  NAND2_X1 U9021 ( .A1(n7763), .A2(n7762), .ZN(n7886) );
  XNOR2_X1 U9022 ( .A(n7886), .B(n8708), .ZN(n8318) );
  XNOR2_X1 U9023 ( .A(n7844), .B(n8318), .ZN(n10690) );
  OR2_X1 U9024 ( .A1(n10672), .A2(n8709), .ZN(n7764) );
  XOR2_X1 U9025 ( .A(n7840), .B(n8318), .Z(n7766) );
  NAND2_X1 U9026 ( .A1(n7766), .A2(n8989), .ZN(n7774) );
  NAND2_X1 U9027 ( .A1(n7587), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7772) );
  NAND2_X1 U9028 ( .A1(n8183), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7771) );
  NAND2_X1 U9029 ( .A1(n7767), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7768) );
  NAND2_X1 U9030 ( .A1(n7830), .A2(n7768), .ZN(n7996) );
  NAND2_X1 U9031 ( .A1(n8159), .A2(n7996), .ZN(n7770) );
  NAND2_X1 U9032 ( .A1(n8291), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7769) );
  NAND4_X1 U9033 ( .A1(n7772), .A2(n7771), .A3(n7770), .A4(n7769), .ZN(n8707)
         );
  AOI22_X1 U9034 ( .A1(n8994), .A2(n8709), .B1(n8707), .B2(n8995), .ZN(n7773)
         );
  OAI211_X1 U9035 ( .C1(n10690), .C2(n8256), .A(n7774), .B(n7773), .ZN(n10692)
         );
  INV_X1 U9036 ( .A(n10692), .ZN(n7779) );
  INV_X1 U9037 ( .A(n10690), .ZN(n7777) );
  INV_X1 U9038 ( .A(n7886), .ZN(n10688) );
  AOI22_X1 U9039 ( .A1(n10580), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n8983), .B2(
        n7897), .ZN(n7775) );
  OAI21_X1 U9040 ( .B1(n10688), .B2(n8937), .A(n7775), .ZN(n7776) );
  AOI21_X1 U9041 ( .B1(n7777), .B2(n8263), .A(n7776), .ZN(n7778) );
  OAI21_X1 U9042 ( .B1(n7779), .B2(n10580), .A(n7778), .ZN(P2_U3223) );
  OR2_X1 U9043 ( .A1(n10680), .A2(n9557), .ZN(n7781) );
  INV_X1 U9044 ( .A(n10703), .ZN(n7903) );
  OR2_X1 U9045 ( .A1(n7802), .A2(n7903), .ZN(n9436) );
  NAND2_X1 U9046 ( .A1(n7802), .A2(n7903), .ZN(n9439) );
  NAND2_X1 U9047 ( .A1(n9436), .A2(n9439), .ZN(n7796) );
  INV_X1 U9048 ( .A(n7796), .ZN(n9372) );
  XNOR2_X1 U9049 ( .A(n7805), .B(n9372), .ZN(n7947) );
  NAND2_X1 U9050 ( .A1(n7798), .A2(n9427), .ZN(n7782) );
  XNOR2_X1 U9051 ( .A(n7782), .B(n9372), .ZN(n7784) );
  INV_X1 U9052 ( .A(n9556), .ZN(n8008) );
  OAI22_X1 U9053 ( .A1(n7878), .A2(n10631), .B1(n8008), .B2(n9880), .ZN(n7783)
         );
  AOI21_X1 U9054 ( .B1(n7784), .B2(n9852), .A(n7783), .ZN(n7785) );
  OAI21_X1 U9055 ( .B1(n7947), .B2(n7786), .A(n7785), .ZN(n7948) );
  NAND2_X1 U9056 ( .A1(n7948), .A2(n10525), .ZN(n7793) );
  AND2_X2 U9057 ( .A1(n7787), .A2(n7955), .ZN(n7809) );
  AOI211_X1 U9058 ( .C1(n7802), .C2(n7788), .A(n9826), .B(n7809), .ZN(n7949)
         );
  NOR2_X1 U9059 ( .A1(n7955), .A2(n9888), .ZN(n7791) );
  OAI22_X1 U9060 ( .A1(n10525), .A2(n7789), .B1(n7877), .B2(n10522), .ZN(n7790) );
  AOI211_X1 U9061 ( .C1(n7949), .C2(n9891), .A(n7791), .B(n7790), .ZN(n7792)
         );
  OAI211_X1 U9062 ( .C1(n7947), .C2(n7794), .A(n7793), .B(n7792), .ZN(P1_U3282) );
  INV_X1 U9063 ( .A(n9427), .ZN(n7795) );
  NOR2_X1 U9064 ( .A1(n7796), .A2(n7795), .ZN(n7797) );
  NAND2_X1 U9065 ( .A1(n7798), .A2(n7797), .ZN(n7799) );
  NAND2_X1 U9066 ( .A1(n7799), .A2(n9436), .ZN(n7908) );
  NAND2_X1 U9067 ( .A1(n10706), .A2(n8008), .ZN(n9440) );
  NAND2_X1 U9068 ( .A1(n9453), .A2(n9440), .ZN(n7917) );
  XNOR2_X1 U9069 ( .A(n7908), .B(n7917), .ZN(n7801) );
  AND2_X1 U9070 ( .A1(n7964), .A2(n10519), .ZN(n7800) );
  AOI21_X1 U9071 ( .B1(n7801), .B2(n9852), .A(n7800), .ZN(n10709) );
  NOR2_X1 U9072 ( .A1(n7802), .A2(n10703), .ZN(n7804) );
  NAND2_X1 U9073 ( .A1(n7802), .A2(n10703), .ZN(n7803) );
  INV_X1 U9074 ( .A(n7917), .ZN(n9374) );
  XNOR2_X1 U9075 ( .A(n7918), .B(n9374), .ZN(n10712) );
  NAND2_X1 U9076 ( .A1(n10712), .A2(n9855), .ZN(n7813) );
  INV_X1 U9077 ( .A(n7902), .ZN(n7806) );
  AOI22_X1 U9078 ( .A1(n9859), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7806), .B2(
        n9857), .ZN(n7807) );
  OAI21_X1 U9079 ( .B1(n9861), .B2(n7903), .A(n7807), .ZN(n7811) );
  INV_X1 U9080 ( .A(n10706), .ZN(n7808) );
  OAI211_X1 U9081 ( .C1(n7809), .C2(n7808), .A(n9884), .B(n7919), .ZN(n10707)
         );
  NOR2_X1 U9082 ( .A1(n10707), .A2(n9865), .ZN(n7810) );
  AOI211_X1 U9083 ( .C1(n9869), .C2(n10706), .A(n7811), .B(n7810), .ZN(n7812)
         );
  OAI211_X1 U9084 ( .C1(n9685), .C2(n10709), .A(n7813), .B(n7812), .ZN(
        P1_U3281) );
  NAND2_X1 U9085 ( .A1(n8174), .A2(n10054), .ZN(n7815) );
  OR2_X1 U9086 ( .A1(n7814), .A2(P1_U3086), .ZN(n9339) );
  OAI211_X1 U9087 ( .C1(n7816), .C2(n10284), .A(n7815), .B(n9339), .ZN(
        P1_U3332) );
  NAND2_X1 U9088 ( .A1(n8174), .A2(n7817), .ZN(n7818) );
  OAI211_X1 U9089 ( .C1(n6477), .C2(n9156), .A(n7818), .B(n8507), .ZN(P2_U3272) );
  NAND2_X1 U9090 ( .A1(n7820), .A2(n7819), .ZN(n7822) );
  XNOR2_X1 U9091 ( .A(n7822), .B(n7821), .ZN(n7829) );
  OAI21_X1 U9092 ( .B1(n9276), .B2(n7903), .A(n7823), .ZN(n7827) );
  OAI22_X1 U9093 ( .A1(n9278), .A2(n7825), .B1(n9275), .B2(n7824), .ZN(n7826)
         );
  AOI211_X1 U9094 ( .C1(n10680), .C2(n9281), .A(n7827), .B(n7826), .ZN(n7828)
         );
  OAI21_X1 U9095 ( .B1(n7829), .B2(n9284), .A(n7828), .ZN(P1_U3217) );
  NAND2_X1 U9096 ( .A1(n8291), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7835) );
  NAND2_X1 U9097 ( .A1(n7587), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7834) );
  NAND2_X1 U9098 ( .A1(n7830), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7831) );
  NAND2_X1 U9099 ( .A1(n7933), .A2(n7831), .ZN(n8077) );
  NAND2_X1 U9100 ( .A1(n8159), .A2(n8077), .ZN(n7833) );
  NAND2_X1 U9101 ( .A1(n8183), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7832) );
  NAND4_X1 U9102 ( .A1(n7835), .A2(n7834), .A3(n7833), .A4(n7832), .ZN(n8706)
         );
  INV_X1 U9103 ( .A(n8706), .ZN(n8513) );
  NAND2_X1 U9104 ( .A1(n7836), .A2(n8288), .ZN(n7838) );
  AOI22_X1 U9105 ( .A1(n8132), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8131), .B2(
        n10371), .ZN(n7837) );
  NAND2_X1 U9106 ( .A1(n7838), .A2(n7837), .ZN(n7986) );
  OR2_X1 U9107 ( .A1(n7986), .A2(n8067), .ZN(n8398) );
  NAND2_X1 U9108 ( .A1(n7986), .A2(n8067), .ZN(n8387) );
  NAND2_X1 U9109 ( .A1(n8398), .A2(n8387), .ZN(n8322) );
  NAND2_X1 U9110 ( .A1(n7886), .A2(n8708), .ZN(n7839) );
  NAND2_X1 U9111 ( .A1(n7840), .A2(n7839), .ZN(n7842) );
  OR2_X1 U9112 ( .A1(n7886), .A2(n8708), .ZN(n7841) );
  XOR2_X1 U9113 ( .A(n8322), .B(n7939), .Z(n7843) );
  OAI222_X1 U9114 ( .A1(n10566), .A2(n8513), .B1(n10564), .B2(n7893), .C1(
        n10562), .C2(n7843), .ZN(n7978) );
  INV_X1 U9115 ( .A(n7978), .ZN(n7851) );
  NOR2_X1 U9116 ( .A1(n7886), .A2(n7893), .ZN(n8394) );
  INV_X1 U9117 ( .A(n8394), .ZN(n7845) );
  NAND2_X1 U9118 ( .A1(n7886), .A2(n7893), .ZN(n8381) );
  NAND2_X1 U9119 ( .A1(n7926), .A2(n8381), .ZN(n7846) );
  XOR2_X1 U9120 ( .A(n7846), .B(n8322), .Z(n7979) );
  INV_X1 U9121 ( .A(n7986), .ZN(n7999) );
  NOR2_X1 U9122 ( .A1(n7999), .A2(n8937), .ZN(n7849) );
  INV_X1 U9123 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10381) );
  INV_X1 U9124 ( .A(n7996), .ZN(n7847) );
  OAI22_X1 U9125 ( .A1(n10577), .A2(n10381), .B1(n7847), .B2(n10570), .ZN(
        n7848) );
  AOI211_X1 U9126 ( .C1(n7979), .C2(n8950), .A(n7849), .B(n7848), .ZN(n7850)
         );
  OAI21_X1 U9127 ( .B1(n7851), .B2(n10580), .A(n7850), .ZN(P2_U3222) );
  NAND2_X1 U9128 ( .A1(n7853), .A2(n7852), .ZN(n7855) );
  NAND2_X1 U9129 ( .A1(n7855), .A2(n7854), .ZN(n7859) );
  OR2_X1 U9130 ( .A1(n9564), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9572) );
  OAI21_X1 U9131 ( .B1(n7857), .B2(n7856), .A(n9572), .ZN(n7858) );
  NOR2_X1 U9132 ( .A1(n7858), .A2(n7859), .ZN(n9570) );
  AOI21_X1 U9133 ( .B1(n7859), .B2(n7858), .A(n9570), .ZN(n7872) );
  NOR2_X1 U9134 ( .A1(n7861), .A2(n7860), .ZN(n7863) );
  NAND2_X1 U9135 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9564), .ZN(n7864) );
  OAI21_X1 U9136 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9564), .A(n7864), .ZN(
        n7865) );
  NOR2_X1 U9137 ( .A1(n7866), .A2(n7865), .ZN(n9563) );
  AOI211_X1 U9138 ( .C1(n7866), .C2(n7865), .A(n9563), .B(n9590), .ZN(n7867)
         );
  INV_X1 U9139 ( .A(n7867), .ZN(n7871) );
  INV_X1 U9140 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7868) );
  NAND2_X1 U9141 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9207) );
  OAI21_X1 U9142 ( .B1(n10370), .B2(n7868), .A(n9207), .ZN(n7869) );
  AOI21_X1 U9143 ( .B1(n9564), .B2(n9609), .A(n7869), .ZN(n7870) );
  OAI211_X1 U9144 ( .C1(n7872), .C2(n10362), .A(n7871), .B(n7870), .ZN(
        P1_U3259) );
  NOR2_X1 U9145 ( .A1(n5023), .A2(n7873), .ZN(n7874) );
  XNOR2_X1 U9146 ( .A(n7875), .B(n7874), .ZN(n7876) );
  NAND2_X1 U9147 ( .A1(n7876), .A2(n9259), .ZN(n7882) );
  OAI22_X1 U9148 ( .A1(n9278), .A2(n7878), .B1(n9275), .B2(n7877), .ZN(n7879)
         );
  AOI211_X1 U9149 ( .C1(n8011), .C2(n9556), .A(n7880), .B(n7879), .ZN(n7881)
         );
  OAI211_X1 U9150 ( .C1(n7955), .C2(n9242), .A(n7882), .B(n7881), .ZN(P1_U3236) );
  INV_X1 U9151 ( .A(n7890), .ZN(n7888) );
  XOR2_X1 U9152 ( .A(n8552), .B(n7886), .Z(n7889) );
  INV_X1 U9153 ( .A(n7889), .ZN(n7887) );
  NAND2_X1 U9154 ( .A1(n7890), .A2(n7889), .ZN(n7891) );
  OAI21_X1 U9155 ( .B1(n7893), .B2(n7892), .A(n7990), .ZN(n7894) );
  NAND2_X1 U9156 ( .A1(n7894), .A2(n8685), .ZN(n7899) );
  INV_X1 U9157 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10234) );
  NOR2_X1 U9158 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10234), .ZN(n8735) );
  AOI21_X1 U9159 ( .B1(n8709), .B2(n8676), .A(n8735), .ZN(n7895) );
  OAI21_X1 U9160 ( .B1(n8067), .B2(n8679), .A(n7895), .ZN(n7896) );
  AOI21_X1 U9161 ( .B1(n8694), .B2(n7897), .A(n7896), .ZN(n7898) );
  OAI211_X1 U9162 ( .C1(n10688), .C2(n8697), .A(n7899), .B(n7898), .ZN(
        P2_U3157) );
  XOR2_X1 U9163 ( .A(n7900), .B(n7901), .Z(n7907) );
  INV_X1 U9164 ( .A(n7964), .ZN(n9167) );
  NAND2_X1 U9165 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n10367) );
  OAI21_X1 U9166 ( .B1(n9276), .B2(n9167), .A(n10367), .ZN(n7905) );
  OAI22_X1 U9167 ( .A1(n9278), .A2(n7903), .B1(n9275), .B2(n7902), .ZN(n7904)
         );
  AOI211_X1 U9168 ( .C1(n10706), .C2(n9281), .A(n7905), .B(n7904), .ZN(n7906)
         );
  OAI21_X1 U9169 ( .B1(n7907), .B2(n9284), .A(n7906), .ZN(P1_U3224) );
  NAND2_X1 U9170 ( .A1(n7908), .A2(n9374), .ZN(n7912) );
  NAND2_X1 U9171 ( .A1(n7912), .A2(n9453), .ZN(n7909) );
  NAND2_X1 U9172 ( .A1(n7958), .A2(n9167), .ZN(n9456) );
  NAND2_X1 U9173 ( .A1(n7909), .A2(n9375), .ZN(n7913) );
  INV_X1 U9174 ( .A(n9453), .ZN(n7910) );
  NOR2_X1 U9175 ( .A1(n9375), .A2(n7910), .ZN(n7911) );
  NAND2_X1 U9176 ( .A1(n7913), .A2(n7960), .ZN(n7914) );
  NAND2_X1 U9177 ( .A1(n7914), .A2(n9852), .ZN(n7916) );
  AOI22_X1 U9178 ( .A1(n10704), .A2(n9556), .B1(n9555), .B2(n10519), .ZN(n7915) );
  NAND2_X1 U9179 ( .A1(n7916), .A2(n7915), .ZN(n8026) );
  INV_X1 U9180 ( .A(n8026), .ZN(n7925) );
  XOR2_X1 U9181 ( .A(n9375), .B(n7959), .Z(n8028) );
  NAND2_X1 U9182 ( .A1(n8028), .A2(n9855), .ZN(n7924) );
  AOI211_X1 U9183 ( .C1(n7958), .C2(n7919), .A(n9826), .B(n7970), .ZN(n8027)
         );
  NOR2_X1 U9184 ( .A1(n8033), .A2(n9888), .ZN(n7922) );
  OAI22_X1 U9185 ( .A1(n10525), .A2(n7920), .B1(n8007), .B2(n10522), .ZN(n7921) );
  AOI211_X1 U9186 ( .C1(n8027), .C2(n9891), .A(n7922), .B(n7921), .ZN(n7923)
         );
  OAI211_X1 U9187 ( .C1(n9685), .C2(n7925), .A(n7924), .B(n7923), .ZN(P1_U3280) );
  AND2_X1 U9188 ( .A1(n8387), .A2(n8381), .ZN(n8395) );
  NAND2_X1 U9189 ( .A1(n7926), .A2(n8395), .ZN(n7931) );
  OR2_X1 U9190 ( .A1(n7927), .A2(n8187), .ZN(n7929) );
  AOI22_X1 U9191 ( .A1(n8132), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8131), .B2(
        n10388), .ZN(n7928) );
  XNOR2_X1 U9192 ( .A(n8401), .B(n8706), .ZN(n8400) );
  INV_X1 U9193 ( .A(n8400), .ZN(n7930) );
  NAND3_X1 U9194 ( .A1(n7931), .A2(n7930), .A3(n8398), .ZN(n7932) );
  NAND2_X1 U9195 ( .A1(n8035), .A2(n7932), .ZN(n10697) );
  NAND2_X1 U9196 ( .A1(n8291), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7938) );
  NAND2_X1 U9197 ( .A1(n7587), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7937) );
  NAND2_X1 U9198 ( .A1(n7933), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7934) );
  NAND2_X1 U9199 ( .A1(n8042), .A2(n7934), .ZN(n8648) );
  NAND2_X1 U9200 ( .A1(n8159), .A2(n8648), .ZN(n7936) );
  NAND2_X1 U9201 ( .A1(n8183), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7935) );
  NAND2_X1 U9202 ( .A1(n7986), .A2(n8707), .ZN(n7940) );
  XOR2_X1 U9203 ( .A(n8400), .B(n8050), .Z(n7941) );
  OAI222_X1 U9204 ( .A1(n10564), .A2(n8067), .B1(n10566), .B2(n8569), .C1(
        n10562), .C2(n7941), .ZN(n10699) );
  NAND2_X1 U9205 ( .A1(n10699), .A2(n10577), .ZN(n7945) );
  INV_X1 U9206 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8801) );
  INV_X1 U9207 ( .A(n8077), .ZN(n7942) );
  OAI22_X1 U9208 ( .A1(n10577), .A2(n8801), .B1(n7942), .B2(n10570), .ZN(n7943) );
  AOI21_X1 U9209 ( .B1(n8401), .B2(n9001), .A(n7943), .ZN(n7944) );
  OAI211_X1 U9210 ( .C1(n9004), .C2(n10697), .A(n7945), .B(n7944), .ZN(
        P2_U3221) );
  INV_X1 U9211 ( .A(n7946), .ZN(n10731) );
  INV_X1 U9212 ( .A(n7947), .ZN(n7950) );
  AOI211_X1 U9213 ( .C1(n10731), .C2(n7950), .A(n7949), .B(n7948), .ZN(n7952)
         );
  MUX2_X1 U9214 ( .A(n6889), .B(n7952), .S(n10736), .Z(n7951) );
  OAI21_X1 U9215 ( .B1(n7955), .B2(n9991), .A(n7951), .ZN(P1_U3533) );
  INV_X1 U9216 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7953) );
  MUX2_X1 U9217 ( .A(n7953), .B(n7952), .S(n10740), .Z(n7954) );
  OAI21_X1 U9218 ( .B1(n7955), .B2(n10040), .A(n7954), .ZN(P1_U3486) );
  INV_X1 U9219 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8189) );
  OAI222_X1 U9220 ( .A1(n9159), .A2(n8188), .B1(P2_U3151), .B2(n7956), .C1(
        n8189), .C2(n9156), .ZN(P2_U3270) );
  INV_X1 U9221 ( .A(n8177), .ZN(n8001) );
  INV_X1 U9222 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8178) );
  OAI222_X1 U9223 ( .A1(n9159), .A2(n8001), .B1(P2_U3151), .B2(n7957), .C1(
        n8178), .C2(n9156), .ZN(P2_U3271) );
  NAND2_X1 U9224 ( .A1(n9171), .A2(n9987), .ZN(n9300) );
  XNOR2_X1 U9225 ( .A(n8016), .B(n7961), .ZN(n10732) );
  NAND2_X1 U9226 ( .A1(n7960), .A2(n9456), .ZN(n7962) );
  NAND2_X1 U9227 ( .A1(n7962), .A2(n7961), .ZN(n7963) );
  NAND3_X1 U9228 ( .A1(n8014), .A2(n9852), .A3(n7963), .ZN(n7966) );
  AOI22_X1 U9229 ( .A1(n10704), .A2(n7964), .B1(n9631), .B2(n10519), .ZN(n7965) );
  NAND2_X1 U9230 ( .A1(n7966), .A2(n7965), .ZN(n7967) );
  AOI21_X1 U9231 ( .B1(n10732), .B2(n7968), .A(n7967), .ZN(n10734) );
  AOI21_X1 U9232 ( .B1(n5206), .B2(n9171), .A(n9826), .ZN(n7971) );
  NAND2_X1 U9233 ( .A1(n7971), .A2(n8019), .ZN(n10728) );
  OAI22_X1 U9234 ( .A1(n10525), .A2(n7972), .B1(n9168), .B2(n10522), .ZN(n7973) );
  AOI21_X1 U9235 ( .B1(n9171), .B2(n9869), .A(n7973), .ZN(n7974) );
  OAI21_X1 U9236 ( .B1(n10728), .B2(n9865), .A(n7974), .ZN(n7975) );
  AOI21_X1 U9237 ( .B1(n10732), .B2(n7976), .A(n7975), .ZN(n7977) );
  OAI21_X1 U9238 ( .B1(n10734), .B2(n9685), .A(n7977), .ZN(P1_U3279) );
  INV_X1 U9239 ( .A(n9141), .ZN(n9119) );
  INV_X1 U9240 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7980) );
  AOI21_X1 U9241 ( .B1(n7979), .B2(n10720), .A(n7978), .ZN(n7982) );
  MUX2_X1 U9242 ( .A(n7980), .B(n7982), .S(n10727), .Z(n7981) );
  OAI21_X1 U9243 ( .B1(n7999), .B2(n9119), .A(n7981), .ZN(P2_U3423) );
  INV_X1 U9244 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7983) );
  MUX2_X1 U9245 ( .A(n7983), .B(n7982), .S(n10723), .Z(n7984) );
  OAI21_X1 U9246 ( .B1(n7999), .B2(n9050), .A(n7984), .ZN(P2_U3470) );
  OAI222_X1 U9247 ( .A1(n6299), .A2(P1_U3086), .B1(n8002), .B2(n8188), .C1(
        n7985), .C2(n10284), .ZN(P1_U3330) );
  INV_X1 U9248 ( .A(n7990), .ZN(n7988) );
  INV_X1 U9249 ( .A(n7989), .ZN(n7987) );
  XNOR2_X1 U9250 ( .A(n7986), .B(n8552), .ZN(n8066) );
  XNOR2_X1 U9251 ( .A(n8066), .B(n8707), .ZN(n7991) );
  NOR3_X1 U9252 ( .A1(n7988), .A2(n7987), .A3(n7991), .ZN(n7993) );
  INV_X1 U9253 ( .A(n8069), .ZN(n7992) );
  OAI21_X1 U9254 ( .B1(n7993), .B2(n7992), .A(n8685), .ZN(n7998) );
  INV_X1 U9255 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10144) );
  NOR2_X1 U9256 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10144), .ZN(n10379) );
  AOI21_X1 U9257 ( .B1(n8708), .B2(n8676), .A(n10379), .ZN(n7994) );
  OAI21_X1 U9258 ( .B1(n8513), .B2(n8679), .A(n7994), .ZN(n7995) );
  AOI21_X1 U9259 ( .B1(n7996), .B2(n8694), .A(n7995), .ZN(n7997) );
  OAI211_X1 U9260 ( .C1(n7999), .C2(n8697), .A(n7998), .B(n7997), .ZN(P2_U3176) );
  OAI222_X1 U9261 ( .A1(n5603), .A2(P1_U3086), .B1(n8002), .B2(n8001), .C1(
        n8000), .C2(n10284), .ZN(P1_U3331) );
  AOI21_X1 U9262 ( .B1(n8004), .B2(n8003), .A(n9284), .ZN(n8006) );
  NAND2_X1 U9263 ( .A1(n8006), .A2(n8005), .ZN(n8013) );
  OAI22_X1 U9264 ( .A1(n9278), .A2(n8008), .B1(n9275), .B2(n8007), .ZN(n8009)
         );
  AOI211_X1 U9265 ( .C1(n8011), .C2(n9555), .A(n8010), .B(n8009), .ZN(n8012)
         );
  OAI211_X1 U9266 ( .C1(n8033), .C2(n9242), .A(n8013), .B(n8012), .ZN(P1_U3234) );
  NAND2_X1 U9267 ( .A1(n9632), .A2(n9879), .ZN(n9464) );
  NAND2_X1 U9268 ( .A1(n9468), .A2(n9464), .ZN(n9633) );
  XNOR2_X1 U9269 ( .A(n9341), .B(n9633), .ZN(n8015) );
  AOI22_X1 U9270 ( .A1(n8015), .A2(n9852), .B1(n10519), .B2(n9554), .ZN(n9986)
         );
  INV_X1 U9271 ( .A(n9633), .ZN(n9378) );
  XNOR2_X1 U9272 ( .A(n9634), .B(n9378), .ZN(n9989) );
  NAND2_X1 U9273 ( .A1(n9989), .A2(n9855), .ZN(n8025) );
  INV_X1 U9274 ( .A(n9274), .ZN(n8017) );
  AOI22_X1 U9275 ( .A1(n9859), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8017), .B2(
        n9857), .ZN(n8018) );
  OAI21_X1 U9276 ( .B1(n9861), .B2(n9987), .A(n8018), .ZN(n8023) );
  INV_X1 U9277 ( .A(n8019), .ZN(n8021) );
  INV_X1 U9278 ( .A(n9883), .ZN(n8020) );
  OAI211_X1 U9279 ( .C1(n5202), .C2(n8021), .A(n8020), .B(n9884), .ZN(n9985)
         );
  NOR2_X1 U9280 ( .A1(n9985), .A2(n9865), .ZN(n8022) );
  AOI211_X1 U9281 ( .C1(n9869), .C2(n9632), .A(n8023), .B(n8022), .ZN(n8024)
         );
  OAI211_X1 U9282 ( .C1(n9685), .C2(n9986), .A(n8025), .B(n8024), .ZN(P1_U3278) );
  INV_X1 U9283 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8029) );
  AOI211_X1 U9284 ( .C1(n8028), .C2(n10711), .A(n8027), .B(n8026), .ZN(n8031)
         );
  MUX2_X1 U9285 ( .A(n8029), .B(n8031), .S(n10740), .Z(n8030) );
  OAI21_X1 U9286 ( .B1(n8033), .B2(n10040), .A(n8030), .ZN(P1_U3492) );
  MUX2_X1 U9287 ( .A(n7164), .B(n8031), .S(n10736), .Z(n8032) );
  OAI21_X1 U9288 ( .B1(n8033), .B2(n9991), .A(n8032), .ZN(P1_U3535) );
  OR2_X1 U9289 ( .A1(n8401), .A2(n8513), .ZN(n8034) );
  OR2_X1 U9290 ( .A1(n8036), .A2(n8187), .ZN(n8038) );
  AOI22_X1 U9291 ( .A1(n8132), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8131), .B2(
        n10406), .ZN(n8037) );
  OR2_X1 U9292 ( .A1(n8652), .A2(n8569), .ZN(n8408) );
  NAND2_X1 U9293 ( .A1(n8652), .A2(n8569), .ZN(n8407) );
  NAND2_X1 U9294 ( .A1(n8039), .A2(n8288), .ZN(n8041) );
  AOI22_X1 U9295 ( .A1(n8132), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8131), .B2(
        n10423), .ZN(n8040) );
  NAND2_X1 U9296 ( .A1(n8291), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8047) );
  NAND2_X1 U9297 ( .A1(n7587), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U9298 ( .A1(n8042), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8043) );
  NAND2_X1 U9299 ( .A1(n8055), .A2(n8043), .ZN(n8572) );
  NAND2_X1 U9300 ( .A1(n8159), .A2(n8572), .ZN(n8045) );
  NAND2_X1 U9301 ( .A1(n8183), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8044) );
  NAND4_X1 U9302 ( .A1(n8047), .A2(n8046), .A3(n8045), .A4(n8044), .ZN(n8993)
         );
  XNOR2_X1 U9303 ( .A(n8514), .B(n8692), .ZN(n8326) );
  INV_X1 U9304 ( .A(n8326), .ZN(n8411) );
  OAI21_X1 U9305 ( .B1(n8048), .B2(n8411), .A(n8230), .ZN(n8092) );
  AND2_X1 U9306 ( .A1(n8401), .A2(n8706), .ZN(n8049) );
  INV_X1 U9307 ( .A(n8051), .ZN(n8082) );
  NAND2_X1 U9308 ( .A1(n8652), .A2(n8705), .ZN(n8053) );
  NAND3_X1 U9309 ( .A1(n8080), .A2(n8411), .A3(n8053), .ZN(n8054) );
  NAND3_X1 U9310 ( .A1(n8105), .A2(n8989), .A3(n8054), .ZN(n8062) );
  NAND2_X1 U9311 ( .A1(n8291), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8060) );
  NAND2_X1 U9312 ( .A1(n7587), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8059) );
  NAND2_X1 U9313 ( .A1(n8055), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8056) );
  NAND2_X1 U9314 ( .A1(n8096), .A2(n8056), .ZN(n8988) );
  NAND2_X1 U9315 ( .A1(n8159), .A2(n8988), .ZN(n8058) );
  NAND2_X1 U9316 ( .A1(n8183), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8057) );
  NAND4_X1 U9317 ( .A1(n8060), .A2(n8059), .A3(n8058), .A4(n8057), .ZN(n8978)
         );
  AOI22_X1 U9318 ( .A1(n8705), .A2(n8994), .B1(n8995), .B2(n8978), .ZN(n8061)
         );
  NAND2_X1 U9319 ( .A1(n8062), .A2(n8061), .ZN(n8091) );
  NOR2_X1 U9320 ( .A1(n8575), .A2(n10571), .ZN(n8063) );
  OAI21_X1 U9321 ( .B1(n8091), .B2(n8063), .A(n10577), .ZN(n8065) );
  AOI22_X1 U9322 ( .A1(n10580), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8983), .B2(
        n8572), .ZN(n8064) );
  OAI211_X1 U9323 ( .C1(n8092), .C2(n9004), .A(n8065), .B(n8064), .ZN(P2_U3219) );
  INV_X1 U9324 ( .A(n8401), .ZN(n10695) );
  NAND2_X1 U9325 ( .A1(n8066), .A2(n8067), .ZN(n8068) );
  NAND2_X1 U9326 ( .A1(n8069), .A2(n8068), .ZN(n8070) );
  XNOR2_X1 U9327 ( .A(n8401), .B(n8552), .ZN(n8512) );
  XOR2_X1 U9328 ( .A(n8706), .B(n8512), .Z(n8071) );
  AOI21_X1 U9329 ( .B1(n8070), .B2(n8071), .A(n8683), .ZN(n8074) );
  INV_X1 U9330 ( .A(n8070), .ZN(n8073) );
  INV_X1 U9331 ( .A(n8071), .ZN(n8072) );
  NAND2_X1 U9332 ( .A1(n8074), .A2(n8511), .ZN(n8079) );
  NOR2_X1 U9333 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10242), .ZN(n10397) );
  AOI21_X1 U9334 ( .B1(n8707), .B2(n8676), .A(n10397), .ZN(n8075) );
  OAI21_X1 U9335 ( .B1(n8569), .B2(n8679), .A(n8075), .ZN(n8076) );
  AOI21_X1 U9336 ( .B1(n8694), .B2(n8077), .A(n8076), .ZN(n8078) );
  OAI211_X1 U9337 ( .C1(n10695), .C2(n8697), .A(n8079), .B(n8078), .ZN(
        P2_U3164) );
  INV_X1 U9338 ( .A(n8652), .ZN(n10716) );
  NOR2_X1 U9339 ( .A1(n10716), .A2(n10571), .ZN(n8085) );
  OAI211_X1 U9340 ( .C1(n8082), .C2(n8081), .A(n8989), .B(n8080), .ZN(n8084)
         );
  AOI22_X1 U9341 ( .A1(n8994), .A2(n8706), .B1(n8993), .B2(n8995), .ZN(n8083)
         );
  NAND2_X1 U9342 ( .A1(n8084), .A2(n8083), .ZN(n10717) );
  AOI211_X1 U9343 ( .C1(n8983), .C2(n8648), .A(n8085), .B(n10717), .ZN(n8088)
         );
  OAI21_X1 U9344 ( .B1(n5011), .B2(n8405), .A(n8086), .ZN(n10719) );
  AOI22_X1 U9345 ( .A1(n10719), .A2(n8950), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n10580), .ZN(n8087) );
  OAI21_X1 U9346 ( .B1(n8088), .B2(n10580), .A(n8087), .ZN(P2_U3220) );
  MUX2_X1 U9347 ( .A(n8091), .B(P2_REG1_REG_14__SCAN_IN), .S(n10721), .Z(n8090) );
  OAI22_X1 U9348 ( .A1(n8092), .A2(n9064), .B1(n8575), .B2(n9050), .ZN(n8089)
         );
  OR2_X1 U9349 ( .A1(n8090), .A2(n8089), .ZN(P2_U3473) );
  MUX2_X1 U9350 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8091), .S(n10727), .Z(n8094) );
  OAI22_X1 U9351 ( .A1(n8092), .A2(n9145), .B1(n8575), .B2(n9119), .ZN(n8093)
         );
  OR2_X1 U9352 ( .A1(n8094), .A2(n8093), .ZN(P2_U3432) );
  OAI222_X1 U9353 ( .A1(n10284), .A2(n8095), .B1(n8002), .B2(n8165), .C1(n9533), .C2(P1_U3086), .ZN(P1_U3333) );
  INV_X1 U9354 ( .A(n8206), .ZN(n10281) );
  INV_X1 U9355 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8207) );
  OAI222_X1 U9356 ( .A1(n8267), .A2(n10281), .B1(n6483), .B2(P2_U3151), .C1(
        n8207), .C2(n9156), .ZN(P2_U3267) );
  NAND2_X1 U9357 ( .A1(n8291), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8101) );
  NAND2_X1 U9358 ( .A1(n7587), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8100) );
  NAND2_X1 U9359 ( .A1(n8096), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8097) );
  NAND2_X1 U9360 ( .A1(n8113), .A2(n8097), .ZN(n8982) );
  NAND2_X1 U9361 ( .A1(n8159), .A2(n8982), .ZN(n8099) );
  NAND2_X1 U9362 ( .A1(n8183), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8098) );
  NAND2_X1 U9363 ( .A1(n8102), .A2(n8288), .ZN(n8104) );
  AOI22_X1 U9364 ( .A1(n8132), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8131), .B2(
        n10457), .ZN(n8103) );
  INV_X1 U9365 ( .A(n9135), .ZN(n8109) );
  NAND2_X1 U9366 ( .A1(n8514), .A2(n8993), .ZN(n8418) );
  OR2_X1 U9367 ( .A1(n8106), .A2(n8187), .ZN(n8108) );
  AOI22_X1 U9368 ( .A1(n8132), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8131), .B2(
        n10440), .ZN(n8107) );
  INV_X1 U9369 ( .A(n8978), .ZN(n8610) );
  NAND2_X1 U9370 ( .A1(n9142), .A2(n8610), .ZN(n8420) );
  NAND2_X1 U9371 ( .A1(n8421), .A2(n8420), .ZN(n8991) );
  INV_X1 U9372 ( .A(n9142), .ZN(n8698) );
  XNOR2_X1 U9373 ( .A(n9135), .B(n8619), .ZN(n8976) );
  NAND2_X1 U9374 ( .A1(n8977), .A2(n8976), .ZN(n8975) );
  NAND2_X1 U9375 ( .A1(n8110), .A2(n8288), .ZN(n8112) );
  INV_X1 U9376 ( .A(n8819), .ZN(n10475) );
  AOI22_X1 U9377 ( .A1(n8132), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8131), .B2(
        n10475), .ZN(n8111) );
  NAND2_X1 U9378 ( .A1(n7587), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8118) );
  NAND2_X1 U9379 ( .A1(n8291), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8117) );
  NAND2_X1 U9380 ( .A1(n8113), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8114) );
  NAND2_X1 U9381 ( .A1(n8122), .A2(n8114), .ZN(n8970) );
  NAND2_X1 U9382 ( .A1(n8159), .A2(n8970), .ZN(n8116) );
  NAND2_X1 U9383 ( .A1(n8183), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8115) );
  XNOR2_X1 U9384 ( .A(n9129), .B(n8668), .ZN(n8965) );
  INV_X1 U9385 ( .A(n9129), .ZN(n8430) );
  OR2_X1 U9386 ( .A1(n8119), .A2(n8187), .ZN(n8121) );
  AOI22_X1 U9387 ( .A1(n8132), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8131), .B2(
        n10510), .ZN(n8120) );
  INV_X1 U9388 ( .A(n9123), .ZN(n8672) );
  NAND2_X1 U9389 ( .A1(n8291), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8127) );
  NAND2_X1 U9390 ( .A1(n7587), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8126) );
  NAND2_X1 U9391 ( .A1(n8122), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8123) );
  NAND2_X1 U9392 ( .A1(n8135), .A2(n8123), .ZN(n8959) );
  NAND2_X1 U9393 ( .A1(n8159), .A2(n8959), .ZN(n8125) );
  NAND2_X1 U9394 ( .A1(n8160), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8124) );
  NAND4_X1 U9395 ( .A1(n8127), .A2(n8126), .A3(n8125), .A4(n8124), .ZN(n8967)
         );
  NAND2_X1 U9396 ( .A1(n8672), .A2(n8945), .ZN(n8129) );
  NAND2_X1 U9397 ( .A1(n8130), .A2(n8288), .ZN(n8134) );
  AOI22_X1 U9398 ( .A1(n8132), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8833), .B2(
        n8131), .ZN(n8133) );
  NAND2_X1 U9399 ( .A1(n8291), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8140) );
  NAND2_X1 U9400 ( .A1(n7587), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8139) );
  NAND2_X1 U9401 ( .A1(n8135), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8136) );
  NAND2_X1 U9402 ( .A1(n8147), .A2(n8136), .ZN(n8946) );
  NAND2_X1 U9403 ( .A1(n8159), .A2(n8946), .ZN(n8138) );
  NAND2_X1 U9404 ( .A1(n8183), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8137) );
  NAND4_X1 U9405 ( .A1(n8140), .A2(n8139), .A3(n8138), .A4(n8137), .ZN(n8957)
         );
  INV_X1 U9406 ( .A(n8957), .ZN(n8931) );
  NAND2_X1 U9407 ( .A1(n8143), .A2(n8288), .ZN(n8146) );
  OR2_X1 U9408 ( .A1(n8208), .A2(n8144), .ZN(n8145) );
  NAND2_X1 U9409 ( .A1(n8291), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8152) );
  NAND2_X1 U9410 ( .A1(n7587), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8151) );
  NAND2_X1 U9411 ( .A1(n8147), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8148) );
  NAND2_X1 U9412 ( .A1(n8157), .A2(n8148), .ZN(n8935) );
  NAND2_X1 U9413 ( .A1(n8159), .A2(n8935), .ZN(n8150) );
  NAND2_X1 U9414 ( .A1(n8160), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8149) );
  NAND4_X1 U9415 ( .A1(n8152), .A2(n8151), .A3(n8150), .A4(n8149), .ZN(n8704)
         );
  XNOR2_X1 U9416 ( .A(n8642), .B(n8944), .ZN(n8934) );
  OR2_X1 U9417 ( .A1(n8153), .A2(n8187), .ZN(n8156) );
  OR2_X1 U9418 ( .A1(n8208), .A2(n8154), .ZN(n8155) );
  NAND2_X1 U9419 ( .A1(n8157), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8158) );
  NAND2_X1 U9420 ( .A1(n8169), .A2(n8158), .ZN(n8923) );
  NAND2_X1 U9421 ( .A1(n8923), .A2(n8159), .ZN(n8164) );
  NAND2_X1 U9422 ( .A1(n7587), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8163) );
  NAND2_X1 U9423 ( .A1(n8291), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8162) );
  NAND2_X1 U9424 ( .A1(n8160), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8161) );
  NAND4_X1 U9425 ( .A1(n8164), .A2(n8163), .A3(n8162), .A4(n8161), .ZN(n8703)
         );
  NAND2_X1 U9426 ( .A1(n8922), .A2(n8703), .ZN(n8448) );
  NAND2_X1 U9427 ( .A1(n8451), .A2(n8448), .ZN(n8309) );
  OR2_X1 U9428 ( .A1(n8208), .A2(n8166), .ZN(n8167) );
  INV_X1 U9429 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9105) );
  NAND2_X1 U9430 ( .A1(n8169), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8170) );
  NAND2_X1 U9431 ( .A1(n8171), .A2(n8170), .ZN(n8910) );
  NAND2_X1 U9432 ( .A1(n8910), .A2(n8159), .ZN(n8173) );
  AOI22_X1 U9433 ( .A1(n8291), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n7587), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n8172) );
  NOR2_X1 U9434 ( .A1(n9035), .A2(n8702), .ZN(n8308) );
  NAND2_X1 U9435 ( .A1(n8174), .A2(n8288), .ZN(n8176) );
  OR2_X1 U9436 ( .A1(n8208), .A2(n6477), .ZN(n8175) );
  INV_X1 U9437 ( .A(n8902), .ZN(n9100) );
  NAND2_X1 U9438 ( .A1(n8177), .A2(n8288), .ZN(n8180) );
  OR2_X1 U9439 ( .A1(n8208), .A2(n8178), .ZN(n8179) );
  NAND2_X1 U9440 ( .A1(n8181), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8182) );
  NAND2_X1 U9441 ( .A1(n8192), .A2(n8182), .ZN(n8889) );
  NAND2_X1 U9442 ( .A1(n8889), .A2(n8159), .ZN(n8186) );
  AOI22_X1 U9443 ( .A1(n8291), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n6990), .B2(
        P2_REG1_REG_24__SCAN_IN), .ZN(n8185) );
  NAND2_X1 U9444 ( .A1(n8183), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8184) );
  NAND2_X1 U9445 ( .A1(n8632), .A2(n8898), .ZN(n8465) );
  NAND2_X1 U9446 ( .A1(n8464), .A2(n8465), .ZN(n8459) );
  INV_X1 U9447 ( .A(n8632), .ZN(n9095) );
  INV_X1 U9448 ( .A(n9026), .ZN(n8880) );
  NAND2_X1 U9449 ( .A1(n8192), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8193) );
  NAND2_X1 U9450 ( .A1(n8194), .A2(n8193), .ZN(n8882) );
  NAND2_X1 U9451 ( .A1(n8882), .A2(n8159), .ZN(n8199) );
  INV_X1 U9452 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9091) );
  NAND2_X1 U9453 ( .A1(n7587), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8196) );
  NAND2_X1 U9454 ( .A1(n8291), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8195) );
  OAI211_X1 U9455 ( .C1(n8215), .C2(n9091), .A(n8196), .B(n8195), .ZN(n8197)
         );
  INV_X1 U9456 ( .A(n8197), .ZN(n8198) );
  NAND2_X1 U9457 ( .A1(n8880), .A2(n8887), .ZN(n8200) );
  AOI22_X1 U9458 ( .A1(n8877), .A2(n8200), .B1(n9026), .B2(n8700), .ZN(n8866)
         );
  NAND2_X1 U9459 ( .A1(n9157), .A2(n8288), .ZN(n8202) );
  INV_X1 U9460 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9160) );
  NAND2_X1 U9461 ( .A1(n9086), .A2(n8859), .ZN(n8203) );
  INV_X1 U9462 ( .A(n9086), .ZN(n9022) );
  NAND2_X1 U9463 ( .A1(n8265), .A2(n8288), .ZN(n8205) );
  INV_X1 U9464 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8266) );
  NAND2_X1 U9465 ( .A1(n9080), .A2(n8869), .ZN(n8476) );
  NAND2_X1 U9466 ( .A1(n8206), .A2(n8288), .ZN(n8210) );
  NAND2_X1 U9467 ( .A1(n8211), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8212) );
  NAND2_X1 U9468 ( .A1(n8260), .A2(n8212), .ZN(n8851) );
  NAND2_X1 U9469 ( .A1(n8851), .A2(n8159), .ZN(n8218) );
  INV_X1 U9470 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9073) );
  NAND2_X1 U9471 ( .A1(n8291), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8214) );
  NAND2_X1 U9472 ( .A1(n7587), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8213) );
  OAI211_X1 U9473 ( .C1(n9073), .C2(n8215), .A(n8214), .B(n8213), .ZN(n8216)
         );
  INV_X1 U9474 ( .A(n8216), .ZN(n8217) );
  NOR2_X1 U9475 ( .A1(n9074), .A2(n8858), .ZN(n8219) );
  INV_X1 U9476 ( .A(n9074), .ZN(n9015) );
  NAND2_X1 U9477 ( .A1(n8221), .A2(n8220), .ZN(n8225) );
  INV_X1 U9478 ( .A(n8222), .ZN(n8223) );
  NAND2_X1 U9479 ( .A1(n8223), .A2(n10062), .ZN(n8224) );
  MUX2_X1 U9480 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n8278), .Z(n8269) );
  INV_X1 U9481 ( .A(SI_29_), .ZN(n8226) );
  NAND2_X1 U9482 ( .A1(n9289), .A2(n8288), .ZN(n8228) );
  OR2_X1 U9483 ( .A1(n8208), .A2(n9155), .ZN(n8227) );
  NAND2_X1 U9484 ( .A1(n8228), .A2(n8227), .ZN(n8259) );
  NAND2_X1 U9485 ( .A1(n8259), .A2(n8846), .ZN(n8478) );
  OR2_X1 U9486 ( .A1(n8514), .A2(n8692), .ZN(n8229) );
  NAND2_X1 U9487 ( .A1(n8230), .A2(n8229), .ZN(n8987) );
  INV_X1 U9488 ( .A(n8965), .ZN(n8963) );
  NAND2_X1 U9489 ( .A1(n9123), .A2(n8945), .ZN(n8429) );
  NAND2_X1 U9490 ( .A1(n8232), .A2(n8434), .ZN(n8948) );
  XNOR2_X1 U9491 ( .A(n8947), .B(n8957), .ZN(n8941) );
  OR2_X1 U9492 ( .A1(n8947), .A2(n8931), .ZN(n8233) );
  INV_X1 U9493 ( .A(n8934), .ZN(n8928) );
  INV_X1 U9494 ( .A(n8703), .ZN(n8932) );
  OR2_X1 U9495 ( .A1(n8922), .A2(n8932), .ZN(n8234) );
  INV_X1 U9496 ( .A(n8702), .ZN(n8919) );
  NOR2_X1 U9497 ( .A1(n9035), .A2(n8919), .ZN(n8455) );
  NAND2_X1 U9498 ( .A1(n9035), .A2(n8919), .ZN(n8453) );
  OR2_X1 U9499 ( .A1(n8902), .A2(n8907), .ZN(n8460) );
  NAND2_X1 U9500 ( .A1(n8902), .A2(n8907), .ZN(n8461) );
  NOR2_X1 U9501 ( .A1(n9026), .A2(n8887), .ZN(n8468) );
  NAND2_X1 U9502 ( .A1(n9026), .A2(n8887), .ZN(n8307) );
  NAND2_X1 U9503 ( .A1(n9086), .A2(n8879), .ZN(n8470) );
  NAND2_X1 U9504 ( .A1(n8235), .A2(n8470), .ZN(n8855) );
  INV_X1 U9505 ( .A(n8476), .ZN(n8236) );
  OR2_X1 U9506 ( .A1(n8855), .A2(n8236), .ZN(n8239) );
  AND2_X1 U9507 ( .A1(n8299), .A2(n8475), .ZN(n8238) );
  NAND2_X1 U9508 ( .A1(n9074), .A2(n8237), .ZN(n8242) );
  INV_X1 U9509 ( .A(n8242), .ZN(n8300) );
  AOI21_X1 U9510 ( .B1(n8239), .B2(n8238), .A(n8300), .ZN(n8248) );
  NAND2_X1 U9511 ( .A1(n8476), .A2(n8470), .ZN(n8240) );
  NAND3_X1 U9512 ( .A1(n8298), .A2(n8247), .A3(n8844), .ZN(n8245) );
  NAND2_X1 U9513 ( .A1(n8475), .A2(n8471), .ZN(n8241) );
  AND2_X1 U9514 ( .A1(n8241), .A2(n8476), .ZN(n8297) );
  NAND2_X1 U9515 ( .A1(n8297), .A2(n8242), .ZN(n8243) );
  OAI21_X2 U9516 ( .B1(n8248), .B2(n8247), .A(n8246), .ZN(n8258) );
  AND2_X1 U9517 ( .A1(n8249), .A2(P2_B_REG_SCAN_IN), .ZN(n8250) );
  NOR2_X1 U9518 ( .A1(n10566), .A2(n8250), .ZN(n8835) );
  NAND2_X1 U9519 ( .A1(n8183), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8253) );
  NAND2_X1 U9520 ( .A1(n8291), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8252) );
  NAND2_X1 U9521 ( .A1(n7587), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8251) );
  AND3_X1 U9522 ( .A1(n8253), .A2(n8252), .A3(n8251), .ZN(n8254) );
  NAND2_X1 U9523 ( .A1(n8296), .A2(n8254), .ZN(n8699) );
  AOI22_X1 U9524 ( .A1(n8858), .A2(n8994), .B1(n8835), .B2(n8699), .ZN(n8255)
         );
  OAI21_X1 U9525 ( .B1(n8258), .B2(n8256), .A(n8255), .ZN(n8257) );
  INV_X1 U9526 ( .A(n8258), .ZN(n9009) );
  INV_X1 U9527 ( .A(n8259), .ZN(n9010) );
  NOR2_X1 U9528 ( .A1(n8260), .A2(n10570), .ZN(n8837) );
  AOI21_X1 U9529 ( .B1(n10580), .B2(P2_REG2_REG_29__SCAN_IN), .A(n8837), .ZN(
        n8261) );
  OAI21_X1 U9530 ( .B1(n9010), .B2(n8937), .A(n8261), .ZN(n8262) );
  AOI21_X1 U9531 ( .B1(n9009), .B2(n8263), .A(n8262), .ZN(n8264) );
  OAI21_X1 U9532 ( .B1(n9013), .B2(n10580), .A(n8264), .ZN(P2_U3204) );
  INV_X1 U9533 ( .A(n8265), .ZN(n10283) );
  OAI222_X1 U9534 ( .A1(n8267), .A2(n10283), .B1(n8825), .B2(P2_U3151), .C1(
        n8266), .C2(n9156), .ZN(P2_U3268) );
  NAND2_X1 U9535 ( .A1(n8268), .A2(SI_29_), .ZN(n8273) );
  INV_X1 U9536 ( .A(n8269), .ZN(n8270) );
  NAND2_X1 U9537 ( .A1(n8273), .A2(n8272), .ZN(n8285) );
  INV_X1 U9538 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9295) );
  MUX2_X1 U9539 ( .A(n9295), .B(n8509), .S(n8278), .Z(n8274) );
  INV_X1 U9540 ( .A(SI_30_), .ZN(n10166) );
  NAND2_X1 U9541 ( .A1(n8274), .A2(n10166), .ZN(n8277) );
  INV_X1 U9542 ( .A(n8274), .ZN(n8275) );
  NAND2_X1 U9543 ( .A1(n8275), .A2(SI_30_), .ZN(n8276) );
  NAND2_X1 U9544 ( .A1(n8277), .A2(n8276), .ZN(n8284) );
  MUX2_X1 U9545 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8278), .Z(n8280) );
  INV_X1 U9546 ( .A(SI_31_), .ZN(n8279) );
  XNOR2_X1 U9547 ( .A(n8280), .B(n8279), .ZN(n8281) );
  NOR2_X1 U9548 ( .A1(n8208), .A2(n6453), .ZN(n8283) );
  NAND2_X1 U9549 ( .A1(n8285), .A2(n8284), .ZN(n8286) );
  NAND2_X1 U9550 ( .A1(n10055), .A2(n8288), .ZN(n8290) );
  OR2_X1 U9551 ( .A1(n8208), .A2(n8509), .ZN(n8289) );
  NAND2_X1 U9552 ( .A1(n8183), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8294) );
  NAND2_X1 U9553 ( .A1(n8291), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8293) );
  NAND2_X1 U9554 ( .A1(n7587), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8292) );
  AND3_X1 U9555 ( .A1(n8294), .A2(n8293), .A3(n8292), .ZN(n8295) );
  NAND2_X1 U9556 ( .A1(n8296), .A2(n8295), .ZN(n8836) );
  AND2_X1 U9557 ( .A1(n9067), .A2(n8836), .ZN(n8496) );
  INV_X1 U9558 ( .A(n8699), .ZN(n8301) );
  NAND2_X1 U9559 ( .A1(n9070), .A2(n8699), .ZN(n8306) );
  AOI21_X1 U9560 ( .B1(n8836), .B2(n8306), .A(n9067), .ZN(n8304) );
  NOR2_X1 U9561 ( .A1(n8305), .A2(n8304), .ZN(n8335) );
  OAI21_X1 U9562 ( .B1(n9067), .B2(n8836), .A(n8306), .ZN(n8488) );
  INV_X1 U9563 ( .A(n8307), .ZN(n8467) );
  NAND2_X1 U9564 ( .A1(n8471), .A2(n8470), .ZN(n8867) );
  INV_X1 U9565 ( .A(n8309), .ZN(n8921) );
  INV_X1 U9566 ( .A(n8941), .ZN(n8949) );
  NAND3_X1 U9567 ( .A1(n8311), .A2(n8310), .A3(n8356), .ZN(n8317) );
  NAND4_X1 U9568 ( .A1(n10557), .A2(n8314), .A3(n8313), .A4(n8312), .ZN(n8316)
         );
  NOR3_X1 U9569 ( .A1(n8317), .A2(n8316), .A3(n8315), .ZN(n8321) );
  NAND4_X1 U9570 ( .A1(n8321), .A2(n8320), .A3(n8319), .A4(n8318), .ZN(n8323)
         );
  NOR2_X1 U9571 ( .A1(n8323), .A2(n8322), .ZN(n8324) );
  NAND3_X1 U9572 ( .A1(n8405), .A2(n8324), .A3(n8400), .ZN(n8325) );
  NOR3_X1 U9573 ( .A1(n8991), .A2(n8326), .A3(n8325), .ZN(n8327) );
  NAND4_X1 U9574 ( .A1(n8955), .A2(n8327), .A3(n8973), .A4(n8963), .ZN(n8328)
         );
  NOR3_X1 U9575 ( .A1(n8921), .A2(n8949), .A3(n8328), .ZN(n8329) );
  NAND4_X1 U9576 ( .A1(n8908), .A2(n8458), .A3(n8329), .A4(n8928), .ZN(n8330)
         );
  NAND4_X1 U9577 ( .A1(n8490), .A2(n8856), .A3(n8844), .A4(n8331), .ZN(n8332)
         );
  NOR4_X1 U9578 ( .A1(n8488), .A2(n8496), .A3(n8480), .A4(n8332), .ZN(n8333)
         );
  NOR2_X1 U9579 ( .A1(n8339), .A2(n8338), .ZN(n8340) );
  NOR2_X1 U9580 ( .A1(n8337), .A2(n8340), .ZN(n8348) );
  INV_X1 U9581 ( .A(n8341), .ZN(n8343) );
  OAI211_X1 U9582 ( .C1(n8345), .C2(n8344), .A(n8343), .B(n8342), .ZN(n8347)
         );
  NAND2_X1 U9583 ( .A1(n8350), .A2(n8349), .ZN(n8353) );
  NAND2_X1 U9584 ( .A1(n8357), .A2(n8351), .ZN(n8352) );
  MUX2_X1 U9585 ( .A(n8353), .B(n8352), .S(n8492), .Z(n8354) );
  INV_X1 U9586 ( .A(n8354), .ZN(n8355) );
  INV_X1 U9587 ( .A(n8357), .ZN(n8359) );
  OAI211_X1 U9588 ( .C1(n8364), .C2(n8359), .A(n8365), .B(n8358), .ZN(n8360)
         );
  NAND3_X1 U9589 ( .A1(n8360), .A2(n8361), .A3(n8369), .ZN(n8368) );
  OAI211_X1 U9590 ( .C1(n8364), .C2(n8363), .A(n8362), .B(n8361), .ZN(n8366)
         );
  NAND3_X1 U9591 ( .A1(n8366), .A2(n8365), .A3(n8370), .ZN(n8367) );
  MUX2_X1 U9592 ( .A(n8368), .B(n8367), .S(n8492), .Z(n8374) );
  MUX2_X1 U9593 ( .A(n8370), .B(n8369), .S(n8492), .Z(n8372) );
  AND2_X1 U9594 ( .A1(n8372), .A2(n8371), .ZN(n8373) );
  NAND2_X1 U9595 ( .A1(n8374), .A2(n8373), .ZN(n8391) );
  NAND2_X1 U9596 ( .A1(n8392), .A2(n8375), .ZN(n8377) );
  NAND2_X1 U9597 ( .A1(n8380), .A2(n8379), .ZN(n8376) );
  MUX2_X1 U9598 ( .A(n8377), .B(n8376), .S(n8491), .Z(n8389) );
  INV_X1 U9599 ( .A(n8389), .ZN(n8384) );
  NAND2_X1 U9600 ( .A1(n8379), .A2(n8378), .ZN(n8383) );
  NAND2_X1 U9601 ( .A1(n8381), .A2(n8380), .ZN(n8382) );
  AOI21_X1 U9602 ( .B1(n8384), .B2(n8383), .A(n8382), .ZN(n8385) );
  OAI21_X1 U9603 ( .B1(n8391), .B2(n8389), .A(n8385), .ZN(n8386) );
  NAND3_X1 U9604 ( .A1(n8386), .A2(n8398), .A3(n7845), .ZN(n8388) );
  NAND2_X1 U9605 ( .A1(n8388), .A2(n8387), .ZN(n8399) );
  AOI21_X1 U9606 ( .B1(n8391), .B2(n8390), .A(n8389), .ZN(n8397) );
  INV_X1 U9607 ( .A(n8392), .ZN(n8393) );
  OR2_X1 U9608 ( .A1(n8394), .A2(n8393), .ZN(n8396) );
  NAND2_X1 U9609 ( .A1(n8706), .A2(n8491), .ZN(n8403) );
  NAND2_X1 U9610 ( .A1(n8513), .A2(n8492), .ZN(n8402) );
  MUX2_X1 U9611 ( .A(n8403), .B(n8402), .S(n8401), .Z(n8404) );
  NAND3_X1 U9612 ( .A1(n8406), .A2(n8405), .A3(n8404), .ZN(n8410) );
  MUX2_X1 U9613 ( .A(n8408), .B(n8407), .S(n8491), .Z(n8409) );
  NAND2_X1 U9614 ( .A1(n8410), .A2(n8409), .ZN(n8417) );
  NAND2_X1 U9615 ( .A1(n8417), .A2(n8411), .ZN(n8416) );
  NAND2_X1 U9616 ( .A1(n8421), .A2(n8692), .ZN(n8413) );
  NAND2_X1 U9617 ( .A1(n8420), .A2(n8575), .ZN(n8412) );
  MUX2_X1 U9618 ( .A(n8413), .B(n8412), .S(n8491), .Z(n8414) );
  INV_X1 U9619 ( .A(n8414), .ZN(n8415) );
  INV_X1 U9620 ( .A(n8417), .ZN(n8419) );
  MUX2_X1 U9621 ( .A(n8421), .B(n8420), .S(n8492), .Z(n8422) );
  OR2_X1 U9622 ( .A1(n9135), .A2(n8491), .ZN(n8424) );
  NAND2_X1 U9623 ( .A1(n9135), .A2(n8491), .ZN(n8423) );
  MUX2_X1 U9624 ( .A(n8424), .B(n8423), .S(n8619), .Z(n8425) );
  INV_X1 U9625 ( .A(n8668), .ZN(n8979) );
  MUX2_X1 U9626 ( .A(n8979), .B(n9129), .S(n8491), .Z(n8426) );
  NAND3_X1 U9627 ( .A1(n8431), .A2(n8668), .A3(n8434), .ZN(n8428) );
  NAND3_X1 U9628 ( .A1(n8432), .A2(n8955), .A3(n9129), .ZN(n8427) );
  NAND3_X1 U9629 ( .A1(n8428), .A2(n8429), .A3(n8427), .ZN(n8437) );
  NAND3_X1 U9630 ( .A1(n8431), .A2(n8430), .A3(n8429), .ZN(n8435) );
  NAND3_X1 U9631 ( .A1(n8432), .A2(n8955), .A3(n8979), .ZN(n8433) );
  NAND3_X1 U9632 ( .A1(n8435), .A2(n8434), .A3(n8433), .ZN(n8436) );
  MUX2_X1 U9633 ( .A(n8437), .B(n8436), .S(n8492), .Z(n8442) );
  AND2_X1 U9634 ( .A1(n8957), .A2(n8491), .ZN(n8439) );
  NOR2_X1 U9635 ( .A1(n8957), .A2(n8491), .ZN(n8438) );
  MUX2_X1 U9636 ( .A(n8439), .B(n8438), .S(n8947), .Z(n8440) );
  NOR2_X1 U9637 ( .A1(n8934), .A2(n8440), .ZN(n8441) );
  OAI21_X1 U9638 ( .B1(n8442), .B2(n8949), .A(n8441), .ZN(n8446) );
  OR2_X1 U9639 ( .A1(n8642), .A2(n8491), .ZN(n8444) );
  NAND2_X1 U9640 ( .A1(n8642), .A2(n8491), .ZN(n8443) );
  MUX2_X1 U9641 ( .A(n8444), .B(n8443), .S(n8944), .Z(n8445) );
  NAND2_X1 U9642 ( .A1(n8446), .A2(n8445), .ZN(n8452) );
  INV_X1 U9643 ( .A(n8452), .ZN(n8449) );
  MUX2_X1 U9644 ( .A(n8703), .B(n8922), .S(n8492), .Z(n8447) );
  OAI21_X1 U9645 ( .B1(n8449), .B2(n8448), .A(n8447), .ZN(n8450) );
  OAI21_X1 U9646 ( .B1(n8452), .B2(n8451), .A(n8450), .ZN(n8457) );
  INV_X1 U9647 ( .A(n8453), .ZN(n8454) );
  MUX2_X1 U9648 ( .A(n8455), .B(n8454), .S(n8492), .Z(n8456) );
  AOI21_X1 U9649 ( .B1(n8457), .B2(n8908), .A(n8456), .ZN(n8463) );
  INV_X1 U9650 ( .A(n8459), .ZN(n8890) );
  MUX2_X1 U9651 ( .A(n8461), .B(n8460), .S(n8491), .Z(n8462) );
  MUX2_X1 U9652 ( .A(n8465), .B(n8464), .S(n8492), .Z(n8466) );
  MUX2_X1 U9653 ( .A(n8468), .B(n8467), .S(n8492), .Z(n8469) );
  INV_X1 U9654 ( .A(n8470), .ZN(n8473) );
  INV_X1 U9655 ( .A(n8471), .ZN(n8472) );
  MUX2_X1 U9656 ( .A(n8473), .B(n8472), .S(n8492), .Z(n8474) );
  MUX2_X1 U9657 ( .A(n8476), .B(n8475), .S(n8492), .Z(n8477) );
  MUX2_X1 U9658 ( .A(n8858), .B(n9074), .S(n8491), .Z(n8482) );
  AND3_X1 U9659 ( .A1(n8490), .A2(n8491), .A3(n8478), .ZN(n8487) );
  AOI22_X1 U9660 ( .A1(n8487), .A2(n8858), .B1(n8492), .B2(n9074), .ZN(n8479)
         );
  AOI21_X1 U9661 ( .B1(n8481), .B2(n8482), .A(n8479), .ZN(n8486) );
  INV_X1 U9662 ( .A(n8481), .ZN(n8484) );
  INV_X1 U9663 ( .A(n8482), .ZN(n8483) );
  INV_X1 U9664 ( .A(n8488), .ZN(n8489) );
  INV_X1 U9665 ( .A(n8496), .ZN(n8497) );
  OAI21_X1 U9666 ( .B1(n8499), .B2(n8498), .A(n8497), .ZN(n8500) );
  NAND3_X1 U9667 ( .A1(n8503), .A2(n8502), .A3(n8825), .ZN(n8504) );
  OAI211_X1 U9668 ( .C1(n8505), .C2(n8507), .A(n8504), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8506) );
  INV_X1 U9669 ( .A(n10055), .ZN(n8510) );
  OAI222_X1 U9670 ( .A1(n8508), .A2(P2_U3151), .B1(n9159), .B2(n8510), .C1(
        n9156), .C2(n8509), .ZN(P2_U3265) );
  XNOR2_X1 U9671 ( .A(n8652), .B(n8552), .ZN(n8645) );
  XNOR2_X1 U9672 ( .A(n8514), .B(n8552), .ZN(n8515) );
  XNOR2_X1 U9673 ( .A(n8515), .B(n8993), .ZN(n8566) );
  AND2_X1 U9674 ( .A1(n8515), .A2(n8692), .ZN(n8516) );
  XNOR2_X1 U9675 ( .A(n9142), .B(n8552), .ZN(n8517) );
  XNOR2_X1 U9676 ( .A(n8517), .B(n8978), .ZN(n8687) );
  INV_X1 U9677 ( .A(n8517), .ZN(n8518) );
  NAND2_X1 U9678 ( .A1(n8518), .A2(n8978), .ZN(n8519) );
  NAND2_X1 U9679 ( .A1(n8686), .A2(n8519), .ZN(n8604) );
  XNOR2_X1 U9680 ( .A(n9135), .B(n8552), .ZN(n8605) );
  NAND2_X1 U9681 ( .A1(n8605), .A2(n8619), .ZN(n8520) );
  NAND2_X1 U9682 ( .A1(n8604), .A2(n8520), .ZN(n8523) );
  INV_X1 U9683 ( .A(n8605), .ZN(n8521) );
  NAND2_X1 U9684 ( .A1(n8521), .A2(n8996), .ZN(n8522) );
  XNOR2_X1 U9685 ( .A(n9129), .B(n8552), .ZN(n8615) );
  NAND2_X1 U9686 ( .A1(n8615), .A2(n8668), .ZN(n8524) );
  XNOR2_X1 U9687 ( .A(n9123), .B(n8552), .ZN(n8525) );
  XOR2_X1 U9688 ( .A(n8967), .B(n8525), .Z(n8663) );
  INV_X1 U9689 ( .A(n8525), .ZN(n8526) );
  XNOR2_X1 U9690 ( .A(n8941), .B(n8552), .ZN(n8583) );
  NAND2_X1 U9691 ( .A1(n8584), .A2(n8583), .ZN(n8582) );
  INV_X1 U9692 ( .A(n8583), .ZN(n8527) );
  NAND2_X1 U9693 ( .A1(n8527), .A2(n8957), .ZN(n8528) );
  NAND2_X1 U9694 ( .A1(n8582), .A2(n8528), .ZN(n8637) );
  INV_X1 U9695 ( .A(n8637), .ZN(n8530) );
  XNOR2_X1 U9696 ( .A(n8642), .B(n8552), .ZN(n8531) );
  XOR2_X1 U9697 ( .A(n8704), .B(n8531), .Z(n8638) );
  NAND2_X1 U9698 ( .A1(n8531), .A2(n8944), .ZN(n8532) );
  NAND2_X1 U9699 ( .A1(n8635), .A2(n8532), .ZN(n8589) );
  XNOR2_X1 U9700 ( .A(n8922), .B(n8552), .ZN(n8533) );
  XNOR2_X1 U9701 ( .A(n9035), .B(n8552), .ZN(n8536) );
  XOR2_X1 U9702 ( .A(n8702), .B(n8536), .Z(n8655) );
  INV_X1 U9703 ( .A(n8536), .ZN(n8537) );
  NAND2_X1 U9704 ( .A1(n8537), .A2(n8702), .ZN(n8538) );
  XNOR2_X1 U9705 ( .A(n8632), .B(n6861), .ZN(n8626) );
  XNOR2_X1 U9706 ( .A(n8902), .B(n6861), .ZN(n8539) );
  OAI22_X1 U9707 ( .A1(n8626), .A2(n8898), .B1(n8907), .B2(n8539), .ZN(n8543)
         );
  INV_X1 U9708 ( .A(n8898), .ZN(n8701) );
  OAI21_X1 U9709 ( .B1(n8623), .B2(n8624), .A(n8701), .ZN(n8541) );
  NOR2_X1 U9710 ( .A1(n8701), .A2(n8624), .ZN(n8540) );
  AOI22_X1 U9711 ( .A1(n8626), .A2(n8541), .B1(n8540), .B2(n8539), .ZN(n8542)
         );
  XNOR2_X1 U9712 ( .A(n9026), .B(n8552), .ZN(n8544) );
  XNOR2_X1 U9713 ( .A(n8544), .B(n8700), .ZN(n8598) );
  NAND2_X1 U9714 ( .A1(n8596), .A2(n8598), .ZN(n8546) );
  NAND2_X1 U9715 ( .A1(n8544), .A2(n8887), .ZN(n8545) );
  NAND2_X1 U9716 ( .A1(n8546), .A2(n8545), .ZN(n8673) );
  INV_X1 U9717 ( .A(n8673), .ZN(n8547) );
  XNOR2_X1 U9718 ( .A(n9086), .B(n6592), .ZN(n8674) );
  NAND2_X1 U9719 ( .A1(n8674), .A2(n8859), .ZN(n8548) );
  XNOR2_X1 U9720 ( .A(n9080), .B(n6861), .ZN(n8550) );
  XNOR2_X1 U9721 ( .A(n8550), .B(n8554), .ZN(n8559) );
  INV_X1 U9722 ( .A(n8550), .ZN(n8551) );
  XNOR2_X1 U9723 ( .A(n8842), .B(n8552), .ZN(n8553) );
  AOI22_X1 U9724 ( .A1(n8554), .A2(n8676), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8556) );
  NAND2_X1 U9725 ( .A1(n8851), .A2(n8694), .ZN(n8555) );
  OAI211_X1 U9726 ( .C1(n8846), .C2(n8679), .A(n8556), .B(n8555), .ZN(n8557)
         );
  AOI21_X1 U9727 ( .B1(n9074), .B2(n8681), .A(n8557), .ZN(n8558) );
  XNOR2_X1 U9728 ( .A(n8560), .B(n8559), .ZN(n8565) );
  AOI22_X1 U9729 ( .A1(n8858), .A2(n8689), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8562) );
  NAND2_X1 U9730 ( .A1(n8862), .A2(n8694), .ZN(n8561) );
  OAI211_X1 U9731 ( .C1(n8879), .C2(n8691), .A(n8562), .B(n8561), .ZN(n8563)
         );
  AOI21_X1 U9732 ( .B1(n9080), .B2(n8681), .A(n8563), .ZN(n8564) );
  OAI21_X1 U9733 ( .B1(n8565), .B2(n8683), .A(n8564), .ZN(P2_U3154) );
  XNOR2_X1 U9734 ( .A(n8567), .B(n8566), .ZN(n8568) );
  NAND2_X1 U9735 ( .A1(n8568), .A2(n8685), .ZN(n8574) );
  NOR2_X1 U9736 ( .A1(n8610), .A2(n8679), .ZN(n8571) );
  INV_X1 U9737 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10115) );
  OAI22_X1 U9738 ( .A1(n8569), .A2(n8691), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10115), .ZN(n8570) );
  AOI211_X1 U9739 ( .C1(n8694), .C2(n8572), .A(n8571), .B(n8570), .ZN(n8573)
         );
  OAI211_X1 U9740 ( .C1(n8575), .C2(n8697), .A(n8574), .B(n8573), .ZN(P2_U3155) );
  XNOR2_X1 U9741 ( .A(n8576), .B(n8623), .ZN(n8625) );
  XNOR2_X1 U9742 ( .A(n8625), .B(n8907), .ZN(n8581) );
  AOI22_X1 U9743 ( .A1(n8701), .A2(n8689), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8578) );
  NAND2_X1 U9744 ( .A1(n8694), .A2(n8901), .ZN(n8577) );
  OAI211_X1 U9745 ( .C1(n8919), .C2(n8691), .A(n8578), .B(n8577), .ZN(n8579)
         );
  AOI21_X1 U9746 ( .B1(n8902), .B2(n8681), .A(n8579), .ZN(n8580) );
  OAI21_X1 U9747 ( .B1(n8581), .B2(n8683), .A(n8580), .ZN(P2_U3156) );
  OAI211_X1 U9748 ( .C1(n8584), .C2(n8583), .A(n8582), .B(n8685), .ZN(n8588)
         );
  NOR2_X1 U9749 ( .A1(n10239), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8783) );
  AOI21_X1 U9750 ( .B1(n8704), .B2(n8689), .A(n8783), .ZN(n8585) );
  OAI21_X1 U9751 ( .B1(n8945), .B2(n8691), .A(n8585), .ZN(n8586) );
  AOI21_X1 U9752 ( .B1(n8694), .B2(n8946), .A(n8586), .ZN(n8587) );
  OAI211_X1 U9753 ( .C1(n9120), .C2(n8697), .A(n8588), .B(n8587), .ZN(P2_U3159) );
  XOR2_X1 U9754 ( .A(n8590), .B(n8589), .Z(n8595) );
  NAND2_X1 U9755 ( .A1(n8694), .A2(n8923), .ZN(n8592) );
  AOI22_X1 U9756 ( .A1(n8702), .A2(n8689), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8591) );
  OAI211_X1 U9757 ( .C1(n8944), .C2(n8691), .A(n8592), .B(n8591), .ZN(n8593)
         );
  AOI21_X1 U9758 ( .B1(n8922), .B2(n8681), .A(n8593), .ZN(n8594) );
  OAI21_X1 U9759 ( .B1(n8595), .B2(n8683), .A(n8594), .ZN(P2_U3163) );
  XOR2_X1 U9760 ( .A(n8598), .B(n8597), .Z(n8603) );
  AOI22_X1 U9761 ( .A1(n8701), .A2(n8676), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8600) );
  NAND2_X1 U9762 ( .A1(n8694), .A2(n8882), .ZN(n8599) );
  OAI211_X1 U9763 ( .C1(n8879), .C2(n8679), .A(n8600), .B(n8599), .ZN(n8601)
         );
  AOI21_X1 U9764 ( .B1(n9026), .B2(n8681), .A(n8601), .ZN(n8602) );
  OAI21_X1 U9765 ( .B1(n8603), .B2(n8683), .A(n8602), .ZN(P2_U3165) );
  XNOR2_X1 U9766 ( .A(n8605), .B(n8996), .ZN(n8606) );
  XNOR2_X1 U9767 ( .A(n8604), .B(n8606), .ZN(n8613) );
  NAND2_X1 U9768 ( .A1(n8694), .A2(n8982), .ZN(n8609) );
  INV_X1 U9769 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8607) );
  NOR2_X1 U9770 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8607), .ZN(n10466) );
  AOI21_X1 U9771 ( .B1(n8979), .B2(n8689), .A(n10466), .ZN(n8608) );
  OAI211_X1 U9772 ( .C1(n8610), .C2(n8691), .A(n8609), .B(n8608), .ZN(n8611)
         );
  AOI21_X1 U9773 ( .B1(n9135), .B2(n8681), .A(n8611), .ZN(n8612) );
  OAI21_X1 U9774 ( .B1(n8613), .B2(n8683), .A(n8612), .ZN(P2_U3166) );
  XNOR2_X1 U9775 ( .A(n8615), .B(n8979), .ZN(n8616) );
  XNOR2_X1 U9776 ( .A(n8614), .B(n8616), .ZN(n8622) );
  NAND2_X1 U9777 ( .A1(n8694), .A2(n8970), .ZN(n8618) );
  NOR2_X1 U9778 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6985), .ZN(n10485) );
  AOI21_X1 U9779 ( .B1(n8967), .B2(n8689), .A(n10485), .ZN(n8617) );
  OAI211_X1 U9780 ( .C1(n8619), .C2(n8691), .A(n8618), .B(n8617), .ZN(n8620)
         );
  AOI21_X1 U9781 ( .B1(n9129), .B2(n8681), .A(n8620), .ZN(n8621) );
  OAI21_X1 U9782 ( .B1(n8622), .B2(n8683), .A(n8621), .ZN(P2_U3168) );
  OAI22_X1 U9783 ( .A1(n8625), .A2(n8624), .B1(n8623), .B2(n8576), .ZN(n8628)
         );
  XNOR2_X1 U9784 ( .A(n8626), .B(n8898), .ZN(n8627) );
  XNOR2_X1 U9785 ( .A(n8628), .B(n8627), .ZN(n8634) );
  AOI22_X1 U9786 ( .A1(n8700), .A2(n8689), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8630) );
  NAND2_X1 U9787 ( .A1(n8694), .A2(n8889), .ZN(n8629) );
  OAI211_X1 U9788 ( .C1(n8907), .C2(n8691), .A(n8630), .B(n8629), .ZN(n8631)
         );
  AOI21_X1 U9789 ( .B1(n8632), .B2(n8681), .A(n8631), .ZN(n8633) );
  OAI21_X1 U9790 ( .B1(n8634), .B2(n8683), .A(n8633), .ZN(P2_U3169) );
  INV_X1 U9791 ( .A(n8635), .ZN(n8636) );
  AOI21_X1 U9792 ( .B1(n8638), .B2(n8637), .A(n8636), .ZN(n8644) );
  NAND2_X1 U9793 ( .A1(n8694), .A2(n8935), .ZN(n8640) );
  AOI22_X1 U9794 ( .A1(n8703), .A2(n8689), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8639) );
  OAI211_X1 U9795 ( .C1(n8931), .C2(n8691), .A(n8640), .B(n8639), .ZN(n8641)
         );
  AOI21_X1 U9796 ( .B1(n8642), .B2(n8681), .A(n8641), .ZN(n8643) );
  OAI21_X1 U9797 ( .B1(n8644), .B2(n8683), .A(n8643), .ZN(P2_U3173) );
  XNOR2_X1 U9798 ( .A(n8645), .B(n8705), .ZN(n8646) );
  XNOR2_X1 U9799 ( .A(n8647), .B(n8646), .ZN(n8654) );
  NAND2_X1 U9800 ( .A1(n8694), .A2(n8648), .ZN(n8650) );
  NOR2_X1 U9801 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6981), .ZN(n10414) );
  AOI21_X1 U9802 ( .B1(n8706), .B2(n8676), .A(n10414), .ZN(n8649) );
  OAI211_X1 U9803 ( .C1(n8692), .C2(n8679), .A(n8650), .B(n8649), .ZN(n8651)
         );
  AOI21_X1 U9804 ( .B1(n8652), .B2(n8681), .A(n8651), .ZN(n8653) );
  OAI21_X1 U9805 ( .B1(n8654), .B2(n8683), .A(n8653), .ZN(P2_U3174) );
  INV_X1 U9806 ( .A(n9035), .ZN(n8912) );
  AOI21_X1 U9807 ( .B1(n8656), .B2(n8655), .A(n8683), .ZN(n8658) );
  NAND2_X1 U9808 ( .A1(n8658), .A2(n8657), .ZN(n8662) );
  AOI22_X1 U9809 ( .A1(n8703), .A2(n8676), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8659) );
  OAI21_X1 U9810 ( .B1(n8907), .B2(n8679), .A(n8659), .ZN(n8660) );
  AOI21_X1 U9811 ( .B1(n8910), .B2(n8694), .A(n8660), .ZN(n8661) );
  OAI211_X1 U9812 ( .C1(n8912), .C2(n8697), .A(n8662), .B(n8661), .ZN(P2_U3175) );
  AOI21_X1 U9813 ( .B1(n8664), .B2(n8663), .A(n8683), .ZN(n8666) );
  NAND2_X1 U9814 ( .A1(n8666), .A2(n8665), .ZN(n8671) );
  INV_X1 U9815 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10153) );
  NOR2_X1 U9816 ( .A1(n10153), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10497) );
  AOI21_X1 U9817 ( .B1(n8957), .B2(n8689), .A(n10497), .ZN(n8667) );
  OAI21_X1 U9818 ( .B1(n8668), .B2(n8691), .A(n8667), .ZN(n8669) );
  AOI21_X1 U9819 ( .B1(n8694), .B2(n8959), .A(n8669), .ZN(n8670) );
  OAI211_X1 U9820 ( .C1(n8672), .C2(n8697), .A(n8671), .B(n8670), .ZN(P2_U3178) );
  XNOR2_X1 U9821 ( .A(n8674), .B(n8859), .ZN(n8675) );
  XNOR2_X1 U9822 ( .A(n8673), .B(n8675), .ZN(n8684) );
  AOI22_X1 U9823 ( .A1(n8700), .A2(n8676), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8678) );
  NAND2_X1 U9824 ( .A1(n8871), .A2(n8694), .ZN(n8677) );
  OAI211_X1 U9825 ( .C1(n8869), .C2(n8679), .A(n8678), .B(n8677), .ZN(n8680)
         );
  AOI21_X1 U9826 ( .B1(n9086), .B2(n8681), .A(n8680), .ZN(n8682) );
  OAI21_X1 U9827 ( .B1(n8684), .B2(n8683), .A(n8682), .ZN(P2_U3180) );
  OAI211_X1 U9828 ( .C1(n8688), .C2(n8687), .A(n8686), .B(n8685), .ZN(n8696)
         );
  NOR2_X1 U9829 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6983), .ZN(n10448) );
  AOI21_X1 U9830 ( .B1(n8996), .B2(n8689), .A(n10448), .ZN(n8690) );
  OAI21_X1 U9831 ( .B1(n8692), .B2(n8691), .A(n8690), .ZN(n8693) );
  AOI21_X1 U9832 ( .B1(n8988), .B2(n8694), .A(n8693), .ZN(n8695) );
  OAI211_X1 U9833 ( .C1(n8698), .C2(n8697), .A(n8696), .B(n8695), .ZN(P2_U3181) );
  MUX2_X1 U9834 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8836), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9835 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8699), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9836 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8858), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9837 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8700), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9838 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8701), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9839 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8702), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9840 ( .A(n8703), .B(P2_DATAO_REG_21__SCAN_IN), .S(n10503), .Z(
        P2_U3512) );
  MUX2_X1 U9841 ( .A(n8704), .B(P2_DATAO_REG_20__SCAN_IN), .S(n10503), .Z(
        P2_U3511) );
  MUX2_X1 U9842 ( .A(n8957), .B(P2_DATAO_REG_19__SCAN_IN), .S(n10503), .Z(
        P2_U3510) );
  MUX2_X1 U9843 ( .A(n8967), .B(P2_DATAO_REG_18__SCAN_IN), .S(n10503), .Z(
        P2_U3509) );
  MUX2_X1 U9844 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8979), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9845 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8996), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9846 ( .A(n8978), .B(P2_DATAO_REG_15__SCAN_IN), .S(n10503), .Z(
        P2_U3506) );
  MUX2_X1 U9847 ( .A(n8993), .B(P2_DATAO_REG_14__SCAN_IN), .S(n10503), .Z(
        P2_U3505) );
  MUX2_X1 U9848 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8705), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9849 ( .A(n8706), .B(P2_DATAO_REG_12__SCAN_IN), .S(n10503), .Z(
        P2_U3503) );
  MUX2_X1 U9850 ( .A(n8707), .B(P2_DATAO_REG_11__SCAN_IN), .S(n10503), .Z(
        P2_U3502) );
  MUX2_X1 U9851 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8708), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U9852 ( .A(n8709), .B(P2_DATAO_REG_9__SCAN_IN), .S(n10503), .Z(
        P2_U3500) );
  MUX2_X1 U9853 ( .A(n8710), .B(P2_DATAO_REG_8__SCAN_IN), .S(n10503), .Z(
        P2_U3499) );
  MUX2_X1 U9854 ( .A(n8711), .B(P2_DATAO_REG_7__SCAN_IN), .S(n10503), .Z(
        P2_U3498) );
  MUX2_X1 U9855 ( .A(n8712), .B(P2_DATAO_REG_6__SCAN_IN), .S(n10503), .Z(
        P2_U3497) );
  MUX2_X1 U9856 ( .A(n8713), .B(P2_DATAO_REG_5__SCAN_IN), .S(n10503), .Z(
        P2_U3496) );
  MUX2_X1 U9857 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8714), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U9858 ( .A(n8715), .B(P2_DATAO_REG_3__SCAN_IN), .S(n10503), .Z(
        P2_U3494) );
  MUX2_X1 U9859 ( .A(n8716), .B(P2_DATAO_REG_2__SCAN_IN), .S(n10503), .Z(
        P2_U3493) );
  MUX2_X1 U9860 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6942), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U9861 ( .A(n8717), .B(P2_DATAO_REG_0__SCAN_IN), .S(n10503), .Z(
        P2_U3491) );
  AOI21_X1 U9862 ( .B1(n8720), .B2(n8719), .A(n8718), .ZN(n8811) );
  INV_X1 U9863 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U9864 ( .A1(n8825), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8721) );
  OAI211_X1 U9865 ( .C1(n8825), .C2(n8722), .A(n8745), .B(n8721), .ZN(n8810)
         );
  INV_X1 U9866 ( .A(n8810), .ZN(n8726) );
  OR2_X1 U9867 ( .A1(n8825), .A2(n8765), .ZN(n8725) );
  INV_X1 U9868 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8746) );
  OR2_X1 U9869 ( .A1(n8745), .A2(n8746), .ZN(n8754) );
  INV_X1 U9870 ( .A(n8754), .ZN(n8723) );
  NAND2_X1 U9871 ( .A1(n8825), .A2(n8723), .ZN(n8724) );
  NAND2_X1 U9872 ( .A1(n8725), .A2(n8724), .ZN(n8809) );
  NOR2_X1 U9873 ( .A1(n8726), .A2(n8809), .ZN(n8728) );
  NAND2_X1 U9874 ( .A1(n8811), .A2(n8728), .ZN(n8727) );
  OAI211_X1 U9875 ( .C1(n8811), .C2(n8728), .A(n10513), .B(n8727), .ZN(n8752)
         );
  OAI21_X1 U9876 ( .B1(n8731), .B2(P2_REG2_REG_10__SCAN_IN), .A(n8765), .ZN(
        n8732) );
  AOI21_X1 U9877 ( .B1(n8733), .B2(n8732), .A(n8767), .ZN(n8734) );
  NOR2_X1 U9878 ( .A1(n10489), .A2(n8734), .ZN(n8740) );
  INV_X1 U9879 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8737) );
  INV_X1 U9880 ( .A(n8735), .ZN(n8736) );
  OAI21_X1 U9881 ( .B1(n8738), .B2(n8737), .A(n8736), .ZN(n8739) );
  AOI211_X1 U9882 ( .C1(n10476), .C2(n8745), .A(n8740), .B(n8739), .ZN(n8751)
         );
  NAND2_X1 U9883 ( .A1(n8742), .A2(n8741), .ZN(n8744) );
  NAND2_X1 U9884 ( .A1(n8744), .A2(n8743), .ZN(n8748) );
  MUX2_X1 U9885 ( .A(n8746), .B(P2_REG1_REG_10__SCAN_IN), .S(n8745), .Z(n8747)
         );
  NAND2_X1 U9886 ( .A1(n8747), .A2(n8748), .ZN(n8753) );
  OAI21_X1 U9887 ( .B1(n8748), .B2(n8747), .A(n8753), .ZN(n8749) );
  NAND2_X1 U9888 ( .A1(n8749), .A2(n10483), .ZN(n8750) );
  NAND3_X1 U9889 ( .A1(n8752), .A2(n8751), .A3(n8750), .ZN(P2_U3192) );
  INV_X1 U9890 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9057) );
  AOI22_X1 U9891 ( .A1(n10457), .A2(n9057), .B1(P2_REG1_REG_16__SCAN_IN), .B2(
        n8787), .ZN(n10460) );
  INV_X1 U9892 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8759) );
  AOI22_X1 U9893 ( .A1(n10423), .A2(n8759), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n8795), .ZN(n10426) );
  INV_X1 U9894 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10700) );
  AOI22_X1 U9895 ( .A1(n10388), .A2(n10700), .B1(P2_REG1_REG_12__SCAN_IN), 
        .B2(n8804), .ZN(n10391) );
  NAND2_X1 U9896 ( .A1(n8754), .A2(n8753), .ZN(n8755) );
  NAND2_X1 U9897 ( .A1(n8808), .A2(n8755), .ZN(n8756) );
  XNOR2_X1 U9898 ( .A(n8755), .B(n10371), .ZN(n10373) );
  NAND2_X1 U9899 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n10373), .ZN(n10372) );
  NAND2_X1 U9900 ( .A1(n8799), .A2(n8757), .ZN(n8758) );
  NAND2_X1 U9901 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n10408), .ZN(n10407) );
  NAND2_X1 U9902 ( .A1(n8791), .A2(n8760), .ZN(n8761) );
  NAND2_X1 U9903 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n10442), .ZN(n10441) );
  NAND2_X1 U9904 ( .A1(n8819), .A2(n8762), .ZN(n8763) );
  NAND2_X1 U9905 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n10478), .ZN(n10477) );
  XNOR2_X1 U9906 ( .A(n10510), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n10494) );
  AOI22_X1 U9907 ( .A1(n10495), .A2(n10494), .B1(P2_REG1_REG_18__SCAN_IN), 
        .B2(n10512), .ZN(n8764) );
  XNOR2_X1 U9908 ( .A(n8833), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8824) );
  XNOR2_X1 U9909 ( .A(n8764), .B(n8824), .ZN(n8834) );
  INV_X1 U9910 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n10486) );
  INV_X1 U9911 ( .A(n8765), .ZN(n8766) );
  NOR2_X1 U9912 ( .A1(n10371), .A2(n8768), .ZN(n8769) );
  MUX2_X1 U9913 ( .A(n8801), .B(P2_REG2_REG_12__SCAN_IN), .S(n10388), .Z(n8770) );
  INV_X1 U9914 ( .A(n8770), .ZN(n10399) );
  NOR2_X1 U9915 ( .A1(n10406), .A2(n8771), .ZN(n8772) );
  INV_X1 U9916 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10416) );
  XNOR2_X1 U9917 ( .A(n8795), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n10433) );
  NOR2_X1 U9918 ( .A1(n10440), .A2(n8773), .ZN(n8774) );
  INV_X1 U9919 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n10450) );
  XNOR2_X1 U9920 ( .A(n10440), .B(n8773), .ZN(n10451) );
  INV_X1 U9921 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8776) );
  NOR2_X1 U9922 ( .A1(n8787), .A2(n8776), .ZN(n8775) );
  AOI21_X1 U9923 ( .B1(n8776), .B2(n8787), .A(n8775), .ZN(n10468) );
  INV_X1 U9924 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8777) );
  MUX2_X1 U9925 ( .A(P2_REG2_REG_18__SCAN_IN), .B(n8777), .S(n10510), .Z(
        n10507) );
  NOR2_X1 U9926 ( .A1(n10505), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8779) );
  INV_X1 U9927 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8780) );
  MUX2_X1 U9928 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8780), .S(n8833), .Z(n8827)
         );
  XOR2_X1 U9929 ( .A(n8781), .B(n8827), .Z(n8782) );
  AOI21_X1 U9930 ( .B1(n10498), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n8783), .ZN(
        n8784) );
  MUX2_X1 U9931 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8825), .Z(n8820) );
  XNOR2_X1 U9932 ( .A(n8820), .B(n10475), .ZN(n10481) );
  OR2_X1 U9933 ( .A1(n8825), .A2(n8776), .ZN(n8786) );
  NAND2_X1 U9934 ( .A1(n8825), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8785) );
  NAND2_X1 U9935 ( .A1(n8786), .A2(n8785), .ZN(n8788) );
  OR2_X1 U9936 ( .A1(n8787), .A2(n8788), .ZN(n8818) );
  XNOR2_X1 U9937 ( .A(n8788), .B(n10457), .ZN(n10463) );
  OR2_X1 U9938 ( .A1(n8825), .A2(n10450), .ZN(n8790) );
  NAND2_X1 U9939 ( .A1(n8825), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8789) );
  NAND2_X1 U9940 ( .A1(n8790), .A2(n8789), .ZN(n8792) );
  OR2_X1 U9941 ( .A1(n8791), .A2(n8792), .ZN(n8817) );
  XNOR2_X1 U9942 ( .A(n8792), .B(n10440), .ZN(n10445) );
  OR2_X1 U9943 ( .A1(n8825), .A2(n5096), .ZN(n8794) );
  NAND2_X1 U9944 ( .A1(n8825), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8793) );
  NAND2_X1 U9945 ( .A1(n8794), .A2(n8793), .ZN(n8796) );
  OR2_X1 U9946 ( .A1(n8795), .A2(n8796), .ZN(n8816) );
  XNOR2_X1 U9947 ( .A(n8796), .B(n10423), .ZN(n10429) );
  OR2_X1 U9948 ( .A1(n8825), .A2(n10416), .ZN(n8798) );
  NAND2_X1 U9949 ( .A1(n8825), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8797) );
  NAND2_X1 U9950 ( .A1(n8798), .A2(n8797), .ZN(n8800) );
  OR2_X1 U9951 ( .A1(n8799), .A2(n8800), .ZN(n8815) );
  XNOR2_X1 U9952 ( .A(n8800), .B(n10406), .ZN(n10411) );
  OR2_X1 U9953 ( .A1(n8825), .A2(n8801), .ZN(n8803) );
  NAND2_X1 U9954 ( .A1(n8825), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8802) );
  NAND2_X1 U9955 ( .A1(n8803), .A2(n8802), .ZN(n8805) );
  OR2_X1 U9956 ( .A1(n8804), .A2(n8805), .ZN(n8814) );
  XNOR2_X1 U9957 ( .A(n8805), .B(n10388), .ZN(n10394) );
  OR2_X1 U9958 ( .A1(n8825), .A2(n10381), .ZN(n8807) );
  NAND2_X1 U9959 ( .A1(n8825), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8806) );
  NAND2_X1 U9960 ( .A1(n8807), .A2(n8806), .ZN(n8812) );
  OR2_X1 U9961 ( .A1(n8808), .A2(n8812), .ZN(n8813) );
  AOI21_X1 U9962 ( .B1(n8811), .B2(n8810), .A(n8809), .ZN(n10375) );
  XNOR2_X1 U9963 ( .A(n8812), .B(n10371), .ZN(n10376) );
  NAND2_X1 U9964 ( .A1(n10375), .A2(n10376), .ZN(n10374) );
  NAND2_X1 U9965 ( .A1(n8813), .A2(n10374), .ZN(n10393) );
  NAND2_X1 U9966 ( .A1(n10394), .A2(n10393), .ZN(n10392) );
  NAND2_X1 U9967 ( .A1(n8814), .A2(n10392), .ZN(n10410) );
  NAND2_X1 U9968 ( .A1(n10411), .A2(n10410), .ZN(n10409) );
  NAND2_X1 U9969 ( .A1(n8815), .A2(n10409), .ZN(n10428) );
  NAND2_X1 U9970 ( .A1(n10429), .A2(n10428), .ZN(n10427) );
  NAND2_X1 U9971 ( .A1(n8816), .A2(n10427), .ZN(n10444) );
  NAND2_X1 U9972 ( .A1(n10445), .A2(n10444), .ZN(n10443) );
  NAND2_X1 U9973 ( .A1(n8817), .A2(n10443), .ZN(n10462) );
  NAND2_X1 U9974 ( .A1(n10463), .A2(n10462), .ZN(n10461) );
  NAND2_X1 U9975 ( .A1(n8818), .A2(n10461), .ZN(n10480) );
  NAND2_X1 U9976 ( .A1(n10481), .A2(n10480), .ZN(n10479) );
  OAI21_X1 U9977 ( .B1(n8820), .B2(n8819), .A(n10479), .ZN(n8823) );
  NOR2_X1 U9978 ( .A1(n8825), .A2(n8777), .ZN(n8821) );
  AOI21_X1 U9979 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n8825), .A(n8821), .ZN(
        n8822) );
  NOR2_X1 U9980 ( .A1(n8823), .A2(n8822), .ZN(n10499) );
  NAND2_X1 U9981 ( .A1(n8823), .A2(n8822), .ZN(n10500) );
  OAI21_X1 U9982 ( .B1(n10499), .B2(n10512), .A(n10500), .ZN(n8829) );
  INV_X1 U9983 ( .A(n8824), .ZN(n8826) );
  MUX2_X1 U9984 ( .A(n8827), .B(n8826), .S(n8825), .Z(n8828) );
  XNOR2_X1 U9985 ( .A(n8829), .B(n8828), .ZN(n8831) );
  NOR2_X1 U9986 ( .A1(n8831), .A2(n8830), .ZN(n8832) );
  NAND2_X1 U9987 ( .A1(n8836), .A2(n8835), .ZN(n9065) );
  INV_X1 U9988 ( .A(n9065), .ZN(n8838) );
  NOR3_X1 U9989 ( .A1(n8838), .A2(n10580), .A3(n8837), .ZN(n8841) );
  NOR2_X1 U9990 ( .A1(n10577), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8839) );
  OAI22_X1 U9991 ( .A1(n9067), .A2(n8937), .B1(n8841), .B2(n8839), .ZN(
        P2_U3202) );
  NOR2_X1 U9992 ( .A1(n10577), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8840) );
  OAI22_X1 U9993 ( .A1(n9070), .A2(n8937), .B1(n8841), .B2(n8840), .ZN(
        P2_U3203) );
  XNOR2_X1 U9994 ( .A(n8843), .B(n8842), .ZN(n9077) );
  INV_X1 U9995 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8850) );
  INV_X1 U9996 ( .A(n9014), .ZN(n9072) );
  MUX2_X1 U9997 ( .A(n8850), .B(n9072), .S(n10577), .Z(n8853) );
  AOI22_X1 U9998 ( .A1(n9074), .A2(n9001), .B1(n8983), .B2(n8851), .ZN(n8852)
         );
  OAI211_X1 U9999 ( .C1(n9077), .C2(n9004), .A(n8853), .B(n8852), .ZN(P2_U3205) );
  XNOR2_X1 U10000 ( .A(n8855), .B(n8854), .ZN(n9083) );
  INV_X1 U10001 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8861) );
  XNOR2_X1 U10002 ( .A(n8857), .B(n8856), .ZN(n8860) );
  AOI222_X1 U10003 ( .A1(n8989), .A2(n8860), .B1(n8859), .B2(n8994), .C1(n8858), .C2(n8995), .ZN(n9078) );
  MUX2_X1 U10004 ( .A(n8861), .B(n9078), .S(n10577), .Z(n8864) );
  AOI22_X1 U10005 ( .A1(n9080), .A2(n9001), .B1(n8983), .B2(n8862), .ZN(n8863)
         );
  OAI211_X1 U10006 ( .C1(n9083), .C2(n9004), .A(n8864), .B(n8863), .ZN(
        P2_U3206) );
  XNOR2_X1 U10007 ( .A(n8865), .B(n8867), .ZN(n9089) );
  INV_X1 U10008 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8870) );
  XOR2_X1 U10009 ( .A(n8867), .B(n8866), .Z(n8868) );
  OAI222_X1 U10010 ( .A1(n10566), .A2(n8869), .B1(n10564), .B2(n8887), .C1(
        n8868), .C2(n10562), .ZN(n9021) );
  INV_X1 U10011 ( .A(n9021), .ZN(n9084) );
  MUX2_X1 U10012 ( .A(n8870), .B(n9084), .S(n10577), .Z(n8873) );
  AOI22_X1 U10013 ( .A1(n9086), .A2(n9001), .B1(n8983), .B2(n8871), .ZN(n8872)
         );
  OAI211_X1 U10014 ( .C1(n9089), .C2(n9004), .A(n8873), .B(n8872), .ZN(
        P2_U3207) );
  XNOR2_X1 U10015 ( .A(n8875), .B(n8874), .ZN(n9093) );
  XNOR2_X1 U10016 ( .A(n8877), .B(n8876), .ZN(n8878) );
  OAI222_X1 U10017 ( .A1(n10564), .A2(n8898), .B1(n10566), .B2(n8879), .C1(
        n10562), .C2(n8878), .ZN(n9025) );
  NOR2_X1 U10018 ( .A1(n8880), .A2(n10571), .ZN(n8881) );
  OAI21_X1 U10019 ( .B1(n9025), .B2(n8881), .A(n10577), .ZN(n8884) );
  AOI22_X1 U10020 ( .A1(n8882), .A2(n8983), .B1(n10580), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8883) );
  OAI211_X1 U10021 ( .C1(n9093), .C2(n9004), .A(n8884), .B(n8883), .ZN(
        P2_U3208) );
  NOR2_X1 U10022 ( .A1(n9095), .A2(n10571), .ZN(n8888) );
  XNOR2_X1 U10023 ( .A(n8885), .B(n8890), .ZN(n8886) );
  OAI222_X1 U10024 ( .A1(n10564), .A2(n8907), .B1(n10566), .B2(n8887), .C1(
        n10562), .C2(n8886), .ZN(n9094) );
  AOI211_X1 U10025 ( .C1(n8983), .C2(n8889), .A(n8888), .B(n9094), .ZN(n8893)
         );
  XNOR2_X1 U10026 ( .A(n8891), .B(n8890), .ZN(n9029) );
  AOI22_X1 U10027 ( .A1(n9029), .A2(n8950), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n10580), .ZN(n8892) );
  OAI21_X1 U10028 ( .B1(n8893), .B2(n10580), .A(n8892), .ZN(P2_U3209) );
  XNOR2_X1 U10029 ( .A(n8894), .B(n8895), .ZN(n9101) );
  INV_X1 U10030 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8900) );
  XNOR2_X1 U10031 ( .A(n8896), .B(n8895), .ZN(n8897) );
  OAI222_X1 U10032 ( .A1(n10564), .A2(n8919), .B1(n10566), .B2(n8898), .C1(
        n10562), .C2(n8897), .ZN(n9099) );
  INV_X1 U10033 ( .A(n9099), .ZN(n8899) );
  MUX2_X1 U10034 ( .A(n8900), .B(n8899), .S(n10577), .Z(n8904) );
  AOI22_X1 U10035 ( .A1(n8902), .A2(n9001), .B1(n8983), .B2(n8901), .ZN(n8903)
         );
  OAI211_X1 U10036 ( .C1(n9101), .C2(n9004), .A(n8904), .B(n8903), .ZN(
        P2_U3210) );
  XNOR2_X1 U10037 ( .A(n8905), .B(n8908), .ZN(n8906) );
  OAI222_X1 U10038 ( .A1(n10564), .A2(n8932), .B1(n10566), .B2(n8907), .C1(
        n8906), .C2(n10562), .ZN(n9034) );
  INV_X1 U10039 ( .A(n9034), .ZN(n8916) );
  XNOR2_X1 U10040 ( .A(n8909), .B(n8908), .ZN(n9107) );
  INV_X1 U10041 ( .A(n9107), .ZN(n8914) );
  AOI22_X1 U10042 ( .A1(n10580), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8983), 
        .B2(n8910), .ZN(n8911) );
  OAI21_X1 U10043 ( .B1(n8912), .B2(n8937), .A(n8911), .ZN(n8913) );
  AOI21_X1 U10044 ( .B1(n8914), .B2(n8950), .A(n8913), .ZN(n8915) );
  OAI21_X1 U10045 ( .B1(n8916), .B2(n10580), .A(n8915), .ZN(P2_U3211) );
  XNOR2_X1 U10046 ( .A(n8917), .B(n8921), .ZN(n8918) );
  OAI222_X1 U10047 ( .A1(n10566), .A2(n8919), .B1(n10564), .B2(n8944), .C1(
        n8918), .C2(n10562), .ZN(n9038) );
  INV_X1 U10048 ( .A(n9038), .ZN(n8927) );
  XNOR2_X1 U10049 ( .A(n8920), .B(n8921), .ZN(n9039) );
  INV_X1 U10050 ( .A(n8922), .ZN(n9111) );
  AOI22_X1 U10051 ( .A1(n10580), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8983), 
        .B2(n8923), .ZN(n8924) );
  OAI21_X1 U10052 ( .B1(n9111), .B2(n8937), .A(n8924), .ZN(n8925) );
  AOI21_X1 U10053 ( .B1(n9039), .B2(n8950), .A(n8925), .ZN(n8926) );
  OAI21_X1 U10054 ( .B1(n8927), .B2(n10580), .A(n8926), .ZN(P2_U3212) );
  XNOR2_X1 U10055 ( .A(n8929), .B(n8928), .ZN(n8930) );
  OAI222_X1 U10056 ( .A1(n10566), .A2(n8932), .B1(n10564), .B2(n8931), .C1(
        n8930), .C2(n10562), .ZN(n9042) );
  INV_X1 U10057 ( .A(n9042), .ZN(n8940) );
  XNOR2_X1 U10058 ( .A(n8933), .B(n8934), .ZN(n9043) );
  AOI22_X1 U10059 ( .A1(n10580), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8983), 
        .B2(n8935), .ZN(n8936) );
  OAI21_X1 U10060 ( .B1(n9115), .B2(n8937), .A(n8936), .ZN(n8938) );
  AOI21_X1 U10061 ( .B1(n9043), .B2(n8950), .A(n8938), .ZN(n8939) );
  OAI21_X1 U10062 ( .B1(n8940), .B2(n10580), .A(n8939), .ZN(P2_U3213) );
  XNOR2_X1 U10063 ( .A(n8942), .B(n8941), .ZN(n8943) );
  OAI222_X1 U10064 ( .A1(n10564), .A2(n8945), .B1(n10566), .B2(n8944), .C1(
        n10562), .C2(n8943), .ZN(n9046) );
  AOI21_X1 U10065 ( .B1(n8983), .B2(n8946), .A(n9046), .ZN(n8953) );
  AOI22_X1 U10066 ( .A1(n8947), .A2(n9001), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n10580), .ZN(n8952) );
  XNOR2_X1 U10067 ( .A(n8948), .B(n8949), .ZN(n9047) );
  NAND2_X1 U10068 ( .A1(n9047), .A2(n8950), .ZN(n8951) );
  OAI211_X1 U10069 ( .C1(n8953), .C2(n10580), .A(n8952), .B(n8951), .ZN(
        P2_U3214) );
  XNOR2_X1 U10070 ( .A(n8954), .B(n8955), .ZN(n9126) );
  XNOR2_X1 U10071 ( .A(n8956), .B(n8955), .ZN(n8958) );
  AOI222_X1 U10072 ( .A1(n8989), .A2(n8958), .B1(n8957), .B2(n8995), .C1(n8979), .C2(n8994), .ZN(n9121) );
  MUX2_X1 U10073 ( .A(n8777), .B(n9121), .S(n10577), .Z(n8961) );
  AOI22_X1 U10074 ( .A1(n9123), .A2(n9001), .B1(n8983), .B2(n8959), .ZN(n8960)
         );
  OAI211_X1 U10075 ( .C1(n9126), .C2(n9004), .A(n8961), .B(n8960), .ZN(
        P2_U3215) );
  XNOR2_X1 U10076 ( .A(n8962), .B(n8963), .ZN(n9132) );
  OAI211_X1 U10077 ( .C1(n8966), .C2(n8965), .A(n8964), .B(n8989), .ZN(n8969)
         );
  AOI22_X1 U10078 ( .A1(n8996), .A2(n8994), .B1(n8995), .B2(n8967), .ZN(n8968)
         );
  MUX2_X1 U10079 ( .A(n9128), .B(n10486), .S(n10580), .Z(n8972) );
  AOI22_X1 U10080 ( .A1(n9129), .A2(n9001), .B1(n8983), .B2(n8970), .ZN(n8971)
         );
  OAI211_X1 U10081 ( .C1(n9132), .C2(n9004), .A(n8972), .B(n8971), .ZN(
        P2_U3216) );
  XNOR2_X1 U10082 ( .A(n8974), .B(n8973), .ZN(n9138) );
  OAI211_X1 U10083 ( .C1(n8977), .C2(n8976), .A(n8975), .B(n8989), .ZN(n8981)
         );
  AOI22_X1 U10084 ( .A1(n8979), .A2(n8995), .B1(n8994), .B2(n8978), .ZN(n8980)
         );
  MUX2_X1 U10085 ( .A(n9134), .B(n8776), .S(n10580), .Z(n8985) );
  AOI22_X1 U10086 ( .A1(n9135), .A2(n9001), .B1(n8983), .B2(n8982), .ZN(n8984)
         );
  OAI211_X1 U10087 ( .C1(n9138), .C2(n9004), .A(n8985), .B(n8984), .ZN(
        P2_U3217) );
  XNOR2_X1 U10088 ( .A(n8987), .B(n8986), .ZN(n9146) );
  INV_X1 U10089 ( .A(n8988), .ZN(n8999) );
  OAI211_X1 U10090 ( .C1(n8992), .C2(n8991), .A(n8990), .B(n8989), .ZN(n8998)
         );
  AOI22_X1 U10091 ( .A1(n8996), .A2(n8995), .B1(n8994), .B2(n8993), .ZN(n8997)
         );
  OAI21_X1 U10092 ( .B1(n8999), .B2(n10570), .A(n9140), .ZN(n9000) );
  NAND2_X1 U10093 ( .A1(n9000), .A2(n10577), .ZN(n9003) );
  AOI22_X1 U10094 ( .A1(n9142), .A2(n9001), .B1(P2_REG2_REG_15__SCAN_IN), .B2(
        n10580), .ZN(n9002) );
  OAI211_X1 U10095 ( .C1(n9146), .C2(n9004), .A(n9003), .B(n9002), .ZN(
        P2_U3218) );
  NOR2_X1 U10096 ( .A1(n9065), .A2(n10721), .ZN(n9006) );
  AOI21_X1 U10097 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10721), .A(n9006), .ZN(
        n9005) );
  OAI21_X1 U10098 ( .B1(n9067), .B2(n9050), .A(n9005), .ZN(P2_U3490) );
  AOI21_X1 U10099 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n10721), .A(n9006), .ZN(
        n9007) );
  OAI21_X1 U10100 ( .B1(n9070), .B2(n9050), .A(n9007), .ZN(P2_U3489) );
  NAND2_X1 U10101 ( .A1(n9009), .A2(n9008), .ZN(n9011) );
  MUX2_X1 U10102 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9071), .S(n10723), .Z(
        P2_U3488) );
  MUX2_X1 U10103 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9014), .S(n10723), .Z(
        n9017) );
  OAI22_X1 U10104 ( .A1(n9077), .A2(n9064), .B1(n9015), .B2(n9050), .ZN(n9016)
         );
  OR2_X1 U10105 ( .A1(n9017), .A2(n9016), .ZN(P2_U3487) );
  INV_X1 U10106 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9018) );
  MUX2_X1 U10107 ( .A(n9018), .B(n9078), .S(n10723), .Z(n9020) );
  NAND2_X1 U10108 ( .A1(n9080), .A2(n9061), .ZN(n9019) );
  OAI211_X1 U10109 ( .C1(n9064), .C2(n9083), .A(n9020), .B(n9019), .ZN(
        P2_U3486) );
  MUX2_X1 U10110 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9021), .S(n10723), .Z(
        n9024) );
  OAI22_X1 U10111 ( .A1(n9089), .A2(n9064), .B1(n9022), .B2(n9050), .ZN(n9023)
         );
  OR2_X1 U10112 ( .A1(n9024), .A2(n9023), .ZN(P2_U3485) );
  INV_X1 U10113 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9027) );
  AOI21_X1 U10114 ( .B1(n10671), .B2(n9026), .A(n9025), .ZN(n9090) );
  MUX2_X1 U10115 ( .A(n9027), .B(n9090), .S(n10723), .Z(n9028) );
  OAI21_X1 U10116 ( .B1(n9093), .B2(n9064), .A(n9028), .ZN(P2_U3484) );
  MUX2_X1 U10117 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9094), .S(n10723), .Z(
        n9031) );
  INV_X1 U10118 ( .A(n9029), .ZN(n9096) );
  OAI22_X1 U10119 ( .A1(n9096), .A2(n9064), .B1(n9095), .B2(n9050), .ZN(n9030)
         );
  OR2_X1 U10120 ( .A1(n9031), .A2(n9030), .ZN(P2_U3483) );
  MUX2_X1 U10121 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9099), .S(n10723), .Z(
        n9033) );
  OAI22_X1 U10122 ( .A1(n9101), .A2(n9064), .B1(n9100), .B2(n9050), .ZN(n9032)
         );
  OR2_X1 U10123 ( .A1(n9033), .A2(n9032), .ZN(P2_U3482) );
  INV_X1 U10124 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9036) );
  AOI21_X1 U10125 ( .B1(n10671), .B2(n9035), .A(n9034), .ZN(n9104) );
  MUX2_X1 U10126 ( .A(n9036), .B(n9104), .S(n10723), .Z(n9037) );
  OAI21_X1 U10127 ( .B1(n9064), .B2(n9107), .A(n9037), .ZN(P2_U3481) );
  INV_X1 U10128 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9040) );
  AOI21_X1 U10129 ( .B1(n9039), .B2(n10720), .A(n9038), .ZN(n9108) );
  MUX2_X1 U10130 ( .A(n9040), .B(n9108), .S(n10723), .Z(n9041) );
  OAI21_X1 U10131 ( .B1(n9111), .B2(n9050), .A(n9041), .ZN(P2_U3480) );
  INV_X1 U10132 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9044) );
  AOI21_X1 U10133 ( .B1(n9043), .B2(n10720), .A(n9042), .ZN(n9112) );
  MUX2_X1 U10134 ( .A(n9044), .B(n9112), .S(n10723), .Z(n9045) );
  OAI21_X1 U10135 ( .B1(n9115), .B2(n9050), .A(n9045), .ZN(P2_U3479) );
  INV_X1 U10136 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9048) );
  AOI21_X1 U10137 ( .B1(n9047), .B2(n10720), .A(n9046), .ZN(n9116) );
  MUX2_X1 U10138 ( .A(n9048), .B(n9116), .S(n10723), .Z(n9049) );
  OAI21_X1 U10139 ( .B1(n9120), .B2(n9050), .A(n9049), .ZN(P2_U3478) );
  INV_X1 U10140 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9051) );
  MUX2_X1 U10141 ( .A(n9051), .B(n9121), .S(n10723), .Z(n9053) );
  NAND2_X1 U10142 ( .A1(n9123), .A2(n9061), .ZN(n9052) );
  OAI211_X1 U10143 ( .C1(n9126), .C2(n9064), .A(n9053), .B(n9052), .ZN(
        P2_U3477) );
  INV_X1 U10144 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9054) );
  MUX2_X1 U10145 ( .A(n9128), .B(n9054), .S(n10721), .Z(n9056) );
  NAND2_X1 U10146 ( .A1(n9129), .A2(n9061), .ZN(n9055) );
  OAI211_X1 U10147 ( .C1(n9064), .C2(n9132), .A(n9056), .B(n9055), .ZN(
        P2_U3476) );
  MUX2_X1 U10148 ( .A(n9134), .B(n9057), .S(n10721), .Z(n9059) );
  NAND2_X1 U10149 ( .A1(n9135), .A2(n9061), .ZN(n9058) );
  OAI211_X1 U10150 ( .C1(n9064), .C2(n9138), .A(n9059), .B(n9058), .ZN(
        P2_U3475) );
  INV_X1 U10151 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9060) );
  MUX2_X1 U10152 ( .A(n9140), .B(n9060), .S(n10721), .Z(n9063) );
  NAND2_X1 U10153 ( .A1(n9142), .A2(n9061), .ZN(n9062) );
  OAI211_X1 U10154 ( .C1(n9146), .C2(n9064), .A(n9063), .B(n9062), .ZN(
        P2_U3474) );
  NOR2_X1 U10155 ( .A1(n9065), .A2(n10724), .ZN(n9068) );
  AOI21_X1 U10156 ( .B1(P2_REG0_REG_31__SCAN_IN), .B2(n10724), .A(n9068), .ZN(
        n9066) );
  OAI21_X1 U10157 ( .B1(n9067), .B2(n9119), .A(n9066), .ZN(P2_U3458) );
  AOI21_X1 U10158 ( .B1(P2_REG0_REG_30__SCAN_IN), .B2(n10724), .A(n9068), .ZN(
        n9069) );
  OAI21_X1 U10159 ( .B1(n9070), .B2(n9119), .A(n9069), .ZN(P2_U3457) );
  MUX2_X1 U10160 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9071), .S(n10727), .Z(
        P2_U3456) );
  MUX2_X1 U10161 ( .A(n9073), .B(n9072), .S(n10727), .Z(n9076) );
  NAND2_X1 U10162 ( .A1(n9074), .A2(n9141), .ZN(n9075) );
  OAI211_X1 U10163 ( .C1(n9077), .C2(n9145), .A(n9076), .B(n9075), .ZN(
        P2_U3455) );
  MUX2_X1 U10164 ( .A(n9079), .B(n9078), .S(n10727), .Z(n9082) );
  NAND2_X1 U10165 ( .A1(n9080), .A2(n9141), .ZN(n9081) );
  OAI211_X1 U10166 ( .C1(n9083), .C2(n9145), .A(n9082), .B(n9081), .ZN(
        P2_U3454) );
  MUX2_X1 U10167 ( .A(n9085), .B(n9084), .S(n10727), .Z(n9088) );
  NAND2_X1 U10168 ( .A1(n9086), .A2(n9141), .ZN(n9087) );
  OAI211_X1 U10169 ( .C1(n9089), .C2(n9145), .A(n9088), .B(n9087), .ZN(
        P2_U3453) );
  MUX2_X1 U10170 ( .A(n9091), .B(n9090), .S(n10727), .Z(n9092) );
  OAI21_X1 U10171 ( .B1(n9093), .B2(n9145), .A(n9092), .ZN(P2_U3452) );
  MUX2_X1 U10172 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9094), .S(n10727), .Z(
        n9098) );
  OAI22_X1 U10173 ( .A1(n9096), .A2(n9145), .B1(n9095), .B2(n9119), .ZN(n9097)
         );
  OR2_X1 U10174 ( .A1(n9098), .A2(n9097), .ZN(P2_U3451) );
  MUX2_X1 U10175 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9099), .S(n10727), .Z(
        n9103) );
  OAI22_X1 U10176 ( .A1(n9101), .A2(n9145), .B1(n9100), .B2(n9119), .ZN(n9102)
         );
  OR2_X1 U10177 ( .A1(n9103), .A2(n9102), .ZN(P2_U3450) );
  MUX2_X1 U10178 ( .A(n9105), .B(n9104), .S(n10727), .Z(n9106) );
  OAI21_X1 U10179 ( .B1(n9107), .B2(n9145), .A(n9106), .ZN(P2_U3449) );
  INV_X1 U10180 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9109) );
  MUX2_X1 U10181 ( .A(n9109), .B(n9108), .S(n10727), .Z(n9110) );
  OAI21_X1 U10182 ( .B1(n9111), .B2(n9119), .A(n9110), .ZN(P2_U3448) );
  INV_X1 U10183 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9113) );
  MUX2_X1 U10184 ( .A(n9113), .B(n9112), .S(n10727), .Z(n9114) );
  OAI21_X1 U10185 ( .B1(n9115), .B2(n9119), .A(n9114), .ZN(P2_U3447) );
  INV_X1 U10186 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9117) );
  MUX2_X1 U10187 ( .A(n9117), .B(n9116), .S(n10727), .Z(n9118) );
  OAI21_X1 U10188 ( .B1(n9120), .B2(n9119), .A(n9118), .ZN(P2_U3446) );
  INV_X1 U10189 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9122) );
  MUX2_X1 U10190 ( .A(n9122), .B(n9121), .S(n10727), .Z(n9125) );
  NAND2_X1 U10191 ( .A1(n9123), .A2(n9141), .ZN(n9124) );
  OAI211_X1 U10192 ( .C1(n9126), .C2(n9145), .A(n9125), .B(n9124), .ZN(
        P2_U3444) );
  INV_X1 U10193 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9127) );
  MUX2_X1 U10194 ( .A(n9128), .B(n9127), .S(n10724), .Z(n9131) );
  NAND2_X1 U10195 ( .A1(n9129), .A2(n9141), .ZN(n9130) );
  OAI211_X1 U10196 ( .C1(n9132), .C2(n9145), .A(n9131), .B(n9130), .ZN(
        P2_U3441) );
  INV_X1 U10197 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9133) );
  MUX2_X1 U10198 ( .A(n9134), .B(n9133), .S(n10724), .Z(n9137) );
  NAND2_X1 U10199 ( .A1(n9135), .A2(n9141), .ZN(n9136) );
  OAI211_X1 U10200 ( .C1(n9138), .C2(n9145), .A(n9137), .B(n9136), .ZN(
        P2_U3438) );
  INV_X1 U10201 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9139) );
  MUX2_X1 U10202 ( .A(n9140), .B(n9139), .S(n10724), .Z(n9144) );
  NAND2_X1 U10203 ( .A1(n9142), .A2(n9141), .ZN(n9143) );
  OAI211_X1 U10204 ( .C1(n9146), .C2(n9145), .A(n9144), .B(n9143), .ZN(
        P2_U3435) );
  INV_X1 U10205 ( .A(n10050), .ZN(n9152) );
  NOR4_X1 U10206 ( .A1(n9148), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n9147), .ZN(n9149) );
  AOI21_X1 U10207 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n9150), .A(n9149), .ZN(
        n9151) );
  OAI21_X1 U10208 ( .B1(n9152), .B2(n9159), .A(n9151), .ZN(P2_U3264) );
  INV_X1 U10209 ( .A(n9289), .ZN(n10277) );
  OAI222_X1 U10210 ( .A1(n9159), .A2(n10277), .B1(n9156), .B2(n9155), .C1(
        P2_U3151), .C2(n9153), .ZN(P2_U3266) );
  INV_X1 U10211 ( .A(n9157), .ZN(n10286) );
  OAI222_X1 U10212 ( .A1(n9156), .A2(n9160), .B1(n9159), .B2(n10286), .C1(
        n9158), .C2(P2_U3151), .ZN(P2_U3269) );
  MUX2_X1 U10213 ( .A(n9161), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10214 ( .A1(n9162), .A2(n9163), .ZN(n9164) );
  XOR2_X1 U10215 ( .A(n9165), .B(n9164), .Z(n9173) );
  OAI21_X1 U10216 ( .B1(n9278), .B2(n9167), .A(n9166), .ZN(n9170) );
  OAI22_X1 U10217 ( .A1(n9276), .A2(n9879), .B1(n9275), .B2(n9168), .ZN(n9169)
         );
  AOI211_X1 U10218 ( .C1(n9171), .C2(n9281), .A(n9170), .B(n9169), .ZN(n9172)
         );
  OAI21_X1 U10219 ( .B1(n9173), .B2(n9284), .A(n9172), .ZN(P1_U3215) );
  AOI21_X1 U10220 ( .B1(n9176), .B2(n9174), .A(n9175), .ZN(n9177) );
  OAI21_X1 U10221 ( .B1(n9223), .B2(n9177), .A(n9259), .ZN(n9181) );
  NOR2_X1 U10222 ( .A1(n9276), .A2(n9729), .ZN(n9179) );
  OAI22_X1 U10223 ( .A1(n9638), .A2(n9278), .B1(n9765), .B2(n9275), .ZN(n9178)
         );
  AOI211_X1 U10224 ( .C1(P1_REG3_REG_23__SCAN_IN), .C2(P1_U3086), .A(n9179), 
        .B(n9178), .ZN(n9180) );
  OAI211_X1 U10225 ( .C1(n10019), .C2(n9242), .A(n9181), .B(n9180), .ZN(
        P1_U3216) );
  AOI21_X1 U10226 ( .B1(n9183), .B2(n9182), .A(n4940), .ZN(n9187) );
  NAND2_X1 U10227 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9606) );
  OAI21_X1 U10228 ( .B1(n9276), .B2(n9949), .A(n9606), .ZN(n9185) );
  OAI22_X1 U10229 ( .A1(n9278), .A2(n9822), .B1(n9275), .B2(n9828), .ZN(n9184)
         );
  AOI211_X1 U10230 ( .C1(n9962), .C2(n9281), .A(n9185), .B(n9184), .ZN(n9186)
         );
  OAI21_X1 U10231 ( .B1(n9187), .B2(n9284), .A(n9186), .ZN(P1_U3219) );
  OAI21_X1 U10232 ( .B1(n9190), .B2(n9189), .A(n9188), .ZN(n9191) );
  NAND2_X1 U10233 ( .A1(n9191), .A2(n9259), .ZN(n9195) );
  NOR2_X1 U10234 ( .A1(n9278), .A2(n9949), .ZN(n9193) );
  OAI22_X1 U10235 ( .A1(n9638), .A2(n9276), .B1(n9275), .B2(n9795), .ZN(n9192)
         );
  AOI211_X1 U10236 ( .C1(P1_REG3_REG_21__SCAN_IN), .C2(P1_U3086), .A(n9193), 
        .B(n9192), .ZN(n9194) );
  OAI211_X1 U10237 ( .C1(n5236), .C2(n9242), .A(n9195), .B(n9194), .ZN(
        P1_U3223) );
  OAI21_X1 U10238 ( .B1(n9198), .B2(n9197), .A(n9196), .ZN(n9199) );
  NAND2_X1 U10239 ( .A1(n9199), .A2(n9259), .ZN(n9203) );
  NOR2_X1 U10240 ( .A1(n9276), .A2(n9730), .ZN(n9201) );
  OAI22_X1 U10241 ( .A1(n9278), .A2(n9729), .B1(n9275), .B2(n9736), .ZN(n9200)
         );
  AOI211_X1 U10242 ( .C1(P1_REG3_REG_25__SCAN_IN), .C2(P1_U3086), .A(n9201), 
        .B(n9200), .ZN(n9202) );
  OAI211_X1 U10243 ( .C1(n10014), .C2(n9242), .A(n9203), .B(n9202), .ZN(
        P1_U3225) );
  AOI21_X1 U10244 ( .B1(n9206), .B2(n9205), .A(n9204), .ZN(n9211) );
  OAI21_X1 U10245 ( .B1(n9276), .B2(n9968), .A(n9207), .ZN(n9209) );
  OAI22_X1 U10246 ( .A1(n9278), .A2(n9879), .B1(n9275), .B2(n9881), .ZN(n9208)
         );
  AOI211_X1 U10247 ( .C1(n9982), .C2(n9281), .A(n9209), .B(n9208), .ZN(n9210)
         );
  OAI21_X1 U10248 ( .B1(n9211), .B2(n9284), .A(n9210), .ZN(P1_U3226) );
  XNOR2_X1 U10249 ( .A(n9213), .B(n9212), .ZN(n9214) );
  XNOR2_X1 U10250 ( .A(n9215), .B(n9214), .ZN(n9219) );
  NAND2_X1 U10251 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9562) );
  OAI21_X1 U10252 ( .B1(n9276), .B2(n9822), .A(n9562), .ZN(n9217) );
  OAI22_X1 U10253 ( .A1(n9278), .A2(n9975), .B1(n9275), .B2(n9856), .ZN(n9216)
         );
  AOI211_X1 U10254 ( .C1(n9868), .C2(n9281), .A(n9217), .B(n9216), .ZN(n9218)
         );
  OAI21_X1 U10255 ( .B1(n9219), .B2(n9284), .A(n9218), .ZN(P1_U3228) );
  INV_X1 U10256 ( .A(n9220), .ZN(n9225) );
  NOR3_X1 U10257 ( .A1(n9223), .A2(n9222), .A3(n9221), .ZN(n9224) );
  OAI21_X1 U10258 ( .B1(n9225), .B2(n9224), .A(n9259), .ZN(n9230) );
  OAI22_X1 U10259 ( .A1(n9276), .A2(n9921), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9226), .ZN(n9228) );
  INV_X1 U10260 ( .A(n9639), .ZN(n9779) );
  OAI22_X1 U10261 ( .A1(n9779), .A2(n9278), .B1(n9747), .B2(n9275), .ZN(n9227)
         );
  AOI211_X1 U10262 ( .C1(n9933), .C2(n9281), .A(n9228), .B(n9227), .ZN(n9229)
         );
  NAND2_X1 U10263 ( .A1(n9230), .A2(n9229), .ZN(P1_U3229) );
  INV_X1 U10264 ( .A(n9231), .ZN(n9235) );
  NOR3_X1 U10265 ( .A1(n4940), .A2(n9233), .A3(n9232), .ZN(n9234) );
  OAI21_X1 U10266 ( .B1(n9235), .B2(n9234), .A(n9259), .ZN(n9241) );
  INV_X1 U10267 ( .A(n9836), .ZN(n9324) );
  NOR2_X1 U10268 ( .A1(n9278), .A2(n9324), .ZN(n9238) );
  OAI22_X1 U10269 ( .A1(n9276), .A2(n9778), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9236), .ZN(n9237) );
  AOI211_X1 U10270 ( .C1(n9239), .C2(n9814), .A(n9238), .B(n9237), .ZN(n9240)
         );
  OAI211_X1 U10271 ( .C1(n9614), .C2(n9242), .A(n9241), .B(n9240), .ZN(
        P1_U3233) );
  NAND2_X1 U10272 ( .A1(n9174), .A2(n9243), .ZN(n9244) );
  XOR2_X1 U10273 ( .A(n9245), .B(n9244), .Z(n9250) );
  INV_X1 U10274 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9246) );
  OAI22_X1 U10275 ( .A1(n9278), .A2(n9778), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9246), .ZN(n9248) );
  OAI22_X1 U10276 ( .A1(n9779), .A2(n9276), .B1(n9275), .B2(n9782), .ZN(n9247)
         );
  AOI211_X1 U10277 ( .C1(n9944), .C2(n9281), .A(n9248), .B(n9247), .ZN(n9249)
         );
  OAI21_X1 U10278 ( .B1(n9250), .B2(n9284), .A(n9249), .ZN(P1_U3235) );
  XNOR2_X1 U10279 ( .A(n9252), .B(n9251), .ZN(n9253) );
  XNOR2_X1 U10280 ( .A(n9254), .B(n9253), .ZN(n9258) );
  NAND2_X1 U10281 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9585) );
  OAI21_X1 U10282 ( .B1(n9276), .B2(n9324), .A(n9585), .ZN(n9256) );
  OAI22_X1 U10283 ( .A1(n9278), .A2(n9968), .B1(n9275), .B2(n9841), .ZN(n9255)
         );
  AOI211_X1 U10284 ( .C1(n9847), .C2(n9281), .A(n9256), .B(n9255), .ZN(n9257)
         );
  OAI21_X1 U10285 ( .B1(n9258), .B2(n9284), .A(n9257), .ZN(P1_U3238) );
  NAND2_X1 U10286 ( .A1(n9260), .A2(n9259), .ZN(n9268) );
  AOI21_X1 U10287 ( .B1(n9196), .B2(n9262), .A(n9261), .ZN(n9267) );
  INV_X1 U10288 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9263) );
  OAI22_X1 U10289 ( .A1(n9278), .A2(n9921), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9263), .ZN(n9265) );
  OAI22_X1 U10290 ( .A1(n9276), .A2(n9911), .B1(n9275), .B2(n9717), .ZN(n9264)
         );
  OAI21_X1 U10291 ( .B1(n9268), .B2(n9267), .A(n9266), .ZN(P1_U3240) );
  INV_X1 U10292 ( .A(n9269), .ZN(n9271) );
  NAND2_X1 U10293 ( .A1(n9271), .A2(n9270), .ZN(n9273) );
  XNOR2_X1 U10294 ( .A(n9273), .B(n9272), .ZN(n9285) );
  OAI22_X1 U10295 ( .A1(n9276), .A2(n9975), .B1(n9275), .B2(n9274), .ZN(n9280)
         );
  OAI21_X1 U10296 ( .B1(n9278), .B2(n9987), .A(n9277), .ZN(n9279) );
  NOR2_X1 U10297 ( .A1(n9280), .A2(n9279), .ZN(n9283) );
  NAND2_X1 U10298 ( .A1(n9632), .A2(n9281), .ZN(n9282) );
  OAI211_X1 U10299 ( .C1(n9285), .C2(n9284), .A(n9283), .B(n9282), .ZN(
        P1_U3241) );
  NOR2_X1 U10300 ( .A1(n9287), .A2(n9286), .ZN(n9552) );
  OAI21_X1 U10301 ( .B1(n9339), .B2(n6319), .A(P1_B_REG_SCAN_IN), .ZN(n9551)
         );
  NAND2_X1 U10302 ( .A1(n9289), .A2(n9335), .ZN(n9291) );
  OR2_X1 U10303 ( .A1(n9296), .A2(n10278), .ZN(n9290) );
  OR2_X1 U10304 ( .A1(n9630), .A2(n9902), .ZN(n9512) );
  AND2_X1 U10305 ( .A1(n9516), .A2(n9512), .ZN(n9294) );
  NAND2_X1 U10306 ( .A1(n9630), .A2(n9902), .ZN(n9662) );
  NAND2_X1 U10307 ( .A1(n9693), .A2(n9911), .ZN(n9354) );
  NAND2_X1 U10308 ( .A1(n9662), .A2(n9354), .ZN(n9389) );
  NAND2_X1 U10309 ( .A1(n9904), .A2(n9682), .ZN(n9517) );
  INV_X1 U10310 ( .A(n9517), .ZN(n9293) );
  NAND2_X1 U10311 ( .A1(n9735), .A2(n9921), .ZN(n9658) );
  NAND3_X1 U10312 ( .A1(n9294), .A2(n9661), .A3(n9504), .ZN(n9327) );
  AOI21_X1 U10313 ( .B1(n9660), .B2(n9658), .A(n9327), .ZN(n9292) );
  AOI211_X1 U10314 ( .C1(n9294), .C2(n9389), .A(n9293), .B(n9292), .ZN(n9347)
         );
  INV_X1 U10315 ( .A(n9666), .ZN(n9333) );
  NAND2_X1 U10316 ( .A1(n10055), .A2(n9335), .ZN(n9298) );
  OR2_X1 U10317 ( .A1(n9296), .A2(n9295), .ZN(n9297) );
  NAND2_X1 U10318 ( .A1(n9800), .A2(n9778), .ZN(n9492) );
  NAND2_X1 U10319 ( .A1(n9813), .A2(n9949), .ZN(n9789) );
  NAND2_X1 U10320 ( .A1(n9492), .A2(n9789), .ZN(n9299) );
  NAND2_X1 U10321 ( .A1(n9764), .A2(n9779), .ZN(n9656) );
  NAND2_X1 U10322 ( .A1(n9944), .A2(n9638), .ZN(n9655) );
  NAND2_X1 U10323 ( .A1(n9656), .A2(n9655), .ZN(n9496) );
  NAND2_X1 U10324 ( .A1(n9933), .A2(n9729), .ZN(n9390) );
  INV_X1 U10325 ( .A(n9390), .ZN(n9330) );
  AOI211_X1 U10326 ( .C1(n9653), .C2(n9299), .A(n9496), .B(n9330), .ZN(n9346)
         );
  OR2_X1 U10327 ( .A1(n9813), .A2(n9949), .ZN(n9488) );
  OR2_X1 U10328 ( .A1(n9962), .A2(n9324), .ZN(n9485) );
  NOR2_X1 U10329 ( .A1(n9847), .A2(n9822), .ZN(n9477) );
  NAND2_X1 U10330 ( .A1(n9847), .A2(n9822), .ZN(n9478) );
  NAND2_X1 U10331 ( .A1(n9868), .A2(n9968), .ZN(n9343) );
  AND2_X1 U10332 ( .A1(n9478), .A2(n9343), .ZN(n9474) );
  AND2_X1 U10333 ( .A1(n9464), .A2(n9300), .ZN(n9458) );
  AOI21_X1 U10334 ( .B1(n5664), .B2(n10539), .A(n9521), .ZN(n9301) );
  NAND2_X1 U10335 ( .A1(n6474), .A2(n5611), .ZN(n9361) );
  AND2_X1 U10336 ( .A1(n9301), .A2(n9361), .ZN(n9303) );
  OAI211_X1 U10337 ( .C1(n9304), .C2(n9303), .A(n9302), .B(n9395), .ZN(n9308)
         );
  INV_X1 U10338 ( .A(n9305), .ZN(n9307) );
  AND2_X1 U10339 ( .A1(n9307), .A2(n9306), .ZN(n9401) );
  OAI211_X1 U10340 ( .C1(n9310), .C2(n9309), .A(n9308), .B(n9401), .ZN(n9312)
         );
  INV_X1 U10341 ( .A(n9409), .ZN(n9311) );
  AOI21_X1 U10342 ( .B1(n9312), .B2(n9403), .A(n9311), .ZN(n9315) );
  INV_X1 U10343 ( .A(n9373), .ZN(n9314) );
  OAI21_X1 U10344 ( .B1(n9315), .B2(n9314), .A(n9313), .ZN(n9316) );
  NAND2_X1 U10345 ( .A1(n9439), .A2(n9427), .ZN(n9433) );
  AOI21_X1 U10346 ( .B1(n9316), .B2(n9431), .A(n9433), .ZN(n9317) );
  NAND2_X1 U10347 ( .A1(n9453), .A2(n9436), .ZN(n9441) );
  AND2_X1 U10348 ( .A1(n9456), .A2(n9440), .ZN(n9448) );
  OAI21_X1 U10349 ( .B1(n9317), .B2(n9441), .A(n9448), .ZN(n9318) );
  NAND3_X1 U10350 ( .A1(n9460), .A2(n9318), .A3(n9454), .ZN(n9320) );
  INV_X1 U10351 ( .A(n9468), .ZN(n9319) );
  AOI21_X1 U10352 ( .B1(n9458), .B2(n9320), .A(n9319), .ZN(n9321) );
  NAND2_X1 U10353 ( .A1(n9982), .A2(n9975), .ZN(n9466) );
  OR2_X1 U10354 ( .A1(n9982), .A2(n9975), .ZN(n9469) );
  OAI211_X1 U10355 ( .C1(n9321), .C2(n5119), .A(n9475), .B(n9469), .ZN(n9322)
         );
  NAND2_X1 U10356 ( .A1(n9474), .A2(n9322), .ZN(n9323) );
  NAND3_X1 U10357 ( .A1(n9485), .A2(n5153), .A3(n9323), .ZN(n9325) );
  NAND2_X1 U10358 ( .A1(n9962), .A2(n9324), .ZN(n9484) );
  NAND2_X1 U10359 ( .A1(n9325), .A2(n9484), .ZN(n9326) );
  NAND3_X1 U10360 ( .A1(n9653), .A2(n9488), .A3(n9326), .ZN(n9331) );
  OR2_X1 U10361 ( .A1(n9764), .A2(n9779), .ZN(n9497) );
  OR2_X1 U10362 ( .A1(n9944), .A2(n9638), .ZN(n9355) );
  NAND2_X1 U10363 ( .A1(n9497), .A2(n9355), .ZN(n9495) );
  OR2_X1 U10364 ( .A1(n9933), .A2(n9729), .ZN(n9657) );
  INV_X1 U10365 ( .A(n9657), .ZN(n9391) );
  AOI21_X1 U10366 ( .B1(n9656), .B2(n9495), .A(n9391), .ZN(n9329) );
  INV_X1 U10367 ( .A(n9327), .ZN(n9328) );
  OR2_X1 U10368 ( .A1(n9735), .A2(n9921), .ZN(n9659) );
  OAI211_X1 U10369 ( .C1(n9330), .C2(n9329), .A(n9328), .B(n9659), .ZN(n9344)
         );
  AOI21_X1 U10370 ( .B1(n9346), .B2(n9331), .A(n9344), .ZN(n9332) );
  AOI21_X1 U10371 ( .B1(n9333), .B2(n9628), .A(n9332), .ZN(n9334) );
  NOR2_X1 U10372 ( .A1(n9628), .A2(n9333), .ZN(n9348) );
  AOI21_X1 U10373 ( .B1(n9347), .B2(n9334), .A(n9348), .ZN(n9338) );
  NAND2_X1 U10374 ( .A1(n10050), .A2(n9335), .ZN(n9337) );
  INV_X1 U10375 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10047) );
  OR2_X1 U10376 ( .A1(n9296), .A2(n10047), .ZN(n9336) );
  NOR2_X1 U10377 ( .A1(n9621), .A2(n9620), .ZN(n9520) );
  NAND2_X1 U10378 ( .A1(n9621), .A2(n9620), .ZN(n9538) );
  OAI21_X1 U10379 ( .B1(n9338), .B2(n9520), .A(n9538), .ZN(n9549) );
  AOI21_X1 U10380 ( .B1(n9549), .B2(n9340), .A(n9339), .ZN(n9548) );
  INV_X1 U10381 ( .A(n9872), .ZN(n9877) );
  NAND2_X1 U10382 ( .A1(n9475), .A2(n9343), .ZN(n9636) );
  XNOR2_X1 U10383 ( .A(n9847), .B(n9851), .ZN(n9840) );
  NAND3_X1 U10384 ( .A1(n9806), .A2(n9653), .A3(n9488), .ZN(n9345) );
  AOI21_X1 U10385 ( .B1(n9346), .B2(n9345), .A(n9344), .ZN(n9351) );
  INV_X1 U10386 ( .A(n9347), .ZN(n9350) );
  INV_X1 U10387 ( .A(n9348), .ZN(n9349) );
  OAI21_X1 U10388 ( .B1(n9351), .B2(n9350), .A(n9523), .ZN(n9353) );
  NAND2_X1 U10389 ( .A1(n9666), .A2(n9525), .ZN(n9352) );
  NAND2_X1 U10390 ( .A1(n9628), .A2(n9352), .ZN(n9524) );
  INV_X1 U10391 ( .A(n9538), .ZN(n9386) );
  AOI211_X1 U10392 ( .C1(n9353), .C2(n9524), .A(n9386), .B(n9522), .ZN(n9387)
         );
  XOR2_X1 U10393 ( .A(n9666), .B(n9628), .Z(n9385) );
  NAND2_X1 U10394 ( .A1(n9512), .A2(n9662), .ZN(n9679) );
  NAND2_X1 U10395 ( .A1(n9504), .A2(n9660), .ZN(n9716) );
  NAND2_X1 U10396 ( .A1(n9657), .A2(n9390), .ZN(n9751) );
  NAND2_X1 U10397 ( .A1(n9659), .A2(n9658), .ZN(n9731) );
  NAND2_X1 U10398 ( .A1(n9355), .A2(n9655), .ZN(n9776) );
  INV_X1 U10399 ( .A(n9776), .ZN(n9771) );
  NAND2_X1 U10400 ( .A1(n9488), .A2(n9789), .ZN(n9803) );
  INV_X1 U10401 ( .A(n9803), .ZN(n9807) );
  INV_X1 U10402 ( .A(n9407), .ZN(n9359) );
  INV_X1 U10403 ( .A(n9356), .ZN(n9357) );
  NAND4_X1 U10404 ( .A1(n9360), .A2(n9359), .A3(n9358), .A4(n9357), .ZN(n9365)
         );
  INV_X1 U10405 ( .A(n9361), .ZN(n9362) );
  NOR2_X1 U10406 ( .A1(n9363), .A2(n9362), .ZN(n10527) );
  NAND3_X1 U10407 ( .A1(n10527), .A2(n9521), .A3(n9409), .ZN(n9364) );
  NOR2_X1 U10408 ( .A1(n9365), .A2(n9364), .ZN(n9368) );
  NAND4_X1 U10409 ( .A1(n9368), .A2(n9367), .A3(n9429), .A4(n9366), .ZN(n9369)
         );
  NOR2_X1 U10410 ( .A1(n9370), .A2(n9369), .ZN(n9371) );
  NAND4_X1 U10411 ( .A1(n9374), .A2(n9373), .A3(n9372), .A4(n9371), .ZN(n9376)
         );
  NOR2_X1 U10412 ( .A1(n9376), .A2(n9375), .ZN(n9377) );
  NAND4_X1 U10413 ( .A1(n9872), .A2(n9378), .A3(n9451), .A4(n9377), .ZN(n9379)
         );
  NOR2_X1 U10414 ( .A1(n9636), .A2(n9379), .ZN(n9380) );
  AND4_X1 U10415 ( .A1(n9793), .A2(n9823), .A3(n9380), .A4(n9840), .ZN(n9381)
         );
  NAND4_X1 U10416 ( .A1(n9760), .A2(n9771), .A3(n9807), .A4(n9381), .ZN(n9382)
         );
  OR4_X1 U10417 ( .A1(n9716), .A2(n9751), .A3(n9731), .A4(n9382), .ZN(n9383)
         );
  OAI21_X1 U10418 ( .B1(n9387), .B2(n9532), .A(n5608), .ZN(n9546) );
  NAND3_X1 U10419 ( .A1(n9538), .A2(n9526), .A3(n9523), .ZN(n9543) );
  OAI21_X1 U10420 ( .B1(n9511), .B2(n9661), .A(n9512), .ZN(n9388) );
  AOI21_X1 U10421 ( .B1(n9511), .B2(n9389), .A(n9388), .ZN(n9510) );
  INV_X1 U10422 ( .A(n9511), .ZN(n9515) );
  AND2_X1 U10423 ( .A1(n9658), .A2(n9390), .ZN(n9393) );
  NOR2_X1 U10424 ( .A1(n9731), .A2(n9391), .ZN(n9392) );
  MUX2_X1 U10425 ( .A(n9393), .B(n9392), .S(n9511), .Z(n9501) );
  OAI211_X1 U10426 ( .C1(n9397), .C2(n9396), .A(n9395), .B(n9394), .ZN(n9399)
         );
  MUX2_X1 U10427 ( .A(n9399), .B(n9398), .S(n9511), .Z(n9408) );
  INV_X1 U10428 ( .A(n9400), .ZN(n9406) );
  INV_X1 U10429 ( .A(n9401), .ZN(n9402) );
  NAND2_X1 U10430 ( .A1(n9402), .A2(n9403), .ZN(n9404) );
  MUX2_X1 U10431 ( .A(n9404), .B(n9403), .S(n9511), .Z(n9405) );
  OAI211_X1 U10432 ( .C1(n9408), .C2(n9407), .A(n9406), .B(n9405), .ZN(n9413)
         );
  MUX2_X1 U10433 ( .A(n9410), .B(n9409), .S(n9511), .Z(n9411) );
  NAND3_X1 U10434 ( .A1(n9413), .A2(n9412), .A3(n9411), .ZN(n9422) );
  INV_X1 U10435 ( .A(n9431), .ZN(n9414) );
  AOI21_X1 U10436 ( .B1(n9422), .B2(n9415), .A(n9414), .ZN(n9424) );
  INV_X1 U10437 ( .A(n9416), .ZN(n9417) );
  NOR2_X1 U10438 ( .A1(n9418), .A2(n9417), .ZN(n9421) );
  NAND3_X1 U10439 ( .A1(n9427), .A2(n9429), .A3(n9419), .ZN(n9420) );
  AOI21_X1 U10440 ( .B1(n9422), .B2(n9421), .A(n9420), .ZN(n9423) );
  MUX2_X1 U10441 ( .A(n9424), .B(n9423), .S(n9511), .Z(n9425) );
  NAND2_X1 U10442 ( .A1(n9425), .A2(n9426), .ZN(n9438) );
  NAND2_X1 U10443 ( .A1(n9431), .A2(n9426), .ZN(n9428) );
  NAND2_X1 U10444 ( .A1(n9428), .A2(n9427), .ZN(n9435) );
  INV_X1 U10445 ( .A(n9429), .ZN(n9430) );
  AND2_X1 U10446 ( .A1(n9431), .A2(n9430), .ZN(n9432) );
  NOR2_X1 U10447 ( .A1(n9433), .A2(n9432), .ZN(n9434) );
  MUX2_X1 U10448 ( .A(n9435), .B(n9434), .S(n9515), .Z(n9443) );
  AND2_X1 U10449 ( .A1(n9443), .A2(n9436), .ZN(n9437) );
  NAND2_X1 U10450 ( .A1(n9438), .A2(n9437), .ZN(n9447) );
  AND2_X1 U10451 ( .A1(n9440), .A2(n9439), .ZN(n9445) );
  AOI21_X1 U10452 ( .B1(n9443), .B2(n9442), .A(n9441), .ZN(n9444) );
  MUX2_X1 U10453 ( .A(n9445), .B(n9444), .S(n9515), .Z(n9446) );
  NAND2_X1 U10454 ( .A1(n9447), .A2(n9446), .ZN(n9455) );
  NAND2_X1 U10455 ( .A1(n9455), .A2(n9448), .ZN(n9449) );
  NAND2_X1 U10456 ( .A1(n9449), .A2(n9454), .ZN(n9452) );
  NAND2_X1 U10457 ( .A1(n9468), .A2(n9460), .ZN(n9450) );
  AOI21_X1 U10458 ( .B1(n9452), .B2(n9451), .A(n9450), .ZN(n9463) );
  NAND3_X1 U10459 ( .A1(n9455), .A2(n9454), .A3(n9453), .ZN(n9457) );
  NAND2_X1 U10460 ( .A1(n9457), .A2(n9456), .ZN(n9461) );
  INV_X1 U10461 ( .A(n9458), .ZN(n9459) );
  AOI21_X1 U10462 ( .B1(n9461), .B2(n9460), .A(n9459), .ZN(n9462) );
  MUX2_X1 U10463 ( .A(n9463), .B(n9462), .S(n9511), .Z(n9467) );
  INV_X1 U10464 ( .A(n9464), .ZN(n9465) );
  INV_X1 U10465 ( .A(n9467), .ZN(n9471) );
  AND2_X1 U10466 ( .A1(n9469), .A2(n9468), .ZN(n9470) );
  AOI21_X1 U10467 ( .B1(n9471), .B2(n9470), .A(n5119), .ZN(n9472) );
  NAND2_X1 U10468 ( .A1(n9823), .A2(n5153), .ZN(n9473) );
  AOI21_X1 U10469 ( .B1(n9481), .B2(n9474), .A(n9473), .ZN(n9483) );
  INV_X1 U10470 ( .A(n9475), .ZN(n9476) );
  NOR2_X1 U10471 ( .A1(n9477), .A2(n9476), .ZN(n9480) );
  NAND2_X1 U10472 ( .A1(n9484), .A2(n9478), .ZN(n9479) );
  AOI21_X1 U10473 ( .B1(n9481), .B2(n9480), .A(n9479), .ZN(n9482) );
  MUX2_X1 U10474 ( .A(n9483), .B(n9482), .S(n9511), .Z(n9491) );
  NAND2_X1 U10475 ( .A1(n9789), .A2(n9484), .ZN(n9487) );
  NAND2_X1 U10476 ( .A1(n9488), .A2(n9485), .ZN(n9486) );
  MUX2_X1 U10477 ( .A(n9487), .B(n9486), .S(n9511), .Z(n9490) );
  MUX2_X1 U10478 ( .A(n9488), .B(n9789), .S(n9511), .Z(n9489) );
  OAI211_X1 U10479 ( .C1(n9491), .C2(n9490), .A(n9793), .B(n9489), .ZN(n9494)
         );
  MUX2_X1 U10480 ( .A(n9492), .B(n9653), .S(n9511), .Z(n9493) );
  AOI21_X1 U10481 ( .B1(n9494), .B2(n9493), .A(n9776), .ZN(n9500) );
  MUX2_X1 U10482 ( .A(n9496), .B(n9495), .S(n9511), .Z(n9499) );
  INV_X1 U10483 ( .A(n9751), .ZN(n9743) );
  MUX2_X1 U10484 ( .A(n9656), .B(n9497), .S(n9515), .Z(n9498) );
  OR2_X1 U10485 ( .A1(n9659), .A2(n9511), .ZN(n9502) );
  NAND2_X1 U10486 ( .A1(n9503), .A2(n9515), .ZN(n9505) );
  INV_X1 U10487 ( .A(n9506), .ZN(n9508) );
  NOR2_X1 U10488 ( .A1(n9716), .A2(n5145), .ZN(n9507) );
  AOI21_X1 U10489 ( .B1(n9508), .B2(n9507), .A(n9698), .ZN(n9509) );
  MUX2_X1 U10490 ( .A(n9662), .B(n9512), .S(n9511), .Z(n9513) );
  INV_X1 U10491 ( .A(n9513), .ZN(n9514) );
  MUX2_X1 U10492 ( .A(n9517), .B(n9516), .S(n9515), .Z(n9518) );
  NAND3_X1 U10493 ( .A1(n9519), .A2(n9524), .A3(n9518), .ZN(n9542) );
  INV_X1 U10494 ( .A(n9520), .ZN(n9537) );
  NOR3_X1 U10495 ( .A1(n9537), .A2(n9521), .A3(n5608), .ZN(n9531) );
  NOR3_X1 U10496 ( .A1(n9621), .A2(n9522), .A3(n9524), .ZN(n9530) );
  INV_X1 U10497 ( .A(n9523), .ZN(n9534) );
  OAI211_X1 U10498 ( .C1(n9534), .C2(n9620), .A(n5608), .B(n9621), .ZN(n9528)
         );
  INV_X1 U10499 ( .A(n9524), .ZN(n9536) );
  NAND3_X1 U10500 ( .A1(n9536), .A2(n9526), .A3(n9525), .ZN(n9527) );
  OAI211_X1 U10501 ( .C1(n9610), .C2(n5609), .A(n9528), .B(n9527), .ZN(n9529)
         );
  NOR4_X1 U10502 ( .A1(n9532), .A2(n9531), .A3(n9530), .A4(n9529), .ZN(n9541)
         );
  AOI21_X1 U10503 ( .B1(n9533), .B2(n5609), .A(n5608), .ZN(n9535) );
  AOI211_X1 U10504 ( .C1(n9536), .C2(n5608), .A(n9535), .B(n9534), .ZN(n9539)
         );
  NAND4_X1 U10505 ( .A1(n9539), .A2(n9542), .A3(n9538), .A4(n9537), .ZN(n9540)
         );
  OAI211_X1 U10506 ( .C1(n9543), .C2(n9542), .A(n9541), .B(n9540), .ZN(n9545)
         );
  NAND3_X1 U10507 ( .A1(n9546), .A2(n9545), .A3(n9544), .ZN(n9547) );
  OAI211_X1 U10508 ( .C1(n9288), .C2(n9549), .A(n9548), .B(n9547), .ZN(n9550)
         );
  OAI21_X1 U10509 ( .B1(n9552), .B2(n9551), .A(n9550), .ZN(P1_U3242) );
  INV_X1 U10510 ( .A(n9902), .ZN(n9703) );
  MUX2_X1 U10511 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9703), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10512 ( .A(n9712), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9561), .Z(
        P1_U3581) );
  MUX2_X1 U10513 ( .A(n9702), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9561), .Z(
        P1_U3580) );
  MUX2_X1 U10514 ( .A(n9642), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9561), .Z(
        P1_U3579) );
  MUX2_X1 U10515 ( .A(n9758), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9561), .Z(
        P1_U3578) );
  MUX2_X1 U10516 ( .A(n9791), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9561), .Z(
        P1_U3576) );
  MUX2_X1 U10517 ( .A(n9809), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9561), .Z(
        P1_U3575) );
  MUX2_X1 U10518 ( .A(n9553), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9561), .Z(
        P1_U3574) );
  MUX2_X1 U10519 ( .A(n9836), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9561), .Z(
        P1_U3573) );
  MUX2_X1 U10520 ( .A(n9635), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9561), .Z(
        P1_U3571) );
  MUX2_X1 U10521 ( .A(n9554), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9561), .Z(
        P1_U3570) );
  MUX2_X1 U10522 ( .A(n9631), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9561), .Z(
        P1_U3569) );
  MUX2_X1 U10523 ( .A(n9555), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9561), .Z(
        P1_U3568) );
  MUX2_X1 U10524 ( .A(n9556), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9561), .Z(
        P1_U3566) );
  MUX2_X1 U10525 ( .A(n10703), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9561), .Z(
        P1_U3565) );
  MUX2_X1 U10526 ( .A(n9557), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9561), .Z(
        P1_U3564) );
  MUX2_X1 U10527 ( .A(n10679), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9561), .Z(
        P1_U3563) );
  MUX2_X1 U10528 ( .A(n10661), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9561), .Z(
        P1_U3562) );
  MUX2_X1 U10529 ( .A(n9558), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9561), .Z(
        P1_U3561) );
  MUX2_X1 U10530 ( .A(n9559), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9561), .Z(
        P1_U3560) );
  MUX2_X1 U10531 ( .A(n9560), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9561), .Z(
        P1_U3558) );
  MUX2_X1 U10532 ( .A(n10598), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9561), .Z(
        P1_U3557) );
  INV_X1 U10533 ( .A(n9562), .ZN(n9569) );
  XNOR2_X1 U10534 ( .A(n9587), .B(n9565), .ZN(n9566) );
  NAND2_X1 U10535 ( .A1(n9567), .A2(n9566), .ZN(n9586) );
  AOI221_X1 U10536 ( .B1(n9567), .B2(n9586), .C1(n9566), .C2(n9586), .A(n9590), 
        .ZN(n9568) );
  AOI211_X1 U10537 ( .C1(n10350), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n9569), .B(
        n9568), .ZN(n9577) );
  XNOR2_X1 U10538 ( .A(n9587), .B(n9978), .ZN(n9574) );
  INV_X1 U10539 ( .A(n9570), .ZN(n9571) );
  NAND2_X1 U10540 ( .A1(n9572), .A2(n9571), .ZN(n9573) );
  NAND2_X1 U10541 ( .A1(n9573), .A2(n9574), .ZN(n9581) );
  OAI21_X1 U10542 ( .B1(n9574), .B2(n9573), .A(n9581), .ZN(n9575) );
  NAND2_X1 U10543 ( .A1(n9582), .A2(n9575), .ZN(n9576) );
  OAI211_X1 U10544 ( .C1(n10360), .C2(n9578), .A(n9577), .B(n9576), .ZN(
        P1_U3260) );
  INV_X1 U10545 ( .A(n9602), .ZN(n9596) );
  INV_X1 U10546 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9971) );
  XNOR2_X1 U10547 ( .A(n9602), .B(n9971), .ZN(n9584) );
  OR2_X1 U10548 ( .A1(n9587), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9579) );
  AND2_X1 U10549 ( .A1(n9581), .A2(n9579), .ZN(n9583) );
  AND2_X1 U10550 ( .A1(n9584), .A2(n9579), .ZN(n9580) );
  NAND2_X1 U10551 ( .A1(n9581), .A2(n9580), .ZN(n9598) );
  OAI211_X1 U10552 ( .C1(n9584), .C2(n9583), .A(n9582), .B(n9598), .ZN(n9595)
         );
  INV_X1 U10553 ( .A(n9585), .ZN(n9594) );
  OAI21_X1 U10554 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n9587), .A(n9586), .ZN(
        n9592) );
  NOR2_X1 U10555 ( .A1(n9602), .A2(n9588), .ZN(n9589) );
  AOI21_X1 U10556 ( .B1(n9602), .B2(n9588), .A(n9589), .ZN(n9591) );
  AOI211_X1 U10557 ( .C1(n9592), .C2(n9591), .A(n9601), .B(n9590), .ZN(n9593)
         );
  NAND2_X1 U10558 ( .A1(n9602), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9597) );
  NAND2_X1 U10559 ( .A1(n9598), .A2(n9597), .ZN(n9600) );
  XNOR2_X1 U10560 ( .A(n5608), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9599) );
  XNOR2_X1 U10561 ( .A(n9600), .B(n9599), .ZN(n9613) );
  MUX2_X1 U10562 ( .A(n9829), .B(P1_REG2_REG_19__SCAN_IN), .S(n5608), .Z(n9603) );
  XNOR2_X1 U10563 ( .A(n9604), .B(n9603), .ZN(n9605) );
  NAND2_X1 U10564 ( .A1(n9605), .A2(n10366), .ZN(n9612) );
  NAND2_X1 U10565 ( .A1(n10350), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n9607) );
  NAND2_X1 U10566 ( .A1(n9607), .A2(n9606), .ZN(n9608) );
  AOI21_X1 U10567 ( .B1(n9610), .B2(n9609), .A(n9608), .ZN(n9611) );
  OAI211_X1 U10568 ( .C1(n9613), .C2(n10362), .A(n9612), .B(n9611), .ZN(
        P1_U3262) );
  INV_X1 U10569 ( .A(n9982), .ZN(n9889) );
  NAND2_X1 U10570 ( .A1(n9883), .A2(n9889), .ZN(n9886) );
  NOR2_X2 U10571 ( .A1(n9886), .A2(n9868), .ZN(n9862) );
  NAND2_X1 U10572 ( .A1(n10031), .A2(n9862), .ZN(n9844) );
  NOR2_X2 U10573 ( .A1(n9933), .A2(n9762), .ZN(n9745) );
  NAND2_X1 U10574 ( .A1(n9999), .A2(n9645), .ZN(n9624) );
  XNOR2_X1 U10575 ( .A(n9621), .B(n9624), .ZN(n9616) );
  NOR2_X1 U10576 ( .A1(n10348), .A2(n9617), .ZN(n9618) );
  NOR2_X1 U10577 ( .A1(n9880), .A2(n9618), .ZN(n9667) );
  INV_X1 U10578 ( .A(n9667), .ZN(n9619) );
  NOR2_X1 U10579 ( .A1(n9685), .A2(n9898), .ZN(n9626) );
  NOR2_X1 U10580 ( .A1(n9995), .A2(n9888), .ZN(n9622) );
  AOI211_X1 U10581 ( .C1(n9685), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9626), .B(
        n9622), .ZN(n9623) );
  OAI21_X1 U10582 ( .B1(n9895), .B2(n9865), .A(n9623), .ZN(P1_U3263) );
  OAI211_X1 U10583 ( .C1(n9999), .C2(n9645), .A(n9884), .B(n9624), .ZN(n9899)
         );
  NOR2_X1 U10584 ( .A1(n10525), .A2(n9625), .ZN(n9627) );
  AOI211_X1 U10585 ( .C1(n9628), .C2(n9869), .A(n9627), .B(n9626), .ZN(n9629)
         );
  OAI21_X1 U10586 ( .B1(n9899), .B2(n9865), .A(n9629), .ZN(P1_U3264) );
  NAND2_X1 U10587 ( .A1(n10019), .A2(n9779), .ZN(n9640) );
  NAND2_X1 U10588 ( .A1(n9933), .A2(n9758), .ZN(n9641) );
  INV_X1 U10589 ( .A(n9933), .ZN(n9746) );
  NAND2_X1 U10590 ( .A1(n10014), .A2(n9921), .ZN(n9643) );
  AOI22_X1 U10591 ( .A1(n9715), .A2(n9716), .B1(n9702), .B2(n9724), .ZN(n9690)
         );
  INV_X1 U10592 ( .A(n9644), .ZN(n9673) );
  OAI22_X1 U10593 ( .A1(n10525), .A2(n9647), .B1(n9646), .B2(n10522), .ZN(
        n9648) );
  AOI21_X1 U10594 ( .B1(n9677), .B2(n9703), .A(n9648), .ZN(n9649) );
  OAI21_X1 U10595 ( .B1(n5499), .B2(n9888), .A(n9649), .ZN(n9669) );
  INV_X1 U10596 ( .A(n9793), .ZN(n9651) );
  INV_X1 U10597 ( .A(n9789), .ZN(n9650) );
  NOR2_X1 U10598 ( .A1(n9651), .A2(n9650), .ZN(n9652) );
  NAND2_X1 U10599 ( .A1(n9805), .A2(n9652), .ZN(n9654) );
  INV_X1 U10600 ( .A(n9662), .ZN(n9663) );
  NOR2_X1 U10601 ( .A1(n9681), .A2(n9663), .ZN(n9665) );
  XNOR2_X1 U10602 ( .A(n9665), .B(n9664), .ZN(n9668) );
  OAI21_X1 U10603 ( .B1(n9671), .B2(n9679), .A(n9670), .ZN(n9908) );
  INV_X1 U10604 ( .A(n9672), .ZN(n9692) );
  OAI211_X1 U10605 ( .C1(n10003), .C2(n9692), .A(n9673), .B(n9884), .ZN(n9909)
         );
  INV_X1 U10606 ( .A(n9909), .ZN(n9688) );
  OAI22_X1 U10607 ( .A1(n10525), .A2(n9675), .B1(n9674), .B2(n10522), .ZN(
        n9676) );
  AOI21_X1 U10608 ( .B1(n9677), .B2(n9712), .A(n9676), .ZN(n9678) );
  OAI21_X1 U10609 ( .B1(n10003), .B2(n9888), .A(n9678), .ZN(n9687) );
  NOR2_X1 U10610 ( .A1(n9682), .A2(n9880), .ZN(n9683) );
  NOR2_X1 U10611 ( .A1(n9910), .A2(n9685), .ZN(n9686) );
  OAI21_X1 U10612 ( .B1(n9908), .B2(n9894), .A(n9689), .ZN(P1_U3265) );
  XNOR2_X1 U10613 ( .A(n9690), .B(n9698), .ZN(n9916) );
  INV_X1 U10614 ( .A(n9916), .ZN(n9708) );
  AOI211_X1 U10615 ( .C1(n9693), .C2(n9721), .A(n9826), .B(n9692), .ZN(n9915)
         );
  NOR2_X1 U10616 ( .A1(n9615), .A2(n9888), .ZN(n9697) );
  OAI22_X1 U10617 ( .A1(n10525), .A2(n9695), .B1(n9694), .B2(n10522), .ZN(
        n9696) );
  AOI211_X1 U10618 ( .C1(n9915), .C2(n9891), .A(n9697), .B(n9696), .ZN(n9707)
         );
  NAND2_X1 U10619 ( .A1(n9699), .A2(n9698), .ZN(n9700) );
  NAND3_X1 U10620 ( .A1(n9701), .A2(n9852), .A3(n9700), .ZN(n9705) );
  AOI22_X1 U10621 ( .A1(n9703), .A2(n10519), .B1(n10704), .B2(n9702), .ZN(
        n9704) );
  NAND2_X1 U10622 ( .A1(n9705), .A2(n9704), .ZN(n9914) );
  NAND2_X1 U10623 ( .A1(n9914), .A2(n10525), .ZN(n9706) );
  OAI211_X1 U10624 ( .C1(n9708), .C2(n9894), .A(n9707), .B(n9706), .ZN(
        P1_U3266) );
  NAND2_X1 U10625 ( .A1(n9709), .A2(n9716), .ZN(n9710) );
  NAND2_X1 U10626 ( .A1(n9711), .A2(n9710), .ZN(n9714) );
  AND2_X1 U10627 ( .A1(n9712), .A2(n10519), .ZN(n9713) );
  AOI21_X1 U10628 ( .B1(n9714), .B2(n9852), .A(n9713), .ZN(n9920) );
  XOR2_X1 U10629 ( .A(n9716), .B(n9715), .Z(n9923) );
  NAND2_X1 U10630 ( .A1(n9923), .A2(n9855), .ZN(n9726) );
  INV_X1 U10631 ( .A(n9717), .ZN(n9718) );
  AOI22_X1 U10632 ( .A1(n9685), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9718), .B2(
        n9857), .ZN(n9719) );
  OAI21_X1 U10633 ( .B1(n9861), .B2(n9921), .A(n9719), .ZN(n9723) );
  INV_X1 U10634 ( .A(n9724), .ZN(n10010) );
  INV_X1 U10635 ( .A(n9720), .ZN(n9733) );
  OAI211_X1 U10636 ( .C1(n10010), .C2(n9733), .A(n9884), .B(n9721), .ZN(n9919)
         );
  NOR2_X1 U10637 ( .A1(n9919), .A2(n9865), .ZN(n9722) );
  AOI211_X1 U10638 ( .C1(n9869), .C2(n9724), .A(n9723), .B(n9722), .ZN(n9725)
         );
  OAI211_X1 U10639 ( .C1(n9685), .C2(n9920), .A(n9726), .B(n9725), .ZN(
        P1_U3267) );
  XOR2_X1 U10640 ( .A(n9731), .B(n9727), .Z(n9728) );
  OAI222_X1 U10641 ( .A1(n9880), .A2(n9730), .B1(n10631), .B2(n9729), .C1(
        n10529), .C2(n9728), .ZN(n9926) );
  INV_X1 U10642 ( .A(n9926), .ZN(n9742) );
  XOR2_X1 U10643 ( .A(n9732), .B(n9731), .Z(n9928) );
  NAND2_X1 U10644 ( .A1(n9928), .A2(n9855), .ZN(n9741) );
  INV_X1 U10645 ( .A(n9745), .ZN(n9734) );
  AOI211_X1 U10646 ( .C1(n9735), .C2(n9734), .A(n9826), .B(n9733), .ZN(n9927)
         );
  NOR2_X1 U10647 ( .A1(n10014), .A2(n9888), .ZN(n9739) );
  OAI22_X1 U10648 ( .A1(n10525), .A2(n9737), .B1(n9736), .B2(n10522), .ZN(
        n9738) );
  AOI211_X1 U10649 ( .C1(n9927), .C2(n9891), .A(n9739), .B(n9738), .ZN(n9740)
         );
  OAI211_X1 U10650 ( .C1(n9859), .C2(n9742), .A(n9741), .B(n9740), .ZN(
        P1_U3268) );
  XNOR2_X1 U10651 ( .A(n9744), .B(n9743), .ZN(n9935) );
  AOI211_X1 U10652 ( .C1(n9933), .C2(n9762), .A(n9826), .B(n9745), .ZN(n9932)
         );
  NOR2_X1 U10653 ( .A1(n9746), .A2(n9888), .ZN(n9750) );
  OAI22_X1 U10654 ( .A1(n10525), .A2(n9748), .B1(n9747), .B2(n10522), .ZN(
        n9749) );
  AOI211_X1 U10655 ( .C1(n9932), .C2(n9891), .A(n9750), .B(n9749), .ZN(n9755)
         );
  XNOR2_X1 U10656 ( .A(n9752), .B(n9751), .ZN(n9753) );
  OAI222_X1 U10657 ( .A1(n9880), .A2(n9921), .B1(n10631), .B2(n9779), .C1(
        n9753), .C2(n10529), .ZN(n9931) );
  NAND2_X1 U10658 ( .A1(n9931), .A2(n10525), .ZN(n9754) );
  OAI211_X1 U10659 ( .C1(n9935), .C2(n9894), .A(n9755), .B(n9754), .ZN(
        P1_U3269) );
  OAI21_X1 U10660 ( .B1(n9760), .B2(n9757), .A(n9756), .ZN(n9759) );
  AOI222_X1 U10661 ( .A1(n9852), .A2(n9759), .B1(n9758), .B2(n10519), .C1(
        n9791), .C2(n10704), .ZN(n9936) );
  XNOR2_X1 U10662 ( .A(n9761), .B(n9760), .ZN(n9939) );
  NAND2_X1 U10663 ( .A1(n9939), .A2(n9855), .ZN(n9770) );
  INV_X1 U10664 ( .A(n9762), .ZN(n9763) );
  AOI211_X1 U10665 ( .C1(n9764), .C2(n9780), .A(n9826), .B(n9763), .ZN(n9938)
         );
  INV_X1 U10666 ( .A(n9765), .ZN(n9766) );
  AOI22_X1 U10667 ( .A1(n9859), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9766), .B2(
        n9857), .ZN(n9767) );
  OAI21_X1 U10668 ( .B1(n10019), .B2(n9888), .A(n9767), .ZN(n9768) );
  AOI21_X1 U10669 ( .B1(n9938), .B2(n9891), .A(n9768), .ZN(n9769) );
  OAI211_X1 U10670 ( .C1(n9685), .C2(n9936), .A(n9770), .B(n9769), .ZN(
        P1_U3270) );
  XNOR2_X1 U10671 ( .A(n9772), .B(n9771), .ZN(n9946) );
  INV_X1 U10672 ( .A(n9773), .ZN(n9774) );
  AOI21_X1 U10673 ( .B1(n9776), .B2(n9775), .A(n9774), .ZN(n9777) );
  OAI222_X1 U10674 ( .A1(n9880), .A2(n9779), .B1(n10631), .B2(n9778), .C1(
        n10529), .C2(n9777), .ZN(n9942) );
  INV_X1 U10675 ( .A(n9780), .ZN(n9781) );
  AOI211_X1 U10676 ( .C1(n9944), .C2(n4951), .A(n9826), .B(n9781), .ZN(n9943)
         );
  NAND2_X1 U10677 ( .A1(n9943), .A2(n9891), .ZN(n9785) );
  INV_X1 U10678 ( .A(n9782), .ZN(n9783) );
  AOI22_X1 U10679 ( .A1(n9859), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9783), .B2(
        n9857), .ZN(n9784) );
  OAI211_X1 U10680 ( .C1(n9786), .C2(n9888), .A(n9785), .B(n9784), .ZN(n9787)
         );
  AOI21_X1 U10681 ( .B1(n9942), .B2(n10525), .A(n9787), .ZN(n9788) );
  OAI21_X1 U10682 ( .B1(n9946), .B2(n9894), .A(n9788), .ZN(P1_U3271) );
  NAND2_X1 U10683 ( .A1(n9805), .A2(n9789), .ZN(n9790) );
  XNOR2_X1 U10684 ( .A(n9790), .B(n9793), .ZN(n9792) );
  AOI22_X1 U10685 ( .A1(n9792), .A2(n9852), .B1(n10519), .B2(n9791), .ZN(n9948) );
  XNOR2_X1 U10686 ( .A(n9794), .B(n9793), .ZN(n9951) );
  NAND2_X1 U10687 ( .A1(n9951), .A2(n9855), .ZN(n9802) );
  INV_X1 U10688 ( .A(n9795), .ZN(n9796) );
  AOI22_X1 U10689 ( .A1(n9859), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9796), .B2(
        n9857), .ZN(n9797) );
  OAI21_X1 U10690 ( .B1(n9861), .B2(n9949), .A(n9797), .ZN(n9799) );
  OAI211_X1 U10691 ( .C1(n5236), .C2(n5005), .A(n4951), .B(n9884), .ZN(n9947)
         );
  NOR2_X1 U10692 ( .A1(n9947), .A2(n9865), .ZN(n9798) );
  AOI211_X1 U10693 ( .C1(n9869), .C2(n9800), .A(n9799), .B(n9798), .ZN(n9801)
         );
  OAI211_X1 U10694 ( .C1(n9685), .C2(n9948), .A(n9802), .B(n9801), .ZN(
        P1_U3272) );
  XNOR2_X1 U10695 ( .A(n9804), .B(n9803), .ZN(n9956) );
  INV_X1 U10696 ( .A(n9956), .ZN(n9819) );
  OAI21_X1 U10697 ( .B1(n9807), .B2(n9806), .A(n9805), .ZN(n9808) );
  NAND2_X1 U10698 ( .A1(n9808), .A2(n9852), .ZN(n9811) );
  AOI22_X1 U10699 ( .A1(n9809), .A2(n10519), .B1(n9836), .B2(n10704), .ZN(
        n9810) );
  NAND2_X1 U10700 ( .A1(n9811), .A2(n9810), .ZN(n9954) );
  INV_X1 U10701 ( .A(n9812), .ZN(n9825) );
  AOI211_X1 U10702 ( .C1(n9813), .C2(n9825), .A(n9826), .B(n5005), .ZN(n9955)
         );
  NAND2_X1 U10703 ( .A1(n9955), .A2(n9891), .ZN(n9816) );
  AOI22_X1 U10704 ( .A1(n9859), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9814), .B2(
        n9857), .ZN(n9815) );
  OAI211_X1 U10705 ( .C1(n9614), .C2(n9888), .A(n9816), .B(n9815), .ZN(n9817)
         );
  AOI21_X1 U10706 ( .B1(n9954), .B2(n10525), .A(n9817), .ZN(n9818) );
  OAI21_X1 U10707 ( .B1(n9819), .B2(n9894), .A(n9818), .ZN(P1_U3273) );
  XOR2_X1 U10708 ( .A(n9823), .B(n9820), .Z(n9821) );
  OAI222_X1 U10709 ( .A1(n9880), .A2(n9949), .B1(n10631), .B2(n9822), .C1(
        n10529), .C2(n9821), .ZN(n9960) );
  INV_X1 U10710 ( .A(n9960), .ZN(n9834) );
  NAND2_X1 U10711 ( .A1(n9824), .A2(n9823), .ZN(n9959) );
  NAND3_X1 U10712 ( .A1(n5089), .A2(n9855), .A3(n9959), .ZN(n9833) );
  AOI211_X1 U10713 ( .C1(n9962), .C2(n9844), .A(n9826), .B(n9812), .ZN(n9961)
         );
  INV_X1 U10714 ( .A(n9962), .ZN(n9827) );
  NOR2_X1 U10715 ( .A1(n9827), .A2(n9888), .ZN(n9831) );
  OAI22_X1 U10716 ( .A1(n10525), .A2(n9829), .B1(n9828), .B2(n10522), .ZN(
        n9830) );
  AOI211_X1 U10717 ( .C1(n9961), .C2(n9891), .A(n9831), .B(n9830), .ZN(n9832)
         );
  OAI211_X1 U10718 ( .C1(n9685), .C2(n9834), .A(n9833), .B(n9832), .ZN(
        P1_U3274) );
  XNOR2_X1 U10719 ( .A(n9835), .B(n5150), .ZN(n9838) );
  AND2_X1 U10720 ( .A1(n9836), .A2(n10519), .ZN(n9837) );
  AOI21_X1 U10721 ( .B1(n9838), .B2(n9852), .A(n9837), .ZN(n9967) );
  XOR2_X1 U10722 ( .A(n9839), .B(n9840), .Z(n9970) );
  NAND2_X1 U10723 ( .A1(n9970), .A2(n9855), .ZN(n9849) );
  INV_X1 U10724 ( .A(n9841), .ZN(n9842) );
  AOI22_X1 U10725 ( .A1(n9859), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9842), .B2(
        n9857), .ZN(n9843) );
  OAI21_X1 U10726 ( .B1(n9861), .B2(n9968), .A(n9843), .ZN(n9846) );
  OAI211_X1 U10727 ( .C1(n10031), .C2(n9862), .A(n9884), .B(n9844), .ZN(n9966)
         );
  NOR2_X1 U10728 ( .A1(n9966), .A2(n9865), .ZN(n9845) );
  AOI211_X1 U10729 ( .C1(n9869), .C2(n9847), .A(n9846), .B(n9845), .ZN(n9848)
         );
  OAI211_X1 U10730 ( .C1(n9685), .C2(n9967), .A(n9849), .B(n9848), .ZN(
        P1_U3275) );
  XNOR2_X1 U10731 ( .A(n9850), .B(n5251), .ZN(n9853) );
  AOI22_X1 U10732 ( .A1(n9853), .A2(n9852), .B1(n10519), .B2(n9851), .ZN(n9974) );
  XNOR2_X1 U10733 ( .A(n9854), .B(n5251), .ZN(n9977) );
  NAND2_X1 U10734 ( .A1(n9977), .A2(n9855), .ZN(n9871) );
  INV_X1 U10735 ( .A(n9856), .ZN(n9858) );
  AOI22_X1 U10736 ( .A1(n9859), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9858), .B2(
        n9857), .ZN(n9860) );
  OAI21_X1 U10737 ( .B1(n9861), .B2(n9975), .A(n9860), .ZN(n9867) );
  INV_X1 U10738 ( .A(n9868), .ZN(n10035) );
  INV_X1 U10739 ( .A(n9886), .ZN(n9864) );
  INV_X1 U10740 ( .A(n9862), .ZN(n9863) );
  OAI211_X1 U10741 ( .C1(n10035), .C2(n9864), .A(n9863), .B(n9884), .ZN(n9973)
         );
  NOR2_X1 U10742 ( .A1(n9973), .A2(n9865), .ZN(n9866) );
  AOI211_X1 U10743 ( .C1(n9869), .C2(n9868), .A(n9867), .B(n9866), .ZN(n9870)
         );
  OAI211_X1 U10744 ( .C1(n9685), .C2(n9974), .A(n9871), .B(n9870), .ZN(
        P1_U3276) );
  XNOR2_X1 U10745 ( .A(n9873), .B(n9872), .ZN(n9984) );
  INV_X1 U10746 ( .A(n9874), .ZN(n9875) );
  AOI21_X1 U10747 ( .B1(n9877), .B2(n9876), .A(n9875), .ZN(n9878) );
  OAI222_X1 U10748 ( .A1(n9880), .A2(n9968), .B1(n10631), .B2(n9879), .C1(
        n10529), .C2(n9878), .ZN(n9980) );
  NOR2_X1 U10749 ( .A1(n10522), .A2(n9881), .ZN(n9882) );
  OAI21_X1 U10750 ( .B1(n9980), .B2(n9882), .A(n10525), .ZN(n9893) );
  OR2_X1 U10751 ( .A1(n9883), .A2(n9889), .ZN(n9885) );
  AND3_X1 U10752 ( .A1(n9886), .A2(n9885), .A3(n9884), .ZN(n9981) );
  OAI22_X1 U10753 ( .A1(n9889), .A2(n9888), .B1(n9887), .B2(n10525), .ZN(n9890) );
  AOI21_X1 U10754 ( .B1(n9981), .B2(n9891), .A(n9890), .ZN(n9892) );
  OAI211_X1 U10755 ( .C1(n9984), .C2(n9894), .A(n9893), .B(n9892), .ZN(
        P1_U3277) );
  MUX2_X1 U10756 ( .A(n9896), .B(n9992), .S(n10736), .Z(n9897) );
  OAI21_X1 U10757 ( .B1(n9995), .B2(n9991), .A(n9897), .ZN(P1_U3553) );
  AND2_X1 U10758 ( .A1(n9899), .A2(n9898), .ZN(n9996) );
  MUX2_X1 U10759 ( .A(n9900), .B(n9996), .S(n10736), .Z(n9901) );
  OAI21_X1 U10760 ( .B1(n9999), .B2(n9991), .A(n9901), .ZN(P1_U3552) );
  MUX2_X1 U10761 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10000), .S(n10736), .Z(
        P1_U3551) );
  INV_X1 U10762 ( .A(n9908), .ZN(n9912) );
  AOI211_X1 U10763 ( .C1(n9916), .C2(n10711), .A(n9915), .B(n9914), .ZN(n10004) );
  MUX2_X1 U10764 ( .A(n9917), .B(n10004), .S(n10736), .Z(n9918) );
  OAI21_X1 U10765 ( .B1(n9615), .B2(n9991), .A(n9918), .ZN(P1_U3549) );
  OAI211_X1 U10766 ( .C1(n9921), .C2(n10631), .A(n9920), .B(n9919), .ZN(n9922)
         );
  AOI21_X1 U10767 ( .B1(n9923), .B2(n10711), .A(n9922), .ZN(n10007) );
  MUX2_X1 U10768 ( .A(n9924), .B(n10007), .S(n10736), .Z(n9925) );
  OAI21_X1 U10769 ( .B1(n10010), .B2(n9991), .A(n9925), .ZN(P1_U3548) );
  INV_X1 U10770 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9929) );
  AOI211_X1 U10771 ( .C1(n9928), .C2(n10711), .A(n9927), .B(n9926), .ZN(n10011) );
  MUX2_X1 U10772 ( .A(n9929), .B(n10011), .S(n10736), .Z(n9930) );
  OAI21_X1 U10773 ( .B1(n10014), .B2(n9991), .A(n9930), .ZN(P1_U3547) );
  AOI211_X1 U10774 ( .C1(n10705), .C2(n9933), .A(n9932), .B(n9931), .ZN(n9934)
         );
  OAI21_X1 U10775 ( .B1(n9935), .B2(n10528), .A(n9934), .ZN(n10015) );
  MUX2_X1 U10776 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10015), .S(n10736), .Z(
        P1_U3546) );
  INV_X1 U10777 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9940) );
  INV_X1 U10778 ( .A(n9936), .ZN(n9937) );
  AOI211_X1 U10779 ( .C1(n9939), .C2(n10711), .A(n9938), .B(n9937), .ZN(n10016) );
  MUX2_X1 U10780 ( .A(n9940), .B(n10016), .S(n10736), .Z(n9941) );
  OAI21_X1 U10781 ( .B1(n10019), .B2(n9991), .A(n9941), .ZN(P1_U3545) );
  AOI211_X1 U10782 ( .C1(n10705), .C2(n9944), .A(n9943), .B(n9942), .ZN(n9945)
         );
  OAI21_X1 U10783 ( .B1(n9946), .B2(n10528), .A(n9945), .ZN(n10020) );
  MUX2_X1 U10784 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10020), .S(n10736), .Z(
        P1_U3544) );
  OAI211_X1 U10785 ( .C1(n9949), .C2(n10631), .A(n9948), .B(n9947), .ZN(n9950)
         );
  AOI21_X1 U10786 ( .B1(n9951), .B2(n10711), .A(n9950), .ZN(n10021) );
  MUX2_X1 U10787 ( .A(n9952), .B(n10021), .S(n10736), .Z(n9953) );
  OAI21_X1 U10788 ( .B1(n5236), .B2(n9991), .A(n9953), .ZN(P1_U3543) );
  AOI211_X1 U10789 ( .C1(n9956), .C2(n10711), .A(n9955), .B(n9954), .ZN(n10024) );
  MUX2_X1 U10790 ( .A(n9957), .B(n10024), .S(n10736), .Z(n9958) );
  OAI21_X1 U10791 ( .B1(n9614), .B2(n9991), .A(n9958), .ZN(P1_U3542) );
  NAND2_X1 U10792 ( .A1(n9959), .A2(n10711), .ZN(n9964) );
  AOI211_X1 U10793 ( .C1(n10705), .C2(n9962), .A(n9961), .B(n9960), .ZN(n9963)
         );
  OAI21_X1 U10794 ( .B1(n9965), .B2(n9964), .A(n9963), .ZN(n10027) );
  MUX2_X1 U10795 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10027), .S(n10736), .Z(
        P1_U3541) );
  OAI211_X1 U10796 ( .C1(n9968), .C2(n10631), .A(n9967), .B(n9966), .ZN(n9969)
         );
  AOI21_X1 U10797 ( .B1(n9970), .B2(n10711), .A(n9969), .ZN(n10028) );
  MUX2_X1 U10798 ( .A(n9971), .B(n10028), .S(n10736), .Z(n9972) );
  OAI21_X1 U10799 ( .B1(n10031), .B2(n9991), .A(n9972), .ZN(P1_U3540) );
  OAI211_X1 U10800 ( .C1(n9975), .C2(n10631), .A(n9974), .B(n9973), .ZN(n9976)
         );
  AOI21_X1 U10801 ( .B1(n9977), .B2(n10711), .A(n9976), .ZN(n10032) );
  MUX2_X1 U10802 ( .A(n9978), .B(n10032), .S(n10736), .Z(n9979) );
  OAI21_X1 U10803 ( .B1(n10035), .B2(n9991), .A(n9979), .ZN(P1_U3539) );
  AOI211_X1 U10804 ( .C1(n10705), .C2(n9982), .A(n9981), .B(n9980), .ZN(n9983)
         );
  OAI21_X1 U10805 ( .B1(n10528), .B2(n9984), .A(n9983), .ZN(n10036) );
  MUX2_X1 U10806 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10036), .S(n10736), .Z(
        P1_U3538) );
  OAI211_X1 U10807 ( .C1(n9987), .C2(n10631), .A(n9986), .B(n9985), .ZN(n9988)
         );
  AOI21_X1 U10808 ( .B1(n9989), .B2(n10711), .A(n9988), .ZN(n10037) );
  MUX2_X1 U10809 ( .A(n6010), .B(n10037), .S(n10736), .Z(n9990) );
  OAI21_X1 U10810 ( .B1(n5202), .B2(n9991), .A(n9990), .ZN(P1_U3537) );
  INV_X1 U10811 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9993) );
  MUX2_X1 U10812 ( .A(n9993), .B(n9992), .S(n10740), .Z(n9994) );
  OAI21_X1 U10813 ( .B1(n9995), .B2(n10040), .A(n9994), .ZN(P1_U3521) );
  INV_X1 U10814 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9997) );
  MUX2_X1 U10815 ( .A(n9997), .B(n9996), .S(n10740), .Z(n9998) );
  OAI21_X1 U10816 ( .B1(n9999), .B2(n10040), .A(n9998), .ZN(P1_U3520) );
  INV_X1 U10817 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10002) );
  INV_X1 U10818 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10005) );
  MUX2_X1 U10819 ( .A(n10005), .B(n10004), .S(n10740), .Z(n10006) );
  OAI21_X1 U10820 ( .B1(n9615), .B2(n10040), .A(n10006), .ZN(P1_U3517) );
  INV_X1 U10821 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10008) );
  MUX2_X1 U10822 ( .A(n10008), .B(n10007), .S(n10740), .Z(n10009) );
  OAI21_X1 U10823 ( .B1(n10010), .B2(n10040), .A(n10009), .ZN(P1_U3516) );
  MUX2_X1 U10824 ( .A(n10012), .B(n10011), .S(n10740), .Z(n10013) );
  OAI21_X1 U10825 ( .B1(n10014), .B2(n10040), .A(n10013), .ZN(P1_U3515) );
  MUX2_X1 U10826 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10015), .S(n10740), .Z(
        P1_U3514) );
  INV_X1 U10827 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10017) );
  MUX2_X1 U10828 ( .A(n10017), .B(n10016), .S(n10740), .Z(n10018) );
  OAI21_X1 U10829 ( .B1(n10019), .B2(n10040), .A(n10018), .ZN(P1_U3513) );
  MUX2_X1 U10830 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10020), .S(n10740), .Z(
        P1_U3512) );
  INV_X1 U10831 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10022) );
  MUX2_X1 U10832 ( .A(n10022), .B(n10021), .S(n10740), .Z(n10023) );
  OAI21_X1 U10833 ( .B1(n5236), .B2(n10040), .A(n10023), .ZN(P1_U3511) );
  MUX2_X1 U10834 ( .A(n10025), .B(n10024), .S(n10740), .Z(n10026) );
  OAI21_X1 U10835 ( .B1(n9614), .B2(n10040), .A(n10026), .ZN(P1_U3510) );
  MUX2_X1 U10836 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10027), .S(n10740), .Z(
        P1_U3509) );
  MUX2_X1 U10837 ( .A(n10029), .B(n10028), .S(n10740), .Z(n10030) );
  OAI21_X1 U10838 ( .B1(n10031), .B2(n10040), .A(n10030), .ZN(P1_U3507) );
  INV_X1 U10839 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10033) );
  MUX2_X1 U10840 ( .A(n10033), .B(n10032), .S(n10740), .Z(n10034) );
  OAI21_X1 U10841 ( .B1(n10035), .B2(n10040), .A(n10034), .ZN(P1_U3504) );
  MUX2_X1 U10842 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10036), .S(n10740), .Z(
        P1_U3501) );
  INV_X1 U10843 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10038) );
  MUX2_X1 U10844 ( .A(n10038), .B(n10037), .S(n10740), .Z(n10039) );
  OAI21_X1 U10845 ( .B1(n5202), .B2(n10040), .A(n10039), .ZN(P1_U3498) );
  INV_X1 U10846 ( .A(n10041), .ZN(n10043) );
  MUX2_X1 U10847 ( .A(n10044), .B(P1_D_REG_1__SCAN_IN), .S(n4930), .Z(P1_U3440) );
  MUX2_X1 U10848 ( .A(n10045), .B(P1_D_REG_0__SCAN_IN), .S(n4930), .Z(P1_U3439) );
  NAND3_X1 U10849 ( .A1(n10046), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n10048) );
  OAI22_X1 U10850 ( .A1(n5265), .A2(n10048), .B1(n10047), .B2(n10284), .ZN(
        n10049) );
  AOI21_X1 U10851 ( .B1(n10050), .B2(n10054), .A(n10049), .ZN(n10051) );
  INV_X1 U10852 ( .A(n10051), .ZN(P1_U3324) );
  AOI222_X1 U10853 ( .A1(n10055), .A2(n10054), .B1(n10052), .B2(
        P1_STATE_REG_SCAN_IN), .C1(P2_DATAO_REG_30__SCAN_IN), .C2(n10053), 
        .ZN(n10276) );
  OAI22_X1 U10854 ( .A1(n10265), .A2(keyinput_62), .B1(keyinput_61), .B2(
        P2_REG3_REG_6__SCAN_IN), .ZN(n10056) );
  AOI221_X1 U10855 ( .B1(n10265), .B2(keyinput_62), .C1(P2_REG3_REG_6__SCAN_IN), .C2(keyinput_61), .A(n10056), .ZN(n10274) );
  INV_X1 U10856 ( .A(keyinput_60), .ZN(n10154) );
  INV_X1 U10857 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10263) );
  INV_X1 U10858 ( .A(keyinput_59), .ZN(n10151) );
  OAI22_X1 U10859 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_51), .B1(
        keyinput_48), .B2(P2_REG3_REG_16__SCAN_IN), .ZN(n10057) );
  AOI221_X1 U10860 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_51), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_48), .A(n10057), .ZN(n10139) );
  OAI22_X1 U10861 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_50), .B1(
        keyinput_52), .B2(P2_REG3_REG_4__SCAN_IN), .ZN(n10058) );
  AOI221_X1 U10862 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_50), .C1(
        P2_REG3_REG_4__SCAN_IN), .C2(keyinput_52), .A(n10058), .ZN(n10138) );
  OAI22_X1 U10863 ( .A1(n6979), .A2(keyinput_53), .B1(n6975), .B2(keyinput_49), 
        .ZN(n10059) );
  AOI221_X1 U10864 ( .B1(n6979), .B2(keyinput_53), .C1(keyinput_49), .C2(n6975), .A(n10059), .ZN(n10137) );
  INV_X1 U10865 ( .A(keyinput_41), .ZN(n10125) );
  INV_X1 U10866 ( .A(keyinput_40), .ZN(n10123) );
  INV_X1 U10867 ( .A(keyinput_39), .ZN(n10121) );
  INV_X1 U10868 ( .A(keyinput_16), .ZN(n10084) );
  OAI22_X1 U10869 ( .A1(n10188), .A2(keyinput_15), .B1(SI_18_), .B2(
        keyinput_14), .ZN(n10060) );
  AOI221_X1 U10870 ( .B1(n10188), .B2(keyinput_15), .C1(keyinput_14), .C2(
        SI_18_), .A(n10060), .ZN(n10081) );
  INV_X1 U10871 ( .A(keyinput_12), .ZN(n10079) );
  INV_X1 U10872 ( .A(keyinput_11), .ZN(n10077) );
  INV_X1 U10873 ( .A(keyinput_10), .ZN(n10075) );
  OAI22_X1 U10874 ( .A1(n10062), .A2(keyinput_4), .B1(SI_29_), .B2(keyinput_3), 
        .ZN(n10061) );
  AOI221_X1 U10875 ( .B1(n10062), .B2(keyinput_4), .C1(keyinput_3), .C2(SI_29_), .A(n10061), .ZN(n10069) );
  INV_X1 U10876 ( .A(keyinput_2), .ZN(n10065) );
  OAI22_X1 U10877 ( .A1(SI_31_), .A2(keyinput_1), .B1(P2_WR_REG_SCAN_IN), .B2(
        keyinput_0), .ZN(n10063) );
  AOI221_X1 U10878 ( .B1(SI_31_), .B2(keyinput_1), .C1(keyinput_0), .C2(
        P2_WR_REG_SCAN_IN), .A(n10063), .ZN(n10064) );
  OAI221_X1 U10879 ( .B1(SI_30_), .B2(keyinput_2), .C1(n10166), .C2(n10065), 
        .A(n10064), .ZN(n10068) );
  AOI22_X1 U10880 ( .A1(SI_27_), .A2(keyinput_5), .B1(n10170), .B2(keyinput_6), 
        .ZN(n10066) );
  OAI221_X1 U10881 ( .B1(SI_27_), .B2(keyinput_5), .C1(n10170), .C2(keyinput_6), .A(n10066), .ZN(n10067) );
  AOI21_X1 U10882 ( .B1(n10069), .B2(n10068), .A(n10067), .ZN(n10072) );
  AOI22_X1 U10883 ( .A1(SI_23_), .A2(keyinput_9), .B1(n10177), .B2(keyinput_8), 
        .ZN(n10070) );
  OAI221_X1 U10884 ( .B1(SI_23_), .B2(keyinput_9), .C1(n10177), .C2(keyinput_8), .A(n10070), .ZN(n10071) );
  AOI211_X1 U10885 ( .C1(n10163), .C2(keyinput_7), .A(n10072), .B(n10071), 
        .ZN(n10073) );
  OAI21_X1 U10886 ( .B1(n10163), .B2(keyinput_7), .A(n10073), .ZN(n10074) );
  OAI221_X1 U10887 ( .B1(SI_22_), .B2(keyinput_10), .C1(n10180), .C2(n10075), 
        .A(n10074), .ZN(n10076) );
  OAI221_X1 U10888 ( .B1(SI_21_), .B2(n10077), .C1(n10183), .C2(keyinput_11), 
        .A(n10076), .ZN(n10078) );
  OAI221_X1 U10889 ( .B1(SI_20_), .B2(keyinput_12), .C1(n10186), .C2(n10079), 
        .A(n10078), .ZN(n10080) );
  OAI211_X1 U10890 ( .C1(SI_19_), .C2(keyinput_13), .A(n10081), .B(n10080), 
        .ZN(n10082) );
  AOI21_X1 U10891 ( .B1(SI_19_), .B2(keyinput_13), .A(n10082), .ZN(n10083) );
  AOI221_X1 U10892 ( .B1(SI_16_), .B2(n10084), .C1(n10195), .C2(keyinput_16), 
        .A(n10083), .ZN(n10087) );
  AOI22_X1 U10893 ( .A1(SI_14_), .A2(keyinput_18), .B1(SI_15_), .B2(
        keyinput_17), .ZN(n10085) );
  OAI221_X1 U10894 ( .B1(SI_14_), .B2(keyinput_18), .C1(SI_15_), .C2(
        keyinput_17), .A(n10085), .ZN(n10086) );
  OAI22_X1 U10895 ( .A1(n10087), .A2(n10086), .B1(SI_13_), .B2(keyinput_19), 
        .ZN(n10091) );
  INV_X1 U10896 ( .A(SI_12_), .ZN(n10089) );
  OAI22_X1 U10897 ( .A1(n10089), .A2(keyinput_20), .B1(SI_9_), .B2(keyinput_23), .ZN(n10088) );
  AOI221_X1 U10898 ( .B1(n10089), .B2(keyinput_20), .C1(keyinput_23), .C2(
        SI_9_), .A(n10088), .ZN(n10090) );
  OAI221_X1 U10899 ( .B1(n10091), .B2(keyinput_19), .C1(n10091), .C2(SI_13_), 
        .A(n10090), .ZN(n10095) );
  INV_X1 U10900 ( .A(SI_11_), .ZN(n10204) );
  AOI22_X1 U10901 ( .A1(n10199), .A2(keyinput_22), .B1(n10204), .B2(
        keyinput_21), .ZN(n10092) );
  OAI221_X1 U10902 ( .B1(n10199), .B2(keyinput_22), .C1(n10204), .C2(
        keyinput_21), .A(n10092), .ZN(n10094) );
  NAND2_X1 U10903 ( .A1(keyinput_25), .A2(SI_7_), .ZN(n10093) );
  OAI221_X1 U10904 ( .B1(n10095), .B2(n10094), .C1(keyinput_25), .C2(SI_7_), 
        .A(n10093), .ZN(n10102) );
  AOI22_X1 U10905 ( .A1(n10210), .A2(keyinput_24), .B1(keyinput_26), .B2(
        n10097), .ZN(n10096) );
  OAI221_X1 U10906 ( .B1(n10210), .B2(keyinput_24), .C1(n10097), .C2(
        keyinput_26), .A(n10096), .ZN(n10101) );
  XNOR2_X1 U10907 ( .A(n10098), .B(keyinput_27), .ZN(n10100) );
  XNOR2_X1 U10908 ( .A(SI_4_), .B(keyinput_28), .ZN(n10099) );
  OAI211_X1 U10909 ( .C1(n10102), .C2(n10101), .A(n10100), .B(n10099), .ZN(
        n10113) );
  INV_X1 U10910 ( .A(keyinput_29), .ZN(n10103) );
  MUX2_X1 U10911 ( .A(n10103), .B(keyinput_29), .S(SI_3_), .Z(n10112) );
  INV_X1 U10912 ( .A(SI_0_), .ZN(n10105) );
  OAI22_X1 U10913 ( .A1(n10105), .A2(keyinput_32), .B1(P2_RD_REG_SCAN_IN), 
        .B2(keyinput_33), .ZN(n10104) );
  AOI221_X1 U10914 ( .B1(n10105), .B2(keyinput_32), .C1(keyinput_33), .C2(
        P2_RD_REG_SCAN_IN), .A(n10104), .ZN(n10106) );
  OAI21_X1 U10915 ( .B1(keyinput_31), .B2(SI_1_), .A(n10106), .ZN(n10111) );
  INV_X1 U10916 ( .A(keyinput_31), .ZN(n10109) );
  XNOR2_X1 U10917 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_34), .ZN(n10108) );
  XNOR2_X1 U10918 ( .A(SI_2_), .B(keyinput_30), .ZN(n10107) );
  OAI211_X1 U10919 ( .C1(n10221), .C2(n10109), .A(n10108), .B(n10107), .ZN(
        n10110) );
  AOI211_X1 U10920 ( .C1(n10113), .C2(n10112), .A(n10111), .B(n10110), .ZN(
        n10119) );
  AOI22_X1 U10921 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_36), .B1(n10115), .B2(keyinput_37), .ZN(n10114) );
  OAI221_X1 U10922 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_36), .C1(
        n10115), .C2(keyinput_37), .A(n10114), .ZN(n10118) );
  INV_X1 U10923 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10228) );
  AOI22_X1 U10924 ( .A1(n6977), .A2(keyinput_35), .B1(n10228), .B2(keyinput_38), .ZN(n10116) );
  OAI221_X1 U10925 ( .B1(n6977), .B2(keyinput_35), .C1(n10228), .C2(
        keyinput_38), .A(n10116), .ZN(n10117) );
  NOR3_X1 U10926 ( .A1(n10119), .A2(n10118), .A3(n10117), .ZN(n10120) );
  AOI221_X1 U10927 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(n10121), .C1(n10234), 
        .C2(keyinput_39), .A(n10120), .ZN(n10122) );
  AOI221_X1 U10928 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_40), .C1(n7084), 
        .C2(n10123), .A(n10122), .ZN(n10124) );
  AOI221_X1 U10929 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_41), .C1(
        n10239), .C2(n10125), .A(n10124), .ZN(n10135) );
  INV_X1 U10930 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10127) );
  AOI22_X1 U10931 ( .A1(n10128), .A2(keyinput_43), .B1(n10127), .B2(
        keyinput_42), .ZN(n10126) );
  OAI221_X1 U10932 ( .B1(n10128), .B2(keyinput_43), .C1(n10127), .C2(
        keyinput_42), .A(n10126), .ZN(n10134) );
  INV_X1 U10933 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10130) );
  OAI22_X1 U10934 ( .A1(n10242), .A2(keyinput_46), .B1(n10130), .B2(
        keyinput_44), .ZN(n10129) );
  AOI221_X1 U10935 ( .B1(n10242), .B2(keyinput_46), .C1(keyinput_44), .C2(
        n10130), .A(n10129), .ZN(n10133) );
  OAI22_X1 U10936 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_47), .B1(
        keyinput_45), .B2(P2_REG3_REG_21__SCAN_IN), .ZN(n10131) );
  AOI221_X1 U10937 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_47), .C1(
        P2_REG3_REG_21__SCAN_IN), .C2(keyinput_45), .A(n10131), .ZN(n10132) );
  OAI211_X1 U10938 ( .C1(n10135), .C2(n10134), .A(n10133), .B(n10132), .ZN(
        n10136) );
  NAND4_X1 U10939 ( .A1(n10139), .A2(n10138), .A3(n10137), .A4(n10136), .ZN(
        n10142) );
  INV_X1 U10940 ( .A(keyinput_54), .ZN(n10140) );
  MUX2_X1 U10941 ( .A(n10140), .B(keyinput_54), .S(P2_REG3_REG_0__SCAN_IN), 
        .Z(n10141) );
  NAND2_X1 U10942 ( .A1(n10142), .A2(n10141), .ZN(n10149) );
  OAI22_X1 U10943 ( .A1(n10144), .A2(keyinput_58), .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_57), .ZN(n10143) );
  AOI221_X1 U10944 ( .B1(n10144), .B2(keyinput_58), .C1(keyinput_57), .C2(
        P2_REG3_REG_22__SCAN_IN), .A(n10143), .ZN(n10148) );
  INV_X1 U10945 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10146) );
  OAI22_X1 U10946 ( .A1(n10146), .A2(keyinput_55), .B1(n6981), .B2(keyinput_56), .ZN(n10145) );
  AOI221_X1 U10947 ( .B1(n10146), .B2(keyinput_55), .C1(keyinput_56), .C2(
        n6981), .A(n10145), .ZN(n10147) );
  NAND3_X1 U10948 ( .A1(n10149), .A2(n10148), .A3(n10147), .ZN(n10150) );
  OAI221_X1 U10949 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_59), .C1(n10263), .C2(n10151), .A(n10150), .ZN(n10152) );
  OAI221_X1 U10950 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(n10154), .C1(n10153), 
        .C2(keyinput_60), .A(n10152), .ZN(n10273) );
  XOR2_X1 U10951 ( .A(keyinput_63), .B(keyinput_127), .Z(n10271) );
  XNOR2_X1 U10952 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_124), .ZN(n10268)
         );
  INV_X1 U10953 ( .A(keyinput_123), .ZN(n10262) );
  OAI22_X1 U10954 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_112), .B1(
        keyinput_113), .B2(P2_REG3_REG_5__SCAN_IN), .ZN(n10155) );
  AOI221_X1 U10955 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_112), .C1(
        P2_REG3_REG_5__SCAN_IN), .C2(keyinput_113), .A(n10155), .ZN(n10251) );
  OAI22_X1 U10956 ( .A1(n6985), .A2(keyinput_114), .B1(keyinput_117), .B2(
        P2_REG3_REG_9__SCAN_IN), .ZN(n10156) );
  AOI221_X1 U10957 ( .B1(n6985), .B2(keyinput_114), .C1(P2_REG3_REG_9__SCAN_IN), .C2(keyinput_117), .A(n10156), .ZN(n10250) );
  OAI22_X1 U10958 ( .A1(n10158), .A2(keyinput_115), .B1(n6866), .B2(
        keyinput_116), .ZN(n10157) );
  AOI221_X1 U10959 ( .B1(n10158), .B2(keyinput_115), .C1(keyinput_116), .C2(
        n6866), .A(n10157), .ZN(n10249) );
  INV_X1 U10960 ( .A(keyinput_105), .ZN(n10238) );
  INV_X1 U10961 ( .A(keyinput_104), .ZN(n10236) );
  INV_X1 U10962 ( .A(keyinput_103), .ZN(n10233) );
  INV_X1 U10963 ( .A(SI_14_), .ZN(n10160) );
  OAI22_X1 U10964 ( .A1(n10160), .A2(keyinput_82), .B1(SI_15_), .B2(
        keyinput_81), .ZN(n10159) );
  AOI221_X1 U10965 ( .B1(n10160), .B2(keyinput_82), .C1(keyinput_81), .C2(
        SI_15_), .A(n10159), .ZN(n10197) );
  INV_X1 U10966 ( .A(keyinput_80), .ZN(n10194) );
  INV_X1 U10967 ( .A(keyinput_76), .ZN(n10185) );
  INV_X1 U10968 ( .A(keyinput_75), .ZN(n10182) );
  INV_X1 U10969 ( .A(keyinput_74), .ZN(n10179) );
  OAI22_X1 U10970 ( .A1(n10163), .A2(keyinput_71), .B1(n10162), .B2(
        keyinput_73), .ZN(n10161) );
  AOI221_X1 U10971 ( .B1(n10163), .B2(keyinput_71), .C1(keyinput_73), .C2(
        n10162), .A(n10161), .ZN(n10175) );
  INV_X1 U10972 ( .A(keyinput_66), .ZN(n10167) );
  AOI22_X1 U10973 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_64), .B1(SI_31_), 
        .B2(keyinput_65), .ZN(n10164) );
  OAI221_X1 U10974 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_64), .C1(SI_31_), 
        .C2(keyinput_65), .A(n10164), .ZN(n10165) );
  AOI221_X1 U10975 ( .B1(SI_30_), .B2(n10167), .C1(n10166), .C2(keyinput_66), 
        .A(n10165), .ZN(n10173) );
  AOI22_X1 U10976 ( .A1(SI_29_), .A2(keyinput_67), .B1(SI_28_), .B2(
        keyinput_68), .ZN(n10168) );
  OAI221_X1 U10977 ( .B1(SI_29_), .B2(keyinput_67), .C1(SI_28_), .C2(
        keyinput_68), .A(n10168), .ZN(n10172) );
  OAI22_X1 U10978 ( .A1(n10170), .A2(keyinput_70), .B1(keyinput_69), .B2(
        SI_27_), .ZN(n10169) );
  AOI221_X1 U10979 ( .B1(n10170), .B2(keyinput_70), .C1(SI_27_), .C2(
        keyinput_69), .A(n10169), .ZN(n10171) );
  OAI21_X1 U10980 ( .B1(n10173), .B2(n10172), .A(n10171), .ZN(n10174) );
  OAI211_X1 U10981 ( .C1(n10177), .C2(keyinput_72), .A(n10175), .B(n10174), 
        .ZN(n10176) );
  AOI21_X1 U10982 ( .B1(n10177), .B2(keyinput_72), .A(n10176), .ZN(n10178) );
  AOI221_X1 U10983 ( .B1(SI_22_), .B2(keyinput_74), .C1(n10180), .C2(n10179), 
        .A(n10178), .ZN(n10181) );
  AOI221_X1 U10984 ( .B1(SI_21_), .B2(keyinput_75), .C1(n10183), .C2(n10182), 
        .A(n10181), .ZN(n10184) );
  AOI221_X1 U10985 ( .B1(SI_20_), .B2(keyinput_76), .C1(n10186), .C2(n10185), 
        .A(n10184), .ZN(n10190) );
  AOI22_X1 U10986 ( .A1(SI_18_), .A2(keyinput_78), .B1(n10188), .B2(
        keyinput_79), .ZN(n10187) );
  OAI221_X1 U10987 ( .B1(SI_18_), .B2(keyinput_78), .C1(n10188), .C2(
        keyinput_79), .A(n10187), .ZN(n10189) );
  AOI211_X1 U10988 ( .C1(n10192), .C2(keyinput_77), .A(n10190), .B(n10189), 
        .ZN(n10191) );
  OAI21_X1 U10989 ( .B1(n10192), .B2(keyinput_77), .A(n10191), .ZN(n10193) );
  OAI221_X1 U10990 ( .B1(SI_16_), .B2(keyinput_80), .C1(n10195), .C2(n10194), 
        .A(n10193), .ZN(n10196) );
  AOI22_X1 U10991 ( .A1(SI_13_), .A2(keyinput_83), .B1(n10197), .B2(n10196), 
        .ZN(n10201) );
  AOI22_X1 U10992 ( .A1(SI_12_), .A2(keyinput_84), .B1(n10199), .B2(
        keyinput_86), .ZN(n10198) );
  OAI221_X1 U10993 ( .B1(SI_12_), .B2(keyinput_84), .C1(n10199), .C2(
        keyinput_86), .A(n10198), .ZN(n10200) );
  AOI221_X1 U10994 ( .B1(SI_13_), .B2(n10201), .C1(keyinput_83), .C2(n10201), 
        .A(n10200), .ZN(n10206) );
  OAI22_X1 U10995 ( .A1(n10204), .A2(keyinput_85), .B1(n10203), .B2(
        keyinput_87), .ZN(n10202) );
  AOI221_X1 U10996 ( .B1(n10204), .B2(keyinput_85), .C1(keyinput_87), .C2(
        n10203), .A(n10202), .ZN(n10205) );
  AOI22_X1 U10997 ( .A1(n10206), .A2(n10205), .B1(keyinput_89), .B2(n10208), 
        .ZN(n10207) );
  OAI21_X1 U10998 ( .B1(keyinput_89), .B2(n10208), .A(n10207), .ZN(n10214) );
  AOI22_X1 U10999 ( .A1(SI_6_), .A2(keyinput_90), .B1(n10210), .B2(keyinput_88), .ZN(n10209) );
  OAI221_X1 U11000 ( .B1(SI_6_), .B2(keyinput_90), .C1(n10210), .C2(
        keyinput_88), .A(n10209), .ZN(n10213) );
  OAI22_X1 U11001 ( .A1(SI_5_), .A2(keyinput_91), .B1(keyinput_92), .B2(SI_4_), 
        .ZN(n10211) );
  AOI221_X1 U11002 ( .B1(SI_5_), .B2(keyinput_91), .C1(SI_4_), .C2(keyinput_92), .A(n10211), .ZN(n10212) );
  OAI21_X1 U11003 ( .B1(n10214), .B2(n10213), .A(n10212), .ZN(n10225) );
  INV_X1 U11004 ( .A(keyinput_93), .ZN(n10215) );
  MUX2_X1 U11005 ( .A(n10215), .B(keyinput_93), .S(SI_3_), .Z(n10224) );
  OAI22_X1 U11006 ( .A1(n5573), .A2(keyinput_97), .B1(SI_0_), .B2(keyinput_96), 
        .ZN(n10216) );
  AOI221_X1 U11007 ( .B1(n5573), .B2(keyinput_97), .C1(keyinput_96), .C2(SI_0_), .A(n10216), .ZN(n10217) );
  OAI21_X1 U11008 ( .B1(keyinput_95), .B2(SI_1_), .A(n10217), .ZN(n10223) );
  INV_X1 U11009 ( .A(keyinput_95), .ZN(n10220) );
  XNOR2_X1 U11010 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_98), .ZN(n10219) );
  XNOR2_X1 U11011 ( .A(SI_2_), .B(keyinput_94), .ZN(n10218) );
  OAI211_X1 U11012 ( .C1(n10221), .C2(n10220), .A(n10219), .B(n10218), .ZN(
        n10222) );
  AOI211_X1 U11013 ( .C1(n10225), .C2(n10224), .A(n10223), .B(n10222), .ZN(
        n10231) );
  AOI22_X1 U11014 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_101), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_100), .ZN(n10226) );
  OAI221_X1 U11015 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_101), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_100), .A(n10226), .ZN(n10230)
         );
  AOI22_X1 U11016 ( .A1(n10228), .A2(keyinput_102), .B1(keyinput_99), .B2(
        n6977), .ZN(n10227) );
  OAI221_X1 U11017 ( .B1(n10228), .B2(keyinput_102), .C1(n6977), .C2(
        keyinput_99), .A(n10227), .ZN(n10229) );
  NOR3_X1 U11018 ( .A1(n10231), .A2(n10230), .A3(n10229), .ZN(n10232) );
  AOI221_X1 U11019 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_103), .C1(
        n10234), .C2(n10233), .A(n10232), .ZN(n10235) );
  AOI221_X1 U11020 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n10236), .C1(n7084), 
        .C2(keyinput_104), .A(n10235), .ZN(n10237) );
  AOI221_X1 U11021 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_105), .C1(
        n10239), .C2(n10238), .A(n10237), .ZN(n10247) );
  AOI22_X1 U11022 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_107), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput_106), .ZN(n10240) );
  OAI221_X1 U11023 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_107), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_106), .A(n10240), .ZN(n10246)
         );
  OAI22_X1 U11024 ( .A1(n10242), .A2(keyinput_110), .B1(keyinput_108), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n10241) );
  AOI221_X1 U11025 ( .B1(n10242), .B2(keyinput_110), .C1(
        P2_REG3_REG_1__SCAN_IN), .C2(keyinput_108), .A(n10241), .ZN(n10245) );
  OAI22_X1 U11026 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_111), .B1(
        P2_REG3_REG_21__SCAN_IN), .B2(keyinput_109), .ZN(n10243) );
  AOI221_X1 U11027 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_111), .C1(
        keyinput_109), .C2(P2_REG3_REG_21__SCAN_IN), .A(n10243), .ZN(n10244)
         );
  OAI211_X1 U11028 ( .C1(n10247), .C2(n10246), .A(n10245), .B(n10244), .ZN(
        n10248) );
  NAND4_X1 U11029 ( .A1(n10251), .A2(n10250), .A3(n10249), .A4(n10248), .ZN(
        n10254) );
  INV_X1 U11030 ( .A(keyinput_118), .ZN(n10252) );
  MUX2_X1 U11031 ( .A(keyinput_118), .B(n10252), .S(P2_REG3_REG_0__SCAN_IN), 
        .Z(n10253) );
  NAND2_X1 U11032 ( .A1(n10254), .A2(n10253), .ZN(n10260) );
  OAI22_X1 U11033 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_119), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_122), .ZN(n10255) );
  AOI221_X1 U11034 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_119), .C1(
        keyinput_122), .C2(P2_REG3_REG_11__SCAN_IN), .A(n10255), .ZN(n10259)
         );
  INV_X1 U11035 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10257) );
  OAI22_X1 U11036 ( .A1(n10257), .A2(keyinput_121), .B1(n6981), .B2(
        keyinput_120), .ZN(n10256) );
  AOI221_X1 U11037 ( .B1(n10257), .B2(keyinput_121), .C1(keyinput_120), .C2(
        n6981), .A(n10256), .ZN(n10258) );
  NAND3_X1 U11038 ( .A1(n10260), .A2(n10259), .A3(n10258), .ZN(n10261) );
  OAI221_X1 U11039 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_123), .C1(
        n10263), .C2(n10262), .A(n10261), .ZN(n10267) );
  AOI22_X1 U11040 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_125), .B1(n10265), .B2(keyinput_126), .ZN(n10264) );
  OAI221_X1 U11041 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_125), .C1(
        n10265), .C2(keyinput_126), .A(n10264), .ZN(n10266) );
  AOI21_X1 U11042 ( .B1(n10268), .B2(n10267), .A(n10266), .ZN(n10270) );
  NAND2_X1 U11043 ( .A1(keyinput_63), .A2(n6983), .ZN(n10269) );
  OAI221_X1 U11044 ( .B1(n10271), .B2(n10270), .C1(keyinput_63), .C2(n6983), 
        .A(n10269), .ZN(n10272) );
  AOI21_X1 U11045 ( .B1(n10274), .B2(n10273), .A(n10272), .ZN(n10275) );
  XNOR2_X1 U11046 ( .A(n10276), .B(n10275), .ZN(P1_U3325) );
  OAI222_X1 U11047 ( .A1(P1_U3086), .A2(n10279), .B1(n10284), .B2(n10278), 
        .C1(n10277), .C2(n8002), .ZN(P1_U3326) );
  OAI222_X1 U11048 ( .A1(P1_U3086), .A2(n10282), .B1(n8002), .B2(n10281), .C1(
        n10280), .C2(n10285), .ZN(P1_U3327) );
  OAI222_X1 U11049 ( .A1(P1_U3086), .A2(n10348), .B1(n10284), .B2(n6258), .C1(
        n10283), .C2(n8002), .ZN(P1_U3328) );
  OAI222_X1 U11050 ( .A1(n10287), .A2(P1_U3086), .B1(n8002), .B2(n10286), .C1(
        n10285), .C2(n6234), .ZN(P1_U3329) );
  MUX2_X1 U11051 ( .A(n10288), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U11052 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n4930), .ZN(P1_U3323) );
  AND2_X1 U11053 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n4930), .ZN(P1_U3322) );
  AND2_X1 U11054 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n4930), .ZN(P1_U3321) );
  AND2_X1 U11055 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n4930), .ZN(P1_U3320) );
  AND2_X1 U11056 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n4930), .ZN(P1_U3319) );
  AND2_X1 U11057 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n4930), .ZN(P1_U3318) );
  AND2_X1 U11058 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n4930), .ZN(P1_U3317) );
  AND2_X1 U11059 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n4930), .ZN(P1_U3316) );
  AND2_X1 U11060 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n4930), .ZN(P1_U3315) );
  AND2_X1 U11061 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n4930), .ZN(P1_U3314) );
  AND2_X1 U11062 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n4930), .ZN(P1_U3313) );
  AND2_X1 U11063 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n4930), .ZN(P1_U3312) );
  AND2_X1 U11064 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n4930), .ZN(P1_U3311) );
  AND2_X1 U11065 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n4930), .ZN(P1_U3310) );
  AND2_X1 U11066 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n4930), .ZN(P1_U3309) );
  AND2_X1 U11067 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n4930), .ZN(P1_U3308) );
  AND2_X1 U11068 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n4930), .ZN(P1_U3307) );
  AND2_X1 U11069 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n4930), .ZN(P1_U3306) );
  AND2_X1 U11070 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n4930), .ZN(P1_U3305) );
  AND2_X1 U11071 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n4930), .ZN(P1_U3304) );
  AND2_X1 U11072 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n4930), .ZN(P1_U3303) );
  AND2_X1 U11073 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n4930), .ZN(P1_U3302) );
  AND2_X1 U11074 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n4930), .ZN(P1_U3301) );
  AND2_X1 U11075 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n4930), .ZN(P1_U3300) );
  AND2_X1 U11076 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n4930), .ZN(P1_U3299) );
  AND2_X1 U11077 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n4930), .ZN(P1_U3298) );
  AND2_X1 U11078 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n4930), .ZN(P1_U3297) );
  AND2_X1 U11079 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n4930), .ZN(P1_U3296) );
  AND2_X1 U11080 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n4930), .ZN(P1_U3295) );
  AND2_X1 U11081 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n4930), .ZN(P1_U3294) );
  XOR2_X1 U11082 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  INV_X1 U11083 ( .A(n10292), .ZN(n10291) );
  OAI222_X1 U11084 ( .A1(n10294), .A2(n10293), .B1(n10294), .B2(n10292), .C1(
        n10291), .C2(n10290), .ZN(ADD_1068_U5) );
  AOI21_X1 U11085 ( .B1(n10297), .B2(n10296), .A(n10295), .ZN(ADD_1068_U54) );
  AOI21_X1 U11086 ( .B1(n10300), .B2(n10299), .A(n10298), .ZN(ADD_1068_U53) );
  OAI21_X1 U11087 ( .B1(n10303), .B2(n10302), .A(n10301), .ZN(ADD_1068_U52) );
  OAI21_X1 U11088 ( .B1(n10306), .B2(n10305), .A(n10304), .ZN(ADD_1068_U51) );
  OAI21_X1 U11089 ( .B1(n10309), .B2(n10308), .A(n10307), .ZN(ADD_1068_U50) );
  OAI21_X1 U11090 ( .B1(n10312), .B2(n10311), .A(n10310), .ZN(ADD_1068_U49) );
  OAI21_X1 U11091 ( .B1(n10315), .B2(n10314), .A(n10313), .ZN(ADD_1068_U48) );
  OAI21_X1 U11092 ( .B1(n10318), .B2(n10317), .A(n10316), .ZN(ADD_1068_U47) );
  OAI21_X1 U11093 ( .B1(n10321), .B2(n10320), .A(n10319), .ZN(ADD_1068_U63) );
  OAI21_X1 U11094 ( .B1(n10324), .B2(n10323), .A(n10322), .ZN(ADD_1068_U62) );
  OAI21_X1 U11095 ( .B1(n10327), .B2(n10326), .A(n10325), .ZN(ADD_1068_U61) );
  OAI21_X1 U11096 ( .B1(n10330), .B2(n10329), .A(n10328), .ZN(ADD_1068_U60) );
  OAI21_X1 U11097 ( .B1(n10333), .B2(n10332), .A(n10331), .ZN(ADD_1068_U59) );
  OAI21_X1 U11098 ( .B1(n10336), .B2(n10335), .A(n10334), .ZN(ADD_1068_U58) );
  OAI21_X1 U11099 ( .B1(n10339), .B2(n10338), .A(n10337), .ZN(ADD_1068_U57) );
  OAI21_X1 U11100 ( .B1(n10342), .B2(n10341), .A(n10340), .ZN(ADD_1068_U56) );
  OAI21_X1 U11101 ( .B1(n10345), .B2(n10344), .A(n10343), .ZN(ADD_1068_U55) );
  NAND2_X1 U11102 ( .A1(n10348), .A2(n10534), .ZN(n10346) );
  OAI211_X1 U11103 ( .C1(P1_REG2_REG_0__SCAN_IN), .C2(n10348), .A(n10347), .B(
        n10346), .ZN(n10349) );
  XOR2_X1 U11104 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10349), .Z(n10352) );
  AOI22_X1 U11105 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10350), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10351) );
  OAI21_X1 U11106 ( .B1(n10353), .B2(n10352), .A(n10351), .ZN(P1_U3243) );
  INV_X1 U11107 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10369) );
  OAI21_X1 U11108 ( .B1(n10356), .B2(n10355), .A(n10354), .ZN(n10365) );
  AOI21_X1 U11109 ( .B1(n10359), .B2(n10358), .A(n10357), .ZN(n10363) );
  OAI22_X1 U11110 ( .A1(n10363), .A2(n10362), .B1(n10361), .B2(n10360), .ZN(
        n10364) );
  AOI21_X1 U11111 ( .B1(n10366), .B2(n10365), .A(n10364), .ZN(n10368) );
  OAI211_X1 U11112 ( .C1(n10370), .C2(n10369), .A(n10368), .B(n10367), .ZN(
        P1_U3255) );
  AOI22_X1 U11113 ( .A1(n10476), .A2(n10371), .B1(n10498), .B2(
        P2_ADDR_REG_11__SCAN_IN), .ZN(n10387) );
  OAI21_X1 U11114 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n10373), .A(n10372), 
        .ZN(n10378) );
  OAI21_X1 U11115 ( .B1(n10376), .B2(n10375), .A(n10374), .ZN(n10377) );
  AOI22_X1 U11116 ( .A1(n10378), .A2(n10483), .B1(n10513), .B2(n10377), .ZN(
        n10386) );
  INV_X1 U11117 ( .A(n10379), .ZN(n10385) );
  AOI21_X1 U11118 ( .B1(n10382), .B2(n10381), .A(n10380), .ZN(n10383) );
  OR2_X1 U11119 ( .A1(n10489), .A2(n10383), .ZN(n10384) );
  NAND4_X1 U11120 ( .A1(n10387), .A2(n10386), .A3(n10385), .A4(n10384), .ZN(
        P2_U3193) );
  AOI22_X1 U11121 ( .A1(n10476), .A2(n10388), .B1(n10498), .B2(
        P2_ADDR_REG_12__SCAN_IN), .ZN(n10405) );
  OAI21_X1 U11122 ( .B1(n10391), .B2(n10390), .A(n10389), .ZN(n10396) );
  OAI21_X1 U11123 ( .B1(n10394), .B2(n10393), .A(n10392), .ZN(n10395) );
  AOI22_X1 U11124 ( .A1(n10396), .A2(n10483), .B1(n10513), .B2(n10395), .ZN(
        n10404) );
  INV_X1 U11125 ( .A(n10397), .ZN(n10403) );
  AOI21_X1 U11126 ( .B1(n10400), .B2(n10399), .A(n10398), .ZN(n10401) );
  OR2_X1 U11127 ( .A1(n10401), .A2(n10489), .ZN(n10402) );
  NAND4_X1 U11128 ( .A1(n10405), .A2(n10404), .A3(n10403), .A4(n10402), .ZN(
        P2_U3194) );
  AOI22_X1 U11129 ( .A1(n10476), .A2(n10406), .B1(n10498), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n10422) );
  OAI21_X1 U11130 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n10408), .A(n10407), 
        .ZN(n10413) );
  OAI21_X1 U11131 ( .B1(n10411), .B2(n10410), .A(n10409), .ZN(n10412) );
  AOI22_X1 U11132 ( .A1(n10413), .A2(n10483), .B1(n10513), .B2(n10412), .ZN(
        n10421) );
  INV_X1 U11133 ( .A(n10414), .ZN(n10420) );
  AOI21_X1 U11134 ( .B1(n10417), .B2(n10416), .A(n10415), .ZN(n10418) );
  OR2_X1 U11135 ( .A1(n10489), .A2(n10418), .ZN(n10419) );
  NAND4_X1 U11136 ( .A1(n10422), .A2(n10421), .A3(n10420), .A4(n10419), .ZN(
        P2_U3195) );
  AOI22_X1 U11137 ( .A1(n10476), .A2(n10423), .B1(n10498), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n10439) );
  OAI21_X1 U11138 ( .B1(n10426), .B2(n10425), .A(n10424), .ZN(n10431) );
  OAI21_X1 U11139 ( .B1(n10429), .B2(n10428), .A(n10427), .ZN(n10430) );
  AOI22_X1 U11140 ( .A1(n10431), .A2(n10483), .B1(n10513), .B2(n10430), .ZN(
        n10438) );
  NAND2_X1 U11141 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n10437)
         );
  AOI21_X1 U11142 ( .B1(n10434), .B2(n10433), .A(n10432), .ZN(n10435) );
  OR2_X1 U11143 ( .A1(n10435), .A2(n10489), .ZN(n10436) );
  NAND4_X1 U11144 ( .A1(n10439), .A2(n10438), .A3(n10437), .A4(n10436), .ZN(
        P2_U3196) );
  AOI22_X1 U11145 ( .A1(n10476), .A2(n10440), .B1(n10498), .B2(
        P2_ADDR_REG_15__SCAN_IN), .ZN(n10456) );
  OAI21_X1 U11146 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n10442), .A(n10441), 
        .ZN(n10447) );
  OAI21_X1 U11147 ( .B1(n10445), .B2(n10444), .A(n10443), .ZN(n10446) );
  AOI22_X1 U11148 ( .A1(n10447), .A2(n10483), .B1(n10513), .B2(n10446), .ZN(
        n10455) );
  INV_X1 U11149 ( .A(n10448), .ZN(n10454) );
  AOI21_X1 U11150 ( .B1(n10451), .B2(n10450), .A(n10449), .ZN(n10452) );
  OR2_X1 U11151 ( .A1(n10489), .A2(n10452), .ZN(n10453) );
  NAND4_X1 U11152 ( .A1(n10456), .A2(n10455), .A3(n10454), .A4(n10453), .ZN(
        P2_U3197) );
  AOI22_X1 U11153 ( .A1(n10476), .A2(n10457), .B1(n10498), .B2(
        P2_ADDR_REG_16__SCAN_IN), .ZN(n10474) );
  OAI21_X1 U11154 ( .B1(n10460), .B2(n10459), .A(n10458), .ZN(n10465) );
  OAI21_X1 U11155 ( .B1(n10463), .B2(n10462), .A(n10461), .ZN(n10464) );
  AOI22_X1 U11156 ( .A1(n10465), .A2(n10483), .B1(n10513), .B2(n10464), .ZN(
        n10473) );
  INV_X1 U11157 ( .A(n10466), .ZN(n10472) );
  AOI21_X1 U11158 ( .B1(n10469), .B2(n10468), .A(n10467), .ZN(n10470) );
  OR2_X1 U11159 ( .A1(n10470), .A2(n10489), .ZN(n10471) );
  NAND4_X1 U11160 ( .A1(n10474), .A2(n10473), .A3(n10472), .A4(n10471), .ZN(
        P2_U3198) );
  AOI22_X1 U11161 ( .A1(n10476), .A2(n10475), .B1(n10498), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n10493) );
  OAI21_X1 U11162 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n10478), .A(n10477), 
        .ZN(n10484) );
  OAI21_X1 U11163 ( .B1(n10481), .B2(n10480), .A(n10479), .ZN(n10482) );
  AOI22_X1 U11164 ( .A1(n10484), .A2(n10483), .B1(n10513), .B2(n10482), .ZN(
        n10492) );
  INV_X1 U11165 ( .A(n10485), .ZN(n10491) );
  AOI21_X1 U11166 ( .B1(n10487), .B2(n10486), .A(n10504), .ZN(n10488) );
  OR2_X1 U11167 ( .A1(n10489), .A2(n10488), .ZN(n10490) );
  NAND4_X1 U11168 ( .A1(n10493), .A2(n10492), .A3(n10491), .A4(n10490), .ZN(
        P2_U3199) );
  INV_X1 U11169 ( .A(n10499), .ZN(n10501) );
  NAND2_X1 U11170 ( .A1(n10501), .A2(n10500), .ZN(n10514) );
  OAI21_X1 U11171 ( .B1(n10514), .B2(n10503), .A(n10502), .ZN(n10511) );
  NOR2_X1 U11172 ( .A1(n10505), .A2(n10504), .ZN(n10506) );
  XNOR2_X1 U11173 ( .A(n10507), .B(n10506), .ZN(n10508) );
  AOI22_X1 U11174 ( .A1(n10511), .A2(n10510), .B1(n10509), .B2(n10508), .ZN(
        n10516) );
  NAND3_X1 U11175 ( .A1(n10514), .A2(n10513), .A3(n10512), .ZN(n10515) );
  NAND3_X1 U11176 ( .A1(n10517), .A2(n10516), .A3(n10515), .ZN(P2_U3200) );
  XNOR2_X1 U11177 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NOR3_X1 U11178 ( .A1(n10527), .A2(n10518), .A3(n10532), .ZN(n10524) );
  AND2_X1 U11179 ( .A1(n5664), .A2(n10519), .ZN(n10531) );
  NAND3_X1 U11180 ( .A1(n10533), .A2(n10532), .A3(n9288), .ZN(n10520) );
  OAI21_X1 U11181 ( .B1(n10522), .B2(n10521), .A(n10520), .ZN(n10523) );
  NOR3_X1 U11182 ( .A1(n10524), .A2(n10531), .A3(n10523), .ZN(n10526) );
  AOI22_X1 U11183 ( .A1(n9685), .A2(n5619), .B1(n10526), .B2(n10525), .ZN(
        P1_U3293) );
  AOI21_X1 U11184 ( .B1(n10529), .B2(n10528), .A(n10527), .ZN(n10530) );
  AOI211_X1 U11185 ( .C1(n10533), .C2(n10532), .A(n10531), .B(n10530), .ZN(
        n10536) );
  AOI22_X1 U11186 ( .A1(n10736), .A2(n10536), .B1(n10534), .B2(n10735), .ZN(
        P1_U3522) );
  INV_X1 U11187 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U11188 ( .A1(n10740), .A2(n10536), .B1(n10535), .B2(n10737), .ZN(
        P1_U3453) );
  NAND2_X1 U11189 ( .A1(n6474), .A2(n10704), .ZN(n10538) );
  OAI211_X1 U11190 ( .C1(n10539), .C2(n10729), .A(n10538), .B(n10537), .ZN(
        n10540) );
  AOI21_X1 U11191 ( .B1(n10541), .B2(n10711), .A(n10540), .ZN(n10542) );
  AND2_X1 U11192 ( .A1(n10543), .A2(n10542), .ZN(n10546) );
  AOI22_X1 U11193 ( .A1(n10736), .A2(n10546), .B1(n10544), .B2(n10735), .ZN(
        P1_U3523) );
  INV_X1 U11194 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10545) );
  AOI22_X1 U11195 ( .A1(n10740), .A2(n10546), .B1(n10545), .B2(n10737), .ZN(
        P1_U3456) );
  OAI21_X1 U11196 ( .B1(n10548), .B2(n10729), .A(n10547), .ZN(n10550) );
  AOI211_X1 U11197 ( .C1(n10731), .C2(n10551), .A(n10550), .B(n10549), .ZN(
        n10554) );
  AOI22_X1 U11198 ( .A1(n10736), .A2(n10554), .B1(n10552), .B2(n10735), .ZN(
        P1_U3524) );
  INV_X1 U11199 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U11200 ( .A1(n10740), .A2(n10554), .B1(n10553), .B2(n10737), .ZN(
        P1_U3459) );
  OAI21_X1 U11201 ( .B1(n8337), .B2(n10557), .A(n10555), .ZN(n10575) );
  NOR2_X1 U11202 ( .A1(n10572), .A2(n10715), .ZN(n10567) );
  NAND3_X1 U11203 ( .A1(n10558), .A2(n10557), .A3(n10556), .ZN(n10559) );
  AND2_X1 U11204 ( .A1(n10560), .A2(n10559), .ZN(n10561) );
  OAI222_X1 U11205 ( .A1(n10566), .A2(n10565), .B1(n10564), .B2(n10563), .C1(
        n10562), .C2(n10561), .ZN(n10573) );
  AOI211_X1 U11206 ( .C1(n10720), .C2(n10575), .A(n10567), .B(n10573), .ZN(
        n10569) );
  AOI22_X1 U11207 ( .A1(n10723), .A2(n10569), .B1(n6500), .B2(n10721), .ZN(
        P2_U3461) );
  INV_X1 U11208 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U11209 ( .A1(n10727), .A2(n10569), .B1(n10568), .B2(n10724), .ZN(
        P2_U3396) );
  OAI22_X1 U11210 ( .A1(n10572), .A2(n10571), .B1(n10570), .B2(n10263), .ZN(
        n10574) );
  AOI211_X1 U11211 ( .C1(n10576), .C2(n10575), .A(n10574), .B(n10573), .ZN(
        n10578) );
  AOI22_X1 U11212 ( .A1(n10580), .A2(n10579), .B1(n10578), .B2(n10577), .ZN(
        P2_U3231) );
  INV_X1 U11213 ( .A(n10581), .ZN(n10585) );
  OAI22_X1 U11214 ( .A1(n10583), .A2(n10696), .B1(n10582), .B2(n10715), .ZN(
        n10584) );
  NOR2_X1 U11215 ( .A1(n10585), .A2(n10584), .ZN(n10588) );
  INV_X1 U11216 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10586) );
  AOI22_X1 U11217 ( .A1(n10723), .A2(n10588), .B1(n10586), .B2(n10721), .ZN(
        P2_U3462) );
  INV_X1 U11218 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10587) );
  AOI22_X1 U11219 ( .A1(n10727), .A2(n10588), .B1(n10587), .B2(n10724), .ZN(
        P2_U3399) );
  INV_X1 U11220 ( .A(n10589), .ZN(n10593) );
  OAI22_X1 U11221 ( .A1(n10591), .A2(n10696), .B1(n10590), .B2(n10715), .ZN(
        n10592) );
  NOR2_X1 U11222 ( .A1(n10593), .A2(n10592), .ZN(n10596) );
  AOI22_X1 U11223 ( .A1(n10723), .A2(n10596), .B1(n10594), .B2(n10721), .ZN(
        P2_U3463) );
  INV_X1 U11224 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10595) );
  AOI22_X1 U11225 ( .A1(n10727), .A2(n10596), .B1(n10595), .B2(n10724), .ZN(
        P2_U3402) );
  AOI22_X1 U11226 ( .A1(n10598), .A2(n10704), .B1(n10705), .B2(n10597), .ZN(
        n10600) );
  NAND3_X1 U11227 ( .A1(n10601), .A2(n10600), .A3(n10599), .ZN(n10602) );
  AOI21_X1 U11228 ( .B1(n10711), .B2(n10603), .A(n10602), .ZN(n10605) );
  AOI22_X1 U11229 ( .A1(n10736), .A2(n10605), .B1(n6646), .B2(n10735), .ZN(
        P1_U3526) );
  INV_X1 U11230 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10604) );
  AOI22_X1 U11231 ( .A1(n10740), .A2(n10605), .B1(n10604), .B2(n10737), .ZN(
        P1_U3465) );
  AND2_X1 U11232 ( .A1(n10606), .A2(n10711), .ZN(n10611) );
  OAI211_X1 U11233 ( .C1(n10609), .C2(n10631), .A(n10608), .B(n10607), .ZN(
        n10610) );
  NOR3_X1 U11234 ( .A1(n10612), .A2(n10611), .A3(n10610), .ZN(n10613) );
  AOI22_X1 U11235 ( .A1(n10736), .A2(n10613), .B1(n6647), .B2(n10735), .ZN(
        P1_U3527) );
  AOI22_X1 U11236 ( .A1(n10740), .A2(n10613), .B1(n5754), .B2(n10737), .ZN(
        P1_U3468) );
  NOR2_X1 U11237 ( .A1(n10614), .A2(n10715), .ZN(n10616) );
  AOI211_X1 U11238 ( .C1(n10720), .C2(n10617), .A(n10616), .B(n10615), .ZN(
        n10620) );
  AOI22_X1 U11239 ( .A1(n10723), .A2(n10620), .B1(n10618), .B2(n10721), .ZN(
        P2_U3465) );
  INV_X1 U11240 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U11241 ( .A1(n10727), .A2(n10620), .B1(n10619), .B2(n10724), .ZN(
        P2_U3408) );
  OAI21_X1 U11242 ( .B1(n10622), .B2(n10729), .A(n10621), .ZN(n10624) );
  AOI211_X1 U11243 ( .C1(n10711), .C2(n10625), .A(n10624), .B(n10623), .ZN(
        n10627) );
  AOI22_X1 U11244 ( .A1(n10736), .A2(n10627), .B1(n6666), .B2(n10735), .ZN(
        P1_U3528) );
  INV_X1 U11245 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10626) );
  AOI22_X1 U11246 ( .A1(n10740), .A2(n10627), .B1(n10626), .B2(n10737), .ZN(
        P1_U3471) );
  INV_X1 U11247 ( .A(n10628), .ZN(n10635) );
  OAI211_X1 U11248 ( .C1(n10632), .C2(n10631), .A(n10630), .B(n10629), .ZN(
        n10634) );
  AOI211_X1 U11249 ( .C1(n10731), .C2(n10635), .A(n10634), .B(n10633), .ZN(
        n10637) );
  AOI22_X1 U11250 ( .A1(n10736), .A2(n10637), .B1(n6663), .B2(n10735), .ZN(
        P1_U3529) );
  INV_X1 U11251 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10636) );
  AOI22_X1 U11252 ( .A1(n10740), .A2(n10637), .B1(n10636), .B2(n10737), .ZN(
        P1_U3474) );
  OAI22_X1 U11253 ( .A1(n10639), .A2(n10689), .B1(n10638), .B2(n10715), .ZN(
        n10640) );
  NOR2_X1 U11254 ( .A1(n10641), .A2(n10640), .ZN(n10644) );
  INV_X1 U11255 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10642) );
  AOI22_X1 U11256 ( .A1(n10723), .A2(n10644), .B1(n10642), .B2(n10721), .ZN(
        P2_U3466) );
  INV_X1 U11257 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10643) );
  AOI22_X1 U11258 ( .A1(n10727), .A2(n10644), .B1(n10643), .B2(n10724), .ZN(
        P2_U3411) );
  NAND2_X1 U11259 ( .A1(n10645), .A2(n10731), .ZN(n10647) );
  OAI211_X1 U11260 ( .C1(n10648), .C2(n10729), .A(n10647), .B(n10646), .ZN(
        n10649) );
  NOR2_X1 U11261 ( .A1(n10650), .A2(n10649), .ZN(n10653) );
  AOI22_X1 U11262 ( .A1(n10736), .A2(n10653), .B1(n10651), .B2(n10735), .ZN(
        P1_U3530) );
  INV_X1 U11263 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U11264 ( .A1(n10740), .A2(n10653), .B1(n10652), .B2(n10737), .ZN(
        P1_U3477) );
  OAI21_X1 U11265 ( .B1(n10655), .B2(n10715), .A(n10654), .ZN(n10656) );
  AOI21_X1 U11266 ( .B1(n10720), .B2(n10657), .A(n10656), .ZN(n10660) );
  AOI22_X1 U11267 ( .A1(n10723), .A2(n10660), .B1(n10658), .B2(n10721), .ZN(
        P2_U3467) );
  INV_X1 U11268 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10659) );
  AOI22_X1 U11269 ( .A1(n10727), .A2(n10660), .B1(n10659), .B2(n10724), .ZN(
        P2_U3414) );
  AOI22_X1 U11270 ( .A1(n10662), .A2(n10705), .B1(n10704), .B2(n10661), .ZN(
        n10663) );
  NAND3_X1 U11271 ( .A1(n10665), .A2(n10664), .A3(n10663), .ZN(n10666) );
  AOI21_X1 U11272 ( .B1(n10711), .B2(n10667), .A(n10666), .ZN(n10669) );
  AOI22_X1 U11273 ( .A1(n10736), .A2(n10669), .B1(n6699), .B2(n10735), .ZN(
        P1_U3531) );
  INV_X1 U11274 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U11275 ( .A1(n10740), .A2(n10669), .B1(n10668), .B2(n10737), .ZN(
        P1_U3480) );
  NAND2_X1 U11276 ( .A1(n10670), .A2(n10720), .ZN(n10674) );
  NAND2_X1 U11277 ( .A1(n10672), .A2(n10671), .ZN(n10673) );
  AOI22_X1 U11278 ( .A1(n10723), .A2(n10678), .B1(n10676), .B2(n10721), .ZN(
        P2_U3468) );
  INV_X1 U11279 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10677) );
  AOI22_X1 U11280 ( .A1(n10727), .A2(n10678), .B1(n10677), .B2(n10724), .ZN(
        P2_U3417) );
  AOI22_X1 U11281 ( .A1(n10680), .A2(n10705), .B1(n10704), .B2(n10679), .ZN(
        n10682) );
  NAND3_X1 U11282 ( .A1(n10683), .A2(n10682), .A3(n10681), .ZN(n10684) );
  AOI21_X1 U11283 ( .B1(n10711), .B2(n10685), .A(n10684), .ZN(n10687) );
  AOI22_X1 U11284 ( .A1(n10736), .A2(n10687), .B1(n6733), .B2(n10735), .ZN(
        P1_U3532) );
  INV_X1 U11285 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U11286 ( .A1(n10740), .A2(n10687), .B1(n10686), .B2(n10737), .ZN(
        P1_U3483) );
  OAI22_X1 U11287 ( .A1(n10690), .A2(n10689), .B1(n10688), .B2(n10715), .ZN(
        n10691) );
  NOR2_X1 U11288 ( .A1(n10692), .A2(n10691), .ZN(n10694) );
  AOI22_X1 U11289 ( .A1(n10723), .A2(n10694), .B1(n8746), .B2(n10721), .ZN(
        P2_U3469) );
  INV_X1 U11290 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U11291 ( .A1(n10727), .A2(n10694), .B1(n10693), .B2(n10724), .ZN(
        P2_U3420) );
  OAI22_X1 U11292 ( .A1(n10697), .A2(n10696), .B1(n10695), .B2(n10715), .ZN(
        n10698) );
  NOR2_X1 U11293 ( .A1(n10699), .A2(n10698), .ZN(n10702) );
  AOI22_X1 U11294 ( .A1(n10723), .A2(n10702), .B1(n10700), .B2(n10721), .ZN(
        P2_U3471) );
  INV_X1 U11295 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10701) );
  AOI22_X1 U11296 ( .A1(n10727), .A2(n10702), .B1(n10701), .B2(n10724), .ZN(
        P2_U3426) );
  AOI22_X1 U11297 ( .A1(n10706), .A2(n10705), .B1(n10704), .B2(n10703), .ZN(
        n10708) );
  NAND3_X1 U11298 ( .A1(n10709), .A2(n10708), .A3(n10707), .ZN(n10710) );
  AOI21_X1 U11299 ( .B1(n10712), .B2(n10711), .A(n10710), .ZN(n10714) );
  AOI22_X1 U11300 ( .A1(n10736), .A2(n10714), .B1(n5932), .B2(n10735), .ZN(
        P1_U3534) );
  INV_X1 U11301 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10713) );
  AOI22_X1 U11302 ( .A1(n10740), .A2(n10714), .B1(n10713), .B2(n10737), .ZN(
        P1_U3489) );
  NOR2_X1 U11303 ( .A1(n10716), .A2(n10715), .ZN(n10718) );
  AOI211_X1 U11304 ( .C1(n10720), .C2(n10719), .A(n10718), .B(n10717), .ZN(
        n10726) );
  INV_X1 U11305 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10722) );
  AOI22_X1 U11306 ( .A1(n10723), .A2(n10726), .B1(n10722), .B2(n10721), .ZN(
        P2_U3472) );
  INV_X1 U11307 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10725) );
  AOI22_X1 U11308 ( .A1(n10727), .A2(n10726), .B1(n10725), .B2(n10724), .ZN(
        P2_U3429) );
  OAI21_X1 U11309 ( .B1(n7969), .B2(n10729), .A(n10728), .ZN(n10730) );
  AOI21_X1 U11310 ( .B1(n10732), .B2(n10731), .A(n10730), .ZN(n10733) );
  AND2_X1 U11311 ( .A1(n10734), .A2(n10733), .ZN(n10739) );
  AOI22_X1 U11312 ( .A1(n10736), .A2(n10739), .B1(n7617), .B2(n10735), .ZN(
        P1_U3536) );
  INV_X1 U11313 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10738) );
  AOI22_X1 U11314 ( .A1(n10740), .A2(n10739), .B1(n10738), .B2(n10737), .ZN(
        P1_U3495) );
  XNOR2_X1 U11315 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  CLKBUF_X1 U5003 ( .A(n5735), .Z(n9296) );
  CLKBUF_X1 U5011 ( .A(n5755), .Z(n6448) );
  CLKBUF_X2 U5013 ( .A(n5648), .Z(n5086) );
  CLKBUF_X1 U5068 ( .A(n5751), .Z(n6337) );
  AND2_X1 U6210 ( .A1(n10043), .A2(n10042), .ZN(n10744) );
endmodule

