

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658;

  NAND2_X1 U2240 ( .A1(n2063), .A2(n2064), .ZN(n3639) );
  NAND2_X1 U2241 ( .A1(n2960), .A2(n2959), .ZN(n4086) );
  NAND2_X1 U2242 ( .A1(n2084), .A2(n2034), .ZN(n4367) );
  INV_X4 U2243 ( .A(n2726), .ZN(n2813) );
  NAND3_X1 U2244 ( .A1(n2164), .A2(n2165), .A3(n2021), .ZN(n2170) );
  INV_X1 U2245 ( .A(n2367), .ZN(n2538) );
  INV_X2 U2246 ( .A(n2726), .ZN(n2769) );
  AND2_X1 U2247 ( .A1(n3126), .A2(n2810), .ZN(n2674) );
  OAI22_X2 U2248 ( .A1(n3297), .A2(n2927), .B1(n2926), .B2(n3310), .ZN(n3109)
         );
  OAI21_X1 U2249 ( .B1(n4086), .B2(n2962), .A(n2961), .ZN(n4068) );
  CLKBUF_X2 U2250 ( .A(n2399), .Z(n2453) );
  AND2_X1 U2251 ( .A1(n2312), .A2(n4570), .ZN(n3020) );
  NAND2_X1 U2252 ( .A1(n2293), .A2(IR_REG_31__SCAN_IN), .ZN(n2294) );
  INV_X2 U2253 ( .A(n2879), .ZN(n4461) );
  XNOR2_X2 U2254 ( .A(n2841), .B(n3062), .ZN(n3056) );
  NAND4_X2 U2255 ( .A1(n2403), .A2(n2402), .A3(n2401), .A4(n2400), .ZN(n3934)
         );
  XNOR2_X2 U2256 ( .A(n2294), .B(IR_REG_24__SCAN_IN), .ZN(n2775) );
  OAI211_X2 U2258 ( .C1(IR_REG_1__SCAN_IN), .C2(IR_REG_31__SCAN_IN), .A(n2160), 
        .B(n2159), .ZN(n2880) );
  OAI21_X1 U2259 ( .B1(n4068), .B2(n2964), .A(n2963), .ZN(n4049) );
  NAND2_X2 U2260 ( .A1(n2920), .A2(n2336), .ZN(n2970) );
  NAND4_X1 U2261 ( .A1(n2423), .A2(n2422), .A3(n2421), .A4(n2420), .ZN(n3933)
         );
  INV_X2 U2262 ( .A(n2921), .ZN(n2920) );
  XNOR2_X1 U2264 ( .A(n2319), .B(n2318), .ZN(n2322) );
  INV_X2 U2265 ( .A(IR_REG_31__SCAN_IN), .ZN(n3033) );
  MUX2_X1 U2266 ( .A(REG1_REG_28__SCAN_IN), .B(n3024), .S(n4658), .Z(n3014) );
  MUX2_X1 U2267 ( .A(REG0_REG_28__SCAN_IN), .B(n3024), .S(n4647), .Z(n3025) );
  AOI21_X1 U2268 ( .B1(n2153), .B2(n2011), .A(n2152), .ZN(n3984) );
  AND2_X1 U2269 ( .A1(n4030), .A2(n4040), .ZN(n4032) );
  AND2_X1 U2270 ( .A1(n3969), .A2(n2862), .ZN(n2863) );
  NOR2_X1 U2271 ( .A1(n4012), .A2(n2095), .ZN(n4303) );
  AND2_X1 U2272 ( .A1(n4013), .A2(n4021), .ZN(n2095) );
  NAND2_X1 U2273 ( .A1(n2951), .A2(n2950), .ZN(n4229) );
  NAND2_X1 U2274 ( .A1(n4496), .A2(n2057), .ZN(n3966) );
  NOR2_X1 U2275 ( .A1(n4484), .A2(n4483), .ZN(n4482) );
  OAI21_X1 U2276 ( .B1(n3181), .B2(n2139), .A(n2135), .ZN(n3263) );
  NAND2_X1 U2277 ( .A1(n2208), .A2(n2206), .ZN(n3368) );
  INV_X1 U2278 ( .A(n3402), .ZN(n2084) );
  NAND3_X1 U2279 ( .A1(n2127), .A2(n2130), .A3(n3792), .ZN(n3331) );
  OAI22_X1 U2280 ( .A1(n3091), .A2(n3257), .B1(n4456), .B2(n2894), .ZN(n3100)
         );
  XNOR2_X1 U2281 ( .A(n2893), .B(n4457), .ZN(n3091) );
  INV_X2 U2282 ( .A(n4581), .ZN(n1998) );
  OAI21_X1 U2283 ( .B1(n2818), .B2(n4563), .A(n4276), .ZN(n3724) );
  AND2_X1 U2284 ( .A1(n3225), .A2(n3342), .ZN(n4636) );
  INV_X1 U2285 ( .A(n2968), .ZN(n4555) );
  AND2_X1 U2286 ( .A1(n2144), .A2(n2143), .ZN(n2889) );
  CLKBUF_X1 U2287 ( .A(n2367), .Z(n2768) );
  INV_X2 U2288 ( .A(n2674), .ZN(n2770) );
  INV_X1 U2289 ( .A(n4562), .ZN(n2336) );
  CLKBUF_X1 U2290 ( .A(n2349), .Z(n3027) );
  AND2_X1 U2291 ( .A1(n2844), .A2(n4474), .ZN(n2845) );
  NAND2_X1 U2292 ( .A1(n3934), .A2(n3117), .ZN(n3779) );
  CLKBUF_X1 U2293 ( .A(n2439), .Z(n2764) );
  NAND2_X1 U2294 ( .A1(n2325), .A2(n2322), .ZN(n2439) );
  NAND2_X1 U2295 ( .A1(n2323), .A2(n2322), .ZN(n2377) );
  OAI21_X1 U2296 ( .B1(n2313), .B2(IR_REG_22__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2794) );
  AND2_X1 U2297 ( .A1(n2292), .A2(n2313), .ZN(n4452) );
  NAND2_X1 U2298 ( .A1(n2839), .A2(n2838), .ZN(n3959) );
  INV_X1 U2299 ( .A(n2322), .ZN(n3037) );
  NAND2_X1 U2300 ( .A1(n2826), .A2(IR_REG_31__SCAN_IN), .ZN(n2875) );
  NAND2_X1 U2301 ( .A1(n3034), .A2(IR_REG_31__SCAN_IN), .ZN(n2316) );
  AND4_X1 U2302 ( .A1(n2303), .A2(n2272), .A3(n2082), .A4(n2083), .ZN(n2317)
         );
  CLKBUF_X1 U2303 ( .A(n2303), .Z(n2297) );
  OAI211_X1 U2304 ( .C1(n2174), .C2(n2368), .A(n2173), .B(n2172), .ZN(n2879)
         );
  INV_X1 U2305 ( .A(IR_REG_23__SCAN_IN), .ZN(n2793) );
  NOR2_X1 U2306 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2284)
         );
  NOR2_X1 U2307 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2275)
         );
  NOR2_X1 U2308 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2274)
         );
  NOR2_X1 U2309 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2273)
         );
  INV_X1 U2310 ( .A(IR_REG_21__SCAN_IN), .ZN(n2290) );
  NOR2_X1 U2311 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2266)
         );
  NOR2_X1 U2312 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2285)
         );
  NOR2_X2 U2313 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2368)
         );
  OAI22_X2 U2314 ( .A1(n3458), .A2(n3459), .B1(n2649), .B2(n2650), .ZN(n3695)
         );
  INV_X4 U2315 ( .A(n2000), .ZN(n2447) );
  NAND4_X4 U2316 ( .A1(n2329), .A2(n2328), .A3(n2327), .A4(n2326), .ZN(n2921)
         );
  OR2_X2 U2317 ( .A1(n2000), .A2(n2324), .ZN(n2327) );
  OAI211_X1 U2318 ( .C1(n2875), .C2(IR_REG_28__SCAN_IN), .A(n2331), .B(n2330), 
        .ZN(n2332) );
  BUF_X4 U2319 ( .A(n2377), .Z(n2000) );
  NAND2_X2 U2320 ( .A1(n2974), .A2(n3781), .ZN(n3181) );
  INV_X1 U2321 ( .A(n3722), .ZN(n2066) );
  INV_X1 U2322 ( .A(n2110), .ZN(n2108) );
  OAI21_X1 U2323 ( .B1(n2197), .B2(n2195), .A(n2041), .ZN(n2194) );
  INV_X1 U2324 ( .A(n2954), .ZN(n2195) );
  INV_X1 U2325 ( .A(IR_REG_22__SCAN_IN), .ZN(n2295) );
  NAND2_X1 U2326 ( .A1(n3959), .A2(n2840), .ZN(n2841) );
  OR2_X1 U2327 ( .A1(n4518), .A2(n2904), .ZN(n2905) );
  NAND2_X1 U2328 ( .A1(n4036), .A2(n4010), .ZN(n4015) );
  AND2_X1 U2329 ( .A1(n2203), .A2(n2202), .ZN(n2214) );
  AND2_X1 U2330 ( .A1(n2940), .A2(n2023), .ZN(n2202) );
  INV_X1 U2331 ( .A(n2217), .ZN(n2213) );
  NAND2_X1 U2332 ( .A1(n2312), .A2(n4452), .ZN(n3126) );
  INV_X1 U2333 ( .A(IR_REG_18__SCAN_IN), .ZN(n2283) );
  INV_X1 U2334 ( .A(IR_REG_17__SCAN_IN), .ZN(n2282) );
  AOI21_X1 U2335 ( .B1(n2065), .B2(n2243), .A(n2043), .ZN(n2064) );
  OR2_X1 U2336 ( .A1(n2718), .A2(n3645), .ZN(n2738) );
  INV_X1 U2337 ( .A(n2437), .ZN(n2820) );
  NAND2_X1 U2338 ( .A1(n4472), .A2(n2168), .ZN(n2164) );
  NOR2_X1 U2339 ( .A1(n3085), .A2(n4471), .ZN(n2168) );
  NAND2_X1 U2340 ( .A1(n2845), .A2(n2166), .ZN(n2165) );
  INV_X1 U2341 ( .A(n3085), .ZN(n2166) );
  INV_X1 U2342 ( .A(IR_REG_7__SCAN_IN), .ZN(n2473) );
  AOI21_X1 U2343 ( .B1(n3203), .B2(n3204), .A(n2141), .ZN(n2898) );
  NOR2_X1 U2344 ( .A1(n3207), .A2(n3554), .ZN(n2141) );
  XNOR2_X1 U2345 ( .A(n2905), .B(n4597), .ZN(n4529) );
  NAND2_X1 U2346 ( .A1(n4529), .A2(n4528), .ZN(n4527) );
  NAND2_X1 U2347 ( .A1(n2119), .A2(n4032), .ZN(n2117) );
  NOR2_X1 U2348 ( .A1(n4307), .A2(n2124), .ZN(n2119) );
  OR2_X1 U2349 ( .A1(n2760), .A2(n2819), .ZN(n4025) );
  NAND3_X1 U2350 ( .A1(n2222), .A2(n2223), .A3(n2224), .ZN(n4009) );
  NAND2_X1 U2351 ( .A1(n2226), .A2(n2037), .ZN(n2223) );
  AOI21_X1 U2352 ( .B1(n2226), .B2(n2225), .A(n2036), .ZN(n2224) );
  OR2_X1 U2353 ( .A1(n2738), .A2(n3743), .ZN(n2750) );
  NOR2_X1 U2354 ( .A1(n2230), .A2(n2040), .ZN(n2229) );
  NAND2_X1 U2355 ( .A1(n2963), .A2(n2964), .ZN(n2221) );
  AOI21_X1 U2356 ( .B1(n2001), .B2(n2189), .A(n2033), .ZN(n2188) );
  INV_X1 U2357 ( .A(n2268), .ZN(n2189) );
  INV_X1 U2358 ( .A(n4144), .ZN(n2191) );
  NAND2_X1 U2359 ( .A1(n3117), .A2(n3221), .ZN(n2085) );
  NAND2_X1 U2360 ( .A1(n4015), .A2(n3828), .ZN(n3898) );
  NOR2_X1 U2361 ( .A1(n2111), .A2(n4256), .ZN(n2110) );
  NOR2_X1 U2362 ( .A1(n2114), .A2(n2112), .ZN(n2111) );
  INV_X1 U2363 ( .A(n2969), .ZN(n2354) );
  OR2_X2 U2364 ( .A1(n3126), .A2(n2335), .ZN(n2397) );
  OR2_X1 U2365 ( .A1(n3982), .A2(n2816), .ZN(n2810) );
  AND2_X1 U2366 ( .A1(n4075), .A2(n4061), .ZN(n3841) );
  INV_X1 U2367 ( .A(n2323), .ZN(n2325) );
  NAND2_X1 U2368 ( .A1(n2843), .A2(n2842), .ZN(n2844) );
  NOR2_X1 U2369 ( .A1(n2227), .A2(n2966), .ZN(n2226) );
  INV_X1 U2370 ( .A(n2229), .ZN(n2227) );
  OR2_X1 U2371 ( .A1(n4149), .A2(n4139), .ZN(n4111) );
  OR2_X1 U2372 ( .A1(n4166), .A2(n4193), .ZN(n4160) );
  OR2_X1 U2373 ( .A1(n3185), .A2(n3931), .ZN(n3782) );
  INV_X1 U2374 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2435) );
  NAND2_X1 U2375 ( .A1(REG3_REG_5__SCAN_IN), .A2(REG3_REG_6__SCAN_IN), .ZN(
        n2103) );
  INV_X1 U2376 ( .A(n3779), .ZN(n2133) );
  INV_X1 U2377 ( .A(n2417), .ZN(n2415) );
  NAND2_X1 U2378 ( .A1(n3775), .A2(n3776), .ZN(n2131) );
  AND2_X1 U2379 ( .A1(n4451), .A2(n4452), .ZN(n3003) );
  NOR2_X1 U2380 ( .A1(n3188), .A2(n3254), .ZN(n2096) );
  INV_X1 U2381 ( .A(n3336), .ZN(n3342) );
  INV_X1 U2382 ( .A(n4451), .ZN(n2816) );
  INV_X1 U2383 ( .A(IR_REG_27__SCAN_IN), .ZN(n2874) );
  AND2_X1 U2384 ( .A1(n2297), .A2(n2296), .ZN(n2299) );
  INV_X1 U2385 ( .A(IR_REG_13__SCAN_IN), .ZN(n3491) );
  INV_X1 U2386 ( .A(n2384), .ZN(n2272) );
  INV_X1 U2387 ( .A(IR_REG_5__SCAN_IN), .ZN(n2258) );
  NAND2_X1 U2388 ( .A1(n2032), .A2(n2238), .ZN(n2237) );
  INV_X1 U2389 ( .A(n3740), .ZN(n2238) );
  INV_X1 U2390 ( .A(IR_REG_8__SCAN_IN), .ZN(n3498) );
  INV_X1 U2391 ( .A(n3274), .ZN(n2252) );
  NAND2_X1 U2392 ( .A1(n3695), .A2(n3696), .ZN(n3694) );
  INV_X1 U2393 ( .A(n2251), .ZN(n2250) );
  OAI21_X1 U2394 ( .B1(n2511), .B2(n2002), .A(n3273), .ZN(n2251) );
  AND2_X1 U2395 ( .A1(n2002), .A2(n2017), .ZN(n2248) );
  INV_X1 U2396 ( .A(n3696), .ZN(n2241) );
  NAND2_X1 U2397 ( .A1(n2068), .A2(n2242), .ZN(n2067) );
  INV_X1 U2398 ( .A(n3695), .ZN(n2068) );
  NAND2_X1 U2399 ( .A1(n2067), .A2(n2065), .ZN(n3720) );
  AND2_X1 U2400 ( .A1(n2622), .A2(n2003), .ZN(n2079) );
  OR2_X1 U2401 ( .A1(n2733), .A2(n3642), .ZN(n2737) );
  NAND2_X1 U2402 ( .A1(n3639), .A2(n2732), .ZN(n2239) );
  AND2_X1 U2403 ( .A1(n2731), .A2(n3640), .ZN(n2732) );
  INV_X1 U2404 ( .A(n4092), .ZN(n3745) );
  OR2_X1 U2405 ( .A1(n3908), .A2(n3907), .ZN(n3909) );
  OR2_X1 U2406 ( .A1(n2453), .A2(n3189), .ZN(n2442) );
  OR2_X1 U2407 ( .A1(n3831), .A2(n2454), .ZN(n2455) );
  NAND2_X1 U2408 ( .A1(n2052), .A2(n2051), .ZN(n2053) );
  NAND2_X1 U2409 ( .A1(n2879), .A2(REG2_REG_2__SCAN_IN), .ZN(n2051) );
  NAND2_X1 U2410 ( .A1(n4461), .A2(n4292), .ZN(n2052) );
  NAND2_X1 U2411 ( .A1(n2879), .A2(n2836), .ZN(n2837) );
  INV_X1 U2412 ( .A(n3082), .ZN(n2149) );
  AND2_X1 U2413 ( .A1(n2888), .A2(n4474), .ZN(n2151) );
  NAND2_X1 U2414 ( .A1(n2054), .A2(n2056), .ZN(n2055) );
  NAND2_X1 U2415 ( .A1(n3064), .A2(REG2_REG_6__SCAN_IN), .ZN(n2054) );
  OR2_X1 U2416 ( .A1(n3076), .A2(n2849), .ZN(n2850) );
  OR2_X1 U2417 ( .A1(n3101), .A2(n2854), .ZN(n2855) );
  NOR2_X1 U2418 ( .A1(n2553), .A2(n2552), .ZN(n2555) );
  OAI21_X1 U2419 ( .B1(n3966), .B2(n3963), .A(n2899), .ZN(n2900) );
  NAND2_X1 U2420 ( .A1(n4527), .A2(n2907), .ZN(n4540) );
  INV_X1 U2421 ( .A(n2870), .ZN(n2180) );
  INV_X1 U2422 ( .A(n4538), .ZN(n2177) );
  AND2_X1 U2423 ( .A1(n4025), .A2(n2761), .ZN(n3434) );
  NAND2_X1 U2424 ( .A1(n2748), .A2(REG3_REG_27__SCAN_IN), .ZN(n2760) );
  INV_X1 U2425 ( .A(n2750), .ZN(n2748) );
  NOR2_X1 U2426 ( .A1(n2965), .A2(n2232), .ZN(n2231) );
  INV_X1 U2427 ( .A(n2963), .ZN(n2232) );
  AND2_X1 U2428 ( .A1(n3828), .A2(n3825), .ZN(n4040) );
  INV_X1 U2429 ( .A(n3919), .ZN(n4058) );
  NAND2_X1 U2430 ( .A1(n4131), .A2(n4120), .ZN(n2958) );
  NAND2_X1 U2431 ( .A1(n2606), .A2(n2008), .ZN(n2666) );
  INV_X1 U2432 ( .A(n2995), .ZN(n4150) );
  OR2_X1 U2433 ( .A1(n2990), .A2(n4176), .ZN(n2955) );
  AOI21_X1 U2434 ( .B1(n2199), .B2(n2198), .A(n2953), .ZN(n2197) );
  INV_X1 U2435 ( .A(n2952), .ZN(n2198) );
  AND2_X1 U2436 ( .A1(n4256), .A2(n4254), .ZN(n2948) );
  AND2_X1 U2437 ( .A1(n2612), .A2(n2611), .ZN(n4242) );
  NAND2_X1 U2438 ( .A1(n2097), .A2(REG3_REG_15__SCAN_IN), .ZN(n2595) );
  OR2_X1 U2439 ( .A1(n2544), .A2(n3713), .ZN(n2564) );
  INV_X1 U2440 ( .A(n2209), .ZN(n2208) );
  NAND2_X1 U2441 ( .A1(n3249), .A2(n2207), .ZN(n2206) );
  OAI22_X1 U2442 ( .A1(n2210), .A2(n2214), .B1(n3283), .B2(n2218), .ZN(n2209)
         );
  NAND2_X1 U2443 ( .A1(n2497), .A2(n2099), .ZN(n2532) );
  AND2_X1 U2444 ( .A1(n2014), .A2(n2220), .ZN(n2217) );
  AOI21_X1 U2445 ( .B1(n2138), .B2(n2137), .A(n2136), .ZN(n2135) );
  INV_X1 U2446 ( .A(n3785), .ZN(n2137) );
  INV_X1 U2447 ( .A(n3784), .ZN(n2136) );
  OR2_X1 U2448 ( .A1(n2466), .A2(n3092), .ZN(n2485) );
  NAND2_X1 U2449 ( .A1(n2102), .A2(n2415), .ZN(n2452) );
  INV_X1 U2450 ( .A(n2103), .ZN(n2102) );
  NAND2_X1 U2451 ( .A1(n2967), .A2(n3987), .ZN(n4172) );
  NAND2_X1 U2452 ( .A1(n2970), .A2(n3768), .ZN(n2968) );
  AND2_X1 U2453 ( .A1(n2969), .A2(n4571), .ZN(n4551) );
  NAND2_X1 U2454 ( .A1(n2968), .A2(n4551), .ZN(n4550) );
  NOR2_X1 U2455 ( .A1(n4451), .A2(n4452), .ZN(n4570) );
  AND2_X1 U2456 ( .A1(n4059), .A2(n2092), .ZN(n4012) );
  NOR2_X1 U2457 ( .A1(n2093), .A2(n4021), .ZN(n2092) );
  INV_X1 U2458 ( .A(n2094), .ZN(n2093) );
  INV_X1 U2459 ( .A(n3460), .ZN(n4193) );
  AND2_X1 U2460 ( .A1(n4172), .A2(n4388), .ZN(n4629) );
  NOR2_X1 U2461 ( .A1(n3033), .A2(n2300), .ZN(n2301) );
  INV_X1 U2462 ( .A(IR_REG_26__SCAN_IN), .ZN(n2300) );
  INV_X1 U2463 ( .A(n2826), .ZN(n2305) );
  XNOR2_X1 U2464 ( .A(n2281), .B(n2280), .ZN(n2312) );
  INV_X1 U2465 ( .A(IR_REG_20__SCAN_IN), .ZN(n2280) );
  NAND2_X1 U2466 ( .A1(n2279), .A2(IR_REG_31__SCAN_IN), .ZN(n2281) );
  NAND2_X1 U2467 ( .A1(n2578), .A2(IR_REG_31__SCAN_IN), .ZN(n2599) );
  OR2_X1 U2468 ( .A1(n2577), .A2(IR_REG_14__SCAN_IN), .ZN(n2578) );
  XNOR2_X1 U2469 ( .A(n2599), .B(IR_REG_15__SCAN_IN), .ZN(n2903) );
  NAND2_X1 U2470 ( .A1(n2555), .A2(n3491), .ZN(n2577) );
  INV_X1 U2471 ( .A(IR_REG_4__SCAN_IN), .ZN(n2405) );
  INV_X1 U2472 ( .A(IR_REG_3__SCAN_IN), .ZN(n2385) );
  OAI21_X1 U2473 ( .B1(n3707), .B2(n3709), .A(n3708), .ZN(n3443) );
  AND2_X1 U2474 ( .A1(n2744), .A2(n2743), .ZN(n4033) );
  AND2_X1 U2475 ( .A1(n2738), .A2(n2719), .ZN(n4081) );
  AND2_X1 U2476 ( .A1(n2253), .A2(n2071), .ZN(n2070) );
  AND2_X1 U2477 ( .A1(n2673), .A2(n2672), .ZN(n4168) );
  OR2_X1 U2478 ( .A1(n4146), .A2(n2453), .ZN(n2673) );
  INV_X1 U2479 ( .A(n4168), .ZN(n4129) );
  INV_X1 U2480 ( .A(n4242), .ZN(n4205) );
  INV_X1 U2481 ( .A(n3316), .ZN(n3928) );
  AND2_X1 U2482 ( .A1(n2914), .A2(n2912), .ZN(n4465) );
  OAI21_X1 U2483 ( .B1(n2880), .B2(REG2_REG_1__SCAN_IN), .A(n2158), .ZN(n3938)
         );
  NAND2_X1 U2484 ( .A1(n2880), .A2(REG2_REG_1__SCAN_IN), .ZN(n2158) );
  NAND2_X1 U2485 ( .A1(n3938), .A2(n3946), .ZN(n3951) );
  XNOR2_X1 U2486 ( .A(n2474), .B(n2473), .ZN(n3076) );
  NAND2_X1 U2487 ( .A1(n4487), .A2(n2142), .ZN(n3203) );
  XNOR2_X1 U2488 ( .A(n2898), .B(n4602), .ZN(n4497) );
  NAND2_X1 U2489 ( .A1(n4497), .A2(REG2_REG_12__SCAN_IN), .ZN(n4496) );
  XNOR2_X1 U2490 ( .A(n2900), .B(n2901), .ZN(n4506) );
  NAND2_X1 U2491 ( .A1(n4526), .A2(n4525), .ZN(n4524) );
  AND4_X1 U2492 ( .A1(n2118), .A2(n2117), .A3(n2116), .A4(n2010), .ZN(n4306)
         );
  NAND2_X1 U2493 ( .A1(n2123), .A2(n2120), .ZN(n2116) );
  AND2_X1 U2494 ( .A1(n2312), .A2(n3982), .ZN(n4572) );
  INV_X1 U2495 ( .A(n3698), .ZN(n2244) );
  AND2_X1 U2496 ( .A1(n2081), .A2(n2080), .ZN(n3650) );
  INV_X1 U2497 ( .A(n2772), .ZN(n2716) );
  OAI21_X1 U2498 ( .B1(n3902), .B2(n3901), .A(n3900), .ZN(n3904) );
  AND2_X1 U2499 ( .A1(n3842), .A2(n4050), .ZN(n3895) );
  NOR2_X1 U2500 ( .A1(n3082), .A2(n2398), .ZN(n2150) );
  INV_X1 U2501 ( .A(n2231), .ZN(n2225) );
  NOR2_X1 U2502 ( .A1(n2689), .A2(n2665), .ZN(n2098) );
  NAND2_X1 U2503 ( .A1(n2109), .A2(n2107), .ZN(n2113) );
  NOR2_X1 U2504 ( .A1(n3887), .A2(n2108), .ZN(n2107) );
  AND2_X1 U2505 ( .A1(n2105), .A2(REG3_REG_19__SCAN_IN), .ZN(n2104) );
  INV_X1 U2506 ( .A(n2666), .ZN(n2664) );
  OAI21_X1 U2507 ( .B1(n4229), .B2(n2196), .A(n2193), .ZN(n2192) );
  NAND2_X1 U2508 ( .A1(n2199), .A2(n2954), .ZN(n2196) );
  INV_X1 U2509 ( .A(n2194), .ZN(n2193) );
  AND2_X1 U2510 ( .A1(n4202), .A2(n4159), .ZN(n4184) );
  NOR2_X1 U2511 ( .A1(n2623), .A2(n2106), .ZN(n2105) );
  INV_X1 U2512 ( .A(n2016), .ZN(n2606) );
  AND2_X1 U2513 ( .A1(n4205), .A2(n4223), .ZN(n4105) );
  NOR2_X1 U2514 ( .A1(n2564), .A2(n2563), .ZN(n2097) );
  NAND2_X1 U2515 ( .A1(n2219), .A2(n2211), .ZN(n2210) );
  INV_X1 U2516 ( .A(n2218), .ZN(n2211) );
  NOR2_X1 U2517 ( .A1(n2210), .A2(n2213), .ZN(n2207) );
  NOR2_X1 U2518 ( .A1(n3205), .A2(n2100), .ZN(n2099) );
  INV_X1 U2519 ( .A(n2498), .ZN(n2497) );
  AND2_X1 U2520 ( .A1(n3191), .A2(n2928), .ZN(n2929) );
  NAND2_X1 U2521 ( .A1(n2931), .A2(n3215), .ZN(n2933) );
  AND2_X1 U2522 ( .A1(n3110), .A2(n2932), .ZN(n3191) );
  INV_X1 U2523 ( .A(n3933), .ZN(n3333) );
  NOR2_X1 U2524 ( .A1(n3420), .A2(n4010), .ZN(n2094) );
  NOR2_X1 U2525 ( .A1(n2089), .A2(n3687), .ZN(n2088) );
  INV_X1 U2526 ( .A(n2090), .ZN(n2089) );
  NOR2_X1 U2527 ( .A1(n4128), .A2(n3845), .ZN(n2090) );
  AND2_X1 U2528 ( .A1(n2259), .A2(n2266), .ZN(n2257) );
  NOR2_X1 U2529 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2259)
         );
  XNOR2_X1 U2530 ( .A(n2388), .B(n2674), .ZN(n2392) );
  OAI22_X1 U2531 ( .A1(n2926), .A2(n2397), .B1(n3310), .B2(n2367), .ZN(n2388)
         );
  NAND2_X1 U2532 ( .A1(n2875), .A2(IR_REG_27__SCAN_IN), .ZN(n2330) );
  NOR2_X1 U2533 ( .A1(n2076), .A2(n2074), .ZN(n2073) );
  INV_X1 U2534 ( .A(n2260), .ZN(n2076) );
  INV_X1 U2535 ( .A(n3659), .ZN(n2074) );
  AND2_X1 U2536 ( .A1(n2254), .A2(n2465), .ZN(n2253) );
  INV_X1 U2537 ( .A(n3172), .ZN(n2254) );
  NAND2_X1 U2538 ( .A1(n2075), .A2(n2260), .ZN(n2071) );
  INV_X1 U2539 ( .A(n2434), .ZN(n2075) );
  NAND2_X1 U2540 ( .A1(n2351), .A2(n2265), .ZN(n3131) );
  OAI21_X1 U2541 ( .B1(n2772), .B2(n2354), .A(n2353), .ZN(n3130) );
  INV_X1 U2542 ( .A(n2352), .ZN(n2353) );
  NAND2_X1 U2543 ( .A1(n2606), .A2(n2104), .ZN(n2651) );
  NAND2_X1 U2544 ( .A1(n3242), .A2(n2511), .ZN(n3239) );
  OR2_X1 U2545 ( .A1(n2828), .A2(n3002), .ZN(n3744) );
  OR2_X1 U2546 ( .A1(n3132), .A2(n3010), .ZN(n2818) );
  OR2_X1 U2547 ( .A1(n2813), .A2(n2812), .ZN(n2825) );
  NAND2_X1 U2548 ( .A1(n3078), .A2(n2892), .ZN(n2893) );
  OR2_X1 U2549 ( .A1(n3076), .A2(n3570), .ZN(n2892) );
  NOR2_X1 U2550 ( .A1(n4482), .A2(n2857), .ZN(n3210) );
  NAND2_X1 U2551 ( .A1(n2183), .A2(REG1_REG_12__SCAN_IN), .ZN(n2181) );
  NAND2_X1 U2552 ( .A1(n2182), .A2(n2181), .ZN(n3968) );
  NAND2_X1 U2553 ( .A1(n3968), .A2(n2861), .ZN(n3969) );
  INV_X1 U2554 ( .A(n3971), .ZN(n2861) );
  NAND2_X1 U2555 ( .A1(n2186), .A2(REG1_REG_14__SCAN_IN), .ZN(n2185) );
  NAND2_X1 U2556 ( .A1(n2864), .A2(n2186), .ZN(n2184) );
  INV_X1 U2557 ( .A(n4515), .ZN(n2186) );
  NOR2_X1 U2558 ( .A1(n4502), .A2(n4503), .ZN(n4501) );
  AOI21_X1 U2559 ( .B1(n2011), .B2(n2155), .A(n3981), .ZN(n2154) );
  INV_X1 U2560 ( .A(n4541), .ZN(n2155) );
  INV_X1 U2561 ( .A(n3839), .ZN(n4021) );
  NAND2_X1 U2562 ( .A1(n4032), .A2(n4014), .ZN(n2122) );
  NOR2_X1 U2563 ( .A1(n4307), .A2(n2121), .ZN(n2120) );
  AND2_X1 U2564 ( .A1(n2767), .A2(n2766), .ZN(n4036) );
  NAND2_X1 U2565 ( .A1(n2664), .A2(n2098), .ZN(n2704) );
  AND2_X1 U2566 ( .A1(n2710), .A2(n2709), .ZN(n4115) );
  AND2_X1 U2567 ( .A1(n2630), .A2(n2629), .ZN(n4186) );
  INV_X1 U2568 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2623) );
  NAND2_X1 U2569 ( .A1(n2606), .A2(n2105), .ZN(n2640) );
  AND2_X1 U2570 ( .A1(n2647), .A2(n2646), .ZN(n4207) );
  NAND2_X1 U2571 ( .A1(n2606), .A2(REG3_REG_17__SCAN_IN), .ZN(n2624) );
  NAND2_X1 U2572 ( .A1(n2115), .A2(n2114), .ZN(n4267) );
  INV_X1 U2573 ( .A(n4270), .ZN(n2115) );
  INV_X1 U2574 ( .A(n2097), .ZN(n2593) );
  AND4_X1 U2575 ( .A1(n2549), .A2(n2548), .A3(n2547), .A4(n2546), .ZN(n3380)
         );
  INV_X1 U2576 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3205) );
  OAI21_X1 U2577 ( .B1(n3249), .B2(n2205), .A(n2204), .ZN(n3284) );
  AOI21_X1 U2578 ( .B1(n2214), .B2(n2213), .A(n2212), .ZN(n2204) );
  INV_X1 U2579 ( .A(n2214), .ZN(n2205) );
  NAND2_X1 U2580 ( .A1(n2497), .A2(REG3_REG_10__SCAN_IN), .ZN(n2516) );
  AND4_X1 U2581 ( .A1(n2490), .A2(n2489), .A3(n2488), .A4(n2487), .ZN(n3316)
         );
  AND4_X1 U2582 ( .A1(n2522), .A2(n2521), .A3(n2520), .A4(n2519), .ZN(n3364)
         );
  NAND2_X1 U2583 ( .A1(n2483), .A2(REG3_REG_9__SCAN_IN), .ZN(n2498) );
  INV_X1 U2584 ( .A(n2485), .ZN(n2483) );
  INV_X1 U2585 ( .A(REG3_REG_8__SCAN_IN), .ZN(n3092) );
  NOR2_X1 U2586 ( .A1(n2103), .A2(n2435), .ZN(n2101) );
  NAND2_X1 U2587 ( .A1(n4636), .A2(n3185), .ZN(n3255) );
  NAND2_X1 U2588 ( .A1(n2131), .A2(n2132), .ZN(n2130) );
  AND2_X1 U2589 ( .A1(n2132), .A2(n3860), .ZN(n2128) );
  NAND2_X1 U2590 ( .A1(n2415), .A2(REG3_REG_5__SCAN_IN), .ZN(n2450) );
  NAND2_X1 U2591 ( .A1(n2129), .A2(n3779), .ZN(n3219) );
  NAND2_X1 U2592 ( .A1(n3301), .A2(n2134), .ZN(n2129) );
  INV_X1 U2593 ( .A(n2131), .ZN(n2134) );
  OR2_X1 U2594 ( .A1(n3116), .A2(n3412), .ZN(n3226) );
  NAND2_X1 U2595 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2417) );
  NAND2_X1 U2596 ( .A1(n3301), .A2(n3775), .ZN(n3111) );
  AND2_X1 U2597 ( .A1(n3003), .A2(n4448), .ZN(n4559) );
  INV_X1 U2598 ( .A(n4576), .ZN(n4557) );
  NAND2_X1 U2599 ( .A1(n3003), .A2(n3002), .ZN(n4576) );
  INV_X1 U2600 ( .A(n4273), .ZN(n4563) );
  AND2_X1 U2601 ( .A1(n4453), .A2(n4570), .ZN(n4273) );
  NAND2_X1 U2602 ( .A1(n4059), .A2(n2094), .ZN(n4013) );
  NAND2_X1 U2603 ( .A1(n4059), .A2(n4041), .ZN(n3017) );
  NOR2_X1 U2604 ( .A1(n4078), .A2(n4055), .ZN(n4059) );
  NAND2_X1 U2605 ( .A1(n4138), .A2(n2086), .ZN(n4078) );
  NOR2_X1 U2606 ( .A1(n2087), .A2(n3016), .ZN(n2086) );
  INV_X1 U2607 ( .A(n2088), .ZN(n2087) );
  NAND2_X1 U2608 ( .A1(n4138), .A2(n2088), .ZN(n4097) );
  INV_X1 U2609 ( .A(n4165), .ZN(n4176) );
  NAND2_X1 U2610 ( .A1(n4174), .A2(n4176), .ZN(n4175) );
  NAND2_X1 U2611 ( .A1(n4274), .A2(n2006), .ZN(n4233) );
  NAND2_X1 U2612 ( .A1(n3321), .A2(n3292), .ZN(n3369) );
  AND2_X1 U2613 ( .A1(n4636), .A2(n2005), .ZN(n3324) );
  NAND2_X1 U2614 ( .A1(n4636), .A2(n2096), .ZN(n4385) );
  INV_X1 U2615 ( .A(n3020), .ZN(n4635) );
  NOR2_X1 U2616 ( .A1(n3013), .A2(n3119), .ZN(n3023) );
  AND2_X1 U2617 ( .A1(n2777), .A2(n4449), .ZN(n3043) );
  AND2_X1 U2618 ( .A1(n2256), .A2(n2026), .ZN(n2082) );
  INV_X1 U2619 ( .A(IR_REG_28__SCAN_IN), .ZN(n2315) );
  INV_X1 U2620 ( .A(IR_REG_29__SCAN_IN), .ZN(n2318) );
  NAND2_X1 U2621 ( .A1(n2310), .A2(n2012), .ZN(n2778) );
  OR2_X1 U2622 ( .A1(n2553), .A2(IR_REG_10__SCAN_IN), .ZN(n2523) );
  INV_X1 U2623 ( .A(IR_REG_11__SCAN_IN), .ZN(n3532) );
  INV_X1 U2624 ( .A(IR_REG_10__SCAN_IN), .ZN(n2551) );
  XNOR2_X1 U2625 ( .A(n2476), .B(n3498), .ZN(n4456) );
  NAND2_X1 U2626 ( .A1(n2369), .A2(n3033), .ZN(n2173) );
  INV_X1 U2627 ( .A(IR_REG_1__SCAN_IN), .ZN(n2156) );
  NAND2_X1 U2628 ( .A1(n2233), .A2(n2237), .ZN(n3419) );
  NAND2_X1 U2629 ( .A1(n2236), .A2(n2234), .ZN(n2798) );
  NAND2_X1 U2630 ( .A1(n3418), .A2(n2235), .ZN(n2234) );
  NAND2_X1 U2631 ( .A1(n2239), .A2(n2031), .ZN(n2236) );
  INV_X1 U2632 ( .A(n2237), .ZN(n2235) );
  NAND2_X1 U2633 ( .A1(n3149), .A2(n2260), .ZN(n2255) );
  NAND2_X1 U2634 ( .A1(n3694), .A2(n3698), .ZN(n3613) );
  OR2_X1 U2635 ( .A1(n3242), .A2(n2002), .ZN(n2245) );
  AOI21_X1 U2636 ( .B1(n3685), .B2(n3682), .A(n3684), .ZN(n3644) );
  NAND2_X1 U2637 ( .A1(n3660), .A2(n3659), .ZN(n3658) );
  INV_X1 U2638 ( .A(n4571), .ZN(n3767) );
  INV_X1 U2639 ( .A(n3724), .ZN(n3702) );
  OR2_X1 U2640 ( .A1(n2828), .A2(n4448), .ZN(n3701) );
  AOI21_X1 U2641 ( .B1(n2250), .B2(n2248), .A(n2247), .ZN(n2246) );
  NOR2_X1 U2642 ( .A1(n3625), .A2(n3624), .ZN(n2247) );
  AND2_X1 U2643 ( .A1(n2067), .A2(n2240), .ZN(n3721) );
  NAND2_X1 U2644 ( .A1(n3239), .A2(n2515), .ZN(n3277) );
  NAND2_X1 U2645 ( .A1(n2621), .A2(n2003), .ZN(n2078) );
  INV_X1 U2646 ( .A(n3744), .ZN(n3757) );
  AND2_X1 U2647 ( .A1(n2750), .A2(n2739), .ZN(n4063) );
  INV_X1 U2648 ( .A(n3762), .ZN(n3747) );
  INV_X1 U2649 ( .A(n3701), .ZN(n3759) );
  INV_X1 U2650 ( .A(n3702), .ZN(n3758) );
  INV_X1 U2651 ( .A(n3750), .ZN(n3764) );
  MUX2_X1 U2652 ( .A(n3912), .B(n3911), .S(n4453), .Z(n3913) );
  AOI21_X1 U2653 ( .B1(n2824), .B2(n2320), .A(n2823), .ZN(n3840) );
  INV_X1 U2654 ( .A(n4036), .ZN(n4022) );
  NAND2_X1 U2655 ( .A1(n2758), .A2(n2757), .ZN(n3919) );
  OR2_X1 U2656 ( .A1(n4044), .A2(n2453), .ZN(n2758) );
  INV_X1 U2657 ( .A(n4033), .ZN(n4075) );
  NAND2_X1 U2658 ( .A1(n2725), .A2(n2724), .ZN(n4092) );
  NAND2_X1 U2659 ( .A1(n2684), .A2(n2683), .ZN(n4149) );
  NAND2_X1 U2660 ( .A1(n2657), .A2(n2656), .ZN(n4188) );
  INV_X1 U2661 ( .A(n4207), .ZN(n4166) );
  INV_X1 U2662 ( .A(n4186), .ZN(n4225) );
  NAND2_X1 U2663 ( .A1(n2588), .A2(n2587), .ZN(n3922) );
  OAI211_X1 U2664 ( .C1(n2764), .C2(n2598), .A(n2597), .B(n2596), .ZN(n3923)
         );
  INV_X1 U2665 ( .A(n3380), .ZN(n3925) );
  NAND4_X1 U2666 ( .A1(n2443), .A2(n2442), .A3(n2441), .A4(n2440), .ZN(n3931)
         );
  NAND4_X1 U2667 ( .A1(n2458), .A2(n2457), .A3(n2456), .A4(n2455), .ZN(n3932)
         );
  INV_X1 U2668 ( .A(n2053), .ZN(n3952) );
  NAND2_X1 U2669 ( .A1(n2165), .A2(n2164), .ZN(n3084) );
  AND2_X1 U2670 ( .A1(n2167), .A2(n2171), .ZN(n3086) );
  INV_X1 U2671 ( .A(n2845), .ZN(n2171) );
  NAND2_X1 U2672 ( .A1(n4472), .A2(REG1_REG_4__SCAN_IN), .ZN(n2167) );
  OAI21_X1 U2673 ( .B1(n2151), .B2(REG2_REG_4__SCAN_IN), .A(n2149), .ZN(n2147)
         );
  NOR2_X1 U2674 ( .A1(n4469), .A2(n2151), .ZN(n2148) );
  AND2_X1 U2675 ( .A1(n2146), .A2(n2145), .ZN(n3083) );
  INV_X1 U2676 ( .A(n2151), .ZN(n2145) );
  NAND2_X1 U2677 ( .A1(n4469), .A2(REG2_REG_4__SCAN_IN), .ZN(n2146) );
  NAND2_X1 U2678 ( .A1(n2055), .A2(n2891), .ZN(n3078) );
  INV_X1 U2679 ( .A(n3073), .ZN(n2891) );
  INV_X1 U2680 ( .A(n2055), .ZN(n3074) );
  INV_X1 U2681 ( .A(n2170), .ZN(n2847) );
  XNOR2_X1 U2682 ( .A(n2896), .B(n2895), .ZN(n4488) );
  NAND2_X1 U2683 ( .A1(n4488), .A2(REG2_REG_10__SCAN_IN), .ZN(n4487) );
  NAND2_X1 U2684 ( .A1(n2182), .A2(n2183), .ZN(n4492) );
  NOR2_X1 U2685 ( .A1(n2859), .A2(n2181), .ZN(n4491) );
  OR2_X1 U2686 ( .A1(n2557), .A2(n2556), .ZN(n3977) );
  NAND2_X1 U2687 ( .A1(n2058), .A2(n4602), .ZN(n2057) );
  INV_X1 U2688 ( .A(n2898), .ZN(n2058) );
  NOR2_X1 U2689 ( .A1(n4506), .A2(n3385), .ZN(n4505) );
  NAND2_X1 U2690 ( .A1(n2163), .A2(REG2_REG_14__SCAN_IN), .ZN(n2162) );
  INV_X1 U2691 ( .A(n4519), .ZN(n2163) );
  AND2_X1 U2692 ( .A1(n4465), .A2(n3993), .ZN(n4545) );
  NAND2_X1 U2693 ( .A1(n2910), .A2(n2911), .ZN(n2061) );
  NAND2_X1 U2694 ( .A1(n4539), .A2(n2909), .ZN(n2910) );
  NAND2_X1 U2695 ( .A1(n4536), .A2(n2870), .ZN(n2877) );
  INV_X1 U2696 ( .A(n4545), .ZN(n4513) );
  AND2_X1 U2697 ( .A1(n4465), .A2(n3947), .ZN(n4543) );
  AOI21_X1 U2698 ( .B1(n2178), .B2(n2177), .A(n2050), .ZN(n2176) );
  NAND2_X1 U2699 ( .A1(n2228), .A2(n2229), .ZN(n4039) );
  NAND2_X1 U2700 ( .A1(n4068), .A2(n2231), .ZN(n2228) );
  AND2_X1 U2701 ( .A1(n2190), .A2(n2029), .ZN(n4136) );
  NAND2_X1 U2702 ( .A1(n2190), .A2(n2001), .ZN(n4135) );
  NAND2_X1 U2703 ( .A1(n2191), .A2(n2268), .ZN(n2190) );
  OAI21_X1 U2704 ( .B1(n4229), .B2(n2200), .A(n2197), .ZN(n4192) );
  NAND2_X1 U2705 ( .A1(n2201), .A2(n2199), .ZN(n4210) );
  AND2_X1 U2706 ( .A1(n2201), .A2(n2018), .ZN(n4212) );
  NAND2_X1 U2707 ( .A1(n4229), .A2(n2952), .ZN(n2201) );
  NAND2_X1 U2708 ( .A1(n3249), .A2(n2217), .ZN(n2215) );
  NAND2_X1 U2709 ( .A1(n2216), .A2(n2220), .ZN(n3270) );
  OR2_X1 U2710 ( .A1(n3249), .A2(n2939), .ZN(n2216) );
  INV_X1 U2711 ( .A(n4283), .ZN(n4258) );
  AND2_X1 U2712 ( .A1(n4581), .A2(n3987), .ZN(n4215) );
  XNOR2_X1 U2713 ( .A(n2338), .B(IR_REG_19__SCAN_IN), .ZN(n3982) );
  OAI21_X1 U2714 ( .B1(n2968), .B2(n4551), .A(n4550), .ZN(n4552) );
  AND2_X1 U2715 ( .A1(n4641), .A2(n2817), .ZN(n4578) );
  AND2_X1 U2716 ( .A1(n4581), .A2(n3127), .ZN(n4579) );
  INV_X1 U2717 ( .A(n4658), .ZN(n4656) );
  NOR2_X1 U2718 ( .A1(n4306), .A2(n4305), .ZN(n4311) );
  AND2_X1 U2719 ( .A1(n4274), .A2(n2030), .ZN(n4194) );
  AND2_X2 U2720 ( .A1(n3023), .A2(n3122), .ZN(n4647) );
  NOR2_X1 U2721 ( .A1(n2305), .A2(n2304), .ZN(n2306) );
  NAND2_X1 U2722 ( .A1(n2012), .A2(n2301), .ZN(n2307) );
  NOR2_X1 U2723 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2304)
         );
  INV_X1 U2724 ( .A(n3046), .ZN(n4449) );
  AND2_X1 U2725 ( .A1(n2873), .A2(STATE_REG_SCAN_IN), .ZN(n4591) );
  XNOR2_X1 U2726 ( .A(n2314), .B(IR_REG_22__SCAN_IN), .ZN(n4451) );
  INV_X1 U2727 ( .A(n3982), .ZN(n3987) );
  XNOR2_X1 U2728 ( .A(n2582), .B(n2581), .ZN(n4597) );
  AND2_X1 U2729 ( .A1(n2404), .A2(n2387), .ZN(n4460) );
  NAND2_X1 U2730 ( .A1(n2062), .A2(n2059), .ZN(U3258) );
  NAND2_X1 U2731 ( .A1(n2878), .A2(n3978), .ZN(n2062) );
  AND2_X1 U2732 ( .A1(n2060), .A2(n2919), .ZN(n2059) );
  NAND2_X1 U2733 ( .A1(n4536), .A2(n2178), .ZN(n3978) );
  AND2_X1 U2734 ( .A1(n2957), .A2(n2029), .ZN(n2001) );
  NAND2_X1 U2735 ( .A1(n3262), .A2(n2976), .ZN(n2220) );
  NAND2_X1 U2736 ( .A1(n4138), .A2(n4139), .ZN(n4119) );
  NAND2_X1 U2737 ( .A1(n2252), .A2(n2515), .ZN(n2002) );
  MUX2_X1 U2738 ( .A(n2370), .B(n2879), .S(n2872), .Z(n4287) );
  NAND2_X1 U2739 ( .A1(n3776), .A2(n3779), .ZN(n3110) );
  AND2_X1 U2740 ( .A1(n2272), .A2(n2256), .ZN(n2426) );
  NAND2_X1 U2741 ( .A1(n3674), .A2(n3673), .ZN(n2003) );
  NAND2_X1 U2742 ( .A1(n3770), .A2(n3772), .ZN(n2971) );
  NAND2_X1 U2743 ( .A1(n2272), .A2(n2266), .ZN(n2424) );
  AND2_X1 U2744 ( .A1(n2125), .A2(n4307), .ZN(n2004) );
  NAND2_X1 U2745 ( .A1(n4138), .A2(n2090), .ZN(n2091) );
  NAND2_X1 U2746 ( .A1(n2323), .A2(n3037), .ZN(n2399) );
  INV_X2 U2747 ( .A(n2399), .ZN(n2320) );
  AND2_X1 U2748 ( .A1(n2096), .A2(n2977), .ZN(n2005) );
  AND2_X1 U2749 ( .A1(n4023), .A2(n4024), .ZN(n2126) );
  AND2_X1 U2750 ( .A1(n4248), .A2(n4223), .ZN(n2006) );
  AND2_X1 U2751 ( .A1(n2215), .A2(n2046), .ZN(n2007) );
  NAND2_X1 U2752 ( .A1(n2696), .A2(n2695), .ZN(n3921) );
  OR2_X1 U2753 ( .A1(n2269), .A2(n2244), .ZN(n2243) );
  AND2_X1 U2754 ( .A1(n2104), .A2(REG3_REG_20__SCAN_IN), .ZN(n2008) );
  AND2_X1 U2755 ( .A1(n2032), .A2(n2264), .ZN(n2009) );
  NAND2_X1 U2756 ( .A1(n2126), .A2(n4288), .ZN(n2010) );
  NOR2_X1 U2757 ( .A1(n2911), .A2(n2908), .ZN(n2011) );
  NAND2_X1 U2758 ( .A1(n3782), .A2(n3785), .ZN(n3180) );
  OR2_X1 U2759 ( .A1(n2308), .A2(IR_REG_25__SCAN_IN), .ZN(n2012) );
  AND3_X1 U2760 ( .A1(n2365), .A2(n2364), .A3(n2363), .ZN(n2013) );
  OAI21_X1 U2761 ( .B1(n2631), .B2(IR_REG_18__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2338) );
  NAND2_X1 U2762 ( .A1(n3316), .A2(n2977), .ZN(n2014) );
  OR3_X1 U2763 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .A3(
        IR_REG_25__SCAN_IN), .ZN(n2015) );
  NAND2_X1 U2764 ( .A1(n4211), .A2(n2018), .ZN(n2200) );
  NOR2_X1 U2765 ( .A1(n4175), .A2(n4150), .ZN(n4138) );
  OR2_X1 U2766 ( .A1(n2595), .A2(n3653), .ZN(n2016) );
  NAND4_X1 U2767 ( .A1(n2345), .A2(n2344), .A3(n2343), .A4(n2342), .ZN(n2969)
         );
  AOI21_X1 U2768 ( .B1(n3729), .B2(n3730), .A(n3731), .ZN(n3458) );
  NAND2_X2 U2769 ( .A1(n3126), .A2(n2349), .ZN(n2367) );
  NAND2_X1 U2770 ( .A1(n3625), .A2(n3624), .ZN(n2017) );
  NAND2_X1 U2771 ( .A1(n4205), .A2(n4231), .ZN(n2018) );
  NAND2_X1 U2772 ( .A1(n2013), .A2(n2366), .ZN(n4558) );
  INV_X1 U2773 ( .A(n2192), .ZN(n4158) );
  NOR2_X1 U2774 ( .A1(n4505), .A2(n2902), .ZN(n2019) );
  NOR2_X1 U2775 ( .A1(n4501), .A2(n2864), .ZN(n2020) );
  OR2_X1 U2776 ( .A1(n2846), .A2(n4653), .ZN(n2021) );
  AND2_X1 U2777 ( .A1(n4267), .A2(n3798), .ZN(n2022) );
  OR2_X1 U2778 ( .A1(n3117), .A2(n3934), .ZN(n3776) );
  INV_X1 U2779 ( .A(IR_REG_2__SCAN_IN), .ZN(n2369) );
  INV_X1 U2780 ( .A(n3285), .ZN(n3927) );
  AND4_X1 U2781 ( .A1(n2503), .A2(n2502), .A3(n2501), .A4(n2500), .ZN(n3285)
         );
  INV_X1 U2782 ( .A(n3262), .ZN(n3930) );
  AND4_X1 U2783 ( .A1(n2472), .A2(n2471), .A3(n2470), .A4(n2469), .ZN(n3262)
         );
  NOR2_X1 U2784 ( .A1(n4225), .A2(n4204), .ZN(n2953) );
  INV_X1 U2785 ( .A(n2200), .ZN(n2199) );
  INV_X1 U2786 ( .A(n2219), .ZN(n2212) );
  NAND2_X1 U2787 ( .A1(n3285), .A2(n3323), .ZN(n2219) );
  OR2_X1 U2788 ( .A1(n3285), .A2(n3323), .ZN(n2023) );
  AND2_X1 U2789 ( .A1(n3030), .A2(REG2_REG_5__SCAN_IN), .ZN(n2024) );
  AND2_X1 U2790 ( .A1(n2099), .A2(REG3_REG_12__SCAN_IN), .ZN(n2025) );
  AND2_X1 U2791 ( .A1(n2874), .A2(n2315), .ZN(n2026) );
  NOR2_X1 U2792 ( .A1(n3217), .A2(n2133), .ZN(n2132) );
  AND2_X1 U2793 ( .A1(n2250), .A2(n2017), .ZN(n2027) );
  NAND2_X1 U2794 ( .A1(n2368), .A2(n2369), .ZN(n2384) );
  NAND2_X1 U2795 ( .A1(n4539), .A2(n2011), .ZN(n2028) );
  INV_X1 U2796 ( .A(n2139), .ZN(n2138) );
  NAND2_X1 U2797 ( .A1(n3786), .A2(n2140), .ZN(n2139) );
  NAND2_X1 U2798 ( .A1(n3658), .A2(n2434), .ZN(n3149) );
  INV_X1 U2799 ( .A(n4269), .ZN(n2114) );
  INV_X1 U2800 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2100) );
  INV_X1 U2801 ( .A(n2243), .ZN(n2242) );
  INV_X1 U2802 ( .A(n4128), .ZN(n4139) );
  OR2_X1 U2803 ( .A1(n4129), .A2(n4150), .ZN(n2029) );
  NAND2_X1 U2804 ( .A1(n2245), .A2(n2250), .ZN(n3623) );
  NAND2_X1 U2805 ( .A1(n4022), .A2(n3018), .ZN(n4014) );
  NAND2_X1 U2806 ( .A1(n2249), .A2(n2246), .ZN(n3707) );
  NAND2_X1 U2807 ( .A1(n2255), .A2(n2465), .ZN(n3170) );
  AND2_X1 U2808 ( .A1(n2006), .A2(n4213), .ZN(n2030) );
  AND2_X1 U2809 ( .A1(n3418), .A2(n2009), .ZN(n2031) );
  OR2_X1 U2810 ( .A1(n2747), .A2(n2746), .ZN(n2032) );
  AND2_X1 U2811 ( .A1(n4149), .A2(n4128), .ZN(n2033) );
  NOR2_X1 U2812 ( .A1(n2858), .A2(n4500), .ZN(n2859) );
  INV_X1 U2813 ( .A(n2859), .ZN(n2182) );
  AND2_X1 U2814 ( .A1(n3394), .A2(n3015), .ZN(n2034) );
  XNOR2_X1 U2815 ( .A(n2540), .B(IR_REG_12__SCAN_IN), .ZN(n4602) );
  OR2_X1 U2816 ( .A1(n4188), .A2(n4165), .ZN(n2035) );
  AND2_X1 U2817 ( .A1(n3919), .A2(n3420), .ZN(n2036) );
  AND2_X1 U2818 ( .A1(n2962), .A2(n2961), .ZN(n2037) );
  OAI21_X1 U2819 ( .B1(n2524), .B2(n3532), .A(n2539), .ZN(n3207) );
  AND2_X1 U2820 ( .A1(n2226), .A2(n2961), .ZN(n2038) );
  AND2_X1 U2821 ( .A1(n3712), .A2(n3925), .ZN(n2039) );
  AND2_X1 U2822 ( .A1(n4033), .A2(n4061), .ZN(n2040) );
  NAND2_X1 U2823 ( .A1(n4207), .A2(n4193), .ZN(n2041) );
  AND2_X1 U2824 ( .A1(n2678), .A2(n3614), .ZN(n2042) );
  NAND2_X1 U2825 ( .A1(n3452), .A2(n3451), .ZN(n2043) );
  AND2_X1 U2826 ( .A1(n4455), .A2(REG2_REG_9__SCAN_IN), .ZN(n2044) );
  OAI21_X1 U2827 ( .B1(n4016), .B2(n3828), .A(n4015), .ZN(n2123) );
  NAND2_X1 U2828 ( .A1(n4274), .A2(n4248), .ZN(n4230) );
  INV_X1 U2829 ( .A(n3798), .ZN(n2112) );
  NOR2_X1 U2830 ( .A1(n2069), .A2(n2066), .ZN(n2065) );
  AOI21_X1 U2831 ( .B1(n2242), .B2(n2241), .A(n2042), .ZN(n2240) );
  AND2_X1 U2832 ( .A1(n2030), .A2(n4193), .ZN(n2045) );
  INV_X1 U2833 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2639) );
  INV_X1 U2834 ( .A(n2126), .ZN(n2121) );
  INV_X1 U2835 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2106) );
  NOR2_X1 U2836 ( .A1(n3116), .A2(n2085), .ZN(n3225) );
  NOR2_X1 U2837 ( .A1(n4565), .A2(n4293), .ZN(n3309) );
  INV_X1 U2838 ( .A(n3420), .ZN(n4041) );
  AND2_X1 U2839 ( .A1(n2203), .A2(n2940), .ZN(n2046) );
  NOR2_X1 U2840 ( .A1(n2148), .A2(n2147), .ZN(n2047) );
  INV_X1 U2841 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3700) );
  NAND2_X1 U2842 ( .A1(n3001), .A2(n3000), .ZN(n4573) );
  AND2_X1 U2843 ( .A1(n2098), .A2(REG3_REG_24__SCAN_IN), .ZN(n2048) );
  INV_X1 U2844 ( .A(n3117), .ZN(n3412) );
  INV_X1 U2845 ( .A(n2179), .ZN(n2178) );
  OR2_X1 U2846 ( .A1(n2876), .A2(n2180), .ZN(n2179) );
  XNOR2_X1 U2847 ( .A(n2459), .B(IR_REG_6__SCAN_IN), .ZN(n4459) );
  INV_X1 U2848 ( .A(n4459), .ZN(n2169) );
  XOR2_X1 U2849 ( .A(n3982), .B(REG1_REG_19__SCAN_IN), .Z(n2049) );
  AND2_X1 U2850 ( .A1(n4592), .A2(REG1_REG_18__SCAN_IN), .ZN(n2050) );
  NAND2_X1 U2851 ( .A1(n3936), .A2(n3937), .ZN(n3935) );
  NAND2_X1 U2852 ( .A1(n2882), .A2(n2053), .ZN(n3954) );
  AOI21_X2 U2853 ( .B1(n3100), .B2(n3099), .A(n2044), .ZN(n2896) );
  NAND2_X1 U2854 ( .A1(n2890), .A2(n4459), .ZN(n2056) );
  NAND3_X1 U2855 ( .A1(n2028), .A2(n4543), .A3(n2061), .ZN(n2060) );
  NAND2_X1 U2856 ( .A1(n3695), .A2(n2065), .ZN(n2063) );
  INV_X1 U2857 ( .A(n2240), .ZN(n2069) );
  NAND2_X1 U2858 ( .A1(n2073), .A2(n3660), .ZN(n2072) );
  NAND2_X1 U2859 ( .A1(n2072), .A2(n2070), .ZN(n2482) );
  NAND3_X1 U2860 ( .A1(n2081), .A2(n2080), .A3(n2079), .ZN(n2077) );
  NAND2_X1 U2861 ( .A1(n2575), .A2(n3441), .ZN(n2080) );
  NAND2_X1 U2862 ( .A1(n2576), .A2(n3440), .ZN(n2081) );
  NAND2_X1 U2863 ( .A1(n2077), .A2(n2078), .ZN(n3729) );
  NAND3_X1 U2864 ( .A1(n2426), .A2(n2083), .A3(n2303), .ZN(n2826) );
  NOR2_X2 U2865 ( .A1(n2286), .A2(n2287), .ZN(n2303) );
  NOR2_X2 U2866 ( .A1(n2015), .A2(n2302), .ZN(n2083) );
  OR2_X2 U2867 ( .A1(n3369), .A2(n3627), .ZN(n3402) );
  NAND2_X1 U2868 ( .A1(n3309), .A2(n3310), .ZN(n3116) );
  INV_X1 U2869 ( .A(n2091), .ZN(n4096) );
  AND2_X2 U2870 ( .A1(n4274), .A2(n2045), .ZN(n4174) );
  INV_X1 U2871 ( .A(n3898), .ZN(n3897) );
  NAND2_X1 U2872 ( .A1(n2664), .A2(n2048), .ZN(n2718) );
  NAND2_X1 U2873 ( .A1(n2664), .A2(REG3_REG_21__SCAN_IN), .ZN(n2690) );
  NAND2_X1 U2874 ( .A1(n2497), .A2(n2025), .ZN(n2544) );
  NAND2_X1 U2875 ( .A1(n2101), .A2(n2415), .ZN(n2466) );
  NAND2_X1 U2876 ( .A1(n4270), .A2(n3798), .ZN(n2109) );
  NAND2_X1 U2877 ( .A1(n2109), .A2(n2110), .ZN(n4243) );
  NAND2_X1 U2878 ( .A1(n2113), .A2(n2998), .ZN(n4088) );
  NAND3_X1 U2879 ( .A1(n2122), .A2(n2004), .A3(n2126), .ZN(n2118) );
  NAND2_X1 U2880 ( .A1(n4014), .A2(n2126), .ZN(n2124) );
  NOR2_X1 U2881 ( .A1(n4032), .A2(n2999), .ZN(n4017) );
  INV_X1 U2882 ( .A(n2123), .ZN(n2125) );
  NAND2_X1 U2883 ( .A1(n2973), .A2(n3860), .ZN(n3301) );
  NAND2_X1 U2884 ( .A1(n2973), .A2(n2128), .ZN(n2127) );
  OAI21_X1 U2885 ( .B1(n3181), .B2(n2975), .A(n3785), .ZN(n3248) );
  NAND2_X1 U2886 ( .A1(n2975), .A2(n3785), .ZN(n2140) );
  OR2_X1 U2887 ( .A1(n2896), .A2(n4604), .ZN(n2142) );
  AOI21_X1 U2888 ( .B1(n2151), .B2(n2149), .A(n2024), .ZN(n2143) );
  NAND2_X1 U2889 ( .A1(n4469), .A2(n2150), .ZN(n2144) );
  XNOR2_X1 U2890 ( .A(n2888), .B(n2887), .ZN(n4469) );
  INV_X1 U2891 ( .A(n4540), .ZN(n2153) );
  NAND2_X1 U2892 ( .A1(n4540), .A2(n4541), .ZN(n4539) );
  INV_X1 U2893 ( .A(n2154), .ZN(n2152) );
  NAND2_X1 U2894 ( .A1(n2157), .A2(n2156), .ZN(n2160) );
  INV_X2 U2895 ( .A(IR_REG_0__SCAN_IN), .ZN(n2157) );
  NAND3_X1 U2896 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .A3(
        IR_REG_0__SCAN_IN), .ZN(n2159) );
  NAND2_X1 U2897 ( .A1(n2902), .A2(n2163), .ZN(n2161) );
  OAI21_X1 U2898 ( .B1(n4506), .B2(n2162), .A(n2161), .ZN(n4518) );
  NAND2_X1 U2899 ( .A1(n2368), .A2(n2369), .ZN(n2172) );
  NAND2_X1 U2900 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2174)
         );
  OR2_X1 U2901 ( .A1(n4537), .A2(n2179), .ZN(n2175) );
  NAND2_X1 U2902 ( .A1(n2175), .A2(n2176), .ZN(n3979) );
  NAND2_X1 U2903 ( .A1(n4537), .A2(n4538), .ZN(n4536) );
  NAND2_X1 U2904 ( .A1(n2858), .A2(n4500), .ZN(n2183) );
  OAI21_X1 U2905 ( .B1(n4502), .B2(n2185), .A(n2184), .ZN(n4514) );
  XNOR2_X2 U2906 ( .A(n2863), .B(n2901), .ZN(n4502) );
  AND2_X1 U2907 ( .A1(n4550), .A2(n2922), .ZN(n4284) );
  NAND2_X1 U2908 ( .A1(n2921), .A2(n4562), .ZN(n3768) );
  NAND2_X1 U2909 ( .A1(n4144), .A2(n2001), .ZN(n2187) );
  NAND2_X1 U2910 ( .A1(n2187), .A2(n2188), .ZN(n4103) );
  NAND3_X1 U2911 ( .A1(n2220), .A2(n2939), .A3(n2014), .ZN(n2203) );
  AND2_X1 U2912 ( .A1(n3364), .A2(n3292), .ZN(n2218) );
  NOR2_X1 U2913 ( .A1(n2965), .A2(n2221), .ZN(n2230) );
  NAND2_X1 U2914 ( .A1(n4086), .A2(n2038), .ZN(n2222) );
  NAND2_X1 U2915 ( .A1(n2239), .A2(n2009), .ZN(n2233) );
  NAND2_X1 U2916 ( .A1(n2239), .A2(n2264), .ZN(n3742) );
  NAND2_X1 U2917 ( .A1(n3242), .A2(n2027), .ZN(n2249) );
  AND2_X1 U2918 ( .A1(n2266), .A2(n2258), .ZN(n2256) );
  AND2_X1 U2919 ( .A1(n2257), .A2(n2272), .ZN(n2298) );
  NAND3_X1 U2920 ( .A1(n2257), .A2(n2272), .A3(n2285), .ZN(n2491) );
  OR2_X1 U2921 ( .A1(n2000), .A2(n2340), .ZN(n2344) );
  NAND2_X2 U2922 ( .A1(n2325), .A2(n3037), .ZN(n2437) );
  OR2_X1 U2923 ( .A1(n2317), .A2(n3033), .ZN(n2319) );
  NAND2_X1 U2924 ( .A1(n2291), .A2(n2290), .ZN(n2313) );
  INV_X1 U2925 ( .A(n2289), .ZN(n2291) );
  NAND2_X1 U2926 ( .A1(n3468), .A2(n2361), .ZN(n3428) );
  NOR2_X1 U2927 ( .A1(n4514), .A2(n2866), .ZN(n2868) );
  NAND2_X1 U2928 ( .A1(n4303), .A2(n3020), .ZN(n4313) );
  OR2_X1 U2929 ( .A1(n2491), .A2(IR_REG_9__SCAN_IN), .ZN(n2553) );
  NOR2_X1 U2930 ( .A1(n2872), .A2(n2685), .ZN(n4128) );
  MUX2_X1 U2931 ( .A(DATAI_3_), .B(n4460), .S(n2872), .Z(n3774) );
  OAI21_X1 U2932 ( .B1(n2872), .B2(n2347), .A(n2346), .ZN(n4571) );
  NAND2_X1 U2933 ( .A1(n2872), .A2(IR_REG_0__SCAN_IN), .ZN(n2346) );
  NAND2_X1 U2934 ( .A1(n2872), .A2(n2881), .ZN(n2334) );
  AND2_X1 U2935 ( .A1(n2463), .A2(n2462), .ZN(n2260) );
  OR2_X1 U2936 ( .A1(n3436), .A2(n4444), .ZN(n2261) );
  OR2_X1 U2937 ( .A1(n3436), .A2(n4379), .ZN(n2262) );
  OR2_X1 U2938 ( .A1(n4458), .A2(REG1_REG_7__SCAN_IN), .ZN(n2263) );
  INV_X1 U2939 ( .A(DATAI_0_), .ZN(n2347) );
  NAND2_X1 U2940 ( .A1(n3928), .A2(n3267), .ZN(n2940) );
  AND2_X1 U2941 ( .A1(n2737), .A2(n2736), .ZN(n2264) );
  OR2_X1 U2942 ( .A1(n3027), .A2(n2350), .ZN(n2265) );
  NOR2_X1 U2943 ( .A1(n2287), .A2(IR_REG_17__SCAN_IN), .ZN(n2267) );
  INV_X1 U2944 ( .A(n4307), .ZN(n4018) );
  INV_X1 U2945 ( .A(n3030), .ZN(n2846) );
  INV_X1 U2946 ( .A(n2976), .ZN(n3254) );
  NAND2_X2 U2947 ( .A1(n3123), .A2(n4276), .ZN(n4581) );
  OR2_X1 U2948 ( .A1(n4168), .A2(n2995), .ZN(n2268) );
  AND2_X1 U2949 ( .A1(n3615), .A2(n2677), .ZN(n2269) );
  INV_X1 U2950 ( .A(n3870), .ZN(n2945) );
  AND2_X1 U2951 ( .A1(n2805), .A2(n3764), .ZN(n2270) );
  AND2_X1 U2952 ( .A1(n2832), .A2(n2831), .ZN(n2271) );
  OR2_X1 U2953 ( .A1(n3156), .A2(n3157), .ZN(n2462) );
  AND2_X1 U2954 ( .A1(n3844), .A2(n4087), .ZN(n3891) );
  INV_X1 U2955 ( .A(IR_REG_24__SCAN_IN), .ZN(n3490) );
  OR2_X1 U2956 ( .A1(n4594), .A2(REG2_REG_17__SCAN_IN), .ZN(n2909) );
  AND2_X1 U2957 ( .A1(n3843), .A2(n4069), .ZN(n3892) );
  INV_X1 U2958 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2836) );
  AOI21_X1 U2959 ( .B1(n4535), .B2(ADDR_REG_18__SCAN_IN), .A(n3734), .ZN(n2915) );
  INV_X1 U2960 ( .A(n3444), .ZN(n3015) );
  INV_X1 U2961 ( .A(n3774), .ZN(n3310) );
  OAI21_X1 U2962 ( .B1(n2920), .B2(n2397), .A(n2337), .ZN(n2339) );
  OR2_X1 U2963 ( .A1(n3143), .A2(n2394), .ZN(n2395) );
  INV_X1 U2964 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U2965 ( .A1(n2320), .A2(REG3_REG_1__SCAN_IN), .ZN(n2329) );
  INV_X1 U2966 ( .A(n2915), .ZN(n2918) );
  OR2_X1 U2967 ( .A1(n3745), .A2(n4079), .ZN(n2963) );
  OR2_X1 U2968 ( .A1(n3132), .A2(n2825), .ZN(n2828) );
  INV_X1 U2969 ( .A(n3926), .ZN(n3714) );
  AND2_X1 U2970 ( .A1(n3044), .A2(n3011), .ZN(n3134) );
  OR2_X1 U2971 ( .A1(n4095), .A2(n2453), .ZN(n2710) );
  NOR2_X1 U2972 ( .A1(n3210), .A2(n3209), .ZN(n3208) );
  INV_X1 U2973 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3713) );
  INV_X1 U2974 ( .A(REG3_REG_16__SCAN_IN), .ZN(n3653) );
  INV_X1 U2975 ( .A(n4559), .ZN(n4264) );
  NAND2_X1 U2976 ( .A1(n4562), .A2(n3767), .ZN(n4565) );
  NOR2_X1 U2977 ( .A1(n2872), .A2(n2658), .ZN(n4165) );
  INV_X1 U2978 ( .A(n4573), .ZN(n4288) );
  NAND2_X1 U2979 ( .A1(n3027), .A2(n4591), .ZN(n3010) );
  NOR2_X1 U2980 ( .A1(n2872), .A2(n2697), .ZN(n3845) );
  XNOR2_X1 U2981 ( .A(n2392), .B(n2391), .ZN(n3143) );
  NAND2_X1 U2982 ( .A1(n3470), .A2(n3469), .ZN(n3468) );
  AND2_X1 U2983 ( .A1(n2815), .A2(n2814), .ZN(n3762) );
  INV_X1 U2984 ( .A(n2818), .ZN(n2797) );
  OR2_X1 U2985 ( .A1(n2000), .A2(n2398), .ZN(n2403) );
  AND2_X1 U2986 ( .A1(n4465), .A2(n3002), .ZN(n4509) );
  AOI21_X1 U2987 ( .B1(n2877), .B2(n2876), .A(n4513), .ZN(n2878) );
  INV_X1 U2988 ( .A(n2977), .ZN(n3267) );
  AND2_X1 U2989 ( .A1(n4215), .A2(n3020), .ZN(n4567) );
  INV_X1 U2990 ( .A(n4578), .ZN(n4276) );
  AOI21_X1 U2991 ( .B1(n3043), .B2(n2781), .A(n2780), .ZN(n3022) );
  OR2_X1 U2992 ( .A1(n4309), .A2(n4308), .ZN(n4310) );
  INV_X1 U2993 ( .A(n4629), .ZN(n4644) );
  AND2_X1 U2994 ( .A1(n4572), .A2(n2816), .ZN(n4641) );
  INV_X1 U2995 ( .A(n3010), .ZN(n3044) );
  NAND2_X1 U2996 ( .A1(n2307), .A2(n2306), .ZN(n3046) );
  XNOR2_X1 U2997 ( .A(n2614), .B(IR_REG_17__SCAN_IN), .ZN(n4594) );
  AND2_X1 U2998 ( .A1(n2914), .A2(n2913), .ZN(n4535) );
  NAND2_X1 U2999 ( .A1(n2797), .A2(n2796), .ZN(n3750) );
  INV_X1 U3000 ( .A(n4115), .ZN(n3920) );
  INV_X1 U3001 ( .A(n4460), .ZN(n3062) );
  INV_X1 U3002 ( .A(n4602), .ZN(n4500) );
  INV_X1 U3003 ( .A(n4509), .ZN(n4548) );
  INV_X1 U3004 ( .A(n4567), .ZN(n4234) );
  NAND2_X1 U3005 ( .A1(n4581), .A2(n3199), .ZN(n4283) );
  NAND2_X1 U3006 ( .A1(n4658), .A2(n3020), .ZN(n4379) );
  AND2_X2 U3007 ( .A1(n3023), .A2(n3022), .ZN(n4658) );
  NAND2_X1 U3008 ( .A1(n4647), .A2(n3020), .ZN(n4444) );
  INV_X1 U3009 ( .A(n4647), .ZN(n4646) );
  INV_X1 U3010 ( .A(n4590), .ZN(n4589) );
  NAND2_X1 U3011 ( .A1(n3045), .A2(n3044), .ZN(n4590) );
  INV_X1 U3012 ( .A(n3929), .ZN(U4043) );
  INV_X2 U3013 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3014 ( .A(n2491), .ZN(n2277) );
  NOR2_X1 U3015 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2276)
         );
  NAND4_X1 U3016 ( .A1(n2276), .A2(n2275), .A3(n2274), .A4(n2273), .ZN(n2287)
         );
  NAND2_X1 U3017 ( .A1(n2277), .A2(n2267), .ZN(n2631) );
  INV_X1 U3018 ( .A(IR_REG_19__SCAN_IN), .ZN(n2278) );
  NAND2_X1 U3019 ( .A1(n2338), .A2(n2278), .ZN(n2279) );
  NAND4_X1 U3020 ( .A1(n2285), .A2(n2284), .A3(n2283), .A4(n2282), .ZN(n2286)
         );
  NAND2_X1 U3021 ( .A1(n2298), .A2(n2297), .ZN(n2289) );
  NAND2_X1 U3022 ( .A1(n2289), .A2(IR_REG_31__SCAN_IN), .ZN(n2288) );
  MUX2_X1 U3023 ( .A(IR_REG_31__SCAN_IN), .B(n2288), .S(IR_REG_21__SCAN_IN), 
        .Z(n2292) );
  NAND2_X1 U3024 ( .A1(n2794), .A2(n2793), .ZN(n2293) );
  NAND4_X1 U3025 ( .A1(n2290), .A2(n2793), .A3(n3490), .A4(n2295), .ZN(n2302)
         );
  INV_X1 U3026 ( .A(n2302), .ZN(n2296) );
  NAND2_X1 U3027 ( .A1(n2299), .A2(n2298), .ZN(n2308) );
  NAND2_X1 U3028 ( .A1(n2308), .A2(IR_REG_31__SCAN_IN), .ZN(n2309) );
  MUX2_X1 U3029 ( .A(IR_REG_31__SCAN_IN), .B(n2309), .S(IR_REG_25__SCAN_IN), 
        .Z(n2310) );
  NOR2_X1 U3030 ( .A1(n3046), .A2(n2778), .ZN(n2311) );
  NAND2_X1 U3031 ( .A1(n2775), .A2(n2311), .ZN(n2349) );
  NAND2_X1 U3032 ( .A1(n2313), .A2(IR_REG_31__SCAN_IN), .ZN(n2314) );
  OR2_X4 U3033 ( .A1(n2367), .A2(n3020), .ZN(n2772) );
  NAND2_X1 U3034 ( .A1(n2317), .A2(n2318), .ZN(n3034) );
  XNOR2_X2 U3035 ( .A(n2316), .B(IR_REG_30__SCAN_IN), .ZN(n2323) );
  INV_X1 U3036 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2321) );
  OR2_X1 U3037 ( .A1(n2439), .A2(n2321), .ZN(n2328) );
  INV_X1 U3038 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2324) );
  INV_X1 U3039 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2835) );
  OR2_X1 U3040 ( .A1(n2437), .A2(n2835), .ZN(n2326) );
  NAND2_X1 U3041 ( .A1(n2874), .A2(IR_REG_28__SCAN_IN), .ZN(n2331) );
  INV_X4 U3042 ( .A(n2332), .ZN(n2872) );
  INV_X1 U3043 ( .A(DATAI_1_), .ZN(n2333) );
  BUF_X1 U3044 ( .A(n2880), .Z(n2881) );
  OAI21_X2 U3045 ( .B1(n2872), .B2(DATAI_1_), .A(n2334), .ZN(n4562) );
  INV_X1 U3046 ( .A(n2349), .ZN(n2335) );
  OAI22_X1 U3047 ( .A1(n2772), .A2(n2920), .B1(n4562), .B2(n2397), .ZN(n2359)
         );
  NAND2_X1 U3048 ( .A1(n2538), .A2(n2336), .ZN(n2337) );
  XNOR2_X1 U3049 ( .A(n2339), .B(n2674), .ZN(n2358) );
  XNOR2_X1 U3050 ( .A(n2359), .B(n2358), .ZN(n3470) );
  NAND2_X1 U3051 ( .A1(n2320), .A2(REG3_REG_0__SCAN_IN), .ZN(n2345) );
  INV_X1 U3052 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2340) );
  INV_X1 U3053 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2341) );
  OR2_X1 U3054 ( .A1(n2439), .A2(n2341), .ZN(n2343) );
  INV_X1 U3055 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2350) );
  OR2_X1 U3056 ( .A1(n2437), .A2(n2350), .ZN(n2342) );
  OR2_X1 U3057 ( .A1(n2367), .A2(n3767), .ZN(n2348) );
  OAI21_X1 U3058 ( .B1(n2397), .B2(n2354), .A(n2348), .ZN(n2355) );
  INV_X1 U3059 ( .A(n2355), .ZN(n2351) );
  OAI22_X1 U3060 ( .A1(n2397), .A2(n3767), .B1(n2157), .B2(n3027), .ZN(n2352)
         );
  NAND2_X1 U3061 ( .A1(n3131), .A2(n3130), .ZN(n2357) );
  OR2_X1 U3062 ( .A1(n2355), .A2(n2770), .ZN(n2356) );
  NAND2_X1 U3063 ( .A1(n2357), .A2(n2356), .ZN(n3469) );
  INV_X1 U3064 ( .A(n2358), .ZN(n2360) );
  NAND2_X1 U3065 ( .A1(n2360), .A2(n2359), .ZN(n2361) );
  INV_X1 U3066 ( .A(n3428), .ZN(n2374) );
  NAND2_X1 U3067 ( .A1(n2320), .A2(REG3_REG_2__SCAN_IN), .ZN(n2365) );
  OR2_X1 U3068 ( .A1(n2437), .A2(n2836), .ZN(n2364) );
  INV_X1 U3069 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2362) );
  OR2_X1 U3070 ( .A1(n2439), .A2(n2362), .ZN(n2363) );
  NAND2_X1 U3071 ( .A1(n2447), .A2(REG2_REG_2__SCAN_IN), .ZN(n2366) );
  INV_X1 U3072 ( .A(DATAI_2_), .ZN(n2370) );
  OR2_X1 U3073 ( .A1(n2367), .A2(n4287), .ZN(n2371) );
  OAI21_X1 U3074 ( .B1(n2397), .B2(n2923), .A(n2371), .ZN(n2372) );
  XNOR2_X1 U3075 ( .A(n2372), .B(n2770), .ZN(n2376) );
  OAI22_X1 U3076 ( .A1(n2772), .A2(n2923), .B1(n4287), .B2(n2397), .ZN(n2375)
         );
  XNOR2_X1 U3077 ( .A(n2376), .B(n2375), .ZN(n3426) );
  INV_X1 U3078 ( .A(n3426), .ZN(n2373) );
  NAND2_X1 U3079 ( .A1(n2374), .A2(n2373), .ZN(n3140) );
  OR2_X1 U3080 ( .A1(n2376), .A2(n2375), .ZN(n3141) );
  INV_X1 U3081 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3308) );
  OR2_X1 U3082 ( .A1(n2000), .A2(n3308), .ZN(n2383) );
  OR2_X1 U3083 ( .A1(n2453), .A2(REG3_REG_3__SCAN_IN), .ZN(n2382) );
  INV_X2 U3084 ( .A(n2439), .ZN(n2752) );
  NAND2_X1 U3085 ( .A1(n2752), .A2(REG0_REG_3__SCAN_IN), .ZN(n2380) );
  CLKBUF_X3 U3086 ( .A(n2437), .Z(n3831) );
  INV_X1 U3087 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2378) );
  OR2_X1 U3088 ( .A1(n3831), .A2(n2378), .ZN(n2379) );
  AND2_X1 U3089 ( .A1(n2380), .A2(n2379), .ZN(n2381) );
  NAND3_X1 U3090 ( .A1(n2383), .A2(n2382), .A3(n2381), .ZN(n2925) );
  INV_X1 U3091 ( .A(n2925), .ZN(n2926) );
  NAND2_X1 U3092 ( .A1(n2384), .A2(IR_REG_31__SCAN_IN), .ZN(n2386) );
  NAND2_X1 U3093 ( .A1(n2386), .A2(n2385), .ZN(n2404) );
  OR2_X1 U3094 ( .A1(n2386), .A2(n2385), .ZN(n2387) );
  OAI22_X1 U3095 ( .A1(n2772), .A2(n2926), .B1(n3310), .B2(n2397), .ZN(n2391)
         );
  INV_X1 U3096 ( .A(n2391), .ZN(n2389) );
  NAND2_X1 U3097 ( .A1(n2389), .A2(n2392), .ZN(n2393) );
  AND2_X1 U3098 ( .A1(n3141), .A2(n2393), .ZN(n2390) );
  NAND2_X1 U3099 ( .A1(n3140), .A2(n2390), .ZN(n2396) );
  INV_X1 U3100 ( .A(n2393), .ZN(n2394) );
  NAND2_X1 U3101 ( .A1(n2396), .A2(n2395), .ZN(n3407) );
  INV_X2 U3102 ( .A(n2397), .ZN(n2726) );
  INV_X1 U3103 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2398) );
  OR2_X1 U3104 ( .A1(n2439), .A2(n4628), .ZN(n2402) );
  OAI21_X1 U3105 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2417), .ZN(n3415) );
  OR2_X1 U3106 ( .A1(n2453), .A2(n3415), .ZN(n2401) );
  INV_X1 U3107 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4471) );
  OR2_X1 U3108 ( .A1(n2437), .A2(n4471), .ZN(n2400) );
  INV_X1 U3109 ( .A(n3934), .ZN(n2410) );
  INV_X1 U3110 ( .A(DATAI_4_), .ZN(n2407) );
  NAND2_X1 U3111 ( .A1(n2404), .A2(IR_REG_31__SCAN_IN), .ZN(n2406) );
  XNOR2_X1 U3112 ( .A(n2406), .B(n2405), .ZN(n2887) );
  MUX2_X1 U3113 ( .A(n2407), .B(n2887), .S(n2872), .Z(n3117) );
  OR2_X1 U3114 ( .A1(n2367), .A2(n3117), .ZN(n2408) );
  OAI21_X1 U3115 ( .B1(n2769), .B2(n2410), .A(n2408), .ZN(n2409) );
  XNOR2_X1 U3116 ( .A(n2409), .B(n2770), .ZN(n2413) );
  OAI22_X1 U3117 ( .A1(n2772), .A2(n2410), .B1(n3117), .B2(n2813), .ZN(n2412)
         );
  XNOR2_X1 U3118 ( .A(n2413), .B(n2412), .ZN(n3411) );
  INV_X1 U3119 ( .A(n3411), .ZN(n2411) );
  NAND2_X1 U3120 ( .A1(n3407), .A2(n2411), .ZN(n3408) );
  NAND2_X1 U3121 ( .A1(n2413), .A2(n2412), .ZN(n2414) );
  NAND2_X1 U3122 ( .A1(n3408), .A2(n2414), .ZN(n3660) );
  NAND2_X1 U3123 ( .A1(n2820), .A2(REG1_REG_5__SCAN_IN), .ZN(n2423) );
  INV_X1 U3124 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3224) );
  OR2_X1 U3125 ( .A1(n2000), .A2(n3224), .ZN(n2422) );
  INV_X1 U3126 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2416) );
  NAND2_X1 U3127 ( .A1(n2417), .A2(n2416), .ZN(n2418) );
  NAND2_X1 U3128 ( .A1(n2450), .A2(n2418), .ZN(n3662) );
  OR2_X1 U3129 ( .A1(n2453), .A2(n3662), .ZN(n2421) );
  INV_X1 U3130 ( .A(REG0_REG_5__SCAN_IN), .ZN(n2419) );
  OR2_X1 U3131 ( .A1(n2439), .A2(n2419), .ZN(n2420) );
  NAND2_X1 U3132 ( .A1(n2424), .A2(IR_REG_31__SCAN_IN), .ZN(n2425) );
  MUX2_X1 U3133 ( .A(IR_REG_31__SCAN_IN), .B(n2425), .S(IR_REG_5__SCAN_IN), 
        .Z(n2428) );
  INV_X1 U3134 ( .A(n2426), .ZN(n2427) );
  AND2_X1 U3135 ( .A1(n2428), .A2(n2427), .ZN(n3030) );
  MUX2_X1 U3136 ( .A(DATAI_5_), .B(n3030), .S(n2872), .Z(n3661) );
  INV_X1 U3137 ( .A(n3661), .ZN(n3221) );
  OR2_X1 U3138 ( .A1(n2367), .A2(n3221), .ZN(n2429) );
  OAI21_X1 U3139 ( .B1(n2769), .B2(n3333), .A(n2429), .ZN(n2430) );
  XNOR2_X1 U3140 ( .A(n2430), .B(n2674), .ZN(n2431) );
  OAI22_X1 U3141 ( .A1(n2772), .A2(n3333), .B1(n3221), .B2(n2769), .ZN(n2432)
         );
  XNOR2_X1 U3142 ( .A(n2431), .B(n2432), .ZN(n3659) );
  INV_X1 U3143 ( .A(n2431), .ZN(n2433) );
  NAND2_X1 U3144 ( .A1(n2433), .A2(n2432), .ZN(n2434) );
  NAND2_X1 U3145 ( .A1(n2447), .A2(REG2_REG_7__SCAN_IN), .ZN(n2443) );
  NAND2_X1 U3146 ( .A1(n2452), .A2(n2435), .ZN(n2436) );
  NAND2_X1 U3147 ( .A1(n2466), .A2(n2436), .ZN(n3189) );
  INV_X1 U31480 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2849) );
  OR2_X1 U31490 ( .A1(n2437), .A2(n2849), .ZN(n2441) );
  INV_X1 U3150 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2438) );
  OR2_X1 U3151 ( .A1(n2439), .A2(n2438), .ZN(n2440) );
  INV_X1 U3152 ( .A(n3931), .ZN(n3334) );
  INV_X1 U3153 ( .A(DATAI_7_), .ZN(n2444) );
  OR2_X1 U3154 ( .A1(n2298), .A2(n3033), .ZN(n2474) );
  MUX2_X1 U3155 ( .A(n2444), .B(n3076), .S(n2872), .Z(n3185) );
  OR2_X1 U3156 ( .A1(n2367), .A2(n3185), .ZN(n2445) );
  OAI21_X1 U3157 ( .B1(n2813), .B2(n3334), .A(n2445), .ZN(n2446) );
  XNOR2_X1 U3158 ( .A(n2446), .B(n2770), .ZN(n3161) );
  OAI22_X1 U3159 ( .A1(n2772), .A2(n3334), .B1(n3185), .B2(n2813), .ZN(n3162)
         );
  OR2_X1 U3160 ( .A1(n3161), .A2(n3162), .ZN(n2463) );
  NAND2_X1 U3161 ( .A1(n2447), .A2(REG2_REG_6__SCAN_IN), .ZN(n2458) );
  INV_X1 U3162 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2448) );
  OR2_X1 U3163 ( .A1(n2439), .A2(n2448), .ZN(n2457) );
  INV_X1 U3164 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2449) );
  NAND2_X1 U3165 ( .A1(n2450), .A2(n2449), .ZN(n2451) );
  NAND2_X1 U3166 ( .A1(n2452), .A2(n2451), .ZN(n3340) );
  OR2_X1 U3167 ( .A1(n2453), .A2(n3340), .ZN(n2456) );
  INV_X1 U3168 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2454) );
  INV_X1 U3169 ( .A(n3932), .ZN(n3196) );
  OR2_X1 U3170 ( .A1(n2426), .A2(n3033), .ZN(n2459) );
  MUX2_X1 U3171 ( .A(DATAI_6_), .B(n4459), .S(n2872), .Z(n3336) );
  OR2_X1 U3172 ( .A1(n2367), .A2(n3342), .ZN(n2460) );
  OAI21_X1 U3173 ( .B1(n2813), .B2(n3196), .A(n2460), .ZN(n2461) );
  XNOR2_X1 U3174 ( .A(n2461), .B(n2770), .ZN(n3156) );
  OAI22_X1 U3175 ( .A1(n2772), .A2(n3196), .B1(n3342), .B2(n2813), .ZN(n3157)
         );
  AND2_X1 U3176 ( .A1(n3156), .A2(n3157), .ZN(n2464) );
  AOI22_X1 U3177 ( .A1(n2464), .A2(n2463), .B1(n3161), .B2(n3162), .ZN(n2465)
         );
  NAND2_X1 U3178 ( .A1(n2820), .A2(REG1_REG_8__SCAN_IN), .ZN(n2472) );
  INV_X1 U3179 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3257) );
  OR2_X1 U3180 ( .A1(n2000), .A2(n3257), .ZN(n2471) );
  NAND2_X1 U3181 ( .A1(n2466), .A2(n3092), .ZN(n2467) );
  NAND2_X1 U3182 ( .A1(n2485), .A2(n2467), .ZN(n3256) );
  OR2_X1 U3183 ( .A1(n2453), .A2(n3256), .ZN(n2470) );
  INV_X1 U3184 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2468) );
  OR2_X1 U3185 ( .A1(n2439), .A2(n2468), .ZN(n2469) );
  INV_X1 U3186 ( .A(DATAI_8_), .ZN(n2477) );
  NAND2_X1 U3187 ( .A1(n2474), .A2(n2473), .ZN(n2475) );
  NAND2_X1 U3188 ( .A1(n2475), .A2(IR_REG_31__SCAN_IN), .ZN(n2476) );
  MUX2_X1 U3189 ( .A(n2477), .B(n4456), .S(n2872), .Z(n2976) );
  OR2_X1 U3190 ( .A1(n2768), .A2(n2976), .ZN(n2478) );
  OAI21_X1 U3191 ( .B1(n2813), .B2(n3262), .A(n2478), .ZN(n2479) );
  XNOR2_X1 U3192 ( .A(n2479), .B(n2770), .ZN(n2481) );
  OAI22_X1 U3193 ( .A1(n2772), .A2(n3262), .B1(n2976), .B2(n2769), .ZN(n2480)
         );
  AND2_X1 U3194 ( .A1(n2481), .A2(n2480), .ZN(n3172) );
  OR2_X1 U3195 ( .A1(n2481), .A2(n2480), .ZN(n3171) );
  NAND2_X1 U3196 ( .A1(n2482), .A2(n3171), .ZN(n3231) );
  NAND2_X1 U3197 ( .A1(n2752), .A2(REG0_REG_9__SCAN_IN), .ZN(n2490) );
  INV_X1 U3198 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3581) );
  OR2_X1 U3199 ( .A1(n2000), .A2(n3581), .ZN(n2489) );
  INV_X1 U3200 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2484) );
  NAND2_X1 U3201 ( .A1(n2485), .A2(n2484), .ZN(n2486) );
  NAND2_X1 U3202 ( .A1(n2498), .A2(n2486), .ZN(n3268) );
  OR2_X1 U3203 ( .A1(n2453), .A2(n3268), .ZN(n2488) );
  INV_X1 U3204 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2854) );
  OR2_X1 U3205 ( .A1(n3831), .A2(n2854), .ZN(n2487) );
  INV_X1 U3206 ( .A(DATAI_9_), .ZN(n2494) );
  NAND2_X1 U3207 ( .A1(n2491), .A2(IR_REG_31__SCAN_IN), .ZN(n2492) );
  MUX2_X1 U3208 ( .A(IR_REG_31__SCAN_IN), .B(n2492), .S(IR_REG_9__SCAN_IN), 
        .Z(n2493) );
  NAND2_X1 U3209 ( .A1(n2493), .A2(n2553), .ZN(n3101) );
  MUX2_X1 U32100 ( .A(n2494), .B(n3101), .S(n2872), .Z(n2977) );
  OR2_X1 U32110 ( .A1(n2367), .A2(n2977), .ZN(n2495) );
  OAI21_X1 U32120 ( .B1(n2813), .B2(n3316), .A(n2495), .ZN(n2496) );
  XNOR2_X1 U32130 ( .A(n2496), .B(n2674), .ZN(n2508) );
  OAI22_X1 U32140 ( .A1(n2772), .A2(n3316), .B1(n2977), .B2(n2769), .ZN(n2509)
         );
  XNOR2_X1 U32150 ( .A(n2508), .B(n2509), .ZN(n3232) );
  NAND2_X1 U32160 ( .A1(n3231), .A2(n3232), .ZN(n3242) );
  NAND2_X1 U32170 ( .A1(n2752), .A2(REG0_REG_10__SCAN_IN), .ZN(n2503) );
  INV_X1 U32180 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4484) );
  OR2_X1 U32190 ( .A1(n3831), .A2(n4484), .ZN(n2502) );
  INV_X1 U32200 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3326) );
  OR2_X1 U32210 ( .A1(n2000), .A2(n3326), .ZN(n2501) );
  NAND2_X1 U32220 ( .A1(n2498), .A2(n2100), .ZN(n2499) );
  NAND2_X1 U32230 ( .A1(n2516), .A2(n2499), .ZN(n3325) );
  OR2_X1 U32240 ( .A1(n2453), .A2(n3325), .ZN(n2500) );
  INV_X1 U32250 ( .A(DATAI_10_), .ZN(n2505) );
  NAND2_X1 U32260 ( .A1(n2553), .A2(IR_REG_31__SCAN_IN), .ZN(n2504) );
  XNOR2_X1 U32270 ( .A(n2504), .B(n2551), .ZN(n4604) );
  MUX2_X1 U32280 ( .A(n2505), .B(n4604), .S(n2872), .Z(n3323) );
  OR2_X1 U32290 ( .A1(n2367), .A2(n3323), .ZN(n2506) );
  OAI21_X1 U32300 ( .B1(n2769), .B2(n3285), .A(n2506), .ZN(n2507) );
  XNOR2_X1 U32310 ( .A(n2507), .B(n2674), .ZN(n2512) );
  OAI22_X1 U32320 ( .A1(n2772), .A2(n3285), .B1(n3323), .B2(n2813), .ZN(n2513)
         );
  XNOR2_X1 U32330 ( .A(n2512), .B(n2513), .ZN(n3240) );
  INV_X1 U32340 ( .A(n2508), .ZN(n2510) );
  OR2_X1 U32350 ( .A1(n2510), .A2(n2509), .ZN(n3241) );
  AND2_X1 U32360 ( .A1(n3240), .A2(n3241), .ZN(n2511) );
  INV_X1 U32370 ( .A(n2512), .ZN(n2514) );
  NAND2_X1 U32380 ( .A1(n2514), .A2(n2513), .ZN(n2515) );
  NAND2_X1 U32390 ( .A1(n2820), .A2(REG1_REG_11__SCAN_IN), .ZN(n2522) );
  INV_X1 U32400 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3554) );
  OR2_X1 U32410 ( .A1(n2000), .A2(n3554), .ZN(n2521) );
  NAND2_X1 U32420 ( .A1(n2516), .A2(n3205), .ZN(n2517) );
  NAND2_X1 U32430 ( .A1(n2532), .A2(n2517), .ZN(n3293) );
  OR2_X1 U32440 ( .A1(n2453), .A2(n3293), .ZN(n2520) );
  INV_X1 U32450 ( .A(REG0_REG_11__SCAN_IN), .ZN(n2518) );
  OR2_X1 U32460 ( .A1(n2764), .A2(n2518), .ZN(n2519) );
  NAND2_X1 U32470 ( .A1(n2523), .A2(IR_REG_31__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U32480 ( .A1(n2524), .A2(n3532), .ZN(n2539) );
  INV_X1 U32490 ( .A(DATAI_11_), .ZN(n2525) );
  MUX2_X1 U32500 ( .A(n3207), .B(n2525), .S(n1999), .Z(n3292) );
  OR2_X1 U32510 ( .A1(n3292), .A2(n2367), .ZN(n2526) );
  OAI21_X1 U32520 ( .B1(n2813), .B2(n3364), .A(n2526), .ZN(n2527) );
  XNOR2_X1 U32530 ( .A(n2527), .B(n2770), .ZN(n2529) );
  OAI22_X1 U32540 ( .A1(n2772), .A2(n3364), .B1(n3292), .B2(n2813), .ZN(n2528)
         );
  AND2_X1 U32550 ( .A1(n2529), .A2(n2528), .ZN(n3274) );
  INV_X1 U32560 ( .A(n2528), .ZN(n2531) );
  INV_X1 U32570 ( .A(n2529), .ZN(n2530) );
  NAND2_X1 U32580 ( .A1(n2531), .A2(n2530), .ZN(n3273) );
  NAND2_X1 U32590 ( .A1(n2447), .A2(REG2_REG_12__SCAN_IN), .ZN(n2537) );
  INV_X1 U32600 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4442) );
  OR2_X1 U32610 ( .A1(n2764), .A2(n4442), .ZN(n2536) );
  INV_X1 U32620 ( .A(REG3_REG_12__SCAN_IN), .ZN(n3628) );
  NAND2_X1 U32630 ( .A1(n2532), .A2(n3628), .ZN(n2533) );
  NAND2_X1 U32640 ( .A1(n2544), .A2(n2533), .ZN(n3629) );
  OR2_X1 U32650 ( .A1(n2453), .A2(n3629), .ZN(n2535) );
  INV_X1 U32660 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4493) );
  OR2_X1 U32670 ( .A1(n3831), .A2(n4493), .ZN(n2534) );
  NAND4_X1 U32680 ( .A1(n2537), .A2(n2536), .A3(n2535), .A4(n2534), .ZN(n3926)
         );
  NAND2_X1 U32690 ( .A1(n2539), .A2(IR_REG_31__SCAN_IN), .ZN(n2540) );
  MUX2_X1 U32700 ( .A(n4602), .B(DATAI_12_), .S(n1999), .Z(n3627) );
  NAND2_X1 U32710 ( .A1(n2538), .A2(n3627), .ZN(n2541) );
  OAI21_X1 U32720 ( .B1(n3714), .B2(n2813), .A(n2541), .ZN(n2542) );
  XNOR2_X1 U32730 ( .A(n2542), .B(n2674), .ZN(n3625) );
  INV_X1 U32740 ( .A(n3627), .ZN(n2979) );
  OAI22_X1 U32750 ( .A1(n2772), .A2(n3714), .B1(n2979), .B2(n2769), .ZN(n2543)
         );
  INV_X1 U32760 ( .A(n2543), .ZN(n3624) );
  NAND2_X1 U32770 ( .A1(n2544), .A2(n3713), .ZN(n2545) );
  AND2_X1 U32780 ( .A1(n2564), .A2(n2545), .ZN(n3716) );
  NAND2_X1 U32790 ( .A1(n3716), .A2(n2320), .ZN(n2549) );
  NAND2_X1 U32800 ( .A1(n2820), .A2(REG1_REG_13__SCAN_IN), .ZN(n2548) );
  INV_X1 U32810 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3571) );
  OR2_X1 U32820 ( .A1(n2000), .A2(n3571), .ZN(n2547) );
  INV_X1 U32830 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4438) );
  OR2_X1 U32840 ( .A1(n2764), .A2(n4438), .ZN(n2546) );
  INV_X1 U32850 ( .A(DATAI_13_), .ZN(n3535) );
  INV_X1 U32860 ( .A(IR_REG_12__SCAN_IN), .ZN(n2550) );
  NAND3_X1 U32870 ( .A1(n3532), .A2(n2551), .A3(n2550), .ZN(n2552) );
  NOR2_X1 U32880 ( .A1(n2555), .A2(n3033), .ZN(n2554) );
  MUX2_X1 U32890 ( .A(n3033), .B(n2554), .S(IR_REG_13__SCAN_IN), .Z(n2557) );
  INV_X1 U32900 ( .A(n2577), .ZN(n2556) );
  MUX2_X1 U32910 ( .A(n3535), .B(n3977), .S(n2872), .Z(n3394) );
  OAI22_X1 U32920 ( .A1(n3380), .A2(n2769), .B1(n2768), .B2(n3394), .ZN(n2558)
         );
  XNOR2_X1 U32930 ( .A(n2558), .B(n2770), .ZN(n2559) );
  OAI22_X1 U32940 ( .A1(n2772), .A2(n3380), .B1(n3394), .B2(n2813), .ZN(n2560)
         );
  AND2_X1 U32950 ( .A1(n2559), .A2(n2560), .ZN(n3709) );
  INV_X1 U32960 ( .A(n2559), .ZN(n2562) );
  INV_X1 U32970 ( .A(n2560), .ZN(n2561) );
  NAND2_X1 U32980 ( .A1(n2562), .A2(n2561), .ZN(n3708) );
  NAND2_X1 U32990 ( .A1(n2564), .A2(n2563), .ZN(n2565) );
  NAND2_X1 U33000 ( .A1(n2593), .A2(n2565), .ZN(n3446) );
  INV_X1 U33010 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3385) );
  OR2_X1 U33020 ( .A1(n2000), .A2(n3385), .ZN(n2568) );
  INV_X1 U33030 ( .A(REG0_REG_14__SCAN_IN), .ZN(n2566) );
  OR2_X1 U33040 ( .A1(n2764), .A2(n2566), .ZN(n2567) );
  AND2_X1 U33050 ( .A1(n2568), .A2(n2567), .ZN(n2570) );
  INV_X1 U33060 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4503) );
  OR2_X1 U33070 ( .A1(n3831), .A2(n4503), .ZN(n2569) );
  OAI211_X1 U33080 ( .C1(n3446), .C2(n2453), .A(n2570), .B(n2569), .ZN(n3924)
         );
  INV_X1 U33090 ( .A(n3924), .ZN(n4265) );
  NAND2_X1 U33100 ( .A1(n2577), .A2(IR_REG_31__SCAN_IN), .ZN(n2571) );
  XNOR2_X1 U33110 ( .A(n2571), .B(IR_REG_14__SCAN_IN), .ZN(n4600) );
  MUX2_X1 U33120 ( .A(DATAI_14_), .B(n4600), .S(n2872), .Z(n3444) );
  NAND2_X1 U33130 ( .A1(n2538), .A2(n3444), .ZN(n2572) );
  OAI21_X1 U33140 ( .B1(n4265), .B2(n2769), .A(n2572), .ZN(n2573) );
  XNOR2_X1 U33150 ( .A(n2573), .B(n2674), .ZN(n2574) );
  NAND2_X1 U33160 ( .A1(n3443), .A2(n2574), .ZN(n2576) );
  OAI22_X1 U33170 ( .A1(n2772), .A2(n4265), .B1(n3015), .B2(n2769), .ZN(n3440)
         );
  INV_X1 U33180 ( .A(n3443), .ZN(n2575) );
  INV_X1 U33190 ( .A(n2574), .ZN(n3441) );
  INV_X1 U33200 ( .A(DATAI_16_), .ZN(n4596) );
  INV_X1 U33210 ( .A(IR_REG_15__SCAN_IN), .ZN(n2579) );
  NAND2_X1 U33220 ( .A1(n2599), .A2(n2579), .ZN(n2580) );
  NAND2_X1 U33230 ( .A1(n2580), .A2(IR_REG_31__SCAN_IN), .ZN(n2582) );
  INV_X1 U33240 ( .A(IR_REG_16__SCAN_IN), .ZN(n2581) );
  MUX2_X1 U33250 ( .A(n4596), .B(n4597), .S(n2872), .Z(n4248) );
  NAND2_X1 U33260 ( .A1(n2595), .A2(n3653), .ZN(n2583) );
  AND2_X1 U33270 ( .A1(n2016), .A2(n2583), .ZN(n4249) );
  NAND2_X1 U33280 ( .A1(n4249), .A2(n2320), .ZN(n2588) );
  INV_X1 U33290 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4525) );
  NAND2_X1 U33300 ( .A1(n2752), .A2(REG0_REG_16__SCAN_IN), .ZN(n2585) );
  NAND2_X1 U33310 ( .A1(n2447), .A2(REG2_REG_16__SCAN_IN), .ZN(n2584) );
  OAI211_X1 U33320 ( .C1(n3831), .C2(n4525), .A(n2585), .B(n2584), .ZN(n2586)
         );
  INV_X1 U33330 ( .A(n2586), .ZN(n2587) );
  NAND2_X1 U33340 ( .A1(n3922), .A2(n2726), .ZN(n2589) );
  OAI21_X1 U33350 ( .B1(n4248), .B2(n2768), .A(n2589), .ZN(n2590) );
  XNOR2_X1 U33360 ( .A(n2590), .B(n2674), .ZN(n3672) );
  INV_X1 U33370 ( .A(n3672), .ZN(n2605) );
  NAND2_X1 U33380 ( .A1(n2716), .A2(n3922), .ZN(n2592) );
  OR2_X1 U33390 ( .A1(n4248), .A2(n2769), .ZN(n2591) );
  NAND2_X1 U33400 ( .A1(n2592), .A2(n2591), .ZN(n2618) );
  INV_X1 U33410 ( .A(REG0_REG_15__SCAN_IN), .ZN(n2598) );
  INV_X1 U33420 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3530) );
  NAND2_X1 U33430 ( .A1(n2593), .A2(n3530), .ZN(n2594) );
  NAND2_X1 U33440 ( .A1(n2595), .A2(n2594), .ZN(n4277) );
  OR2_X1 U33450 ( .A1(n4277), .A2(n2453), .ZN(n2597) );
  AOI22_X1 U33460 ( .A1(n2820), .A2(REG1_REG_15__SCAN_IN), .B1(n2447), .B2(
        REG2_REG_15__SCAN_IN), .ZN(n2596) );
  NAND2_X1 U33470 ( .A1(n2716), .A2(n3923), .ZN(n2601) );
  MUX2_X1 U33480 ( .A(DATAI_15_), .B(n2903), .S(n2872), .Z(n4275) );
  NAND2_X1 U33490 ( .A1(n2726), .A2(n4275), .ZN(n2600) );
  NAND2_X1 U33500 ( .A1(n2601), .A2(n2600), .ZN(n3669) );
  NAND2_X1 U33510 ( .A1(n2726), .A2(n3923), .ZN(n2603) );
  NAND2_X1 U33520 ( .A1(n2538), .A2(n4275), .ZN(n2602) );
  NAND2_X1 U3353 ( .A1(n2603), .A2(n2602), .ZN(n2604) );
  XNOR2_X1 U33540 ( .A(n2604), .B(n2770), .ZN(n2617) );
  AOI22_X1 U3355 ( .A1(n2605), .A2(n2618), .B1(n3669), .B2(n2617), .ZN(n2622)
         );
  NAND2_X1 U3356 ( .A1(n2016), .A2(n2106), .ZN(n2607) );
  NAND2_X1 U3357 ( .A1(n2624), .A2(n2607), .ZN(n4235) );
  OR2_X1 U3358 ( .A1(n4235), .A2(n2453), .ZN(n2612) );
  INV_X1 U3359 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4356) );
  NAND2_X1 U3360 ( .A1(n2752), .A2(REG0_REG_17__SCAN_IN), .ZN(n2609) );
  INV_X1 U3361 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4236) );
  OR2_X1 U3362 ( .A1(n2000), .A2(n4236), .ZN(n2608) );
  OAI211_X1 U3363 ( .C1(n4356), .C2(n3831), .A(n2609), .B(n2608), .ZN(n2610)
         );
  INV_X1 U3364 ( .A(n2610), .ZN(n2611) );
  OR2_X1 U3365 ( .A1(n2491), .A2(n2287), .ZN(n2613) );
  NAND2_X1 U3366 ( .A1(n2613), .A2(IR_REG_31__SCAN_IN), .ZN(n2614) );
  MUX2_X1 U3367 ( .A(DATAI_17_), .B(n4594), .S(n2872), .Z(n4231) );
  INV_X1 U3368 ( .A(n4231), .ZN(n4223) );
  OAI22_X1 U3369 ( .A1(n4242), .A2(n2769), .B1(n4223), .B2(n2768), .ZN(n2615)
         );
  XNOR2_X1 U3370 ( .A(n2615), .B(n2770), .ZN(n3674) );
  OAI22_X1 U3371 ( .A1(n4242), .A2(n2772), .B1(n4223), .B2(n2813), .ZN(n3673)
         );
  OAI21_X1 U3372 ( .B1(n2617), .B2(n3669), .A(n2618), .ZN(n2616) );
  NAND2_X1 U3373 ( .A1(n2616), .A2(n3672), .ZN(n2620) );
  INV_X1 U3374 ( .A(n2617), .ZN(n3651) );
  INV_X1 U3375 ( .A(n2618), .ZN(n3671) );
  INV_X1 U3376 ( .A(n3669), .ZN(n3755) );
  NAND3_X1 U3377 ( .A1(n3651), .A2(n3671), .A3(n3755), .ZN(n2619) );
  OAI211_X1 U3378 ( .C1(n3674), .C2(n3673), .A(n2620), .B(n2619), .ZN(n2621)
         );
  NAND2_X1 U3379 ( .A1(n2624), .A2(n2623), .ZN(n2625) );
  NAND2_X1 U3380 ( .A1(n2640), .A2(n2625), .ZN(n4217) );
  OR2_X1 U3381 ( .A1(n4217), .A2(n2453), .ZN(n2630) );
  INV_X1 U3382 ( .A(REG1_REG_18__SCAN_IN), .ZN(n2871) );
  NAND2_X1 U3383 ( .A1(n2447), .A2(REG2_REG_18__SCAN_IN), .ZN(n2627) );
  INV_X1 U3384 ( .A(REG0_REG_18__SCAN_IN), .ZN(n3534) );
  OR2_X1 U3385 ( .A1(n2764), .A2(n3534), .ZN(n2626) );
  OAI211_X1 U3386 ( .C1(n2871), .C2(n3831), .A(n2627), .B(n2626), .ZN(n2628)
         );
  INV_X1 U3387 ( .A(n2628), .ZN(n2629) );
  NAND2_X1 U3388 ( .A1(n2631), .A2(IR_REG_31__SCAN_IN), .ZN(n2632) );
  XNOR2_X1 U3389 ( .A(n2632), .B(IR_REG_18__SCAN_IN), .ZN(n4592) );
  MUX2_X1 U3390 ( .A(DATAI_18_), .B(n4592), .S(n2872), .Z(n4204) );
  INV_X1 U3391 ( .A(n4204), .ZN(n4213) );
  OAI22_X1 U3392 ( .A1(n4186), .A2(n2813), .B1(n4213), .B2(n2367), .ZN(n2633)
         );
  XNOR2_X1 U3393 ( .A(n2633), .B(n2674), .ZN(n2638) );
  INV_X1 U3394 ( .A(n2638), .ZN(n2636) );
  NOR2_X1 U3395 ( .A1(n2769), .A2(n4213), .ZN(n2634) );
  AOI21_X1 U3396 ( .B1(n4225), .B2(n2716), .A(n2634), .ZN(n2637) );
  INV_X1 U3397 ( .A(n2637), .ZN(n2635) );
  NAND2_X1 U3398 ( .A1(n2636), .A2(n2635), .ZN(n3730) );
  AND2_X1 U3399 ( .A1(n2638), .A2(n2637), .ZN(n3731) );
  NAND2_X1 U3400 ( .A1(n2640), .A2(n2639), .ZN(n2641) );
  NAND2_X1 U3401 ( .A1(n2651), .A2(n2641), .ZN(n3462) );
  INV_X1 U3402 ( .A(n3462), .ZN(n4196) );
  NAND2_X1 U3403 ( .A1(n4196), .A2(n2320), .ZN(n2647) );
  INV_X1 U3404 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2644) );
  NAND2_X1 U3405 ( .A1(n2820), .A2(REG1_REG_19__SCAN_IN), .ZN(n2643) );
  NAND2_X1 U3406 ( .A1(n2752), .A2(REG0_REG_19__SCAN_IN), .ZN(n2642) );
  OAI211_X1 U3407 ( .C1(n2000), .C2(n2644), .A(n2643), .B(n2642), .ZN(n2645)
         );
  INV_X1 U3408 ( .A(n2645), .ZN(n2646) );
  MUX2_X1 U3409 ( .A(DATAI_19_), .B(n3982), .S(n2872), .Z(n3460) );
  OAI22_X1 U3410 ( .A1(n4207), .A2(n2769), .B1(n4193), .B2(n2768), .ZN(n2648)
         );
  XNOR2_X1 U3411 ( .A(n2648), .B(n2770), .ZN(n2650) );
  OAI22_X1 U3412 ( .A1(n4207), .A2(n2772), .B1(n4193), .B2(n2769), .ZN(n2649)
         );
  XNOR2_X1 U3413 ( .A(n2650), .B(n2649), .ZN(n3459) );
  NAND2_X1 U3414 ( .A1(n2651), .A2(n3700), .ZN(n2652) );
  AND2_X1 U3415 ( .A1(n2666), .A2(n2652), .ZN(n4177) );
  NAND2_X1 U3416 ( .A1(n4177), .A2(n2320), .ZN(n2657) );
  INV_X1 U3417 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4344) );
  NAND2_X1 U3418 ( .A1(n2752), .A2(REG0_REG_20__SCAN_IN), .ZN(n2654) );
  NAND2_X1 U3419 ( .A1(n2447), .A2(REG2_REG_20__SCAN_IN), .ZN(n2653) );
  OAI211_X1 U3420 ( .C1(n3831), .C2(n4344), .A(n2654), .B(n2653), .ZN(n2655)
         );
  INV_X1 U3421 ( .A(n2655), .ZN(n2656) );
  INV_X1 U3422 ( .A(DATAI_20_), .ZN(n2658) );
  NOR2_X1 U3423 ( .A1(n2768), .A2(n4176), .ZN(n2659) );
  AOI21_X1 U3424 ( .B1(n4188), .B2(n2726), .A(n2659), .ZN(n2660) );
  XNOR2_X1 U3425 ( .A(n2660), .B(n2770), .ZN(n2663) );
  NOR2_X1 U3426 ( .A1(n2813), .A2(n4176), .ZN(n2661) );
  AOI21_X1 U3427 ( .B1(n4188), .B2(n2716), .A(n2661), .ZN(n2662) );
  OR2_X1 U3428 ( .A1(n2663), .A2(n2662), .ZN(n3696) );
  NAND2_X1 U3429 ( .A1(n2663), .A2(n2662), .ZN(n3698) );
  INV_X1 U3430 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2665) );
  NAND2_X1 U3431 ( .A1(n2666), .A2(n2665), .ZN(n2667) );
  NAND2_X1 U3432 ( .A1(n2690), .A2(n2667), .ZN(n4146) );
  INV_X1 U3433 ( .A(REG0_REG_21__SCAN_IN), .ZN(n2670) );
  NAND2_X1 U3434 ( .A1(n2820), .A2(REG1_REG_21__SCAN_IN), .ZN(n2669) );
  NAND2_X1 U3435 ( .A1(n2447), .A2(REG2_REG_21__SCAN_IN), .ZN(n2668) );
  OAI211_X1 U3436 ( .C1(n2670), .C2(n2764), .A(n2669), .B(n2668), .ZN(n2671)
         );
  INV_X1 U3437 ( .A(n2671), .ZN(n2672) );
  NAND2_X1 U3438 ( .A1(n1999), .A2(DATAI_21_), .ZN(n2995) );
  OAI22_X1 U3439 ( .A1(n4168), .A2(n2769), .B1(n2995), .B2(n2768), .ZN(n2675)
         );
  XNOR2_X1 U3440 ( .A(n2675), .B(n2674), .ZN(n3615) );
  NOR2_X1 U3441 ( .A1(n2769), .A2(n2995), .ZN(n2676) );
  AOI21_X1 U3442 ( .B1(n4129), .B2(n2716), .A(n2676), .ZN(n2677) );
  INV_X1 U3443 ( .A(n3615), .ZN(n2678) );
  INV_X1 U3444 ( .A(n2677), .ZN(n3614) );
  XNOR2_X1 U3445 ( .A(n2690), .B(REG3_REG_22__SCAN_IN), .ZN(n4137) );
  NAND2_X1 U3446 ( .A1(n4137), .A2(n2320), .ZN(n2684) );
  INV_X1 U3447 ( .A(REG1_REG_22__SCAN_IN), .ZN(n2681) );
  NAND2_X1 U3448 ( .A1(n2752), .A2(REG0_REG_22__SCAN_IN), .ZN(n2680) );
  NAND2_X1 U3449 ( .A1(n2447), .A2(REG2_REG_22__SCAN_IN), .ZN(n2679) );
  OAI211_X1 U3450 ( .C1(n3831), .C2(n2681), .A(n2680), .B(n2679), .ZN(n2682)
         );
  INV_X1 U3451 ( .A(n2682), .ZN(n2683) );
  INV_X1 U3452 ( .A(DATAI_22_), .ZN(n2685) );
  AOI22_X1 U3453 ( .A1(n4149), .A2(n2716), .B1(n4128), .B2(n2726), .ZN(n2702)
         );
  AOI22_X1 U3454 ( .A1(n4149), .A2(n2726), .B1(n4128), .B2(n2538), .ZN(n2686)
         );
  XNOR2_X1 U3455 ( .A(n2686), .B(n2770), .ZN(n2703) );
  XOR2_X1 U3456 ( .A(n2702), .B(n2703), .Z(n3722) );
  INV_X1 U3457 ( .A(REG3_REG_22__SCAN_IN), .ZN(n2688) );
  INV_X1 U34580 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2687) );
  OAI21_X1 U34590 ( .B1(n2690), .B2(n2688), .A(n2687), .ZN(n2691) );
  NAND2_X1 U3460 ( .A1(REG3_REG_23__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2689) );
  AND2_X1 U3461 ( .A1(n2691), .A2(n2704), .ZN(n4122) );
  NAND2_X1 U3462 ( .A1(n4122), .A2(n2320), .ZN(n2696) );
  INV_X1 U3463 ( .A(REG2_REG_23__SCAN_IN), .ZN(n3558) );
  NAND2_X1 U3464 ( .A1(n2820), .A2(REG1_REG_23__SCAN_IN), .ZN(n2693) );
  NAND2_X1 U3465 ( .A1(n2752), .A2(REG0_REG_23__SCAN_IN), .ZN(n2692) );
  OAI211_X1 U3466 ( .C1(n2000), .C2(n3558), .A(n2693), .B(n2692), .ZN(n2694)
         );
  INV_X1 U34670 ( .A(n2694), .ZN(n2695) );
  NAND2_X1 U3468 ( .A1(n3921), .A2(n2726), .ZN(n2699) );
  INV_X1 U34690 ( .A(DATAI_23_), .ZN(n2697) );
  INV_X1 U3470 ( .A(n3845), .ZN(n4120) );
  OR2_X1 U34710 ( .A1(n2768), .A2(n4120), .ZN(n2698) );
  NAND2_X1 U3472 ( .A1(n2699), .A2(n2698), .ZN(n2700) );
  XNOR2_X1 U34730 ( .A(n2700), .B(n2770), .ZN(n2714) );
  NOR2_X1 U3474 ( .A1(n2769), .A2(n4120), .ZN(n2701) );
  AOI21_X1 U34750 ( .B1(n3921), .B2(n2716), .A(n2701), .ZN(n2712) );
  XNOR2_X1 U3476 ( .A(n2714), .B(n2712), .ZN(n3452) );
  NAND2_X1 U34770 ( .A1(n2703), .A2(n2702), .ZN(n3451) );
  INV_X1 U3478 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3688) );
  NAND2_X1 U34790 ( .A1(n2704), .A2(n3688), .ZN(n2705) );
  NAND2_X1 U3480 ( .A1(n2718), .A2(n2705), .ZN(n4095) );
  INV_X1 U34810 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4328) );
  NAND2_X1 U3482 ( .A1(n2752), .A2(REG0_REG_24__SCAN_IN), .ZN(n2707) );
  NAND2_X1 U34830 ( .A1(n2447), .A2(REG2_REG_24__SCAN_IN), .ZN(n2706) );
  OAI211_X1 U3484 ( .C1(n3831), .C2(n4328), .A(n2707), .B(n2706), .ZN(n2708)
         );
  INV_X1 U34850 ( .A(n2708), .ZN(n2709) );
  NAND2_X1 U3486 ( .A1(n1999), .A2(DATAI_24_), .ZN(n4098) );
  OAI22_X1 U34870 ( .A1(n4115), .A2(n2813), .B1(n4098), .B2(n2367), .ZN(n2711)
         );
  XNOR2_X1 U3488 ( .A(n2711), .B(n2770), .ZN(n3685) );
  INV_X1 U34890 ( .A(n2712), .ZN(n2713) );
  NAND2_X1 U3490 ( .A1(n2714), .A2(n2713), .ZN(n3638) );
  INV_X1 U34910 ( .A(n3638), .ZN(n2717) );
  NOR2_X1 U3492 ( .A1(n2769), .A2(n4098), .ZN(n2715) );
  AOI21_X1 U34930 ( .B1(n3920), .B2(n2716), .A(n2715), .ZN(n3637) );
  NAND2_X1 U3494 ( .A1(n3637), .A2(n3638), .ZN(n3635) );
  OAI21_X1 U34950 ( .B1(n3685), .B2(n2717), .A(n3635), .ZN(n2731) );
  INV_X1 U3496 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3645) );
  NAND2_X1 U34970 ( .A1(n2718), .A2(n3645), .ZN(n2719) );
  NAND2_X1 U3498 ( .A1(n4081), .A2(n2320), .ZN(n2725) );
  INV_X1 U34990 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2722) );
  NAND2_X1 U3500 ( .A1(n2820), .A2(REG1_REG_25__SCAN_IN), .ZN(n2721) );
  NAND2_X1 U35010 ( .A1(n2752), .A2(REG0_REG_25__SCAN_IN), .ZN(n2720) );
  OAI211_X1 U3502 ( .C1(n2000), .C2(n2722), .A(n2721), .B(n2720), .ZN(n2723)
         );
  INV_X1 U35030 ( .A(n2723), .ZN(n2724) );
  NAND2_X1 U3504 ( .A1(n4092), .A2(n2726), .ZN(n2729) );
  INV_X1 U35050 ( .A(DATAI_25_), .ZN(n2727) );
  NOR2_X1 U35060 ( .A1(n2872), .A2(n2727), .ZN(n3016) );
  INV_X1 U35070 ( .A(n3016), .ZN(n4079) );
  OR2_X1 U35080 ( .A1(n2367), .A2(n4079), .ZN(n2728) );
  NAND2_X1 U35090 ( .A1(n2729), .A2(n2728), .ZN(n2730) );
  XNOR2_X1 U35100 ( .A(n2730), .B(n2770), .ZN(n3642) );
  OAI22_X1 U35110 ( .A1(n3745), .A2(n2772), .B1(n4079), .B2(n2769), .ZN(n3641)
         );
  NAND2_X1 U35120 ( .A1(n3642), .A2(n3641), .ZN(n3640) );
  INV_X1 U35130 ( .A(n3685), .ZN(n2735) );
  INV_X1 U35140 ( .A(n3641), .ZN(n2734) );
  AOI21_X1 U35150 ( .B1(n2735), .B2(n3637), .A(n2734), .ZN(n2733) );
  NAND3_X1 U35160 ( .A1(n2735), .A2(n3637), .A3(n2734), .ZN(n2736) );
  INV_X1 U35170 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3743) );
  NAND2_X1 U35180 ( .A1(n2738), .A2(n3743), .ZN(n2739) );
  NAND2_X1 U35190 ( .A1(n4063), .A2(n2320), .ZN(n2744) );
  INV_X1 U35200 ( .A(REG2_REG_26__SCAN_IN), .ZN(n3557) );
  NAND2_X1 U35210 ( .A1(n2820), .A2(REG1_REG_26__SCAN_IN), .ZN(n2741) );
  NAND2_X1 U35220 ( .A1(n2752), .A2(REG0_REG_26__SCAN_IN), .ZN(n2740) );
  OAI211_X1 U35230 ( .C1(n2000), .C2(n3557), .A(n2741), .B(n2740), .ZN(n2742)
         );
  INV_X1 U35240 ( .A(n2742), .ZN(n2743) );
  NAND2_X1 U35250 ( .A1(n1999), .A2(DATAI_26_), .ZN(n4061) );
  OAI22_X1 U35260 ( .A1(n4033), .A2(n2769), .B1(n4061), .B2(n2768), .ZN(n2745)
         );
  XNOR2_X1 U35270 ( .A(n2745), .B(n2770), .ZN(n2747) );
  OAI22_X1 U35280 ( .A1(n4033), .A2(n2772), .B1(n4061), .B2(n2769), .ZN(n2746)
         );
  NAND2_X1 U35290 ( .A1(n2747), .A2(n2746), .ZN(n3740) );
  INV_X1 U35300 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2749) );
  NAND2_X1 U35310 ( .A1(n2750), .A2(n2749), .ZN(n2751) );
  NAND2_X1 U35320 ( .A1(n2760), .A2(n2751), .ZN(n4044) );
  INV_X1 U35330 ( .A(REG1_REG_27__SCAN_IN), .ZN(n2755) );
  NAND2_X1 U35340 ( .A1(n2447), .A2(REG2_REG_27__SCAN_IN), .ZN(n2754) );
  NAND2_X1 U35350 ( .A1(n2752), .A2(REG0_REG_27__SCAN_IN), .ZN(n2753) );
  OAI211_X1 U35360 ( .C1(n2755), .C2(n3831), .A(n2754), .B(n2753), .ZN(n2756)
         );
  INV_X1 U35370 ( .A(n2756), .ZN(n2757) );
  INV_X1 U35380 ( .A(DATAI_27_), .ZN(n3516) );
  NOR2_X1 U35390 ( .A1(n2872), .A2(n3516), .ZN(n3420) );
  OAI22_X1 U35400 ( .A1(n4058), .A2(n2772), .B1(n4041), .B2(n2813), .ZN(n2799)
         );
  OAI22_X1 U35410 ( .A1(n4058), .A2(n2813), .B1(n4041), .B2(n2367), .ZN(n2759)
         );
  XNOR2_X1 U35420 ( .A(n2759), .B(n2770), .ZN(n2800) );
  XOR2_X1 U35430 ( .A(n2799), .B(n2800), .Z(n3418) );
  INV_X1 U35440 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2819) );
  NAND2_X1 U35450 ( .A1(n2760), .A2(n2819), .ZN(n2761) );
  NAND2_X1 U35460 ( .A1(n3434), .A2(n2320), .ZN(n2767) );
  INV_X1 U35470 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3529) );
  NAND2_X1 U35480 ( .A1(n2820), .A2(REG1_REG_28__SCAN_IN), .ZN(n2763) );
  NAND2_X1 U35490 ( .A1(n2447), .A2(REG2_REG_28__SCAN_IN), .ZN(n2762) );
  OAI211_X1 U35500 ( .C1(n2764), .C2(n3529), .A(n2763), .B(n2762), .ZN(n2765)
         );
  INV_X1 U35510 ( .A(n2765), .ZN(n2766) );
  INV_X1 U35520 ( .A(DATAI_28_), .ZN(n3524) );
  NOR2_X1 U35530 ( .A1(n2872), .A2(n3524), .ZN(n4010) );
  INV_X1 U35540 ( .A(n4010), .ZN(n3018) );
  OAI22_X1 U35550 ( .A1(n4036), .A2(n2769), .B1(n3018), .B2(n2768), .ZN(n2771)
         );
  XNOR2_X1 U35560 ( .A(n2771), .B(n2770), .ZN(n2774) );
  OAI22_X1 U35570 ( .A1(n4036), .A2(n2772), .B1(n3018), .B2(n2813), .ZN(n2773)
         );
  XNOR2_X1 U35580 ( .A(n2774), .B(n2773), .ZN(n2805) );
  INV_X1 U35590 ( .A(n2775), .ZN(n3047) );
  INV_X1 U35600 ( .A(n2778), .ZN(n4450) );
  OR2_X1 U35610 ( .A1(n2775), .A2(n4450), .ZN(n2776) );
  MUX2_X1 U35620 ( .A(n3047), .B(n2776), .S(B_REG_SCAN_IN), .Z(n2777) );
  NAND2_X1 U35630 ( .A1(n3043), .A2(n3503), .ZN(n2779) );
  NAND2_X1 U35640 ( .A1(n3046), .A2(n2778), .ZN(n3049) );
  NAND2_X1 U35650 ( .A1(n2779), .A2(n3049), .ZN(n3009) );
  INV_X1 U35660 ( .A(n3009), .ZN(n3120) );
  INV_X1 U35670 ( .A(D_REG_0__SCAN_IN), .ZN(n2781) );
  NOR2_X1 U35680 ( .A1(n2775), .A2(n4449), .ZN(n2780) );
  INV_X1 U35690 ( .A(D_REG_4__SCAN_IN), .ZN(n4587) );
  INV_X1 U35700 ( .A(D_REG_22__SCAN_IN), .ZN(n4585) );
  NAND2_X1 U35710 ( .A1(n4587), .A2(n4585), .ZN(n3479) );
  INV_X1 U35720 ( .A(n3479), .ZN(n2785) );
  NOR4_X1 U35730 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_31__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n2784) );
  NOR4_X1 U35740 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2783) );
  NOR4_X1 U35750 ( .A1(D_REG_3__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2782) );
  AND4_X1 U35760 ( .A1(n2785), .A2(n2784), .A3(n2783), .A4(n2782), .ZN(n2791)
         );
  NOR4_X1 U35770 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n2789) );
  NOR4_X1 U35780 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2788) );
  NOR4_X1 U35790 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n2787) );
  NOR4_X1 U35800 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2786) );
  AND4_X1 U35810 ( .A1(n2789), .A2(n2788), .A3(n2787), .A4(n2786), .ZN(n2790)
         );
  NAND2_X1 U3582 ( .A1(n2791), .A2(n2790), .ZN(n2792) );
  NAND2_X1 U3583 ( .A1(n3043), .A2(n2792), .ZN(n3012) );
  NAND3_X1 U3584 ( .A1(n3120), .A2(n3022), .A3(n3012), .ZN(n3132) );
  XNOR2_X1 U3585 ( .A(n2794), .B(n2793), .ZN(n2873) );
  INV_X1 U3586 ( .A(n2312), .ZN(n4453) );
  AOI21_X1 U3587 ( .B1(n3982), .B2(n4570), .A(n3003), .ZN(n2806) );
  INV_X1 U3588 ( .A(n2806), .ZN(n2795) );
  NOR2_X1 U3589 ( .A1(n4273), .A2(n2795), .ZN(n2796) );
  NAND2_X1 U3590 ( .A1(n2798), .A2(n2270), .ZN(n2834) );
  NAND2_X1 U3591 ( .A1(n3419), .A2(n3418), .ZN(n2802) );
  INV_X1 U3592 ( .A(n2805), .ZN(n2801) );
  NAND2_X1 U3593 ( .A1(n2800), .A2(n2799), .ZN(n2803) );
  NAND4_X1 U3594 ( .A1(n2802), .A2(n3764), .A3(n2801), .A4(n2803), .ZN(n2833)
         );
  INV_X1 U3595 ( .A(n2803), .ZN(n2804) );
  NAND3_X1 U3596 ( .A1(n2805), .A2(n3764), .A3(n2804), .ZN(n2832) );
  OR2_X1 U3597 ( .A1(n4273), .A2(n2806), .ZN(n3133) );
  NAND2_X1 U3598 ( .A1(n2312), .A2(n3987), .ZN(n2807) );
  NAND2_X1 U3599 ( .A1(n2807), .A2(n3003), .ZN(n3011) );
  NAND3_X1 U3600 ( .A1(n3011), .A2(n3027), .A3(n2873), .ZN(n2808) );
  AOI21_X1 U3601 ( .B1(n3132), .B2(n3133), .A(n2808), .ZN(n2809) );
  OR2_X1 U3602 ( .A1(n2809), .A2(U3149), .ZN(n2815) );
  INV_X1 U3603 ( .A(n2810), .ZN(n2811) );
  NAND2_X1 U3604 ( .A1(n2811), .A2(n4591), .ZN(n2812) );
  INV_X1 U3605 ( .A(n2825), .ZN(n3914) );
  NAND2_X1 U3606 ( .A1(n3132), .A2(n3914), .ZN(n2814) );
  NOR2_X1 U3607 ( .A1(n3010), .A2(n4452), .ZN(n2817) );
  OAI22_X1 U3608 ( .A1(n3702), .A2(n3018), .B1(STATE_REG_SCAN_IN), .B2(n2819), 
        .ZN(n2830) );
  INV_X1 U3609 ( .A(n4025), .ZN(n2824) );
  INV_X1 U3610 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3527) );
  NAND2_X1 U3611 ( .A1(n2447), .A2(REG2_REG_29__SCAN_IN), .ZN(n2822) );
  NAND2_X1 U3612 ( .A1(n2820), .A2(REG1_REG_29__SCAN_IN), .ZN(n2821) );
  OAI211_X1 U3613 ( .C1(n3527), .C2(n2764), .A(n2822), .B(n2821), .ZN(n2823)
         );
  OAI21_X1 U3614 ( .B1(n2826), .B2(IR_REG_27__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2827) );
  XNOR2_X1 U3615 ( .A(n2827), .B(IR_REG_28__SCAN_IN), .ZN(n4448) );
  INV_X1 U3616 ( .A(n4448), .ZN(n3002) );
  OAI22_X1 U3617 ( .A1(n3840), .A2(n3701), .B1(n4058), .B2(n3744), .ZN(n2829)
         );
  AOI211_X1 U3618 ( .C1(n3434), .C2(n3747), .A(n2830), .B(n2829), .ZN(n2831)
         );
  NAND3_X1 U3619 ( .A1(n2834), .A2(n2833), .A3(n2271), .ZN(U3217) );
  INV_X1 U3620 ( .A(n3207), .ZN(n2897) );
  MUX2_X1 U3621 ( .A(n2835), .B(REG1_REG_1__SCAN_IN), .S(n2880), .Z(n3936) );
  AND2_X1 U3622 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3937)
         );
  OR2_X1 U3623 ( .A1(n2881), .A2(n2835), .ZN(n3956) );
  NAND2_X1 U3624 ( .A1(n3935), .A2(n3956), .ZN(n2839) );
  OAI21_X1 U3625 ( .B1(n2879), .B2(n2836), .A(n2837), .ZN(n3957) );
  INV_X1 U3626 ( .A(n3957), .ZN(n2838) );
  NAND2_X1 U3627 ( .A1(n4461), .A2(REG1_REG_2__SCAN_IN), .ZN(n2840) );
  NAND2_X1 U3628 ( .A1(n3056), .A2(REG1_REG_3__SCAN_IN), .ZN(n2843) );
  NAND2_X1 U3629 ( .A1(n2841), .A2(n4460), .ZN(n2842) );
  XNOR2_X2 U3630 ( .A(n2844), .B(n2887), .ZN(n4472) );
  INV_X1 U3631 ( .A(n2887), .ZN(n4474) );
  INV_X1 U3632 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4653) );
  MUX2_X1 U3633 ( .A(n4653), .B(REG1_REG_5__SCAN_IN), .S(n3030), .Z(n3085) );
  INV_X1 U3634 ( .A(n2847), .ZN(n2848) );
  AOI22_X2 U3635 ( .A1(n3063), .A2(REG1_REG_6__SCAN_IN), .B1(n4459), .B2(n2848), .ZN(n3072) );
  NAND2_X1 U3636 ( .A1(n3072), .A2(n2850), .ZN(n2851) );
  INV_X1 U3637 ( .A(n3076), .ZN(n4458) );
  NAND2_X1 U3638 ( .A1(n2851), .A2(n2263), .ZN(n2852) );
  XNOR2_X1 U3639 ( .A(n2852), .B(n4457), .ZN(n3095) );
  NAND2_X1 U3640 ( .A1(n3095), .A2(REG1_REG_8__SCAN_IN), .ZN(n3094) );
  OR2_X1 U3641 ( .A1(n2852), .A2(n4456), .ZN(n2853) );
  NAND2_X1 U3642 ( .A1(n3094), .A2(n2853), .ZN(n3105) );
  XNOR2_X1 U3643 ( .A(n3101), .B(REG1_REG_9__SCAN_IN), .ZN(n3104) );
  NAND2_X1 U3644 ( .A1(n3105), .A2(n3104), .ZN(n3103) );
  NAND2_X1 U3645 ( .A1(n3103), .A2(n2855), .ZN(n2856) );
  INV_X1 U3646 ( .A(n4604), .ZN(n2895) );
  XNOR2_X1 U3647 ( .A(n2856), .B(n2895), .ZN(n4483) );
  AND2_X1 U3648 ( .A1(n2856), .A2(n2895), .ZN(n2857) );
  XNOR2_X1 U3649 ( .A(n2897), .B(REG1_REG_11__SCAN_IN), .ZN(n3209) );
  AOI21_X2 U3650 ( .B1(REG1_REG_11__SCAN_IN), .B2(n2897), .A(n3208), .ZN(n2858) );
  INV_X1 U3651 ( .A(n3977), .ZN(n4454) );
  NAND2_X1 U3652 ( .A1(n4454), .A2(REG1_REG_13__SCAN_IN), .ZN(n2862) );
  INV_X1 U3653 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4374) );
  NAND2_X1 U3654 ( .A1(n3977), .A2(n4374), .ZN(n2860) );
  NAND2_X1 U3655 ( .A1(n2862), .A2(n2860), .ZN(n3971) );
  INV_X1 U3656 ( .A(n4600), .ZN(n2901) );
  NOR2_X1 U3657 ( .A1(n2863), .A2(n2901), .ZN(n2864) );
  INV_X1 U3658 ( .A(n2903), .ZN(n4599) );
  INV_X1 U3659 ( .A(REG1_REG_15__SCAN_IN), .ZN(n2865) );
  AOI22_X1 U3660 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4599), .B1(n2903), .B2(
        n2865), .ZN(n4515) );
  AND2_X1 U3661 ( .A1(n2903), .A2(REG1_REG_15__SCAN_IN), .ZN(n2866) );
  INV_X1 U3662 ( .A(n4597), .ZN(n2867) );
  XNOR2_X1 U3663 ( .A(n2868), .B(n2867), .ZN(n4526) );
  NAND2_X1 U3664 ( .A1(n2868), .A2(n4597), .ZN(n2869) );
  NAND2_X1 U3665 ( .A1(n4524), .A2(n2869), .ZN(n4537) );
  INV_X1 U3666 ( .A(n4594), .ZN(n4549) );
  AOI22_X1 U3667 ( .A1(n4594), .A2(REG1_REG_17__SCAN_IN), .B1(n4356), .B2(
        n4549), .ZN(n4538) );
  OR2_X1 U3668 ( .A1(n4594), .A2(REG1_REG_17__SCAN_IN), .ZN(n2870) );
  INV_X1 U3669 ( .A(n4592), .ZN(n2916) );
  AOI22_X1 U3670 ( .A1(REG1_REG_18__SCAN_IN), .A2(n2916), .B1(n4592), .B2(
        n2871), .ZN(n2876) );
  OR2_X1 U3671 ( .A1(n2873), .A2(U3149), .ZN(n3917) );
  NAND2_X1 U3672 ( .A1(n3010), .A2(n3917), .ZN(n2914) );
  AOI21_X1 U3673 ( .B1(n2873), .B2(n3003), .A(n2872), .ZN(n2912) );
  XNOR2_X1 U3674 ( .A(n2875), .B(n2874), .ZN(n3993) );
  INV_X1 U3675 ( .A(n3993), .ZN(n4463) );
  AND2_X1 U3676 ( .A1(n4463), .A2(n4448), .ZN(n3947) );
  NAND2_X1 U3677 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4592), .ZN(n3980) );
  OAI21_X1 U3678 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4592), .A(n3980), .ZN(n2911) );
  INV_X1 U3679 ( .A(REG2_REG_2__SCAN_IN), .ZN(n4292) );
  AND2_X1 U3680 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3946)
         );
  OR2_X1 U3681 ( .A1(n2881), .A2(n2324), .ZN(n3950) );
  NAND2_X1 U3682 ( .A1(n3951), .A2(n3950), .ZN(n2882) );
  NAND2_X1 U3683 ( .A1(n4461), .A2(REG2_REG_2__SCAN_IN), .ZN(n2883) );
  NAND2_X1 U3684 ( .A1(n3954), .A2(n2883), .ZN(n2884) );
  XNOR2_X1 U3685 ( .A(n2884), .B(n3062), .ZN(n3057) );
  NAND2_X1 U3686 ( .A1(n3057), .A2(REG2_REG_3__SCAN_IN), .ZN(n2886) );
  NAND2_X1 U3687 ( .A1(n2884), .A2(n4460), .ZN(n2885) );
  NAND2_X1 U3688 ( .A1(n2886), .A2(n2885), .ZN(n2888) );
  MUX2_X1 U3689 ( .A(n3224), .B(REG2_REG_5__SCAN_IN), .S(n3030), .Z(n3082) );
  XNOR2_X1 U3690 ( .A(n2889), .B(n4459), .ZN(n3064) );
  INV_X1 U3691 ( .A(n2889), .ZN(n2890) );
  INV_X1 U3692 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3570) );
  MUX2_X1 U3693 ( .A(REG2_REG_7__SCAN_IN), .B(n3570), .S(n3076), .Z(n3073) );
  INV_X1 U3694 ( .A(n2893), .ZN(n2894) );
  XNOR2_X1 U3695 ( .A(n3101), .B(REG2_REG_9__SCAN_IN), .ZN(n3099) );
  INV_X1 U3696 ( .A(n3101), .ZN(n4455) );
  XNOR2_X1 U3697 ( .A(n3207), .B(REG2_REG_11__SCAN_IN), .ZN(n3204) );
  NOR2_X1 U3698 ( .A1(n3977), .A2(n3571), .ZN(n3963) );
  NOR2_X1 U3699 ( .A1(n4454), .A2(REG2_REG_13__SCAN_IN), .ZN(n3964) );
  INV_X1 U3700 ( .A(n3964), .ZN(n2899) );
  NOR2_X1 U3701 ( .A1(n2901), .A2(n2900), .ZN(n2902) );
  INV_X1 U3702 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4278) );
  AOI22_X1 U3703 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4599), .B1(n2903), .B2(
        n4278), .ZN(n4519) );
  AND2_X1 U3704 ( .A1(n2903), .A2(REG2_REG_15__SCAN_IN), .ZN(n2904) );
  INV_X1 U3705 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4528) );
  INV_X1 U3706 ( .A(n2905), .ZN(n2906) );
  NAND2_X1 U3707 ( .A1(n2906), .A2(n4597), .ZN(n2907) );
  NOR2_X1 U3708 ( .A1(n4594), .A2(REG2_REG_17__SCAN_IN), .ZN(n2908) );
  AOI21_X1 U3709 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4594), .A(n2908), .ZN(n4541) );
  INV_X1 U3710 ( .A(n2912), .ZN(n2913) );
  AND2_X1 U3711 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n3734) );
  NOR2_X1 U3712 ( .A1(n4548), .A2(n2916), .ZN(n2917) );
  NOR2_X1 U3713 ( .A1(n2918), .A2(n2917), .ZN(n2919) );
  NAND2_X1 U3714 ( .A1(n2921), .A2(n2336), .ZN(n2922) );
  INV_X1 U3715 ( .A(n4558), .ZN(n2923) );
  NAND2_X2 U3716 ( .A1(n2923), .A2(n4293), .ZN(n3770) );
  NAND2_X1 U3717 ( .A1(n4558), .A2(n4287), .ZN(n3772) );
  NAND2_X1 U3718 ( .A1(n4284), .A2(n2971), .ZN(n4285) );
  NAND2_X1 U3719 ( .A1(n2923), .A2(n4287), .ZN(n2924) );
  NAND2_X1 U3720 ( .A1(n4285), .A2(n2924), .ZN(n3297) );
  NOR2_X1 U3721 ( .A1(n2925), .A2(n3774), .ZN(n2927) );
  NAND2_X1 U3722 ( .A1(n3333), .A2(n3221), .ZN(n2932) );
  NAND2_X1 U3723 ( .A1(n3931), .A2(n3185), .ZN(n3785) );
  OAI21_X1 U3724 ( .B1(n3336), .B2(n3932), .A(n3180), .ZN(n2934) );
  INV_X1 U3725 ( .A(n2934), .ZN(n2928) );
  NAND2_X1 U3726 ( .A1(n3109), .A2(n2929), .ZN(n2938) );
  AND2_X1 U3727 ( .A1(n3932), .A2(n3336), .ZN(n2930) );
  INV_X1 U3728 ( .A(n3185), .ZN(n3188) );
  AOI22_X1 U3729 ( .A1(n3180), .A2(n2930), .B1(n3188), .B2(n3931), .ZN(n2936)
         );
  NAND2_X1 U3730 ( .A1(n3933), .A2(n3661), .ZN(n2931) );
  NAND2_X1 U3731 ( .A1(n3934), .A2(n3412), .ZN(n3215) );
  NAND2_X1 U3732 ( .A1(n2933), .A2(n2932), .ZN(n3192) );
  OR2_X1 U3733 ( .A1(n2934), .A2(n3192), .ZN(n2935) );
  AND2_X1 U3734 ( .A1(n2936), .A2(n2935), .ZN(n2937) );
  NAND2_X1 U3735 ( .A1(n2938), .A2(n2937), .ZN(n3249) );
  NOR2_X1 U3736 ( .A1(n3262), .A2(n2976), .ZN(n2939) );
  INV_X1 U3737 ( .A(n3323), .ZN(n3318) );
  INV_X1 U3738 ( .A(n3292), .ZN(n3287) );
  NAND2_X1 U3739 ( .A1(n3364), .A2(n3287), .ZN(n3361) );
  INV_X1 U3740 ( .A(n3364), .ZN(n3631) );
  NAND2_X1 U3741 ( .A1(n3631), .A2(n3292), .ZN(n3803) );
  NAND2_X1 U3742 ( .A1(n3361), .A2(n3803), .ZN(n3283) );
  OR2_X1 U3743 ( .A1(n3926), .A2(n3627), .ZN(n2941) );
  NAND2_X1 U3744 ( .A1(n3368), .A2(n2941), .ZN(n2943) );
  NAND2_X1 U3745 ( .A1(n3627), .A2(n3926), .ZN(n2942) );
  NAND2_X1 U3746 ( .A1(n2943), .A2(n2942), .ZN(n3396) );
  NAND2_X1 U3747 ( .A1(n3394), .A2(n3380), .ZN(n2944) );
  INV_X1 U3748 ( .A(n3394), .ZN(n3712) );
  AOI21_X1 U3749 ( .B1(n3396), .B2(n2944), .A(n2039), .ZN(n3376) );
  NAND2_X1 U3750 ( .A1(n3015), .A2(n3924), .ZN(n3797) );
  NAND2_X1 U3751 ( .A1(n4265), .A2(n3444), .ZN(n3808) );
  NAND2_X1 U3752 ( .A1(n3797), .A2(n3808), .ZN(n3870) );
  NAND2_X1 U3753 ( .A1(n3923), .A2(n4275), .ZN(n4253) );
  NOR2_X1 U3754 ( .A1(n2945), .A2(n4255), .ZN(n2946) );
  NAND2_X1 U3755 ( .A1(n3376), .A2(n2946), .ZN(n2949) );
  OR2_X1 U3756 ( .A1(n4248), .A2(n3922), .ZN(n3885) );
  NAND2_X1 U3757 ( .A1(n4248), .A2(n3922), .ZN(n4104) );
  NAND2_X1 U3758 ( .A1(n3885), .A2(n4104), .ZN(n4256) );
  OR2_X1 U3759 ( .A1(n3444), .A2(n3924), .ZN(n4261) );
  INV_X1 U3760 ( .A(n4261), .ZN(n2947) );
  INV_X1 U3761 ( .A(n4275), .ZN(n2988) );
  INV_X1 U3762 ( .A(n3923), .ZN(n4241) );
  AOI22_X1 U3763 ( .A1(n2947), .A2(n4253), .B1(n2988), .B2(n4241), .ZN(n4254)
         );
  NAND2_X1 U3764 ( .A1(n2949), .A2(n2948), .ZN(n2951) );
  INV_X1 U3765 ( .A(n3922), .ZN(n4266) );
  OR2_X1 U3766 ( .A1(n4266), .A2(n4248), .ZN(n2950) );
  NAND2_X1 U3767 ( .A1(n4242), .A2(n4223), .ZN(n2952) );
  NAND2_X1 U3768 ( .A1(n4186), .A2(n4204), .ZN(n2989) );
  NAND2_X1 U3769 ( .A1(n4225), .A2(n4213), .ZN(n4182) );
  NAND2_X1 U3770 ( .A1(n2989), .A2(n4182), .ZN(n4211) );
  NAND2_X1 U3771 ( .A1(n4166), .A2(n3460), .ZN(n2954) );
  NAND2_X1 U3772 ( .A1(n4158), .A2(n2035), .ZN(n2956) );
  INV_X1 U3773 ( .A(n4188), .ZN(n2990) );
  NAND2_X1 U3774 ( .A1(n2956), .A2(n2955), .ZN(n4144) );
  XNOR2_X1 U3775 ( .A(n4149), .B(n4128), .ZN(n4134) );
  INV_X1 U3776 ( .A(n4134), .ZN(n2957) );
  NAND2_X1 U3777 ( .A1(n4103), .A2(n2958), .ZN(n2960) );
  NAND2_X1 U3778 ( .A1(n3921), .A2(n3845), .ZN(n2959) );
  NOR2_X1 U3779 ( .A1(n4115), .A2(n4098), .ZN(n2962) );
  NAND2_X1 U3780 ( .A1(n4115), .A2(n4098), .ZN(n2961) );
  NOR2_X1 U3781 ( .A1(n4092), .A2(n3016), .ZN(n2964) );
  NOR2_X1 U3782 ( .A1(n4033), .A2(n4061), .ZN(n2965) );
  NOR2_X1 U3783 ( .A1(n3919), .A2(n3420), .ZN(n2966) );
  NAND2_X1 U3784 ( .A1(n4015), .A2(n4014), .ZN(n4008) );
  XNOR2_X1 U3785 ( .A(n4009), .B(n4008), .ZN(n3432) );
  XNOR2_X1 U3786 ( .A(n3126), .B(n4451), .ZN(n2967) );
  INV_X1 U3787 ( .A(n4641), .ZN(n4388) );
  NOR2_X1 U3788 ( .A1(n2969), .A2(n3767), .ZN(n4554) );
  NAND2_X1 U3789 ( .A1(n4555), .A2(n4554), .ZN(n4553) );
  NAND2_X1 U3790 ( .A1(n4553), .A2(n2970), .ZN(n2972) );
  INV_X1 U3791 ( .A(n2971), .ZN(n3850) );
  NAND2_X1 U3792 ( .A1(n2972), .A2(n3850), .ZN(n3298) );
  NAND2_X1 U3793 ( .A1(n3298), .A2(n3770), .ZN(n2973) );
  XNOR2_X1 U3794 ( .A(n2925), .B(n3774), .ZN(n3860) );
  OR2_X1 U3795 ( .A1(n3310), .A2(n2925), .ZN(n3775) );
  AND2_X1 U3796 ( .A1(n3933), .A2(n3221), .ZN(n3217) );
  OR2_X1 U3797 ( .A1(n3221), .A2(n3933), .ZN(n3792) );
  NAND2_X1 U3798 ( .A1(n3932), .A2(n3342), .ZN(n3791) );
  NAND2_X1 U3799 ( .A1(n3331), .A2(n3791), .ZN(n2974) );
  OR2_X1 U3800 ( .A1(n3342), .A2(n3932), .ZN(n3781) );
  INV_X1 U3801 ( .A(n3782), .ZN(n2975) );
  OR2_X1 U3802 ( .A1(n2976), .A2(n3930), .ZN(n3786) );
  NAND2_X1 U3803 ( .A1(n3930), .A2(n2976), .ZN(n3784) );
  AND2_X1 U3804 ( .A1(n3928), .A2(n2977), .ZN(n3793) );
  OR2_X1 U3805 ( .A1(n2977), .A2(n3928), .ZN(n3787) );
  OAI21_X2 U3806 ( .B1(n3263), .B2(n3793), .A(n3787), .ZN(n3315) );
  NAND2_X1 U3807 ( .A1(n3927), .A2(n3323), .ZN(n3802) );
  NAND2_X1 U3808 ( .A1(n3315), .A2(n3802), .ZN(n2978) );
  OR2_X1 U3809 ( .A1(n3323), .A2(n3927), .ZN(n3796) );
  NAND2_X1 U3810 ( .A1(n2978), .A2(n3796), .ZN(n3363) );
  NAND2_X1 U3811 ( .A1(n2979), .A2(n3926), .ZN(n3390) );
  NAND2_X1 U3812 ( .A1(n3394), .A2(n3925), .ZN(n2980) );
  NAND2_X1 U3813 ( .A1(n3390), .A2(n2980), .ZN(n2983) );
  INV_X1 U3814 ( .A(n3803), .ZN(n2981) );
  NOR2_X1 U3815 ( .A1(n2983), .A2(n2981), .ZN(n2982) );
  NAND2_X1 U3816 ( .A1(n3363), .A2(n2982), .ZN(n2986) );
  INV_X1 U3817 ( .A(n2983), .ZN(n3804) );
  NAND2_X1 U3818 ( .A1(n3627), .A2(n3714), .ZN(n3392) );
  NAND2_X1 U3819 ( .A1(n3392), .A2(n3361), .ZN(n2985) );
  NOR2_X1 U3820 ( .A1(n3394), .A2(n3925), .ZN(n2984) );
  AOI21_X1 U3821 ( .B1(n3804), .B2(n2985), .A(n2984), .ZN(n3812) );
  NAND2_X1 U3822 ( .A1(n2986), .A2(n3812), .ZN(n3379) );
  NAND2_X1 U3823 ( .A1(n3379), .A2(n2945), .ZN(n2987) );
  NAND2_X1 U3824 ( .A1(n2987), .A2(n3808), .ZN(n4270) );
  NAND2_X1 U3825 ( .A1(n2988), .A2(n3923), .ZN(n3798) );
  NAND2_X1 U3826 ( .A1(n4241), .A2(n4275), .ZN(n3809) );
  NAND2_X1 U3827 ( .A1(n3798), .A2(n3809), .ZN(n4269) );
  NAND2_X1 U3828 ( .A1(n4168), .A2(n4150), .ZN(n4110) );
  NAND2_X1 U3829 ( .A1(n4111), .A2(n4110), .ZN(n3820) );
  NAND2_X1 U3830 ( .A1(n4166), .A2(n4193), .ZN(n3847) );
  NAND2_X1 U3831 ( .A1(n3847), .A2(n4182), .ZN(n4161) );
  NAND2_X1 U3832 ( .A1(n4242), .A2(n4231), .ZN(n4201) );
  AND2_X1 U3833 ( .A1(n2989), .A2(n4201), .ZN(n4159) );
  NAND2_X1 U3834 ( .A1(n2990), .A2(n4165), .ZN(n2991) );
  OAI211_X1 U3835 ( .C1(n4161), .C2(n4159), .A(n4160), .B(n2991), .ZN(n4106)
         );
  OR2_X1 U3836 ( .A1(n3820), .A2(n4106), .ZN(n3887) );
  OR2_X1 U3837 ( .A1(n4161), .A2(n4105), .ZN(n3815) );
  INV_X1 U3838 ( .A(n4104), .ZN(n2992) );
  NOR2_X1 U3839 ( .A1(n3815), .A2(n2992), .ZN(n2997) );
  NAND2_X1 U3840 ( .A1(n4188), .A2(n4176), .ZN(n4108) );
  OR2_X1 U3841 ( .A1(n3820), .A2(n4108), .ZN(n2994) );
  AOI22_X1 U3842 ( .A1(n3921), .A2(n4120), .B1(n4149), .B2(n4139), .ZN(n2993)
         );
  AND2_X1 U3843 ( .A1(n2994), .A2(n2993), .ZN(n3819) );
  AND2_X1 U3844 ( .A1(n4129), .A2(n2995), .ZN(n3818) );
  NAND2_X1 U3845 ( .A1(n4111), .A2(n3818), .ZN(n2996) );
  OAI211_X1 U3846 ( .C1(n3887), .C2(n2997), .A(n3819), .B(n2996), .ZN(n3888)
         );
  INV_X1 U3847 ( .A(n3888), .ZN(n2998) );
  INV_X1 U3848 ( .A(n4098), .ZN(n3687) );
  NAND2_X1 U3849 ( .A1(n4115), .A2(n3687), .ZN(n3844) );
  INV_X1 U3850 ( .A(n3921), .ZN(n4131) );
  NAND2_X1 U3851 ( .A1(n4131), .A2(n3845), .ZN(n4087) );
  NAND2_X1 U3852 ( .A1(n4088), .A2(n3891), .ZN(n4070) );
  NAND2_X1 U3853 ( .A1(n4092), .A2(n4079), .ZN(n3843) );
  NAND2_X1 U3854 ( .A1(n3920), .A2(n4098), .ZN(n4069) );
  NAND2_X1 U3855 ( .A1(n4070), .A2(n3892), .ZN(n4051) );
  OR2_X1 U3856 ( .A1(n4075), .A2(n4061), .ZN(n3842) );
  NAND2_X1 U3857 ( .A1(n3745), .A2(n3016), .ZN(n4050) );
  AOI21_X1 U3858 ( .B1(n4051), .B2(n3895), .A(n3841), .ZN(n4030) );
  NAND2_X1 U3859 ( .A1(n4058), .A2(n3420), .ZN(n3828) );
  NAND2_X1 U3860 ( .A1(n3919), .A2(n4041), .ZN(n3825) );
  INV_X1 U3861 ( .A(n3828), .ZN(n2999) );
  XNOR2_X1 U3862 ( .A(n4017), .B(n4008), .ZN(n3006) );
  NAND2_X1 U3863 ( .A1(n4453), .A2(n4452), .ZN(n3001) );
  NAND2_X1 U3864 ( .A1(n3982), .A2(n4451), .ZN(n3000) );
  AOI22_X1 U3865 ( .A1(n3919), .A2(n4559), .B1(n4010), .B2(n4273), .ZN(n3004)
         );
  OAI21_X1 U3866 ( .B1(n3840), .B2(n4576), .A(n3004), .ZN(n3005) );
  AOI21_X1 U3867 ( .B1(n3006), .B2(n4573), .A(n3005), .ZN(n3433) );
  OAI21_X1 U3868 ( .B1(n3432), .B2(n4629), .A(n3433), .ZN(n3024) );
  INV_X1 U3869 ( .A(n4452), .ZN(n3007) );
  NAND2_X1 U3870 ( .A1(n4641), .A2(n3007), .ZN(n3008) );
  NAND2_X1 U3871 ( .A1(n3009), .A2(n3008), .ZN(n3013) );
  NAND2_X1 U3872 ( .A1(n3012), .A2(n3134), .ZN(n3119) );
  INV_X1 U3873 ( .A(n3014), .ZN(n3021) );
  INV_X1 U3874 ( .A(n4287), .ZN(n4293) );
  AND2_X2 U3875 ( .A1(n3324), .A2(n3323), .ZN(n3321) );
  NOR2_X4 U3876 ( .A1(n4367), .A2(n4275), .ZN(n4274) );
  INV_X1 U3877 ( .A(n4061), .ZN(n4055) );
  INV_X1 U3878 ( .A(n3017), .ZN(n3019) );
  OAI21_X1 U3879 ( .B1(n3019), .B2(n3018), .A(n4013), .ZN(n3436) );
  NAND2_X1 U3880 ( .A1(n3021), .A2(n2262), .ZN(U3546) );
  INV_X1 U3881 ( .A(n3022), .ZN(n3122) );
  INV_X1 U3882 ( .A(n3025), .ZN(n3026) );
  NAND2_X1 U3883 ( .A1(n3026), .A2(n2261), .ZN(U3514) );
  INV_X1 U3884 ( .A(n4591), .ZN(n3028) );
  OR2_X2 U3885 ( .A1(n3028), .A2(n3027), .ZN(n3929) );
  MUX2_X1 U3886 ( .A(n2881), .B(n2333), .S(U3149), .Z(n3029) );
  INV_X1 U3887 ( .A(n3029), .ZN(U3351) );
  INV_X1 U3888 ( .A(DATAI_5_), .ZN(n3031) );
  MUX2_X1 U3889 ( .A(n2846), .B(n3031), .S(U3149), .Z(n3032) );
  INV_X1 U3890 ( .A(n3032), .ZN(U3347) );
  INV_X1 U3891 ( .A(DATAI_31_), .ZN(n3036) );
  OR4_X1 U3892 ( .A1(n3034), .A2(IR_REG_30__SCAN_IN), .A3(n3033), .A4(U3149), 
        .ZN(n3035) );
  OAI21_X1 U3893 ( .B1(STATE_REG_SCAN_IN), .B2(n3036), .A(n3035), .ZN(U3321)
         );
  INV_X1 U3894 ( .A(DATAI_29_), .ZN(n3039) );
  NAND2_X1 U3895 ( .A1(n3037), .A2(STATE_REG_SCAN_IN), .ZN(n3038) );
  OAI21_X1 U3896 ( .B1(STATE_REG_SCAN_IN), .B2(n3039), .A(n3038), .ZN(U3323)
         );
  MUX2_X1 U3897 ( .A(n3207), .B(n2525), .S(U3149), .Z(n3040) );
  INV_X1 U3898 ( .A(n3040), .ZN(U3341) );
  INV_X1 U3899 ( .A(DATAI_19_), .ZN(n3041) );
  MUX2_X1 U3900 ( .A(n3041), .B(n3987), .S(STATE_REG_SCAN_IN), .Z(n3042) );
  INV_X1 U3901 ( .A(n3042), .ZN(U3333) );
  INV_X1 U3902 ( .A(n3043), .ZN(n3045) );
  AND2_X1 U3903 ( .A1(n4591), .A2(n3046), .ZN(n3048) );
  AOI22_X1 U3904 ( .A1(n4590), .A2(n2781), .B1(n3048), .B2(n3047), .ZN(U3458)
         );
  INV_X1 U3905 ( .A(D_REG_1__SCAN_IN), .ZN(n3503) );
  INV_X1 U3906 ( .A(n3049), .ZN(n3050) );
  AOI22_X1 U3907 ( .A1(n4590), .A2(n3503), .B1(n4591), .B2(n3050), .ZN(U3459)
         );
  NOR2_X1 U3908 ( .A1(n4535), .A2(U4043), .ZN(U3148) );
  INV_X1 U3909 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n3517) );
  NAND2_X1 U3910 ( .A1(U4043), .A2(n3631), .ZN(n3051) );
  OAI21_X1 U3911 ( .B1(U4043), .B2(n3517), .A(n3051), .ZN(U3561) );
  INV_X1 U3912 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n3552) );
  INV_X1 U3913 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3505) );
  NAND2_X1 U3914 ( .A1(n2447), .A2(REG2_REG_31__SCAN_IN), .ZN(n3053) );
  INV_X1 U3915 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4390) );
  OR2_X1 U3916 ( .A1(n2764), .A2(n4390), .ZN(n3052) );
  OAI211_X1 U3917 ( .C1(n3831), .C2(n3505), .A(n3053), .B(n3052), .ZN(n3995)
         );
  NAND2_X1 U3918 ( .A1(U4043), .A2(n3995), .ZN(n3054) );
  OAI21_X1 U3919 ( .B1(U4043), .B2(n3552), .A(n3054), .ZN(U3581) );
  INV_X1 U3920 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n3545) );
  NAND2_X1 U3921 ( .A1(U4043), .A2(n2969), .ZN(n3055) );
  OAI21_X1 U3922 ( .B1(U4043), .B2(n3545), .A(n3055), .ZN(U3550) );
  XOR2_X1 U3923 ( .A(n3056), .B(REG1_REG_3__SCAN_IN), .Z(n3059) );
  XNOR2_X1 U3924 ( .A(n3057), .B(n3308), .ZN(n3058) );
  AOI22_X1 U3925 ( .A1(n4545), .A2(n3059), .B1(n4543), .B2(n3058), .ZN(n3061)
         );
  INV_X1 U3926 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3513) );
  NOR2_X1 U3927 ( .A1(STATE_REG_SCAN_IN), .A2(n3513), .ZN(n3145) );
  AOI21_X1 U3928 ( .B1(n4535), .B2(ADDR_REG_3__SCAN_IN), .A(n3145), .ZN(n3060)
         );
  OAI211_X1 U3929 ( .C1(n3062), .C2(n4548), .A(n3061), .B(n3060), .ZN(U3243)
         );
  XNOR2_X1 U3930 ( .A(n3063), .B(REG1_REG_6__SCAN_IN), .ZN(n3069) );
  INV_X1 U3931 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3341) );
  XNOR2_X1 U3932 ( .A(n3064), .B(n3341), .ZN(n3067) );
  AND2_X1 U3933 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3152) );
  AOI21_X1 U3934 ( .B1(n4535), .B2(ADDR_REG_6__SCAN_IN), .A(n3152), .ZN(n3065)
         );
  OAI21_X1 U3935 ( .B1(n4548), .B2(n2169), .A(n3065), .ZN(n3066) );
  AOI21_X1 U3936 ( .B1(n3067), .B2(n4543), .A(n3066), .ZN(n3068) );
  OAI21_X1 U3937 ( .B1(n3069), .B2(n4513), .A(n3068), .ZN(U3246) );
  INV_X1 U3938 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n3523) );
  NAND2_X1 U3939 ( .A1(n4205), .A2(U4043), .ZN(n3070) );
  OAI21_X1 U3940 ( .B1(U4043), .B2(n3523), .A(n3070), .ZN(U3567) );
  MUX2_X1 U3941 ( .A(REG1_REG_7__SCAN_IN), .B(n2849), .S(n3076), .Z(n3071) );
  XNOR2_X1 U3942 ( .A(n3072), .B(n3071), .ZN(n3081) );
  INV_X1 U3943 ( .A(n4543), .ZN(n4504) );
  AOI21_X1 U3944 ( .B1(n3074), .B2(n3073), .A(n4504), .ZN(n3079) );
  AND2_X1 U3945 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3166) );
  AOI21_X1 U3946 ( .B1(n4535), .B2(ADDR_REG_7__SCAN_IN), .A(n3166), .ZN(n3075)
         );
  OAI21_X1 U3947 ( .B1(n4548), .B2(n3076), .A(n3075), .ZN(n3077) );
  AOI21_X1 U3948 ( .B1(n3079), .B2(n3078), .A(n3077), .ZN(n3080) );
  OAI21_X1 U3949 ( .B1(n4513), .B2(n3081), .A(n3080), .ZN(U3247) );
  AOI211_X1 U3950 ( .C1(n3083), .C2(n3082), .A(n2047), .B(n4504), .ZN(n3090)
         );
  AOI211_X1 U3951 ( .C1(n3086), .C2(n3085), .A(n3084), .B(n4513), .ZN(n3089)
         );
  AND2_X1 U3952 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3664) );
  AOI21_X1 U3953 ( .B1(n4535), .B2(ADDR_REG_5__SCAN_IN), .A(n3664), .ZN(n3087)
         );
  OAI21_X1 U3954 ( .B1(n4548), .B2(n2846), .A(n3087), .ZN(n3088) );
  OR3_X1 U3955 ( .A1(n3090), .A2(n3089), .A3(n3088), .ZN(U3245) );
  XNOR2_X1 U3956 ( .A(n3091), .B(n3257), .ZN(n3098) );
  NOR2_X1 U3957 ( .A1(STATE_REG_SCAN_IN), .A2(n3092), .ZN(n3176) );
  NOR2_X1 U3958 ( .A1(n4548), .A2(n4456), .ZN(n3093) );
  AOI211_X1 U3959 ( .C1(n4535), .C2(ADDR_REG_8__SCAN_IN), .A(n3176), .B(n3093), 
        .ZN(n3097) );
  OAI211_X1 U3960 ( .C1(n3095), .C2(REG1_REG_8__SCAN_IN), .A(n3094), .B(n4545), 
        .ZN(n3096) );
  OAI211_X1 U3961 ( .C1(n3098), .C2(n4504), .A(n3097), .B(n3096), .ZN(U3248)
         );
  XNOR2_X1 U3962 ( .A(n3100), .B(n3099), .ZN(n3108) );
  AND2_X1 U3963 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3233) );
  NOR2_X1 U3964 ( .A1(n4548), .A2(n3101), .ZN(n3102) );
  AOI211_X1 U3965 ( .C1(n4535), .C2(ADDR_REG_9__SCAN_IN), .A(n3233), .B(n3102), 
        .ZN(n3107) );
  OAI211_X1 U3966 ( .C1(n3105), .C2(n3104), .A(n3103), .B(n4545), .ZN(n3106)
         );
  OAI211_X1 U3967 ( .C1(n3108), .C2(n4504), .A(n3107), .B(n3106), .ZN(U3249)
         );
  XNOR2_X1 U3968 ( .A(n3109), .B(n3110), .ZN(n3125) );
  XOR2_X1 U3969 ( .A(n3110), .B(n3111), .Z(n3114) );
  AOI22_X1 U3970 ( .A1(n4559), .A2(n2925), .B1(n3933), .B2(n4557), .ZN(n3112)
         );
  OAI21_X1 U3971 ( .B1(n4563), .B2(n3117), .A(n3112), .ZN(n3113) );
  AOI21_X1 U3972 ( .B1(n3114), .B2(n4573), .A(n3113), .ZN(n3115) );
  OAI21_X1 U3973 ( .B1(n4172), .B2(n3125), .A(n3115), .ZN(n4625) );
  INV_X1 U3974 ( .A(n3116), .ZN(n3118) );
  OAI211_X1 U3975 ( .C1(n3118), .C2(n3117), .A(n3020), .B(n3226), .ZN(n4624)
         );
  OAI22_X1 U3976 ( .A1(n4624), .A2(n3982), .B1(n4276), .B2(n3415), .ZN(n3124)
         );
  INV_X1 U3977 ( .A(n3119), .ZN(n3121) );
  NAND3_X1 U3978 ( .A1(n3122), .A2(n3121), .A3(n3120), .ZN(n3123) );
  OAI21_X1 U3979 ( .B1(n4625), .B2(n3124), .A(n4581), .ZN(n3129) );
  INV_X1 U3980 ( .A(n3125), .ZN(n4627) );
  OR2_X1 U3981 ( .A1(n3126), .A2(n3987), .ZN(n3198) );
  INV_X1 U3982 ( .A(n3198), .ZN(n3127) );
  AOI22_X1 U3983 ( .A1(n4627), .A2(n4579), .B1(REG2_REG_4__SCAN_IN), .B2(n1998), .ZN(n3128) );
  NAND2_X1 U3984 ( .A1(n3129), .A2(n3128), .ZN(U3286) );
  XNOR2_X1 U3985 ( .A(n3131), .B(n3130), .ZN(n3944) );
  OAI22_X1 U3986 ( .A1(n3702), .A2(n3767), .B1(n3750), .B2(n3944), .ZN(n3139)
         );
  OAI21_X1 U3987 ( .B1(n3914), .B2(n3133), .A(n3132), .ZN(n3135) );
  NAND2_X1 U3988 ( .A1(n3135), .A2(n3134), .ZN(n3467) );
  INV_X1 U3989 ( .A(n3467), .ZN(n3137) );
  INV_X1 U3990 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3136) );
  OAI22_X1 U3991 ( .A1(n3701), .A2(n2920), .B1(n3137), .B2(n3136), .ZN(n3138)
         );
  OR2_X1 U3992 ( .A1(n3139), .A2(n3138), .ZN(U3229) );
  NAND2_X1 U3993 ( .A1(n3140), .A2(n3141), .ZN(n3142) );
  XOR2_X1 U3994 ( .A(n3143), .B(n3142), .Z(n3148) );
  NOR2_X1 U3995 ( .A1(n3762), .A2(REG3_REG_3__SCAN_IN), .ZN(n3144) );
  AOI211_X1 U3996 ( .C1(n3757), .C2(n4558), .A(n3145), .B(n3144), .ZN(n3147)
         );
  AOI22_X1 U3997 ( .A1(n3774), .A2(n3724), .B1(n3759), .B2(n3934), .ZN(n3146)
         );
  OAI211_X1 U3998 ( .C1(n3148), .C2(n3750), .A(n3147), .B(n3146), .ZN(U3215)
         );
  INV_X1 U3999 ( .A(n3157), .ZN(n3159) );
  XNOR2_X1 U4000 ( .A(n3156), .B(n3159), .ZN(n3150) );
  XNOR2_X1 U4001 ( .A(n3149), .B(n3150), .ZN(n3155) );
  AOI22_X1 U4002 ( .A1(n3336), .A2(n3724), .B1(n3759), .B2(n3931), .ZN(n3154)
         );
  NOR2_X1 U4003 ( .A1(n3762), .A2(n3340), .ZN(n3151) );
  AOI211_X1 U4004 ( .C1(n3757), .C2(n3933), .A(n3152), .B(n3151), .ZN(n3153)
         );
  OAI211_X1 U4005 ( .C1(n3155), .C2(n3750), .A(n3154), .B(n3153), .ZN(U3236)
         );
  INV_X1 U4006 ( .A(n3149), .ZN(n3160) );
  OAI21_X1 U4007 ( .B1(n3149), .B2(n3157), .A(n3156), .ZN(n3158) );
  OAI21_X1 U4008 ( .B1(n3160), .B2(n3159), .A(n3158), .ZN(n3164) );
  XOR2_X1 U4009 ( .A(n3162), .B(n3161), .Z(n3163) );
  XNOR2_X1 U4010 ( .A(n3164), .B(n3163), .ZN(n3169) );
  AOI22_X1 U4011 ( .A1(n3188), .A2(n3724), .B1(n3759), .B2(n3930), .ZN(n3168)
         );
  NOR2_X1 U4012 ( .A1(n3762), .A2(n3189), .ZN(n3165) );
  AOI211_X1 U4013 ( .C1(n3757), .C2(n3932), .A(n3166), .B(n3165), .ZN(n3167)
         );
  OAI211_X1 U4014 ( .C1(n3169), .C2(n3750), .A(n3168), .B(n3167), .ZN(U3210)
         );
  INV_X1 U4015 ( .A(n3171), .ZN(n3173) );
  NOR2_X1 U4016 ( .A1(n3173), .A2(n3172), .ZN(n3174) );
  XNOR2_X1 U4017 ( .A(n3170), .B(n3174), .ZN(n3179) );
  AOI22_X1 U4018 ( .A1(n3254), .A2(n3724), .B1(n3757), .B2(n3931), .ZN(n3178)
         );
  NOR2_X1 U4019 ( .A1(n3762), .A2(n3256), .ZN(n3175) );
  AOI211_X1 U4020 ( .C1(n3759), .C2(n3928), .A(n3176), .B(n3175), .ZN(n3177)
         );
  OAI211_X1 U4021 ( .C1(n3179), .C2(n3750), .A(n3178), .B(n3177), .ZN(U3218)
         );
  INV_X1 U4022 ( .A(n3180), .ZN(n3864) );
  XNOR2_X1 U4023 ( .A(n3181), .B(n3864), .ZN(n3182) );
  NAND2_X1 U4024 ( .A1(n3182), .A2(n4573), .ZN(n3184) );
  AOI22_X1 U4025 ( .A1(n3930), .A2(n4557), .B1(n4559), .B2(n3932), .ZN(n3183)
         );
  OAI211_X1 U4026 ( .C1(n4563), .C2(n3185), .A(n3184), .B(n3183), .ZN(n4642)
         );
  INV_X1 U4027 ( .A(n4642), .ZN(n3202) );
  INV_X1 U4028 ( .A(n4636), .ZN(n3187) );
  INV_X1 U4029 ( .A(n3255), .ZN(n3186) );
  AOI211_X1 U4030 ( .C1(n3188), .C2(n3187), .A(n4635), .B(n3186), .ZN(n4643)
         );
  OAI22_X1 U4031 ( .A1(n4581), .A2(n3570), .B1(n3189), .B2(n4276), .ZN(n3190)
         );
  AOI21_X1 U4032 ( .B1(n4643), .B2(n4215), .A(n3190), .ZN(n3201) );
  NAND2_X1 U4033 ( .A1(n3109), .A2(n3191), .ZN(n3193) );
  AND2_X1 U4034 ( .A1(n3193), .A2(n3192), .ZN(n3332) );
  INV_X1 U4035 ( .A(n3332), .ZN(n3194) );
  OAI21_X1 U4036 ( .B1(n3194), .B2(n3932), .A(n3336), .ZN(n3195) );
  OAI21_X1 U4037 ( .B1(n3196), .B2(n3332), .A(n3195), .ZN(n3197) );
  XNOR2_X1 U4038 ( .A(n3197), .B(n3864), .ZN(n4645) );
  NAND2_X1 U4039 ( .A1(n4172), .A2(n3198), .ZN(n3199) );
  NAND2_X1 U4040 ( .A1(n4645), .A2(n4258), .ZN(n3200) );
  OAI211_X1 U4041 ( .C1(n3202), .C2(n1998), .A(n3201), .B(n3200), .ZN(U3283)
         );
  XOR2_X1 U4042 ( .A(n3204), .B(n3203), .Z(n3213) );
  NOR2_X1 U40430 ( .A1(n3205), .A2(STATE_REG_SCAN_IN), .ZN(n3279) );
  AOI21_X1 U4044 ( .B1(n4535), .B2(ADDR_REG_11__SCAN_IN), .A(n3279), .ZN(n3206) );
  OAI21_X1 U4045 ( .B1(n4548), .B2(n3207), .A(n3206), .ZN(n3212) );
  AOI211_X1 U4046 ( .C1(n3210), .C2(n3209), .A(n4513), .B(n3208), .ZN(n3211)
         );
  AOI211_X1 U4047 ( .C1(n4543), .C2(n3213), .A(n3212), .B(n3211), .ZN(n3214)
         );
  INV_X1 U4048 ( .A(n3214), .ZN(U3251) );
  NAND2_X1 U4049 ( .A1(n3109), .A2(n3110), .ZN(n3216) );
  NAND2_X1 U4050 ( .A1(n3216), .A2(n3215), .ZN(n3218) );
  INV_X1 U4051 ( .A(n3217), .ZN(n3778) );
  NAND2_X1 U4052 ( .A1(n3778), .A2(n3792), .ZN(n3856) );
  XNOR2_X1 U4053 ( .A(n3218), .B(n3856), .ZN(n4630) );
  XNOR2_X1 U4054 ( .A(n3219), .B(n3856), .ZN(n3223) );
  AOI22_X1 U4055 ( .A1(n4557), .A2(n3932), .B1(n3934), .B2(n4559), .ZN(n3220)
         );
  OAI21_X1 U4056 ( .B1(n4563), .B2(n3221), .A(n3220), .ZN(n3222) );
  AOI21_X1 U4057 ( .B1(n3223), .B2(n4573), .A(n3222), .ZN(n4631) );
  MUX2_X1 U4058 ( .A(n4631), .B(n3224), .S(n1998), .Z(n3229) );
  AOI21_X1 U4059 ( .B1(n3661), .B2(n3226), .A(n3225), .ZN(n4634) );
  INV_X1 U4060 ( .A(n3662), .ZN(n3227) );
  AOI22_X1 U4061 ( .A1(n4567), .A2(n4634), .B1(n3227), .B2(n4578), .ZN(n3228)
         );
  OAI211_X1 U4062 ( .C1(n4283), .C2(n4630), .A(n3229), .B(n3228), .ZN(U3285)
         );
  NAND2_X1 U4063 ( .A1(n3929), .A2(DATAO_REG_29__SCAN_IN), .ZN(n3230) );
  OAI21_X1 U4064 ( .B1(n3840), .B2(n3929), .A(n3230), .ZN(U3579) );
  OAI21_X1 U4065 ( .B1(n3232), .B2(n3231), .A(n3242), .ZN(n3237) );
  AOI22_X1 U4066 ( .A1(n3267), .A2(n3758), .B1(n3759), .B2(n3927), .ZN(n3235)
         );
  AOI21_X1 U4067 ( .B1(n3757), .B2(n3930), .A(n3233), .ZN(n3234) );
  OAI211_X1 U4068 ( .C1(n3762), .C2(n3268), .A(n3235), .B(n3234), .ZN(n3236)
         );
  AOI21_X1 U4069 ( .B1(n3237), .B2(n3764), .A(n3236), .ZN(n3238) );
  INV_X1 U4070 ( .A(n3238), .ZN(U3228) );
  NAND2_X1 U4071 ( .A1(n3239), .A2(n3764), .ZN(n3247) );
  AOI21_X1 U4072 ( .B1(n3242), .B2(n3241), .A(n3240), .ZN(n3246) );
  AOI22_X1 U4073 ( .A1(n3318), .A2(n3724), .B1(n3757), .B2(n3928), .ZN(n3245)
         );
  NOR2_X1 U4074 ( .A1(STATE_REG_SCAN_IN), .A2(n2100), .ZN(n4485) );
  NOR2_X1 U4075 ( .A1(n3762), .A2(n3325), .ZN(n3243) );
  AOI211_X1 U4076 ( .C1(n3759), .C2(n3631), .A(n4485), .B(n3243), .ZN(n3244)
         );
  OAI211_X1 U4077 ( .C1(n3247), .C2(n3246), .A(n3245), .B(n3244), .ZN(U3214)
         );
  NAND2_X1 U4078 ( .A1(n3786), .A2(n3784), .ZN(n3857) );
  XNOR2_X1 U4079 ( .A(n3248), .B(n3857), .ZN(n3253) );
  XNOR2_X1 U4080 ( .A(n3249), .B(n3857), .ZN(n4389) );
  OAI22_X1 U4081 ( .A1(n3334), .A2(n4264), .B1(n3316), .B2(n4576), .ZN(n3250)
         );
  AOI21_X1 U4082 ( .B1(n3254), .B2(n4273), .A(n3250), .ZN(n3251) );
  OAI21_X1 U4083 ( .B1(n4389), .B2(n4172), .A(n3251), .ZN(n3252) );
  AOI21_X1 U4084 ( .B1(n4573), .B2(n3253), .A(n3252), .ZN(n4387) );
  INV_X1 U4085 ( .A(n4389), .ZN(n3260) );
  NAND2_X1 U4086 ( .A1(n3255), .A2(n3254), .ZN(n4384) );
  AND3_X1 U4087 ( .A1(n4567), .A2(n4385), .A3(n4384), .ZN(n3259) );
  OAI22_X1 U4088 ( .A1(n4581), .A2(n3257), .B1(n3256), .B2(n4276), .ZN(n3258)
         );
  AOI211_X1 U4089 ( .C1(n3260), .C2(n4579), .A(n3259), .B(n3258), .ZN(n3261)
         );
  OAI21_X1 U4090 ( .B1(n4387), .B2(n1998), .A(n3261), .ZN(U3282) );
  OAI22_X1 U4091 ( .A1(n3262), .A2(n4264), .B1(n3285), .B2(n4576), .ZN(n3266)
         );
  INV_X1 U4092 ( .A(n3793), .ZN(n3789) );
  AND2_X1 U4093 ( .A1(n3789), .A2(n3787), .ZN(n3852) );
  XNOR2_X1 U4094 ( .A(n3263), .B(n3852), .ZN(n3264) );
  NOR2_X1 U4095 ( .A1(n3264), .A2(n4288), .ZN(n3265) );
  AOI211_X1 U4096 ( .C1(n4273), .C2(n3267), .A(n3266), .B(n3265), .ZN(n3354)
         );
  AOI21_X1 U4097 ( .B1(n3267), .B2(n4385), .A(n3324), .ZN(n3358) );
  OAI22_X1 U4098 ( .A1(n4581), .A2(n3581), .B1(n3268), .B2(n4276), .ZN(n3269)
         );
  AOI21_X1 U4099 ( .B1(n3358), .B2(n4567), .A(n3269), .ZN(n3272) );
  XOR2_X1 U4100 ( .A(n3270), .B(n3852), .Z(n3356) );
  NAND2_X1 U4101 ( .A1(n3356), .A2(n4258), .ZN(n3271) );
  OAI211_X1 U4102 ( .C1(n3354), .C2(n1998), .A(n3272), .B(n3271), .ZN(U3281)
         );
  INV_X1 U4103 ( .A(n3273), .ZN(n3275) );
  NOR2_X1 U4104 ( .A1(n3275), .A2(n3274), .ZN(n3276) );
  XNOR2_X1 U4105 ( .A(n3277), .B(n3276), .ZN(n3282) );
  AOI22_X1 U4106 ( .A1(n3287), .A2(n3724), .B1(n3757), .B2(n3927), .ZN(n3281)
         );
  NOR2_X1 U4107 ( .A1(n3762), .A2(n3293), .ZN(n3278) );
  AOI211_X1 U4108 ( .C1(n3759), .C2(n3926), .A(n3279), .B(n3278), .ZN(n3280)
         );
  OAI211_X1 U4109 ( .C1(n3282), .C2(n3750), .A(n3281), .B(n3280), .ZN(U3233)
         );
  INV_X1 U4110 ( .A(n3283), .ZN(n3851) );
  XNOR2_X1 U4111 ( .A(n3363), .B(n3851), .ZN(n3290) );
  XNOR2_X1 U4112 ( .A(n3284), .B(n3851), .ZN(n3291) );
  OAI22_X1 U4113 ( .A1(n3714), .A2(n4576), .B1(n3285), .B2(n4264), .ZN(n3286)
         );
  AOI21_X1 U4114 ( .B1(n3287), .B2(n4273), .A(n3286), .ZN(n3288) );
  OAI21_X1 U4115 ( .B1(n3291), .B2(n4172), .A(n3288), .ZN(n3289) );
  AOI21_X1 U4116 ( .B1(n3290), .B2(n4573), .A(n3289), .ZN(n4382) );
  INV_X1 U4117 ( .A(n3291), .ZN(n4380) );
  OAI21_X1 U4118 ( .B1(n3321), .B2(n3292), .A(n3369), .ZN(n4383) );
  NOR2_X1 U4119 ( .A1(n4383), .A2(n4234), .ZN(n3295) );
  OAI22_X1 U4120 ( .A1(n4581), .A2(n3554), .B1(n3293), .B2(n4276), .ZN(n3294)
         );
  AOI211_X1 U4121 ( .C1(n4380), .C2(n4579), .A(n3295), .B(n3294), .ZN(n3296)
         );
  OAI21_X1 U4122 ( .B1(n4382), .B2(n1998), .A(n3296), .ZN(U3279) );
  INV_X1 U4123 ( .A(n3860), .ZN(n3299) );
  XNOR2_X1 U4124 ( .A(n3297), .B(n3299), .ZN(n4620) );
  INV_X1 U4125 ( .A(n4172), .ZN(n4574) );
  NAND2_X1 U4126 ( .A1(n4620), .A2(n4574), .ZN(n3307) );
  NAND3_X1 U4127 ( .A1(n3298), .A2(n3770), .A3(n3299), .ZN(n3300) );
  NAND2_X1 U4128 ( .A1(n3301), .A2(n3300), .ZN(n3305) );
  AOI22_X1 U4129 ( .A1(n4559), .A2(n4558), .B1(n3934), .B2(n4557), .ZN(n3303)
         );
  NAND2_X1 U4130 ( .A1(n4273), .A2(n3774), .ZN(n3302) );
  NAND2_X1 U4131 ( .A1(n3303), .A2(n3302), .ZN(n3304) );
  AOI21_X1 U4132 ( .B1(n3305), .B2(n4573), .A(n3304), .ZN(n3306) );
  AND2_X1 U4133 ( .A1(n3307), .A2(n3306), .ZN(n4622) );
  OAI22_X1 U4134 ( .A1(n4581), .A2(n3308), .B1(n4276), .B2(REG3_REG_3__SCAN_IN), .ZN(n3313) );
  OR2_X1 U4135 ( .A1(n3309), .A2(n3310), .ZN(n3311) );
  NAND2_X1 U4136 ( .A1(n3116), .A2(n3311), .ZN(n4618) );
  NOR2_X1 U4137 ( .A1(n4234), .A2(n4618), .ZN(n3312) );
  AOI211_X1 U4138 ( .C1(n4579), .C2(n4620), .A(n3313), .B(n3312), .ZN(n3314)
         );
  OAI21_X1 U4139 ( .B1(n1998), .B2(n4622), .A(n3314), .ZN(U3287) );
  NAND2_X1 U4140 ( .A1(n3796), .A2(n3802), .ZN(n3855) );
  XNOR2_X1 U4141 ( .A(n3315), .B(n3855), .ZN(n3320) );
  OAI22_X1 U4142 ( .A1(n3316), .A2(n4264), .B1(n3364), .B2(n4576), .ZN(n3317)
         );
  AOI21_X1 U4143 ( .B1(n3318), .B2(n4273), .A(n3317), .ZN(n3319) );
  OAI21_X1 U4144 ( .B1(n3320), .B2(n4288), .A(n3319), .ZN(n3347) );
  INV_X1 U4145 ( .A(n3347), .ZN(n3330) );
  XNOR2_X1 U4146 ( .A(n2007), .B(n3855), .ZN(n3348) );
  INV_X1 U4147 ( .A(n3321), .ZN(n3322) );
  OAI21_X1 U4148 ( .B1(n3324), .B2(n3323), .A(n3322), .ZN(n3353) );
  NOR2_X1 U4149 ( .A1(n3353), .A2(n4234), .ZN(n3328) );
  OAI22_X1 U4150 ( .A1(n4581), .A2(n3326), .B1(n3325), .B2(n4276), .ZN(n3327)
         );
  AOI211_X1 U4151 ( .C1(n3348), .C2(n4258), .A(n3328), .B(n3327), .ZN(n3329)
         );
  OAI21_X1 U4152 ( .B1(n1998), .B2(n3330), .A(n3329), .ZN(U3280) );
  NAND2_X1 U4153 ( .A1(n3781), .A2(n3791), .ZN(n3858) );
  XNOR2_X1 U4154 ( .A(n3331), .B(n3858), .ZN(n3339) );
  XNOR2_X1 U4155 ( .A(n3332), .B(n3858), .ZN(n4640) );
  NAND2_X1 U4156 ( .A1(n4640), .A2(n4574), .ZN(n3338) );
  OAI22_X1 U4157 ( .A1(n3334), .A2(n4576), .B1(n3333), .B2(n4264), .ZN(n3335)
         );
  AOI21_X1 U4158 ( .B1(n3336), .B2(n4273), .A(n3335), .ZN(n3337) );
  OAI211_X1 U4159 ( .C1(n3339), .C2(n4288), .A(n3338), .B(n3337), .ZN(n4638)
         );
  INV_X1 U4160 ( .A(n4638), .ZN(n3346) );
  OAI22_X1 U4161 ( .A1(n4581), .A2(n3341), .B1(n3340), .B2(n4276), .ZN(n3344)
         );
  NOR2_X1 U4162 ( .A1(n3225), .A2(n3342), .ZN(n4637) );
  NOR3_X1 U4163 ( .A1(n4234), .A2(n4636), .A3(n4637), .ZN(n3343) );
  AOI211_X1 U4164 ( .C1(n4579), .C2(n4640), .A(n3344), .B(n3343), .ZN(n3345)
         );
  OAI21_X1 U4165 ( .B1(n1998), .B2(n3346), .A(n3345), .ZN(U3284) );
  INV_X1 U4166 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3349) );
  AOI21_X1 U4167 ( .B1(n3348), .B2(n4644), .A(n3347), .ZN(n3351) );
  MUX2_X1 U4168 ( .A(n3349), .B(n3351), .S(n4647), .Z(n3350) );
  OAI21_X1 U4169 ( .B1(n3353), .B2(n4444), .A(n3350), .ZN(U3487) );
  MUX2_X1 U4170 ( .A(n4484), .B(n3351), .S(n4658), .Z(n3352) );
  OAI21_X1 U4171 ( .B1(n4379), .B2(n3353), .A(n3352), .ZN(U3528) );
  INV_X1 U4172 ( .A(n3354), .ZN(n3355) );
  AOI21_X1 U4173 ( .B1(n4644), .B2(n3356), .A(n3355), .ZN(n3360) );
  INV_X1 U4174 ( .A(n4444), .ZN(n4395) );
  AOI22_X1 U4175 ( .A1(n3358), .A2(n4395), .B1(REG0_REG_9__SCAN_IN), .B2(n4646), .ZN(n3357) );
  OAI21_X1 U4176 ( .B1(n3360), .B2(n4646), .A(n3357), .ZN(U3485) );
  INV_X1 U4177 ( .A(n4379), .ZN(n4299) );
  AOI22_X1 U4178 ( .A1(n3358), .A2(n4299), .B1(REG1_REG_9__SCAN_IN), .B2(n4656), .ZN(n3359) );
  OAI21_X1 U4179 ( .B1(n3360), .B2(n4656), .A(n3359), .ZN(U3527) );
  NAND2_X1 U4180 ( .A1(n3390), .A2(n3392), .ZN(n3848) );
  INV_X1 U4181 ( .A(n3361), .ZN(n3362) );
  AOI21_X1 U4182 ( .B1(n3363), .B2(n3803), .A(n3362), .ZN(n3393) );
  XOR2_X1 U4183 ( .A(n3848), .B(n3393), .Z(n3367) );
  OAI22_X1 U4184 ( .A1(n3380), .A2(n4576), .B1(n3364), .B2(n4264), .ZN(n3365)
         );
  AOI21_X1 U4185 ( .B1(n3627), .B2(n4273), .A(n3365), .ZN(n3366) );
  OAI21_X1 U4186 ( .B1(n3367), .B2(n4288), .A(n3366), .ZN(n4376) );
  INV_X1 U4187 ( .A(n4376), .ZN(n3375) );
  XOR2_X1 U4188 ( .A(n3368), .B(n3848), .Z(n4377) );
  NAND2_X1 U4189 ( .A1(n3369), .A2(n3627), .ZN(n3370) );
  NAND2_X1 U4190 ( .A1(n3402), .A2(n3370), .ZN(n4445) );
  NOR2_X1 U4191 ( .A1(n4445), .A2(n4234), .ZN(n3373) );
  INV_X1 U4192 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3371) );
  OAI22_X1 U4193 ( .A1(n4581), .A2(n3371), .B1(n3629), .B2(n4276), .ZN(n3372)
         );
  AOI211_X1 U4194 ( .C1(n4377), .C2(n4258), .A(n3373), .B(n3372), .ZN(n3374)
         );
  OAI21_X1 U4195 ( .B1(n1998), .B2(n3375), .A(n3374), .ZN(U3278) );
  INV_X1 U4196 ( .A(n3376), .ZN(n3378) );
  NAND2_X1 U4197 ( .A1(n3376), .A2(n3870), .ZN(n4262) );
  INV_X1 U4198 ( .A(n4262), .ZN(n3377) );
  AOI21_X1 U4199 ( .B1(n2945), .B2(n3378), .A(n3377), .ZN(n4371) );
  INV_X1 U4200 ( .A(n4371), .ZN(n3388) );
  XNOR2_X1 U4201 ( .A(n3379), .B(n3870), .ZN(n3383) );
  OAI22_X1 U4202 ( .A1(n4241), .A2(n4576), .B1(n3380), .B2(n4264), .ZN(n3381)
         );
  AOI21_X1 U4203 ( .B1(n3444), .B2(n4273), .A(n3381), .ZN(n3382) );
  OAI21_X1 U4204 ( .B1(n3383), .B2(n4288), .A(n3382), .ZN(n3384) );
  AOI21_X1 U4205 ( .B1(n3388), .B2(n4574), .A(n3384), .ZN(n4370) );
  OAI21_X1 U4206 ( .B1(n3402), .B2(n3712), .A(n3444), .ZN(n4368) );
  AND3_X1 U4207 ( .A1(n4368), .A2(n4567), .A3(n4367), .ZN(n3387) );
  OAI22_X1 U4208 ( .A1(n4581), .A2(n3385), .B1(n3446), .B2(n4276), .ZN(n3386)
         );
  AOI211_X1 U4209 ( .C1(n3388), .C2(n4579), .A(n3387), .B(n3386), .ZN(n3389)
         );
  OAI21_X1 U4210 ( .B1(n1998), .B2(n4370), .A(n3389), .ZN(U3276) );
  INV_X1 U4211 ( .A(n3390), .ZN(n3391) );
  AOI21_X1 U4212 ( .B1(n3393), .B2(n3392), .A(n3391), .ZN(n3395) );
  XNOR2_X1 U4213 ( .A(n3394), .B(n3925), .ZN(n3869) );
  XNOR2_X1 U4214 ( .A(n3395), .B(n3869), .ZN(n3400) );
  OAI22_X1 U4215 ( .A1(n4265), .A2(n4576), .B1(n3714), .B2(n4264), .ZN(n3398)
         );
  XNOR2_X1 U4216 ( .A(n3396), .B(n3869), .ZN(n3401) );
  NOR2_X1 U4217 ( .A1(n3401), .A2(n4172), .ZN(n3397) );
  AOI211_X1 U4218 ( .C1(n4273), .C2(n3712), .A(n3398), .B(n3397), .ZN(n3399)
         );
  OAI21_X1 U4219 ( .B1(n4288), .B2(n3400), .A(n3399), .ZN(n4372) );
  INV_X1 U4220 ( .A(n4372), .ZN(n3406) );
  INV_X1 U4221 ( .A(n3401), .ZN(n4373) );
  XNOR2_X1 U4222 ( .A(n3402), .B(n3712), .ZN(n4440) );
  AOI22_X1 U4223 ( .A1(n1998), .A2(REG2_REG_13__SCAN_IN), .B1(n3716), .B2(
        n4578), .ZN(n3403) );
  OAI21_X1 U4224 ( .B1(n4440), .B2(n4234), .A(n3403), .ZN(n3404) );
  AOI21_X1 U4225 ( .B1(n4373), .B2(n4579), .A(n3404), .ZN(n3405) );
  OAI21_X1 U4226 ( .B1(n3406), .B2(n1998), .A(n3405), .ZN(U3277) );
  INV_X1 U4227 ( .A(n3407), .ZN(n3410) );
  INV_X1 U4228 ( .A(n3408), .ZN(n3409) );
  AOI211_X1 U4229 ( .C1(n3411), .C2(n3410), .A(n3750), .B(n3409), .ZN(n3417)
         );
  AOI22_X1 U4230 ( .A1(n3412), .A2(n3758), .B1(n3759), .B2(n3933), .ZN(n3414)
         );
  AND2_X1 U4231 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4475) );
  AOI21_X1 U4232 ( .B1(n3757), .B2(n2925), .A(n4475), .ZN(n3413) );
  OAI211_X1 U4233 ( .C1(n3762), .C2(n3415), .A(n3414), .B(n3413), .ZN(n3416)
         );
  OR2_X1 U4234 ( .A1(n3417), .A2(n3416), .ZN(U3227) );
  XNOR2_X1 U4235 ( .A(n3419), .B(n3418), .ZN(n3425) );
  AOI22_X1 U4236 ( .A1(n4075), .A2(n3757), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3422) );
  NAND2_X1 U4237 ( .A1(n3758), .A2(n3420), .ZN(n3421) );
  OAI211_X1 U4238 ( .C1(n3762), .C2(n4044), .A(n3422), .B(n3421), .ZN(n3423)
         );
  AOI21_X1 U4239 ( .B1(n3759), .B2(n4022), .A(n3423), .ZN(n3424) );
  OAI21_X1 U4240 ( .B1(n3425), .B2(n3750), .A(n3424), .ZN(U3211) );
  INV_X1 U4241 ( .A(n3140), .ZN(n3427) );
  AOI21_X1 U4242 ( .B1(n3426), .B2(n3428), .A(n3427), .ZN(n3431) );
  AOI22_X1 U4243 ( .A1(n3757), .A2(n2921), .B1(REG3_REG_2__SCAN_IN), .B2(n3467), .ZN(n3430) );
  AOI22_X1 U4244 ( .A1(n4293), .A2(n3758), .B1(n3759), .B2(n2925), .ZN(n3429)
         );
  OAI211_X1 U4245 ( .C1(n3431), .C2(n3750), .A(n3430), .B(n3429), .ZN(U3234)
         );
  INV_X1 U4246 ( .A(n3433), .ZN(n3438) );
  AOI22_X1 U4247 ( .A1(n3434), .A2(n4578), .B1(REG2_REG_28__SCAN_IN), .B2(
        n1998), .ZN(n3435) );
  OAI21_X1 U4248 ( .B1(n3436), .B2(n4234), .A(n3435), .ZN(n3437) );
  AOI21_X1 U4249 ( .B1(n3438), .B2(n4581), .A(n3437), .ZN(n3439) );
  OAI21_X1 U4250 ( .B1(n3432), .B2(n4283), .A(n3439), .ZN(U3262) );
  XNOR2_X1 U4251 ( .A(n3441), .B(n3440), .ZN(n3442) );
  XNOR2_X1 U4252 ( .A(n3443), .B(n3442), .ZN(n3450) );
  AOI22_X1 U4253 ( .A1(n3444), .A2(n3758), .B1(n3759), .B2(n3923), .ZN(n3449)
         );
  NAND2_X1 U4254 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n4510) );
  NAND2_X1 U4255 ( .A1(n3757), .A2(n3925), .ZN(n3445) );
  OAI211_X1 U4256 ( .C1(n3762), .C2(n3446), .A(n4510), .B(n3445), .ZN(n3447)
         );
  INV_X1 U4257 ( .A(n3447), .ZN(n3448) );
  OAI211_X1 U4258 ( .C1(n3450), .C2(n3750), .A(n3449), .B(n3448), .ZN(U3212)
         );
  AND2_X1 U4259 ( .A1(n3720), .A2(n3451), .ZN(n3453) );
  OAI211_X1 U4260 ( .C1(n3453), .C2(n3452), .A(n3764), .B(n3639), .ZN(n3457)
         );
  AOI22_X1 U4261 ( .A1(n4149), .A2(n3757), .B1(n3845), .B2(n3724), .ZN(n3456)
         );
  AOI22_X1 U4262 ( .A1(n3920), .A2(n3759), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3455) );
  NAND2_X1 U4263 ( .A1(n3747), .A2(n4122), .ZN(n3454) );
  NAND4_X1 U4264 ( .A1(n3457), .A2(n3456), .A3(n3455), .A4(n3454), .ZN(U3213)
         );
  XOR2_X1 U4265 ( .A(n3459), .B(n3458), .Z(n3466) );
  AOI22_X1 U4266 ( .A1(n3460), .A2(n3758), .B1(n3757), .B2(n4225), .ZN(n3465)
         );
  NAND2_X1 U4267 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3986) );
  NAND2_X1 U4268 ( .A1(n3759), .A2(n4188), .ZN(n3461) );
  OAI211_X1 U4269 ( .C1(n3762), .C2(n3462), .A(n3986), .B(n3461), .ZN(n3463)
         );
  INV_X1 U4270 ( .A(n3463), .ZN(n3464) );
  OAI211_X1 U4271 ( .C1(n3466), .C2(n3750), .A(n3465), .B(n3464), .ZN(U3216)
         );
  AOI22_X1 U4272 ( .A1(n2336), .A2(n3758), .B1(n3759), .B2(n4558), .ZN(n3473)
         );
  AOI22_X1 U4273 ( .A1(n3757), .A2(n2969), .B1(n3467), .B2(REG3_REG_1__SCAN_IN), .ZN(n3472) );
  OAI211_X1 U4274 ( .C1(n3470), .C2(n3469), .A(n3764), .B(n3468), .ZN(n3471)
         );
  NAND3_X1 U4275 ( .A1(n3473), .A2(n3472), .A3(n3471), .ZN(U3219) );
  NAND3_X1 U4276 ( .A1(IR_REG_23__SCAN_IN), .A2(REG3_REG_24__SCAN_IN), .A3(
        REG3_REG_15__SCAN_IN), .ZN(n3476) );
  NAND4_X1 U4277 ( .A1(IR_REG_3__SCAN_IN), .A2(REG0_REG_28__SCAN_IN), .A3(
        REG0_REG_12__SCAN_IN), .A4(n3527), .ZN(n3475) );
  INV_X1 U4278 ( .A(DATAI_15_), .ZN(n4598) );
  NAND4_X1 U4279 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        REG0_REG_21__SCAN_IN), .A4(n4598), .ZN(n3474) );
  OR4_X1 U4280 ( .A1(REG0_REG_18__SCAN_IN), .A2(n3476), .A3(n3475), .A4(n3474), 
        .ZN(n3497) );
  NAND4_X1 U4281 ( .A1(REG1_REG_3__SCAN_IN), .A2(REG1_REG_17__SCAN_IN), .A3(
        DATAO_REG_0__SCAN_IN), .A4(n2835), .ZN(n3496) );
  NOR4_X1 U4282 ( .A1(REG3_REG_12__SCAN_IN), .A2(REG2_REG_26__SCAN_IN), .A3(
        REG2_REG_23__SCAN_IN), .A4(n3570), .ZN(n3486) );
  INV_X1 U4283 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3515) );
  NAND4_X1 U4284 ( .A1(DATAI_27_), .A2(REG2_REG_4__SCAN_IN), .A3(n3515), .A4(
        n3571), .ZN(n3478) );
  INV_X1 U4285 ( .A(ADDR_REG_11__SCAN_IN), .ZN(n3501) );
  NAND4_X1 U4286 ( .A1(REG1_REG_5__SCAN_IN), .A2(REG1_REG_31__SCAN_IN), .A3(
        n3503), .A4(n3501), .ZN(n3477) );
  NOR4_X1 U4287 ( .A1(DATAO_REG_11__SCAN_IN), .A2(n3479), .A3(n3478), .A4(
        n3477), .ZN(n3485) );
  NOR4_X1 U4288 ( .A1(REG3_REG_5__SCAN_IN), .A2(REG2_REG_25__SCAN_IN), .A3(
        REG1_REG_12__SCAN_IN), .A4(REG2_REG_10__SCAN_IN), .ZN(n3484) );
  NAND4_X1 U4289 ( .A1(REG2_REG_9__SCAN_IN), .A2(D_REG_0__SCAN_IN), .A3(
        DATAI_8_), .A4(n3385), .ZN(n3482) );
  NAND3_X1 U4290 ( .A1(REG3_REG_17__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        DATAO_REG_31__SCAN_IN), .ZN(n3481) );
  NAND4_X1 U4291 ( .A1(D_REG_5__SCAN_IN), .A2(REG2_REG_11__SCAN_IN), .A3(
        REG0_REG_0__SCAN_IN), .A4(DATAI_30_), .ZN(n3480) );
  NOR4_X1 U4292 ( .A1(ADDR_REG_8__SCAN_IN), .A2(n3482), .A3(n3481), .A4(n3480), 
        .ZN(n3483) );
  NAND4_X1 U4293 ( .A1(n3486), .A2(n3485), .A3(n3484), .A4(n3483), .ZN(n3495)
         );
  NAND3_X1 U4294 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .ZN(n3488) );
  NAND2_X1 U4295 ( .A1(REG2_REG_3__SCAN_IN), .A2(DATAI_2_), .ZN(n3487) );
  OR4_X1 U4296 ( .A1(n3488), .A2(n3487), .A3(DATAI_28_), .A4(DATAI_13_), .ZN(
        n3493) );
  NOR4_X1 U4297 ( .A1(IR_REG_11__SCAN_IN), .A2(DATAI_16_), .A3(
        REG2_REG_24__SCAN_IN), .A4(n4328), .ZN(n3489) );
  NAND4_X1 U4298 ( .A1(n3491), .A2(n3490), .A3(IR_REG_27__SCAN_IN), .A4(n3489), 
        .ZN(n3492) );
  OR4_X1 U4299 ( .A1(n3493), .A2(REG0_REG_13__SCAN_IN), .A3(
        DATAO_REG_17__SCAN_IN), .A4(n3492), .ZN(n3494) );
  NOR4_X1 U4300 ( .A1(n3497), .A2(n3496), .A3(n3495), .A4(n3494), .ZN(n3499)
         );
  OAI21_X1 U4301 ( .B1(n3499), .B2(n3498), .A(keyinput52), .ZN(n3612) );
  AOI22_X1 U4302 ( .A1(n3628), .A2(keyinput34), .B1(keyinput28), .B2(n3501), 
        .ZN(n3500) );
  OAI221_X1 U4303 ( .B1(n3628), .B2(keyinput34), .C1(n3501), .C2(keyinput28), 
        .A(n3500), .ZN(n3510) );
  AOI22_X1 U4304 ( .A1(n4653), .A2(keyinput24), .B1(n3503), .B2(keyinput26), 
        .ZN(n3502) );
  OAI221_X1 U4305 ( .B1(n4653), .B2(keyinput24), .C1(n3503), .C2(keyinput26), 
        .A(n3502), .ZN(n3509) );
  AOI22_X1 U4306 ( .A1(n3505), .A2(keyinput30), .B1(n3385), .B2(keyinput20), 
        .ZN(n3504) );
  OAI221_X1 U4307 ( .B1(n3505), .B2(keyinput30), .C1(n3385), .C2(keyinput20), 
        .A(n3504), .ZN(n3508) );
  AOI22_X1 U4308 ( .A1(n2477), .A2(keyinput22), .B1(n4587), .B2(keyinput25), 
        .ZN(n3506) );
  OAI221_X1 U4309 ( .B1(n2477), .B2(keyinput22), .C1(n4587), .C2(keyinput25), 
        .A(n3506), .ZN(n3507) );
  NOR4_X1 U4310 ( .A1(n3510), .A2(n3509), .A3(n3508), .A4(n3507), .ZN(n3611)
         );
  AOI22_X1 U4311 ( .A1(n4596), .A2(keyinput6), .B1(n2835), .B2(keyinput8), 
        .ZN(n3511) );
  OAI221_X1 U4312 ( .B1(n4596), .B2(keyinput6), .C1(n2835), .C2(keyinput8), 
        .A(n3511), .ZN(n3521) );
  AOI22_X1 U4313 ( .A1(n2106), .A2(keyinput23), .B1(keyinput3), .B2(n3513), 
        .ZN(n3512) );
  OAI221_X1 U4314 ( .B1(n2106), .B2(keyinput23), .C1(n3513), .C2(keyinput3), 
        .A(n3512), .ZN(n3520) );
  AOI22_X1 U4315 ( .A1(n3516), .A2(keyinput36), .B1(keyinput40), .B2(n3515), 
        .ZN(n3514) );
  OAI221_X1 U4316 ( .B1(n3516), .B2(keyinput36), .C1(n3515), .C2(keyinput40), 
        .A(n3514), .ZN(n3519) );
  XNOR2_X1 U4317 ( .A(n3517), .B(keyinput56), .ZN(n3518) );
  OR4_X1 U4318 ( .A1(n3521), .A2(n3520), .A3(n3519), .A4(n3518), .ZN(n3543) );
  AOI22_X1 U4319 ( .A1(n3524), .A2(keyinput46), .B1(keyinput58), .B2(n3523), 
        .ZN(n3522) );
  OAI221_X1 U4320 ( .B1(n3524), .B2(keyinput46), .C1(n3523), .C2(keyinput58), 
        .A(n3522), .ZN(n3542) );
  INV_X1 U4321 ( .A(D_REG_3__SCAN_IN), .ZN(n4588) );
  INV_X1 U4322 ( .A(D_REG_29__SCAN_IN), .ZN(n4583) );
  AOI22_X1 U4323 ( .A1(n4588), .A2(keyinput53), .B1(keyinput50), .B2(n4583), 
        .ZN(n3525) );
  OAI221_X1 U4324 ( .B1(n4588), .B2(keyinput53), .C1(n4583), .C2(keyinput50), 
        .A(n3525), .ZN(n3541) );
  AOI22_X1 U4325 ( .A1(n3527), .A2(keyinput60), .B1(keyinput49), .B2(n4442), 
        .ZN(n3526) );
  OAI221_X1 U4326 ( .B1(n3527), .B2(keyinput60), .C1(n4442), .C2(keyinput49), 
        .A(n3526), .ZN(n3539) );
  AOI22_X1 U4327 ( .A1(n3530), .A2(keyinput54), .B1(keyinput61), .B2(n3529), 
        .ZN(n3528) );
  OAI221_X1 U4328 ( .B1(n3530), .B2(keyinput54), .C1(n3529), .C2(keyinput61), 
        .A(n3528), .ZN(n3538) );
  AOI22_X1 U4329 ( .A1(n3532), .A2(keyinput5), .B1(keyinput4), .B2(n4328), 
        .ZN(n3531) );
  OAI221_X1 U4330 ( .B1(n3532), .B2(keyinput5), .C1(n4328), .C2(keyinput4), 
        .A(n3531), .ZN(n3537) );
  AOI22_X1 U4331 ( .A1(n3535), .A2(keyinput17), .B1(keyinput18), .B2(n3534), 
        .ZN(n3533) );
  OAI221_X1 U4332 ( .B1(n3535), .B2(keyinput17), .C1(n3534), .C2(keyinput18), 
        .A(n3533), .ZN(n3536) );
  OR4_X1 U4333 ( .A1(n3539), .A2(n3538), .A3(n3537), .A4(n3536), .ZN(n3540) );
  NOR4_X1 U4334 ( .A1(n3543), .A2(n3542), .A3(n3541), .A4(n3540), .ZN(n3610)
         );
  AOI22_X1 U4335 ( .A1(n3545), .A2(keyinput9), .B1(n2378), .B2(keyinput10), 
        .ZN(n3544) );
  OAI221_X1 U4336 ( .B1(n3545), .B2(keyinput9), .C1(n2378), .C2(keyinput10), 
        .A(n3544), .ZN(n3549) );
  INV_X1 U4337 ( .A(D_REG_5__SCAN_IN), .ZN(n4586) );
  AOI22_X1 U4338 ( .A1(n2341), .A2(keyinput31), .B1(n4586), .B2(keyinput59), 
        .ZN(n3546) );
  OAI221_X1 U4339 ( .B1(n2341), .B2(keyinput31), .C1(n4586), .C2(keyinput59), 
        .A(n3546), .ZN(n3548) );
  INV_X1 U4340 ( .A(D_REG_23__SCAN_IN), .ZN(n4584) );
  XNOR2_X1 U4341 ( .A(n4584), .B(keyinput27), .ZN(n3547) );
  NOR3_X1 U4342 ( .A1(n3549), .A2(n3548), .A3(n3547), .ZN(n3568) );
  INV_X1 U4343 ( .A(ADDR_REG_8__SCAN_IN), .ZN(n3551) );
  AOI22_X1 U4344 ( .A1(n3552), .A2(keyinput39), .B1(keyinput19), .B2(n3551), 
        .ZN(n3550) );
  OAI221_X1 U4345 ( .B1(n3552), .B2(keyinput39), .C1(n3551), .C2(keyinput19), 
        .A(n3550), .ZN(n3561) );
  INV_X1 U4346 ( .A(DATAI_30_), .ZN(n3555) );
  AOI22_X1 U4347 ( .A1(n3555), .A2(keyinput7), .B1(n3554), .B2(keyinput15), 
        .ZN(n3553) );
  OAI221_X1 U4348 ( .B1(n3555), .B2(keyinput7), .C1(n3554), .C2(keyinput15), 
        .A(n3553), .ZN(n3560) );
  AOI22_X1 U4349 ( .A1(n3558), .A2(keyinput33), .B1(n3557), .B2(keyinput37), 
        .ZN(n3556) );
  OAI221_X1 U4350 ( .B1(n3558), .B2(keyinput33), .C1(n3557), .C2(keyinput37), 
        .A(n3556), .ZN(n3559) );
  NOR3_X1 U4351 ( .A1(n3561), .A2(n3560), .A3(n3559), .ZN(n3567) );
  AOI22_X1 U4352 ( .A1(n4356), .A2(keyinput13), .B1(keyinput14), .B2(n3308), 
        .ZN(n3562) );
  OAI221_X1 U4353 ( .B1(n4356), .B2(keyinput13), .C1(n3308), .C2(keyinput14), 
        .A(n3562), .ZN(n3565) );
  AOI22_X1 U4354 ( .A1(n4493), .A2(keyinput35), .B1(keyinput51), .B2(n3326), 
        .ZN(n3563) );
  OAI221_X1 U4355 ( .B1(n4493), .B2(keyinput35), .C1(n3326), .C2(keyinput51), 
        .A(n3563), .ZN(n3564) );
  NOR2_X1 U4356 ( .A1(n3565), .A2(n3564), .ZN(n3566) );
  NAND3_X1 U4357 ( .A1(n3568), .A2(n3567), .A3(n3566), .ZN(n3608) );
  AOI22_X1 U4358 ( .A1(n3571), .A2(keyinput41), .B1(keyinput32), .B2(n3570), 
        .ZN(n3569) );
  OAI221_X1 U4359 ( .B1(n3571), .B2(keyinput41), .C1(n3570), .C2(keyinput32), 
        .A(n3569), .ZN(n3607) );
  AOI22_X1 U4360 ( .A1(n4585), .A2(keyinput11), .B1(keyinput0), .B2(n4438), 
        .ZN(n3572) );
  OAI221_X1 U4361 ( .B1(n4585), .B2(keyinput11), .C1(n4438), .C2(keyinput0), 
        .A(n3572), .ZN(n3573) );
  INV_X1 U4362 ( .A(n3573), .ZN(n3579) );
  XNOR2_X1 U4363 ( .A(keyinput45), .B(n4598), .ZN(n3575) );
  XNOR2_X1 U4364 ( .A(keyinput47), .B(n2722), .ZN(n3574) );
  NOR2_X1 U4365 ( .A1(n3575), .A2(n3574), .ZN(n3578) );
  XNOR2_X1 U4366 ( .A(DATAI_2_), .B(keyinput44), .ZN(n3577) );
  XNOR2_X1 U4367 ( .A(IR_REG_13__SCAN_IN), .B(keyinput12), .ZN(n3576) );
  NAND4_X1 U4368 ( .A1(n3579), .A2(n3578), .A3(n3577), .A4(n3576), .ZN(n3606)
         );
  AOI22_X1 U4369 ( .A1(n2781), .A2(keyinput29), .B1(keyinput43), .B2(n3581), 
        .ZN(n3580) );
  OAI221_X1 U4370 ( .B1(n2781), .B2(keyinput29), .C1(n3581), .C2(keyinput43), 
        .A(n3580), .ZN(n3582) );
  INV_X1 U4371 ( .A(n3582), .ZN(n3604) );
  XNOR2_X1 U4372 ( .A(IR_REG_5__SCAN_IN), .B(keyinput63), .ZN(n3588) );
  NAND2_X1 U4373 ( .A1(n2398), .A2(keyinput38), .ZN(n3587) );
  INV_X1 U4374 ( .A(keyinput38), .ZN(n3583) );
  NAND2_X1 U4375 ( .A1(n3583), .A2(REG2_REG_4__SCAN_IN), .ZN(n3586) );
  INV_X1 U4376 ( .A(keyinput52), .ZN(n3584) );
  NAND2_X1 U4377 ( .A1(n3584), .A2(IR_REG_8__SCAN_IN), .ZN(n3585) );
  NAND4_X1 U4378 ( .A1(n3588), .A2(n3587), .A3(n3586), .A4(n3585), .ZN(n3591)
         );
  INV_X1 U4379 ( .A(REG2_REG_24__SCAN_IN), .ZN(n3589) );
  XNOR2_X1 U4380 ( .A(keyinput2), .B(n3589), .ZN(n3590) );
  NOR2_X1 U4381 ( .A1(n3591), .A2(n3590), .ZN(n3603) );
  XNOR2_X1 U4382 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput55), .ZN(n3595) );
  XNOR2_X1 U4383 ( .A(REG3_REG_24__SCAN_IN), .B(keyinput42), .ZN(n3594) );
  XNOR2_X1 U4384 ( .A(IR_REG_21__SCAN_IN), .B(keyinput1), .ZN(n3593) );
  XNOR2_X1 U4385 ( .A(IR_REG_3__SCAN_IN), .B(keyinput62), .ZN(n3592) );
  NAND4_X1 U4386 ( .A1(n3595), .A2(n3594), .A3(n3593), .A4(n3592), .ZN(n3601)
         );
  XNOR2_X1 U4387 ( .A(REG0_REG_21__SCAN_IN), .B(keyinput48), .ZN(n3599) );
  XNOR2_X1 U4388 ( .A(IR_REG_23__SCAN_IN), .B(keyinput21), .ZN(n3598) );
  XNOR2_X1 U4389 ( .A(IR_REG_24__SCAN_IN), .B(keyinput57), .ZN(n3597) );
  XNOR2_X1 U4390 ( .A(IR_REG_27__SCAN_IN), .B(keyinput16), .ZN(n3596) );
  NAND4_X1 U4391 ( .A1(n3599), .A2(n3598), .A3(n3597), .A4(n3596), .ZN(n3600)
         );
  NOR2_X1 U4392 ( .A1(n3601), .A2(n3600), .ZN(n3602) );
  NAND3_X1 U4393 ( .A1(n3604), .A2(n3603), .A3(n3602), .ZN(n3605) );
  NOR4_X1 U4394 ( .A1(n3608), .A2(n3607), .A3(n3606), .A4(n3605), .ZN(n3609)
         );
  NAND4_X1 U4395 ( .A1(n3612), .A2(n3611), .A3(n3610), .A4(n3609), .ZN(n3622)
         );
  XNOR2_X1 U4396 ( .A(n3615), .B(n3614), .ZN(n3616) );
  XNOR2_X1 U4397 ( .A(n3613), .B(n3616), .ZN(n3620) );
  AOI22_X1 U4398 ( .A1(n4149), .A2(n3759), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3618) );
  AOI22_X1 U4399 ( .A1(n4150), .A2(n3758), .B1(n3757), .B2(n4188), .ZN(n3617)
         );
  OAI211_X1 U4400 ( .C1(n3762), .C2(n4146), .A(n3618), .B(n3617), .ZN(n3619)
         );
  AOI21_X1 U4401 ( .B1(n3620), .B2(n3764), .A(n3619), .ZN(n3621) );
  XOR2_X1 U4402 ( .A(n3622), .B(n3621), .Z(U3220) );
  XNOR2_X1 U4403 ( .A(n3625), .B(n3624), .ZN(n3626) );
  XNOR2_X1 U4404 ( .A(n3623), .B(n3626), .ZN(n3634) );
  AOI22_X1 U4405 ( .A1(n3627), .A2(n3758), .B1(n3759), .B2(n3925), .ZN(n3633)
         );
  NOR2_X1 U4406 ( .A1(n3628), .A2(STATE_REG_SCAN_IN), .ZN(n4494) );
  NOR2_X1 U4407 ( .A1(n3762), .A2(n3629), .ZN(n3630) );
  AOI211_X1 U4408 ( .C1(n3757), .C2(n3631), .A(n4494), .B(n3630), .ZN(n3632)
         );
  OAI211_X1 U4409 ( .C1(n3634), .C2(n3750), .A(n3633), .B(n3632), .ZN(U3221)
         );
  INV_X1 U4410 ( .A(n3635), .ZN(n3636) );
  NAND2_X1 U4411 ( .A1(n3639), .A2(n3636), .ZN(n3682) );
  AOI21_X1 U4412 ( .B1(n3639), .B2(n3638), .A(n3637), .ZN(n3684) );
  OAI21_X1 U4413 ( .B1(n3642), .B2(n3641), .A(n3640), .ZN(n3643) );
  XNOR2_X1 U4414 ( .A(n3644), .B(n3643), .ZN(n3649) );
  OAI22_X1 U4415 ( .A1(n4115), .A2(n3744), .B1(n3702), .B2(n4079), .ZN(n3647)
         );
  OAI22_X1 U4416 ( .A1(n4033), .A2(n3701), .B1(STATE_REG_SCAN_IN), .B2(n3645), 
        .ZN(n3646) );
  AOI211_X1 U4417 ( .C1(n4081), .C2(n3747), .A(n3647), .B(n3646), .ZN(n3648)
         );
  OAI21_X1 U4418 ( .B1(n3649), .B2(n3750), .A(n3648), .ZN(U3222) );
  NOR2_X1 U4419 ( .A1(n3650), .A2(n3651), .ZN(n3754) );
  NAND2_X1 U4420 ( .A1(n3650), .A2(n3651), .ZN(n3752) );
  OAI21_X1 U4421 ( .B1(n3754), .B2(n3669), .A(n3752), .ZN(n3652) );
  XNOR2_X1 U4422 ( .A(n3672), .B(n3671), .ZN(n3668) );
  XNOR2_X1 U4423 ( .A(n3652), .B(n3668), .ZN(n3657) );
  INV_X1 U4424 ( .A(n4248), .ZN(n4247) );
  AOI22_X1 U4425 ( .A1(n4247), .A2(n3758), .B1(n3757), .B2(n3923), .ZN(n3656)
         );
  NOR2_X1 U4426 ( .A1(n3653), .A2(STATE_REG_SCAN_IN), .ZN(n4523) );
  NOR2_X1 U4427 ( .A1(n3701), .A2(n4242), .ZN(n3654) );
  AOI211_X1 U4428 ( .C1(n4249), .C2(n3747), .A(n4523), .B(n3654), .ZN(n3655)
         );
  OAI211_X1 U4429 ( .C1(n3657), .C2(n3750), .A(n3656), .B(n3655), .ZN(U3223)
         );
  OAI211_X1 U4430 ( .C1(n3660), .C2(n3659), .A(n3658), .B(n3764), .ZN(n3667)
         );
  AOI22_X1 U4431 ( .A1(n3661), .A2(n3758), .B1(n3759), .B2(n3932), .ZN(n3666)
         );
  NOR2_X1 U4432 ( .A1(n3762), .A2(n3662), .ZN(n3663) );
  AOI211_X1 U4433 ( .C1(n3757), .C2(n3934), .A(n3664), .B(n3663), .ZN(n3665)
         );
  NAND3_X1 U4434 ( .A1(n3667), .A2(n3666), .A3(n3665), .ZN(U3224) );
  AOI211_X1 U4435 ( .C1(n3669), .C2(n3752), .A(n3668), .B(n3754), .ZN(n3670)
         );
  AOI21_X1 U4436 ( .B1(n3672), .B2(n3671), .A(n3670), .ZN(n3676) );
  XNOR2_X1 U4437 ( .A(n3674), .B(n3673), .ZN(n3675) );
  XNOR2_X1 U4438 ( .A(n3676), .B(n3675), .ZN(n3680) );
  AOI22_X1 U4439 ( .A1(n4231), .A2(n3758), .B1(n3759), .B2(n4225), .ZN(n3678)
         );
  AND2_X1 U4440 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4534) );
  AOI21_X1 U4441 ( .B1(n3757), .B2(n3922), .A(n4534), .ZN(n3677) );
  OAI211_X1 U4442 ( .C1(n3762), .C2(n4235), .A(n3678), .B(n3677), .ZN(n3679)
         );
  AOI21_X1 U4443 ( .B1(n3680), .B2(n3764), .A(n3679), .ZN(n3681) );
  INV_X1 U4444 ( .A(n3681), .ZN(U3225) );
  INV_X1 U4445 ( .A(n3682), .ZN(n3683) );
  NOR2_X1 U4446 ( .A1(n3684), .A2(n3683), .ZN(n3686) );
  XNOR2_X1 U4447 ( .A(n3686), .B(n3685), .ZN(n3693) );
  AOI22_X1 U4448 ( .A1(n3921), .A2(n3757), .B1(n3687), .B2(n3724), .ZN(n3692)
         );
  INV_X1 U4449 ( .A(n4095), .ZN(n3690) );
  OAI22_X1 U4450 ( .A1(n3745), .A2(n3701), .B1(STATE_REG_SCAN_IN), .B2(n3688), 
        .ZN(n3689) );
  AOI21_X1 U4451 ( .B1(n3690), .B2(n3747), .A(n3689), .ZN(n3691) );
  OAI211_X1 U4452 ( .C1(n3693), .C2(n3750), .A(n3692), .B(n3691), .ZN(U3226)
         );
  INV_X1 U4453 ( .A(n3694), .ZN(n3699) );
  AOI21_X1 U4454 ( .B1(n3698), .B2(n3696), .A(n3695), .ZN(n3697) );
  AOI21_X1 U4455 ( .B1(n3699), .B2(n3698), .A(n3697), .ZN(n3706) );
  OAI22_X1 U4456 ( .A1(n3701), .A2(n4168), .B1(STATE_REG_SCAN_IN), .B2(n3700), 
        .ZN(n3704) );
  OAI22_X1 U4457 ( .A1(n3702), .A2(n4176), .B1(n3744), .B2(n4207), .ZN(n3703)
         );
  AOI211_X1 U4458 ( .C1(n4177), .C2(n3747), .A(n3704), .B(n3703), .ZN(n3705)
         );
  OAI21_X1 U4459 ( .B1(n3706), .B2(n3750), .A(n3705), .ZN(U3230) );
  INV_X1 U4460 ( .A(n3708), .ZN(n3710) );
  NOR2_X1 U4461 ( .A1(n3710), .A2(n3709), .ZN(n3711) );
  XNOR2_X1 U4462 ( .A(n3707), .B(n3711), .ZN(n3719) );
  AOI22_X1 U4463 ( .A1(n3712), .A2(n3724), .B1(n3759), .B2(n3924), .ZN(n3718)
         );
  NOR2_X1 U4464 ( .A1(n3713), .A2(STATE_REG_SCAN_IN), .ZN(n3974) );
  NOR2_X1 U4465 ( .A1(n3744), .A2(n3714), .ZN(n3715) );
  AOI211_X1 U4466 ( .C1(n3716), .C2(n3747), .A(n3974), .B(n3715), .ZN(n3717)
         );
  OAI211_X1 U4467 ( .C1(n3719), .C2(n3750), .A(n3718), .B(n3717), .ZN(U3231)
         );
  OAI21_X1 U4468 ( .B1(n3722), .B2(n3721), .A(n3720), .ZN(n3723) );
  NAND2_X1 U4469 ( .A1(n3723), .A2(n3764), .ZN(n3728) );
  AOI22_X1 U4470 ( .A1(n4129), .A2(n3757), .B1(n4128), .B2(n3724), .ZN(n3727)
         );
  AOI22_X1 U4471 ( .A1(n3921), .A2(n3759), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3726) );
  NAND2_X1 U4472 ( .A1(n3747), .A2(n4137), .ZN(n3725) );
  NAND4_X1 U4473 ( .A1(n3728), .A2(n3727), .A3(n3726), .A4(n3725), .ZN(U3232)
         );
  INV_X1 U4474 ( .A(n3730), .ZN(n3732) );
  NOR2_X1 U4475 ( .A1(n3732), .A2(n3731), .ZN(n3733) );
  XNOR2_X1 U4476 ( .A(n3729), .B(n3733), .ZN(n3738) );
  AOI22_X1 U4477 ( .A1(n4204), .A2(n3758), .B1(n3759), .B2(n4166), .ZN(n3736)
         );
  AOI21_X1 U4478 ( .B1(n3757), .B2(n4205), .A(n3734), .ZN(n3735) );
  OAI211_X1 U4479 ( .C1(n3762), .C2(n4217), .A(n3736), .B(n3735), .ZN(n3737)
         );
  AOI21_X1 U4480 ( .B1(n3738), .B2(n3764), .A(n3737), .ZN(n3739) );
  INV_X1 U4481 ( .A(n3739), .ZN(U3235) );
  NAND2_X1 U4482 ( .A1(n2032), .A2(n3740), .ZN(n3741) );
  XNOR2_X1 U4483 ( .A(n3742), .B(n3741), .ZN(n3751) );
  OAI22_X1 U4484 ( .A1(n3745), .A2(n3744), .B1(STATE_REG_SCAN_IN), .B2(n3743), 
        .ZN(n3746) );
  AOI21_X1 U4485 ( .B1(n4055), .B2(n3758), .A(n3746), .ZN(n3749) );
  AOI22_X1 U4486 ( .A1(n3919), .A2(n3759), .B1(n4063), .B2(n3747), .ZN(n3748)
         );
  OAI211_X1 U4487 ( .C1(n3751), .C2(n3750), .A(n3749), .B(n3748), .ZN(U3237)
         );
  INV_X1 U4488 ( .A(n3752), .ZN(n3753) );
  NOR2_X1 U4489 ( .A1(n3754), .A2(n3753), .ZN(n3756) );
  XNOR2_X1 U4490 ( .A(n3756), .B(n3755), .ZN(n3765) );
  AOI22_X1 U4491 ( .A1(n4275), .A2(n3758), .B1(n3757), .B2(n3924), .ZN(n3761)
         );
  AND2_X1 U4492 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4517) );
  AOI21_X1 U4493 ( .B1(n3759), .B2(n3922), .A(n4517), .ZN(n3760) );
  OAI211_X1 U4494 ( .C1(n3762), .C2(n4277), .A(n3761), .B(n3760), .ZN(n3763)
         );
  AOI21_X1 U4495 ( .B1(n3765), .B2(n3764), .A(n3763), .ZN(n3766) );
  INV_X1 U4496 ( .A(n3766), .ZN(U3238) );
  AND2_X1 U4497 ( .A1(n2969), .A2(n3767), .ZN(n3863) );
  INV_X1 U4498 ( .A(n3863), .ZN(n3769) );
  OAI211_X1 U4499 ( .C1(n4554), .C2(n4452), .A(n3769), .B(n3768), .ZN(n3771)
         );
  NAND3_X1 U4500 ( .A1(n3771), .A2(n3770), .A3(n2970), .ZN(n3773) );
  OAI211_X1 U4501 ( .C1(n3774), .C2(n2926), .A(n3773), .B(n3772), .ZN(n3777)
         );
  NAND3_X1 U4502 ( .A1(n3777), .A2(n3776), .A3(n3775), .ZN(n3780) );
  NAND4_X1 U4503 ( .A1(n3780), .A2(n3779), .A3(n3778), .A4(n3791), .ZN(n3783)
         );
  AND3_X1 U4504 ( .A1(n3783), .A2(n3782), .A3(n3781), .ZN(n3788) );
  NAND2_X1 U4505 ( .A1(n3785), .A2(n3784), .ZN(n3794) );
  OAI211_X1 U4506 ( .C1(n3788), .C2(n3794), .A(n3787), .B(n3786), .ZN(n3790)
         );
  NAND4_X1 U4507 ( .A1(n3790), .A2(n3797), .A3(n3798), .A4(n3789), .ZN(n3807)
         );
  INV_X1 U4508 ( .A(n3791), .ZN(n3795) );
  NOR4_X1 U4509 ( .A1(n3795), .A2(n3794), .A3(n3793), .A4(n3792), .ZN(n3801)
         );
  INV_X1 U4510 ( .A(n3796), .ZN(n3800) );
  NAND2_X1 U4511 ( .A1(n3798), .A2(n3797), .ZN(n3799) );
  NAND2_X1 U4512 ( .A1(n3799), .A2(n3809), .ZN(n3883) );
  OAI21_X1 U4513 ( .B1(n3801), .B2(n3800), .A(n3883), .ZN(n3806) );
  NAND3_X1 U4514 ( .A1(n3804), .A2(n3803), .A3(n3802), .ZN(n3805) );
  AOI21_X1 U4515 ( .B1(n3807), .B2(n3806), .A(n3805), .ZN(n3814) );
  NAND2_X1 U4516 ( .A1(n3809), .A2(n3808), .ZN(n3884) );
  INV_X1 U4517 ( .A(n3884), .ZN(n3811) );
  INV_X1 U4518 ( .A(n3883), .ZN(n3810) );
  AOI21_X1 U4519 ( .B1(n3812), .B2(n3811), .A(n3810), .ZN(n3813) );
  OAI21_X1 U4520 ( .B1(n3814), .B2(n3813), .A(n4104), .ZN(n3816) );
  AOI21_X1 U4521 ( .B1(n3816), .B2(n3885), .A(n3815), .ZN(n3817) );
  NOR2_X1 U4522 ( .A1(n3817), .A2(n3887), .ZN(n3822) );
  INV_X1 U4523 ( .A(n3818), .ZN(n3846) );
  OAI21_X1 U4524 ( .B1(n3820), .B2(n3846), .A(n3819), .ZN(n3821) );
  OAI21_X1 U4525 ( .B1(n3822), .B2(n3821), .A(n3891), .ZN(n3824) );
  INV_X1 U4526 ( .A(n3895), .ZN(n3823) );
  AOI21_X1 U4527 ( .B1(n3892), .B2(n3824), .A(n3823), .ZN(n3827) );
  NAND2_X1 U4528 ( .A1(n1999), .A2(DATAI_29_), .ZN(n3839) );
  OAI21_X1 U4529 ( .B1(n3840), .B2(n4021), .A(n4014), .ZN(n3901) );
  INV_X1 U4530 ( .A(n3825), .ZN(n3826) );
  NOR4_X1 U4531 ( .A1(n3827), .A2(n3901), .A3(n3841), .A4(n3826), .ZN(n3838)
         );
  NAND2_X1 U4532 ( .A1(n1999), .A2(DATAI_31_), .ZN(n3996) );
  NAND2_X1 U4533 ( .A1(n3995), .A2(n3996), .ZN(n3833) );
  INV_X1 U4534 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4302) );
  NAND2_X1 U4535 ( .A1(n2447), .A2(REG2_REG_30__SCAN_IN), .ZN(n3830) );
  INV_X1 U4536 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4400) );
  OR2_X1 U4537 ( .A1(n2764), .A2(n4400), .ZN(n3829) );
  OAI211_X1 U4538 ( .C1(n3831), .C2(n4302), .A(n3830), .B(n3829), .ZN(n4019)
         );
  NAND2_X1 U4539 ( .A1(n1999), .A2(DATAI_30_), .ZN(n4000) );
  OR2_X1 U4540 ( .A1(n4019), .A2(n4000), .ZN(n3832) );
  NAND2_X1 U4541 ( .A1(n3833), .A2(n3832), .ZN(n3854) );
  AOI21_X1 U4542 ( .B1(n3840), .B2(n4021), .A(n3854), .ZN(n3900) );
  OAI21_X1 U4543 ( .B1(n3897), .B2(n3901), .A(n3900), .ZN(n3837) );
  INV_X1 U4544 ( .A(n3833), .ZN(n3836) );
  NAND2_X1 U4545 ( .A1(n4019), .A2(n4000), .ZN(n3906) );
  OR2_X1 U4546 ( .A1(n3995), .A2(n3996), .ZN(n3834) );
  NAND2_X1 U4547 ( .A1(n3906), .A2(n3834), .ZN(n3853) );
  INV_X1 U4548 ( .A(n3853), .ZN(n3835) );
  OAI22_X1 U4549 ( .A1(n3838), .A2(n3837), .B1(n3836), .B2(n3835), .ZN(n3912)
         );
  INV_X1 U4550 ( .A(n4008), .ZN(n3882) );
  XNOR2_X1 U4551 ( .A(n3840), .B(n3839), .ZN(n4307) );
  INV_X1 U4552 ( .A(n3841), .ZN(n3899) );
  NAND2_X1 U4553 ( .A1(n3899), .A2(n3842), .ZN(n4053) );
  NAND2_X1 U4554 ( .A1(n4050), .A2(n3843), .ZN(n4071) );
  INV_X1 U4555 ( .A(n4071), .ZN(n3878) );
  NAND2_X1 U4556 ( .A1(n3844), .A2(n4069), .ZN(n4089) );
  INV_X1 U4557 ( .A(n4089), .ZN(n3877) );
  XNOR2_X1 U4558 ( .A(n3921), .B(n3845), .ZN(n4113) );
  NAND2_X1 U4559 ( .A1(n3846), .A2(n4110), .ZN(n4147) );
  NAND2_X1 U4560 ( .A1(n4160), .A2(n3847), .ZN(n4191) );
  NOR2_X1 U4561 ( .A1(n4191), .A2(n3848), .ZN(n3873) );
  INV_X1 U4562 ( .A(n4105), .ZN(n3849) );
  NAND2_X1 U4563 ( .A1(n3849), .A2(n4201), .ZN(n4228) );
  NAND4_X1 U4564 ( .A1(n3852), .A2(n3851), .A3(n3850), .A4(n4555), .ZN(n3868)
         );
  NOR3_X1 U4565 ( .A1(n3855), .A2(n3854), .A3(n3853), .ZN(n3862) );
  NOR2_X1 U4566 ( .A1(n3856), .A2(n3110), .ZN(n3861) );
  NOR2_X1 U4567 ( .A1(n3858), .A2(n3857), .ZN(n3859) );
  NAND4_X1 U4568 ( .A1(n3862), .A2(n3861), .A3(n3860), .A4(n3859), .ZN(n3867)
         );
  OR2_X1 U4569 ( .A1(n3863), .A2(n4554), .ZN(n4607) );
  INV_X1 U4570 ( .A(n4607), .ZN(n3865) );
  NAND2_X1 U4571 ( .A1(n3865), .A2(n3864), .ZN(n3866) );
  NOR4_X1 U4572 ( .A1(n4228), .A2(n3868), .A3(n3867), .A4(n3866), .ZN(n3872)
         );
  NOR3_X1 U4573 ( .A1(n4211), .A2(n3870), .A3(n3869), .ZN(n3871) );
  NAND4_X1 U4574 ( .A1(n3873), .A2(n2114), .A3(n3872), .A4(n3871), .ZN(n3874)
         );
  OR3_X1 U4575 ( .A1(n4147), .A2(n4256), .A3(n3874), .ZN(n3875) );
  XNOR2_X1 U4576 ( .A(n4188), .B(n4176), .ZN(n4162) );
  NOR2_X1 U4577 ( .A1(n3875), .A2(n4162), .ZN(n3876) );
  NAND4_X1 U4578 ( .A1(n3878), .A2(n3877), .A3(n4113), .A4(n3876), .ZN(n3879)
         );
  NOR2_X1 U4579 ( .A1(n4053), .A2(n3879), .ZN(n3881) );
  AND2_X1 U4580 ( .A1(n4040), .A2(n4134), .ZN(n3880) );
  NAND4_X1 U4581 ( .A1(n3882), .A2(n4307), .A3(n3881), .A4(n3880), .ZN(n3910)
         );
  OAI21_X1 U4582 ( .B1(n3379), .B2(n3884), .A(n3883), .ZN(n3890) );
  INV_X1 U4583 ( .A(n3885), .ZN(n3886) );
  NOR2_X1 U4584 ( .A1(n3887), .A2(n3886), .ZN(n3889) );
  AOI21_X1 U4585 ( .B1(n3890), .B2(n3889), .A(n3888), .ZN(n3894) );
  INV_X1 U4586 ( .A(n3891), .ZN(n3893) );
  OAI21_X1 U4587 ( .B1(n3894), .B2(n3893), .A(n3892), .ZN(n3896) );
  NAND4_X1 U4588 ( .A1(n3896), .A2(n3897), .A3(n3895), .A4(n3900), .ZN(n3905)
         );
  AOI21_X1 U4589 ( .B1(n4040), .B2(n3899), .A(n3898), .ZN(n3902) );
  INV_X1 U4590 ( .A(n4000), .ZN(n4002) );
  INV_X1 U4591 ( .A(n3995), .ZN(n3903) );
  AOI22_X1 U4592 ( .A1(n3905), .A2(n3904), .B1(n4002), .B2(n3903), .ZN(n3908)
         );
  AOI21_X1 U4593 ( .B1(n3906), .B2(n3995), .A(n3996), .ZN(n3907) );
  MUX2_X1 U4594 ( .A(n3910), .B(n3909), .S(n4452), .Z(n3911) );
  XNOR2_X1 U4595 ( .A(n3913), .B(n3987), .ZN(n3918) );
  NAND2_X1 U4596 ( .A1(n3914), .A2(n3947), .ZN(n3915) );
  OAI211_X1 U4597 ( .C1(n4451), .C2(n3917), .A(n3915), .B(B_REG_SCAN_IN), .ZN(
        n3916) );
  OAI21_X1 U4598 ( .B1(n3918), .B2(n3917), .A(n3916), .ZN(U3239) );
  MUX2_X1 U4599 ( .A(n4019), .B(DATAO_REG_30__SCAN_IN), .S(n3929), .Z(U3580)
         );
  MUX2_X1 U4600 ( .A(DATAO_REG_28__SCAN_IN), .B(n4022), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4601 ( .A(n3919), .B(DATAO_REG_27__SCAN_IN), .S(n3929), .Z(U3577)
         );
  MUX2_X1 U4602 ( .A(n4075), .B(DATAO_REG_26__SCAN_IN), .S(n3929), .Z(U3576)
         );
  MUX2_X1 U4603 ( .A(n4092), .B(DATAO_REG_25__SCAN_IN), .S(n3929), .Z(U3575)
         );
  MUX2_X1 U4604 ( .A(n3920), .B(DATAO_REG_24__SCAN_IN), .S(n3929), .Z(U3574)
         );
  MUX2_X1 U4605 ( .A(n3921), .B(DATAO_REG_23__SCAN_IN), .S(n3929), .Z(U3573)
         );
  MUX2_X1 U4606 ( .A(n4149), .B(DATAO_REG_22__SCAN_IN), .S(n3929), .Z(U3572)
         );
  MUX2_X1 U4607 ( .A(n4129), .B(DATAO_REG_21__SCAN_IN), .S(n3929), .Z(U3571)
         );
  MUX2_X1 U4608 ( .A(n4188), .B(DATAO_REG_20__SCAN_IN), .S(n3929), .Z(U3570)
         );
  MUX2_X1 U4609 ( .A(n4166), .B(DATAO_REG_19__SCAN_IN), .S(n3929), .Z(U3569)
         );
  MUX2_X1 U4610 ( .A(n4225), .B(DATAO_REG_18__SCAN_IN), .S(n3929), .Z(U3568)
         );
  MUX2_X1 U4611 ( .A(n3922), .B(DATAO_REG_16__SCAN_IN), .S(n3929), .Z(U3566)
         );
  MUX2_X1 U4612 ( .A(n3923), .B(DATAO_REG_15__SCAN_IN), .S(n3929), .Z(U3565)
         );
  MUX2_X1 U4613 ( .A(n3924), .B(DATAO_REG_14__SCAN_IN), .S(n3929), .Z(U3564)
         );
  MUX2_X1 U4614 ( .A(n3925), .B(DATAO_REG_13__SCAN_IN), .S(n3929), .Z(U3563)
         );
  MUX2_X1 U4615 ( .A(n3926), .B(DATAO_REG_12__SCAN_IN), .S(n3929), .Z(U3562)
         );
  MUX2_X1 U4616 ( .A(n3927), .B(DATAO_REG_10__SCAN_IN), .S(n3929), .Z(U3560)
         );
  MUX2_X1 U4617 ( .A(n3928), .B(DATAO_REG_9__SCAN_IN), .S(n3929), .Z(U3559) );
  MUX2_X1 U4618 ( .A(n3930), .B(DATAO_REG_8__SCAN_IN), .S(n3929), .Z(U3558) );
  MUX2_X1 U4619 ( .A(n3931), .B(DATAO_REG_7__SCAN_IN), .S(n3929), .Z(U3557) );
  MUX2_X1 U4620 ( .A(n3932), .B(DATAO_REG_6__SCAN_IN), .S(n3929), .Z(U3556) );
  MUX2_X1 U4621 ( .A(n3933), .B(DATAO_REG_5__SCAN_IN), .S(n3929), .Z(U3555) );
  MUX2_X1 U4622 ( .A(n3934), .B(DATAO_REG_4__SCAN_IN), .S(n3929), .Z(U3554) );
  MUX2_X1 U4623 ( .A(n2925), .B(DATAO_REG_3__SCAN_IN), .S(n3929), .Z(U3553) );
  MUX2_X1 U4624 ( .A(n4558), .B(DATAO_REG_2__SCAN_IN), .S(n3929), .Z(U3552) );
  MUX2_X1 U4625 ( .A(n2921), .B(DATAO_REG_1__SCAN_IN), .S(n3929), .Z(U3551) );
  OAI211_X1 U4626 ( .C1(n3937), .C2(n3936), .A(n4545), .B(n3935), .ZN(n3943)
         );
  OAI211_X1 U4627 ( .C1(n3946), .C2(n3938), .A(n4543), .B(n3951), .ZN(n3942)
         );
  AOI22_X1 U4628 ( .A1(n4535), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3941) );
  INV_X1 U4629 ( .A(n2881), .ZN(n3939) );
  NAND2_X1 U4630 ( .A1(n4509), .A2(n3939), .ZN(n3940) );
  NAND4_X1 U4631 ( .A1(n3943), .A2(n3942), .A3(n3941), .A4(n3940), .ZN(U3241)
         );
  NAND3_X1 U4632 ( .A1(n3944), .A2(n4448), .A3(n3993), .ZN(n3949) );
  OR2_X1 U4633 ( .A1(n3993), .A2(REG2_REG_0__SCAN_IN), .ZN(n3945) );
  NAND2_X1 U4634 ( .A1(n4448), .A2(n3945), .ZN(n4464) );
  AOI22_X1 U4635 ( .A1(n3947), .A2(n3946), .B1(n4464), .B2(n2157), .ZN(n3948)
         );
  NAND3_X1 U4636 ( .A1(n3949), .A2(U4043), .A3(n3948), .ZN(n4480) );
  AOI22_X1 U4637 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4535), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3962) );
  NAND3_X1 U4638 ( .A1(n3952), .A2(n3951), .A3(n3950), .ZN(n3953) );
  AND3_X1 U4639 ( .A1(n4543), .A2(n3954), .A3(n3953), .ZN(n3955) );
  AOI21_X1 U4640 ( .B1(n4509), .B2(n4461), .A(n3955), .ZN(n3961) );
  NAND3_X1 U4641 ( .A1(n3957), .A2(n3935), .A3(n3956), .ZN(n3958) );
  NAND3_X1 U4642 ( .A1(n4545), .A2(n3959), .A3(n3958), .ZN(n3960) );
  NAND4_X1 U4643 ( .A1(n4480), .A2(n3962), .A3(n3961), .A4(n3960), .ZN(U3242)
         );
  NOR2_X1 U4644 ( .A1(n3964), .A2(n3963), .ZN(n3967) );
  AOI21_X1 U4645 ( .B1(n3967), .B2(n3966), .A(n4504), .ZN(n3965) );
  OAI21_X1 U4646 ( .B1(n3967), .B2(n3966), .A(n3965), .ZN(n3976) );
  INV_X1 U4647 ( .A(n3968), .ZN(n3972) );
  INV_X1 U4648 ( .A(n3969), .ZN(n3970) );
  AOI211_X1 U4649 ( .C1(n3972), .C2(n3971), .A(n3970), .B(n4513), .ZN(n3973)
         );
  AOI211_X1 U4650 ( .C1(n4535), .C2(ADDR_REG_13__SCAN_IN), .A(n3974), .B(n3973), .ZN(n3975) );
  OAI211_X1 U4651 ( .C1(n4548), .C2(n3977), .A(n3976), .B(n3975), .ZN(U3253)
         );
  XNOR2_X1 U4652 ( .A(n3979), .B(n2049), .ZN(n3991) );
  INV_X1 U4653 ( .A(n3980), .ZN(n3981) );
  MUX2_X1 U4654 ( .A(REG2_REG_19__SCAN_IN), .B(n2644), .S(n3982), .Z(n3983) );
  XNOR2_X1 U4655 ( .A(n3984), .B(n3983), .ZN(n3989) );
  NAND2_X1 U4656 ( .A1(n4535), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3985) );
  OAI211_X1 U4657 ( .C1(n4548), .C2(n3987), .A(n3986), .B(n3985), .ZN(n3988)
         );
  AOI21_X1 U4658 ( .B1(n3989), .B2(n4543), .A(n3988), .ZN(n3990) );
  OAI21_X1 U4659 ( .B1(n3991), .B2(n4513), .A(n3990), .ZN(U3259) );
  NAND2_X1 U4660 ( .A1(n4012), .A2(n4000), .ZN(n3999) );
  XOR2_X1 U4661 ( .A(n3996), .B(n3999), .Z(n4394) );
  INV_X1 U4662 ( .A(B_REG_SCAN_IN), .ZN(n3992) );
  NOR2_X1 U4663 ( .A1(n3993), .A2(n3992), .ZN(n3994) );
  NOR2_X1 U4664 ( .A1(n4576), .A2(n3994), .ZN(n4020) );
  NAND2_X1 U4665 ( .A1(n4020), .A2(n3995), .ZN(n4003) );
  OAI21_X1 U4666 ( .B1(n4563), .B2(n3996), .A(n4003), .ZN(n4392) );
  NAND2_X1 U4667 ( .A1(n4581), .A2(n4392), .ZN(n3998) );
  NAND2_X1 U4668 ( .A1(n1998), .A2(REG2_REG_31__SCAN_IN), .ZN(n3997) );
  OAI211_X1 U4669 ( .C1(n4394), .C2(n4234), .A(n3998), .B(n3997), .ZN(U3260)
         );
  INV_X1 U4670 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4007) );
  OAI21_X1 U4671 ( .B1(n4012), .B2(n4000), .A(n3999), .ZN(n4001) );
  INV_X1 U4672 ( .A(n4001), .ZN(n4396) );
  NAND2_X1 U4673 ( .A1(n4396), .A2(n4567), .ZN(n4006) );
  NAND2_X1 U4674 ( .A1(n4273), .A2(n4002), .ZN(n4004) );
  NAND2_X1 U4675 ( .A1(n4004), .A2(n4003), .ZN(n4397) );
  NAND2_X1 U4676 ( .A1(n4581), .A2(n4397), .ZN(n4005) );
  OAI211_X1 U4677 ( .C1(n4581), .C2(n4007), .A(n4006), .B(n4005), .ZN(U3261)
         );
  NAND2_X1 U4678 ( .A1(n4009), .A2(n4008), .ZN(n4309) );
  NAND2_X1 U4679 ( .A1(n4022), .A2(n4010), .ZN(n4304) );
  NAND2_X1 U4680 ( .A1(n4309), .A2(n4304), .ZN(n4011) );
  XOR2_X1 U4681 ( .A(n4307), .B(n4011), .Z(n4029) );
  AOI22_X1 U4682 ( .A1(n4303), .A2(n4567), .B1(REG2_REG_29__SCAN_IN), .B2(
        n1998), .ZN(n4028) );
  INV_X1 U4683 ( .A(n4014), .ZN(n4016) );
  AOI22_X1 U4684 ( .A1(n4273), .A2(n4021), .B1(n4020), .B2(n4019), .ZN(n4024)
         );
  NAND2_X1 U4685 ( .A1(n4022), .A2(n4559), .ZN(n4023) );
  NOR2_X1 U4686 ( .A1(n4025), .A2(n4276), .ZN(n4026) );
  OAI21_X1 U4687 ( .B1(n4306), .B2(n4026), .A(n4581), .ZN(n4027) );
  OAI211_X1 U4688 ( .C1(n4029), .C2(n4283), .A(n4028), .B(n4027), .ZN(U3354)
         );
  NOR2_X1 U4689 ( .A1(n4030), .A2(n4040), .ZN(n4031) );
  OR2_X1 U4690 ( .A1(n4032), .A2(n4031), .ZN(n4038) );
  OAI22_X1 U4691 ( .A1(n4033), .A2(n4264), .B1(n4041), .B2(n4563), .ZN(n4034)
         );
  INV_X1 U4692 ( .A(n4034), .ZN(n4035) );
  OAI21_X1 U4693 ( .B1(n4036), .B2(n4576), .A(n4035), .ZN(n4037) );
  AOI21_X1 U4694 ( .B1(n4038), .B2(n4573), .A(n4037), .ZN(n4315) );
  XOR2_X1 U4695 ( .A(n4040), .B(n4039), .Z(n4314) );
  NAND2_X1 U4696 ( .A1(n4314), .A2(n4258), .ZN(n4048) );
  OR2_X1 U4697 ( .A1(n4059), .A2(n4041), .ZN(n4042) );
  NAND2_X1 U4698 ( .A1(n3017), .A2(n4042), .ZN(n4317) );
  INV_X1 U4699 ( .A(n4317), .ZN(n4046) );
  INV_X1 U4700 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4043) );
  OAI22_X1 U4701 ( .A1(n4044), .A2(n4276), .B1(n4043), .B2(n4581), .ZN(n4045)
         );
  AOI21_X1 U4702 ( .B1(n4046), .B2(n4567), .A(n4045), .ZN(n4047) );
  OAI211_X1 U4703 ( .C1(n4315), .C2(n1998), .A(n4048), .B(n4047), .ZN(U3263)
         );
  XOR2_X1 U4704 ( .A(n4053), .B(n4049), .Z(n4319) );
  INV_X1 U4705 ( .A(n4319), .ZN(n4067) );
  NAND2_X1 U4706 ( .A1(n4051), .A2(n4050), .ZN(n4052) );
  XOR2_X1 U4707 ( .A(n4053), .B(n4052), .Z(n4054) );
  NAND2_X1 U4708 ( .A1(n4054), .A2(n4573), .ZN(n4057) );
  AOI22_X1 U4709 ( .A1(n4092), .A2(n4559), .B1(n4055), .B2(n4273), .ZN(n4056)
         );
  OAI211_X1 U4710 ( .C1(n4058), .C2(n4576), .A(n4057), .B(n4056), .ZN(n4318)
         );
  INV_X1 U4711 ( .A(n4078), .ZN(n4062) );
  INV_X1 U4712 ( .A(n4059), .ZN(n4060) );
  OAI21_X1 U4713 ( .B1(n4062), .B2(n4061), .A(n4060), .ZN(n4406) );
  AOI22_X1 U4714 ( .A1(n4063), .A2(n4578), .B1(REG2_REG_26__SCAN_IN), .B2(
        n1998), .ZN(n4064) );
  OAI21_X1 U4715 ( .B1(n4406), .B2(n4234), .A(n4064), .ZN(n4065) );
  AOI21_X1 U4716 ( .B1(n4318), .B2(n4581), .A(n4065), .ZN(n4066) );
  OAI21_X1 U4717 ( .B1(n4067), .B2(n4283), .A(n4066), .ZN(U3264) );
  XNOR2_X1 U4718 ( .A(n4068), .B(n4071), .ZN(n4323) );
  INV_X1 U4719 ( .A(n4323), .ZN(n4085) );
  NAND2_X1 U4720 ( .A1(n4070), .A2(n4069), .ZN(n4072) );
  XNOR2_X1 U4721 ( .A(n4072), .B(n4071), .ZN(n4073) );
  NAND2_X1 U4722 ( .A1(n4073), .A2(n4573), .ZN(n4077) );
  OAI22_X1 U4723 ( .A1(n4115), .A2(n4264), .B1(n4079), .B2(n4563), .ZN(n4074)
         );
  AOI21_X1 U4724 ( .B1(n4075), .B2(n4557), .A(n4074), .ZN(n4076) );
  NAND2_X1 U4725 ( .A1(n4077), .A2(n4076), .ZN(n4322) );
  INV_X1 U4726 ( .A(n4097), .ZN(n4080) );
  OAI21_X1 U4727 ( .B1(n4080), .B2(n4079), .A(n4078), .ZN(n4410) );
  AOI22_X1 U4728 ( .A1(n4081), .A2(n4578), .B1(REG2_REG_25__SCAN_IN), .B2(
        n1998), .ZN(n4082) );
  OAI21_X1 U4729 ( .B1(n4410), .B2(n4234), .A(n4082), .ZN(n4083) );
  AOI21_X1 U4730 ( .B1(n4581), .B2(n4322), .A(n4083), .ZN(n4084) );
  OAI21_X1 U4731 ( .B1(n4085), .B2(n4283), .A(n4084), .ZN(U3265) );
  XOR2_X1 U4732 ( .A(n4089), .B(n4086), .Z(n4327) );
  INV_X1 U4733 ( .A(n4327), .ZN(n4102) );
  NAND2_X1 U4734 ( .A1(n4088), .A2(n4087), .ZN(n4090) );
  XNOR2_X1 U4735 ( .A(n4090), .B(n4089), .ZN(n4094) );
  OAI22_X1 U4736 ( .A1(n4131), .A2(n4264), .B1(n4098), .B2(n4563), .ZN(n4091)
         );
  AOI21_X1 U4737 ( .B1(n4557), .B2(n4092), .A(n4091), .ZN(n4093) );
  OAI21_X1 U4738 ( .B1(n4094), .B2(n4288), .A(n4093), .ZN(n4326) );
  OAI22_X1 U4739 ( .A1(n4095), .A2(n4276), .B1(n3589), .B2(n4581), .ZN(n4100)
         );
  OAI21_X1 U4740 ( .B1(n4096), .B2(n4098), .A(n4097), .ZN(n4414) );
  NOR2_X1 U4741 ( .A1(n4414), .A2(n4234), .ZN(n4099) );
  AOI211_X1 U4742 ( .C1(n4581), .C2(n4326), .A(n4100), .B(n4099), .ZN(n4101)
         );
  OAI21_X1 U4743 ( .B1(n4102), .B2(n4283), .A(n4101), .ZN(U3266) );
  XNOR2_X1 U4744 ( .A(n4103), .B(n4113), .ZN(n4331) );
  INV_X1 U4745 ( .A(n4331), .ZN(n4126) );
  NAND2_X1 U4746 ( .A1(n4243), .A2(n4104), .ZN(n4222) );
  OR2_X2 U4747 ( .A1(n4222), .A2(n4105), .ZN(n4202) );
  INV_X1 U4748 ( .A(n4106), .ZN(n4107) );
  OAI21_X1 U4749 ( .B1(n4202), .B2(n4161), .A(n4107), .ZN(n4109) );
  NAND2_X1 U4750 ( .A1(n4109), .A2(n4108), .ZN(n4148) );
  OAI21_X1 U4751 ( .B1(n4148), .B2(n4147), .A(n4110), .ZN(n4127) );
  INV_X1 U4752 ( .A(n4111), .ZN(n4112) );
  AOI21_X1 U4753 ( .B1(n4127), .B2(n4134), .A(n4112), .ZN(n4114) );
  XNOR2_X1 U4754 ( .A(n4114), .B(n4113), .ZN(n4118) );
  OAI22_X1 U4755 ( .A1(n4115), .A2(n4576), .B1(n4563), .B2(n4120), .ZN(n4116)
         );
  AOI21_X1 U4756 ( .B1(n4559), .B2(n4149), .A(n4116), .ZN(n4117) );
  OAI21_X1 U4757 ( .B1(n4118), .B2(n4288), .A(n4117), .ZN(n4330) );
  INV_X1 U4758 ( .A(n4119), .ZN(n4121) );
  OAI21_X1 U4759 ( .B1(n4121), .B2(n4120), .A(n2091), .ZN(n4418) );
  AOI22_X1 U4760 ( .A1(n4122), .A2(n4578), .B1(REG2_REG_23__SCAN_IN), .B2(
        n1998), .ZN(n4123) );
  OAI21_X1 U4761 ( .B1(n4418), .B2(n4234), .A(n4123), .ZN(n4124) );
  AOI21_X1 U4762 ( .B1(n4330), .B2(n4581), .A(n4124), .ZN(n4125) );
  OAI21_X1 U4763 ( .B1(n4126), .B2(n4283), .A(n4125), .ZN(U3267) );
  XNOR2_X1 U4764 ( .A(n4127), .B(n4134), .ZN(n4133) );
  AOI22_X1 U4765 ( .A1(n4129), .A2(n4559), .B1(n4128), .B2(n4273), .ZN(n4130)
         );
  OAI21_X1 U4766 ( .B1(n4131), .B2(n4576), .A(n4130), .ZN(n4132) );
  AOI21_X1 U4767 ( .B1(n4133), .B2(n4573), .A(n4132), .ZN(n4336) );
  OAI21_X1 U4768 ( .B1(n4136), .B2(n2957), .A(n4135), .ZN(n4337) );
  AOI22_X1 U4769 ( .A1(n4137), .A2(n4578), .B1(n1998), .B2(
        REG2_REG_22__SCAN_IN), .ZN(n4141) );
  OR2_X1 U4770 ( .A1(n4138), .A2(n4139), .ZN(n4334) );
  NAND3_X1 U4771 ( .A1(n4119), .A2(n4334), .A3(n4567), .ZN(n4140) );
  OAI211_X1 U4772 ( .C1(n4337), .C2(n4283), .A(n4141), .B(n4140), .ZN(n4142)
         );
  INV_X1 U4773 ( .A(n4142), .ZN(n4143) );
  OAI21_X1 U4774 ( .B1(n1998), .B2(n4336), .A(n4143), .ZN(U3268) );
  XNOR2_X1 U4775 ( .A(n4144), .B(n4147), .ZN(n4341) );
  AOI21_X1 U4776 ( .B1(n4150), .B2(n4175), .A(n4138), .ZN(n4338) );
  INV_X1 U4777 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4145) );
  OAI22_X1 U4778 ( .A1(n4146), .A2(n4276), .B1(n4581), .B2(n4145), .ZN(n4156)
         );
  XNOR2_X1 U4779 ( .A(n4148), .B(n4147), .ZN(n4154) );
  NAND2_X1 U4780 ( .A1(n4149), .A2(n4557), .ZN(n4152) );
  AOI22_X1 U4781 ( .A1(n4188), .A2(n4559), .B1(n4150), .B2(n4273), .ZN(n4151)
         );
  NAND2_X1 U4782 ( .A1(n4152), .A2(n4151), .ZN(n4153) );
  AOI21_X1 U4783 ( .B1(n4154), .B2(n4573), .A(n4153), .ZN(n4340) );
  NOR2_X1 U4784 ( .A1(n4340), .A2(n1998), .ZN(n4155) );
  AOI211_X1 U4785 ( .C1(n4338), .C2(n4567), .A(n4156), .B(n4155), .ZN(n4157)
         );
  OAI21_X1 U4786 ( .B1(n4341), .B2(n4283), .A(n4157), .ZN(U3269) );
  XNOR2_X1 U4787 ( .A(n4158), .B(n4162), .ZN(n4173) );
  OAI21_X1 U4788 ( .B1(n4184), .B2(n4161), .A(n4160), .ZN(n4164) );
  INV_X1 U4789 ( .A(n4162), .ZN(n4163) );
  XNOR2_X1 U4790 ( .A(n4164), .B(n4163), .ZN(n4170) );
  AOI22_X1 U4791 ( .A1(n4166), .A2(n4559), .B1(n4165), .B2(n4273), .ZN(n4167)
         );
  OAI21_X1 U4792 ( .B1(n4168), .B2(n4576), .A(n4167), .ZN(n4169) );
  AOI21_X1 U4793 ( .B1(n4170), .B2(n4573), .A(n4169), .ZN(n4171) );
  OAI21_X1 U4794 ( .B1(n4173), .B2(n4172), .A(n4171), .ZN(n4342) );
  INV_X1 U4795 ( .A(n4342), .ZN(n4181) );
  INV_X1 U4796 ( .A(n4173), .ZN(n4343) );
  OAI21_X1 U4797 ( .B1(n4174), .B2(n4176), .A(n4175), .ZN(n4424) );
  AOI22_X1 U4798 ( .A1(n1998), .A2(REG2_REG_20__SCAN_IN), .B1(n4177), .B2(
        n4578), .ZN(n4178) );
  OAI21_X1 U4799 ( .B1(n4424), .B2(n4234), .A(n4178), .ZN(n4179) );
  AOI21_X1 U4800 ( .B1(n4343), .B2(n4579), .A(n4179), .ZN(n4180) );
  OAI21_X1 U4801 ( .B1(n4181), .B2(n1998), .A(n4180), .ZN(U3270) );
  INV_X1 U4802 ( .A(n4182), .ZN(n4183) );
  NOR2_X1 U4803 ( .A1(n4184), .A2(n4183), .ZN(n4185) );
  XNOR2_X1 U4804 ( .A(n4185), .B(n4191), .ZN(n4190) );
  OAI22_X1 U4805 ( .A1(n4186), .A2(n4264), .B1(n4563), .B2(n4193), .ZN(n4187)
         );
  AOI21_X1 U4806 ( .B1(n4188), .B2(n4557), .A(n4187), .ZN(n4189) );
  OAI21_X1 U4807 ( .B1(n4190), .B2(n4288), .A(n4189), .ZN(n4346) );
  INV_X1 U4808 ( .A(n4346), .ZN(n4200) );
  XNOR2_X1 U4809 ( .A(n4192), .B(n4191), .ZN(n4347) );
  NOR2_X1 U4810 ( .A1(n4194), .A2(n4193), .ZN(n4195) );
  OR2_X1 U4811 ( .A1(n4174), .A2(n4195), .ZN(n4428) );
  AOI22_X1 U4812 ( .A1(n1998), .A2(REG2_REG_19__SCAN_IN), .B1(n4196), .B2(
        n4578), .ZN(n4197) );
  OAI21_X1 U4813 ( .B1(n4428), .B2(n4234), .A(n4197), .ZN(n4198) );
  AOI21_X1 U4814 ( .B1(n4347), .B2(n4258), .A(n4198), .ZN(n4199) );
  OAI21_X1 U4815 ( .B1(n1998), .B2(n4200), .A(n4199), .ZN(U3271) );
  NAND2_X1 U4816 ( .A1(n4202), .A2(n4201), .ZN(n4203) );
  XOR2_X1 U4817 ( .A(n4203), .B(n4211), .Z(n4209) );
  AOI22_X1 U4818 ( .A1(n4205), .A2(n4559), .B1(n4204), .B2(n4273), .ZN(n4206)
         );
  OAI21_X1 U4819 ( .B1(n4207), .B2(n4576), .A(n4206), .ZN(n4208) );
  AOI21_X1 U4820 ( .B1(n4209), .B2(n4573), .A(n4208), .ZN(n4352) );
  OAI21_X1 U4821 ( .B1(n4212), .B2(n4211), .A(n4210), .ZN(n4350) );
  XNOR2_X1 U4822 ( .A(n4233), .B(n4213), .ZN(n4214) );
  NAND2_X1 U4823 ( .A1(n4214), .A2(n3020), .ZN(n4351) );
  INV_X1 U4824 ( .A(n4215), .ZN(n4216) );
  NOR2_X1 U4825 ( .A1(n4351), .A2(n4216), .ZN(n4220) );
  INV_X1 U4826 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4218) );
  OAI22_X1 U4827 ( .A1(n4581), .A2(n4218), .B1(n4217), .B2(n4276), .ZN(n4219)
         );
  AOI211_X1 U4828 ( .C1(n4350), .C2(n4258), .A(n4220), .B(n4219), .ZN(n4221)
         );
  OAI21_X1 U4829 ( .B1(n1998), .B2(n4352), .A(n4221), .ZN(U3272) );
  XOR2_X1 U4830 ( .A(n4228), .B(n4222), .Z(n4227) );
  OAI22_X1 U4831 ( .A1(n4266), .A2(n4264), .B1(n4563), .B2(n4223), .ZN(n4224)
         );
  AOI21_X1 U4832 ( .B1(n4225), .B2(n4557), .A(n4224), .ZN(n4226) );
  OAI21_X1 U4833 ( .B1(n4227), .B2(n4288), .A(n4226), .ZN(n4354) );
  INV_X1 U4834 ( .A(n4354), .ZN(n4240) );
  XOR2_X1 U4835 ( .A(n4229), .B(n4228), .Z(n4355) );
  NAND2_X1 U4836 ( .A1(n4230), .A2(n4231), .ZN(n4232) );
  NAND2_X1 U4837 ( .A1(n4233), .A2(n4232), .ZN(n4433) );
  NOR2_X1 U4838 ( .A1(n4433), .A2(n4234), .ZN(n4238) );
  OAI22_X1 U4839 ( .A1(n4581), .A2(n4236), .B1(n4235), .B2(n4276), .ZN(n4237)
         );
  AOI211_X1 U4840 ( .C1(n4355), .C2(n4258), .A(n4238), .B(n4237), .ZN(n4239)
         );
  OAI21_X1 U4841 ( .B1(n1998), .B2(n4240), .A(n4239), .ZN(U3273) );
  OAI22_X1 U4842 ( .A1(n4242), .A2(n4576), .B1(n4241), .B2(n4264), .ZN(n4246)
         );
  INV_X1 U4843 ( .A(n4243), .ZN(n4244) );
  AOI211_X1 U4844 ( .C1(n2022), .C2(n4256), .A(n4288), .B(n4244), .ZN(n4245)
         );
  AOI211_X1 U4845 ( .C1(n4273), .C2(n4247), .A(n4246), .B(n4245), .ZN(n4360)
         );
  OAI21_X1 U4846 ( .B1(n4274), .B2(n4248), .A(n4230), .ZN(n4361) );
  INV_X1 U4847 ( .A(n4361), .ZN(n4252) );
  INV_X1 U4848 ( .A(n4249), .ZN(n4250) );
  OAI22_X1 U4849 ( .A1(n4581), .A2(n4528), .B1(n4250), .B2(n4276), .ZN(n4251)
         );
  AOI21_X1 U4850 ( .B1(n4252), .B2(n4567), .A(n4251), .ZN(n4260) );
  INV_X1 U4851 ( .A(n4253), .ZN(n4255) );
  OAI21_X1 U4852 ( .B1(n4262), .B2(n4255), .A(n4254), .ZN(n4257) );
  XNOR2_X1 U4853 ( .A(n4257), .B(n4256), .ZN(n4358) );
  NAND2_X1 U4854 ( .A1(n4358), .A2(n4258), .ZN(n4259) );
  OAI211_X1 U4855 ( .C1(n4360), .C2(n1998), .A(n4260), .B(n4259), .ZN(U3274)
         );
  NAND2_X1 U4856 ( .A1(n4262), .A2(n4261), .ZN(n4263) );
  XNOR2_X1 U4857 ( .A(n4263), .B(n2114), .ZN(n4366) );
  OAI22_X1 U4858 ( .A1(n4266), .A2(n4576), .B1(n4265), .B2(n4264), .ZN(n4272)
         );
  INV_X1 U4859 ( .A(n4267), .ZN(n4268) );
  AOI211_X1 U4860 ( .C1(n4270), .C2(n4269), .A(n4288), .B(n4268), .ZN(n4271)
         );
  AOI211_X1 U4861 ( .C1(n4273), .C2(n4275), .A(n4272), .B(n4271), .ZN(n4365)
         );
  INV_X1 U4862 ( .A(n4365), .ZN(n4281) );
  INV_X1 U4863 ( .A(n4274), .ZN(n4363) );
  NAND2_X1 U4864 ( .A1(n4367), .A2(n4275), .ZN(n4362) );
  AND3_X1 U4865 ( .A1(n4363), .A2(n4567), .A3(n4362), .ZN(n4280) );
  OAI22_X1 U4866 ( .A1(n4581), .A2(n4278), .B1(n4277), .B2(n4276), .ZN(n4279)
         );
  AOI211_X1 U4867 ( .C1(n4281), .C2(n4581), .A(n4280), .B(n4279), .ZN(n4282)
         );
  OAI21_X1 U4868 ( .B1(n4366), .B2(n4283), .A(n4282), .ZN(U3275) );
  OAI21_X1 U4869 ( .B1(n4284), .B2(n2971), .A(n4285), .ZN(n4617) );
  AOI22_X1 U4870 ( .A1(n4559), .A2(n2921), .B1(n2925), .B2(n4557), .ZN(n4286)
         );
  OAI21_X1 U4871 ( .B1(n4563), .B2(n4287), .A(n4286), .ZN(n4291) );
  NAND3_X1 U4872 ( .A1(n4553), .A2(n2971), .A3(n2970), .ZN(n4289) );
  AOI21_X1 U4873 ( .B1(n3298), .B2(n4289), .A(n4288), .ZN(n4290) );
  AOI211_X1 U4874 ( .C1(n4574), .C2(n4617), .A(n4291), .B(n4290), .ZN(n4614)
         );
  MUX2_X1 U4875 ( .A(n4292), .B(n4614), .S(n4581), .Z(n4296) );
  AOI22_X1 U4876 ( .A1(n4579), .A2(n4617), .B1(REG3_REG_2__SCAN_IN), .B2(n4578), .ZN(n4295) );
  INV_X1 U4877 ( .A(n3309), .ZN(n4613) );
  NAND2_X1 U4878 ( .A1(n4565), .A2(n4293), .ZN(n4612) );
  NAND3_X1 U4879 ( .A1(n4567), .A2(n4613), .A3(n4612), .ZN(n4294) );
  NAND3_X1 U4880 ( .A1(n4296), .A2(n4295), .A3(n4294), .ZN(U3288) );
  NAND2_X1 U4881 ( .A1(n4658), .A2(n4392), .ZN(n4298) );
  NAND2_X1 U4882 ( .A1(n4656), .A2(REG1_REG_31__SCAN_IN), .ZN(n4297) );
  OAI211_X1 U4883 ( .C1(n4394), .C2(n4379), .A(n4298), .B(n4297), .ZN(U3549)
         );
  NAND2_X1 U4884 ( .A1(n4396), .A2(n4299), .ZN(n4301) );
  NAND2_X1 U4885 ( .A1(n4658), .A2(n4397), .ZN(n4300) );
  OAI211_X1 U4886 ( .C1(n4658), .C2(n4302), .A(n4301), .B(n4300), .ZN(U3548)
         );
  NAND4_X1 U4887 ( .A1(n4309), .A2(n4644), .A3(n4018), .A4(n4304), .ZN(n4312)
         );
  NOR3_X1 U4888 ( .A1(n4018), .A2(n4304), .A3(n4629), .ZN(n4305) );
  NAND2_X1 U4889 ( .A1(n4307), .A2(n4644), .ZN(n4308) );
  NAND4_X1 U4890 ( .A1(n4313), .A2(n4312), .A3(n4311), .A4(n4310), .ZN(n4401)
         );
  MUX2_X1 U4891 ( .A(REG1_REG_29__SCAN_IN), .B(n4401), .S(n4658), .Z(U3547) );
  NAND2_X1 U4892 ( .A1(n4314), .A2(n4644), .ZN(n4316) );
  OAI211_X1 U4893 ( .C1(n4635), .C2(n4317), .A(n4316), .B(n4315), .ZN(n4402)
         );
  MUX2_X1 U4894 ( .A(REG1_REG_27__SCAN_IN), .B(n4402), .S(n4658), .Z(U3545) );
  INV_X1 U4895 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4320) );
  AOI21_X1 U4896 ( .B1(n4319), .B2(n4644), .A(n4318), .ZN(n4403) );
  MUX2_X1 U4897 ( .A(n4320), .B(n4403), .S(n4658), .Z(n4321) );
  OAI21_X1 U4898 ( .B1(n4379), .B2(n4406), .A(n4321), .ZN(U3544) );
  INV_X1 U4899 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4324) );
  AOI21_X1 U4900 ( .B1(n4323), .B2(n4644), .A(n4322), .ZN(n4407) );
  MUX2_X1 U4901 ( .A(n4324), .B(n4407), .S(n4658), .Z(n4325) );
  OAI21_X1 U4902 ( .B1(n4379), .B2(n4410), .A(n4325), .ZN(U3543) );
  AOI21_X1 U4903 ( .B1(n4327), .B2(n4644), .A(n4326), .ZN(n4411) );
  MUX2_X1 U4904 ( .A(n4328), .B(n4411), .S(n4658), .Z(n4329) );
  OAI21_X1 U4905 ( .B1(n4379), .B2(n4414), .A(n4329), .ZN(U3542) );
  INV_X1 U4906 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4332) );
  AOI21_X1 U4907 ( .B1(n4331), .B2(n4644), .A(n4330), .ZN(n4415) );
  MUX2_X1 U4908 ( .A(n4332), .B(n4415), .S(n4658), .Z(n4333) );
  OAI21_X1 U4909 ( .B1(n4379), .B2(n4418), .A(n4333), .ZN(U3541) );
  NAND3_X1 U4910 ( .A1(n4119), .A2(n4334), .A3(n3020), .ZN(n4335) );
  OAI211_X1 U4911 ( .C1(n4337), .C2(n4629), .A(n4336), .B(n4335), .ZN(n4419)
         );
  MUX2_X1 U4912 ( .A(REG1_REG_22__SCAN_IN), .B(n4419), .S(n4658), .Z(U3540) );
  NAND2_X1 U4913 ( .A1(n4338), .A2(n3020), .ZN(n4339) );
  OAI211_X1 U4914 ( .C1(n4341), .C2(n4629), .A(n4340), .B(n4339), .ZN(n4420)
         );
  MUX2_X1 U4915 ( .A(REG1_REG_21__SCAN_IN), .B(n4420), .S(n4658), .Z(U3539) );
  AOI21_X1 U4916 ( .B1(n4641), .B2(n4343), .A(n4342), .ZN(n4421) );
  MUX2_X1 U4917 ( .A(n4344), .B(n4421), .S(n4658), .Z(n4345) );
  OAI21_X1 U4918 ( .B1(n4379), .B2(n4424), .A(n4345), .ZN(U3538) );
  INV_X1 U4919 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4348) );
  AOI21_X1 U4920 ( .B1(n4347), .B2(n4644), .A(n4346), .ZN(n4425) );
  MUX2_X1 U4921 ( .A(n4348), .B(n4425), .S(n4658), .Z(n4349) );
  OAI21_X1 U4922 ( .B1(n4379), .B2(n4428), .A(n4349), .ZN(U3537) );
  INV_X1 U4923 ( .A(n4350), .ZN(n4353) );
  OAI211_X1 U4924 ( .C1(n4353), .C2(n4629), .A(n4352), .B(n4351), .ZN(n4429)
         );
  MUX2_X1 U4925 ( .A(REG1_REG_18__SCAN_IN), .B(n4429), .S(n4658), .Z(U3536) );
  AOI21_X1 U4926 ( .B1(n4355), .B2(n4644), .A(n4354), .ZN(n4430) );
  MUX2_X1 U4927 ( .A(n4356), .B(n4430), .S(n4658), .Z(n4357) );
  OAI21_X1 U4928 ( .B1(n4379), .B2(n4433), .A(n4357), .ZN(U3535) );
  NAND2_X1 U4929 ( .A1(n4358), .A2(n4644), .ZN(n4359) );
  OAI211_X1 U4930 ( .C1(n4635), .C2(n4361), .A(n4360), .B(n4359), .ZN(n4434)
         );
  MUX2_X1 U4931 ( .A(REG1_REG_16__SCAN_IN), .B(n4434), .S(n4658), .Z(U3534) );
  NAND3_X1 U4932 ( .A1(n4363), .A2(n3020), .A3(n4362), .ZN(n4364) );
  OAI211_X1 U4933 ( .C1(n4366), .C2(n4629), .A(n4365), .B(n4364), .ZN(n4435)
         );
  MUX2_X1 U4934 ( .A(REG1_REG_15__SCAN_IN), .B(n4435), .S(n4658), .Z(U3533) );
  NAND3_X1 U4935 ( .A1(n4368), .A2(n3020), .A3(n4367), .ZN(n4369) );
  OAI211_X1 U4936 ( .C1(n4371), .C2(n4388), .A(n4370), .B(n4369), .ZN(n4436)
         );
  MUX2_X1 U4937 ( .A(REG1_REG_14__SCAN_IN), .B(n4436), .S(n4658), .Z(U3532) );
  AOI21_X1 U4938 ( .B1(n4641), .B2(n4373), .A(n4372), .ZN(n4437) );
  MUX2_X1 U4939 ( .A(n4374), .B(n4437), .S(n4658), .Z(n4375) );
  OAI21_X1 U4940 ( .B1(n4440), .B2(n4379), .A(n4375), .ZN(U3531) );
  AOI21_X1 U4941 ( .B1(n4377), .B2(n4644), .A(n4376), .ZN(n4441) );
  MUX2_X1 U4942 ( .A(n4493), .B(n4441), .S(n4658), .Z(n4378) );
  OAI21_X1 U4943 ( .B1(n4379), .B2(n4445), .A(n4378), .ZN(U3530) );
  NAND2_X1 U4944 ( .A1(n4380), .A2(n4641), .ZN(n4381) );
  OAI211_X1 U4945 ( .C1(n4635), .C2(n4383), .A(n4382), .B(n4381), .ZN(n4446)
         );
  MUX2_X1 U4946 ( .A(REG1_REG_11__SCAN_IN), .B(n4446), .S(n4658), .Z(U3529) );
  NAND3_X1 U4947 ( .A1(n4385), .A2(n3020), .A3(n4384), .ZN(n4386) );
  OAI211_X1 U4948 ( .C1(n4389), .C2(n4388), .A(n4387), .B(n4386), .ZN(n4447)
         );
  MUX2_X1 U4949 ( .A(REG1_REG_8__SCAN_IN), .B(n4447), .S(n4658), .Z(U3526) );
  NOR2_X1 U4950 ( .A1(n4647), .A2(n4390), .ZN(n4391) );
  AOI21_X1 U4951 ( .B1(n4647), .B2(n4392), .A(n4391), .ZN(n4393) );
  OAI21_X1 U4952 ( .B1(n4394), .B2(n4444), .A(n4393), .ZN(U3517) );
  NAND2_X1 U4953 ( .A1(n4396), .A2(n4395), .ZN(n4399) );
  NAND2_X1 U4954 ( .A1(n4647), .A2(n4397), .ZN(n4398) );
  OAI211_X1 U4955 ( .C1(n4647), .C2(n4400), .A(n4399), .B(n4398), .ZN(U3516)
         );
  MUX2_X1 U4956 ( .A(REG0_REG_29__SCAN_IN), .B(n4401), .S(n4647), .Z(U3515) );
  MUX2_X1 U4957 ( .A(REG0_REG_27__SCAN_IN), .B(n4402), .S(n4647), .Z(U3513) );
  INV_X1 U4958 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4404) );
  MUX2_X1 U4959 ( .A(n4404), .B(n4403), .S(n4647), .Z(n4405) );
  OAI21_X1 U4960 ( .B1(n4406), .B2(n4444), .A(n4405), .ZN(U3512) );
  INV_X1 U4961 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4408) );
  MUX2_X1 U4962 ( .A(n4408), .B(n4407), .S(n4647), .Z(n4409) );
  OAI21_X1 U4963 ( .B1(n4410), .B2(n4444), .A(n4409), .ZN(U3511) );
  INV_X1 U4964 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4412) );
  MUX2_X1 U4965 ( .A(n4412), .B(n4411), .S(n4647), .Z(n4413) );
  OAI21_X1 U4966 ( .B1(n4414), .B2(n4444), .A(n4413), .ZN(U3510) );
  INV_X1 U4967 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4416) );
  MUX2_X1 U4968 ( .A(n4416), .B(n4415), .S(n4647), .Z(n4417) );
  OAI21_X1 U4969 ( .B1(n4418), .B2(n4444), .A(n4417), .ZN(U3509) );
  MUX2_X1 U4970 ( .A(REG0_REG_22__SCAN_IN), .B(n4419), .S(n4647), .Z(U3508) );
  MUX2_X1 U4971 ( .A(REG0_REG_21__SCAN_IN), .B(n4420), .S(n4647), .Z(U3507) );
  INV_X1 U4972 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4422) );
  MUX2_X1 U4973 ( .A(n4422), .B(n4421), .S(n4647), .Z(n4423) );
  OAI21_X1 U4974 ( .B1(n4424), .B2(n4444), .A(n4423), .ZN(U3506) );
  INV_X1 U4975 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4426) );
  MUX2_X1 U4976 ( .A(n4426), .B(n4425), .S(n4647), .Z(n4427) );
  OAI21_X1 U4977 ( .B1(n4428), .B2(n4444), .A(n4427), .ZN(U3505) );
  MUX2_X1 U4978 ( .A(REG0_REG_18__SCAN_IN), .B(n4429), .S(n4647), .Z(U3503) );
  INV_X1 U4979 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4431) );
  MUX2_X1 U4980 ( .A(n4431), .B(n4430), .S(n4647), .Z(n4432) );
  OAI21_X1 U4981 ( .B1(n4433), .B2(n4444), .A(n4432), .ZN(U3501) );
  MUX2_X1 U4982 ( .A(REG0_REG_16__SCAN_IN), .B(n4434), .S(n4647), .Z(U3499) );
  MUX2_X1 U4983 ( .A(REG0_REG_15__SCAN_IN), .B(n4435), .S(n4647), .Z(U3497) );
  MUX2_X1 U4984 ( .A(REG0_REG_14__SCAN_IN), .B(n4436), .S(n4647), .Z(U3495) );
  MUX2_X1 U4985 ( .A(n4438), .B(n4437), .S(n4647), .Z(n4439) );
  OAI21_X1 U4986 ( .B1(n4440), .B2(n4444), .A(n4439), .ZN(U3493) );
  MUX2_X1 U4987 ( .A(n4442), .B(n4441), .S(n4647), .Z(n4443) );
  OAI21_X1 U4988 ( .B1(n4445), .B2(n4444), .A(n4443), .ZN(U3491) );
  MUX2_X1 U4989 ( .A(REG0_REG_11__SCAN_IN), .B(n4446), .S(n4647), .Z(U3489) );
  MUX2_X1 U4990 ( .A(REG0_REG_8__SCAN_IN), .B(n4447), .S(n4647), .Z(U3483) );
  MUX2_X1 U4991 ( .A(DATAI_30_), .B(n2323), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4992 ( .A(n4448), .B(DATAI_28_), .S(U3149), .Z(U3324) );
  MUX2_X1 U4993 ( .A(DATAI_27_), .B(n4463), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U4994 ( .A(n4449), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4995 ( .A(DATAI_25_), .B(n4450), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U4996 ( .A(DATAI_24_), .B(n2775), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U4997 ( .A(DATAI_22_), .B(n4451), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4998 ( .A(n4452), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U4999 ( .A(DATAI_20_), .B(n4453), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5000 ( .A(n4454), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U5001 ( .A(n4455), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  INV_X1 U5002 ( .A(n4456), .ZN(n4457) );
  MUX2_X1 U5003 ( .A(DATAI_8_), .B(n4457), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5004 ( .A(n4458), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5005 ( .A(n4459), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5006 ( .A(DATAI_4_), .B(n4474), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5007 ( .A(n4460), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5008 ( .A(n4461), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  INV_X1 U5009 ( .A(n4464), .ZN(n4462) );
  OAI211_X1 U5010 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4463), .A(n4465), .B(n4462), 
        .ZN(n4468) );
  AOI22_X1 U5011 ( .A1(n4465), .A2(n4464), .B1(n4545), .B2(n2350), .ZN(n4467)
         );
  AOI22_X1 U5012 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4535), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4466) );
  OAI221_X1 U5013 ( .B1(IR_REG_0__SCAN_IN), .B2(n4468), .C1(n2157), .C2(n4467), 
        .A(n4466), .ZN(U3240) );
  XNOR2_X1 U5014 ( .A(n4469), .B(n2398), .ZN(n4470) );
  NAND2_X1 U5015 ( .A1(n4543), .A2(n4470), .ZN(n4479) );
  XNOR2_X1 U5016 ( .A(n4472), .B(n4471), .ZN(n4473) );
  NAND2_X1 U5017 ( .A1(n4545), .A2(n4473), .ZN(n4478) );
  NAND2_X1 U5018 ( .A1(n4509), .A2(n4474), .ZN(n4477) );
  AOI21_X1 U5019 ( .B1(n4535), .B2(ADDR_REG_4__SCAN_IN), .A(n4475), .ZN(n4476)
         );
  AND4_X1 U5020 ( .A1(n4479), .A2(n4478), .A3(n4477), .A4(n4476), .ZN(n4481)
         );
  NAND2_X1 U5021 ( .A1(n4481), .A2(n4480), .ZN(U3244) );
  AOI211_X1 U5022 ( .C1(n4484), .C2(n4483), .A(n4482), .B(n4513), .ZN(n4486)
         );
  AOI211_X1 U5023 ( .C1(n4535), .C2(ADDR_REG_10__SCAN_IN), .A(n4486), .B(n4485), .ZN(n4490) );
  OAI211_X1 U5024 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4488), .A(n4543), .B(n4487), .ZN(n4489) );
  OAI211_X1 U5025 ( .C1(n4548), .C2(n4604), .A(n4490), .B(n4489), .ZN(U3250)
         );
  AOI211_X1 U5026 ( .C1(n4493), .C2(n4492), .A(n4491), .B(n4513), .ZN(n4495)
         );
  AOI211_X1 U5027 ( .C1(n4535), .C2(ADDR_REG_12__SCAN_IN), .A(n4495), .B(n4494), .ZN(n4499) );
  OAI211_X1 U5028 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4497), .A(n4543), .B(n4496), .ZN(n4498) );
  OAI211_X1 U5029 ( .C1(n4548), .C2(n4500), .A(n4499), .B(n4498), .ZN(U3252)
         );
  NAND2_X1 U5030 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4535), .ZN(n4512) );
  AOI211_X1 U5031 ( .C1(n4503), .C2(n4502), .A(n4501), .B(n4513), .ZN(n4508)
         );
  AOI211_X1 U5032 ( .C1(n3385), .C2(n4506), .A(n4505), .B(n4504), .ZN(n4507)
         );
  AOI211_X1 U5033 ( .C1(n4509), .C2(n4600), .A(n4508), .B(n4507), .ZN(n4511)
         );
  NAND3_X1 U5034 ( .A1(n4512), .A2(n4511), .A3(n4510), .ZN(U3254) );
  AOI211_X1 U5035 ( .C1(n2020), .C2(n4515), .A(n4514), .B(n4513), .ZN(n4516)
         );
  AOI211_X1 U5036 ( .C1(n4535), .C2(ADDR_REG_15__SCAN_IN), .A(n4517), .B(n4516), .ZN(n4522) );
  AOI21_X1 U5037 ( .B1(n4519), .B2(n2019), .A(n4518), .ZN(n4520) );
  NAND2_X1 U5038 ( .A1(n4543), .A2(n4520), .ZN(n4521) );
  OAI211_X1 U5039 ( .C1(n4548), .C2(n4599), .A(n4522), .B(n4521), .ZN(U3255)
         );
  AOI21_X1 U5040 ( .B1(n4535), .B2(ADDR_REG_16__SCAN_IN), .A(n4523), .ZN(n4533) );
  OAI21_X1 U5041 ( .B1(n4526), .B2(n4525), .A(n4524), .ZN(n4531) );
  OAI21_X1 U5042 ( .B1(n4529), .B2(n4528), .A(n4527), .ZN(n4530) );
  AOI22_X1 U5043 ( .A1(n4545), .A2(n4531), .B1(n4543), .B2(n4530), .ZN(n4532)
         );
  OAI211_X1 U5044 ( .C1(n4597), .C2(n4548), .A(n4533), .B(n4532), .ZN(U3256)
         );
  AOI21_X1 U5045 ( .B1(n4535), .B2(ADDR_REG_17__SCAN_IN), .A(n4534), .ZN(n4547) );
  OAI21_X1 U5046 ( .B1(n4538), .B2(n4537), .A(n4536), .ZN(n4544) );
  OAI21_X1 U5047 ( .B1(n4541), .B2(n4540), .A(n4539), .ZN(n4542) );
  AOI22_X1 U5048 ( .A1(n4545), .A2(n4544), .B1(n4543), .B2(n4542), .ZN(n4546)
         );
  OAI211_X1 U5049 ( .C1(n4549), .C2(n4548), .A(n4547), .B(n4546), .ZN(U3257)
         );
  INV_X1 U5050 ( .A(n4552), .ZN(n4609) );
  OAI21_X1 U5051 ( .B1(n4555), .B2(n4554), .A(n4553), .ZN(n4556) );
  NAND2_X1 U5052 ( .A1(n4556), .A2(n4573), .ZN(n4561) );
  AOI22_X1 U5053 ( .A1(n4559), .A2(n2969), .B1(n4558), .B2(n4557), .ZN(n4560)
         );
  OAI211_X1 U5054 ( .C1(n4563), .C2(n4562), .A(n4561), .B(n4560), .ZN(n4564)
         );
  AOI21_X1 U5055 ( .B1(n4574), .B2(n4609), .A(n4564), .ZN(n4611) );
  AOI22_X1 U5056 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1998), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4578), .ZN(n4569) );
  INV_X1 U5057 ( .A(n4565), .ZN(n4566) );
  AOI21_X1 U5058 ( .B1(n4571), .B2(n2336), .A(n4566), .ZN(n4608) );
  AOI22_X1 U5059 ( .A1(n4567), .A2(n4608), .B1(n4579), .B2(n4609), .ZN(n4568)
         );
  OAI211_X1 U5060 ( .C1(n1998), .C2(n4611), .A(n4569), .B(n4568), .ZN(U3289)
         );
  AND2_X1 U5061 ( .A1(n4571), .A2(n4570), .ZN(n4606) );
  INV_X1 U5062 ( .A(n4572), .ZN(n4577) );
  OAI21_X1 U5063 ( .B1(n4574), .B2(n4573), .A(n4607), .ZN(n4575) );
  OAI21_X1 U5064 ( .B1(n2920), .B2(n4576), .A(n4575), .ZN(n4605) );
  AOI21_X1 U5065 ( .B1(n4606), .B2(n4577), .A(n4605), .ZN(n4582) );
  AOI22_X1 U5066 ( .A1(n4579), .A2(n4607), .B1(REG3_REG_0__SCAN_IN), .B2(n4578), .ZN(n4580) );
  OAI221_X1 U5067 ( .B1(n1998), .B2(n4582), .C1(n4581), .C2(n2340), .A(n4580), 
        .ZN(U3290) );
  AND2_X1 U5068 ( .A1(D_REG_31__SCAN_IN), .A2(n4590), .ZN(U3291) );
  AND2_X1 U5069 ( .A1(D_REG_30__SCAN_IN), .A2(n4590), .ZN(U3292) );
  NOR2_X1 U5070 ( .A1(n4589), .A2(n4583), .ZN(U3293) );
  AND2_X1 U5071 ( .A1(D_REG_28__SCAN_IN), .A2(n4590), .ZN(U3294) );
  AND2_X1 U5072 ( .A1(D_REG_27__SCAN_IN), .A2(n4590), .ZN(U3295) );
  AND2_X1 U5073 ( .A1(D_REG_26__SCAN_IN), .A2(n4590), .ZN(U3296) );
  AND2_X1 U5074 ( .A1(D_REG_25__SCAN_IN), .A2(n4590), .ZN(U3297) );
  AND2_X1 U5075 ( .A1(D_REG_24__SCAN_IN), .A2(n4590), .ZN(U3298) );
  NOR2_X1 U5076 ( .A1(n4589), .A2(n4584), .ZN(U3299) );
  NOR2_X1 U5077 ( .A1(n4589), .A2(n4585), .ZN(U3300) );
  AND2_X1 U5078 ( .A1(D_REG_21__SCAN_IN), .A2(n4590), .ZN(U3301) );
  AND2_X1 U5079 ( .A1(D_REG_20__SCAN_IN), .A2(n4590), .ZN(U3302) );
  AND2_X1 U5080 ( .A1(D_REG_19__SCAN_IN), .A2(n4590), .ZN(U3303) );
  AND2_X1 U5081 ( .A1(D_REG_18__SCAN_IN), .A2(n4590), .ZN(U3304) );
  AND2_X1 U5082 ( .A1(D_REG_17__SCAN_IN), .A2(n4590), .ZN(U3305) );
  AND2_X1 U5083 ( .A1(D_REG_16__SCAN_IN), .A2(n4590), .ZN(U3306) );
  AND2_X1 U5084 ( .A1(D_REG_15__SCAN_IN), .A2(n4590), .ZN(U3307) );
  AND2_X1 U5085 ( .A1(D_REG_14__SCAN_IN), .A2(n4590), .ZN(U3308) );
  AND2_X1 U5086 ( .A1(D_REG_13__SCAN_IN), .A2(n4590), .ZN(U3309) );
  AND2_X1 U5087 ( .A1(D_REG_12__SCAN_IN), .A2(n4590), .ZN(U3310) );
  AND2_X1 U5088 ( .A1(D_REG_11__SCAN_IN), .A2(n4590), .ZN(U3311) );
  AND2_X1 U5089 ( .A1(D_REG_10__SCAN_IN), .A2(n4590), .ZN(U3312) );
  AND2_X1 U5090 ( .A1(D_REG_9__SCAN_IN), .A2(n4590), .ZN(U3313) );
  AND2_X1 U5091 ( .A1(D_REG_8__SCAN_IN), .A2(n4590), .ZN(U3314) );
  AND2_X1 U5092 ( .A1(D_REG_7__SCAN_IN), .A2(n4590), .ZN(U3315) );
  AND2_X1 U5093 ( .A1(D_REG_6__SCAN_IN), .A2(n4590), .ZN(U3316) );
  NOR2_X1 U5094 ( .A1(n4589), .A2(n4586), .ZN(U3317) );
  NOR2_X1 U5095 ( .A1(n4589), .A2(n4587), .ZN(U3318) );
  NOR2_X1 U5096 ( .A1(n4589), .A2(n4588), .ZN(U3319) );
  AND2_X1 U5097 ( .A1(D_REG_2__SCAN_IN), .A2(n4590), .ZN(U3320) );
  AOI21_X1 U5098 ( .B1(U3149), .B2(n2697), .A(n4591), .ZN(U3329) );
  OAI22_X1 U5099 ( .A1(U3149), .A2(n4592), .B1(DATAI_18_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4593) );
  INV_X1 U5100 ( .A(n4593), .ZN(U3334) );
  OAI22_X1 U5101 ( .A1(U3149), .A2(n4594), .B1(DATAI_17_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4595) );
  INV_X1 U5102 ( .A(n4595), .ZN(U3335) );
  AOI22_X1 U5103 ( .A1(STATE_REG_SCAN_IN), .A2(n4597), .B1(n4596), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5104 ( .A1(STATE_REG_SCAN_IN), .A2(n4599), .B1(n4598), .B2(U3149), 
        .ZN(U3337) );
  OAI22_X1 U5105 ( .A1(U3149), .A2(n4600), .B1(DATAI_14_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4601) );
  INV_X1 U5106 ( .A(n4601), .ZN(U3338) );
  OAI22_X1 U5107 ( .A1(U3149), .A2(n4602), .B1(DATAI_12_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4603) );
  INV_X1 U5108 ( .A(n4603), .ZN(U3340) );
  AOI22_X1 U5109 ( .A1(STATE_REG_SCAN_IN), .A2(n4604), .B1(n2505), .B2(U3149), 
        .ZN(U3342) );
  AOI22_X1 U5110 ( .A1(STATE_REG_SCAN_IN), .A2(n2157), .B1(n2347), .B2(U3149), 
        .ZN(U3352) );
  AOI211_X1 U5111 ( .C1(n4641), .C2(n4607), .A(n4606), .B(n4605), .ZN(n4648)
         );
  AOI22_X1 U5112 ( .A1(n4647), .A2(n4648), .B1(n2341), .B2(n4646), .ZN(U3467)
         );
  AOI22_X1 U5113 ( .A1(n4609), .A2(n4641), .B1(n3020), .B2(n4608), .ZN(n4610)
         );
  AND2_X1 U5114 ( .A1(n4611), .A2(n4610), .ZN(n4649) );
  AOI22_X1 U5115 ( .A1(n4647), .A2(n4649), .B1(n2321), .B2(n4646), .ZN(U3469)
         );
  AND3_X1 U5116 ( .A1(n4613), .A2(n3020), .A3(n4612), .ZN(n4616) );
  INV_X1 U5117 ( .A(n4614), .ZN(n4615) );
  AOI211_X1 U5118 ( .C1(n4641), .C2(n4617), .A(n4616), .B(n4615), .ZN(n4650)
         );
  AOI22_X1 U5119 ( .A1(n4647), .A2(n4650), .B1(n2362), .B2(n4646), .ZN(U3471)
         );
  NOR2_X1 U5120 ( .A1(n4618), .A2(n4635), .ZN(n4619) );
  AOI21_X1 U5121 ( .B1(n4620), .B2(n4641), .A(n4619), .ZN(n4621) );
  AND2_X1 U5122 ( .A1(n4622), .A2(n4621), .ZN(n4651) );
  INV_X1 U5123 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4623) );
  AOI22_X1 U5124 ( .A1(n4647), .A2(n4651), .B1(n4623), .B2(n4646), .ZN(U3473)
         );
  INV_X1 U5125 ( .A(n4624), .ZN(n4626) );
  AOI211_X1 U5126 ( .C1(n4627), .C2(n4641), .A(n4626), .B(n4625), .ZN(n4652)
         );
  INV_X1 U5127 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4628) );
  AOI22_X1 U5128 ( .A1(n4647), .A2(n4652), .B1(n4628), .B2(n4646), .ZN(U3475)
         );
  NOR2_X1 U5129 ( .A1(n4630), .A2(n4629), .ZN(n4633) );
  INV_X1 U5130 ( .A(n4631), .ZN(n4632) );
  AOI211_X1 U5131 ( .C1(n3020), .C2(n4634), .A(n4633), .B(n4632), .ZN(n4654)
         );
  AOI22_X1 U5132 ( .A1(n4647), .A2(n4654), .B1(n2419), .B2(n4646), .ZN(U3477)
         );
  NOR3_X1 U5133 ( .A1(n4637), .A2(n4636), .A3(n4635), .ZN(n4639) );
  AOI211_X1 U5134 ( .C1(n4641), .C2(n4640), .A(n4639), .B(n4638), .ZN(n4655)
         );
  AOI22_X1 U5135 ( .A1(n4647), .A2(n4655), .B1(n2448), .B2(n4646), .ZN(U3479)
         );
  AOI211_X1 U5136 ( .C1(n4645), .C2(n4644), .A(n4643), .B(n4642), .ZN(n4657)
         );
  AOI22_X1 U5137 ( .A1(n4647), .A2(n4657), .B1(n2438), .B2(n4646), .ZN(U3481)
         );
  AOI22_X1 U5138 ( .A1(n4658), .A2(n4648), .B1(n2350), .B2(n4656), .ZN(U3518)
         );
  AOI22_X1 U5139 ( .A1(n4658), .A2(n4649), .B1(n2835), .B2(n4656), .ZN(U3519)
         );
  AOI22_X1 U5140 ( .A1(n4658), .A2(n4650), .B1(n2836), .B2(n4656), .ZN(U3520)
         );
  AOI22_X1 U5141 ( .A1(n4658), .A2(n4651), .B1(n2378), .B2(n4656), .ZN(U3521)
         );
  AOI22_X1 U5142 ( .A1(n4658), .A2(n4652), .B1(n4471), .B2(n4656), .ZN(U3522)
         );
  AOI22_X1 U5143 ( .A1(n4658), .A2(n4654), .B1(n4653), .B2(n4656), .ZN(U3523)
         );
  AOI22_X1 U5144 ( .A1(n4658), .A2(n4655), .B1(n2454), .B2(n4656), .ZN(U3524)
         );
  AOI22_X1 U5145 ( .A1(n4658), .A2(n4657), .B1(n2849), .B2(n4656), .ZN(U3525)
         );
  CLKBUF_X1 U2257 ( .A(n2332), .Z(n1999) );
  XNOR2_X1 U2263 ( .A(n2170), .B(n2169), .ZN(n3063) );
endmodule

