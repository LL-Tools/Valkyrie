

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2961, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793;

  AND2_X1 U3409 ( .A1(n5190), .A2(n5189), .ZN(n5504) );
  XNOR2_X1 U3410 ( .A(n5188), .B(n4263), .ZN(n5514) );
  NAND2_X1 U3411 ( .A1(n3929), .A2(n3930), .ZN(n5188) );
  NAND2_X1 U3412 ( .A1(n4418), .A2(n3016), .ZN(n6778) );
  AND2_X1 U3413 ( .A1(n3835), .A2(n3534), .ZN(n3812) );
  CLKBUF_X2 U3414 ( .A(n4282), .Z(n4310) );
  CLKBUF_X2 U3415 ( .A(n3361), .Z(n4308) );
  CLKBUF_X2 U3416 ( .A(n3475), .Z(n3499) );
  CLKBUF_X2 U3417 ( .A(n3255), .Z(n3569) );
  CLKBUF_X2 U3418 ( .A(n3345), .Z(n3469) );
  BUF_X2 U3419 ( .A(n4283), .Z(n4318) );
  AND4_X1 U3421 ( .A1(n3200), .A2(n3199), .A3(n3198), .A4(n3197), .ZN(n3206)
         );
  AND2_X1 U3422 ( .A1(n3155), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5070)
         );
  NOR2_X2 U3423 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3160) );
  AND2_X1 U3424 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4615) );
  XNOR2_X1 U3425 ( .A(n3512), .B(n3516), .ZN(n3804) );
  OAI21_X1 U3426 ( .B1(n4633), .B2(n3780), .A(n3776), .ZN(n6174) );
  NAND2_X1 U3427 ( .A1(n3467), .A2(n3466), .ZN(n4638) );
  NAND2_X1 U3428 ( .A1(n3409), .A2(n3410), .ZN(n3443) );
  NAND2_X1 U3429 ( .A1(n4138), .A2(n4068), .ZN(n4489) );
  OR2_X1 U3430 ( .A1(n3940), .A2(n3053), .ZN(n5189) );
  INV_X1 U3431 ( .A(n4963), .ZN(n3109) );
  NAND2_X1 U3432 ( .A1(n6154), .A2(n6156), .ZN(n6155) );
  CLKBUF_X3 U3433 ( .A(n4635), .Z(n2964) );
  INV_X1 U3434 ( .A(n6778), .ZN(n6054) );
  BUF_X1 U3435 ( .A(n3253), .Z(n4656) );
  OAI211_X1 U3436 ( .C1(n3546), .C2(n3822), .A(n3041), .B(n3036), .ZN(n4963)
         );
  INV_X1 U3437 ( .A(n6025), .ZN(n6790) );
  XNOR2_X1 U3438 ( .A(n3415), .B(n3414), .ZN(n4635) );
  NAND4_X4 U3439 ( .A1(n3208), .A2(n3207), .A3(n3206), .A4(n3205), .ZN(n3273)
         );
  INV_X1 U3440 ( .A(n3347), .ZN(n2961) );
  NAND2_X2 U3442 ( .A1(n5357), .A2(n3110), .ZN(n3940) );
  NAND2_X2 U3443 ( .A1(n5414), .A2(n3650), .ZN(n5357) );
  NAND2_X1 U3444 ( .A1(n6067), .A2(n4566), .ZN(n5371) );
  NOR2_X1 U34450 ( .A1(n3371), .A2(n6509), .ZN(n3426) );
  MUX2_X1 U34460 ( .A(n3832), .B(n3370), .S(n3784), .Z(n3371) );
  NOR2_X2 U34470 ( .A1(n4090), .A2(n3253), .ZN(n4076) );
  INV_X2 U34480 ( .A(n4068), .ZN(n5224) );
  INV_X4 U3449 ( .A(n4237), .ZN(n3253) );
  INV_X1 U3450 ( .A(n3759), .ZN(n3275) );
  NAND3_X2 U34510 ( .A1(n3218), .A2(n3217), .A3(n3216), .ZN(n4566) );
  CLKBUF_X2 U34520 ( .A(n3398), .Z(n4317) );
  BUF_X2 U34530 ( .A(n3254), .Z(n3454) );
  AND2_X2 U3454 ( .A1(n4600), .A2(n4593), .ZN(n3357) );
  AND2_X2 U34550 ( .A1(n4593), .A2(n3160), .ZN(n3340) );
  NAND2_X1 U34560 ( .A1(n5115), .A2(n5114), .ZN(n5382) );
  OAI21_X1 U3457 ( .B1(n5441), .B2(n6157), .A(n5440), .ZN(n5442) );
  AND2_X1 U3458 ( .A1(n4067), .A2(n3042), .ZN(n5478) );
  OAI21_X1 U34590 ( .B1(n4395), .B2(n4396), .A(n4361), .ZN(n5441) );
  AOI21_X1 U34600 ( .B1(n5080), .B2(n6262), .A(n3095), .ZN(n4262) );
  AND2_X1 U34610 ( .A1(n3131), .A2(n2994), .ZN(n3127) );
  XNOR2_X1 U34620 ( .A(n4230), .B(n4232), .ZN(n5080) );
  NAND2_X1 U34630 ( .A1(n3034), .A2(n2985), .ZN(n5634) );
  XNOR2_X1 U34640 ( .A(n6146), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5913)
         );
  NAND2_X1 U34650 ( .A1(n3101), .A2(n3104), .ZN(n5120) );
  AND2_X1 U3466 ( .A1(n3107), .A2(n4583), .ZN(n4745) );
  NAND2_X1 U3467 ( .A1(n3009), .A2(n3531), .ZN(n3835) );
  OR2_X1 U34680 ( .A1(n5250), .A2(n6554), .ZN(n5244) );
  OR2_X1 U34690 ( .A1(n4266), .A2(n3090), .ZN(n5150) );
  NAND2_X1 U34700 ( .A1(n4157), .A2(n4156), .ZN(n4266) );
  CLKBUF_X1 U34710 ( .A(n5374), .Z(n6076) );
  NAND2_X1 U34720 ( .A1(n5359), .A2(n5360), .ZN(n5362) );
  CLKBUF_X1 U34730 ( .A(n4599), .Z(n5866) );
  AND2_X1 U34740 ( .A1(n4215), .A2(n4214), .ZN(n4239) );
  NOR2_X1 U3475 ( .A1(n4682), .A2(n4656), .ZN(n6417) );
  NOR2_X1 U3476 ( .A1(n4682), .A2(n3274), .ZN(n6435) );
  NOR2_X1 U3477 ( .A1(n4682), .A2(n4069), .ZN(n6423) );
  NOR2_X1 U3478 ( .A1(n4682), .A2(n5373), .ZN(n6456) );
  NOR2_X1 U3479 ( .A1(n4682), .A2(n3275), .ZN(n6441) );
  NOR2_X1 U3480 ( .A1(n4683), .A2(n5010), .ZN(n6413) );
  NOR2_X1 U3481 ( .A1(n4682), .A2(n4660), .ZN(n6447) );
  NAND2_X2 U3482 ( .A1(n3430), .A2(n3429), .ZN(n6275) );
  OR2_X1 U3483 ( .A1(n5276), .A2(n5986), .ZN(n5987) );
  NAND2_X1 U3484 ( .A1(n3299), .A2(n3382), .ZN(n3322) );
  AOI21_X1 U3485 ( .B1(n3446), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3389), 
        .ZN(n3390) );
  AND2_X1 U3486 ( .A1(n3429), .A2(n3373), .ZN(n3374) );
  AOI21_X1 U3487 ( .B1(n3314), .B2(n3313), .A(n3312), .ZN(n4081) );
  INV_X1 U3488 ( .A(n3302), .ZN(n3902) );
  CLKBUF_X1 U3489 ( .A(n4082), .Z(n4561) );
  NAND2_X1 U3490 ( .A1(n3070), .A2(n3069), .ZN(n3302) );
  AND2_X1 U3491 ( .A1(n3272), .A2(n4084), .ZN(n3309) );
  AOI21_X1 U3492 ( .B1(n3275), .B2(n3283), .A(n4078), .ZN(n3276) );
  CLKBUF_X1 U3493 ( .A(n3303), .Z(n6605) );
  NAND2_X1 U3494 ( .A1(n4068), .A2(n4549), .ZN(n4223) );
  AND2_X1 U3495 ( .A1(n3266), .A2(n4077), .ZN(n3774) );
  AND2_X1 U3496 ( .A1(n4069), .A2(n4077), .ZN(n3786) );
  CLKBUF_X1 U3497 ( .A(n3307), .Z(n4660) );
  NOR2_X1 U3498 ( .A1(n4212), .A2(n4077), .ZN(n4092) );
  NAND2_X1 U3499 ( .A1(n3307), .A2(n3759), .ZN(n3289) );
  INV_X2 U3500 ( .A(n5224), .ZN(n2963) );
  INV_X2 U3501 ( .A(n4090), .ZN(n4681) );
  NAND2_X4 U3502 ( .A1(n4077), .A2(n4237), .ZN(n4068) );
  OR2_X1 U3503 ( .A1(n3353), .A2(n3352), .ZN(n3784) );
  NAND3_X1 U3504 ( .A1(n3367), .A2(n3144), .A3(n3152), .ZN(n3837) );
  INV_X1 U3505 ( .A(n3286), .ZN(n3307) );
  NAND2_X2 U3506 ( .A1(n3165), .A2(n2975), .ZN(n3759) );
  NAND2_X1 U3507 ( .A1(n3185), .A2(n3184), .ZN(n3284) );
  AND2_X1 U3508 ( .A1(n3232), .A2(n3231), .ZN(n3242) );
  AND4_X1 U3509 ( .A1(n3159), .A2(n3158), .A3(n3157), .A4(n3156), .ZN(n3165)
         );
  AND3_X1 U3510 ( .A1(n3215), .A2(n3214), .A3(n3213), .ZN(n3217) );
  AND4_X1 U3511 ( .A1(n3212), .A2(n3211), .A3(n3210), .A4(n3209), .ZN(n3218)
         );
  AND4_X1 U3512 ( .A1(n3230), .A2(n3229), .A3(n3228), .A4(n3227), .ZN(n3231)
         );
  AND4_X1 U3513 ( .A1(n3226), .A2(n3225), .A3(n3224), .A4(n3223), .ZN(n3232)
         );
  AND4_X1 U3514 ( .A1(n3196), .A2(n3195), .A3(n3194), .A4(n3193), .ZN(n3207)
         );
  AND4_X1 U3515 ( .A1(n3183), .A2(n3182), .A3(n3181), .A4(n3180), .ZN(n3184)
         );
  AND4_X1 U3516 ( .A1(n3179), .A2(n3178), .A3(n3177), .A4(n3176), .ZN(n3185)
         );
  CLKBUF_X1 U3517 ( .A(n6598), .Z(n6579) );
  CLKBUF_X2 U3518 ( .A(n3357), .Z(n4316) );
  AND2_X2 U3519 ( .A1(n5229), .A2(n6509), .ZN(n6233) );
  AND2_X2 U3520 ( .A1(n5070), .A2(n3160), .ZN(n3398) );
  NOR2_X1 U3521 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6524), .ZN(n6615) );
  AND2_X2 U3522 ( .A1(n4593), .A2(n4615), .ZN(n3346) );
  AND2_X2 U3523 ( .A1(n4618), .A2(n3160), .ZN(n4283) );
  AND2_X2 U3524 ( .A1(n3416), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5068)
         );
  INV_X2 U3525 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6509) );
  NOR2_X2 U3526 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4618) );
  AND2_X2 U3527 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4593) );
  AND2_X2 U3528 ( .A1(n4615), .A2(n5070), .ZN(n3393) );
  INV_X1 U3529 ( .A(n3532), .ZN(n3531) );
  INV_X1 U3530 ( .A(n3533), .ZN(n3009) );
  NOR2_X1 U3531 ( .A1(n3051), .A2(n3050), .ZN(n3049) );
  INV_X1 U3532 ( .A(n5367), .ZN(n3050) );
  NOR2_X1 U3534 ( .A1(n4088), .A2(n6509), .ZN(n4354) );
  INV_X1 U3535 ( .A(n4023), .ZN(n4357) );
  AND2_X2 U3536 ( .A1(n3278), .A2(n3273), .ZN(n3871) );
  INV_X1 U3537 ( .A(n3864), .ZN(n3278) );
  NOR3_X1 U3538 ( .A1(n4426), .A2(n4425), .A3(n4424), .ZN(n4427) );
  INV_X1 U3539 ( .A(n4417), .ZN(n4426) );
  OAI21_X1 U3540 ( .B1(n3888), .B2(n3511), .A(n3510), .ZN(n3516) );
  NAND2_X1 U3541 ( .A1(n4090), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3864) );
  AND2_X1 U3542 ( .A1(n3253), .A2(n4090), .ZN(n3303) );
  AND2_X1 U3543 ( .A1(n3148), .A2(n3118), .ZN(n3117) );
  INV_X1 U3544 ( .A(n5113), .ZN(n3118) );
  NOR2_X1 U3545 ( .A1(n5260), .A2(n3114), .ZN(n3113) );
  INV_X1 U3546 ( .A(n5356), .ZN(n3114) );
  NAND2_X1 U3547 ( .A1(n3108), .A2(n3052), .ZN(n3051) );
  INV_X1 U3548 ( .A(n5419), .ZN(n3052) );
  INV_X1 U3549 ( .A(n4746), .ZN(n3041) );
  XNOR2_X1 U3550 ( .A(n3835), .B(n3543), .ZN(n3822) );
  INV_X1 U3551 ( .A(n3627), .ZN(n3678) );
  NAND2_X1 U3552 ( .A1(n4660), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3627) );
  OR2_X1 U3553 ( .A1(n5262), .A2(n5349), .ZN(n3098) );
  NOR2_X2 U3554 ( .A1(n5987), .A2(n4136), .ZN(n5363) );
  AND2_X1 U3555 ( .A1(n3902), .A2(n3903), .ZN(n4219) );
  NAND2_X1 U3556 ( .A1(n3274), .A2(n3837), .ZN(n3832) );
  INV_X1 U3557 ( .A(n3871), .ZN(n3888) );
  NAND2_X1 U3558 ( .A1(n3871), .A2(n3870), .ZN(n3900) );
  AND4_X1 U3559 ( .A1(n3204), .A2(n3203), .A3(n3202), .A4(n3201), .ZN(n3205)
         );
  AND4_X1 U3560 ( .A1(n3192), .A2(n3191), .A3(n3190), .A4(n3189), .ZN(n3208)
         );
  INV_X1 U3561 ( .A(n3636), .ZN(n3634) );
  NAND2_X1 U3562 ( .A1(n4044), .A2(n4043), .ZN(n5148) );
  NAND2_X1 U3563 ( .A1(n3044), .A2(n3043), .ZN(n4067) );
  INV_X1 U3564 ( .A(n5148), .ZN(n3043) );
  NAND2_X1 U3565 ( .A1(n3980), .A2(n3055), .ZN(n3054) );
  INV_X1 U3566 ( .A(n5172), .ZN(n3055) );
  INV_X1 U3567 ( .A(n5434), .ZN(n3120) );
  NAND2_X1 U3568 ( .A1(n3068), .A2(n3067), .ZN(n5446) );
  AND2_X1 U3569 ( .A1(n5462), .A2(n3001), .ZN(n3067) );
  NAND2_X1 U3570 ( .A1(n3030), .A2(n3029), .ZN(n4214) );
  AND2_X1 U3571 ( .A1(n5307), .A2(n4399), .ZN(n6025) );
  NOR2_X1 U3572 ( .A1(n4418), .A2(n6749), .ZN(n4399) );
  NOR2_X1 U3573 ( .A1(n3017), .A2(n6749), .ZN(n3016) );
  INV_X1 U3574 ( .A(n6250), .ZN(n6262) );
  BUF_X1 U3575 ( .A(n3453), .Z(n4307) );
  AND2_X1 U3576 ( .A1(n3516), .A2(n3515), .ZN(n3517) );
  OR2_X1 U3577 ( .A1(n3528), .A2(n3527), .ZN(n3824) );
  OR2_X1 U3578 ( .A1(n3509), .A2(n3508), .ZN(n3813) );
  AND2_X1 U3579 ( .A1(n3280), .A2(n3279), .ZN(n3295) );
  OR2_X1 U3580 ( .A1(n3890), .A2(n3889), .ZN(n3892) );
  AND2_X1 U3581 ( .A1(n6478), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3889)
         );
  AND2_X1 U3582 ( .A1(n4203), .A2(n4198), .ZN(n3895) );
  AOI22_X1 U3584 ( .A1(n3398), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3357), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3173) );
  NOR2_X1 U3585 ( .A1(n3979), .A2(n5187), .ZN(n3980) );
  AND2_X1 U3586 ( .A1(n3596), .A2(n3581), .ZN(n3108) );
  NOR2_X1 U3587 ( .A1(n5130), .A2(n5118), .ZN(n3104) );
  INV_X1 U3588 ( .A(n5472), .ZN(n3068) );
  OAI21_X1 U3589 ( .B1(n3846), .B2(n3062), .A(n3002), .ZN(n3004) );
  INV_X1 U3590 ( .A(n3127), .ZN(n3003) );
  NOR2_X1 U3591 ( .A1(n3138), .A2(n3063), .ZN(n3135) );
  OR2_X1 U3592 ( .A1(n3093), .A2(n3092), .ZN(n3091) );
  INV_X1 U3593 ( .A(n5175), .ZN(n3092) );
  INV_X1 U3594 ( .A(n4838), .ZN(n4119) );
  NAND2_X1 U3595 ( .A1(n4599), .A2(n6509), .ZN(n3467) );
  AND2_X1 U3596 ( .A1(n3447), .A2(n4685), .ZN(n5009) );
  INV_X1 U3597 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6474) );
  INV_X1 U3598 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4936) );
  OR2_X2 U3599 ( .A1(n3265), .A2(n3264), .ZN(n4077) );
  OAI21_X1 U3600 ( .B1(n6610), .B2(n4627), .A(n6502), .ZN(n4649) );
  INV_X1 U3601 ( .A(n3899), .ZN(n4202) );
  NAND2_X1 U3602 ( .A1(n3028), .A2(n3872), .ZN(n3873) );
  OAI211_X1 U3603 ( .C1(n2966), .C2(n2987), .A(n3024), .B(n2980), .ZN(n3028)
         );
  INV_X1 U3604 ( .A(n3486), .ZN(n3489) );
  OR2_X1 U3605 ( .A1(n6233), .A2(n6508), .ZN(n4398) );
  AND4_X1 U3606 ( .A1(n3236), .A2(n3235), .A3(n3234), .A4(n3233), .ZN(n3241)
         );
  AND4_X1 U3607 ( .A1(n3240), .A2(n3239), .A3(n3238), .A4(n3237), .ZN(n3150)
         );
  AND2_X1 U3608 ( .A1(n4152), .A2(n5223), .ZN(n5226) );
  OAI21_X1 U3609 ( .B1(n3492), .B2(n5450), .A(n4351), .ZN(n5113) );
  BUF_X1 U3610 ( .A(n3759), .Z(n5372) );
  MUX2_X1 U3611 ( .A(n5183), .B(n4520), .S(n4519), .Z(n4570) );
  OR2_X1 U3612 ( .A1(n4456), .A2(READY_N), .ZN(n4457) );
  INV_X1 U3613 ( .A(n4021), .ZN(n4384) );
  NAND2_X1 U3614 ( .A1(n3715), .A2(n3022), .ZN(n3914) );
  AND2_X1 U3615 ( .A1(n2969), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3022)
         );
  NAND2_X1 U3616 ( .A1(n3715), .A2(n2969), .ZN(n3750) );
  NAND2_X1 U3617 ( .A1(n3715), .A2(n3714), .ZN(n3722) );
  NOR2_X1 U3618 ( .A1(n3112), .A2(n3111), .ZN(n3110) );
  INV_X1 U3619 ( .A(n5347), .ZN(n3111) );
  INV_X1 U3620 ( .A(n3113), .ZN(n3112) );
  NAND2_X1 U3621 ( .A1(n3681), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3717)
         );
  NAND2_X1 U3622 ( .A1(n3597), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3598)
         );
  NOR2_X1 U3623 ( .A1(n6673), .A2(n3598), .ZN(n3629) );
  AND2_X1 U3624 ( .A1(n3592), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3597)
         );
  OR2_X1 U3625 ( .A1(n3557), .A2(n6011), .ZN(n3558) );
  NOR2_X1 U3626 ( .A1(n4753), .A2(n2977), .ZN(n3036) );
  OR2_X1 U3627 ( .A1(n3546), .A2(n3678), .ZN(n3038) );
  NAND2_X1 U3628 ( .A1(n3041), .A2(n3040), .ZN(n5000) );
  AND2_X1 U3629 ( .A1(n3037), .A2(n3039), .ZN(n4999) );
  NAND2_X1 U3630 ( .A1(n3822), .A2(n3678), .ZN(n3037) );
  NOR2_X1 U3631 ( .A1(n3535), .A2(n3012), .ZN(n3011) );
  INV_X1 U3632 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3012) );
  AOI21_X1 U3633 ( .B1(n4546), .B2(n4547), .A(n3792), .ZN(n6175) );
  NAND2_X1 U3634 ( .A1(n3068), .A2(n5462), .ZN(n5454) );
  NOR2_X1 U3635 ( .A1(n5150), .A2(n5149), .ZN(n5152) );
  NAND2_X1 U3636 ( .A1(n3065), .A2(n3064), .ZN(n3139) );
  AOI21_X1 U3637 ( .B1(n3082), .B2(n3851), .A(n2968), .ZN(n3065) );
  NAND2_X1 U3638 ( .A1(n3125), .A2(n3066), .ZN(n3064) );
  NAND2_X1 U3639 ( .A1(n3139), .A2(n3137), .ZN(n5472) );
  OR2_X1 U3640 ( .A1(n3091), .A2(n4377), .ZN(n3090) );
  XNOR2_X1 U3641 ( .A(n3076), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3074)
         );
  AND2_X1 U3642 ( .A1(n3078), .A2(n2998), .ZN(n3076) );
  NAND2_X1 U3643 ( .A1(n5533), .A2(n6707), .ZN(n3078) );
  NAND2_X1 U3644 ( .A1(n3035), .A2(n4245), .ZN(n5653) );
  OAI21_X1 U3645 ( .B1(n2990), .B2(n5678), .A(n5489), .ZN(n3035) );
  NAND2_X1 U3646 ( .A1(n3080), .A2(n3079), .ZN(n4375) );
  AOI21_X1 U3647 ( .B1(n2967), .B2(n3063), .A(n2984), .ZN(n3079) );
  NAND2_X1 U3648 ( .A1(n3097), .A2(n5248), .ZN(n3096) );
  INV_X1 U3649 ( .A(n3098), .ZN(n3097) );
  INV_X1 U3650 ( .A(n6196), .ZN(n5718) );
  INV_X1 U3651 ( .A(n3846), .ZN(n3130) );
  AOI21_X1 U3652 ( .B1(n5913), .B2(n3132), .A(n2982), .ZN(n3131) );
  INV_X1 U3653 ( .A(n5552), .ZN(n3132) );
  NAND2_X1 U3654 ( .A1(n3122), .A2(n3124), .ZN(n3121) );
  OR2_X1 U3655 ( .A1(n6146), .A2(n5751), .ZN(n5553) );
  NOR2_X1 U3656 ( .A1(n6192), .A2(n4242), .ZN(n5713) );
  NOR2_X1 U3657 ( .A1(n2965), .A2(n3087), .ZN(n3086) );
  INV_X1 U3658 ( .A(n5277), .ZN(n3087) );
  INV_X1 U3659 ( .A(n6264), .ZN(n6200) );
  AOI22_X1 U3660 ( .A1(n3871), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3406), 
        .B2(n3405), .ZN(n3407) );
  NAND2_X1 U3661 ( .A1(n3005), .A2(n2988), .ZN(n3408) );
  INV_X1 U3662 ( .A(n6313), .ZN(n3119) );
  NAND2_X1 U3663 ( .A1(n4539), .A2(n4538), .ZN(n6469) );
  AND2_X1 U3664 ( .A1(n6316), .A2(n6315), .ZN(n6320) );
  INV_X1 U3665 ( .A(n5866), .ZN(n6278) );
  NAND2_X1 U3666 ( .A1(n4637), .A2(n4633), .ZN(n6403) );
  OAI21_X1 U3667 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6588), .A(n4891), 
        .ZN(n6405) );
  NAND2_X1 U3668 ( .A1(n6509), .A2(n4649), .ZN(n5010) );
  AND2_X1 U3669 ( .A1(n6749), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3901) );
  AOI21_X1 U3670 ( .B1(n5251), .B2(REIP_REG_18__SCAN_IN), .A(n3015), .ZN(n3014) );
  OAI22_X1 U3671 ( .A1(n6029), .A2(n5343), .B1(n5694), .B2(n6044), .ZN(n3015)
         );
  AND2_X1 U3672 ( .A1(n5307), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6779) );
  INV_X1 U3673 ( .A(n6781), .ZN(n6033) );
  NAND2_X1 U3674 ( .A1(n6067), .A2(n5373), .ZN(n5369) );
  NAND2_X1 U3675 ( .A1(n3757), .A2(n3756), .ZN(n5407) );
  NAND2_X1 U3676 ( .A1(n3754), .A2(n3755), .ZN(n3756) );
  AND2_X1 U3677 ( .A1(n5416), .A2(n4568), .ZN(n5422) );
  XNOR2_X1 U3678 ( .A(n4389), .B(n5092), .ZN(n4418) );
  INV_X1 U3679 ( .A(n4387), .ZN(n4388) );
  AOI21_X1 U3680 ( .B1(n4067), .B2(n4066), .A(n5128), .ZN(n5469) );
  NOR2_X1 U3681 ( .A1(n4061), .A2(n3145), .ZN(n4066) );
  OR2_X2 U3682 ( .A1(n4558), .A2(n6481), .ZN(n6159) );
  NAND2_X1 U3683 ( .A1(n3120), .A2(n3000), .ZN(n4188) );
  NOR2_X1 U3684 ( .A1(n5601), .A2(n3033), .ZN(n5593) );
  AND2_X1 U3685 ( .A1(n6196), .A2(n5589), .ZN(n3033) );
  NOR2_X1 U3686 ( .A1(n5634), .A2(n4248), .ZN(n5621) );
  AND2_X1 U3687 ( .A1(n5919), .A2(n5717), .ZN(n5732) );
  OR2_X1 U3688 ( .A1(n4239), .A2(n4221), .ZN(n6184) );
  OR2_X1 U3689 ( .A1(n4239), .A2(n4236), .ZN(n6250) );
  NAND2_X1 U3690 ( .A1(n3428), .A2(n3427), .ZN(n3430) );
  INV_X1 U3691 ( .A(n3426), .ZN(n3427) );
  INV_X1 U3692 ( .A(n6401), .ZN(n6406) );
  NOR2_X2 U3693 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6401) );
  INV_X1 U3694 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6478) );
  AND2_X1 U3695 ( .A1(n4089), .A2(n4566), .ZN(n3069) );
  AOI22_X1 U3696 ( .A1(n3361), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3453), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3166) );
  AOI22_X1 U3697 ( .A1(n4282), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3169) );
  AOI22_X1 U3698 ( .A1(n3340), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3170) );
  OAI21_X1 U3699 ( .B1(n3888), .B2(n3483), .A(n3482), .ZN(n3515) );
  NAND2_X1 U3700 ( .A1(n3835), .A2(n3834), .ZN(n3848) );
  NOR2_X1 U3701 ( .A1(n3833), .A2(n3832), .ZN(n3834) );
  NAND2_X1 U3702 ( .A1(n4681), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3452) );
  OR2_X1 U3703 ( .A1(n3465), .A2(n3464), .ZN(n3764) );
  AOI22_X1 U3704 ( .A1(n3361), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4282), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3179) );
  OR2_X1 U3705 ( .A1(n3866), .A2(n3867), .ZN(n3026) );
  NAND2_X1 U3706 ( .A1(n3900), .A2(n3869), .ZN(n3025) );
  NAND2_X1 U3708 ( .A1(n4089), .A2(n3269), .ZN(n4073) );
  INV_X1 U3709 ( .A(n4431), .ZN(n3103) );
  NAND2_X1 U3710 ( .A1(n3346), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3202)
         );
  AOI22_X1 U3711 ( .A1(n3355), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3398), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3209) );
  OR2_X1 U3712 ( .A1(n4058), .A2(n4057), .ZN(n4305) );
  NOR2_X1 U3713 ( .A1(n4018), .A2(n3019), .ZN(n3018) );
  INV_X1 U3714 ( .A(n3717), .ZN(n3715) );
  XNOR2_X1 U3715 ( .A(n3498), .B(n3515), .ZN(n3761) );
  OR2_X1 U3716 ( .A1(n4265), .A2(n3094), .ZN(n3093) );
  INV_X1 U3717 ( .A(n5193), .ZN(n3094) );
  NAND2_X1 U3718 ( .A1(n3851), .A2(n3082), .ZN(n3081) );
  NAND2_X1 U3719 ( .A1(n5573), .A2(n3123), .ZN(n3061) );
  INV_X1 U3720 ( .A(n3841), .ZN(n3123) );
  NAND2_X1 U3721 ( .A1(n3060), .A2(n5582), .ZN(n3058) );
  AND2_X1 U3722 ( .A1(n3061), .A2(n3843), .ZN(n3122) );
  INV_X1 U3723 ( .A(n5573), .ZN(n3124) );
  NAND2_X1 U3724 ( .A1(n3089), .A2(n4119), .ZN(n3088) );
  INV_X1 U3725 ( .A(n5001), .ZN(n3089) );
  NAND2_X1 U3726 ( .A1(n3819), .A2(n3818), .ZN(n3820) );
  NAND2_X1 U3727 ( .A1(n3812), .A2(n3870), .ZN(n3819) );
  NAND2_X1 U3728 ( .A1(n3809), .A2(n3808), .ZN(n3810) );
  NOR2_X1 U3729 ( .A1(n4213), .A2(n4212), .ZN(n3029) );
  OR2_X1 U3730 ( .A1(n3332), .A2(n3331), .ZN(n3785) );
  OR2_X1 U3731 ( .A1(n3404), .A2(n3403), .ZN(n3405) );
  OR2_X1 U3732 ( .A1(n3273), .A2(n6509), .ZN(n3451) );
  INV_X1 U3733 ( .A(n3405), .ZN(n3772) );
  OR2_X1 U3734 ( .A1(n3685), .A2(n3686), .ZN(n4088) );
  AND2_X2 U3735 ( .A1(n3856), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4600)
         );
  INV_X1 U3736 ( .A(n4068), .ZN(n3271) );
  NAND2_X1 U3737 ( .A1(n3450), .A2(n3449), .ZN(n4621) );
  AND2_X1 U3738 ( .A1(n6398), .A2(n3388), .ZN(n4849) );
  NOR2_X1 U3739 ( .A1(n4633), .A2(n4634), .ZN(n4643) );
  AND2_X1 U3740 ( .A1(n3282), .A2(n3281), .ZN(n4209) );
  AND3_X1 U3741 ( .A1(n3786), .A2(n3307), .A3(n3289), .ZN(n3282) );
  INV_X1 U3742 ( .A(n4073), .ZN(n3281) );
  NAND2_X1 U3743 ( .A1(n4209), .A2(n4090), .ZN(n4444) );
  OR2_X1 U3744 ( .A1(n4558), .A2(n4444), .ZN(n4456) );
  NAND2_X1 U3745 ( .A1(n6510), .A2(n6509), .ZN(n3904) );
  AND2_X1 U3746 ( .A1(n4204), .A2(n4203), .ZN(n4447) );
  AND2_X1 U3747 ( .A1(n5980), .A2(n5307), .ZN(n5274) );
  AND2_X1 U3748 ( .A1(n5152), .A2(n3099), .ZN(n4364) );
  NOR2_X1 U3749 ( .A1(n3102), .A2(n3100), .ZN(n3099) );
  INV_X1 U3750 ( .A(n4175), .ZN(n3100) );
  NAND2_X1 U3751 ( .A1(n3104), .A2(n3103), .ZN(n3102) );
  AND2_X1 U3752 ( .A1(n4146), .A2(n4145), .ZN(n5349) );
  NOR2_X1 U3753 ( .A1(n3085), .A2(n3083), .ZN(n4585) );
  OAI21_X1 U3754 ( .B1(n4223), .B2(EBX_REG_3__SCAN_IN), .A(n3084), .ZN(n3083)
         );
  NOR2_X1 U3755 ( .A1(n4489), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3085)
         );
  NAND2_X1 U3756 ( .A1(n5224), .A2(EBX_REG_3__SCAN_IN), .ZN(n3084) );
  NAND2_X1 U3757 ( .A1(n4271), .A2(n2972), .ZN(n4387) );
  AND2_X1 U3758 ( .A1(n4343), .A2(n3115), .ZN(n4386) );
  AND2_X1 U3759 ( .A1(n2978), .A2(n3116), .ZN(n3115) );
  INV_X1 U3760 ( .A(n4362), .ZN(n3116) );
  NAND2_X1 U3761 ( .A1(n4271), .A2(n2971), .ZN(n4358) );
  OR2_X1 U3762 ( .A1(n3021), .A2(n3020), .ZN(n4337) );
  NAND2_X1 U3763 ( .A1(n3956), .A2(n3018), .ZN(n4045) );
  NOR2_X1 U3764 ( .A1(n3976), .A2(n3972), .ZN(n3956) );
  NAND2_X1 U3765 ( .A1(n3956), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4019)
         );
  INV_X1 U3766 ( .A(n3980), .ZN(n3053) );
  OR2_X1 U3767 ( .A1(n3914), .A2(n5210), .ZN(n3976) );
  AND2_X1 U3768 ( .A1(n3720), .A2(n3719), .ZN(n5246) );
  AND3_X1 U3769 ( .A1(n3684), .A2(n3683), .A3(n3682), .ZN(n5260) );
  INV_X1 U3770 ( .A(n3653), .ZN(n3654) );
  AND2_X1 U3771 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n3654), .ZN(n3681)
         );
  AND2_X1 U3772 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n3629), .ZN(n3630)
         );
  NAND2_X1 U3773 ( .A1(n3630), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3653)
         );
  AND2_X1 U3774 ( .A1(n3614), .A2(n3613), .ZN(n5419) );
  INV_X1 U3775 ( .A(n3051), .ZN(n3048) );
  AND3_X1 U3776 ( .A1(n3595), .A2(n3594), .A3(n3593), .ZN(n5270) );
  NOR2_X1 U3777 ( .A1(n6706), .A2(n3558), .ZN(n3592) );
  INV_X1 U3778 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6706) );
  NAND2_X1 U3779 ( .A1(n3491), .A2(n2979), .ZN(n3557) );
  NAND2_X1 U3780 ( .A1(n3105), .A2(n3514), .ZN(n4748) );
  CLKBUF_X1 U3781 ( .A(n4746), .Z(n4747) );
  NAND2_X1 U3782 ( .A1(n3491), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3536)
         );
  AND2_X1 U3783 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3489), .ZN(n3491)
         );
  NAND2_X1 U3784 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3486) );
  AND3_X2 U3785 ( .A1(n3106), .A2(n3441), .A3(n3442), .ZN(n4744) );
  NAND2_X1 U3786 ( .A1(n4581), .A2(n3154), .ZN(n3106) );
  AOI21_X1 U3787 ( .B1(n4489), .B2(EBX_REG_30__SCAN_IN), .A(n4222), .ZN(n4365)
         );
  INV_X1 U3788 ( .A(n5446), .ZN(n5426) );
  NAND2_X1 U3789 ( .A1(n5621), .A2(n2981), .ZN(n5601) );
  INV_X1 U3790 ( .A(n4225), .ZN(n3101) );
  AOI21_X1 U3791 ( .B1(n3137), .B2(n2968), .A(n2983), .ZN(n3136) );
  NAND2_X1 U3792 ( .A1(n3004), .A2(n3135), .ZN(n3134) );
  AND2_X1 U3793 ( .A1(n4164), .A2(n4163), .ZN(n5175) );
  INV_X1 U3794 ( .A(n4155), .ZN(n4156) );
  INV_X1 U3795 ( .A(n5211), .ZN(n4157) );
  INV_X1 U3796 ( .A(n5917), .ZN(n4140) );
  INV_X1 U3797 ( .A(n5363), .ZN(n5916) );
  AND2_X1 U3798 ( .A1(n5562), .A2(n5574), .ZN(n6145) );
  NAND2_X1 U3799 ( .A1(n3057), .A2(n3831), .ZN(n3056) );
  INV_X1 U3800 ( .A(n5045), .ZN(n3057) );
  AND2_X1 U3801 ( .A1(n4129), .A2(n4128), .ZN(n5056) );
  NAND2_X1 U3802 ( .A1(n6264), .A2(n6201), .ZN(n6192) );
  AND2_X1 U3803 ( .A1(n4118), .A2(n4117), .ZN(n4838) );
  NAND2_X1 U3804 ( .A1(n4120), .A2(n4119), .ZN(n5002) );
  AND2_X1 U3805 ( .A1(n6401), .A2(n6749), .ZN(n5229) );
  INV_X1 U3806 ( .A(n4737), .ZN(n4114) );
  XNOR2_X1 U3807 ( .A(n3810), .B(n4734), .ZN(n4729) );
  AND2_X1 U3808 ( .A1(n5085), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6164)
         );
  AND2_X1 U3809 ( .A1(n3796), .A2(n3795), .ZN(n5086) );
  AND2_X2 U3810 ( .A1(n4237), .A2(n4090), .ZN(n4549) );
  NAND2_X1 U3811 ( .A1(n5738), .A2(n5737), .ZN(n6196) );
  INV_X1 U3812 ( .A(n4549), .ZN(n4231) );
  INV_X1 U3813 ( .A(n4209), .ZN(n4540) );
  AND2_X1 U3814 ( .A1(n3286), .A2(n4566), .ZN(n4233) );
  NAND2_X1 U3815 ( .A1(n4138), .A2(EBX_REG_0__SCAN_IN), .ZN(n4105) );
  OAI21_X1 U3816 ( .B1(n6275), .B2(n3780), .A(n3779), .ZN(n4487) );
  OAI211_X1 U3817 ( .C1(n3888), .C2(n3369), .A(n3368), .B(n3832), .ZN(n3424)
         );
  OR2_X1 U3818 ( .A1(n3413), .A2(n3412), .ZN(n3380) );
  NAND2_X1 U3819 ( .A1(n3008), .A2(n3007), .ZN(n3006) );
  INV_X1 U3820 ( .A(n3391), .ZN(n3007) );
  XNOR2_X1 U3821 ( .A(n4620), .B(n4621), .ZN(n4599) );
  INV_X1 U3822 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3416) );
  INV_X1 U3823 ( .A(n3383), .ZN(n3321) );
  INV_X1 U3824 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3155) );
  CLKBUF_X1 U3825 ( .A(n3444), .Z(n4620) );
  AOI21_X1 U3826 ( .B1(n4768), .B2(n6401), .A(n4842), .ZN(n4847) );
  AND2_X1 U3827 ( .A1(n4590), .A2(n5759), .ZN(n5831) );
  AOI21_X1 U3828 ( .B1(n5864), .B2(STATEBS16_REG_SCAN_IN), .A(n6406), .ZN(
        n5872) );
  OR2_X1 U3829 ( .A1(n5907), .A2(n6449), .ZN(n5864) );
  AND2_X1 U3830 ( .A1(n2964), .A2(n5767), .ZN(n5821) );
  NAND2_X1 U3831 ( .A1(n4643), .A2(n4758), .ZN(n4811) );
  NAND3_X1 U3832 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6509), .A3(n4649), .ZN(
        n4682) );
  AND2_X1 U3833 ( .A1(n4849), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6279) );
  INV_X1 U3834 ( .A(n3032), .ZN(n3031) );
  AOI21_X1 U3835 ( .B1(n3898), .B2(n3897), .A(n3896), .ZN(n3032) );
  AND2_X1 U3836 ( .A1(n6509), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4397) );
  INV_X1 U3837 ( .A(n6503), .ZN(n6610) );
  OR2_X1 U3838 ( .A1(n5146), .A2(n4415), .ZN(n5116) );
  NOR2_X1 U3839 ( .A1(n5976), .A2(n4403), .ZN(n5960) );
  NAND2_X1 U3840 ( .A1(n6775), .A2(n4407), .ZN(n5976) );
  INV_X1 U3841 ( .A(n6779), .ZN(n6047) );
  INV_X1 U3842 ( .A(n5274), .ZN(n6030) );
  INV_X1 U3843 ( .A(n4395), .ZN(n5115) );
  NOR2_X2 U3844 ( .A1(n6075), .A2(n5100), .ZN(n6072) );
  NAND2_X1 U3845 ( .A1(n3650), .A2(n3638), .ZN(n3047) );
  AOI21_X1 U3846 ( .B1(n3030), .B2(n4564), .A(n4563), .ZN(n4565) );
  INV_X2 U3847 ( .A(n6073), .ZN(n5424) );
  INV_X1 U3848 ( .A(n5422), .ZN(n5417) );
  NOR2_X1 U3849 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4629), .ZN(n6085) );
  INV_X1 U3850 ( .A(n6085), .ZN(n6111) );
  OR3_X1 U3851 ( .A1(n4558), .A2(n4497), .A3(n6603), .ZN(n6114) );
  AND2_X1 U3852 ( .A1(n5073), .A2(n6492), .ZN(n4497) );
  INV_X1 U3853 ( .A(n6111), .ZN(n6601) );
  INV_X2 U3854 ( .A(n6108), .ZN(n6112) );
  INV_X2 U3855 ( .A(n6142), .ZN(n6136) );
  OR2_X1 U3856 ( .A1(n4457), .A2(n4656), .ZN(n6125) );
  AOI21_X1 U3857 ( .B1(n4362), .B2(n4361), .A(n4386), .ZN(n5432) );
  NAND2_X1 U3858 ( .A1(n5162), .A2(n5148), .ZN(n3042) );
  AOI21_X1 U3859 ( .B1(n5164), .B2(n5163), .A(n3044), .ZN(n5484) );
  AOI21_X1 U3860 ( .B1(n5189), .B2(n5172), .A(n5161), .ZN(n5496) );
  NOR2_X1 U3861 ( .A1(n5000), .A2(n4999), .ZN(n4965) );
  NAND2_X1 U3862 ( .A1(n3120), .A2(n4185), .ZN(n5427) );
  AOI21_X1 U3863 ( .B1(n5611), .B2(n5434), .A(n5448), .ZN(n5617) );
  NOR2_X1 U3864 ( .A1(n5629), .A2(n5630), .ZN(n5623) );
  AND2_X1 U3865 ( .A1(n3139), .A2(n2973), .ZN(n5471) );
  INV_X1 U3866 ( .A(n5644), .ZN(n3034) );
  XNOR2_X1 U3867 ( .A(n3077), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3075)
         );
  NAND2_X1 U3868 ( .A1(n5506), .A2(n3074), .ZN(n3073) );
  NAND2_X1 U3869 ( .A1(n5498), .A2(n5649), .ZN(n3077) );
  AND2_X1 U3870 ( .A1(n5667), .A2(n5490), .ZN(n5650) );
  OAI22_X1 U3871 ( .A1(n5506), .A2(n3010), .B1(n5535), .B2(n5491), .ZN(n5492)
         );
  INV_X1 U3872 ( .A(n5498), .ZN(n3010) );
  NAND2_X1 U3873 ( .A1(n5506), .A2(n3078), .ZN(n5500) );
  NAND2_X1 U3874 ( .A1(n5732), .A2(n4256), .ZN(n5695) );
  NAND2_X1 U3875 ( .A1(n3130), .A2(n3129), .ZN(n3128) );
  OR2_X1 U3876 ( .A1(n5738), .A2(n5714), .ZN(n4253) );
  CLKBUF_X1 U3877 ( .A(n5554), .Z(n5555) );
  NOR2_X1 U3878 ( .A1(n4239), .A2(n4592), .ZN(n6264) );
  OR2_X1 U3879 ( .A1(n4239), .A2(n5073), .ZN(n5738) );
  INV_X1 U3880 ( .A(n6184), .ZN(n6266) );
  NAND2_X1 U3881 ( .A1(n3006), .A2(n3444), .ZN(n4590) );
  OAI21_X1 U3882 ( .B1(n4628), .B2(n6586), .A(n5010), .ZN(n6274) );
  CLKBUF_X1 U3883 ( .A(n3416), .Z(n3417) );
  CLKBUF_X1 U3884 ( .A(n3856), .Z(n3857) );
  INV_X1 U3885 ( .A(n4768), .ZN(n4767) );
  OAI21_X1 U3886 ( .B1(n6286), .B2(n6302), .A(n6285), .ZN(n6305) );
  INV_X1 U3887 ( .A(n6346), .ZN(n6336) );
  OAI21_X1 U3888 ( .B1(n6321), .B2(n6318), .A(n6317), .ZN(n6343) );
  INV_X1 U3889 ( .A(n5775), .ZN(n5819) );
  INV_X1 U3890 ( .A(n4994), .ZN(n6350) );
  INV_X1 U3891 ( .A(n6396), .ZN(n6382) );
  AOI22_X1 U3892 ( .A1(n5872), .A2(n6404), .B1(n6279), .B2(n5867), .ZN(n5910)
         );
  INV_X1 U3893 ( .A(n6464), .ZN(n6449) );
  INV_X1 U3894 ( .A(n6453), .ZN(n6458) );
  OAI21_X1 U3895 ( .B1(n6412), .B2(n6408), .A(n6407), .ZN(n6461) );
  NOR2_X1 U3896 ( .A1(n6657), .A2(n5010), .ZN(n6419) );
  NOR2_X1 U3897 ( .A1(n4665), .A2(n5010), .ZN(n6425) );
  NOR2_X1 U3898 ( .A1(n4670), .A2(n5010), .ZN(n6431) );
  NOR2_X1 U3899 ( .A1(n4757), .A2(n5010), .ZN(n6437) );
  NOR2_X1 U3900 ( .A1(n4752), .A2(n5010), .ZN(n6443) );
  NOR2_X1 U3901 ( .A1(n4661), .A2(n5010), .ZN(n6450) );
  NOR2_X1 U3902 ( .A1(n4674), .A2(n5010), .ZN(n6460) );
  OAI22_X1 U3903 ( .A1(n4810), .A2(n4809), .B1(n5874), .B2(n5011), .ZN(n4826)
         );
  OAI21_X1 U3904 ( .B1(n4809), .B2(n4808), .A(n4807), .ZN(n4827) );
  INV_X1 U3905 ( .A(n6369), .ZN(n6400) );
  INV_X1 U3906 ( .A(n6419), .ZN(n5882) );
  INV_X1 U3907 ( .A(n6425), .ZN(n5886) );
  INV_X1 U3908 ( .A(n6431), .ZN(n5890) );
  INV_X1 U3909 ( .A(n6443), .ZN(n5898) );
  INV_X1 U3910 ( .A(n6450), .ZN(n5902) );
  OR2_X1 U3911 ( .A1(n4648), .A2(n5767), .ZN(n4928) );
  INV_X1 U3912 ( .A(n6460), .ZN(n5909) );
  NAND2_X1 U3913 ( .A1(n4531), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6502) );
  AND2_X1 U3914 ( .A1(n6490), .A2(n6489), .ZN(n6497) );
  NOR2_X1 U3915 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6510) );
  AND2_X1 U3916 ( .A1(n3901), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6511) );
  INV_X1 U3917 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6588) );
  OAI21_X1 U3918 ( .B1(n5441), .B2(n6790), .A(n4427), .ZN(n4428) );
  OR2_X1 U3919 ( .A1(n3013), .A2(n5245), .ZN(U2809) );
  OAI211_X1 U3920 ( .C1(n5518), .C2(n6790), .A(n3014), .B(n2992), .ZN(n3013)
         );
  OAI21_X1 U3921 ( .B1(n5387), .B2(n5371), .A(n4179), .ZN(U2833) );
  AND2_X1 U3922 ( .A1(n4178), .A2(n3147), .ZN(n4179) );
  OR2_X1 U3923 ( .A1(n5626), .A2(n5369), .ZN(n4178) );
  NAND2_X1 U3924 ( .A1(n4270), .A2(n4269), .ZN(U2838) );
  NAND2_X1 U3925 ( .A1(n5514), .A2(n4264), .ZN(n4270) );
  NAND2_X1 U3926 ( .A1(n3931), .A2(n6177), .ZN(n3939) );
  OAI21_X1 U3927 ( .B1(n5684), .B2(n6159), .A(n3936), .ZN(n3937) );
  NAND2_X1 U3928 ( .A1(n3913), .A2(n3912), .ZN(U2967) );
  AOI21_X1 U3929 ( .B1(n3911), .B2(n3910), .A(n3909), .ZN(n3912) );
  NAND2_X1 U3930 ( .A1(n3758), .A2(n6177), .ZN(n3913) );
  INV_X1 U3931 ( .A(n4261), .ZN(n3095) );
  CLKBUF_X3 U3933 ( .A(n3470), .Z(n4311) );
  AND2_X2 U3934 ( .A1(n4603), .A2(n5070), .ZN(n3355) );
  CLKBUF_X3 U3935 ( .A(n3355), .Z(n3356) );
  INV_X1 U3936 ( .A(n3851), .ZN(n3063) );
  NAND2_X1 U3937 ( .A1(n3109), .A2(n3108), .ZN(n5269) );
  AND2_X2 U3938 ( .A1(n4603), .A2(n4618), .ZN(n3459) );
  CLKBUF_X3 U3939 ( .A(n3459), .Z(n3362) );
  INV_X1 U3940 ( .A(n3273), .ZN(n3354) );
  CLKBUF_X3 U3941 ( .A(n3393), .Z(n4309) );
  OR2_X1 U3942 ( .A1(n2989), .A2(n3088), .ZN(n2965) );
  NAND2_X1 U3943 ( .A1(n5357), .A2(n5356), .ZN(n5258) );
  AND2_X1 U3944 ( .A1(n3858), .A2(n5372), .ZN(n2966) );
  AND2_X1 U3945 ( .A1(n3146), .A2(n3081), .ZN(n2967) );
  OAI21_X1 U3946 ( .B1(n3929), .B2(n3930), .A(n5188), .ZN(n5208) );
  AND2_X1 U3947 ( .A1(n6146), .A2(n4180), .ZN(n2968) );
  OAI211_X1 U3948 ( .C1(n5043), .C2(n3060), .A(n5582), .B(n3056), .ZN(n5581)
         );
  AND2_X1 U3949 ( .A1(n3109), .A2(n3048), .ZN(n5366) );
  OR2_X2 U3950 ( .A1(n3252), .A2(n3251), .ZN(n4237) );
  INV_X1 U3951 ( .A(n3133), .ZN(n3129) );
  INV_X1 U3952 ( .A(n5913), .ZN(n3133) );
  NOR2_X1 U3953 ( .A1(n4736), .A2(n2965), .ZN(n5055) );
  OR2_X1 U3954 ( .A1(n5362), .A2(n5262), .ZN(n5261) );
  AND2_X1 U3955 ( .A1(n3714), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n2969)
         );
  AND2_X1 U3956 ( .A1(n3018), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n2970)
         );
  AND2_X1 U3957 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n2971) );
  AND2_X1 U3958 ( .A1(n2971), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n2972)
         );
  NAND2_X2 U3959 ( .A1(n3443), .A2(n3411), .ZN(n4633) );
  OR2_X1 U3960 ( .A1(n5310), .A2(n4423), .ZN(n6029) );
  NAND2_X1 U3961 ( .A1(n3125), .A2(n3126), .ZN(n5487) );
  OR2_X1 U3962 ( .A1(n5533), .A2(n4181), .ZN(n2973) );
  INV_X1 U3963 ( .A(n3847), .ZN(n3082) );
  NOR2_X1 U3964 ( .A1(n5713), .A2(n4252), .ZN(n2974) );
  AND4_X1 U3965 ( .A1(n3164), .A2(n3163), .A3(n3162), .A4(n3161), .ZN(n2975)
         );
  NOR2_X1 U3966 ( .A1(n4266), .A2(n4265), .ZN(n2976) );
  NAND2_X1 U3967 ( .A1(n3038), .A2(n4964), .ZN(n2977) );
  AND2_X1 U3968 ( .A1(n5357), .A2(n3113), .ZN(n5259) );
  OAI21_X1 U3969 ( .B1(n3125), .B2(n3082), .A(n3066), .ZN(n4182) );
  NAND2_X1 U3970 ( .A1(n5581), .A2(n3841), .ZN(n5572) );
  NAND2_X1 U3971 ( .A1(n3846), .A2(n5552), .ZN(n5912) );
  NAND2_X1 U3972 ( .A1(n3128), .A2(n3131), .ZN(n5546) );
  NOR2_X1 U3973 ( .A1(n4266), .A2(n3093), .ZN(n5174) );
  AND2_X1 U3974 ( .A1(n3117), .A2(n4396), .ZN(n2978) );
  NAND2_X1 U3975 ( .A1(n5572), .A2(n5573), .ZN(n5562) );
  INV_X1 U3976 ( .A(n5533), .ZN(n3933) );
  NAND2_X1 U3977 ( .A1(n5161), .A2(n4062), .ZN(n5162) );
  INV_X1 U3978 ( .A(n5162), .ZN(n3044) );
  AND2_X1 U3979 ( .A1(n3011), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n2979)
         );
  NAND2_X1 U3980 ( .A1(n3759), .A2(n3354), .ZN(n3865) );
  INV_X1 U3981 ( .A(n3865), .ZN(n3270) );
  INV_X1 U3982 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3445) );
  OR2_X1 U3983 ( .A1(n3900), .A2(n4200), .ZN(n2980) );
  OR2_X1 U3984 ( .A1(n5718), .A2(n5611), .ZN(n2981) );
  AND2_X1 U3985 ( .A1(n6146), .A2(n5924), .ZN(n2982) );
  AND2_X1 U3986 ( .A1(n6146), .A2(n5640), .ZN(n2983) );
  AND2_X1 U3987 ( .A1(n3933), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n2984)
         );
  OR2_X1 U3988 ( .A1(n4258), .A2(n4247), .ZN(n2985) );
  OR2_X1 U3989 ( .A1(n3900), .A2(n4202), .ZN(n2986) );
  NAND2_X1 U3990 ( .A1(n4200), .A2(STATE2_REG_0__SCAN_IN), .ZN(n2987) );
  OR2_X1 U3991 ( .A1(n3772), .A2(n3451), .ZN(n2988) );
  OR2_X1 U3992 ( .A1(n5057), .A2(n5056), .ZN(n2989) );
  INV_X1 U3993 ( .A(n3138), .ZN(n3137) );
  NAND2_X1 U3994 ( .A1(n5473), .A2(n2973), .ZN(n3138) );
  NOR2_X1 U3995 ( .A1(n6191), .A2(n5680), .ZN(n2990) );
  NOR2_X1 U3996 ( .A1(n6146), .A2(n5740), .ZN(n2991) );
  NAND2_X1 U3997 ( .A1(n4229), .A2(n3153), .ZN(n4429) );
  OR2_X1 U3998 ( .A1(n5244), .A2(REIP_REG_18__SCAN_IN), .ZN(n2992) );
  OR2_X1 U3999 ( .A1(n4225), .A2(n5130), .ZN(n2993) );
  INV_X1 U4000 ( .A(n3289), .ZN(n3071) );
  NAND2_X1 U4001 ( .A1(n6146), .A2(n5740), .ZN(n2994) );
  AND2_X1 U4002 ( .A1(n5372), .A2(n2987), .ZN(n2995) );
  NAND2_X1 U4003 ( .A1(n6146), .A2(n3845), .ZN(n2996) );
  OR3_X2 U4004 ( .A1(n6599), .A2(n6500), .A3(n4398), .ZN(n5307) );
  INV_X1 U4005 ( .A(n5307), .ZN(n3017) );
  NOR2_X1 U4006 ( .A1(n4736), .A2(n3088), .ZN(n4966) );
  NAND2_X1 U4007 ( .A1(n3109), .A2(n3581), .ZN(n5051) );
  NAND2_X1 U4008 ( .A1(n4531), .A2(n6511), .ZN(n4558) );
  INV_X1 U4009 ( .A(n4558), .ZN(n3030) );
  NOR2_X1 U4010 ( .A1(n5362), .A2(n3098), .ZN(n5247) );
  AOI21_X1 U4011 ( .B1(n3761), .B2(n3678), .A(n3488), .ZN(n4755) );
  NAND2_X1 U4012 ( .A1(n3769), .A2(n3768), .ZN(n5085) );
  NOR2_X1 U4013 ( .A1(n4109), .A2(n4584), .ZN(n4587) );
  NAND2_X1 U4014 ( .A1(n3271), .A2(n3270), .ZN(n4084) );
  NOR2_X1 U4015 ( .A1(n5362), .A2(n3096), .ZN(n5222) );
  INV_X1 U4016 ( .A(n4736), .ZN(n4120) );
  NAND2_X1 U4017 ( .A1(n4114), .A2(n4113), .ZN(n4736) );
  AND2_X1 U4018 ( .A1(n5363), .A2(n4140), .ZN(n5359) );
  NAND2_X1 U4019 ( .A1(n4271), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n2997)
         );
  NAND2_X1 U4020 ( .A1(n3956), .A2(n2970), .ZN(n3021) );
  AND3_X1 U4021 ( .A1(n6146), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n2998) );
  OR2_X1 U4022 ( .A1(n4266), .A2(n3091), .ZN(n4376) );
  INV_X2 U4023 ( .A(n6157), .ZN(n6177) );
  INV_X1 U4024 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6755) );
  INV_X1 U4025 ( .A(n3546), .ZN(n3039) );
  AND2_X1 U4026 ( .A1(n3491), .A2(n3011), .ZN(n2999) );
  INV_X1 U4027 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3019) );
  INV_X1 U4028 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6749) );
  AND2_X1 U4029 ( .A1(n4185), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3000)
         );
  INV_X1 U4030 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3020) );
  AND2_X1 U4031 ( .A1(n6756), .A2(n5444), .ZN(n3001) );
  NOR2_X2 U4032 ( .A1(n4768), .A2(n6275), .ZN(n6303) );
  NAND2_X2 U4033 ( .A1(n6155), .A2(n3821), .ZN(n5043) );
  AOI21_X1 U4034 ( .B1(n3003), .B2(n3126), .A(n3082), .ZN(n3002) );
  NAND2_X2 U4035 ( .A1(n3846), .A2(n3127), .ZN(n3125) );
  NAND3_X1 U4036 ( .A1(n3006), .A2(n3444), .A3(n6509), .ZN(n3005) );
  INV_X1 U4037 ( .A(n3392), .ZN(n3008) );
  NAND2_X2 U4038 ( .A1(n5554), .A2(n5553), .ZN(n3846) );
  NAND3_X1 U4039 ( .A1(n3072), .A2(n3121), .A3(n2996), .ZN(n5554) );
  NAND2_X2 U4040 ( .A1(n5508), .A2(n5507), .ZN(n5506) );
  INV_X1 U4041 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3023) );
  NAND3_X1 U4042 ( .A1(n3025), .A2(n3026), .A3(n3027), .ZN(n3024) );
  NAND2_X1 U4043 ( .A1(n3858), .A2(n2995), .ZN(n3027) );
  NAND2_X2 U4044 ( .A1(n3031), .A2(n2986), .ZN(n4531) );
  INV_X1 U4045 ( .A(n4753), .ZN(n3040) );
  NAND3_X1 U4046 ( .A1(n3650), .A2(n5415), .A3(n3638), .ZN(n5414) );
  NAND2_X1 U4047 ( .A1(n5414), .A2(n3045), .ZN(n5911) );
  NAND2_X1 U4048 ( .A1(n3047), .A2(n3046), .ZN(n3045) );
  INV_X1 U4049 ( .A(n5415), .ZN(n3046) );
  NAND2_X1 U4050 ( .A1(n3109), .A2(n3049), .ZN(n3637) );
  INV_X1 U4051 ( .A(n3637), .ZN(n3635) );
  NOR2_X1 U4052 ( .A1(n3940), .A2(n3054), .ZN(n5161) );
  NAND4_X1 U4053 ( .A1(n3059), .A2(n3061), .A3(n3843), .A4(n3058), .ZN(n3072)
         );
  NAND3_X1 U4054 ( .A1(n5043), .A2(n5045), .A3(n5582), .ZN(n3059) );
  INV_X1 U4055 ( .A(n3831), .ZN(n3060) );
  NAND2_X1 U4056 ( .A1(n5044), .A2(n3831), .ZN(n5580) );
  NAND2_X1 U4057 ( .A1(n5043), .A2(n5045), .ZN(n5044) );
  AOI21_X2 U4058 ( .B1(n3062), .B2(n3847), .A(n3063), .ZN(n3066) );
  INV_X1 U4059 ( .A(n3126), .ZN(n3062) );
  NAND2_X1 U4060 ( .A1(n3275), .A2(n3286), .ZN(n4089) );
  NAND2_X1 U4061 ( .A1(n3071), .A2(n3274), .ZN(n3070) );
  OAI21_X1 U4062 ( .B1(n5506), .B2(n3075), .A(n3073), .ZN(n5486) );
  NAND2_X1 U4063 ( .A1(n5487), .A2(n2967), .ZN(n3080) );
  NAND2_X1 U4064 ( .A1(n4120), .A2(n3086), .ZN(n5276) );
  NAND2_X1 U4065 ( .A1(n5152), .A2(n4175), .ZN(n4225) );
  NAND3_X1 U4066 ( .A1(n4745), .A2(n4744), .A3(n4748), .ZN(n4746) );
  NAND2_X1 U4067 ( .A1(n3804), .A2(n3678), .ZN(n3105) );
  INV_X1 U4068 ( .A(n4755), .ZN(n3107) );
  NAND2_X1 U4069 ( .A1(n4343), .A2(n2978), .ZN(n4361) );
  AND2_X1 U4070 ( .A1(n4343), .A2(n3117), .ZN(n4395) );
  NAND2_X1 U4071 ( .A1(n4343), .A2(n3148), .ZN(n5112) );
  NAND3_X1 U4072 ( .A1(n3339), .A2(n3383), .A3(n6509), .ZN(n3425) );
  NAND2_X1 U4073 ( .A1(n3339), .A2(n3383), .ZN(n6313) );
  NAND2_X1 U4074 ( .A1(n5778), .A2(n3119), .ZN(n6357) );
  AOI22_X1 U4075 ( .A1(n5067), .A2(n3119), .B1(n3861), .B2(n5069), .ZN(n6467)
         );
  AND2_X1 U4076 ( .A1(n5866), .A2(n3119), .ZN(n4938) );
  NAND3_X1 U4077 ( .A1(n6278), .A2(n3119), .A3(n5831), .ZN(n4761) );
  AOI21_X1 U4078 ( .B1(n6404), .B2(n3119), .A(n6455), .ZN(n6411) );
  AOI21_X2 U4079 ( .B1(n3127), .B2(n3133), .A(n2991), .ZN(n3126) );
  NAND2_X1 U4080 ( .A1(n3134), .A2(n3136), .ZN(n5464) );
  NAND2_X1 U4081 ( .A1(n3154), .A2(n4580), .ZN(n3442) );
  INV_X1 U4082 ( .A(n3335), .ZN(n3338) );
  OAI22_X2 U4083 ( .A1(n4375), .A2(n4374), .B1(n3933), .B2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5508) );
  AND2_X2 U4084 ( .A1(n5068), .A2(n4600), .ZN(n3470) );
  AND2_X2 U4085 ( .A1(n4615), .A2(n4618), .ZN(n3255) );
  NOR2_X2 U4086 ( .A1(n4943), .A2(n6275), .ZN(n5907) );
  OR2_X1 U4087 ( .A1(n4648), .A2(n6275), .ZN(n4885) );
  INV_X1 U4088 ( .A(n6275), .ZN(n5767) );
  AOI21_X1 U4089 ( .B1(n6275), .B2(n4660), .A(n5874), .ZN(n4520) );
  OAI21_X1 U4090 ( .B1(n5446), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5427), 
        .ZN(n5428) );
  AOI22_X1 U4091 ( .A1(n4282), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3249) );
  XNOR2_X1 U4092 ( .A(n3443), .B(n4638), .ZN(n3763) );
  OR2_X1 U4093 ( .A1(n3410), .A2(n3409), .ZN(n3411) );
  AND2_X1 U4094 ( .A1(n3310), .A2(n3309), .ZN(n3140) );
  NAND2_X1 U4095 ( .A1(n6159), .A2(n3905), .ZN(n5576) );
  INV_X2 U4096 ( .A(n5416), .ZN(n6075) );
  INV_X1 U4097 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U4098 ( .A1(n4095), .A2(n6511), .ZN(n5337) );
  INV_X2 U4099 ( .A(n5337), .ZN(n6067) );
  INV_X1 U4100 ( .A(n6159), .ZN(n3910) );
  OR2_X1 U4101 ( .A1(n5599), .A2(n6044), .ZN(n3141) );
  INV_X1 U4102 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6409) );
  INV_X1 U4103 ( .A(n3959), .ZN(n3755) );
  OR2_X1 U4104 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3492) );
  AND2_X1 U4105 ( .A1(n3496), .A2(n3495), .ZN(n3142) );
  NOR2_X1 U4106 ( .A1(n3318), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3143)
         );
  AND3_X1 U4107 ( .A1(n3360), .A2(n3359), .A3(n3358), .ZN(n3144) );
  AND2_X1 U4108 ( .A1(n4064), .A2(n3492), .ZN(n3145) );
  OR2_X1 U4109 ( .A1(n3933), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3146)
         );
  OR2_X1 U4110 ( .A1(n6067), .A2(n4177), .ZN(n3147) );
  AND2_X1 U4111 ( .A1(n4342), .A2(n4341), .ZN(n3148) );
  AND2_X1 U4112 ( .A1(n5186), .A2(n5185), .ZN(n3149) );
  INV_X1 U4113 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5210) );
  INV_X1 U4114 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3884) );
  INV_X1 U4115 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3861) );
  INV_X1 U4116 ( .A(n5371), .ZN(n4264) );
  INV_X1 U4117 ( .A(n5462), .ZN(n4186) );
  BUF_X1 U4118 ( .A(n3763), .Z(n4637) );
  AND2_X1 U4119 ( .A1(n3760), .A2(n6605), .ZN(n3151) );
  AND4_X1 U4120 ( .A1(n3366), .A2(n3365), .A3(n3364), .A4(n3363), .ZN(n3152)
         );
  INV_X1 U4121 ( .A(n4233), .ZN(n5100) );
  OR2_X1 U4122 ( .A1(n5120), .A2(n4430), .ZN(n3153) );
  NAND2_X1 U4123 ( .A1(n4569), .A2(n4570), .ZN(n3154) );
  INV_X1 U4124 ( .A(n3848), .ZN(n3844) );
  INV_X2 U4125 ( .A(n3844), .ZN(n5533) );
  INV_X1 U4126 ( .A(n3799), .ZN(n6166) );
  AND2_X2 U4127 ( .A1(n4593), .A2(n4603), .ZN(n3345) );
  AND2_X1 U4128 ( .A1(n4937), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3863)
         );
  NOR2_X1 U4129 ( .A1(n5148), .A2(n5164), .ZN(n4340) );
  OR2_X1 U4130 ( .A1(n3481), .A2(n3480), .ZN(n3814) );
  NAND2_X1 U4131 ( .A1(n3871), .A2(n3685), .ZN(n3316) );
  AOI22_X1 U4132 ( .A1(n3340), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3162) );
  AND2_X1 U4133 ( .A1(n5127), .A2(n4340), .ZN(n4341) );
  AND4_X1 U4134 ( .A1(n5502), .A2(n5183), .A3(n5209), .A4(n5520), .ZN(n3960)
         );
  AOI21_X2 U4135 ( .B1(n3761), .B2(n3870), .A(n3151), .ZN(n3799) );
  OR2_X1 U4136 ( .A1(n6146), .A2(n3842), .ZN(n3843) );
  INV_X1 U4137 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3972) );
  AND2_X1 U4138 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3714) );
  INV_X1 U4139 ( .A(n5270), .ZN(n3596) );
  NAND2_X1 U4140 ( .A1(n6166), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3800)
         );
  NAND2_X1 U4141 ( .A1(n3425), .A2(n3374), .ZN(n3413) );
  AND2_X1 U4142 ( .A1(n3892), .A2(n3891), .ZN(n3899) );
  INV_X1 U4143 ( .A(n4192), .ZN(n4193) );
  OR2_X1 U4144 ( .A1(n5231), .A2(n3492), .ZN(n3752) );
  AND2_X1 U4145 ( .A1(n3530), .A2(n3529), .ZN(n3532) );
  NAND2_X1 U4146 ( .A1(n4282), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3235)
         );
  INV_X1 U4147 ( .A(n4354), .ZN(n4349) );
  INV_X1 U4148 ( .A(n5052), .ZN(n3581) );
  INV_X1 U4149 ( .A(n3418), .ZN(n4023) );
  AND2_X1 U4150 ( .A1(n6780), .A2(EBX_REG_29__SCAN_IN), .ZN(n4424) );
  AND2_X1 U4151 ( .A1(n4169), .A2(n4168), .ZN(n4377) );
  AND2_X1 U4152 ( .A1(n4149), .A2(n4148), .ZN(n5248) );
  AND2_X1 U4153 ( .A1(n3753), .A2(n3752), .ZN(n3959) );
  INV_X1 U4154 ( .A(n3492), .ZN(n5183) );
  INV_X1 U4155 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3535) );
  NOR2_X1 U4156 ( .A1(n5435), .A2(n5589), .ZN(n4185) );
  AND2_X1 U4157 ( .A1(n5372), .A2(n4237), .ZN(n3870) );
  INV_X1 U4158 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4613) );
  INV_X1 U4159 ( .A(n4848), .ZN(n4880) );
  OAI21_X1 U4160 ( .B1(n5782), .B2(n6588), .A(n5781), .ZN(n5813) );
  INV_X1 U4161 ( .A(n5010), .ZN(n4891) );
  OAI211_X1 U4162 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n5874), .A(n6285), .B(n5873), .ZN(n5903) );
  INV_X1 U4163 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6011) );
  AND2_X1 U4164 ( .A1(n4219), .A2(n4218), .ZN(n4564) );
  INV_X1 U4165 ( .A(n5187), .ZN(n4263) );
  INV_X1 U4166 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6673) );
  AND2_X1 U4167 ( .A1(n4975), .A2(n4974), .ZN(n6347) );
  OR2_X1 U4168 ( .A1(n4633), .A2(n4638), .ZN(n4694) );
  OR2_X1 U4169 ( .A1(n6403), .A2(n2964), .ZN(n4943) );
  INV_X1 U4170 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6397) );
  NOR2_X1 U4171 ( .A1(n4590), .A2(n5759), .ZN(n6359) );
  NAND2_X1 U4172 ( .A1(n5307), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5310) );
  INV_X1 U4173 ( .A(n6044), .ZN(n6787) );
  INV_X1 U4174 ( .A(n6029), .ZN(n6780) );
  OAI22_X1 U4175 ( .A1(n5663), .A2(n5369), .B1(n5204), .B2(n6067), .ZN(n4268)
         );
  INV_X1 U4176 ( .A(n5369), .ZN(n6065) );
  AND2_X1 U4177 ( .A1(n5416), .A2(n4567), .ZN(n6073) );
  INV_X1 U4178 ( .A(n6114), .ZN(n6098) );
  INV_X1 U4179 ( .A(n6125), .ZN(n6122) );
  NOR2_X1 U4180 ( .A1(n5695), .A2(n4257), .ZN(n5667) );
  NAND2_X1 U4181 ( .A1(n2974), .A2(n4253), .ZN(n5919) );
  OAI21_X1 U4182 ( .B1(n4847), .B2(n4846), .A(n4845), .ZN(n4887) );
  OAI22_X1 U4183 ( .A1(n6321), .A2(n6320), .B1(n6319), .B2(n6409), .ZN(n6342)
         );
  OAI21_X1 U4184 ( .B1(n4700), .B2(n4699), .A(n4698), .ZN(n4723) );
  OR4_X1 U4185 ( .A1(n4972), .A2(n6279), .A3(n5868), .A4(n4971), .ZN(n6351) );
  INV_X1 U4186 ( .A(n4694), .ZN(n5822) );
  OAI211_X1 U4187 ( .C1(n5829), .C2(n5828), .A(n5827), .B(n5826), .ZN(n5856)
         );
  OAI21_X1 U4188 ( .B1(n4942), .B2(n4940), .A(n4939), .ZN(n4959) );
  AND2_X1 U4189 ( .A1(n6277), .A2(n5866), .ZN(n6404) );
  INV_X1 U4190 ( .A(n6308), .ZN(n6457) );
  NAND3_X1 U4191 ( .A1(n5013), .A2(n5827), .A3(n5012), .ZN(n5036) );
  NOR2_X2 U4192 ( .A1(n4811), .A2(n5767), .ZN(n5040) );
  NOR2_X1 U4193 ( .A1(n6749), .A2(n5874), .ZN(n4627) );
  INV_X1 U4194 ( .A(n6573), .ZN(n6575) );
  NAND2_X1 U4195 ( .A1(n4456), .A2(n4453), .ZN(n6599) );
  INV_X1 U4196 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6604) );
  INV_X1 U4197 ( .A(n6615), .ZN(n6598) );
  OR2_X1 U4198 ( .A1(n5310), .A2(n4435), .ZN(n6044) );
  AND2_X1 U4199 ( .A1(n6790), .A2(n5298), .ZN(n6051) );
  INV_X1 U4200 ( .A(n4268), .ZN(n4269) );
  INV_X1 U4201 ( .A(n5514), .ZN(n5402) );
  INV_X1 U4202 ( .A(n5569), .ZN(n5425) );
  NAND2_X1 U4203 ( .A1(n6125), .A2(n4565), .ZN(n5416) );
  OR2_X1 U4204 ( .A1(n6114), .A2(n4681), .ZN(n6079) );
  OR2_X1 U4205 ( .A1(n6098), .A2(n6601), .ZN(n6108) );
  OR2_X1 U4206 ( .A1(n4558), .A2(n6492), .ZN(n6142) );
  INV_X1 U4207 ( .A(n3937), .ZN(n3938) );
  OR2_X2 U4208 ( .A1(n5565), .A2(n4522), .ZN(n6182) );
  OR2_X1 U4209 ( .A1(n6516), .A2(n6406), .ZN(n6157) );
  AND2_X1 U4210 ( .A1(n4382), .A2(n4381), .ZN(n4383) );
  INV_X1 U4211 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4937) );
  INV_X1 U4212 ( .A(n4765), .ZN(n4803) );
  OR2_X1 U4213 ( .A1(n4637), .A2(n6276), .ZN(n6346) );
  OR2_X1 U4214 ( .A1(n4637), .A2(n5768), .ZN(n6339) );
  AOI22_X1 U4215 ( .A1(n4697), .A2(n4699), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4693), .ZN(n4726) );
  NAND2_X1 U4216 ( .A1(n5822), .A2(n5821), .ZN(n6385) );
  NAND2_X1 U4217 ( .A1(n5822), .A2(n4969), .ZN(n6396) );
  NAND2_X1 U4218 ( .A1(n4935), .A2(n6275), .ZN(n5862) );
  INV_X1 U4219 ( .A(n6437), .ZN(n5894) );
  OR2_X1 U4220 ( .A1(n6403), .A2(n5863), .ZN(n6464) );
  OR2_X1 U4221 ( .A1(n6403), .A2(n5006), .ZN(n6453) );
  OR2_X1 U4222 ( .A1(n4811), .A2(n6275), .ZN(n4927) );
  NOR2_X1 U4223 ( .A1(n4895), .A2(n4894), .ZN(n4934) );
  INV_X1 U4224 ( .A(n6585), .ZN(n6581) );
  INV_X1 U4225 ( .A(READY_N), .ZN(n6606) );
  INV_X1 U4226 ( .A(n6567), .ZN(n6577) );
  NAND2_X1 U4227 ( .A1(n4436), .A2(n3141), .ZN(U2798) );
  OAI21_X1 U4228 ( .B1(n5377), .B2(n5371), .A(n4373), .ZN(U2829) );
  NAND2_X1 U4229 ( .A1(n3939), .A2(n3938), .ZN(U2966) );
  AND2_X4 U4230 ( .A1(n5068), .A2(n4615), .ZN(n4282) );
  AOI22_X1 U4231 ( .A1(n4282), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3159) );
  AND2_X2 U4232 ( .A1(n3445), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4603)
         );
  INV_X1 U4233 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3856) );
  AND2_X2 U4234 ( .A1(n4600), .A2(n4618), .ZN(n3254) );
  AOI22_X1 U4235 ( .A1(n3345), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3158) );
  AND2_X2 U4236 ( .A1(n4600), .A2(n5070), .ZN(n3361) );
  AND2_X4 U4237 ( .A1(n5068), .A2(n3160), .ZN(n3453) );
  AOI22_X1 U4238 ( .A1(n3361), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3453), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3157) );
  AOI22_X1 U4239 ( .A1(n3470), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3156) );
  AOI22_X1 U4240 ( .A1(n3355), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4283), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3164) );
  AND2_X4 U4241 ( .A1(n5068), .A2(n4603), .ZN(n3475) );
  AOI22_X1 U4242 ( .A1(n3475), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3163) );
  AOI22_X1 U4243 ( .A1(n3398), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3357), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3161) );
  AOI22_X1 U4244 ( .A1(n3345), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3168) );
  AOI22_X1 U4245 ( .A1(n3470), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3167) );
  NAND4_X1 U4246 ( .A1(n3169), .A2(n3168), .A3(n3167), .A4(n3166), .ZN(n3175)
         );
  AOI22_X1 U4247 ( .A1(n3355), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4283), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3172) );
  AOI22_X1 U4248 ( .A1(n3475), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3171) );
  NAND4_X1 U4249 ( .A1(n3173), .A2(n3172), .A3(n3171), .A4(n3170), .ZN(n3174)
         );
  OR2_X2 U4250 ( .A1(n3175), .A2(n3174), .ZN(n3286) );
  NAND2_X1 U4251 ( .A1(n3759), .A2(n3286), .ZN(n3186) );
  AOI22_X1 U4252 ( .A1(n3355), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3178) );
  AOI22_X1 U4253 ( .A1(n3357), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3177) );
  AOI22_X1 U4254 ( .A1(n3340), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3176) );
  AOI22_X1 U4255 ( .A1(n3345), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3453), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3183) );
  AOI22_X1 U4256 ( .A1(n3393), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3182) );
  AOI22_X1 U4257 ( .A1(n3475), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3398), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U4258 ( .A1(n3470), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4283), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3180) );
  INV_X2 U4259 ( .A(n3284), .ZN(n4069) );
  NAND2_X1 U4260 ( .A1(n3186), .A2(n4069), .ZN(n3188) );
  NAND2_X1 U4261 ( .A1(n3759), .A2(n3284), .ZN(n3187) );
  NAND2_X1 U4262 ( .A1(n3188), .A2(n3187), .ZN(n3222) );
  NAND2_X1 U4263 ( .A1(n4282), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3192)
         );
  NAND2_X1 U4264 ( .A1(n3355), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3191) );
  NAND2_X1 U4265 ( .A1(n3345), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3190) );
  NAND2_X1 U4266 ( .A1(n4283), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3189) );
  NAND2_X1 U4267 ( .A1(n3361), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3196)
         );
  NAND2_X1 U4268 ( .A1(n3453), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3195) );
  NAND2_X1 U4269 ( .A1(n3393), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3194)
         );
  NAND2_X1 U4270 ( .A1(n3254), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3193) );
  NAND2_X1 U4271 ( .A1(n3398), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3200) );
  NAND2_X1 U4272 ( .A1(n3475), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3199) );
  NAND2_X1 U4273 ( .A1(n3357), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3198)
         );
  NAND2_X1 U4274 ( .A1(n3255), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3197)
         );
  NAND2_X1 U4275 ( .A1(n3470), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3204) );
  NAND2_X1 U4276 ( .A1(n3459), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3203) );
  NAND2_X1 U4277 ( .A1(n3340), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3201) );
  NAND2_X1 U4278 ( .A1(n3273), .A2(n3284), .ZN(n3219) );
  AOI22_X1 U4279 ( .A1(n3361), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3212) );
  AOI22_X1 U4280 ( .A1(n3393), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3211) );
  AOI22_X1 U4281 ( .A1(n3255), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3210) );
  AOI22_X1 U4282 ( .A1(n3453), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3215) );
  AOI22_X1 U4283 ( .A1(n3475), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3214) );
  AOI22_X1 U4284 ( .A1(n3357), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4283), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3213) );
  AOI22_X1 U4285 ( .A1(n3470), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4282), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3216) );
  OAI211_X1 U4286 ( .C1(n3286), .C2(n3273), .A(n3219), .B(n4566), .ZN(n3220)
         );
  INV_X1 U4287 ( .A(n3220), .ZN(n3221) );
  NAND2_X1 U4288 ( .A1(n3222), .A2(n3221), .ZN(n3288) );
  NAND2_X1 U4289 ( .A1(n3355), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3226) );
  NAND2_X1 U4290 ( .A1(n3398), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3225) );
  NAND2_X1 U4291 ( .A1(n3357), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3224)
         );
  NAND2_X1 U4292 ( .A1(n4283), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3223) );
  NAND2_X1 U4293 ( .A1(n3475), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3230) );
  NAND2_X1 U4294 ( .A1(n3255), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3229)
         );
  NAND2_X1 U4295 ( .A1(n3340), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3228) );
  NAND2_X1 U4296 ( .A1(n3346), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3227)
         );
  NAND2_X1 U4297 ( .A1(n3393), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3236)
         );
  NAND2_X1 U4298 ( .A1(n3470), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3234) );
  NAND2_X1 U4299 ( .A1(n3459), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3233) );
  NAND2_X1 U4300 ( .A1(n3361), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3240)
         );
  NAND2_X1 U4301 ( .A1(n3345), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3239) );
  NAND2_X1 U4302 ( .A1(n3254), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3238) );
  NAND2_X1 U4303 ( .A1(n3453), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3237) );
  NAND3_X4 U4304 ( .A1(n3242), .A2(n3241), .A3(n3150), .ZN(n4090) );
  NAND2_X1 U4305 ( .A1(n3288), .A2(n4681), .ZN(n3268) );
  AOI22_X1 U4306 ( .A1(n3453), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3246) );
  AOI22_X1 U4307 ( .A1(n3470), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3357), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3245) );
  AOI22_X1 U4308 ( .A1(n3475), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3398), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3244) );
  AOI22_X1 U4309 ( .A1(n3340), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3243) );
  NAND4_X1 U4310 ( .A1(n3246), .A2(n3245), .A3(n3244), .A4(n3243), .ZN(n3252)
         );
  AOI22_X1 U4311 ( .A1(n3361), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3250) );
  AOI22_X1 U4312 ( .A1(n3459), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4283), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3248) );
  AOI22_X1 U4313 ( .A1(n3355), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3247) );
  NAND4_X1 U4314 ( .A1(n3250), .A2(n3249), .A3(n3248), .A4(n3247), .ZN(n3251)
         );
  INV_X1 U4315 ( .A(n4090), .ZN(n3266) );
  AOI22_X1 U4316 ( .A1(n3254), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4283), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3259) );
  AOI22_X1 U4317 ( .A1(n3355), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3357), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3258) );
  AOI22_X1 U4318 ( .A1(n3345), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3453), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4319 ( .A1(n3255), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3256) );
  NAND4_X1 U4320 ( .A1(n3259), .A2(n3258), .A3(n3257), .A4(n3256), .ZN(n3265)
         );
  AOI22_X1 U4321 ( .A1(n3361), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4282), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U4322 ( .A1(n3470), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3262) );
  AOI22_X1 U4323 ( .A1(n3398), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3261) );
  AOI22_X1 U4324 ( .A1(n3475), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3260) );
  NAND4_X1 U4325 ( .A1(n3263), .A2(n3262), .A3(n3261), .A4(n3260), .ZN(n3264)
         );
  NAND2_X1 U4326 ( .A1(n3774), .A2(n3289), .ZN(n3267) );
  AND3_X2 U4327 ( .A1(n3268), .A2(n5309), .A3(n3267), .ZN(n3311) );
  AND2_X1 U4328 ( .A1(n3354), .A2(n4566), .ZN(n3269) );
  NAND2_X1 U4329 ( .A1(n4073), .A2(n3303), .ZN(n3272) );
  INV_X1 U4330 ( .A(n3273), .ZN(n3274) );
  XNOR2_X1 U4331 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n4195) );
  NAND2_X1 U4332 ( .A1(n3253), .A2(n4195), .ZN(n3283) );
  INV_X1 U4333 ( .A(n3786), .ZN(n4078) );
  NAND4_X1 U4334 ( .A1(n3311), .A2(n3309), .A3(n3902), .A4(n3276), .ZN(n3277)
         );
  NAND2_X1 U4335 ( .A1(n3277), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3320) );
  NAND2_X1 U4336 ( .A1(n3320), .A2(n3316), .ZN(n3385) );
  NAND2_X1 U4337 ( .A1(n3385), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3294) );
  NAND2_X1 U4338 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3387) );
  OAI21_X1 U4339 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n3387), .ZN(n5008) );
  OR2_X1 U4340 ( .A1(n3904), .A2(n5008), .ZN(n3280) );
  INV_X1 U4341 ( .A(n3901), .ZN(n6493) );
  NAND2_X1 U4342 ( .A1(n6493), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3279) );
  INV_X1 U4343 ( .A(n3283), .ZN(n3292) );
  INV_X1 U4344 ( .A(n5297), .ZN(n4218) );
  AND2_X1 U4345 ( .A1(n4092), .A2(n3275), .ZN(n3285) );
  NAND2_X1 U4346 ( .A1(n4218), .A2(n3285), .ZN(n4082) );
  INV_X1 U4347 ( .A(n4082), .ZN(n3287) );
  NAND2_X1 U4348 ( .A1(n3287), .A2(n4233), .ZN(n4216) );
  INV_X1 U4349 ( .A(n3288), .ZN(n3291) );
  NAND2_X1 U4350 ( .A1(n3289), .A2(n4077), .ZN(n3304) );
  NOR2_X1 U4351 ( .A1(n3865), .A2(n4090), .ZN(n3290) );
  AND3_X2 U4352 ( .A1(n3291), .A2(n3304), .A3(n3290), .ZN(n4192) );
  NAND2_X2 U4353 ( .A1(n4192), .A2(n4656), .ZN(n5927) );
  OAI211_X1 U4354 ( .C1(n4444), .C2(n3292), .A(n4216), .B(n5927), .ZN(n3293)
         );
  NAND2_X1 U4355 ( .A1(n3293), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3298) );
  NAND3_X1 U4356 ( .A1(n3294), .A2(n3295), .A3(n3298), .ZN(n3381) );
  INV_X1 U4358 ( .A(n3295), .ZN(n3296) );
  NOR2_X1 U4359 ( .A1(n3296), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3297)
         );
  OR2_X2 U4360 ( .A1(n3298), .A2(n3297), .ZN(n3382) );
  NAND2_X1 U4361 ( .A1(n3685), .A2(n3273), .ZN(n3300) );
  NAND2_X1 U4362 ( .A1(n3300), .A2(n4077), .ZN(n3301) );
  OAI21_X1 U4363 ( .B1(n3302), .B2(n3301), .A(n4237), .ZN(n3306) );
  NAND2_X1 U4364 ( .A1(n3304), .A2(n3303), .ZN(n3305) );
  AND2_X1 U4365 ( .A1(n3306), .A2(n3305), .ZN(n3315) );
  AND2_X1 U4366 ( .A1(n4092), .A2(n4681), .ZN(n4083) );
  NAND2_X1 U4367 ( .A1(n6510), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3308) );
  AOI21_X1 U4368 ( .B1(n4083), .B2(n4660), .A(n3308), .ZN(n3310) );
  INV_X1 U4369 ( .A(n3311), .ZN(n3314) );
  NAND2_X1 U4370 ( .A1(n3270), .A2(n4237), .ZN(n3313) );
  AND2_X1 U4371 ( .A1(n4212), .A2(n4090), .ZN(n3312) );
  NAND3_X1 U4372 ( .A1(n3315), .A2(n3140), .A3(n4081), .ZN(n3335) );
  MUX2_X1 U4373 ( .A(n3904), .B(n3901), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3317) );
  AND2_X1 U4374 ( .A1(n3316), .A2(n3317), .ZN(n3319) );
  INV_X1 U4375 ( .A(n3317), .ZN(n3318) );
  AOI21_X2 U4376 ( .B1(n3320), .B2(n3319), .A(n3143), .ZN(n3336) );
  NAND2_X1 U4377 ( .A1(n3335), .A2(n3336), .ZN(n3383) );
  XNOR2_X2 U4378 ( .A(n3322), .B(n3321), .ZN(n5865) );
  NAND2_X1 U4379 ( .A1(n5865), .A2(n6509), .ZN(n3334) );
  INV_X1 U4380 ( .A(n3451), .ZN(n3376) );
  AOI22_X1 U4381 ( .A1(n3469), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3453), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4382 ( .A1(n4309), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U4383 ( .A1(n3499), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4384 ( .A1(n4288), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3323) );
  NAND4_X1 U4385 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), .ZN(n3332)
         );
  AOI22_X1 U4386 ( .A1(n3361), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4310), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4387 ( .A1(n3356), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3329) );
  AOI22_X1 U4388 ( .A1(n4311), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3328) );
  AOI22_X1 U4389 ( .A1(n4317), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3327) );
  NAND4_X1 U4390 ( .A1(n3330), .A2(n3329), .A3(n3328), .A4(n3327), .ZN(n3331)
         );
  NAND2_X1 U4391 ( .A1(n3376), .A2(n3785), .ZN(n3333) );
  NAND2_X2 U4392 ( .A1(n3334), .A2(n3333), .ZN(n3415) );
  INV_X1 U4393 ( .A(n3336), .ZN(n3337) );
  NAND2_X1 U4394 ( .A1(n3338), .A2(n3337), .ZN(n3339) );
  INV_X1 U4395 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4396 ( .A1(n4308), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3453), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3344) );
  AOI22_X1 U4397 ( .A1(n4311), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4310), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3343) );
  AOI22_X1 U4398 ( .A1(n3398), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3342) );
  AOI22_X1 U4399 ( .A1(n3499), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3341) );
  NAND4_X1 U4400 ( .A1(n3344), .A2(n3343), .A3(n3342), .A4(n3341), .ZN(n3353)
         );
  AOI22_X1 U4401 ( .A1(n3469), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3351) );
  AOI22_X1 U4402 ( .A1(n4309), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3350) );
  AOI22_X1 U4403 ( .A1(n3356), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3349) );
  INV_X1 U4404 ( .A(n3346), .ZN(n3347) );
  AOI22_X1 U4405 ( .A1(n3357), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n2961), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3348) );
  NAND4_X1 U4406 ( .A1(n3351), .A2(n3350), .A3(n3349), .A4(n3348), .ZN(n3352)
         );
  AOI21_X1 U4407 ( .B1(n4681), .B2(n3784), .A(n6509), .ZN(n3368) );
  AOI22_X1 U4408 ( .A1(n3499), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4409 ( .A1(n3356), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4410 ( .A1(n4288), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n2961), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4411 ( .A1(n3398), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3357), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4412 ( .A1(n3361), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3453), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4413 ( .A1(n3469), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3365) );
  AOI22_X1 U4414 ( .A1(n4282), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4415 ( .A1(n4311), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3363) );
  INV_X1 U4416 ( .A(n3837), .ZN(n3375) );
  NAND2_X1 U4417 ( .A1(n3375), .A2(n3274), .ZN(n3370) );
  NAND2_X1 U4418 ( .A1(n3424), .A2(n3426), .ZN(n3429) );
  INV_X1 U4419 ( .A(n3832), .ZN(n3372) );
  NAND2_X1 U4420 ( .A1(n3372), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3373) );
  INV_X1 U4421 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3379) );
  NAND2_X1 U4422 ( .A1(n3376), .A2(n3375), .ZN(n3378) );
  INV_X1 U4423 ( .A(n3452), .ZN(n3406) );
  NAND2_X1 U4424 ( .A1(n3406), .A2(n3785), .ZN(n3377) );
  OAI211_X1 U4425 ( .C1(n3888), .C2(n3379), .A(n3378), .B(n3377), .ZN(n3412)
         );
  AND2_X2 U4426 ( .A1(n3415), .A2(n3380), .ZN(n3409) );
  INV_X1 U4427 ( .A(n3381), .ZN(n3384) );
  OAI21_X2 U4428 ( .B1(n3384), .B2(n3383), .A(n3382), .ZN(n3392) );
  INV_X1 U4430 ( .A(n3387), .ZN(n3386) );
  NAND2_X1 U4431 ( .A1(n3386), .A2(n6474), .ZN(n6398) );
  NAND2_X1 U4432 ( .A1(n3387), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3388) );
  OAI22_X1 U4433 ( .A1(n4849), .A2(n3904), .B1(n3901), .B2(n6474), .ZN(n3389)
         );
  INV_X1 U4434 ( .A(n3390), .ZN(n3391) );
  NAND2_X1 U4435 ( .A1(n3392), .A2(n3391), .ZN(n3444) );
  AOI22_X1 U4436 ( .A1(n4308), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3453), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3397) );
  AOI22_X1 U4437 ( .A1(n3469), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3396) );
  AOI22_X1 U4438 ( .A1(n4282), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3395) );
  INV_X1 U4439 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n6655) );
  AOI22_X1 U4440 ( .A1(n4311), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3394) );
  NAND4_X1 U4441 ( .A1(n3397), .A2(n3396), .A3(n3395), .A4(n3394), .ZN(n3404)
         );
  AOI22_X1 U4442 ( .A1(n4317), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3402) );
  AOI22_X1 U4443 ( .A1(n3356), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3401) );
  AOI22_X1 U4444 ( .A1(n3499), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4445 ( .A1(n4288), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3399) );
  NAND4_X1 U4446 ( .A1(n3402), .A2(n3401), .A3(n3400), .A4(n3399), .ZN(n3403)
         );
  XNOR2_X1 U4447 ( .A(n3408), .B(n3407), .ZN(n3410) );
  NOR2_X1 U4448 ( .A1(n4633), .A2(n3627), .ZN(n3440) );
  NAND2_X1 U4449 ( .A1(n5874), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4021) );
  NOR2_X1 U4450 ( .A1(n3440), .A2(n4384), .ZN(n4581) );
  XNOR2_X1 U4451 ( .A(n3413), .B(n3412), .ZN(n3414) );
  NAND2_X1 U4452 ( .A1(n4635), .A2(n3678), .ZN(n3423) );
  AND2_X1 U4453 ( .A1(n4233), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3436) );
  INV_X1 U4454 ( .A(n3436), .ZN(n3494) );
  NOR2_X2 U4455 ( .A1(n4566), .A2(n5874), .ZN(n3418) );
  NAND2_X1 U4456 ( .A1(n4357), .A2(EAX_REG_1__SCAN_IN), .ZN(n3420) );
  NAND2_X1 U4457 ( .A1(n6409), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3419)
         );
  OAI211_X1 U4458 ( .C1(n3494), .C2(n3417), .A(n3420), .B(n3419), .ZN(n3421)
         );
  INV_X1 U4459 ( .A(n3421), .ZN(n3422) );
  NAND2_X1 U4460 ( .A1(n3423), .A2(n3422), .ZN(n4569) );
  NAND2_X1 U4461 ( .A1(n3425), .A2(n3424), .ZN(n3428) );
  AOI22_X1 U4462 ( .A1(n3418), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6409), .ZN(n3432) );
  NAND2_X1 U4463 ( .A1(n3436), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3431) );
  OAI211_X1 U4464 ( .C1(n6313), .C2(n3627), .A(n3432), .B(n3431), .ZN(n4519)
         );
  INV_X1 U4465 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3434) );
  OAI21_X1 U4466 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3486), .ZN(n6181) );
  NAND2_X1 U4467 ( .A1(n5183), .A2(n6181), .ZN(n3433) );
  OAI21_X1 U4468 ( .B1(n4021), .B2(n3434), .A(n3433), .ZN(n3435) );
  AOI21_X1 U4469 ( .B1(n4357), .B2(EAX_REG_2__SCAN_IN), .A(n3435), .ZN(n3438)
         );
  NAND2_X1 U4470 ( .A1(n3436), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3437) );
  AND2_X1 U4471 ( .A1(n3438), .A2(n3437), .ZN(n4580) );
  INV_X1 U4472 ( .A(n4580), .ZN(n3439) );
  OR2_X1 U4473 ( .A1(n3440), .A2(n3439), .ZN(n3441) );
  INV_X1 U4474 ( .A(n3443), .ZN(n3468) );
  NAND2_X1 U4475 ( .A1(n3446), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3450) );
  INV_X1 U4476 ( .A(n3904), .ZN(n3448) );
  NAND3_X1 U4477 ( .A1(n6397), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6364) );
  INV_X1 U4478 ( .A(n6364), .ZN(n6363) );
  NAND2_X1 U4479 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6363), .ZN(n6354) );
  NAND2_X1 U4480 ( .A1(n6397), .A2(n6354), .ZN(n3447) );
  NAND3_X1 U4481 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4890) );
  INV_X1 U4482 ( .A(n4890), .ZN(n4651) );
  NAND2_X1 U4483 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4651), .ZN(n4685) );
  AOI22_X1 U4484 ( .A1(n3448), .A2(n5009), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6493), .ZN(n3449) );
  AOI22_X1 U4485 ( .A1(n4308), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3453), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3458) );
  AOI22_X1 U4486 ( .A1(n4282), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3457) );
  AOI22_X1 U4487 ( .A1(n3356), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3456) );
  AOI22_X1 U4488 ( .A1(n4317), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4288), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3455) );
  NAND4_X1 U4489 ( .A1(n3458), .A2(n3457), .A3(n3456), .A4(n3455), .ZN(n3465)
         );
  AOI22_X1 U4490 ( .A1(n4311), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3463) );
  AOI22_X1 U4491 ( .A1(n3362), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3462) );
  AOI22_X1 U4492 ( .A1(n4316), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3461) );
  AOI22_X1 U4493 ( .A1(n3499), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3460) );
  NAND4_X1 U4494 ( .A1(n3463), .A2(n3462), .A3(n3461), .A4(n3460), .ZN(n3464)
         );
  AOI22_X1 U4495 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n3871), .B1(n3893), 
        .B2(n3764), .ZN(n3466) );
  NAND2_X1 U4496 ( .A1(n3468), .A2(n4638), .ZN(n3498) );
  INV_X1 U4497 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4498 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4308), .B1(n3453), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3474) );
  INV_X1 U4499 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6750) );
  AOI22_X1 U4500 ( .A1(n3469), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4501 ( .A1(n4310), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4502 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4311), .B1(n3362), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3471) );
  NAND4_X1 U4503 ( .A1(n3474), .A2(n3473), .A3(n3472), .A4(n3471), .ZN(n3481)
         );
  AOI22_X1 U4504 ( .A1(n4317), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4505 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3356), .B1(n4318), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4506 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3499), .B1(n3569), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3477) );
  AOI22_X1 U4507 ( .A1(n4288), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3476) );
  NAND4_X1 U4508 ( .A1(n3479), .A2(n3478), .A3(n3477), .A4(n3476), .ZN(n3480)
         );
  NAND2_X1 U4509 ( .A1(n3893), .A2(n3814), .ZN(n3482) );
  NAND2_X1 U4510 ( .A1(n5874), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3485)
         );
  NAND2_X1 U4511 ( .A1(n4357), .A2(EAX_REG_4__SCAN_IN), .ZN(n3484) );
  OAI211_X1 U4512 ( .C1(n3494), .C2(n3884), .A(n3485), .B(n3484), .ZN(n3487)
         );
  OAI21_X1 U4513 ( .B1(n3491), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3536), 
        .ZN(n6172) );
  MUX2_X1 U4514 ( .A(n3487), .B(n6172), .S(n5183), .Z(n3488) );
  NAND2_X1 U4515 ( .A1(n3763), .A2(n3678), .ZN(n3497) );
  NOR2_X1 U4516 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3489), .ZN(n3490)
         );
  NOR2_X1 U4517 ( .A1(n3491), .A2(n3490), .ZN(n6055) );
  INV_X1 U4518 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6046) );
  OAI22_X1 U4519 ( .A1(n6055), .A2(n3492), .B1(n4021), .B2(n6046), .ZN(n3493)
         );
  AOI21_X1 U4520 ( .B1(n4357), .B2(EAX_REG_3__SCAN_IN), .A(n3493), .ZN(n3496)
         );
  NAND2_X1 U4521 ( .A1(n3436), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3495) );
  NAND2_X1 U4522 ( .A1(n3497), .A2(n3142), .ZN(n4583) );
  INV_X1 U4523 ( .A(n3498), .ZN(n3518) );
  NAND2_X1 U4524 ( .A1(n3518), .A2(n3515), .ZN(n3512) );
  INV_X1 U4525 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U4526 ( .A1(n4308), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3503) );
  AOI22_X1 U4527 ( .A1(n4316), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3502) );
  AOI22_X1 U4528 ( .A1(n3499), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3501) );
  INV_X2 U4529 ( .A(n3347), .ZN(n4319) );
  AOI22_X1 U4530 ( .A1(n4288), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3500) );
  NAND4_X1 U4531 ( .A1(n3503), .A2(n3502), .A3(n3501), .A4(n3500), .ZN(n3509)
         );
  AOI22_X1 U4532 ( .A1(n4310), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3453), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3507) );
  AOI22_X1 U4533 ( .A1(n4311), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3506) );
  AOI22_X1 U4534 ( .A1(n3362), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3505) );
  AOI22_X1 U4535 ( .A1(n3356), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3504) );
  NAND4_X1 U4536 ( .A1(n3507), .A2(n3506), .A3(n3505), .A4(n3504), .ZN(n3508)
         );
  NAND2_X1 U4537 ( .A1(n3893), .A2(n3813), .ZN(n3510) );
  XNOR2_X1 U4538 ( .A(n3536), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5300) );
  OAI22_X1 U4539 ( .A1(n5300), .A2(n3492), .B1(n4021), .B2(n3535), .ZN(n3513)
         );
  AOI21_X1 U4540 ( .B1(n4357), .B2(EAX_REG_5__SCAN_IN), .A(n3513), .ZN(n3514)
         );
  NAND2_X1 U4541 ( .A1(n3518), .A2(n3517), .ZN(n3533) );
  AOI22_X1 U4542 ( .A1(n4308), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3453), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4543 ( .A1(n3469), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3521) );
  AOI22_X1 U4544 ( .A1(n4310), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3520) );
  AOI22_X1 U4545 ( .A1(n4311), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3519) );
  NAND4_X1 U4546 ( .A1(n3522), .A2(n3521), .A3(n3520), .A4(n3519), .ZN(n3528)
         );
  INV_X1 U4547 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n6703) );
  AOI22_X1 U4548 ( .A1(n4317), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3526) );
  AOI22_X1 U4549 ( .A1(n3356), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3525) );
  AOI22_X1 U4550 ( .A1(n3499), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3524) );
  AOI22_X1 U4551 ( .A1(n4288), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3523) );
  NAND4_X1 U4552 ( .A1(n3526), .A2(n3525), .A3(n3524), .A4(n3523), .ZN(n3527)
         );
  NAND2_X1 U4553 ( .A1(n3893), .A2(n3824), .ZN(n3530) );
  NAND2_X1 U4554 ( .A1(n3871), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3529) );
  NAND2_X1 U4555 ( .A1(n3533), .A2(n3532), .ZN(n3534) );
  OR2_X1 U4556 ( .A1(n2999), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3537) );
  NAND2_X1 U4557 ( .A1(n3557), .A2(n3537), .ZN(n6163) );
  INV_X1 U4558 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4754) );
  INV_X1 U4559 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3538) );
  OAI22_X1 U4560 ( .A1(n4023), .A2(n4754), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3538), .ZN(n3539) );
  MUX2_X1 U4561 ( .A(n6163), .B(n3539), .S(n3492), .Z(n3540) );
  AOI21_X2 U4562 ( .B1(n3812), .B2(n3678), .A(n3540), .ZN(n4753) );
  INV_X1 U4563 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3542) );
  NAND2_X1 U4564 ( .A1(n3893), .A2(n3837), .ZN(n3541) );
  OAI21_X1 U4565 ( .B1(n3542), .B2(n3888), .A(n3541), .ZN(n3543) );
  INV_X1 U4566 ( .A(EAX_REG_7__SCAN_IN), .ZN(n5050) );
  XNOR2_X1 U4567 ( .A(n3557), .B(n6011), .ZN(n6008) );
  NAND2_X1 U4568 ( .A1(n6008), .A2(n5183), .ZN(n3545) );
  NAND2_X1 U4569 ( .A1(n4384), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3544)
         );
  OAI211_X1 U4570 ( .C1(n4023), .C2(n5050), .A(n3545), .B(n3544), .ZN(n3546)
         );
  AOI22_X1 U4571 ( .A1(n4308), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4572 ( .A1(n4282), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4573 ( .A1(n4316), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4574 ( .A1(n3569), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4288), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3547) );
  NAND4_X1 U4575 ( .A1(n3550), .A2(n3549), .A3(n3548), .A4(n3547), .ZN(n3556)
         );
  AOI22_X1 U4576 ( .A1(n4307), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4577 ( .A1(n3356), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4578 ( .A1(n4311), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3552) );
  AOI22_X1 U4579 ( .A1(n3499), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3551) );
  NAND4_X1 U4580 ( .A1(n3554), .A2(n3553), .A3(n3552), .A4(n3551), .ZN(n3555)
         );
  NOR2_X1 U4581 ( .A1(n3556), .A2(n3555), .ZN(n3564) );
  NAND2_X1 U4582 ( .A1(n3558), .A2(n6706), .ZN(n3560) );
  INV_X1 U4583 ( .A(n3592), .ZN(n3559) );
  NAND2_X1 U4584 ( .A1(n3560), .A2(n3559), .ZN(n5584) );
  NOR2_X1 U4585 ( .A1(n4021), .A2(n6706), .ZN(n3561) );
  AOI21_X1 U4586 ( .B1(n5584), .B2(n5183), .A(n3561), .ZN(n3563) );
  NAND2_X1 U4587 ( .A1(n3418), .A2(EAX_REG_8__SCAN_IN), .ZN(n3562) );
  OAI211_X1 U4588 ( .C1(n3627), .C2(n3564), .A(n3563), .B(n3562), .ZN(n4964)
         );
  INV_X1 U4589 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6001) );
  XNOR2_X1 U4590 ( .A(n6001), .B(n3592), .ZN(n5996) );
  INV_X1 U4591 ( .A(n5996), .ZN(n3580) );
  AOI22_X1 U4592 ( .A1(n4308), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4593 ( .A1(n4311), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3567) );
  AOI22_X1 U4594 ( .A1(n4317), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4595 ( .A1(n3499), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3565) );
  NAND4_X1 U4596 ( .A1(n3568), .A2(n3567), .A3(n3566), .A4(n3565), .ZN(n3575)
         );
  AOI22_X1 U4597 ( .A1(n3469), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3573) );
  AOI22_X1 U4598 ( .A1(n3356), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3572) );
  AOI22_X1 U4599 ( .A1(n4310), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3571) );
  AOI22_X1 U4600 ( .A1(n3569), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4288), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3570) );
  NAND4_X1 U4601 ( .A1(n3573), .A2(n3572), .A3(n3571), .A4(n3570), .ZN(n3574)
         );
  NOR2_X1 U4602 ( .A1(n3575), .A2(n3574), .ZN(n3578) );
  NAND2_X1 U4603 ( .A1(n3418), .A2(EAX_REG_9__SCAN_IN), .ZN(n3577) );
  NAND2_X1 U4604 ( .A1(n4384), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3576)
         );
  OAI211_X1 U4605 ( .C1(n3627), .C2(n3578), .A(n3577), .B(n3576), .ZN(n3579)
         );
  AOI21_X1 U4606 ( .B1(n3580), .B2(n5183), .A(n3579), .ZN(n5052) );
  AOI22_X1 U4607 ( .A1(n4308), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4608 ( .A1(n4316), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4609 ( .A1(n3499), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4610 ( .A1(n4288), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3582) );
  NAND4_X1 U4611 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(n3591)
         );
  AOI22_X1 U4612 ( .A1(n4307), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3589) );
  AOI22_X1 U4613 ( .A1(n4310), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3588) );
  AOI22_X1 U4614 ( .A1(n3356), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4615 ( .A1(n4311), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3586) );
  NAND4_X1 U4616 ( .A1(n3589), .A2(n3588), .A3(n3587), .A4(n3586), .ZN(n3590)
         );
  OAI21_X1 U4617 ( .B1(n3591), .B2(n3590), .A(n3678), .ZN(n3595) );
  XNOR2_X1 U4618 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3597), .ZN(n5567)
         );
  AOI22_X1 U4619 ( .A1(n5183), .A2(n5567), .B1(n4384), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3594) );
  NAND2_X1 U4620 ( .A1(n3418), .A2(EAX_REG_10__SCAN_IN), .ZN(n3593) );
  AOI21_X1 U4621 ( .B1(n6673), .B2(n3598), .A(n3629), .ZN(n6149) );
  OR2_X1 U4622 ( .A1(n6149), .A2(n3492), .ZN(n3614) );
  AOI22_X1 U4623 ( .A1(n4309), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4624 ( .A1(n4311), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4625 ( .A1(n4317), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4626 ( .A1(n3499), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3599) );
  NAND4_X1 U4627 ( .A1(n3602), .A2(n3601), .A3(n3600), .A4(n3599), .ZN(n3608)
         );
  AOI22_X1 U4628 ( .A1(n4308), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3606) );
  AOI22_X1 U4629 ( .A1(n4310), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3605) );
  AOI22_X1 U4630 ( .A1(n3356), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3604) );
  AOI22_X1 U4631 ( .A1(n4288), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3603) );
  NAND4_X1 U4632 ( .A1(n3606), .A2(n3605), .A3(n3604), .A4(n3603), .ZN(n3607)
         );
  NOR2_X1 U4633 ( .A1(n3608), .A2(n3607), .ZN(n3611) );
  NAND2_X1 U4634 ( .A1(n3418), .A2(EAX_REG_11__SCAN_IN), .ZN(n3610) );
  NAND2_X1 U4635 ( .A1(n4384), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3609)
         );
  OAI211_X1 U4636 ( .C1(n3627), .C2(n3611), .A(n3610), .B(n3609), .ZN(n3612)
         );
  INV_X1 U4637 ( .A(n3612), .ZN(n3613) );
  AOI22_X1 U4638 ( .A1(n3469), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4639 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4311), .B1(n4309), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4640 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3362), .B1(n4317), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4641 ( .A1(n3569), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3615) );
  NAND4_X1 U4642 ( .A1(n3618), .A2(n3617), .A3(n3616), .A4(n3615), .ZN(n3624)
         );
  AOI22_X1 U4643 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4308), .B1(n4307), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4644 ( .A1(n3356), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4645 ( .A1(n4310), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4646 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3499), .B1(n4288), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3619) );
  NAND4_X1 U4647 ( .A1(n3622), .A2(n3621), .A3(n3620), .A4(n3619), .ZN(n3623)
         );
  NOR2_X1 U4648 ( .A1(n3624), .A2(n3623), .ZN(n3628) );
  XNOR2_X1 U4649 ( .A(n3629), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6777)
         );
  NAND2_X1 U4650 ( .A1(n6777), .A2(n5183), .ZN(n3626) );
  AOI22_X1 U4651 ( .A1(n3418), .A2(EAX_REG_12__SCAN_IN), .B1(n4384), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3625) );
  OAI211_X1 U4652 ( .C1(n3628), .C2(n3627), .A(n3626), .B(n3625), .ZN(n5367)
         );
  INV_X1 U4653 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3632) );
  OAI21_X1 U4654 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3630), .A(n3653), 
        .ZN(n5984) );
  NAND2_X1 U4655 ( .A1(n5984), .A2(n5183), .ZN(n3631) );
  OAI21_X1 U4656 ( .B1(n3632), .B2(n4021), .A(n3631), .ZN(n3633) );
  AOI21_X1 U4657 ( .B1(n4357), .B2(EAX_REG_13__SCAN_IN), .A(n3633), .ZN(n3636)
         );
  NAND2_X2 U4658 ( .A1(n3635), .A2(n3634), .ZN(n3650) );
  NAND2_X1 U4659 ( .A1(n3637), .A2(n3636), .ZN(n3638) );
  AOI22_X1 U4660 ( .A1(n3469), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4661 ( .A1(n4310), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4662 ( .A1(n3356), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4663 ( .A1(n4316), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3639) );
  NAND4_X1 U4664 ( .A1(n3642), .A2(n3641), .A3(n3640), .A4(n3639), .ZN(n3648)
         );
  AOI22_X1 U4665 ( .A1(n4308), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4666 ( .A1(n4311), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4667 ( .A1(n4317), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4668 ( .A1(n3499), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4288), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3643) );
  NAND4_X1 U4669 ( .A1(n3646), .A2(n3645), .A3(n3644), .A4(n3643), .ZN(n3647)
         );
  OR2_X1 U4670 ( .A1(n3648), .A2(n3647), .ZN(n3649) );
  AND2_X1 U4671 ( .A1(n3678), .A2(n3649), .ZN(n5415) );
  INV_X1 U4672 ( .A(EAX_REG_14__SCAN_IN), .ZN(n3652) );
  OAI21_X1 U4673 ( .B1(PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n6604), .A(n5874), 
        .ZN(n3651) );
  OAI21_X1 U4674 ( .B1(n4023), .B2(n3652), .A(n3651), .ZN(n3657) );
  NOR2_X1 U4675 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n3654), .ZN(n3655)
         );
  NOR2_X1 U4676 ( .A1(n3681), .A2(n3655), .ZN(n5970) );
  NAND2_X1 U4677 ( .A1(n5970), .A2(n5183), .ZN(n3656) );
  NAND2_X1 U4678 ( .A1(n3657), .A2(n3656), .ZN(n3669) );
  AOI22_X1 U4679 ( .A1(n4308), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U4680 ( .A1(n3356), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4681 ( .A1(n3362), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3659) );
  AOI22_X1 U4682 ( .A1(n4288), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3658) );
  NAND4_X1 U4683 ( .A1(n3661), .A2(n3660), .A3(n3659), .A4(n3658), .ZN(n3667)
         );
  AOI22_X1 U4684 ( .A1(n3469), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4685 ( .A1(n4310), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4686 ( .A1(n4311), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4687 ( .A1(n3475), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3662) );
  NAND4_X1 U4688 ( .A1(n3665), .A2(n3664), .A3(n3663), .A4(n3662), .ZN(n3666)
         );
  OAI21_X1 U4689 ( .B1(n3667), .B2(n3666), .A(n3678), .ZN(n3668) );
  NAND2_X1 U4690 ( .A1(n3669), .A2(n3668), .ZN(n5356) );
  AOI22_X1 U4691 ( .A1(n3469), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3673) );
  AOI22_X1 U4692 ( .A1(n4311), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4693 ( .A1(n3356), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4694 ( .A1(n4288), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3670) );
  NAND4_X1 U4695 ( .A1(n3673), .A2(n3672), .A3(n3671), .A4(n3670), .ZN(n3680)
         );
  AOI22_X1 U4696 ( .A1(n4308), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4310), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3677) );
  AOI22_X1 U4697 ( .A1(n4309), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4698 ( .A1(n3499), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3675) );
  AOI22_X1 U4699 ( .A1(n4316), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3674) );
  NAND4_X1 U4700 ( .A1(n3677), .A2(n3676), .A3(n3675), .A4(n3674), .ZN(n3679)
         );
  OAI21_X1 U4701 ( .B1(n3680), .B2(n3679), .A(n3678), .ZN(n3684) );
  OAI21_X1 U4702 ( .B1(n3681), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n3717), 
        .ZN(n5542) );
  AOI22_X1 U4703 ( .A1(n5542), .A2(n5183), .B1(PHYADDRPOINTER_REG_15__SCAN_IN), 
        .B2(n4384), .ZN(n3683) );
  NAND2_X1 U4704 ( .A1(n3418), .A2(EAX_REG_15__SCAN_IN), .ZN(n3682) );
  NAND2_X1 U4705 ( .A1(n3273), .A2(n4566), .ZN(n3686) );
  AOI22_X1 U4706 ( .A1(n4310), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4707 ( .A1(n4311), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4708 ( .A1(n3356), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4709 ( .A1(n3475), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3687) );
  NAND4_X1 U4710 ( .A1(n3690), .A2(n3689), .A3(n3688), .A4(n3687), .ZN(n3696)
         );
  AOI22_X1 U4711 ( .A1(n4308), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4712 ( .A1(n3454), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3693) );
  AOI22_X1 U4713 ( .A1(n4316), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4714 ( .A1(n3569), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4288), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3691) );
  NAND4_X1 U4715 ( .A1(n3694), .A2(n3693), .A3(n3692), .A4(n3691), .ZN(n3695)
         );
  OR2_X1 U4716 ( .A1(n3696), .A2(n3695), .ZN(n3697) );
  NAND2_X1 U4717 ( .A1(n4354), .A2(n3697), .ZN(n3700) );
  XNOR2_X1 U4718 ( .A(n3717), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5955)
         );
  INV_X1 U4719 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3716) );
  OAI22_X1 U4720 ( .A1(n5955), .A2(n3492), .B1(n3716), .B2(n4021), .ZN(n3698)
         );
  AOI21_X1 U4721 ( .B1(n4357), .B2(EAX_REG_16__SCAN_IN), .A(n3698), .ZN(n3699)
         );
  NAND2_X1 U4722 ( .A1(n3700), .A2(n3699), .ZN(n5347) );
  AOI22_X1 U4723 ( .A1(n4308), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4724 ( .A1(n4310), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4725 ( .A1(n3499), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4726 ( .A1(n4288), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3701) );
  NAND4_X1 U4727 ( .A1(n3704), .A2(n3703), .A3(n3702), .A4(n3701), .ZN(n3710)
         );
  AOI22_X1 U4728 ( .A1(n4307), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3708) );
  AOI22_X1 U4729 ( .A1(n4311), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3707) );
  AOI22_X1 U4730 ( .A1(n3356), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4731 ( .A1(n4317), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3705) );
  NAND4_X1 U4732 ( .A1(n3708), .A2(n3707), .A3(n3706), .A4(n3705), .ZN(n3709)
         );
  NOR2_X1 U4733 ( .A1(n3710), .A2(n3709), .ZN(n3713) );
  INV_X1 U4734 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6743) );
  AOI21_X1 U4735 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n6743), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3711) );
  AOI21_X1 U4736 ( .B1(n4357), .B2(EAX_REG_17__SCAN_IN), .A(n3711), .ZN(n3712)
         );
  OAI21_X1 U4737 ( .B1(n4349), .B2(n3713), .A(n3712), .ZN(n3720) );
  OAI21_X1 U4738 ( .B1(n3717), .B2(n3716), .A(n6743), .ZN(n3718) );
  AND2_X1 U4739 ( .A1(n3722), .A2(n3718), .ZN(n5527) );
  NAND2_X1 U4740 ( .A1(n5527), .A2(n5183), .ZN(n3719) );
  INV_X1 U4741 ( .A(n5246), .ZN(n3721) );
  NOR2_X2 U4742 ( .A1(n3940), .A2(n3721), .ZN(n5240) );
  NAND2_X1 U4743 ( .A1(n3722), .A2(n3023), .ZN(n3723) );
  NAND2_X1 U4744 ( .A1(n3750), .A2(n3723), .ZN(n5520) );
  AOI22_X1 U4745 ( .A1(n4308), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4746 ( .A1(n4310), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4747 ( .A1(n4309), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4748 ( .A1(n3356), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3724) );
  NAND4_X1 U4749 ( .A1(n3727), .A2(n3726), .A3(n3725), .A4(n3724), .ZN(n3733)
         );
  AOI22_X1 U4750 ( .A1(n4311), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4751 ( .A1(n4316), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3730) );
  AOI22_X1 U4752 ( .A1(n3475), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3729) );
  AOI22_X1 U4753 ( .A1(n4288), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3728) );
  NAND4_X1 U4754 ( .A1(n3731), .A2(n3730), .A3(n3729), .A4(n3728), .ZN(n3732)
         );
  OR2_X1 U4755 ( .A1(n3733), .A2(n3732), .ZN(n3734) );
  NAND2_X1 U4756 ( .A1(n4354), .A2(n3734), .ZN(n3736) );
  AOI22_X1 U4757 ( .A1(n3418), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6409), .ZN(n3735) );
  NAND2_X1 U4758 ( .A1(n3736), .A2(n3735), .ZN(n3955) );
  MUX2_X1 U4759 ( .A(n5520), .B(n3955), .S(n3492), .Z(n5239) );
  NAND2_X1 U4760 ( .A1(n5240), .A2(n5239), .ZN(n3754) );
  AOI22_X1 U4761 ( .A1(n4308), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4762 ( .A1(n3469), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4763 ( .A1(n4310), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4764 ( .A1(n4311), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3737) );
  NAND4_X1 U4765 ( .A1(n3740), .A2(n3739), .A3(n3738), .A4(n3737), .ZN(n3746)
         );
  AOI22_X1 U4766 ( .A1(n4317), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4767 ( .A1(n3356), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4768 ( .A1(n3499), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4769 ( .A1(n4288), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3741) );
  NAND4_X1 U4770 ( .A1(n3744), .A2(n3743), .A3(n3742), .A4(n3741), .ZN(n3745)
         );
  NOR2_X1 U4771 ( .A1(n3746), .A2(n3745), .ZN(n3749) );
  AOI21_X1 U4772 ( .B1(n6755), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3747) );
  AOI21_X1 U4773 ( .B1(n4357), .B2(EAX_REG_19__SCAN_IN), .A(n3747), .ZN(n3748)
         );
  OAI21_X1 U4774 ( .B1(n4349), .B2(n3749), .A(n3748), .ZN(n3753) );
  NAND2_X1 U4775 ( .A1(n3750), .A2(n6755), .ZN(n3751) );
  NAND2_X1 U4776 ( .A1(n3914), .A2(n3751), .ZN(n5231) );
  NOR2_X2 U4777 ( .A1(n3754), .A2(n3755), .ZN(n3929) );
  INV_X1 U4778 ( .A(n3929), .ZN(n3757) );
  INV_X1 U4779 ( .A(n5407), .ZN(n3758) );
  NAND2_X1 U4780 ( .A1(n4397), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6516) );
  NAND2_X1 U4781 ( .A1(n3785), .A2(n3784), .ZN(n3773) );
  NAND2_X1 U4782 ( .A1(n3773), .A2(n3772), .ZN(n3766) );
  NAND2_X1 U4783 ( .A1(n3766), .A2(n3764), .ZN(n3816) );
  XNOR2_X1 U4784 ( .A(n3816), .B(n3814), .ZN(n3760) );
  INV_X1 U4785 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3762) );
  NAND2_X1 U4786 ( .A1(n3799), .A2(n3762), .ZN(n3798) );
  NAND2_X1 U4787 ( .A1(n3763), .A2(n3870), .ZN(n3769) );
  INV_X1 U4788 ( .A(n3764), .ZN(n3765) );
  XNOR2_X1 U4789 ( .A(n3766), .B(n3765), .ZN(n3767) );
  NAND2_X1 U4790 ( .A1(n3767), .A2(n6605), .ZN(n3768) );
  INV_X1 U4791 ( .A(n5085), .ZN(n3770) );
  NAND2_X1 U4792 ( .A1(n3770), .A2(n6256), .ZN(n3771) );
  AND2_X1 U4793 ( .A1(n3798), .A2(n3771), .ZN(n3797) );
  INV_X1 U4794 ( .A(n3870), .ZN(n3780) );
  XNOR2_X1 U4795 ( .A(n3773), .B(n3772), .ZN(n3775) );
  AOI21_X1 U4796 ( .B1(n3775), .B2(n6605), .A(n3774), .ZN(n3776) );
  NAND2_X1 U4797 ( .A1(n6174), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3793)
         );
  INV_X1 U4798 ( .A(n6605), .ZN(n4072) );
  INV_X1 U4799 ( .A(n3774), .ZN(n3777) );
  OAI21_X1 U4800 ( .B1(n4072), .B2(n3784), .A(n3777), .ZN(n3778) );
  INV_X1 U4801 ( .A(n3778), .ZN(n3779) );
  NAND2_X1 U4802 ( .A1(n4487), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3781)
         );
  INV_X1 U4803 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U4804 ( .A1(n3781), .A2(n6269), .ZN(n3783) );
  AND2_X1 U4805 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3782) );
  NAND2_X1 U4806 ( .A1(n4487), .A2(n3782), .ZN(n3791) );
  AND2_X1 U4807 ( .A1(n3783), .A2(n3791), .ZN(n4546) );
  NAND2_X1 U4808 ( .A1(n2964), .A2(n3870), .ZN(n3790) );
  XNOR2_X1 U4809 ( .A(n3785), .B(n3784), .ZN(n3787) );
  OAI211_X1 U4810 ( .C1(n3787), .C2(n4072), .A(n3786), .B(n5372), .ZN(n3788)
         );
  INV_X1 U4811 ( .A(n3788), .ZN(n3789) );
  NAND2_X1 U4812 ( .A1(n3790), .A2(n3789), .ZN(n4547) );
  INV_X1 U4813 ( .A(n3791), .ZN(n3792) );
  NAND2_X1 U4814 ( .A1(n3793), .A2(n6175), .ZN(n3796) );
  INV_X1 U4815 ( .A(n6174), .ZN(n3794) );
  INV_X1 U4816 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U4817 ( .A1(n3794), .A2(n6173), .ZN(n3795) );
  NAND2_X1 U4818 ( .A1(n3797), .A2(n5086), .ZN(n3803) );
  NAND2_X1 U4819 ( .A1(n3798), .A2(n6164), .ZN(n3801) );
  AND2_X1 U4820 ( .A1(n3801), .A2(n3800), .ZN(n3802) );
  NAND2_X1 U4821 ( .A1(n3803), .A2(n3802), .ZN(n4727) );
  NAND2_X1 U4822 ( .A1(n3804), .A2(n3870), .ZN(n3809) );
  INV_X1 U4823 ( .A(n3814), .ZN(n3805) );
  OR2_X1 U4824 ( .A1(n3816), .A2(n3805), .ZN(n3806) );
  XNOR2_X1 U4825 ( .A(n3806), .B(n3813), .ZN(n3807) );
  NAND2_X1 U4826 ( .A1(n3807), .A2(n6605), .ZN(n3808) );
  INV_X1 U4827 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4734) );
  NAND2_X1 U4828 ( .A1(n4727), .A2(n4729), .ZN(n4728) );
  NAND2_X1 U4829 ( .A1(n3810), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3811)
         );
  NAND2_X1 U4830 ( .A1(n4728), .A2(n3811), .ZN(n6154) );
  NAND2_X1 U4831 ( .A1(n3814), .A2(n3813), .ZN(n3815) );
  OR2_X1 U4832 ( .A1(n3816), .A2(n3815), .ZN(n3823) );
  XNOR2_X1 U4833 ( .A(n3823), .B(n3824), .ZN(n3817) );
  NAND2_X1 U4834 ( .A1(n3817), .A2(n6605), .ZN(n3818) );
  INV_X1 U4835 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6236) );
  XNOR2_X1 U4836 ( .A(n3820), .B(n6236), .ZN(n6156) );
  NAND2_X1 U4837 ( .A1(n3820), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3821)
         );
  NAND2_X1 U4838 ( .A1(n3822), .A2(n3870), .ZN(n3828) );
  INV_X1 U4839 ( .A(n3823), .ZN(n3825) );
  NAND2_X1 U4840 ( .A1(n3825), .A2(n3824), .ZN(n3836) );
  XNOR2_X1 U4841 ( .A(n3836), .B(n3837), .ZN(n3826) );
  NAND2_X1 U4842 ( .A1(n3826), .A2(n6605), .ZN(n3827) );
  NAND2_X1 U4843 ( .A1(n3828), .A2(n3827), .ZN(n3830) );
  INV_X1 U4844 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3829) );
  XNOR2_X1 U4845 ( .A(n3830), .B(n3829), .ZN(n5045) );
  NAND2_X1 U4846 ( .A1(n3830), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3831)
         );
  NAND2_X1 U4847 ( .A1(n3870), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3833) );
  INV_X1 U4848 ( .A(n3836), .ZN(n3838) );
  NAND3_X1 U4849 ( .A1(n3838), .A2(n6605), .A3(n3837), .ZN(n3839) );
  NAND2_X1 U4850 ( .A1(n3848), .A2(n3839), .ZN(n3840) );
  INV_X1 U4851 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4125) );
  XNOR2_X1 U4852 ( .A(n3840), .B(n4125), .ZN(n5582) );
  NAND2_X1 U4853 ( .A1(n3840), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3841)
         );
  INV_X1 U4854 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6735) );
  NAND2_X1 U4855 ( .A1(n5533), .A2(n6735), .ZN(n5573) );
  NOR3_X1 U4856 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .A3(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .ZN(n3842) );
  INV_X4 U4857 ( .A(n3844), .ZN(n6146) );
  NAND2_X1 U4858 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3845) );
  INV_X1 U4859 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U4860 ( .A1(n6146), .A2(n5751), .ZN(n5552) );
  INV_X1 U4861 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5924) );
  INV_X1 U4862 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U4863 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4244) );
  NAND2_X1 U4864 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4255) );
  OAI21_X1 U4865 ( .B1(n4244), .B2(n4255), .A(n5533), .ZN(n3847) );
  INV_X1 U4866 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3849) );
  INV_X1 U4867 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5707) );
  INV_X1 U4868 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5721) );
  INV_X1 U4869 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5731) );
  NAND4_X1 U4870 ( .A1(n3849), .A2(n5707), .A3(n5721), .A4(n5731), .ZN(n3850)
         );
  NAND2_X1 U4871 ( .A1(n3933), .A2(n3850), .ZN(n3851) );
  XNOR2_X1 U4872 ( .A(n6146), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3852)
         );
  XNOR2_X1 U4873 ( .A(n4182), .B(n3852), .ZN(n5693) );
  INV_X1 U4874 ( .A(n5693), .ZN(n3911) );
  NAND2_X1 U4875 ( .A1(n4656), .A2(n5372), .ZN(n3853) );
  NAND2_X1 U4876 ( .A1(n5297), .A2(n3853), .ZN(n3866) );
  INV_X1 U4877 ( .A(n3866), .ZN(n3875) );
  XNOR2_X1 U4878 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3859) );
  NAND2_X1 U4879 ( .A1(n3863), .A2(n3859), .ZN(n3855) );
  NAND2_X1 U4880 ( .A1(n4936), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3854) );
  NAND2_X1 U4881 ( .A1(n3855), .A2(n3854), .ZN(n3878) );
  XNOR2_X1 U4882 ( .A(n3857), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3876)
         );
  XNOR2_X1 U4883 ( .A(n3878), .B(n3876), .ZN(n4199) );
  NAND2_X1 U4884 ( .A1(n3893), .A2(n4199), .ZN(n3874) );
  NAND2_X1 U4885 ( .A1(n3893), .A2(n4237), .ZN(n3858) );
  INV_X1 U4886 ( .A(n3859), .ZN(n3860) );
  XNOR2_X1 U4887 ( .A(n3860), .B(n3863), .ZN(n4200) );
  AND2_X1 U4888 ( .A1(n3861), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3862)
         );
  NOR2_X1 U4889 ( .A1(n3863), .A2(n3862), .ZN(n3868) );
  AOI21_X1 U4890 ( .B1(n3865), .B2(n3868), .A(n3864), .ZN(n3867) );
  NAND2_X1 U4891 ( .A1(n3893), .A2(n3868), .ZN(n3869) );
  OAI211_X1 U4892 ( .C1(n4199), .C2(n3888), .A(n3874), .B(n3875), .ZN(n3872)
         );
  OAI21_X1 U4893 ( .B1(n3875), .B2(n3874), .A(n3873), .ZN(n3898) );
  INV_X1 U4894 ( .A(n3876), .ZN(n3877) );
  NAND2_X1 U4895 ( .A1(n3878), .A2(n3877), .ZN(n3880) );
  NAND2_X1 U4896 ( .A1(n6474), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3879) );
  NAND2_X1 U4897 ( .A1(n3880), .A2(n3879), .ZN(n3886) );
  XNOR2_X1 U4898 ( .A(n4613), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3885)
         );
  INV_X1 U4899 ( .A(n3885), .ZN(n3881) );
  NAND2_X1 U4900 ( .A1(n3886), .A2(n3881), .ZN(n3883) );
  NAND2_X1 U4901 ( .A1(n6397), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3882) );
  NAND2_X1 U4902 ( .A1(n3883), .A2(n3882), .ZN(n3890) );
  NAND2_X1 U4903 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3884), .ZN(n3891) );
  OR2_X1 U4904 ( .A1(n3890), .A2(n3891), .ZN(n4203) );
  XNOR2_X1 U4905 ( .A(n3886), .B(n3885), .ZN(n4198) );
  INV_X1 U4906 ( .A(n3895), .ZN(n3887) );
  NAND2_X1 U4907 ( .A1(n3888), .A2(n3887), .ZN(n3897) );
  AOI22_X1 U4908 ( .A1(n3893), .A2(n3899), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6509), .ZN(n3894) );
  OAI21_X1 U4909 ( .B1(n3900), .B2(n3895), .A(n3894), .ZN(n3896) );
  AOI21_X1 U4910 ( .B1(n4088), .B2(n4681), .A(n4078), .ZN(n3903) );
  NAND2_X1 U4911 ( .A1(n4219), .A2(n3270), .ZN(n6481) );
  NAND2_X1 U4912 ( .A1(n6406), .A2(n3904), .ZN(n6600) );
  NAND2_X1 U4913 ( .A1(n6600), .A2(n6509), .ZN(n3905) );
  NAND2_X1 U4914 ( .A1(n6509), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3907) );
  NAND2_X1 U4915 ( .A1(n6604), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3906) );
  AND2_X1 U4916 ( .A1(n3907), .A2(n3906), .ZN(n4522) );
  INV_X2 U4917 ( .A(n5576), .ZN(n5565) );
  AND2_X1 U4918 ( .A1(n6233), .A2(REIP_REG_19__SCAN_IN), .ZN(n5686) );
  AOI21_X1 U4919 ( .B1(n5565), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5686), 
        .ZN(n3908) );
  OAI21_X1 U4920 ( .B1(n6182), .B2(n5231), .A(n3908), .ZN(n3909) );
  NAND2_X1 U4921 ( .A1(n3914), .A2(n5210), .ZN(n3915) );
  NAND2_X1 U4922 ( .A1(n3976), .A2(n3915), .ZN(n5209) );
  AOI22_X1 U4923 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4308), .B1(n3469), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4924 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4311), .B1(n4310), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4925 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3362), .B1(n4316), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4926 ( .A1(n4288), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3916) );
  NAND4_X1 U4927 ( .A1(n3919), .A2(n3918), .A3(n3917), .A4(n3916), .ZN(n3925)
         );
  AOI22_X1 U4928 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3454), .B1(n4307), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4929 ( .A1(n3356), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4930 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4309), .B1(n4318), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4931 ( .A1(n3475), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3920) );
  NAND4_X1 U4932 ( .A1(n3923), .A2(n3922), .A3(n3921), .A4(n3920), .ZN(n3924)
         );
  OR2_X1 U4933 ( .A1(n3925), .A2(n3924), .ZN(n3926) );
  NAND2_X1 U4934 ( .A1(n4354), .A2(n3926), .ZN(n3928) );
  AOI22_X1 U4935 ( .A1(n3418), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6409), .ZN(n3927) );
  NAND2_X1 U4936 ( .A1(n3928), .A2(n3927), .ZN(n3954) );
  MUX2_X1 U4937 ( .A(n5209), .B(n3954), .S(n3492), .Z(n3930) );
  INV_X1 U4938 ( .A(n5208), .ZN(n3931) );
  INV_X1 U4939 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3932) );
  XNOR2_X1 U4940 ( .A(n5533), .B(n3932), .ZN(n4374) );
  XOR2_X1 U4941 ( .A(n4374), .B(n4375), .Z(n5684) );
  AND2_X1 U4942 ( .A1(n6233), .A2(REIP_REG_20__SCAN_IN), .ZN(n5676) );
  AOI21_X1 U4943 ( .B1(n5565), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5676), 
        .ZN(n3934) );
  OAI21_X1 U4944 ( .B1(n6182), .B2(n5209), .A(n3934), .ZN(n3935) );
  INV_X1 U4945 ( .A(n3935), .ZN(n3936) );
  AOI22_X1 U4946 ( .A1(n4308), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4947 ( .A1(n4310), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4948 ( .A1(n4316), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4949 ( .A1(n4288), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3941) );
  NAND4_X1 U4950 ( .A1(n3944), .A2(n3943), .A3(n3942), .A4(n3941), .ZN(n3950)
         );
  AOI22_X1 U4951 ( .A1(n3469), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4952 ( .A1(n3356), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4953 ( .A1(n4311), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4954 ( .A1(n3475), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3945) );
  NAND4_X1 U4955 ( .A1(n3948), .A2(n3947), .A3(n3946), .A4(n3945), .ZN(n3949)
         );
  OR2_X1 U4956 ( .A1(n3950), .A2(n3949), .ZN(n3951) );
  NAND2_X1 U4957 ( .A1(n4354), .A2(n3951), .ZN(n3953) );
  AOI22_X1 U4958 ( .A1(n3418), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6409), .ZN(n3952) );
  NAND2_X1 U4959 ( .A1(n3953), .A2(n3952), .ZN(n5184) );
  AND4_X1 U4960 ( .A1(n3955), .A2(n3954), .A3(n5184), .A4(n3492), .ZN(n3961)
         );
  INV_X1 U4961 ( .A(n3956), .ZN(n3957) );
  NAND2_X1 U4962 ( .A1(n3957), .A2(n3019), .ZN(n3958) );
  NAND2_X1 U4963 ( .A1(n4019), .A2(n3958), .ZN(n5502) );
  OAI211_X1 U4964 ( .C1(n3961), .C2(n3960), .A(n5246), .B(n3959), .ZN(n3979)
         );
  AOI22_X1 U4965 ( .A1(n4308), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4966 ( .A1(n3469), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4967 ( .A1(n4282), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4968 ( .A1(n4311), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3962) );
  NAND4_X1 U4969 ( .A1(n3965), .A2(n3964), .A3(n3963), .A4(n3962), .ZN(n3971)
         );
  AOI22_X1 U4970 ( .A1(n4317), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U4971 ( .A1(n3356), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4972 ( .A1(n3499), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4973 ( .A1(n4288), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3966) );
  NAND4_X1 U4974 ( .A1(n3969), .A2(n3968), .A3(n3967), .A4(n3966), .ZN(n3970)
         );
  NOR2_X1 U4975 ( .A1(n3971), .A2(n3970), .ZN(n3975) );
  AOI21_X1 U4976 ( .B1(n3972), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3973) );
  AOI21_X1 U4977 ( .B1(n4357), .B2(EAX_REG_21__SCAN_IN), .A(n3973), .ZN(n3974)
         );
  OAI21_X1 U4978 ( .B1(n4349), .B2(n3975), .A(n3974), .ZN(n3978) );
  XNOR2_X1 U4979 ( .A(n3976), .B(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5510)
         );
  NAND2_X1 U4980 ( .A1(n5510), .A2(n5183), .ZN(n3977) );
  NAND2_X1 U4981 ( .A1(n3978), .A2(n3977), .ZN(n5187) );
  AOI22_X1 U4982 ( .A1(n4309), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4983 ( .A1(n4311), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4984 ( .A1(n3356), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4985 ( .A1(n3569), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3981) );
  NAND4_X1 U4986 ( .A1(n3984), .A2(n3983), .A3(n3982), .A4(n3981), .ZN(n3990)
         );
  AOI22_X1 U4987 ( .A1(n4308), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U4988 ( .A1(n4310), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U4989 ( .A1(n4317), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U4990 ( .A1(n3499), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4288), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3985) );
  NAND4_X1 U4991 ( .A1(n3988), .A2(n3987), .A3(n3986), .A4(n3985), .ZN(n3989)
         );
  NOR2_X1 U4992 ( .A1(n3990), .A2(n3989), .ZN(n4006) );
  AOI22_X1 U4993 ( .A1(n4308), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4994 ( .A1(n3469), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U4995 ( .A1(n4310), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4996 ( .A1(n4311), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3991) );
  NAND4_X1 U4997 ( .A1(n3994), .A2(n3993), .A3(n3992), .A4(n3991), .ZN(n4000)
         );
  AOI22_X1 U4998 ( .A1(n4317), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4999 ( .A1(n3356), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U5000 ( .A1(n3499), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U5001 ( .A1(n4288), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3995) );
  NAND4_X1 U5002 ( .A1(n3998), .A2(n3997), .A3(n3996), .A4(n3995), .ZN(n3999)
         );
  NOR2_X1 U5003 ( .A1(n4000), .A2(n3999), .ZN(n4007) );
  XOR2_X1 U5004 ( .A(n4006), .B(n4007), .Z(n4003) );
  INV_X1 U5005 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4001) );
  INV_X1 U5006 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5173) );
  OAI22_X1 U5007 ( .A1(n4023), .A2(n4001), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5173), .ZN(n4002) );
  AOI21_X1 U5008 ( .B1(n4354), .B2(n4003), .A(n4002), .ZN(n4063) );
  NAND2_X1 U5009 ( .A1(n4063), .A2(n3492), .ZN(n4005) );
  XNOR2_X1 U5010 ( .A(n4019), .B(n5173), .ZN(n5494) );
  OR2_X1 U5011 ( .A1(n5494), .A2(n3492), .ZN(n4004) );
  NAND2_X1 U5012 ( .A1(n4005), .A2(n4004), .ZN(n5172) );
  OR2_X1 U5013 ( .A1(n4007), .A2(n4006), .ZN(n4028) );
  AOI22_X1 U5014 ( .A1(n3499), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U5015 ( .A1(n4310), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U5016 ( .A1(n4311), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U5017 ( .A1(n3569), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4008) );
  NAND4_X1 U5018 ( .A1(n4011), .A2(n4010), .A3(n4009), .A4(n4008), .ZN(n4017)
         );
  AOI22_X1 U5019 ( .A1(n3356), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U5020 ( .A1(n4308), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4014) );
  INV_X1 U5021 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n6640) );
  AOI22_X1 U5022 ( .A1(n4317), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U5023 ( .A1(n4307), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4288), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4012) );
  NAND4_X1 U5024 ( .A1(n4015), .A2(n4014), .A3(n4013), .A4(n4012), .ZN(n4016)
         );
  NOR2_X1 U5025 ( .A1(n4017), .A2(n4016), .ZN(n4027) );
  XNOR2_X1 U5026 ( .A(n4028), .B(n4027), .ZN(n4026) );
  INV_X1 U5027 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6638) );
  OAI21_X1 U5028 ( .B1(n4019), .B2(n5173), .A(n6638), .ZN(n4020) );
  NAND2_X1 U5029 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4018) );
  NAND2_X1 U5030 ( .A1(n4020), .A2(n4045), .ZN(n5482) );
  INV_X1 U5031 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4022) );
  OAI22_X1 U5032 ( .A1(n4023), .A2(n4022), .B1(n6638), .B2(n4021), .ZN(n4024)
         );
  AOI21_X1 U5033 ( .B1(n5482), .B2(n5183), .A(n4024), .ZN(n4025) );
  OAI21_X1 U5034 ( .B1(n4026), .B2(n4349), .A(n4025), .ZN(n4062) );
  OR2_X1 U5035 ( .A1(n4028), .A2(n4027), .ZN(n4047) );
  AOI22_X1 U5036 ( .A1(n3469), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U5037 ( .A1(n4309), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U5038 ( .A1(n4317), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U5039 ( .A1(n3569), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4029) );
  NAND4_X1 U5040 ( .A1(n4032), .A2(n4031), .A3(n4030), .A4(n4029), .ZN(n4038)
         );
  AOI22_X1 U5041 ( .A1(n4308), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U5042 ( .A1(n4311), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4310), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U5043 ( .A1(n3356), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U5044 ( .A1(n3499), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4288), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4033) );
  NAND4_X1 U5045 ( .A1(n4036), .A2(n4035), .A3(n4034), .A4(n4033), .ZN(n4037)
         );
  NOR2_X1 U5046 ( .A1(n4038), .A2(n4037), .ZN(n4048) );
  XOR2_X1 U5047 ( .A(n4047), .B(n4048), .Z(n4039) );
  NAND2_X1 U5048 ( .A1(n4039), .A2(n4354), .ZN(n4042) );
  INV_X1 U5049 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5154) );
  AOI21_X1 U5050 ( .B1(n5154), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4040) );
  AOI21_X1 U5051 ( .B1(n4357), .B2(EAX_REG_25__SCAN_IN), .A(n4040), .ZN(n4041)
         );
  NAND2_X1 U5052 ( .A1(n4042), .A2(n4041), .ZN(n4044) );
  XNOR2_X1 U5053 ( .A(n4045), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5153)
         );
  NAND2_X1 U5054 ( .A1(n5153), .A2(n5183), .ZN(n4043) );
  NAND2_X1 U5055 ( .A1(n3021), .A2(n3020), .ZN(n4046) );
  NAND2_X1 U5056 ( .A1(n4337), .A2(n4046), .ZN(n5467) );
  AND2_X1 U5057 ( .A1(n5467), .A2(n5183), .ZN(n4061) );
  NOR2_X1 U5058 ( .A1(n4048), .A2(n4047), .ZN(n4306) );
  AOI22_X1 U5059 ( .A1(n4308), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U5060 ( .A1(n3469), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U5061 ( .A1(n4282), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4050) );
  AOI22_X1 U5062 ( .A1(n4311), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4049) );
  NAND4_X1 U5063 ( .A1(n4052), .A2(n4051), .A3(n4050), .A4(n4049), .ZN(n4058)
         );
  AOI22_X1 U5064 ( .A1(n4317), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U5065 ( .A1(n3356), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U5066 ( .A1(n3499), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U5067 ( .A1(n4288), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4053) );
  NAND4_X1 U5068 ( .A1(n4056), .A2(n4055), .A3(n4054), .A4(n4053), .ZN(n4057)
         );
  XNOR2_X1 U5069 ( .A(n4306), .B(n4305), .ZN(n4060) );
  AOI22_X1 U5070 ( .A1(n3418), .A2(EAX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6409), .ZN(n4059) );
  OAI21_X1 U5071 ( .B1(n4060), .B2(n4349), .A(n4059), .ZN(n4064) );
  INV_X1 U5072 ( .A(n4062), .ZN(n5164) );
  INV_X1 U5073 ( .A(n4063), .ZN(n4065) );
  NAND2_X1 U5074 ( .A1(n4065), .A2(n4064), .ZN(n4332) );
  NOR4_X2 U5075 ( .A1(n5189), .A2(n5164), .A3(n4332), .A4(n5148), .ZN(n5128)
         );
  INV_X1 U5076 ( .A(n5469), .ZN(n5387) );
  OAI22_X1 U5077 ( .A1(n3902), .A2(n2963), .B1(n4069), .B2(n4233), .ZN(n4070)
         );
  INV_X1 U5078 ( .A(n4070), .ZN(n4080) );
  NAND2_X1 U5079 ( .A1(n3685), .A2(n4090), .ZN(n4071) );
  NAND2_X1 U5080 ( .A1(n4072), .A2(n4071), .ZN(n4075) );
  OR2_X1 U5081 ( .A1(n4073), .A2(n3071), .ZN(n4074) );
  NAND2_X1 U5082 ( .A1(n4075), .A2(n4074), .ZN(n4191) );
  AND2_X1 U5083 ( .A1(n4076), .A2(n4069), .ZN(n4533) );
  INV_X1 U5084 ( .A(n4077), .ZN(n4669) );
  NAND2_X2 U5085 ( .A1(n4669), .A2(n4090), .ZN(n4138) );
  OAI21_X1 U5086 ( .B1(n4533), .B2(n4489), .A(n4078), .ZN(n4079) );
  NAND4_X1 U5087 ( .A1(n4081), .A2(n4080), .A3(n4191), .A4(n4079), .ZN(n4542)
         );
  INV_X1 U5088 ( .A(n4088), .ZN(n5069) );
  NAND2_X1 U5089 ( .A1(n5069), .A2(n4083), .ZN(n4607) );
  INV_X1 U5090 ( .A(n4084), .ZN(n4085) );
  NAND2_X1 U5091 ( .A1(n4085), .A2(n4681), .ZN(n4086) );
  OAI211_X1 U5092 ( .C1(n4561), .C2(n3286), .A(n4607), .B(n4086), .ZN(n4087)
         );
  NOR2_X1 U5093 ( .A1(n4542), .A2(n4087), .ZN(n4238) );
  NOR2_X1 U5094 ( .A1(n4088), .A2(n4656), .ZN(n4190) );
  NAND2_X1 U5095 ( .A1(n4238), .A2(n4190), .ZN(n4592) );
  INV_X1 U5096 ( .A(n4089), .ZN(n4093) );
  NOR2_X1 U5097 ( .A1(n4566), .A2(n3273), .ZN(n4091) );
  NAND4_X1 U5098 ( .A1(n4093), .A2(n4092), .A3(n4549), .A4(n4091), .ZN(n4094)
         );
  OAI21_X1 U5099 ( .B1(n4531), .B2(n4592), .A(n4094), .ZN(n4095) );
  NAND2_X1 U5100 ( .A1(n4138), .A2(n6173), .ZN(n4097) );
  INV_X1 U5101 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U5102 ( .A1(n4549), .A2(n6068), .ZN(n4096) );
  NAND3_X1 U5103 ( .A1(n4097), .A2(n4068), .A3(n4096), .ZN(n4099) );
  NAND2_X1 U5104 ( .A1(n5224), .A2(n6068), .ZN(n4098) );
  NAND2_X1 U5105 ( .A1(n4099), .A2(n4098), .ZN(n5308) );
  NAND2_X1 U5106 ( .A1(n4585), .A2(n5308), .ZN(n4109) );
  NAND2_X1 U5107 ( .A1(n4138), .A2(n6269), .ZN(n4101) );
  INV_X1 U5108 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4571) );
  NAND2_X1 U5109 ( .A1(n4549), .A2(n4571), .ZN(n4100) );
  NAND3_X1 U5110 ( .A1(n4101), .A2(n4068), .A3(n4100), .ZN(n4103) );
  NAND2_X1 U5111 ( .A1(n5224), .A2(n4571), .ZN(n4102) );
  NAND2_X1 U5112 ( .A1(n4103), .A2(n4102), .ZN(n4106) );
  INV_X1 U5113 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U5114 ( .A1(n4068), .A2(n5327), .ZN(n4104) );
  NAND2_X1 U5115 ( .A1(n4105), .A2(n4104), .ZN(n4490) );
  XNOR2_X1 U5116 ( .A(n4106), .B(n4490), .ZN(n4548) );
  NAND2_X1 U5117 ( .A1(n4548), .A2(n4549), .ZN(n4551) );
  INV_X1 U5118 ( .A(n4106), .ZN(n4107) );
  NAND2_X1 U5119 ( .A1(n4107), .A2(n4490), .ZN(n4108) );
  NAND2_X1 U5120 ( .A1(n4551), .A2(n4108), .ZN(n4584) );
  MUX2_X1 U5121 ( .A(n2963), .B(n4138), .S(EBX_REG_4__SCAN_IN), .Z(n4111) );
  NAND2_X1 U5122 ( .A1(n4231), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4110)
         );
  NAND2_X1 U5123 ( .A1(n4111), .A2(n4110), .ZN(n4804) );
  NAND2_X1 U5124 ( .A1(n4587), .A2(n4804), .ZN(n4737) );
  MUX2_X1 U5125 ( .A(n4223), .B(n2963), .S(EBX_REG_5__SCAN_IN), .Z(n4112) );
  OAI21_X1 U5126 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4489), .A(n4112), 
        .ZN(n4738) );
  INV_X1 U5127 ( .A(n4738), .ZN(n4113) );
  NAND2_X1 U5128 ( .A1(n4138), .A2(n6236), .ZN(n4116) );
  INV_X1 U5129 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U5130 ( .A1(n4549), .A2(n6023), .ZN(n4115) );
  NAND3_X1 U5131 ( .A1(n4116), .A2(n2963), .A3(n4115), .ZN(n4118) );
  NAND2_X1 U5132 ( .A1(n5224), .A2(n6023), .ZN(n4117) );
  NAND2_X1 U5133 ( .A1(n2963), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4121)
         );
  OAI211_X1 U5134 ( .C1(n4231), .C2(EBX_REG_7__SCAN_IN), .A(n4138), .B(n4121), 
        .ZN(n4122) );
  OAI21_X1 U5135 ( .B1(n4223), .B2(EBX_REG_7__SCAN_IN), .A(n4122), .ZN(n5001)
         );
  MUX2_X1 U5136 ( .A(n4223), .B(n2963), .S(EBX_REG_9__SCAN_IN), .Z(n4124) );
  OR2_X1 U5137 ( .A1(n4489), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4123)
         );
  NAND2_X1 U5138 ( .A1(n4124), .A2(n4123), .ZN(n5057) );
  NAND2_X1 U5139 ( .A1(n4138), .A2(n4125), .ZN(n4127) );
  INV_X1 U5140 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U5141 ( .A1(n4549), .A2(n5291), .ZN(n4126) );
  NAND3_X1 U5142 ( .A1(n4127), .A2(n2963), .A3(n4126), .ZN(n4129) );
  NAND2_X1 U5143 ( .A1(n5224), .A2(n5291), .ZN(n4128) );
  MUX2_X1 U5144 ( .A(n2963), .B(n4138), .S(EBX_REG_10__SCAN_IN), .Z(n4131) );
  NAND2_X1 U5145 ( .A1(n4231), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4130) );
  NAND2_X1 U5146 ( .A1(n4131), .A2(n4130), .ZN(n5277) );
  NAND2_X1 U5147 ( .A1(n2963), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4132) );
  OAI211_X1 U5148 ( .C1(n4231), .C2(EBX_REG_11__SCAN_IN), .A(n4138), .B(n4132), 
        .ZN(n4133) );
  OAI21_X1 U5149 ( .B1(n4223), .B2(EBX_REG_11__SCAN_IN), .A(n4133), .ZN(n5986)
         );
  MUX2_X1 U5150 ( .A(n2963), .B(n4138), .S(EBX_REG_12__SCAN_IN), .Z(n4135) );
  NAND2_X1 U5151 ( .A1(n4231), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4134) );
  NAND2_X1 U5152 ( .A1(n4135), .A2(n4134), .ZN(n5364) );
  INV_X1 U5153 ( .A(n5364), .ZN(n4136) );
  NAND2_X1 U5154 ( .A1(n2963), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4137) );
  OAI211_X1 U5155 ( .C1(n4231), .C2(EBX_REG_13__SCAN_IN), .A(n4138), .B(n4137), 
        .ZN(n4139) );
  OAI21_X1 U5156 ( .B1(n4223), .B2(EBX_REG_13__SCAN_IN), .A(n4139), .ZN(n5917)
         );
  MUX2_X1 U5157 ( .A(n2963), .B(n4138), .S(EBX_REG_14__SCAN_IN), .Z(n4142) );
  NAND2_X1 U5158 ( .A1(n4231), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4141) );
  NAND2_X1 U5159 ( .A1(n4142), .A2(n4141), .ZN(n5360) );
  NAND2_X1 U5160 ( .A1(n2963), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4143) );
  OAI211_X1 U5161 ( .C1(n4231), .C2(EBX_REG_15__SCAN_IN), .A(n4138), .B(n4143), 
        .ZN(n4144) );
  OAI21_X1 U5162 ( .B1(n4223), .B2(EBX_REG_15__SCAN_IN), .A(n4144), .ZN(n5262)
         );
  MUX2_X1 U5163 ( .A(n2963), .B(n4138), .S(EBX_REG_16__SCAN_IN), .Z(n4146) );
  NAND2_X1 U5164 ( .A1(n4231), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4145) );
  INV_X1 U5165 ( .A(n4223), .ZN(n4161) );
  INV_X1 U5166 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5344) );
  NAND2_X1 U5167 ( .A1(n4161), .A2(n5344), .ZN(n4149) );
  NAND2_X1 U5168 ( .A1(n2963), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4147) );
  OAI211_X1 U5169 ( .C1(n4231), .C2(EBX_REG_17__SCAN_IN), .A(n4138), .B(n4147), 
        .ZN(n4148) );
  MUX2_X1 U5170 ( .A(n2963), .B(n4138), .S(EBX_REG_19__SCAN_IN), .Z(n4151) );
  NAND2_X1 U5171 ( .A1(n4231), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4150) );
  NAND2_X1 U5172 ( .A1(n4151), .A2(n4150), .ZN(n5227) );
  NAND2_X1 U5173 ( .A1(n5222), .A2(n5227), .ZN(n5211) );
  OR2_X1 U5174 ( .A1(n4489), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4152)
         );
  INV_X1 U5175 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U5176 ( .A1(n4549), .A2(n5343), .ZN(n5223) );
  OAI22_X1 U5177 ( .A1(n4489), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n4231), .ZN(n5213) );
  NAND2_X1 U5178 ( .A1(n5226), .A2(n5213), .ZN(n4154) );
  NAND2_X1 U5179 ( .A1(n5224), .A2(EBX_REG_20__SCAN_IN), .ZN(n4153) );
  OAI211_X1 U5180 ( .C1(n5226), .C2(n5224), .A(n4154), .B(n4153), .ZN(n4155)
         );
  MUX2_X1 U5181 ( .A(n4223), .B(n2963), .S(EBX_REG_21__SCAN_IN), .Z(n4158) );
  OAI21_X1 U5182 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n4489), .A(n4158), 
        .ZN(n4265) );
  MUX2_X1 U5183 ( .A(n2963), .B(n4138), .S(EBX_REG_22__SCAN_IN), .Z(n4160) );
  NAND2_X1 U5184 ( .A1(n4231), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4159) );
  NAND2_X1 U5185 ( .A1(n4160), .A2(n4159), .ZN(n5193) );
  INV_X1 U5186 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U5187 ( .A1(n4161), .A2(n5340), .ZN(n4164) );
  NAND2_X1 U5188 ( .A1(n2963), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4162) );
  OAI211_X1 U5189 ( .C1(n4231), .C2(EBX_REG_23__SCAN_IN), .A(n4138), .B(n4162), 
        .ZN(n4163) );
  INV_X1 U5190 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4165) );
  NAND2_X1 U5191 ( .A1(n4138), .A2(n4165), .ZN(n4166) );
  OAI211_X1 U5192 ( .C1(EBX_REG_24__SCAN_IN), .C2(n4231), .A(n4166), .B(n2963), 
        .ZN(n4169) );
  INV_X1 U5193 ( .A(EBX_REG_24__SCAN_IN), .ZN(n4167) );
  NAND2_X1 U5194 ( .A1(n5224), .A2(n4167), .ZN(n4168) );
  MUX2_X1 U5195 ( .A(n4223), .B(n2963), .S(EBX_REG_25__SCAN_IN), .Z(n4170) );
  OAI21_X1 U5196 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n4489), .A(n4170), 
        .ZN(n5149) );
  INV_X1 U5197 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4171) );
  NAND2_X1 U5198 ( .A1(n4138), .A2(n4171), .ZN(n4172) );
  OAI211_X1 U5199 ( .C1(EBX_REG_26__SCAN_IN), .C2(n4231), .A(n4172), .B(n2963), 
        .ZN(n4174) );
  INV_X1 U5200 ( .A(EBX_REG_26__SCAN_IN), .ZN(n4177) );
  NAND2_X1 U5201 ( .A1(n5224), .A2(n4177), .ZN(n4173) );
  NAND2_X1 U5202 ( .A1(n4174), .A2(n4173), .ZN(n4175) );
  OR2_X1 U5203 ( .A1(n5152), .A2(n4175), .ZN(n4176) );
  NAND2_X1 U5204 ( .A1(n4225), .A2(n4176), .ZN(n5626) );
  INV_X1 U5205 ( .A(n4566), .ZN(n5373) );
  AND2_X1 U5206 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5490) );
  AND2_X1 U5207 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5674) );
  AND2_X1 U5208 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4258) );
  NAND3_X1 U5209 ( .A1(n5490), .A2(n5674), .A3(n4258), .ZN(n4180) );
  NOR2_X1 U5210 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5657) );
  NOR2_X1 U5211 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4379) );
  NOR2_X1 U5212 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5673) );
  AND3_X1 U5213 ( .A1(n5657), .A2(n4379), .A3(n5673), .ZN(n4181) );
  XNOR2_X1 U5214 ( .A(n6146), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5473)
         );
  INV_X1 U5215 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5640) );
  INV_X1 U5216 ( .A(n5464), .ZN(n4184) );
  NAND2_X1 U5217 ( .A1(n6146), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5463) );
  INV_X1 U5218 ( .A(n5463), .ZN(n4183) );
  NAND2_X1 U5219 ( .A1(n4184), .A2(n4183), .ZN(n5434) );
  NAND2_X1 U5220 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5435) );
  INV_X1 U5221 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5589) );
  INV_X1 U5222 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5592) );
  NOR2_X1 U5223 ( .A1(n5533), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5462)
         );
  INV_X1 U5224 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6756) );
  INV_X1 U5225 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5444) );
  NAND3_X1 U5226 ( .A1(n5426), .A2(n5592), .A3(n5589), .ZN(n4187) );
  NAND2_X1 U5227 ( .A1(n4188), .A2(n4187), .ZN(n4189) );
  XNOR2_X1 U5228 ( .A(n4189), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4394)
         );
  INV_X1 U5229 ( .A(n4190), .ZN(n4207) );
  NAND2_X1 U5230 ( .A1(n4219), .A2(n4191), .ZN(n4194) );
  NAND2_X1 U5231 ( .A1(n4194), .A2(n4193), .ZN(n4535) );
  INV_X1 U5232 ( .A(n4195), .ZN(n4197) );
  INV_X1 U5233 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4196) );
  NAND2_X1 U5234 ( .A1(n4197), .A2(n4196), .ZN(n6603) );
  NAND2_X1 U5235 ( .A1(n4237), .A2(n6603), .ZN(n4205) );
  NAND3_X1 U5236 ( .A1(n4200), .A2(n4199), .A3(n4198), .ZN(n4201) );
  NAND2_X1 U5237 ( .A1(n4202), .A2(n4201), .ZN(n4204) );
  NOR2_X1 U5238 ( .A1(n4447), .A2(READY_N), .ZN(n4559) );
  NAND3_X1 U5239 ( .A1(n4205), .A2(n4559), .A3(n4212), .ZN(n4206) );
  OAI211_X1 U5240 ( .C1(n4531), .C2(n4207), .A(n4535), .B(n4206), .ZN(n4208)
         );
  NAND2_X1 U5241 ( .A1(n4208), .A2(n6511), .ZN(n4215) );
  NAND2_X1 U5242 ( .A1(n4656), .A2(n6603), .ZN(n4401) );
  NAND2_X1 U5243 ( .A1(n4401), .A2(n6606), .ZN(n4210) );
  OAI211_X1 U5244 ( .C1(n4540), .C2(n4210), .A(n4090), .B(n5100), .ZN(n4211)
         );
  INV_X1 U5245 ( .A(n4211), .ZN(n4213) );
  OAI22_X1 U5246 ( .A1(n3274), .A2(n4216), .B1(n4540), .B2(n4231), .ZN(n4217)
         );
  INV_X1 U5247 ( .A(n4217), .ZN(n4220) );
  INV_X1 U5248 ( .A(n4564), .ZN(n4591) );
  AND4_X1 U5249 ( .A1(n5927), .A2(n4220), .A3(n4591), .A4(n6481), .ZN(n4221)
         );
  AND2_X1 U5250 ( .A1(n4231), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4222)
         );
  MUX2_X1 U5251 ( .A(n4223), .B(n2963), .S(EBX_REG_27__SCAN_IN), .Z(n4224) );
  OAI21_X1 U5252 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n4489), .A(n4224), 
        .ZN(n5130) );
  NAND2_X1 U5253 ( .A1(n4138), .A2(n5444), .ZN(n4226) );
  OAI211_X1 U5254 ( .C1(EBX_REG_28__SCAN_IN), .C2(n4231), .A(n4226), .B(n2963), 
        .ZN(n4228) );
  INV_X1 U5255 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U5256 ( .A1(n5224), .A2(n5334), .ZN(n4227) );
  AND2_X1 U5257 ( .A1(n4228), .A2(n4227), .ZN(n5118) );
  OAI22_X1 U5258 ( .A1(n4489), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n4231), .ZN(n4431) );
  NAND2_X1 U5259 ( .A1(n4364), .A2(n2963), .ZN(n4229) );
  INV_X1 U5260 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U5261 ( .A1(n5224), .A2(n5333), .ZN(n4430) );
  NOR2_X1 U5262 ( .A1(n4364), .A2(n5224), .ZN(n4370) );
  AOI21_X1 U5263 ( .B1(n4365), .B2(n4429), .A(n4370), .ZN(n4230) );
  OAI22_X1 U5264 ( .A1(n4489), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4231), .ZN(n4232) );
  NAND2_X1 U5265 ( .A1(n4209), .A2(n6605), .ZN(n6492) );
  NAND2_X1 U5266 ( .A1(n4233), .A2(n3274), .ZN(n4234) );
  OR2_X1 U5267 ( .A1(n4561), .A2(n4234), .ZN(n4235) );
  AND2_X1 U5268 ( .A1(n6492), .A2(n4235), .ZN(n4236) );
  NAND2_X1 U5269 ( .A1(n4192), .A2(n4237), .ZN(n5073) );
  OR2_X1 U5270 ( .A1(n4239), .A2(n4238), .ZN(n4250) );
  NAND2_X1 U5271 ( .A1(n6200), .A2(n4250), .ZN(n4240) );
  INV_X1 U5272 ( .A(n4240), .ZN(n5737) );
  INV_X1 U5273 ( .A(n5435), .ZN(n5611) );
  INV_X1 U5274 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U5275 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6259) );
  OR3_X1 U5276 ( .A1(n3762), .A2(n6256), .A3(n6259), .ZN(n4740) );
  NAND2_X1 U5277 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4241) );
  OR2_X1 U5278 ( .A1(n4740), .A2(n4241), .ZN(n6194) );
  INV_X1 U5279 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6710) );
  NAND2_X1 U5280 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6213) );
  OR3_X1 U5281 ( .A1(n6710), .A2(n6735), .A3(n6213), .ZN(n4242) );
  NOR2_X1 U5282 ( .A1(n6194), .A2(n4242), .ZN(n4249) );
  AND2_X1 U5283 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5736) );
  AND2_X1 U5284 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5736), .ZN(n5741)
         );
  NAND2_X1 U5285 ( .A1(n5741), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4254) );
  NOR2_X1 U5286 ( .A1(n4255), .A2(n4254), .ZN(n4243) );
  NAND2_X1 U5287 ( .A1(n4249), .A2(n4243), .ZN(n5680) );
  INV_X1 U5288 ( .A(n6233), .ZN(n6248) );
  NAND2_X1 U5289 ( .A1(n4239), .A2(n6248), .ZN(n4488) );
  INV_X1 U5290 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U5291 ( .A1(n6260), .A2(n4240), .ZN(n4493) );
  NAND2_X1 U5292 ( .A1(n4488), .A2(n4493), .ZN(n4730) );
  NOR2_X1 U5293 ( .A1(n6264), .A2(n4730), .ZN(n5712) );
  INV_X1 U5294 ( .A(n5712), .ZN(n6191) );
  OAI21_X1 U5295 ( .B1(n6269), .B2(n6260), .A(n6173), .ZN(n6258) );
  NAND3_X1 U5296 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n6258), .ZN(n4733) );
  NOR2_X1 U5297 ( .A1(n4241), .A2(n4733), .ZN(n6201) );
  AND2_X1 U5298 ( .A1(n5713), .A2(n4243), .ZN(n5678) );
  INV_X1 U5299 ( .A(n4244), .ZN(n5672) );
  NAND2_X1 U5300 ( .A1(n5672), .A2(n5674), .ZN(n4257) );
  INV_X1 U5301 ( .A(n4257), .ZN(n5489) );
  NAND2_X1 U5302 ( .A1(n5738), .A2(n4250), .ZN(n6193) );
  OR2_X1 U5303 ( .A1(n6193), .A2(n6191), .ZN(n4245) );
  INV_X1 U5304 ( .A(n5490), .ZN(n5659) );
  NAND2_X1 U5305 ( .A1(n6196), .A2(n5659), .ZN(n4246) );
  NAND2_X1 U5306 ( .A1(n5653), .A2(n4246), .ZN(n5644) );
  NAND2_X1 U5307 ( .A1(n5738), .A2(n6260), .ZN(n4553) );
  NAND2_X1 U5308 ( .A1(n6193), .A2(n4553), .ZN(n6268) );
  AND2_X1 U5309 ( .A1(n6200), .A2(n6268), .ZN(n4247) );
  NAND2_X1 U5310 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5630) );
  AND2_X1 U5311 ( .A1(n6196), .A2(n5630), .ZN(n4248) );
  OAI21_X1 U5312 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5718), .A(n5593), 
        .ZN(n4260) );
  AND2_X1 U5313 ( .A1(n6233), .A2(REIP_REG_31__SCAN_IN), .ZN(n4390) );
  INV_X1 U5314 ( .A(n4249), .ZN(n5714) );
  NOR2_X1 U5315 ( .A1(n5714), .A2(n4250), .ZN(n4251) );
  AND2_X1 U5316 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n4251), .ZN(n4252)
         );
  INV_X1 U5317 ( .A(n4254), .ZN(n5717) );
  INV_X1 U5318 ( .A(n4255), .ZN(n4256) );
  NAND2_X1 U5319 ( .A1(n5650), .A2(n4258), .ZN(n5629) );
  NAND2_X1 U5320 ( .A1(n5623), .A2(n5611), .ZN(n5603) );
  NOR4_X1 U5321 ( .A1(n5603), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5589), 
        .A4(n5592), .ZN(n4259) );
  AOI211_X1 U5322 ( .C1(INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n4260), .A(n4390), .B(n4259), .ZN(n4261) );
  OAI21_X1 U5323 ( .B1(n4394), .B2(n6184), .A(n4262), .ZN(U2987) );
  AND2_X1 U5324 ( .A1(n4266), .A2(n4265), .ZN(n4267) );
  OR2_X1 U5325 ( .A1(n4267), .A2(n2976), .ZN(n5663) );
  INV_X1 U5326 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5204) );
  INV_X1 U5327 ( .A(n4337), .ZN(n4271) );
  INV_X1 U5328 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4420) );
  INV_X1 U5329 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5104) );
  XNOR2_X1 U5330 ( .A(n4387), .B(n5104), .ZN(n5430) );
  AOI22_X1 U5331 ( .A1(n4310), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4275) );
  AOI22_X1 U5332 ( .A1(n4311), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4274) );
  AOI22_X1 U5333 ( .A1(n4317), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4273) );
  AOI22_X1 U5334 ( .A1(n3499), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4272) );
  NAND4_X1 U5335 ( .A1(n4275), .A2(n4274), .A3(n4273), .A4(n4272), .ZN(n4281)
         );
  AOI22_X1 U5336 ( .A1(n4308), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4279) );
  AOI22_X1 U5337 ( .A1(n3469), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4278) );
  AOI22_X1 U5338 ( .A1(n3356), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4277) );
  AOI22_X1 U5339 ( .A1(n4288), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4276) );
  NAND4_X1 U5340 ( .A1(n4279), .A2(n4278), .A3(n4277), .A4(n4276), .ZN(n4280)
         );
  NOR2_X1 U5341 ( .A1(n4281), .A2(n4280), .ZN(n4327) );
  AOI22_X1 U5342 ( .A1(n4282), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4287) );
  AOI22_X1 U5343 ( .A1(n4311), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4286) );
  AOI22_X1 U5344 ( .A1(n4317), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4285) );
  AOI22_X1 U5345 ( .A1(n3356), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4283), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4284) );
  NAND4_X1 U5346 ( .A1(n4287), .A2(n4286), .A3(n4285), .A4(n4284), .ZN(n4294)
         );
  AOI22_X1 U5347 ( .A1(n4308), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4292) );
  AOI22_X1 U5348 ( .A1(n4309), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4291) );
  AOI22_X1 U5349 ( .A1(n3475), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4290) );
  AOI22_X1 U5350 ( .A1(n4288), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4289) );
  NAND4_X1 U5351 ( .A1(n4292), .A2(n4291), .A3(n4290), .A4(n4289), .ZN(n4293)
         );
  NOR2_X1 U5352 ( .A1(n4294), .A2(n4293), .ZN(n4352) );
  AOI22_X1 U5353 ( .A1(n4308), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4298) );
  AOI22_X1 U5354 ( .A1(n4310), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4297) );
  AOI22_X1 U5355 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n4309), .B1(n4316), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4296) );
  AOI22_X1 U5356 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4288), .B1(n3569), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4295) );
  NAND4_X1 U5357 ( .A1(n4298), .A2(n4297), .A3(n4296), .A4(n4295), .ZN(n4304)
         );
  AOI22_X1 U5358 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4311), .B1(n4307), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4302) );
  AOI22_X1 U5359 ( .A1(n3356), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4301) );
  AOI22_X1 U5360 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3362), .B1(n4318), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4300) );
  AOI22_X1 U5361 ( .A1(n3475), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4299) );
  NAND4_X1 U5362 ( .A1(n4302), .A2(n4301), .A3(n4300), .A4(n4299), .ZN(n4303)
         );
  NOR2_X1 U5363 ( .A1(n4304), .A2(n4303), .ZN(n4333) );
  NAND2_X1 U5364 ( .A1(n4306), .A2(n4305), .ZN(n4334) );
  NOR2_X1 U5365 ( .A1(n4333), .A2(n4334), .ZN(n4346) );
  AOI22_X1 U5366 ( .A1(n4308), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4315) );
  AOI22_X1 U5367 ( .A1(n3469), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4314) );
  AOI22_X1 U5368 ( .A1(n4310), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4309), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4313) );
  AOI22_X1 U5369 ( .A1(n4311), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4312) );
  NAND4_X1 U5370 ( .A1(n4315), .A2(n4314), .A3(n4313), .A4(n4312), .ZN(n4325)
         );
  AOI22_X1 U5371 ( .A1(n4317), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4323) );
  AOI22_X1 U5372 ( .A1(n3356), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4322) );
  AOI22_X1 U5373 ( .A1(n3475), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3569), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4321) );
  AOI22_X1 U5374 ( .A1(n4288), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4320) );
  NAND4_X1 U5375 ( .A1(n4323), .A2(n4322), .A3(n4321), .A4(n4320), .ZN(n4324)
         );
  OR2_X1 U5376 ( .A1(n4325), .A2(n4324), .ZN(n4345) );
  NAND2_X1 U5377 ( .A1(n4346), .A2(n4345), .ZN(n4353) );
  NOR2_X1 U5378 ( .A1(n4352), .A2(n4353), .ZN(n4326) );
  XOR2_X1 U5379 ( .A(n4327), .B(n4326), .Z(n4330) );
  AOI21_X1 U5380 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6409), .A(n5183), 
        .ZN(n4329) );
  NAND2_X1 U5381 ( .A1(n4357), .A2(EAX_REG_30__SCAN_IN), .ZN(n4328) );
  OAI211_X1 U5382 ( .C1(n4330), .C2(n4349), .A(n4329), .B(n4328), .ZN(n4331)
         );
  OAI21_X1 U5383 ( .B1(n3492), .B2(n5430), .A(n4331), .ZN(n4362) );
  INV_X1 U5384 ( .A(n5189), .ZN(n4343) );
  INV_X1 U5385 ( .A(n4332), .ZN(n4342) );
  XOR2_X1 U5386 ( .A(n4334), .B(n4333), .Z(n4335) );
  NAND2_X1 U5387 ( .A1(n4335), .A2(n4354), .ZN(n4339) );
  INV_X1 U5388 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5133) );
  NOR2_X1 U5389 ( .A1(n5133), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4336) );
  AOI211_X1 U5390 ( .C1(n4357), .C2(EAX_REG_27__SCAN_IN), .A(n5183), .B(n4336), 
        .ZN(n4338) );
  XNOR2_X1 U5391 ( .A(n4337), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5132)
         );
  AOI22_X1 U5392 ( .A1(n4339), .A2(n4338), .B1(n5183), .B2(n5132), .ZN(n5127)
         );
  INV_X1 U5393 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6734) );
  NAND2_X1 U5394 ( .A1(n2997), .A2(n6734), .ZN(n4344) );
  NAND2_X1 U5395 ( .A1(n4358), .A2(n4344), .ZN(n5450) );
  XNOR2_X1 U5396 ( .A(n4346), .B(n4345), .ZN(n4350) );
  NOR2_X1 U5397 ( .A1(n6734), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4347) );
  AOI211_X1 U5398 ( .C1(n4357), .C2(EAX_REG_28__SCAN_IN), .A(n5183), .B(n4347), 
        .ZN(n4348) );
  OAI21_X1 U5399 ( .B1(n4350), .B2(n4349), .A(n4348), .ZN(n4351) );
  XOR2_X1 U5400 ( .A(n4353), .B(n4352), .Z(n4355) );
  NAND2_X1 U5401 ( .A1(n4355), .A2(n4354), .ZN(n4360) );
  NOR2_X1 U5402 ( .A1(n4420), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4356) );
  AOI211_X1 U5403 ( .C1(n4357), .C2(EAX_REG_29__SCAN_IN), .A(n5183), .B(n4356), 
        .ZN(n4359) );
  XNOR2_X1 U5404 ( .A(n4358), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4419)
         );
  AOI22_X1 U5405 ( .A1(n4360), .A2(n4359), .B1(n5183), .B2(n4419), .ZN(n4396)
         );
  INV_X1 U5406 ( .A(n5432), .ZN(n5377) );
  INV_X1 U5407 ( .A(n4365), .ZN(n4363) );
  OAI21_X1 U5408 ( .B1(n4364), .B2(n5120), .A(n4363), .ZN(n4369) );
  INV_X1 U5409 ( .A(n5120), .ZN(n4367) );
  INV_X1 U5410 ( .A(n4364), .ZN(n4366) );
  OAI211_X1 U5411 ( .C1(n4367), .C2(n4068), .A(n4366), .B(n4365), .ZN(n4368)
         );
  OAI21_X1 U5412 ( .B1(n4370), .B2(n4369), .A(n4368), .ZN(n5103) );
  INV_X1 U5413 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4371) );
  OAI22_X1 U5414 ( .A1(n5103), .A2(n5369), .B1(n4371), .B2(n6067), .ZN(n4372)
         );
  INV_X1 U5415 ( .A(n4372), .ZN(n4373) );
  XNOR2_X1 U5416 ( .A(n6146), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5507)
         );
  NOR2_X1 U5417 ( .A1(n5533), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5498)
         );
  NAND2_X1 U5418 ( .A1(n4376), .A2(n4377), .ZN(n4378) );
  AND2_X1 U5419 ( .A1(n5150), .A2(n4378), .ZN(n5338) );
  AND2_X1 U5420 ( .A1(n6233), .A2(REIP_REG_24__SCAN_IN), .ZN(n5480) );
  AOI21_X1 U5421 ( .B1(n5338), .B2(n6262), .A(n5480), .ZN(n4382) );
  INV_X1 U5422 ( .A(n4379), .ZN(n4380) );
  OAI211_X1 U5423 ( .C1(n5650), .C2(INSTADDRPOINTER_REG_24__SCAN_IN), .A(n5634), .B(n4380), .ZN(n4381) );
  OAI21_X1 U5424 ( .B1(n5486), .B2(n6184), .A(n4383), .ZN(U2994) );
  AOI22_X1 U5425 ( .A1(n3418), .A2(EAX_REG_31__SCAN_IN), .B1(n4384), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4385) );
  XNOR2_X1 U5426 ( .A(n4386), .B(n4385), .ZN(n5099) );
  NAND2_X1 U5427 ( .A1(n4388), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4389)
         );
  INV_X1 U5428 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5092) );
  AOI21_X1 U5429 ( .B1(n5565), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n4390), 
        .ZN(n4391) );
  OAI21_X1 U5430 ( .B1(n6182), .B2(n4418), .A(n4391), .ZN(n4392) );
  AOI21_X1 U5431 ( .B1(n5099), .B2(n6177), .A(n4392), .ZN(n4393) );
  OAI21_X1 U5432 ( .B1(n4394), .B2(n6159), .A(n4393), .ZN(U2955) );
  NOR2_X1 U5433 ( .A1(n4193), .A2(n4447), .ZN(n4439) );
  NAND2_X1 U5434 ( .A1(n4439), .A2(n6511), .ZN(n4453) );
  NAND2_X1 U5435 ( .A1(n6749), .A2(n5874), .ZN(n6503) );
  NOR3_X1 U5436 ( .A1(n6509), .A2(n6588), .A3(n6503), .ZN(n6500) );
  AND2_X1 U5437 ( .A1(n4397), .A2(n5183), .ZN(n6508) );
  NAND2_X1 U5438 ( .A1(n6606), .A2(n6604), .ZN(n4434) );
  INV_X1 U5439 ( .A(n4434), .ZN(n4400) );
  NAND3_X1 U5440 ( .A1(n4401), .A2(n4090), .A3(n4400), .ZN(n4402) );
  OR2_X2 U5441 ( .A1(n5310), .A2(n4402), .ZN(n5980) );
  INV_X2 U5442 ( .A(n5980), .ZN(n6775) );
  INV_X1 U5443 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6784) );
  INV_X1 U5444 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6667) );
  INV_X1 U5445 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6740) );
  NAND3_X1 U5446 ( .A1(REIP_REG_3__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6031) );
  NOR3_X1 U5447 ( .A1(n6667), .A2(n6740), .A3(n6031), .ZN(n5272) );
  NAND2_X1 U5448 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_8__SCAN_IN), .ZN(
        n5283) );
  INV_X1 U5449 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6538) );
  NOR2_X1 U5450 ( .A1(n5283), .A2(n6538), .ZN(n5275) );
  INV_X1 U5451 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6542) );
  INV_X1 U5452 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6543) );
  NOR2_X1 U5453 ( .A1(n6542), .A2(n6543), .ZN(n5985) );
  NAND4_X1 U5454 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5272), .A3(n5275), .A4(
        n5985), .ZN(n6773) );
  NOR2_X1 U5455 ( .A1(n6784), .A2(n6773), .ZN(n4407) );
  NAND2_X1 U5456 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .ZN(
        n4403) );
  AND2_X1 U5457 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n4404) );
  NAND2_X1 U5458 ( .A1(n5960), .A2(n4404), .ZN(n5250) );
  INV_X1 U5459 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U5460 ( .A1(REIP_REG_18__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .ZN(
        n5233) );
  INV_X1 U5461 ( .A(n5233), .ZN(n5191) );
  NAND2_X1 U5462 ( .A1(n5191), .A2(REIP_REG_20__SCAN_IN), .ZN(n4405) );
  NOR2_X2 U5463 ( .A1(n5244), .A2(n4405), .ZN(n5201) );
  AND2_X1 U5464 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5171) );
  NAND2_X1 U5465 ( .A1(n5171), .A2(REIP_REG_23__SCAN_IN), .ZN(n4409) );
  INV_X1 U5466 ( .A(n4409), .ZN(n4406) );
  NAND2_X1 U5467 ( .A1(n5201), .A2(n4406), .ZN(n5167) );
  NAND3_X1 U5468 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4412) );
  NOR2_X1 U5469 ( .A1(n5167), .A2(n4412), .ZN(n5129) );
  NAND3_X1 U5470 ( .A1(n5129), .A2(REIP_REG_27__SCAN_IN), .A3(
        REIP_REG_28__SCAN_IN), .ZN(n5105) );
  NAND2_X1 U5471 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n4408) );
  NAND4_X1 U5472 ( .A1(n4407), .A2(REIP_REG_14__SCAN_IN), .A3(
        REIP_REG_13__SCAN_IN), .A4(n5307), .ZN(n5965) );
  NOR3_X1 U5473 ( .A1(n6554), .A2(n4408), .A3(n5965), .ZN(n5221) );
  AND2_X1 U5474 ( .A1(n5221), .A2(REIP_REG_20__SCAN_IN), .ZN(n5192) );
  NOR2_X1 U5475 ( .A1(n4409), .A2(n5233), .ZN(n4410) );
  NAND2_X1 U5476 ( .A1(n5192), .A2(n4410), .ZN(n4411) );
  NAND2_X1 U5477 ( .A1(n4411), .A2(n6030), .ZN(n5181) );
  NAND2_X1 U5478 ( .A1(n6030), .A2(n4412), .ZN(n4413) );
  NAND2_X1 U5479 ( .A1(n5181), .A2(n4413), .ZN(n5146) );
  AND2_X1 U5480 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4414) );
  NOR2_X1 U5481 ( .A1(n5980), .A2(n4414), .ZN(n4415) );
  INV_X1 U5482 ( .A(n5116), .ZN(n4416) );
  MUX2_X1 U5483 ( .A(n5105), .B(n4416), .S(REIP_REG_29__SCAN_IN), .Z(n4417) );
  INV_X1 U5484 ( .A(n4419), .ZN(n5438) );
  OAI22_X1 U5485 ( .A1(n4420), .A2(n6047), .B1(n6778), .B2(n5438), .ZN(n4425)
         );
  NOR3_X1 U5486 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .A3(n6603), .ZN(
        n6495) );
  INV_X1 U5487 ( .A(n6495), .ZN(n4421) );
  AND2_X1 U5488 ( .A1(n6605), .A2(n4421), .ZN(n5090) );
  INV_X1 U5489 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5081) );
  AND3_X1 U5490 ( .A1(n4090), .A2(n5081), .A3(n4434), .ZN(n4422) );
  NOR2_X1 U5491 ( .A1(n5090), .A2(n4422), .ZN(n4423) );
  INV_X1 U5492 ( .A(n4428), .ZN(n4436) );
  INV_X1 U5493 ( .A(n4429), .ZN(n4433) );
  OAI211_X1 U5494 ( .C1(n5224), .C2(n4431), .A(n5120), .B(n4430), .ZN(n4432)
         );
  NAND2_X1 U5495 ( .A1(n4433), .A2(n4432), .ZN(n5599) );
  NAND3_X1 U5496 ( .A1(n4549), .A2(EBX_REG_31__SCAN_IN), .A3(n4434), .ZN(n4435) );
  INV_X1 U5497 ( .A(n5229), .ZN(n4437) );
  NAND2_X1 U5498 ( .A1(n4456), .A2(n4437), .ZN(n4452) );
  AOI21_X1 U5499 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n4453), .A(n4452), .ZN(
        n4438) );
  INV_X1 U5500 ( .A(n4438), .ZN(U2788) );
  OR2_X1 U5501 ( .A1(n4531), .A2(n4218), .ZN(n4442) );
  INV_X1 U5502 ( .A(n4439), .ZN(n4440) );
  NAND2_X1 U5503 ( .A1(n4440), .A2(n4444), .ZN(n4441) );
  NAND2_X1 U5504 ( .A1(n4442), .A2(n4441), .ZN(n5933) );
  OR2_X1 U5505 ( .A1(n6605), .A2(n4076), .ZN(n6602) );
  AOI21_X1 U5506 ( .B1(n6602), .B2(n6603), .A(READY_N), .ZN(n4443) );
  OR2_X1 U5507 ( .A1(n5933), .A2(n4443), .ZN(n6483) );
  AND2_X1 U5508 ( .A1(n6483), .A2(n6511), .ZN(n5940) );
  INV_X1 U5509 ( .A(MORE_REG_SCAN_IN), .ZN(n4451) );
  NAND2_X1 U5510 ( .A1(n6481), .A2(n4444), .ZN(n4445) );
  NOR2_X1 U5511 ( .A1(n4445), .A2(n4564), .ZN(n4446) );
  MUX2_X1 U5512 ( .A(n4446), .B(n4592), .S(n4531), .Z(n4449) );
  NAND2_X1 U5513 ( .A1(n4192), .A2(n4447), .ZN(n4448) );
  NAND2_X1 U5514 ( .A1(n4449), .A2(n4448), .ZN(n6485) );
  NAND2_X1 U5515 ( .A1(n5940), .A2(n6485), .ZN(n4450) );
  OAI21_X1 U5516 ( .B1(n5940), .B2(n4451), .A(n4450), .ZN(U3471) );
  NOR2_X1 U5517 ( .A1(n4452), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4454) );
  AND2_X1 U5518 ( .A1(n4454), .A2(n4453), .ZN(n4455) );
  OAI22_X1 U5519 ( .A1(n4455), .A2(n6602), .B1(n4454), .B2(n6599), .ZN(U3474)
         );
  INV_X1 U5520 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4459) );
  AND2_X2 U5521 ( .A1(n4457), .A2(n6142), .ZN(n6140) );
  INV_X1 U5522 ( .A(DATAI_15_), .ZN(n6753) );
  INV_X1 U5523 ( .A(EAX_REG_15__SCAN_IN), .ZN(n4458) );
  OAI222_X1 U5524 ( .A1(n4459), .A2(n6118), .B1(n6125), .B2(n6753), .C1(n4458), 
        .C2(n6142), .ZN(U2954) );
  AOI22_X1 U5525 ( .A1(n6140), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6136), .ZN(n4460) );
  INV_X1 U5526 ( .A(DATAI_6_), .ZN(n4661) );
  OR2_X1 U5527 ( .A1(n6125), .A2(n4661), .ZN(n4463) );
  NAND2_X1 U5528 ( .A1(n4460), .A2(n4463), .ZN(U2945) );
  AOI22_X1 U5529 ( .A1(n6140), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n6136), .ZN(n4461) );
  INV_X1 U5530 ( .A(DATAI_14_), .ZN(n6757) );
  OR2_X1 U5531 ( .A1(n6125), .A2(n6757), .ZN(n4465) );
  NAND2_X1 U5532 ( .A1(n4461), .A2(n4465), .ZN(U2953) );
  AOI22_X1 U5533 ( .A1(n6140), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6136), .ZN(n4462) );
  INV_X1 U5534 ( .A(DATAI_7_), .ZN(n4674) );
  OR2_X1 U5535 ( .A1(n6125), .A2(n4674), .ZN(n4467) );
  NAND2_X1 U5536 ( .A1(n4462), .A2(n4467), .ZN(U2931) );
  AOI22_X1 U5537 ( .A1(n6140), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6136), .ZN(n4464) );
  NAND2_X1 U5538 ( .A1(n4464), .A2(n4463), .ZN(U2930) );
  AOI22_X1 U5539 ( .A1(n6140), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n6136), .ZN(n4466) );
  NAND2_X1 U5540 ( .A1(n4466), .A2(n4465), .ZN(U2938) );
  AOI22_X1 U5541 ( .A1(n6140), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6136), .ZN(n4468) );
  NAND2_X1 U5542 ( .A1(n4468), .A2(n4467), .ZN(U2946) );
  AOI22_X1 U5543 ( .A1(n6140), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6136), .ZN(n4469) );
  NAND2_X1 U5544 ( .A1(n6122), .A2(DATAI_0_), .ZN(n4470) );
  NAND2_X1 U5545 ( .A1(n4469), .A2(n4470), .ZN(U2939) );
  AOI22_X1 U5546 ( .A1(n6140), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6136), .ZN(n4471) );
  NAND2_X1 U5547 ( .A1(n4471), .A2(n4470), .ZN(U2924) );
  AOI22_X1 U5548 ( .A1(n6140), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6136), .ZN(n4472) );
  NAND2_X1 U5549 ( .A1(n6122), .A2(DATAI_1_), .ZN(n4474) );
  NAND2_X1 U5550 ( .A1(n4472), .A2(n4474), .ZN(U2940) );
  AOI22_X1 U5551 ( .A1(n6140), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6136), .ZN(n4473) );
  NAND2_X1 U5552 ( .A1(n6122), .A2(DATAI_2_), .ZN(n4481) );
  NAND2_X1 U5553 ( .A1(n4473), .A2(n4481), .ZN(U2941) );
  AOI22_X1 U5554 ( .A1(n6140), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n6136), .ZN(n4475) );
  NAND2_X1 U5555 ( .A1(n4475), .A2(n4474), .ZN(U2925) );
  AOI22_X1 U5556 ( .A1(n6140), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6136), .ZN(n4476) );
  NAND2_X1 U5557 ( .A1(n6122), .A2(DATAI_3_), .ZN(n4483) );
  NAND2_X1 U5558 ( .A1(n4476), .A2(n4483), .ZN(U2927) );
  AOI22_X1 U5559 ( .A1(n6140), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6136), .ZN(n4477) );
  NAND2_X1 U5560 ( .A1(n6122), .A2(DATAI_4_), .ZN(n4479) );
  NAND2_X1 U5561 ( .A1(n4477), .A2(n4479), .ZN(U2943) );
  AOI22_X1 U5562 ( .A1(n6140), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6136), .ZN(n4478) );
  NAND2_X1 U5563 ( .A1(n6122), .A2(DATAI_5_), .ZN(n4485) );
  NAND2_X1 U5564 ( .A1(n4478), .A2(n4485), .ZN(U2944) );
  AOI22_X1 U5565 ( .A1(n6140), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6136), .ZN(n4480) );
  NAND2_X1 U5566 ( .A1(n4480), .A2(n4479), .ZN(U2928) );
  AOI22_X1 U5567 ( .A1(n6140), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6136), .ZN(n4482) );
  NAND2_X1 U5568 ( .A1(n4482), .A2(n4481), .ZN(U2926) );
  AOI22_X1 U5569 ( .A1(n6140), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6136), .ZN(n4484) );
  NAND2_X1 U5570 ( .A1(n4484), .A2(n4483), .ZN(U2942) );
  AOI22_X1 U5571 ( .A1(n6140), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6136), .ZN(n4486) );
  NAND2_X1 U5572 ( .A1(n4486), .A2(n4485), .ZN(U2929) );
  XOR2_X1 U5573 ( .A(n4487), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n4525) );
  AOI21_X1 U5574 ( .B1(n5738), .B2(n4488), .A(n6260), .ZN(n4495) );
  OR2_X1 U5575 ( .A1(n4489), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4491)
         );
  NAND2_X1 U5576 ( .A1(n4491), .A2(n4490), .ZN(n5326) );
  AND2_X1 U5577 ( .A1(n6233), .A2(REIP_REG_0__SCAN_IN), .ZN(n4524) );
  INV_X1 U5578 ( .A(n4524), .ZN(n4492) );
  OAI211_X1 U5579 ( .C1(n6250), .C2(n5326), .A(n4493), .B(n4492), .ZN(n4494)
         );
  AOI211_X1 U5580 ( .C1(n4525), .C2(n6266), .A(n4495), .B(n4494), .ZN(n4496)
         );
  INV_X1 U5581 ( .A(n4496), .ZN(U3018) );
  INV_X1 U5582 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4499) );
  INV_X1 U5583 ( .A(n4627), .ZN(n4629) );
  AOI22_X1 U5584 ( .A1(UWORD_REG_14__SCAN_IN), .A2(n6601), .B1(n6112), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4498) );
  OAI21_X1 U5585 ( .B1(n4499), .B2(n6079), .A(n4498), .ZN(U2893) );
  INV_X1 U5586 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4501) );
  AOI22_X1 U5587 ( .A1(UWORD_REG_10__SCAN_IN), .A2(n6601), .B1(n6112), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4500) );
  OAI21_X1 U5588 ( .B1(n4501), .B2(n6079), .A(n4500), .ZN(U2897) );
  INV_X1 U5589 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4503) );
  AOI22_X1 U5590 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n6601), .B1(n6112), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4502) );
  OAI21_X1 U5591 ( .B1(n4503), .B2(n6079), .A(n4502), .ZN(U2895) );
  INV_X1 U5592 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4505) );
  AOI22_X1 U5593 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n6085), .B1(n6112), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4504) );
  OAI21_X1 U5594 ( .B1(n4505), .B2(n6079), .A(n4504), .ZN(U2904) );
  INV_X1 U5595 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4507) );
  AOI22_X1 U5596 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n6085), .B1(n6112), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4506) );
  OAI21_X1 U5597 ( .B1(n4507), .B2(n6079), .A(n4506), .ZN(U2902) );
  INV_X1 U5598 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4509) );
  AOI22_X1 U5599 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n6085), .B1(n6112), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4508) );
  OAI21_X1 U5600 ( .B1(n4509), .B2(n6079), .A(n4508), .ZN(U2901) );
  AOI22_X1 U5601 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n6085), .B1(n6112), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4510) );
  OAI21_X1 U5602 ( .B1(n4001), .B2(n6079), .A(n4510), .ZN(U2900) );
  INV_X1 U5603 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4512) );
  AOI22_X1 U5604 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n6085), .B1(n6112), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4511) );
  OAI21_X1 U5605 ( .B1(n4512), .B2(n6079), .A(n4511), .ZN(U2898) );
  INV_X1 U5606 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4514) );
  AOI22_X1 U5607 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n6085), .B1(n6112), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4513) );
  OAI21_X1 U5608 ( .B1(n4514), .B2(n6079), .A(n4513), .ZN(U2906) );
  INV_X1 U5609 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4516) );
  AOI22_X1 U5610 ( .A1(UWORD_REG_11__SCAN_IN), .A2(n6085), .B1(n6112), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4515) );
  OAI21_X1 U5611 ( .B1(n4516), .B2(n6079), .A(n4515), .ZN(U2896) );
  INV_X1 U5612 ( .A(EAX_REG_20__SCAN_IN), .ZN(n6704) );
  AOI22_X1 U5613 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6085), .B1(n6112), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4517) );
  OAI21_X1 U5614 ( .B1(n6704), .B2(n6079), .A(n4517), .ZN(U2903) );
  INV_X1 U5615 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6652) );
  AOI22_X1 U5616 ( .A1(UWORD_REG_13__SCAN_IN), .A2(n6085), .B1(n6112), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4518) );
  OAI21_X1 U5617 ( .B1(n6652), .B2(n6079), .A(n4518), .ZN(U2894) );
  XNOR2_X1 U5618 ( .A(n4520), .B(n4519), .ZN(n5332) );
  INV_X1 U5619 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4521) );
  AOI21_X1 U5620 ( .B1(n5576), .B2(n4522), .A(n4521), .ZN(n4523) );
  AOI211_X1 U5621 ( .C1(n4525), .C2(n3910), .A(n4524), .B(n4523), .ZN(n4526)
         );
  OAI21_X1 U5622 ( .B1(n5332), .B2(n6157), .A(n4526), .ZN(U2986) );
  INV_X1 U5623 ( .A(n5073), .ZN(n4527) );
  NAND2_X1 U5624 ( .A1(n4527), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6466) );
  INV_X1 U5625 ( .A(n6510), .ZN(n5926) );
  INV_X1 U5626 ( .A(n6502), .ZN(n5074) );
  INV_X1 U5627 ( .A(n6603), .ZN(n4528) );
  NOR2_X1 U5628 ( .A1(n4549), .A2(n4528), .ZN(n4529) );
  OAI22_X1 U5629 ( .A1(n5073), .A2(n6603), .B1(n4529), .B2(n4540), .ZN(n4530)
         );
  AOI21_X1 U5630 ( .B1(n4530), .B2(n6606), .A(n4564), .ZN(n4532) );
  MUX2_X1 U5631 ( .A(n4592), .B(n4532), .S(n4531), .Z(n4539) );
  INV_X1 U5632 ( .A(n4559), .ZN(n4536) );
  INV_X1 U5633 ( .A(n4533), .ZN(n4534) );
  OAI211_X1 U5634 ( .C1(n5927), .C2(n4536), .A(n4535), .B(n4534), .ZN(n4537)
         );
  INV_X1 U5635 ( .A(n4537), .ZN(n4538) );
  NAND2_X1 U5636 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4627), .ZN(n6586) );
  INV_X1 U5637 ( .A(n6586), .ZN(n6518) );
  AOI22_X1 U5638 ( .A1(n6469), .A2(n6511), .B1(FLUSH_REG_SCAN_IN), .B2(n6518), 
        .ZN(n5928) );
  OAI21_X1 U5639 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6588), .A(n5928), .ZN(
        n5930) );
  INV_X1 U5640 ( .A(n5930), .ZN(n5078) );
  AOI21_X1 U5641 ( .B1(n5074), .B2(n3861), .A(n5078), .ZN(n5077) );
  INV_X1 U5642 ( .A(n5077), .ZN(n4544) );
  NAND4_X1 U5643 ( .A1(n5927), .A2(n4540), .A3(n4561), .A4(n4084), .ZN(n4541)
         );
  OR2_X1 U5644 ( .A1(n4542), .A2(n4541), .ZN(n5067) );
  OAI22_X1 U5645 ( .A1(n6467), .A2(n5926), .B1(n6749), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4543) );
  OAI22_X1 U5646 ( .A1(n4544), .A2(n4543), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5930), .ZN(n4545) );
  OAI21_X1 U5647 ( .B1(n6466), .B2(n5926), .A(n4545), .ZN(U3461) );
  OAI222_X1 U5648 ( .A1(n5326), .A2(n5369), .B1(n5327), .B2(n6067), .C1(n5371), 
        .C2(n5332), .ZN(U2859) );
  XNOR2_X1 U5649 ( .A(n4547), .B(n4546), .ZN(n4579) );
  OR2_X1 U5650 ( .A1(n4548), .A2(n4549), .ZN(n4550) );
  AND2_X1 U5651 ( .A1(n4551), .A2(n4550), .ZN(n4572) );
  INV_X1 U5652 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6589) );
  OAI22_X1 U5653 ( .A1(n6250), .A2(n4572), .B1(n6589), .B2(n6248), .ZN(n4552)
         );
  INV_X1 U5654 ( .A(n4552), .ZN(n4557) );
  NAND2_X1 U5655 ( .A1(n6196), .A2(n4553), .ZN(n4555) );
  INV_X1 U5656 ( .A(n4730), .ZN(n4554) );
  MUX2_X1 U5657 ( .A(n4555), .B(n4554), .S(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .Z(n4556) );
  OAI211_X1 U5658 ( .C1(n4579), .C2(n6184), .A(n4557), .B(n4556), .ZN(U3017)
         );
  NAND2_X1 U5659 ( .A1(n6511), .A2(n4559), .ZN(n4562) );
  NAND4_X1 U5660 ( .A1(n5373), .A2(n3274), .A3(n6511), .A4(n3286), .ZN(n4560)
         );
  OAI22_X1 U5661 ( .A1(n5927), .A2(n4562), .B1(n4561), .B2(n4560), .ZN(n4563)
         );
  NAND2_X1 U5662 ( .A1(n3685), .A2(n4566), .ZN(n4567) );
  INV_X1 U5663 ( .A(n4567), .ZN(n4568) );
  INV_X1 U5664 ( .A(DATAI_0_), .ZN(n4683) );
  INV_X1 U5665 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6115) );
  OAI222_X1 U5666 ( .A1(n5424), .A2(n5332), .B1(n5417), .B2(n4683), .C1(n5416), 
        .C2(n6115), .ZN(U2891) );
  OAI21_X1 U5667 ( .B1(n4570), .B2(n4569), .A(n3154), .ZN(n5325) );
  INV_X1 U5668 ( .A(n5325), .ZN(n4577) );
  OAI22_X1 U5669 ( .A1(n5369), .A2(n4572), .B1(n4571), .B2(n6067), .ZN(n4573)
         );
  AOI21_X1 U5670 ( .B1(n4577), .B2(n4264), .A(n4573), .ZN(n4574) );
  INV_X1 U5671 ( .A(n4574), .ZN(U2858) );
  INV_X1 U5672 ( .A(DATAI_1_), .ZN(n6657) );
  INV_X1 U5673 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6109) );
  OAI222_X1 U5674 ( .A1(n5325), .A2(n5424), .B1(n5417), .B2(n6657), .C1(n5416), 
        .C2(n6109), .ZN(U2890) );
  INV_X1 U5675 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5320) );
  AOI22_X1 U5676 ( .A1(n5565), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6233), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4575) );
  OAI21_X1 U5677 ( .B1(n6182), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4575), 
        .ZN(n4576) );
  AOI21_X1 U5678 ( .B1(n4577), .B2(n6177), .A(n4576), .ZN(n4578) );
  OAI21_X1 U5679 ( .B1(n4579), .B2(n6159), .A(n4578), .ZN(U2985) );
  AND3_X1 U5680 ( .A1(n3154), .A2(n4581), .A3(n4580), .ZN(n4582) );
  NOR2_X1 U5681 ( .A1(n4744), .A2(n4582), .ZN(n6178) );
  INV_X1 U5682 ( .A(n6178), .ZN(n5318) );
  INV_X1 U5683 ( .A(DATAI_2_), .ZN(n4665) );
  INV_X1 U5684 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6107) );
  OAI222_X1 U5685 ( .A1(n5318), .A2(n5424), .B1(n5417), .B2(n4665), .C1(n5416), 
        .C2(n6107), .ZN(U2889) );
  NAND2_X1 U5686 ( .A1(n4744), .A2(n4583), .ZN(n4756) );
  OAI21_X1 U5687 ( .B1(n4744), .B2(n4583), .A(n4756), .ZN(n6052) );
  INV_X1 U5688 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4589) );
  INV_X1 U5689 ( .A(n4584), .ZN(n4586) );
  AOI21_X1 U5690 ( .B1(n4586), .B2(n5308), .A(n4585), .ZN(n4588) );
  OR2_X1 U5691 ( .A1(n4588), .A2(n4587), .ZN(n6249) );
  OAI222_X1 U5692 ( .A1(n6052), .A2(n5371), .B1(n4589), .B2(n6067), .C1(n6249), 
        .C2(n5369), .ZN(U2856) );
  INV_X1 U5693 ( .A(DATAI_3_), .ZN(n4670) );
  INV_X1 U5694 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6105) );
  OAI222_X1 U5695 ( .A1(n6052), .A2(n5424), .B1(n5417), .B2(n4670), .C1(n5416), 
        .C2(n6105), .ZN(U2888) );
  INV_X1 U5696 ( .A(n5067), .ZN(n4598) );
  NAND2_X1 U5697 ( .A1(n4592), .A2(n4591), .ZN(n4601) );
  XNOR2_X1 U5698 ( .A(n4593), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4596)
         );
  XNOR2_X1 U5699 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4594) );
  OAI22_X1 U5700 ( .A1(n5073), .A2(n4594), .B1(n4607), .B2(n4596), .ZN(n4595)
         );
  AOI21_X1 U5701 ( .B1(n4601), .B2(n4596), .A(n4595), .ZN(n4597) );
  OAI21_X1 U5702 ( .B1(n4590), .B2(n4598), .A(n4597), .ZN(n5063) );
  MUX2_X1 U5703 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n5063), .S(n6469), 
        .Z(n6473) );
  MUX2_X1 U5704 ( .A(n4600), .B(n4613), .S(n4593), .Z(n4602) );
  OAI21_X1 U5705 ( .B1(n4603), .B2(n4602), .A(n4601), .ZN(n4611) );
  NAND2_X1 U5706 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4604) );
  XNOR2_X1 U5707 ( .A(n4613), .B(n4604), .ZN(n4608) );
  NAND2_X1 U5708 ( .A1(n4593), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4605) );
  NAND2_X1 U5709 ( .A1(n4605), .A2(n4613), .ZN(n4606) );
  NAND2_X1 U5710 ( .A1(n3347), .A2(n4606), .ZN(n5764) );
  OAI22_X1 U5711 ( .A1(n5073), .A2(n4608), .B1(n4607), .B2(n5764), .ZN(n4609)
         );
  INV_X1 U5712 ( .A(n4609), .ZN(n4610) );
  NAND2_X1 U5713 ( .A1(n4611), .A2(n4610), .ZN(n4612) );
  AOI21_X1 U5714 ( .B1(n5866), .B2(n5067), .A(n4612), .ZN(n5765) );
  MUX2_X1 U5715 ( .A(n4613), .B(n5765), .S(n6469), .Z(n6475) );
  INV_X1 U5716 ( .A(n6475), .ZN(n4614) );
  NAND3_X1 U5717 ( .A1(n6473), .A2(n4614), .A3(n6749), .ZN(n4617) );
  NOR2_X1 U5718 ( .A1(n6749), .A2(FLUSH_REG_SCAN_IN), .ZN(n4624) );
  NAND2_X1 U5719 ( .A1(n4615), .A2(n4624), .ZN(n4616) );
  NAND2_X1 U5720 ( .A1(n4617), .A2(n4616), .ZN(n6488) );
  INV_X1 U5721 ( .A(n6488), .ZN(n4619) );
  NOR2_X1 U5722 ( .A1(n4619), .A2(n4618), .ZN(n4630) );
  INV_X1 U5723 ( .A(n4621), .ZN(n5778) );
  NOR2_X1 U5724 ( .A1(n4620), .A2(n5778), .ZN(n4622) );
  XNOR2_X1 U5725 ( .A(n4622), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6036)
         );
  OAI22_X1 U5726 ( .A1(n6036), .A2(n5927), .B1(n6469), .B2(n3884), .ZN(n4623)
         );
  NAND2_X1 U5727 ( .A1(n4623), .A2(n6749), .ZN(n4626) );
  NAND2_X1 U5728 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n4624), .ZN(n4625) );
  NAND2_X1 U5729 ( .A1(n4626), .A2(n4625), .ZN(n6486) );
  NOR3_X1 U5730 ( .A1(n4630), .A2(n6486), .A3(FLUSH_REG_SCAN_IN), .ZN(n4628)
         );
  NOR3_X1 U5731 ( .A1(n4630), .A2(n6486), .A3(n4629), .ZN(n6491) );
  NAND2_X1 U5732 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6588), .ZN(n4639) );
  INV_X1 U5733 ( .A(n4639), .ZN(n5761) );
  OAI22_X1 U5734 ( .A1(n6275), .A2(n6406), .B1(n6313), .B2(n5761), .ZN(n4631)
         );
  OAI21_X1 U5735 ( .B1(n6491), .B2(n4631), .A(n6274), .ZN(n4632) );
  OAI21_X1 U5736 ( .B1(n6274), .B2(n4937), .A(n4632), .ZN(U3465) );
  INV_X1 U5737 ( .A(n6274), .ZN(n4642) );
  INV_X1 U5738 ( .A(n4638), .ZN(n4634) );
  INV_X1 U5739 ( .A(n2964), .ZN(n4758) );
  INV_X1 U5740 ( .A(n4811), .ZN(n4636) );
  NAND2_X1 U5741 ( .A1(n4636), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4806) );
  AND2_X1 U5742 ( .A1(n2964), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6310) );
  NAND2_X1 U5743 ( .A1(n5822), .A2(n6310), .ZN(n6356) );
  NAND3_X1 U5744 ( .A1(n4806), .A2(n6403), .A3(n6356), .ZN(n6312) );
  AND2_X1 U5745 ( .A1(n6401), .A2(n6604), .ZN(n4842) );
  AOI222_X1 U5746 ( .A1(n6312), .A2(n6401), .B1(n5866), .B2(n4639), .C1(n4637), 
        .C2(n4842), .ZN(n4641) );
  NAND2_X1 U5747 ( .A1(n4642), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4640) );
  OAI21_X1 U5748 ( .B1(n4642), .B2(n4641), .A(n4640), .ZN(U3462) );
  NAND2_X1 U5749 ( .A1(n4643), .A2(n2964), .ZN(n4648) );
  INV_X1 U5750 ( .A(n4648), .ZN(n4644) );
  INV_X1 U5751 ( .A(n4842), .ZN(n6283) );
  OAI21_X1 U5752 ( .B1(n4644), .B2(n6157), .A(n6283), .ZN(n4646) );
  INV_X1 U5753 ( .A(n5865), .ZN(n5759) );
  INV_X1 U5754 ( .A(n4685), .ZN(n4645) );
  AOI21_X1 U5755 ( .B1(n4938), .B2(n6359), .A(n4645), .ZN(n4650) );
  NAND2_X1 U5756 ( .A1(n4646), .A2(n4650), .ZN(n4647) );
  INV_X1 U5757 ( .A(n6405), .ZN(n6361) );
  OAI211_X1 U5758 ( .C1(n6401), .C2(n4651), .A(n4647), .B(n6361), .ZN(n4688)
         );
  NAND2_X1 U5759 ( .A1(n6177), .A2(DATAI_29_), .ZN(n5849) );
  NAND2_X1 U5760 ( .A1(n6177), .A2(DATAI_21_), .ZN(n6446) );
  OAI22_X1 U5761 ( .A1(n5849), .A2(n4928), .B1(n4885), .B2(n6446), .ZN(n4654)
         );
  INV_X1 U5762 ( .A(n6441), .ZN(n5805) );
  INV_X1 U5763 ( .A(n4650), .ZN(n4652) );
  AOI22_X1 U5764 ( .A1(n4652), .A2(n6401), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4651), .ZN(n4684) );
  INV_X1 U5765 ( .A(DATAI_5_), .ZN(n4752) );
  OAI22_X1 U5766 ( .A1(n5805), .A2(n4685), .B1(n4684), .B2(n5898), .ZN(n4653)
         );
  AOI211_X1 U5767 ( .C1(INSTQUEUE_REG_15__5__SCAN_IN), .C2(n4688), .A(n4654), 
        .B(n4653), .ZN(n4655) );
  INV_X1 U5768 ( .A(n4655), .ZN(U3145) );
  NAND2_X1 U5769 ( .A1(n6177), .A2(DATAI_25_), .ZN(n6422) );
  NAND2_X1 U5770 ( .A1(n6177), .A2(DATAI_17_), .ZN(n6373) );
  OAI22_X1 U5771 ( .A1(n6422), .A2(n4928), .B1(n4885), .B2(n6373), .ZN(n4658)
         );
  INV_X1 U5772 ( .A(n6417), .ZN(n5788) );
  OAI22_X1 U5773 ( .A1(n5788), .A2(n4685), .B1(n4684), .B2(n5882), .ZN(n4657)
         );
  AOI211_X1 U5774 ( .C1(INSTQUEUE_REG_15__1__SCAN_IN), .C2(n4688), .A(n4658), 
        .B(n4657), .ZN(n4659) );
  INV_X1 U5775 ( .A(n4659), .ZN(U3141) );
  NAND2_X1 U5776 ( .A1(n6177), .A2(DATAI_30_), .ZN(n6389) );
  NAND2_X1 U5777 ( .A1(n6177), .A2(DATAI_22_), .ZN(n6454) );
  OAI22_X1 U5778 ( .A1(n6389), .A2(n4928), .B1(n4885), .B2(n6454), .ZN(n4663)
         );
  INV_X1 U5779 ( .A(n6447), .ZN(n5810) );
  OAI22_X1 U5780 ( .A1(n5810), .A2(n4685), .B1(n4684), .B2(n5902), .ZN(n4662)
         );
  AOI211_X1 U5781 ( .C1(INSTQUEUE_REG_15__6__SCAN_IN), .C2(n4688), .A(n4663), 
        .B(n4662), .ZN(n4664) );
  INV_X1 U5782 ( .A(n4664), .ZN(U3146) );
  NAND2_X1 U5783 ( .A1(n6177), .A2(DATAI_26_), .ZN(n6428) );
  NAND2_X1 U5784 ( .A1(n6177), .A2(DATAI_18_), .ZN(n6329) );
  OAI22_X1 U5785 ( .A1(n6428), .A2(n4928), .B1(n4885), .B2(n6329), .ZN(n4667)
         );
  INV_X1 U5786 ( .A(n6423), .ZN(n5792) );
  OAI22_X1 U5787 ( .A1(n5792), .A2(n4685), .B1(n4684), .B2(n5886), .ZN(n4666)
         );
  AOI211_X1 U5788 ( .C1(INSTQUEUE_REG_15__2__SCAN_IN), .C2(n4688), .A(n4667), 
        .B(n4666), .ZN(n4668) );
  INV_X1 U5789 ( .A(n4668), .ZN(U3142) );
  NAND2_X1 U5790 ( .A1(n6177), .A2(DATAI_27_), .ZN(n5842) );
  NAND2_X1 U5791 ( .A1(n6177), .A2(DATAI_19_), .ZN(n6434) );
  OAI22_X1 U5792 ( .A1(n5842), .A2(n4928), .B1(n4885), .B2(n6434), .ZN(n4672)
         );
  NOR2_X1 U5793 ( .A1(n4682), .A2(n4669), .ZN(n6429) );
  INV_X1 U5794 ( .A(n6429), .ZN(n5796) );
  OAI22_X1 U5795 ( .A1(n5796), .A2(n4685), .B1(n4684), .B2(n5890), .ZN(n4671)
         );
  AOI211_X1 U5796 ( .C1(INSTQUEUE_REG_15__3__SCAN_IN), .C2(n4688), .A(n4672), 
        .B(n4671), .ZN(n4673) );
  INV_X1 U5797 ( .A(n4673), .ZN(U3143) );
  NAND2_X1 U5798 ( .A1(n6177), .A2(DATAI_31_), .ZN(n6465) );
  NAND2_X1 U5799 ( .A1(n6177), .A2(DATAI_23_), .ZN(n6308) );
  OAI22_X1 U5800 ( .A1(n6465), .A2(n4928), .B1(n4885), .B2(n6308), .ZN(n4676)
         );
  INV_X1 U5801 ( .A(n6456), .ZN(n5817) );
  OAI22_X1 U5802 ( .A1(n5817), .A2(n4685), .B1(n4684), .B2(n5909), .ZN(n4675)
         );
  AOI211_X1 U5803 ( .C1(INSTQUEUE_REG_15__7__SCAN_IN), .C2(n4688), .A(n4676), 
        .B(n4675), .ZN(n4677) );
  INV_X1 U5804 ( .A(n4677), .ZN(U3147) );
  NAND2_X1 U5805 ( .A1(n6177), .A2(DATAI_28_), .ZN(n6440) );
  NAND2_X1 U5806 ( .A1(n6177), .A2(DATAI_20_), .ZN(n6381) );
  OAI22_X1 U5807 ( .A1(n6440), .A2(n4928), .B1(n4885), .B2(n6381), .ZN(n4679)
         );
  INV_X1 U5808 ( .A(n6435), .ZN(n5801) );
  INV_X1 U5809 ( .A(DATAI_4_), .ZN(n4757) );
  OAI22_X1 U5810 ( .A1(n5801), .A2(n4685), .B1(n4684), .B2(n5894), .ZN(n4678)
         );
  AOI211_X1 U5811 ( .C1(INSTQUEUE_REG_15__4__SCAN_IN), .C2(n4688), .A(n4679), 
        .B(n4678), .ZN(n4680) );
  INV_X1 U5812 ( .A(n4680), .ZN(U3144) );
  NAND2_X1 U5813 ( .A1(n6177), .A2(DATAI_24_), .ZN(n6416) );
  NAND2_X1 U5814 ( .A1(n6177), .A2(DATAI_16_), .ZN(n6369) );
  OAI22_X1 U5815 ( .A1(n6416), .A2(n4928), .B1(n4885), .B2(n6369), .ZN(n4687)
         );
  NOR2_X2 U5816 ( .A1(n4682), .A2(n4681), .ZN(n6399) );
  INV_X1 U5817 ( .A(n6399), .ZN(n5784) );
  INV_X1 U5818 ( .A(n6413), .ZN(n5878) );
  OAI22_X1 U5819 ( .A1(n5784), .A2(n4685), .B1(n4684), .B2(n5878), .ZN(n4686)
         );
  AOI211_X1 U5820 ( .C1(INSTQUEUE_REG_15__0__SCAN_IN), .C2(n4688), .A(n4687), 
        .B(n4686), .ZN(n4689) );
  INV_X1 U5821 ( .A(n4689), .ZN(U3140) );
  NOR3_X1 U5822 ( .A1(n4694), .A2(n2964), .A3(n6604), .ZN(n4690) );
  NOR2_X1 U5823 ( .A1(n4690), .A2(n6406), .ZN(n4697) );
  INV_X1 U5824 ( .A(n4590), .ZN(n4691) );
  NAND2_X1 U5825 ( .A1(n4691), .A2(n5759), .ZN(n5773) );
  OR2_X1 U5826 ( .A1(n5773), .A2(n6357), .ZN(n4692) );
  NAND3_X1 U5827 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6397), .A3(n4936), .ZN(n5769) );
  OR2_X1 U5828 ( .A1(n4937), .A2(n5769), .ZN(n4721) );
  NAND2_X1 U5829 ( .A1(n4692), .A2(n4721), .ZN(n4699) );
  INV_X1 U5830 ( .A(n5769), .ZN(n4693) );
  INV_X1 U5831 ( .A(n6373), .ZN(n6418) );
  NOR2_X1 U5832 ( .A1(n4694), .A2(n2964), .ZN(n4695) );
  NAND2_X1 U5833 ( .A1(n4695), .A2(n5767), .ZN(n4994) );
  NAND2_X1 U5834 ( .A1(n4695), .A2(n6275), .ZN(n5775) );
  OAI22_X1 U5835 ( .A1(n5788), .A2(n4721), .B1(n5775), .B2(n6422), .ZN(n4696)
         );
  AOI21_X1 U5836 ( .B1(n6418), .B2(n6350), .A(n4696), .ZN(n4702) );
  INV_X1 U5837 ( .A(n4697), .ZN(n4700) );
  AOI21_X1 U5838 ( .B1(n6406), .B2(n5769), .A(n6405), .ZN(n4698) );
  NAND2_X1 U5839 ( .A1(n4723), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4701) );
  OAI211_X1 U5840 ( .C1(n4726), .C2(n5882), .A(n4702), .B(n4701), .ZN(U3061)
         );
  INV_X1 U5841 ( .A(n6381), .ZN(n6436) );
  OAI22_X1 U5842 ( .A1(n5801), .A2(n4721), .B1(n5775), .B2(n6440), .ZN(n4703)
         );
  AOI21_X1 U5843 ( .B1(n6436), .B2(n6350), .A(n4703), .ZN(n4705) );
  NAND2_X1 U5844 ( .A1(n4723), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4704) );
  OAI211_X1 U5845 ( .C1(n4726), .C2(n5894), .A(n4705), .B(n4704), .ZN(U3064)
         );
  INV_X1 U5846 ( .A(n6329), .ZN(n6424) );
  OAI22_X1 U5847 ( .A1(n5792), .A2(n4721), .B1(n5775), .B2(n6428), .ZN(n4706)
         );
  AOI21_X1 U5848 ( .B1(n6424), .B2(n6350), .A(n4706), .ZN(n4708) );
  NAND2_X1 U5849 ( .A1(n4723), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4707) );
  OAI211_X1 U5850 ( .C1(n4726), .C2(n5886), .A(n4708), .B(n4707), .ZN(U3062)
         );
  INV_X1 U5851 ( .A(n6454), .ZN(n6386) );
  OAI22_X1 U5852 ( .A1(n5810), .A2(n4721), .B1(n5775), .B2(n6389), .ZN(n4709)
         );
  AOI21_X1 U5853 ( .B1(n6386), .B2(n6350), .A(n4709), .ZN(n4711) );
  NAND2_X1 U5854 ( .A1(n4723), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4710) );
  OAI211_X1 U5855 ( .C1(n4726), .C2(n5902), .A(n4711), .B(n4710), .ZN(U3066)
         );
  INV_X1 U5856 ( .A(n6434), .ZN(n5798) );
  OAI22_X1 U5857 ( .A1(n5796), .A2(n4721), .B1(n5775), .B2(n5842), .ZN(n4712)
         );
  AOI21_X1 U5858 ( .B1(n5798), .B2(n6350), .A(n4712), .ZN(n4714) );
  NAND2_X1 U5859 ( .A1(n4723), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4713) );
  OAI211_X1 U5860 ( .C1(n4726), .C2(n5890), .A(n4714), .B(n4713), .ZN(U3063)
         );
  INV_X1 U5861 ( .A(n6446), .ZN(n5807) );
  OAI22_X1 U5862 ( .A1(n5805), .A2(n4721), .B1(n5775), .B2(n5849), .ZN(n4715)
         );
  AOI21_X1 U5863 ( .B1(n5807), .B2(n6350), .A(n4715), .ZN(n4717) );
  NAND2_X1 U5864 ( .A1(n4723), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4716) );
  OAI211_X1 U5865 ( .C1(n4726), .C2(n5898), .A(n4717), .B(n4716), .ZN(U3065)
         );
  OAI22_X1 U5866 ( .A1(n5784), .A2(n4721), .B1(n5775), .B2(n6416), .ZN(n4718)
         );
  AOI21_X1 U5867 ( .B1(n6400), .B2(n6350), .A(n4718), .ZN(n4720) );
  NAND2_X1 U5868 ( .A1(n4723), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4719) );
  OAI211_X1 U5869 ( .C1(n4726), .C2(n5878), .A(n4720), .B(n4719), .ZN(U3060)
         );
  OAI22_X1 U5870 ( .A1(n5817), .A2(n4721), .B1(n5775), .B2(n6465), .ZN(n4722)
         );
  AOI21_X1 U5871 ( .B1(n6457), .B2(n6350), .A(n4722), .ZN(n4725) );
  NAND2_X1 U5872 ( .A1(n4723), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4724) );
  OAI211_X1 U5873 ( .C1(n4726), .C2(n5909), .A(n4725), .B(n4724), .ZN(U3067)
         );
  OAI21_X1 U5874 ( .B1(n4729), .B2(n4727), .A(n4728), .ZN(n4837) );
  NOR2_X1 U5875 ( .A1(n4734), .A2(n4733), .ZN(n6229) );
  INV_X1 U5876 ( .A(n6229), .ZN(n4732) );
  AOI22_X1 U5877 ( .A1(n6259), .A2(n6193), .B1(n6200), .B2(n4730), .ZN(n4731)
         );
  INV_X1 U5878 ( .A(n4731), .ZN(n6267) );
  AOI21_X1 U5879 ( .B1(n6196), .B2(n4732), .A(n6267), .ZN(n6235) );
  AOI221_X1 U5880 ( .B1(n6200), .B2(n4734), .C1(n4733), .C2(n4734), .A(n6235), 
        .ZN(n4735) );
  INV_X1 U5881 ( .A(n4735), .ZN(n4743) );
  NAND2_X1 U5882 ( .A1(n4737), .A2(n4738), .ZN(n4739) );
  AND2_X1 U5883 ( .A1(n4736), .A2(n4739), .ZN(n5301) );
  AND2_X1 U5884 ( .A1(n6233), .A2(REIP_REG_5__SCAN_IN), .ZN(n4831) );
  NOR3_X1 U5885 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4740), .A3(n6268), 
        .ZN(n4741) );
  AOI211_X1 U5886 ( .C1(n6262), .C2(n5301), .A(n4831), .B(n4741), .ZN(n4742)
         );
  OAI211_X1 U5887 ( .C1(n6184), .C2(n4837), .A(n4743), .B(n4742), .ZN(U3013)
         );
  AND2_X1 U5888 ( .A1(n4745), .A2(n4744), .ZN(n4749) );
  OAI21_X1 U5889 ( .B1(n4749), .B2(n4748), .A(n4747), .ZN(n5304) );
  INV_X1 U5890 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4751) );
  INV_X1 U5891 ( .A(n5301), .ZN(n4750) );
  OAI222_X1 U5892 ( .A1(n5304), .A2(n5371), .B1(n6067), .B2(n4751), .C1(n4750), 
        .C2(n5369), .ZN(U2854) );
  INV_X1 U5893 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6101) );
  OAI222_X1 U5894 ( .A1(n5304), .A2(n5424), .B1(n5417), .B2(n4752), .C1(n5416), 
        .C2(n6101), .ZN(U2886) );
  XNOR2_X1 U5895 ( .A(n4747), .B(n4753), .ZN(n6158) );
  OAI222_X1 U5896 ( .A1(n5417), .A2(n4661), .B1(n5424), .B2(n6158), .C1(n4754), 
        .C2(n5416), .ZN(U2885) );
  XOR2_X1 U5897 ( .A(n4755), .B(n4756), .Z(n6169) );
  INV_X1 U5898 ( .A(n6169), .ZN(n6037) );
  INV_X1 U5899 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6103) );
  OAI222_X1 U5900 ( .A1(n5424), .A2(n6037), .B1(n5417), .B2(n4757), .C1(n5416), 
        .C2(n6103), .ZN(U2887) );
  NAND3_X1 U5901 ( .A1(n6397), .A2(n6474), .A3(n4936), .ZN(n4843) );
  INV_X1 U5902 ( .A(n4843), .ZN(n4764) );
  NAND2_X1 U5903 ( .A1(n4633), .A2(n4758), .ZN(n4759) );
  OR2_X1 U5904 ( .A1(n4637), .A2(n4759), .ZN(n4768) );
  INV_X1 U5905 ( .A(n4847), .ZN(n4762) );
  NOR2_X1 U5906 ( .A1(n4937), .A2(n4843), .ZN(n4797) );
  INV_X1 U5907 ( .A(n4797), .ZN(n4760) );
  AND2_X1 U5908 ( .A1(n4761), .A2(n4760), .ZN(n4766) );
  AOI21_X1 U5909 ( .B1(n4762), .B2(n4766), .A(n6405), .ZN(n4763) );
  OAI21_X1 U5910 ( .B1(n6401), .B2(n4764), .A(n4763), .ZN(n4765) );
  INV_X1 U5911 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4772) );
  OAI22_X1 U5912 ( .A1(n4847), .A2(n4766), .B1(n4843), .B2(n6409), .ZN(n4800)
         );
  NAND2_X1 U5913 ( .A1(n4767), .A2(n6275), .ZN(n4848) );
  AOI22_X1 U5914 ( .A1(n6303), .A2(n5798), .B1(n6429), .B2(n4797), .ZN(n4769)
         );
  OAI21_X1 U5915 ( .B1(n5842), .B2(n4848), .A(n4769), .ZN(n4770) );
  AOI21_X1 U5916 ( .B1(n6431), .B2(n4800), .A(n4770), .ZN(n4771) );
  OAI21_X1 U5917 ( .B1(n4803), .B2(n4772), .A(n4771), .ZN(U3031) );
  INV_X1 U5918 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4776) );
  AOI22_X1 U5919 ( .A1(n6303), .A2(n6400), .B1(n6399), .B2(n4797), .ZN(n4773)
         );
  OAI21_X1 U5920 ( .B1(n6416), .B2(n4848), .A(n4773), .ZN(n4774) );
  AOI21_X1 U5921 ( .B1(n6413), .B2(n4800), .A(n4774), .ZN(n4775) );
  OAI21_X1 U5922 ( .B1(n4803), .B2(n4776), .A(n4775), .ZN(U3028) );
  INV_X1 U5923 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4780) );
  AOI22_X1 U5924 ( .A1(n6303), .A2(n6424), .B1(n6423), .B2(n4797), .ZN(n4777)
         );
  OAI21_X1 U5925 ( .B1(n6428), .B2(n4848), .A(n4777), .ZN(n4778) );
  AOI21_X1 U5926 ( .B1(n6425), .B2(n4800), .A(n4778), .ZN(n4779) );
  OAI21_X1 U5927 ( .B1(n4803), .B2(n4780), .A(n4779), .ZN(U3030) );
  INV_X1 U5928 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4784) );
  AOI22_X1 U5929 ( .A1(n6303), .A2(n6457), .B1(n6456), .B2(n4797), .ZN(n4781)
         );
  OAI21_X1 U5930 ( .B1(n6465), .B2(n4848), .A(n4781), .ZN(n4782) );
  AOI21_X1 U5931 ( .B1(n6460), .B2(n4800), .A(n4782), .ZN(n4783) );
  OAI21_X1 U5932 ( .B1(n4803), .B2(n4784), .A(n4783), .ZN(U3035) );
  INV_X1 U5933 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4788) );
  AOI22_X1 U5934 ( .A1(n6303), .A2(n6386), .B1(n6447), .B2(n4797), .ZN(n4785)
         );
  OAI21_X1 U5935 ( .B1(n6389), .B2(n4848), .A(n4785), .ZN(n4786) );
  AOI21_X1 U5936 ( .B1(n6450), .B2(n4800), .A(n4786), .ZN(n4787) );
  OAI21_X1 U5937 ( .B1(n4803), .B2(n4788), .A(n4787), .ZN(U3034) );
  INV_X1 U5938 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4792) );
  AOI22_X1 U5939 ( .A1(n6303), .A2(n5807), .B1(n6441), .B2(n4797), .ZN(n4789)
         );
  OAI21_X1 U5940 ( .B1(n5849), .B2(n4848), .A(n4789), .ZN(n4790) );
  AOI21_X1 U5941 ( .B1(n6443), .B2(n4800), .A(n4790), .ZN(n4791) );
  OAI21_X1 U5942 ( .B1(n4803), .B2(n4792), .A(n4791), .ZN(U3033) );
  INV_X1 U5943 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4796) );
  AOI22_X1 U5944 ( .A1(n6303), .A2(n6418), .B1(n6417), .B2(n4797), .ZN(n4793)
         );
  OAI21_X1 U5945 ( .B1(n6422), .B2(n4848), .A(n4793), .ZN(n4794) );
  AOI21_X1 U5946 ( .B1(n6419), .B2(n4800), .A(n4794), .ZN(n4795) );
  OAI21_X1 U5947 ( .B1(n4803), .B2(n4796), .A(n4795), .ZN(U3029) );
  INV_X1 U5948 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4802) );
  AOI22_X1 U5949 ( .A1(n6303), .A2(n6436), .B1(n6435), .B2(n4797), .ZN(n4798)
         );
  OAI21_X1 U5950 ( .B1(n6440), .B2(n4848), .A(n4798), .ZN(n4799) );
  AOI21_X1 U5951 ( .B1(n6437), .B2(n4800), .A(n4799), .ZN(n4801) );
  OAI21_X1 U5952 ( .B1(n4803), .B2(n4802), .A(n4801), .ZN(U3032) );
  OR2_X1 U5953 ( .A1(n4587), .A2(n4804), .ZN(n4805) );
  NAND2_X1 U5954 ( .A1(n4737), .A2(n4805), .ZN(n6241) );
  INV_X1 U5955 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6028) );
  OAI222_X1 U5956 ( .A1(n6241), .A2(n5369), .B1(n6067), .B2(n6028), .C1(n5371), 
        .C2(n6037), .ZN(U2855) );
  NAND2_X1 U5957 ( .A1(n6401), .A2(n4806), .ZN(n4809) );
  INV_X1 U5958 ( .A(n5773), .ZN(n5777) );
  NAND3_X1 U5959 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n4936), .ZN(n5011) );
  NOR2_X1 U5960 ( .A1(n4937), .A2(n5011), .ZN(n4828) );
  AOI21_X1 U5961 ( .B1(n5777), .B2(n4938), .A(n4828), .ZN(n4810) );
  INV_X1 U5962 ( .A(n4810), .ZN(n4808) );
  AOI21_X1 U5963 ( .B1(n6406), .B2(n5011), .A(n6405), .ZN(n4807) );
  AOI22_X1 U5964 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4827), .B1(n6437), 
        .B2(n4826), .ZN(n4813) );
  INV_X1 U5965 ( .A(n6440), .ZN(n6378) );
  AOI22_X1 U5966 ( .A1(n5040), .A2(n6378), .B1(n6435), .B2(n4828), .ZN(n4812)
         );
  OAI211_X1 U5967 ( .C1(n6381), .C2(n4927), .A(n4813), .B(n4812), .ZN(U3128)
         );
  AOI22_X1 U5968 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4827), .B1(n6443), 
        .B2(n4826), .ZN(n4815) );
  INV_X1 U5969 ( .A(n5849), .ZN(n6442) );
  AOI22_X1 U5970 ( .A1(n5040), .A2(n6442), .B1(n6441), .B2(n4828), .ZN(n4814)
         );
  OAI211_X1 U5971 ( .C1(n6446), .C2(n4927), .A(n4815), .B(n4814), .ZN(U3129)
         );
  AOI22_X1 U5972 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4827), .B1(n6413), 
        .B2(n4826), .ZN(n4817) );
  INV_X1 U5973 ( .A(n6416), .ZN(n6355) );
  AOI22_X1 U5974 ( .A1(n5040), .A2(n6355), .B1(n6399), .B2(n4828), .ZN(n4816)
         );
  OAI211_X1 U5975 ( .C1(n6369), .C2(n4927), .A(n4817), .B(n4816), .ZN(U3124)
         );
  AOI22_X1 U5976 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4827), .B1(n6425), 
        .B2(n4826), .ZN(n4819) );
  INV_X1 U5977 ( .A(n6428), .ZN(n6326) );
  AOI22_X1 U5978 ( .A1(n5040), .A2(n6326), .B1(n6423), .B2(n4828), .ZN(n4818)
         );
  OAI211_X1 U5979 ( .C1(n6329), .C2(n4927), .A(n4819), .B(n4818), .ZN(U3126)
         );
  AOI22_X1 U5980 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4827), .B1(n6419), 
        .B2(n4826), .ZN(n4821) );
  INV_X1 U5981 ( .A(n6422), .ZN(n6370) );
  AOI22_X1 U5982 ( .A1(n5040), .A2(n6370), .B1(n6417), .B2(n4828), .ZN(n4820)
         );
  OAI211_X1 U5983 ( .C1(n6373), .C2(n4927), .A(n4821), .B(n4820), .ZN(U3125)
         );
  AOI22_X1 U5984 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4827), .B1(n6460), 
        .B2(n4826), .ZN(n4823) );
  INV_X1 U5985 ( .A(n6465), .ZN(n6304) );
  AOI22_X1 U5986 ( .A1(n5040), .A2(n6304), .B1(n6456), .B2(n4828), .ZN(n4822)
         );
  OAI211_X1 U5987 ( .C1(n6308), .C2(n4927), .A(n4823), .B(n4822), .ZN(U3131)
         );
  AOI22_X1 U5988 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4827), .B1(n6450), 
        .B2(n4826), .ZN(n4825) );
  INV_X1 U5989 ( .A(n6389), .ZN(n6448) );
  AOI22_X1 U5990 ( .A1(n5040), .A2(n6448), .B1(n6447), .B2(n4828), .ZN(n4824)
         );
  OAI211_X1 U5991 ( .C1(n6454), .C2(n4927), .A(n4825), .B(n4824), .ZN(U3130)
         );
  AOI22_X1 U5992 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4827), .B1(n6431), 
        .B2(n4826), .ZN(n4830) );
  INV_X1 U5993 ( .A(n5842), .ZN(n6430) );
  AOI22_X1 U5994 ( .A1(n5040), .A2(n6430), .B1(n6429), .B2(n4828), .ZN(n4829)
         );
  OAI211_X1 U5995 ( .C1(n6434), .C2(n4927), .A(n4830), .B(n4829), .ZN(U3127)
         );
  INV_X1 U5996 ( .A(n5304), .ZN(n4835) );
  INV_X1 U5997 ( .A(n5300), .ZN(n4833) );
  AOI21_X1 U5998 ( .B1(n5565), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4831), 
        .ZN(n4832) );
  OAI21_X1 U5999 ( .B1(n6182), .B2(n4833), .A(n4832), .ZN(n4834) );
  AOI21_X1 U6000 ( .B1(n4835), .B2(n6177), .A(n4834), .ZN(n4836) );
  OAI21_X1 U6001 ( .B1(n6159), .B2(n4837), .A(n4836), .ZN(U2981) );
  INV_X1 U6002 ( .A(n6158), .ZN(n6026) );
  NAND2_X1 U6003 ( .A1(n4736), .A2(n4838), .ZN(n4839) );
  AND2_X1 U6004 ( .A1(n5002), .A2(n4839), .ZN(n6232) );
  INV_X1 U6005 ( .A(n6232), .ZN(n6018) );
  OAI22_X1 U6006 ( .A1(n5369), .A2(n6018), .B1(n6023), .B2(n6067), .ZN(n4840)
         );
  AOI21_X1 U6007 ( .B1(n6026), .B2(n4264), .A(n4840), .ZN(n4841) );
  INV_X1 U6008 ( .A(n4841), .ZN(U2853) );
  INV_X1 U6009 ( .A(n5831), .ZN(n5823) );
  OAI22_X1 U6010 ( .A1(n4885), .A2(n4842), .B1(n5866), .B2(n5823), .ZN(n4846)
         );
  NOR2_X1 U6011 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4843), .ZN(n4882)
         );
  INV_X1 U6012 ( .A(n4882), .ZN(n4844) );
  NOR2_X1 U6013 ( .A1(n4849), .A2(n6409), .ZN(n5869) );
  INV_X1 U6014 ( .A(n5008), .ZN(n4892) );
  NOR2_X1 U6015 ( .A1(n4892), .A2(n5009), .ZN(n5770) );
  OAI21_X1 U6016 ( .B1(n5770), .B2(n5874), .A(n4891), .ZN(n5779) );
  AOI211_X1 U6017 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4844), .A(n5869), .B(
        n5779), .ZN(n4845) );
  NAND2_X1 U6018 ( .A1(n4880), .A2(n5807), .ZN(n4853) );
  OR2_X1 U6019 ( .A1(n5866), .A2(n6406), .ZN(n5774) );
  INV_X1 U6020 ( .A(n5774), .ZN(n4973) );
  NAND2_X1 U6021 ( .A1(n4973), .A2(n5831), .ZN(n4851) );
  NAND2_X1 U6022 ( .A1(n5770), .A2(n6279), .ZN(n4850) );
  NAND2_X1 U6023 ( .A1(n4851), .A2(n4850), .ZN(n4881) );
  AOI22_X1 U6024 ( .A1(n6441), .A2(n4882), .B1(n6443), .B2(n4881), .ZN(n4852)
         );
  OAI211_X1 U6025 ( .C1(n4885), .C2(n5849), .A(n4853), .B(n4852), .ZN(n4854)
         );
  AOI21_X1 U6026 ( .B1(n4887), .B2(INSTQUEUE_REG_0__5__SCAN_IN), .A(n4854), 
        .ZN(n4855) );
  INV_X1 U6027 ( .A(n4855), .ZN(U3025) );
  NAND2_X1 U6028 ( .A1(n4880), .A2(n6418), .ZN(n4857) );
  AOI22_X1 U6029 ( .A1(n6417), .A2(n4882), .B1(n6419), .B2(n4881), .ZN(n4856)
         );
  OAI211_X1 U6030 ( .C1(n4885), .C2(n6422), .A(n4857), .B(n4856), .ZN(n4858)
         );
  AOI21_X1 U6031 ( .B1(n4887), .B2(INSTQUEUE_REG_0__1__SCAN_IN), .A(n4858), 
        .ZN(n4859) );
  INV_X1 U6032 ( .A(n4859), .ZN(U3021) );
  NAND2_X1 U6033 ( .A1(n4880), .A2(n6457), .ZN(n4861) );
  AOI22_X1 U6034 ( .A1(n6456), .A2(n4882), .B1(n6460), .B2(n4881), .ZN(n4860)
         );
  OAI211_X1 U6035 ( .C1(n4885), .C2(n6465), .A(n4861), .B(n4860), .ZN(n4862)
         );
  AOI21_X1 U6036 ( .B1(n4887), .B2(INSTQUEUE_REG_0__7__SCAN_IN), .A(n4862), 
        .ZN(n4863) );
  INV_X1 U6037 ( .A(n4863), .ZN(U3027) );
  NAND2_X1 U6038 ( .A1(n4880), .A2(n6424), .ZN(n4865) );
  AOI22_X1 U6039 ( .A1(n6423), .A2(n4882), .B1(n6425), .B2(n4881), .ZN(n4864)
         );
  OAI211_X1 U6040 ( .C1(n4885), .C2(n6428), .A(n4865), .B(n4864), .ZN(n4866)
         );
  AOI21_X1 U6041 ( .B1(n4887), .B2(INSTQUEUE_REG_0__2__SCAN_IN), .A(n4866), 
        .ZN(n4867) );
  INV_X1 U6042 ( .A(n4867), .ZN(U3022) );
  NAND2_X1 U6043 ( .A1(n4880), .A2(n5798), .ZN(n4869) );
  AOI22_X1 U6044 ( .A1(n6429), .A2(n4882), .B1(n6431), .B2(n4881), .ZN(n4868)
         );
  OAI211_X1 U6045 ( .C1(n4885), .C2(n5842), .A(n4869), .B(n4868), .ZN(n4870)
         );
  AOI21_X1 U6046 ( .B1(n4887), .B2(INSTQUEUE_REG_0__3__SCAN_IN), .A(n4870), 
        .ZN(n4871) );
  INV_X1 U6047 ( .A(n4871), .ZN(U3023) );
  NAND2_X1 U6048 ( .A1(n4880), .A2(n6386), .ZN(n4873) );
  AOI22_X1 U6049 ( .A1(n6447), .A2(n4882), .B1(n6450), .B2(n4881), .ZN(n4872)
         );
  OAI211_X1 U6050 ( .C1(n4885), .C2(n6389), .A(n4873), .B(n4872), .ZN(n4874)
         );
  AOI21_X1 U6051 ( .B1(n4887), .B2(INSTQUEUE_REG_0__6__SCAN_IN), .A(n4874), 
        .ZN(n4875) );
  INV_X1 U6052 ( .A(n4875), .ZN(U3026) );
  NAND2_X1 U6053 ( .A1(n4880), .A2(n6436), .ZN(n4877) );
  AOI22_X1 U6054 ( .A1(n6435), .A2(n4882), .B1(n6437), .B2(n4881), .ZN(n4876)
         );
  OAI211_X1 U6055 ( .C1(n4885), .C2(n6440), .A(n4877), .B(n4876), .ZN(n4878)
         );
  AOI21_X1 U6056 ( .B1(n4887), .B2(INSTQUEUE_REG_0__4__SCAN_IN), .A(n4878), 
        .ZN(n4879) );
  INV_X1 U6057 ( .A(n4879), .ZN(U3024) );
  NAND2_X1 U6058 ( .A1(n4880), .A2(n6400), .ZN(n4884) );
  AOI22_X1 U6059 ( .A1(n6399), .A2(n4882), .B1(n6413), .B2(n4881), .ZN(n4883)
         );
  OAI211_X1 U6060 ( .C1(n4885), .C2(n6416), .A(n4884), .B(n4883), .ZN(n4886)
         );
  AOI21_X1 U6061 ( .B1(n4887), .B2(INSTQUEUE_REG_0__0__SCAN_IN), .A(n4886), 
        .ZN(n4888) );
  INV_X1 U6062 ( .A(n4888), .ZN(U3020) );
  AOI21_X1 U6063 ( .B1(n4927), .B2(n4928), .A(n6604), .ZN(n4889) );
  NOR3_X1 U6064 ( .A1(n4889), .A2(n6359), .A3(n6406), .ZN(n4895) );
  NOR2_X1 U6065 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4890), .ZN(n4926)
         );
  OAI21_X1 U6066 ( .B1(n4892), .B2(n6409), .A(n4891), .ZN(n5868) );
  NOR3_X1 U6067 ( .A1(n5868), .A2(n6397), .A3(n6279), .ZN(n4893) );
  OAI21_X1 U6068 ( .B1(n6588), .B2(n4926), .A(n4893), .ZN(n4894) );
  INV_X1 U6069 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4899) );
  NOR2_X1 U6070 ( .A1(n6278), .A2(n6406), .ZN(n5832) );
  NOR2_X1 U6071 ( .A1(n5008), .A2(n6397), .ZN(n5867) );
  AOI22_X1 U6072 ( .A1(n5832), .A2(n6359), .B1(n5867), .B2(n5869), .ZN(n4924)
         );
  NOR2_X1 U6073 ( .A1(n4924), .A2(n5890), .ZN(n4897) );
  OAI22_X1 U6074 ( .A1(n5842), .A2(n4927), .B1(n4928), .B2(n6434), .ZN(n4896)
         );
  AOI211_X1 U6075 ( .C1(n4926), .C2(n6429), .A(n4897), .B(n4896), .ZN(n4898)
         );
  OAI21_X1 U6076 ( .B1(n4934), .B2(n4899), .A(n4898), .ZN(U3135) );
  INV_X1 U6077 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4903) );
  NOR2_X1 U6078 ( .A1(n4924), .A2(n5902), .ZN(n4901) );
  OAI22_X1 U6079 ( .A1(n6389), .A2(n4927), .B1(n4928), .B2(n6454), .ZN(n4900)
         );
  AOI211_X1 U6080 ( .C1(n4926), .C2(n6447), .A(n4901), .B(n4900), .ZN(n4902)
         );
  OAI21_X1 U6081 ( .B1(n4934), .B2(n4903), .A(n4902), .ZN(U3138) );
  INV_X1 U6082 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4907) );
  NOR2_X1 U6083 ( .A1(n4924), .A2(n5909), .ZN(n4905) );
  OAI22_X1 U6084 ( .A1(n6465), .A2(n4927), .B1(n4928), .B2(n6308), .ZN(n4904)
         );
  AOI211_X1 U6085 ( .C1(n4926), .C2(n6456), .A(n4905), .B(n4904), .ZN(n4906)
         );
  OAI21_X1 U6086 ( .B1(n4934), .B2(n4907), .A(n4906), .ZN(U3139) );
  INV_X1 U6087 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4911) );
  NOR2_X1 U6088 ( .A1(n4924), .A2(n5882), .ZN(n4909) );
  OAI22_X1 U6089 ( .A1(n6422), .A2(n4927), .B1(n4928), .B2(n6373), .ZN(n4908)
         );
  AOI211_X1 U6090 ( .C1(n4926), .C2(n6417), .A(n4909), .B(n4908), .ZN(n4910)
         );
  OAI21_X1 U6091 ( .B1(n4934), .B2(n4911), .A(n4910), .ZN(U3133) );
  INV_X1 U6092 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4915) );
  NOR2_X1 U6093 ( .A1(n4924), .A2(n5898), .ZN(n4913) );
  OAI22_X1 U6094 ( .A1(n5849), .A2(n4927), .B1(n4928), .B2(n6446), .ZN(n4912)
         );
  AOI211_X1 U6095 ( .C1(n4926), .C2(n6441), .A(n4913), .B(n4912), .ZN(n4914)
         );
  OAI21_X1 U6096 ( .B1(n4934), .B2(n4915), .A(n4914), .ZN(U3137) );
  INV_X1 U6097 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4919) );
  NOR2_X1 U6098 ( .A1(n4924), .A2(n5894), .ZN(n4917) );
  OAI22_X1 U6099 ( .A1(n6440), .A2(n4927), .B1(n4928), .B2(n6381), .ZN(n4916)
         );
  AOI211_X1 U6100 ( .C1(n4926), .C2(n6435), .A(n4917), .B(n4916), .ZN(n4918)
         );
  OAI21_X1 U6101 ( .B1(n4934), .B2(n4919), .A(n4918), .ZN(U3136) );
  INV_X1 U6102 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4923) );
  NOR2_X1 U6103 ( .A1(n4924), .A2(n5886), .ZN(n4921) );
  OAI22_X1 U6104 ( .A1(n6428), .A2(n4927), .B1(n4928), .B2(n6329), .ZN(n4920)
         );
  AOI211_X1 U6105 ( .C1(n4926), .C2(n6423), .A(n4921), .B(n4920), .ZN(n4922)
         );
  OAI21_X1 U6106 ( .B1(n4934), .B2(n4923), .A(n4922), .ZN(U3134) );
  INV_X1 U6107 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4933) );
  INV_X1 U6108 ( .A(n4924), .ZN(n4925) );
  AOI22_X1 U6109 ( .A1(n6399), .A2(n4926), .B1(n6413), .B2(n4925), .ZN(n4932)
         );
  INV_X1 U6110 ( .A(n4927), .ZN(n4930) );
  INV_X1 U6111 ( .A(n4928), .ZN(n4929) );
  AOI22_X1 U6112 ( .A1(n6355), .A2(n4930), .B1(n4929), .B2(n6400), .ZN(n4931)
         );
  OAI211_X1 U6113 ( .C1(n4934), .C2(n4933), .A(n4932), .B(n4931), .ZN(U3132)
         );
  INV_X1 U6114 ( .A(n4943), .ZN(n4935) );
  OAI21_X1 U6115 ( .B1(n4943), .B2(n6604), .A(n6401), .ZN(n4942) );
  NAND3_X1 U6116 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6474), .A3(n4936), .ZN(n5824) );
  NOR2_X1 U6117 ( .A1(n4937), .A2(n5824), .ZN(n4960) );
  AOI21_X1 U6118 ( .B1(n4938), .B2(n5831), .A(n4960), .ZN(n4941) );
  INV_X1 U6119 ( .A(n4941), .ZN(n4940) );
  AOI21_X1 U6120 ( .B1(n6406), .B2(n5824), .A(n6405), .ZN(n4939) );
  OAI22_X1 U6121 ( .A1(n4942), .A2(n4941), .B1(n5874), .B2(n5824), .ZN(n4958)
         );
  AOI22_X1 U6122 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4959), .B1(n6460), 
        .B2(n4958), .ZN(n4945) );
  AOI22_X1 U6123 ( .A1(n5907), .A2(n6457), .B1(n4960), .B2(n6456), .ZN(n4944)
         );
  OAI211_X1 U6124 ( .C1(n5862), .C2(n6465), .A(n4945), .B(n4944), .ZN(U3099)
         );
  AOI22_X1 U6125 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4959), .B1(n6419), 
        .B2(n4958), .ZN(n4947) );
  AOI22_X1 U6126 ( .A1(n5907), .A2(n6418), .B1(n4960), .B2(n6417), .ZN(n4946)
         );
  OAI211_X1 U6127 ( .C1(n5862), .C2(n6422), .A(n4947), .B(n4946), .ZN(U3093)
         );
  AOI22_X1 U6128 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4959), .B1(n6443), 
        .B2(n4958), .ZN(n4949) );
  AOI22_X1 U6129 ( .A1(n5907), .A2(n5807), .B1(n4960), .B2(n6441), .ZN(n4948)
         );
  OAI211_X1 U6130 ( .C1(n5862), .C2(n5849), .A(n4949), .B(n4948), .ZN(U3097)
         );
  AOI22_X1 U6131 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4959), .B1(n6437), 
        .B2(n4958), .ZN(n4951) );
  AOI22_X1 U6132 ( .A1(n5907), .A2(n6436), .B1(n4960), .B2(n6435), .ZN(n4950)
         );
  OAI211_X1 U6133 ( .C1(n5862), .C2(n6440), .A(n4951), .B(n4950), .ZN(U3096)
         );
  AOI22_X1 U6134 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4959), .B1(n6431), 
        .B2(n4958), .ZN(n4953) );
  AOI22_X1 U6135 ( .A1(n5907), .A2(n5798), .B1(n4960), .B2(n6429), .ZN(n4952)
         );
  OAI211_X1 U6136 ( .C1(n5862), .C2(n5842), .A(n4953), .B(n4952), .ZN(U3095)
         );
  AOI22_X1 U6137 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4959), .B1(n6425), 
        .B2(n4958), .ZN(n4955) );
  AOI22_X1 U6138 ( .A1(n5907), .A2(n6424), .B1(n4960), .B2(n6423), .ZN(n4954)
         );
  OAI211_X1 U6139 ( .C1(n5862), .C2(n6428), .A(n4955), .B(n4954), .ZN(U3094)
         );
  AOI22_X1 U6140 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4959), .B1(n6450), 
        .B2(n4958), .ZN(n4957) );
  AOI22_X1 U6141 ( .A1(n5907), .A2(n6386), .B1(n4960), .B2(n6447), .ZN(n4956)
         );
  OAI211_X1 U6142 ( .C1(n5862), .C2(n6389), .A(n4957), .B(n4956), .ZN(U3098)
         );
  AOI22_X1 U6143 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4959), .B1(n6413), 
        .B2(n4958), .ZN(n4962) );
  AOI22_X1 U6144 ( .A1(n5907), .A2(n6400), .B1(n6399), .B2(n4960), .ZN(n4961)
         );
  OAI211_X1 U6145 ( .C1(n5862), .C2(n6416), .A(n4962), .B(n4961), .ZN(U3092)
         );
  OAI21_X1 U6146 ( .B1(n4965), .B2(n4964), .A(n4963), .ZN(n5588) );
  XNOR2_X1 U6147 ( .A(n4966), .B(n5056), .ZN(n6215) );
  AOI22_X1 U6148 ( .A1(n6215), .A2(n6065), .B1(EBX_REG_8__SCAN_IN), .B2(n5337), 
        .ZN(n4967) );
  OAI21_X1 U6149 ( .B1(n5588), .B2(n5371), .A(n4967), .ZN(U2851) );
  AOI22_X1 U6150 ( .A1(n5422), .A2(DATAI_8_), .B1(n6075), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4968) );
  OAI21_X1 U6151 ( .B1(n5588), .B2(n5424), .A(n4968), .ZN(U2883) );
  NAND2_X1 U6152 ( .A1(n2964), .A2(n6275), .ZN(n5863) );
  INV_X1 U6153 ( .A(n5863), .ZN(n4969) );
  NAND3_X1 U6154 ( .A1(n4994), .A2(n6401), .A3(n6396), .ZN(n4970) );
  AOI21_X1 U6155 ( .B1(n6283), .B2(n4970), .A(n6359), .ZN(n4972) );
  NOR2_X1 U6156 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6364), .ZN(n6349)
         );
  OAI21_X1 U6157 ( .B1(n6588), .B2(n6349), .A(n6397), .ZN(n4971) );
  NAND2_X1 U6158 ( .A1(n4973), .A2(n6359), .ZN(n4975) );
  NOR2_X1 U6159 ( .A1(n5008), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6280)
         );
  NAND2_X1 U6160 ( .A1(n5869), .A2(n6280), .ZN(n4974) );
  OAI22_X1 U6161 ( .A1(n6396), .A2(n6329), .B1(n6347), .B2(n5886), .ZN(n4977)
         );
  INV_X1 U6162 ( .A(n6349), .ZN(n4995) );
  OAI22_X1 U6163 ( .A1(n5792), .A2(n4995), .B1(n4994), .B2(n6428), .ZN(n4976)
         );
  AOI211_X1 U6164 ( .C1(n6351), .C2(INSTQUEUE_REG_6__2__SCAN_IN), .A(n4977), 
        .B(n4976), .ZN(n4978) );
  INV_X1 U6165 ( .A(n4978), .ZN(U3070) );
  OAI22_X1 U6166 ( .A1(n6396), .A2(n6373), .B1(n6347), .B2(n5882), .ZN(n4980)
         );
  OAI22_X1 U6167 ( .A1(n5788), .A2(n4995), .B1(n4994), .B2(n6422), .ZN(n4979)
         );
  AOI211_X1 U6168 ( .C1(n6351), .C2(INSTQUEUE_REG_6__1__SCAN_IN), .A(n4980), 
        .B(n4979), .ZN(n4981) );
  INV_X1 U6169 ( .A(n4981), .ZN(U3069) );
  OAI22_X1 U6170 ( .A1(n6396), .A2(n6308), .B1(n6347), .B2(n5909), .ZN(n4983)
         );
  OAI22_X1 U6171 ( .A1(n5817), .A2(n4995), .B1(n4994), .B2(n6465), .ZN(n4982)
         );
  AOI211_X1 U6172 ( .C1(n6351), .C2(INSTQUEUE_REG_6__7__SCAN_IN), .A(n4983), 
        .B(n4982), .ZN(n4984) );
  INV_X1 U6173 ( .A(n4984), .ZN(U3075) );
  OAI22_X1 U6174 ( .A1(n6396), .A2(n6381), .B1(n6347), .B2(n5894), .ZN(n4986)
         );
  OAI22_X1 U6175 ( .A1(n5801), .A2(n4995), .B1(n4994), .B2(n6440), .ZN(n4985)
         );
  AOI211_X1 U6176 ( .C1(n6351), .C2(INSTQUEUE_REG_6__4__SCAN_IN), .A(n4986), 
        .B(n4985), .ZN(n4987) );
  INV_X1 U6177 ( .A(n4987), .ZN(U3072) );
  OAI22_X1 U6178 ( .A1(n6396), .A2(n6434), .B1(n6347), .B2(n5890), .ZN(n4989)
         );
  OAI22_X1 U6179 ( .A1(n5796), .A2(n4995), .B1(n4994), .B2(n5842), .ZN(n4988)
         );
  AOI211_X1 U6180 ( .C1(n6351), .C2(INSTQUEUE_REG_6__3__SCAN_IN), .A(n4989), 
        .B(n4988), .ZN(n4990) );
  INV_X1 U6181 ( .A(n4990), .ZN(U3071) );
  OAI22_X1 U6182 ( .A1(n6396), .A2(n6454), .B1(n6347), .B2(n5902), .ZN(n4992)
         );
  OAI22_X1 U6183 ( .A1(n5810), .A2(n4995), .B1(n4994), .B2(n6389), .ZN(n4991)
         );
  AOI211_X1 U6184 ( .C1(n6351), .C2(INSTQUEUE_REG_6__6__SCAN_IN), .A(n4992), 
        .B(n4991), .ZN(n4993) );
  INV_X1 U6185 ( .A(n4993), .ZN(U3074) );
  OAI22_X1 U6186 ( .A1(n6396), .A2(n6446), .B1(n6347), .B2(n5898), .ZN(n4997)
         );
  OAI22_X1 U6187 ( .A1(n5805), .A2(n4995), .B1(n4994), .B2(n5849), .ZN(n4996)
         );
  AOI211_X1 U6188 ( .C1(n6351), .C2(INSTQUEUE_REG_6__5__SCAN_IN), .A(n4997), 
        .B(n4996), .ZN(n4998) );
  INV_X1 U6189 ( .A(n4998), .ZN(U3073) );
  INV_X1 U6190 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6693) );
  XOR2_X1 U6191 ( .A(n5000), .B(n4999), .Z(n5049) );
  NAND2_X1 U6192 ( .A1(n5049), .A2(n4264), .ZN(n5005) );
  AND2_X1 U6193 ( .A1(n5002), .A2(n5001), .ZN(n5003) );
  NOR2_X1 U6194 ( .A1(n4966), .A2(n5003), .ZN(n6222) );
  NAND2_X1 U6195 ( .A1(n6065), .A2(n6222), .ZN(n5004) );
  OAI211_X1 U6196 ( .C1(n6693), .C2(n6067), .A(n5005), .B(n5004), .ZN(U2852)
         );
  INV_X1 U6197 ( .A(n5821), .ZN(n5006) );
  OAI21_X1 U6198 ( .B1(n5040), .B2(n6458), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5007) );
  OAI211_X1 U6199 ( .C1(n5778), .C2(n5773), .A(n5007), .B(n6401), .ZN(n5013)
         );
  NAND2_X1 U6200 ( .A1(n5009), .A2(n5008), .ZN(n5014) );
  AOI21_X1 U6201 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5014), .A(n5010), .ZN(
        n5827) );
  OR2_X1 U6202 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5011), .ZN(n5038)
         );
  AOI21_X1 U6203 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5038), .A(n6279), .ZN(
        n5012) );
  NAND2_X1 U6204 ( .A1(n5036), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5017)
         );
  INV_X1 U6205 ( .A(n5014), .ZN(n5830) );
  AOI22_X1 U6206 ( .A1(n5832), .A2(n5777), .B1(n5830), .B2(n5869), .ZN(n5037)
         );
  OAI22_X1 U6207 ( .A1(n5792), .A2(n5038), .B1(n5037), .B2(n5886), .ZN(n5015)
         );
  AOI21_X1 U6208 ( .B1(n6424), .B2(n5040), .A(n5015), .ZN(n5016) );
  OAI211_X1 U6209 ( .C1(n6453), .C2(n6428), .A(n5017), .B(n5016), .ZN(U3118)
         );
  NAND2_X1 U6210 ( .A1(n5036), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5020)
         );
  OAI22_X1 U6211 ( .A1(n5805), .A2(n5038), .B1(n5037), .B2(n5898), .ZN(n5018)
         );
  AOI21_X1 U6212 ( .B1(n5807), .B2(n5040), .A(n5018), .ZN(n5019) );
  OAI211_X1 U6213 ( .C1(n6453), .C2(n5849), .A(n5020), .B(n5019), .ZN(U3121)
         );
  NAND2_X1 U6214 ( .A1(n5036), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5023)
         );
  OAI22_X1 U6215 ( .A1(n5784), .A2(n5038), .B1(n5037), .B2(n5878), .ZN(n5021)
         );
  AOI21_X1 U6216 ( .B1(n6400), .B2(n5040), .A(n5021), .ZN(n5022) );
  OAI211_X1 U6217 ( .C1(n6453), .C2(n6416), .A(n5023), .B(n5022), .ZN(U3116)
         );
  NAND2_X1 U6218 ( .A1(n5036), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5026)
         );
  OAI22_X1 U6219 ( .A1(n5817), .A2(n5038), .B1(n5037), .B2(n5909), .ZN(n5024)
         );
  AOI21_X1 U6220 ( .B1(n6457), .B2(n5040), .A(n5024), .ZN(n5025) );
  OAI211_X1 U6221 ( .C1(n6453), .C2(n6465), .A(n5026), .B(n5025), .ZN(U3123)
         );
  NAND2_X1 U6222 ( .A1(n5036), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5029)
         );
  OAI22_X1 U6223 ( .A1(n5788), .A2(n5038), .B1(n5037), .B2(n5882), .ZN(n5027)
         );
  AOI21_X1 U6224 ( .B1(n6418), .B2(n5040), .A(n5027), .ZN(n5028) );
  OAI211_X1 U6225 ( .C1(n6453), .C2(n6422), .A(n5029), .B(n5028), .ZN(U3117)
         );
  NAND2_X1 U6226 ( .A1(n5036), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5032)
         );
  OAI22_X1 U6227 ( .A1(n5801), .A2(n5038), .B1(n5037), .B2(n5894), .ZN(n5030)
         );
  AOI21_X1 U6228 ( .B1(n6436), .B2(n5040), .A(n5030), .ZN(n5031) );
  OAI211_X1 U6229 ( .C1(n6453), .C2(n6440), .A(n5032), .B(n5031), .ZN(U3120)
         );
  NAND2_X1 U6230 ( .A1(n5036), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5035)
         );
  OAI22_X1 U6231 ( .A1(n5810), .A2(n5038), .B1(n5037), .B2(n5902), .ZN(n5033)
         );
  AOI21_X1 U6232 ( .B1(n6386), .B2(n5040), .A(n5033), .ZN(n5034) );
  OAI211_X1 U6233 ( .C1(n6453), .C2(n6389), .A(n5035), .B(n5034), .ZN(U3122)
         );
  NAND2_X1 U6234 ( .A1(n5036), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5042)
         );
  OAI22_X1 U6235 ( .A1(n5796), .A2(n5038), .B1(n5037), .B2(n5890), .ZN(n5039)
         );
  AOI21_X1 U6236 ( .B1(n5798), .B2(n5040), .A(n5039), .ZN(n5041) );
  OAI211_X1 U6237 ( .C1(n6453), .C2(n5842), .A(n5042), .B(n5041), .ZN(U3119)
         );
  OAI21_X1 U6238 ( .B1(n5043), .B2(n5045), .A(n5044), .ZN(n6223) );
  NAND2_X1 U6239 ( .A1(n6233), .A2(REIP_REG_7__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U6240 ( .A1(n5565), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5046)
         );
  OAI211_X1 U6241 ( .C1(n6182), .C2(n6008), .A(n6220), .B(n5046), .ZN(n5047)
         );
  AOI21_X1 U6242 ( .B1(n5049), .B2(n6177), .A(n5047), .ZN(n5048) );
  OAI21_X1 U6243 ( .B1(n6159), .B2(n6223), .A(n5048), .ZN(U2979) );
  INV_X1 U6244 ( .A(n5049), .ZN(n6013) );
  OAI222_X1 U6245 ( .A1(n5417), .A2(n4674), .B1(n5424), .B2(n6013), .C1(n5050), 
        .C2(n5416), .ZN(U2884) );
  NAND2_X1 U6246 ( .A1(n4963), .A2(n5052), .ZN(n5053) );
  NAND2_X1 U6247 ( .A1(n5051), .A2(n5053), .ZN(n5995) );
  AOI22_X1 U6248 ( .A1(n5422), .A2(DATAI_9_), .B1(n6075), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n5054) );
  OAI21_X1 U6249 ( .B1(n5995), .B2(n5424), .A(n5054), .ZN(U2882) );
  INV_X1 U6250 ( .A(n5056), .ZN(n5059) );
  INV_X1 U6251 ( .A(n5057), .ZN(n5058) );
  AOI21_X1 U6252 ( .B1(n4966), .B2(n5059), .A(n5058), .ZN(n5060) );
  OR2_X1 U6253 ( .A1(n5055), .A2(n5060), .ZN(n6204) );
  INV_X1 U6254 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5998) );
  OAI222_X1 U6255 ( .A1(n6204), .A2(n5369), .B1(n5998), .B2(n6067), .C1(n5995), 
        .C2(n5371), .ZN(U2850) );
  INV_X1 U6256 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6668) );
  AOI22_X1 U6257 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6668), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6269), .ZN(n5076) );
  NOR3_X1 U6258 ( .A1(n6749), .A2(n6260), .A3(n5076), .ZN(n5062) );
  INV_X1 U6259 ( .A(n4593), .ZN(n5064) );
  NOR3_X1 U6260 ( .A1(n6502), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n5064), 
        .ZN(n5061) );
  AOI211_X1 U6261 ( .C1(n6510), .C2(n5063), .A(n5062), .B(n5061), .ZN(n5066)
         );
  AOI21_X1 U6262 ( .B1(n5074), .B2(n5064), .A(n5078), .ZN(n5065) );
  OAI22_X1 U6263 ( .A1(n5066), .A2(n5078), .B1(n5065), .B2(n3857), .ZN(U3459)
         );
  NAND2_X1 U6264 ( .A1(n5865), .A2(n5067), .ZN(n5072) );
  OAI21_X1 U6265 ( .B1(n5068), .B2(n5070), .A(n5069), .ZN(n5071) );
  OAI211_X1 U6266 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n5073), .A(n5072), .B(n5071), .ZN(n6468) );
  NOR2_X1 U6267 ( .A1(n6749), .A2(n6260), .ZN(n5075) );
  AOI222_X1 U6268 ( .A1(n6468), .A2(n6510), .B1(n5076), .B2(n5075), .C1(n5068), 
        .C2(n5074), .ZN(n5079) );
  OAI22_X1 U6269 ( .A1(n5079), .A2(n5078), .B1(n5077), .B2(n3417), .ZN(U3460)
         );
  INV_X1 U6270 ( .A(n5080), .ZN(n5098) );
  OAI22_X1 U6271 ( .A1(n5098), .A2(n5369), .B1(n6067), .B2(n5081), .ZN(U2828)
         );
  INV_X1 U6272 ( .A(n6055), .ZN(n5083) );
  AOI22_X1 U6273 ( .A1(n5565), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n6233), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n5082) );
  OAI21_X1 U6274 ( .B1(n6182), .B2(n5083), .A(n5082), .ZN(n5084) );
  INV_X1 U6275 ( .A(n5084), .ZN(n5089) );
  XNOR2_X1 U6276 ( .A(n5085), .B(n6256), .ZN(n5087) );
  OR2_X1 U6277 ( .A1(n5086), .A2(n5087), .ZN(n6247) );
  NAND2_X1 U6278 ( .A1(n5087), .A2(n5086), .ZN(n6246) );
  NAND3_X1 U6279 ( .A1(n6247), .A2(n3910), .A3(n6246), .ZN(n5088) );
  OAI211_X1 U6280 ( .C1(n6052), .C2(n6157), .A(n5089), .B(n5088), .ZN(U2983)
         );
  NAND2_X1 U6281 ( .A1(n5099), .A2(n6025), .ZN(n5097) );
  INV_X1 U6282 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6571) );
  AOI21_X1 U6283 ( .B1(n6775), .B2(n6571), .A(n5116), .ZN(n5109) );
  OAI21_X1 U6284 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5980), .A(n5109), .ZN(n5095) );
  INV_X1 U6285 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6660) );
  NOR4_X1 U6286 ( .A1(n5105), .A2(REIP_REG_31__SCAN_IN), .A3(n6660), .A4(n6571), .ZN(n5094) );
  NAND2_X1 U6287 ( .A1(n5090), .A2(EBX_REG_31__SCAN_IN), .ZN(n5091) );
  OAI22_X1 U6288 ( .A1(n6047), .A2(n5092), .B1(n5310), .B2(n5091), .ZN(n5093)
         );
  AOI211_X1 U6289 ( .C1(n5095), .C2(REIP_REG_31__SCAN_IN), .A(n5094), .B(n5093), .ZN(n5096) );
  OAI211_X1 U6290 ( .C1(n5098), .C2(n6044), .A(n5097), .B(n5096), .ZN(U2796)
         );
  NAND3_X1 U6291 ( .A1(n5099), .A2(n5373), .A3(n5416), .ZN(n5102) );
  AOI22_X1 U6292 ( .A1(n6072), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6075), .ZN(n5101) );
  NAND2_X1 U6293 ( .A1(n5102), .A2(n5101), .ZN(U2860) );
  INV_X1 U6294 ( .A(n5103), .ZN(n5596) );
  OAI22_X1 U6295 ( .A1(n5104), .A2(n6047), .B1(n6778), .B2(n5430), .ZN(n5107)
         );
  NOR3_X1 U6296 ( .A1(n5105), .A2(REIP_REG_30__SCAN_IN), .A3(n6571), .ZN(n5106) );
  AOI211_X1 U6297 ( .C1(n6780), .C2(EBX_REG_30__SCAN_IN), .A(n5107), .B(n5106), 
        .ZN(n5108) );
  OAI21_X1 U6298 ( .B1(n5109), .B2(n6660), .A(n5108), .ZN(n5110) );
  AOI21_X1 U6299 ( .B1(n5596), .B2(n6787), .A(n5110), .ZN(n5111) );
  OAI21_X1 U6300 ( .B1(n5377), .B2(n6790), .A(n5111), .ZN(U2797) );
  NAND2_X1 U6301 ( .A1(n5112), .A2(n5113), .ZN(n5114) );
  INV_X1 U6302 ( .A(n5382), .ZN(n5452) );
  AND2_X1 U6303 ( .A1(n5129), .A2(REIP_REG_27__SCAN_IN), .ZN(n5117) );
  MUX2_X1 U6304 ( .A(n5117), .B(n5116), .S(REIP_REG_28__SCAN_IN), .Z(n5125) );
  NAND2_X1 U6305 ( .A1(n2993), .A2(n5118), .ZN(n5119) );
  NAND2_X1 U6306 ( .A1(n5120), .A2(n5119), .ZN(n5610) );
  INV_X1 U6307 ( .A(n5450), .ZN(n5121) );
  AOI22_X1 U6308 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n6779), .B1(n6054), 
        .B2(n5121), .ZN(n5123) );
  NAND2_X1 U6309 ( .A1(n6780), .A2(EBX_REG_28__SCAN_IN), .ZN(n5122) );
  OAI211_X1 U6310 ( .C1(n5610), .C2(n6044), .A(n5123), .B(n5122), .ZN(n5124)
         );
  AOI211_X1 U6311 ( .C1(n5452), .C2(n6025), .A(n5125), .B(n5124), .ZN(n5126)
         );
  INV_X1 U6312 ( .A(n5126), .ZN(U2799) );
  OAI21_X1 U6313 ( .B1(n5128), .B2(n5127), .A(n5112), .ZN(n5456) );
  INV_X1 U6314 ( .A(n5129), .ZN(n5137) );
  NAND2_X1 U6315 ( .A1(n4225), .A2(n5130), .ZN(n5131) );
  AND2_X1 U6316 ( .A1(n2993), .A2(n5131), .ZN(n5619) );
  NAND2_X1 U6317 ( .A1(n5619), .A2(n6787), .ZN(n5136) );
  INV_X1 U6318 ( .A(n5132), .ZN(n5458) );
  OAI22_X1 U6319 ( .A1(n5133), .A2(n6047), .B1(n6778), .B2(n5458), .ZN(n5134)
         );
  AOI21_X1 U6320 ( .B1(n6780), .B2(EBX_REG_27__SCAN_IN), .A(n5134), .ZN(n5135)
         );
  OAI211_X1 U6321 ( .C1(REIP_REG_27__SCAN_IN), .C2(n5137), .A(n5136), .B(n5135), .ZN(n5138) );
  AOI21_X1 U6322 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5146), .A(n5138), .ZN(n5139) );
  OAI21_X1 U6323 ( .B1(n5456), .B2(n6790), .A(n5139), .ZN(U2800) );
  NAND2_X1 U6324 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5140) );
  INV_X1 U6325 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6569) );
  OAI21_X1 U6326 ( .B1(n5167), .B2(n5140), .A(n6569), .ZN(n5145) );
  INV_X1 U6327 ( .A(n5467), .ZN(n5141) );
  AOI22_X1 U6328 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6779), .B1(n6054), 
        .B2(n5141), .ZN(n5143) );
  NAND2_X1 U6329 ( .A1(n6780), .A2(EBX_REG_26__SCAN_IN), .ZN(n5142) );
  OAI211_X1 U6330 ( .C1(n5626), .C2(n6044), .A(n5143), .B(n5142), .ZN(n5144)
         );
  AOI21_X1 U6331 ( .B1(n5146), .B2(n5145), .A(n5144), .ZN(n5147) );
  OAI21_X1 U6332 ( .B1(n5387), .B2(n6790), .A(n5147), .ZN(U2801) );
  INV_X1 U6333 ( .A(n5478), .ZN(n5390) );
  AND2_X1 U6334 ( .A1(n5150), .A2(n5149), .ZN(n5151) );
  NOR2_X1 U6335 ( .A1(n5152), .A2(n5151), .ZN(n5636) );
  INV_X1 U6336 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6566) );
  NOR2_X1 U6337 ( .A1(n5181), .A2(n6566), .ZN(n5159) );
  XNOR2_X1 U6338 ( .A(REIP_REG_24__SCAN_IN), .B(REIP_REG_25__SCAN_IN), .ZN(
        n5157) );
  INV_X1 U6339 ( .A(n5153), .ZN(n5476) );
  OAI22_X1 U6340 ( .A1(n5154), .A2(n6047), .B1(n6778), .B2(n5476), .ZN(n5155)
         );
  AOI21_X1 U6341 ( .B1(n6780), .B2(EBX_REG_25__SCAN_IN), .A(n5155), .ZN(n5156)
         );
  OAI21_X1 U6342 ( .B1(n5167), .B2(n5157), .A(n5156), .ZN(n5158) );
  AOI211_X1 U6343 ( .C1(n5636), .C2(n6787), .A(n5159), .B(n5158), .ZN(n5160)
         );
  OAI21_X1 U6344 ( .B1(n5390), .B2(n6790), .A(n5160), .ZN(U2802) );
  INV_X1 U6345 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6564) );
  INV_X1 U6346 ( .A(n5161), .ZN(n5163) );
  NAND2_X1 U6347 ( .A1(n5484), .A2(n6025), .ZN(n5170) );
  OAI22_X1 U6348 ( .A1(n6638), .A2(n6047), .B1(n6778), .B2(n5482), .ZN(n5165)
         );
  AOI21_X1 U6349 ( .B1(n6780), .B2(EBX_REG_24__SCAN_IN), .A(n5165), .ZN(n5166)
         );
  OAI21_X1 U6350 ( .B1(n5167), .B2(REIP_REG_24__SCAN_IN), .A(n5166), .ZN(n5168) );
  AOI21_X1 U6351 ( .B1(n5338), .B2(n6787), .A(n5168), .ZN(n5169) );
  OAI211_X1 U6352 ( .C1(n5181), .C2(n6564), .A(n5170), .B(n5169), .ZN(U2803)
         );
  AOI21_X1 U6353 ( .B1(n5201), .B2(n5171), .A(REIP_REG_23__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U6354 ( .A1(n5496), .A2(n6025), .ZN(n5180) );
  OAI22_X1 U6355 ( .A1(n5173), .A2(n6047), .B1(n6778), .B2(n5494), .ZN(n5178)
         );
  OR2_X1 U6356 ( .A1(n5174), .A2(n5175), .ZN(n5176) );
  NAND2_X1 U6357 ( .A1(n4376), .A2(n5176), .ZN(n5647) );
  NOR2_X1 U6358 ( .A1(n5647), .A2(n6044), .ZN(n5177) );
  AOI211_X1 U6359 ( .C1(EBX_REG_23__SCAN_IN), .C2(n6780), .A(n5178), .B(n5177), 
        .ZN(n5179) );
  OAI211_X1 U6360 ( .C1(n5182), .C2(n5181), .A(n5180), .B(n5179), .ZN(U2804)
         );
  NAND2_X1 U6361 ( .A1(n5502), .A2(n5183), .ZN(n5186) );
  NAND2_X1 U6362 ( .A1(n5184), .A2(n3492), .ZN(n5185) );
  INV_X1 U6364 ( .A(n5504), .ZN(n5399) );
  AOI21_X1 U6365 ( .B1(n5192), .B2(n5191), .A(n5274), .ZN(n5217) );
  NOR2_X1 U6366 ( .A1(n2976), .A2(n5193), .ZN(n5194) );
  OR2_X1 U6367 ( .A1(n5174), .A2(n5194), .ZN(n5654) );
  OAI22_X1 U6368 ( .A1(n3019), .A2(n6047), .B1(n6778), .B2(n5502), .ZN(n5195)
         );
  AOI21_X1 U6369 ( .B1(n6780), .B2(EBX_REG_22__SCAN_IN), .A(n5195), .ZN(n5198)
         );
  XOR2_X1 U6370 ( .A(REIP_REG_22__SCAN_IN), .B(REIP_REG_21__SCAN_IN), .Z(n5196) );
  NAND2_X1 U6371 ( .A1(n5201), .A2(n5196), .ZN(n5197) );
  OAI211_X1 U6372 ( .C1(n5654), .C2(n6044), .A(n5198), .B(n5197), .ZN(n5199)
         );
  AOI21_X1 U6373 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5217), .A(n5199), .ZN(n5200) );
  OAI21_X1 U6374 ( .B1(n5399), .B2(n6790), .A(n5200), .ZN(U2805) );
  INV_X1 U6375 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6670) );
  NAND2_X1 U6376 ( .A1(n5201), .A2(n6670), .ZN(n5203) );
  AOI22_X1 U6377 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n6779), .B1(n6054), 
        .B2(n5510), .ZN(n5202) );
  OAI211_X1 U6378 ( .C1(n5204), .C2(n6029), .A(n5203), .B(n5202), .ZN(n5206)
         );
  NOR2_X1 U6379 ( .A1(n5663), .A2(n6044), .ZN(n5205) );
  AOI211_X1 U6380 ( .C1(n5217), .C2(REIP_REG_21__SCAN_IN), .A(n5206), .B(n5205), .ZN(n5207) );
  OAI21_X1 U6381 ( .B1(n5402), .B2(n6790), .A(n5207), .ZN(U2806) );
  OAI22_X1 U6382 ( .A1(n5210), .A2(n6047), .B1(n6778), .B2(n5209), .ZN(n5216)
         );
  INV_X1 U6383 ( .A(n5226), .ZN(n5212) );
  MUX2_X1 U6384 ( .A(n5212), .B(n2963), .S(n5211), .Z(n5214) );
  XNOR2_X1 U6385 ( .A(n5214), .B(n5213), .ZN(n5671) );
  NOR2_X1 U6386 ( .A1(n5671), .A2(n6044), .ZN(n5215) );
  AOI211_X1 U6387 ( .C1(n6780), .C2(EBX_REG_20__SCAN_IN), .A(n5216), .B(n5215), 
        .ZN(n5220) );
  NOR2_X1 U6388 ( .A1(n5244), .A2(n5233), .ZN(n5218) );
  OAI21_X1 U6389 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5218), .A(n5217), .ZN(n5219) );
  OAI211_X1 U6390 ( .C1(n5208), .C2(n6790), .A(n5220), .B(n5219), .ZN(U2807)
         );
  NOR2_X1 U6391 ( .A1(n5221), .A2(n5274), .ZN(n5251) );
  INV_X1 U6392 ( .A(n5223), .ZN(n5225) );
  MUX2_X1 U6393 ( .A(n5226), .B(n5225), .S(n5224), .Z(n5242) );
  NAND2_X1 U6394 ( .A1(n5222), .A2(n5242), .ZN(n5241) );
  INV_X1 U6395 ( .A(n5227), .ZN(n5228) );
  XNOR2_X1 U6396 ( .A(n5241), .B(n5228), .ZN(n5685) );
  NAND2_X1 U6397 ( .A1(n5307), .A2(n5229), .ZN(n6781) );
  AOI21_X1 U6398 ( .B1(n6779), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6033), 
        .ZN(n5230) );
  OAI21_X1 U6399 ( .B1(n5231), .B2(n6778), .A(n5230), .ZN(n5232) );
  AOI21_X1 U6400 ( .B1(EBX_REG_19__SCAN_IN), .B2(n6780), .A(n5232), .ZN(n5236)
         );
  INV_X1 U6401 ( .A(n5244), .ZN(n5234) );
  OAI211_X1 U6402 ( .C1(REIP_REG_18__SCAN_IN), .C2(REIP_REG_19__SCAN_IN), .A(
        n5234), .B(n5233), .ZN(n5235) );
  OAI211_X1 U6403 ( .C1(n5685), .C2(n6044), .A(n5236), .B(n5235), .ZN(n5237)
         );
  AOI21_X1 U6404 ( .B1(n5251), .B2(REIP_REG_19__SCAN_IN), .A(n5237), .ZN(n5238) );
  OAI21_X1 U6405 ( .B1(n5407), .B2(n6790), .A(n5238), .ZN(U2808) );
  OAI21_X1 U6406 ( .B1(n5240), .B2(n5239), .A(n3754), .ZN(n5518) );
  OAI21_X1 U6407 ( .B1(n5222), .B2(n5242), .A(n5241), .ZN(n5694) );
  AOI21_X1 U6408 ( .B1(n6779), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6033), 
        .ZN(n5243) );
  OAI21_X1 U6409 ( .B1(n5520), .B2(n6778), .A(n5243), .ZN(n5245) );
  XNOR2_X1 U6410 ( .A(n3940), .B(n5246), .ZN(n6069) );
  NOR2_X1 U6411 ( .A1(n5247), .A2(n5248), .ZN(n5249) );
  OR2_X1 U6412 ( .A1(n5222), .A2(n5249), .ZN(n5703) );
  INV_X1 U6413 ( .A(n5250), .ZN(n5252) );
  OAI21_X1 U6414 ( .B1(REIP_REG_17__SCAN_IN), .B2(n5252), .A(n5251), .ZN(n5255) );
  OAI22_X1 U6415 ( .A1(n5344), .A2(n6029), .B1(n6743), .B2(n6047), .ZN(n5253)
         );
  AOI211_X1 U6416 ( .C1(n6054), .C2(n5527), .A(n5253), .B(n6033), .ZN(n5254)
         );
  OAI211_X1 U6417 ( .C1(n6044), .C2(n5703), .A(n5255), .B(n5254), .ZN(n5256)
         );
  AOI21_X1 U6418 ( .B1(n6069), .B2(n6025), .A(n5256), .ZN(n5257) );
  INV_X1 U6419 ( .A(n5257), .ZN(U2810) );
  AOI21_X1 U6420 ( .B1(n5260), .B2(n5258), .A(n5259), .ZN(n5544) );
  INV_X1 U6421 ( .A(n5544), .ZN(n5411) );
  NAND2_X1 U6422 ( .A1(n5362), .A2(n5262), .ZN(n5263) );
  AND2_X1 U6423 ( .A1(n5261), .A2(n5263), .ZN(n5726) );
  NAND3_X1 U6424 ( .A1(n6030), .A2(REIP_REG_15__SCAN_IN), .A3(n5965), .ZN(
        n5264) );
  OAI21_X1 U6425 ( .B1(n6778), .B2(n5542), .A(n5264), .ZN(n5267) );
  INV_X1 U6426 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5353) );
  INV_X1 U6427 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6551) );
  AOI22_X1 U6428 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n6779), .B1(n5960), 
        .B2(n6551), .ZN(n5265) );
  OAI211_X1 U6429 ( .C1(n6029), .C2(n5353), .A(n5265), .B(n6781), .ZN(n5266)
         );
  AOI211_X1 U6430 ( .C1(n5726), .C2(n6787), .A(n5267), .B(n5266), .ZN(n5268)
         );
  OAI21_X1 U6431 ( .B1(n5411), .B2(n6790), .A(n5268), .ZN(U2812) );
  NAND2_X1 U6432 ( .A1(n5051), .A2(n5270), .ZN(n5271) );
  AND2_X1 U6433 ( .A1(n5269), .A2(n5271), .ZN(n5569) );
  INV_X1 U6434 ( .A(n5272), .ZN(n5273) );
  OAI21_X1 U6435 ( .B1(n3017), .B2(n5273), .A(n6030), .ZN(n6019) );
  OAI21_X1 U6436 ( .B1(n5275), .B2(n5274), .A(n6019), .ZN(n6003) );
  OAI21_X1 U6437 ( .B1(n5055), .B2(n5277), .A(n5276), .ZN(n6197) );
  INV_X1 U6438 ( .A(n6197), .ZN(n5278) );
  AOI22_X1 U6439 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6780), .B1(n6787), .B2(n5278), .ZN(n5280) );
  AOI21_X1 U6440 ( .B1(n6779), .B2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6033), 
        .ZN(n5279) );
  OAI211_X1 U6441 ( .C1(n5567), .C2(n6778), .A(n5280), .B(n5279), .ZN(n5281)
         );
  AOI21_X1 U6442 ( .B1(n6003), .B2(REIP_REG_10__SCAN_IN), .A(n5281), .ZN(n5286) );
  NOR2_X1 U6443 ( .A1(n5980), .A2(n6031), .ZN(n6040) );
  INV_X1 U6444 ( .A(n6040), .ZN(n5282) );
  NOR3_X1 U6445 ( .A1(n5282), .A2(n6740), .A3(n6667), .ZN(n6007) );
  NAND2_X1 U6446 ( .A1(n6007), .A2(REIP_REG_6__SCAN_IN), .ZN(n6012) );
  NOR2_X1 U6447 ( .A1(n5283), .A2(n6012), .ZN(n6004) );
  AOI21_X1 U6448 ( .B1(n6542), .B2(n6543), .A(n5985), .ZN(n5284) );
  NAND2_X1 U6449 ( .A1(n6004), .A2(n5284), .ZN(n5285) );
  OAI211_X1 U6450 ( .C1(n5425), .C2(n6790), .A(n5286), .B(n5285), .ZN(U2817)
         );
  INV_X1 U6451 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6017) );
  INV_X1 U6452 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6541) );
  OAI21_X1 U6453 ( .B1(n6017), .B2(n6012), .A(n6541), .ZN(n5287) );
  NAND2_X1 U6454 ( .A1(n6003), .A2(n5287), .ZN(n5295) );
  INV_X1 U6455 ( .A(n5584), .ZN(n5288) );
  NAND2_X1 U6456 ( .A1(n6054), .A2(n5288), .ZN(n5290) );
  NAND2_X1 U6457 ( .A1(n6779), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5289)
         );
  NAND3_X1 U6458 ( .A1(n5290), .A2(n5289), .A3(n6781), .ZN(n5293) );
  NOR2_X1 U6459 ( .A1(n6029), .A2(n5291), .ZN(n5292) );
  AOI211_X1 U6460 ( .C1(n6787), .C2(n6215), .A(n5293), .B(n5292), .ZN(n5294)
         );
  OAI211_X1 U6461 ( .C1(n5588), .C2(n6790), .A(n5295), .B(n5294), .ZN(U2819)
         );
  NAND2_X1 U6462 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6040), .ZN(n5296) );
  AOI21_X1 U6463 ( .B1(n6667), .B2(n5296), .A(n6019), .ZN(n5306) );
  OR2_X1 U6464 ( .A1(n5310), .A2(n5297), .ZN(n5298) );
  OAI21_X1 U6465 ( .B1(n6047), .B2(n3535), .A(n6781), .ZN(n5299) );
  AOI21_X1 U6466 ( .B1(n5300), .B2(n6054), .A(n5299), .ZN(n5303) );
  AOI22_X1 U6467 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6780), .B1(n6787), .B2(n5301), 
        .ZN(n5302) );
  OAI211_X1 U6468 ( .C1(n5304), .C2(n6051), .A(n5303), .B(n5302), .ZN(n5305)
         );
  OR2_X1 U6469 ( .A1(n5306), .A2(n5305), .ZN(U2822) );
  OAI21_X1 U6470 ( .B1(n5980), .B2(REIP_REG_1__SCAN_IN), .A(n5307), .ZN(n6043)
         );
  XNOR2_X1 U6471 ( .A(n4584), .B(n5308), .ZN(n6261) );
  INV_X1 U6472 ( .A(n6261), .ZN(n5311) );
  INV_X1 U6473 ( .A(n4076), .ZN(n5309) );
  OR2_X1 U6474 ( .A1(n5310), .A2(n5309), .ZN(n6045) );
  OAI22_X1 U6475 ( .A1(n5311), .A2(n6044), .B1(n6045), .B2(n4590), .ZN(n5316)
         );
  INV_X1 U6476 ( .A(n6181), .ZN(n5312) );
  AOI22_X1 U6477 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6779), .B1(n6054), 
        .B2(n5312), .ZN(n5314) );
  INV_X1 U6478 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6042) );
  NAND3_X1 U6479 ( .A1(n6775), .A2(REIP_REG_1__SCAN_IN), .A3(n6042), .ZN(n5313) );
  OAI211_X1 U6480 ( .C1(n6068), .C2(n6029), .A(n5314), .B(n5313), .ZN(n5315)
         );
  AOI211_X1 U6481 ( .C1(REIP_REG_2__SCAN_IN), .C2(n6043), .A(n5316), .B(n5315), 
        .ZN(n5317) );
  OAI21_X1 U6482 ( .B1(n5318), .B2(n6051), .A(n5317), .ZN(U2825) );
  AOI22_X1 U6483 ( .A1(EBX_REG_1__SCAN_IN), .A2(n6780), .B1(n3017), .B2(
        REIP_REG_1__SCAN_IN), .ZN(n5324) );
  INV_X1 U6484 ( .A(n4548), .ZN(n5319) );
  OAI22_X1 U6485 ( .A1(n5319), .A2(n6044), .B1(n6045), .B2(n5759), .ZN(n5322)
         );
  OAI22_X1 U6486 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n6778), .B1(n6047), 
        .B2(n5320), .ZN(n5321) );
  AOI211_X1 U6487 ( .C1(n6775), .C2(n6589), .A(n5322), .B(n5321), .ZN(n5323)
         );
  OAI211_X1 U6488 ( .C1(n6051), .C2(n5325), .A(n5324), .B(n5323), .ZN(U2826)
         );
  OAI22_X1 U6489 ( .A1(n5327), .A2(n6029), .B1(n6044), .B2(n5326), .ZN(n5330)
         );
  OAI21_X1 U6490 ( .B1(n6779), .B2(n6054), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5328) );
  OAI21_X1 U6491 ( .B1(n6045), .B2(n6313), .A(n5328), .ZN(n5329) );
  AOI211_X1 U6492 ( .C1(REIP_REG_0__SCAN_IN), .C2(n6030), .A(n5330), .B(n5329), 
        .ZN(n5331) );
  OAI21_X1 U6493 ( .B1(n6051), .B2(n5332), .A(n5331), .ZN(U2827) );
  OAI222_X1 U6494 ( .A1(n5371), .A2(n5441), .B1(n5333), .B2(n6067), .C1(n5599), 
        .C2(n5369), .ZN(U2830) );
  OAI222_X1 U6495 ( .A1(n5371), .A2(n5382), .B1(n5334), .B2(n6067), .C1(n5610), 
        .C2(n5369), .ZN(U2831) );
  AOI22_X1 U6496 ( .A1(n5619), .A2(n6065), .B1(EBX_REG_27__SCAN_IN), .B2(n5337), .ZN(n5335) );
  OAI21_X1 U6497 ( .B1(n5456), .B2(n5371), .A(n5335), .ZN(U2832) );
  AOI22_X1 U6498 ( .A1(n5636), .A2(n6065), .B1(EBX_REG_25__SCAN_IN), .B2(n5337), .ZN(n5336) );
  OAI21_X1 U6499 ( .B1(n5390), .B2(n5371), .A(n5336), .ZN(U2834) );
  INV_X1 U6500 ( .A(n5484), .ZN(n5393) );
  AOI22_X1 U6501 ( .A1(n5338), .A2(n6065), .B1(EBX_REG_24__SCAN_IN), .B2(n5337), .ZN(n5339) );
  OAI21_X1 U6502 ( .B1(n5393), .B2(n5371), .A(n5339), .ZN(U2835) );
  INV_X1 U6503 ( .A(n5496), .ZN(n5396) );
  OAI222_X1 U6504 ( .A1(n5371), .A2(n5396), .B1(n5340), .B2(n6067), .C1(n5647), 
        .C2(n5369), .ZN(U2836) );
  INV_X1 U6505 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5341) );
  OAI222_X1 U6506 ( .A1(n5371), .A2(n5399), .B1(n5341), .B2(n6067), .C1(n5654), 
        .C2(n5369), .ZN(U2837) );
  INV_X1 U6507 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5342) );
  OAI222_X1 U6508 ( .A1(n5371), .A2(n5208), .B1(n5342), .B2(n6067), .C1(n5671), 
        .C2(n5369), .ZN(U2839) );
  INV_X1 U6509 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6651) );
  OAI222_X1 U6510 ( .A1(n5407), .A2(n5371), .B1(n6067), .B2(n6651), .C1(n5369), 
        .C2(n5685), .ZN(U2840) );
  OAI222_X1 U6511 ( .A1(n5371), .A2(n5518), .B1(n5343), .B2(n6067), .C1(n5694), 
        .C2(n5369), .ZN(U2841) );
  OAI22_X1 U6512 ( .A1(n5703), .A2(n5369), .B1(n5344), .B2(n6067), .ZN(n5345)
         );
  AOI21_X1 U6513 ( .B1(n6069), .B2(n4264), .A(n5345), .ZN(n5346) );
  INV_X1 U6514 ( .A(n5346), .ZN(U2842) );
  OR2_X1 U6515 ( .A1(n5259), .A2(n5347), .ZN(n5348) );
  AND2_X1 U6516 ( .A1(n3940), .A2(n5348), .ZN(n6074) );
  INV_X1 U6517 ( .A(n6074), .ZN(n5352) );
  INV_X1 U6518 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5351) );
  AND2_X1 U6519 ( .A1(n5261), .A2(n5349), .ZN(n5350) );
  OR2_X1 U6520 ( .A1(n5350), .A2(n5247), .ZN(n5957) );
  OAI222_X1 U6521 ( .A1(n5371), .A2(n5352), .B1(n5351), .B2(n6067), .C1(n5957), 
        .C2(n5369), .ZN(U2843) );
  NOR2_X1 U6522 ( .A1(n6067), .A2(n5353), .ZN(n5354) );
  AOI21_X1 U6523 ( .B1(n5726), .B2(n6065), .A(n5354), .ZN(n5355) );
  OAI21_X1 U6524 ( .B1(n5411), .B2(n5371), .A(n5355), .ZN(U2844) );
  OR2_X1 U6525 ( .A1(n5357), .A2(n5356), .ZN(n5358) );
  AND2_X1 U6526 ( .A1(n5258), .A2(n5358), .ZN(n5971) );
  INV_X1 U6527 ( .A(n5971), .ZN(n5413) );
  INV_X1 U6528 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6692) );
  OR2_X1 U6529 ( .A1(n5359), .A2(n5360), .ZN(n5361) );
  NAND2_X1 U6530 ( .A1(n5362), .A2(n5361), .ZN(n5967) );
  OAI222_X1 U6531 ( .A1(n5413), .A2(n5371), .B1(n6067), .B2(n6692), .C1(n5967), 
        .C2(n5369), .ZN(U2845) );
  INV_X1 U6532 ( .A(n5987), .ZN(n5365) );
  OAI21_X1 U6533 ( .B1(n5365), .B2(n5364), .A(n5916), .ZN(n6772) );
  INV_X1 U6534 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5368) );
  XOR2_X1 U6535 ( .A(n5367), .B(n5366), .Z(n5559) );
  INV_X1 U6536 ( .A(n5559), .ZN(n6791) );
  OAI222_X1 U6537 ( .A1(n5369), .A2(n6772), .B1(n6067), .B2(n5368), .C1(n5371), 
        .C2(n6791), .ZN(U2847) );
  INV_X1 U6538 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5370) );
  OAI222_X1 U6539 ( .A1(n5425), .A2(n5371), .B1(n6067), .B2(n5370), .C1(n6197), 
        .C2(n5369), .ZN(U2849) );
  AOI22_X1 U6540 ( .A1(n6072), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6075), .ZN(n5376) );
  NOR3_X1 U6541 ( .A1(n6075), .A2(n5373), .A3(n5372), .ZN(n5374) );
  NAND2_X1 U6542 ( .A1(n6076), .A2(DATAI_14_), .ZN(n5375) );
  OAI211_X1 U6543 ( .C1(n5377), .C2(n5424), .A(n5376), .B(n5375), .ZN(U2861)
         );
  AOI22_X1 U6544 ( .A1(n6072), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6075), .ZN(n5379) );
  NAND2_X1 U6545 ( .A1(n6076), .A2(DATAI_13_), .ZN(n5378) );
  OAI211_X1 U6546 ( .C1(n5441), .C2(n5424), .A(n5379), .B(n5378), .ZN(U2862)
         );
  AOI22_X1 U6547 ( .A1(n6072), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6075), .ZN(n5381) );
  NAND2_X1 U6548 ( .A1(n6076), .A2(DATAI_12_), .ZN(n5380) );
  OAI211_X1 U6549 ( .C1(n5382), .C2(n5424), .A(n5381), .B(n5380), .ZN(U2863)
         );
  AOI22_X1 U6550 ( .A1(n6072), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6075), .ZN(n5384) );
  NAND2_X1 U6551 ( .A1(n6076), .A2(DATAI_11_), .ZN(n5383) );
  OAI211_X1 U6552 ( .C1(n5456), .C2(n5424), .A(n5384), .B(n5383), .ZN(U2864)
         );
  AOI22_X1 U6553 ( .A1(n6072), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6075), .ZN(n5386) );
  NAND2_X1 U6554 ( .A1(n6076), .A2(DATAI_10_), .ZN(n5385) );
  OAI211_X1 U6555 ( .C1(n5387), .C2(n5424), .A(n5386), .B(n5385), .ZN(U2865)
         );
  AOI22_X1 U6556 ( .A1(n6072), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6075), .ZN(n5389) );
  NAND2_X1 U6557 ( .A1(n6076), .A2(DATAI_9_), .ZN(n5388) );
  OAI211_X1 U6558 ( .C1(n5390), .C2(n5424), .A(n5389), .B(n5388), .ZN(U2866)
         );
  AOI22_X1 U6559 ( .A1(n6072), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6075), .ZN(n5392) );
  NAND2_X1 U6560 ( .A1(n6076), .A2(DATAI_8_), .ZN(n5391) );
  OAI211_X1 U6561 ( .C1(n5393), .C2(n5424), .A(n5392), .B(n5391), .ZN(U2867)
         );
  AOI22_X1 U6562 ( .A1(n6072), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6075), .ZN(n5395) );
  NAND2_X1 U6563 ( .A1(n6076), .A2(DATAI_7_), .ZN(n5394) );
  OAI211_X1 U6564 ( .C1(n5396), .C2(n5424), .A(n5395), .B(n5394), .ZN(U2868)
         );
  AOI22_X1 U6565 ( .A1(n6072), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n6075), .ZN(n5398) );
  NAND2_X1 U6566 ( .A1(n6076), .A2(DATAI_6_), .ZN(n5397) );
  OAI211_X1 U6567 ( .C1(n5399), .C2(n5424), .A(n5398), .B(n5397), .ZN(U2869)
         );
  AOI22_X1 U6568 ( .A1(n6072), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n6075), .ZN(n5401) );
  NAND2_X1 U6569 ( .A1(n6076), .A2(DATAI_5_), .ZN(n5400) );
  OAI211_X1 U6570 ( .C1(n5402), .C2(n5424), .A(n5401), .B(n5400), .ZN(U2870)
         );
  AOI22_X1 U6571 ( .A1(n6072), .A2(DATAI_20_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n6075), .ZN(n5404) );
  NAND2_X1 U6572 ( .A1(n6076), .A2(DATAI_4_), .ZN(n5403) );
  OAI211_X1 U6573 ( .C1(n5208), .C2(n5424), .A(n5404), .B(n5403), .ZN(U2871)
         );
  AOI22_X1 U6574 ( .A1(n6072), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6075), .ZN(n5406) );
  NAND2_X1 U6575 ( .A1(n6076), .A2(DATAI_3_), .ZN(n5405) );
  OAI211_X1 U6576 ( .C1(n5407), .C2(n5424), .A(n5406), .B(n5405), .ZN(U2872)
         );
  AOI22_X1 U6577 ( .A1(n6072), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n6075), .ZN(n5409) );
  NAND2_X1 U6578 ( .A1(n6076), .A2(DATAI_2_), .ZN(n5408) );
  OAI211_X1 U6579 ( .C1(n5518), .C2(n5424), .A(n5409), .B(n5408), .ZN(U2873)
         );
  AOI22_X1 U6580 ( .A1(n5422), .A2(DATAI_15_), .B1(n6075), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5410) );
  OAI21_X1 U6581 ( .B1(n5411), .B2(n5424), .A(n5410), .ZN(U2876) );
  AOI22_X1 U6582 ( .A1(n5422), .A2(DATAI_14_), .B1(n6075), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5412) );
  OAI21_X1 U6583 ( .B1(n5413), .B2(n5424), .A(n5412), .ZN(U2877) );
  INV_X1 U6584 ( .A(DATAI_13_), .ZN(n6124) );
  INV_X1 U6585 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6641) );
  OAI222_X1 U6586 ( .A1(n5417), .A2(n6124), .B1(n5416), .B2(n6641), .C1(n5424), 
        .C2(n5911), .ZN(U2878) );
  AOI22_X1 U6587 ( .A1(n5422), .A2(DATAI_12_), .B1(n6075), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5418) );
  OAI21_X1 U6588 ( .B1(n6791), .B2(n5424), .A(n5418), .ZN(U2879) );
  AOI21_X1 U6589 ( .B1(n5419), .B2(n5269), .A(n5366), .ZN(n6151) );
  INV_X1 U6590 ( .A(n6151), .ZN(n5421) );
  AOI22_X1 U6591 ( .A1(n5422), .A2(DATAI_11_), .B1(n6075), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5420) );
  OAI21_X1 U6592 ( .B1(n5421), .B2(n5424), .A(n5420), .ZN(U2880) );
  AOI22_X1 U6593 ( .A1(n5422), .A2(DATAI_10_), .B1(n6075), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5423) );
  OAI21_X1 U6594 ( .B1(n5425), .B2(n5424), .A(n5423), .ZN(U2881) );
  XNOR2_X1 U6595 ( .A(n5428), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5598)
         );
  AND2_X1 U6596 ( .A1(n6233), .A2(REIP_REG_30__SCAN_IN), .ZN(n5590) );
  AOI21_X1 U6597 ( .B1(n5565), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5590), 
        .ZN(n5429) );
  OAI21_X1 U6598 ( .B1(n6182), .B2(n5430), .A(n5429), .ZN(n5431) );
  AOI21_X1 U6599 ( .B1(n5432), .B2(n6177), .A(n5431), .ZN(n5433) );
  OAI21_X1 U6600 ( .B1(n5598), .B2(n6159), .A(n5433), .ZN(U2956) );
  OAI21_X1 U6601 ( .B1(n5434), .B2(n5435), .A(n5446), .ZN(n5436) );
  XNOR2_X1 U6602 ( .A(n5436), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5607)
         );
  AND2_X1 U6603 ( .A1(n6233), .A2(REIP_REG_29__SCAN_IN), .ZN(n5600) );
  AOI21_X1 U6604 ( .B1(n5565), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5600), 
        .ZN(n5437) );
  OAI21_X1 U6605 ( .B1(n6182), .B2(n5438), .A(n5437), .ZN(n5439) );
  INV_X1 U6606 ( .A(n5439), .ZN(n5440) );
  INV_X1 U6607 ( .A(n5442), .ZN(n5443) );
  OAI21_X1 U6608 ( .B1(n5607), .B2(n6159), .A(n5443), .ZN(U2957) );
  NAND2_X1 U6609 ( .A1(n5444), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5447) );
  NAND3_X1 U6610 ( .A1(n5454), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n6756), .ZN(n5445) );
  OAI211_X1 U6611 ( .C1(n5434), .C2(n5447), .A(n5446), .B(n5445), .ZN(n5448)
         );
  AND2_X1 U6612 ( .A1(n6233), .A2(REIP_REG_28__SCAN_IN), .ZN(n5608) );
  AOI21_X1 U6613 ( .B1(n5565), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5608), 
        .ZN(n5449) );
  OAI21_X1 U6614 ( .B1(n6182), .B2(n5450), .A(n5449), .ZN(n5451) );
  AOI21_X1 U6615 ( .B1(n5452), .B2(n6177), .A(n5451), .ZN(n5453) );
  OAI21_X1 U6616 ( .B1(n5617), .B2(n6159), .A(n5453), .ZN(U2958) );
  NAND2_X1 U6617 ( .A1(n5434), .A2(n5454), .ZN(n5455) );
  XNOR2_X1 U6618 ( .A(n5455), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5625)
         );
  INV_X1 U6619 ( .A(n5456), .ZN(n5460) );
  AND2_X1 U6620 ( .A1(n6233), .A2(REIP_REG_27__SCAN_IN), .ZN(n5618) );
  AOI21_X1 U6621 ( .B1(n5565), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5618), 
        .ZN(n5457) );
  OAI21_X1 U6622 ( .B1(n6182), .B2(n5458), .A(n5457), .ZN(n5459) );
  AOI21_X1 U6623 ( .B1(n5460), .B2(n6177), .A(n5459), .ZN(n5461) );
  OAI21_X1 U6624 ( .B1(n5625), .B2(n6159), .A(n5461), .ZN(U2959) );
  NAND2_X1 U6625 ( .A1(n4186), .A2(n5463), .ZN(n5465) );
  XOR2_X1 U6626 ( .A(n5465), .B(n5464), .Z(n5633) );
  AND2_X1 U6627 ( .A1(n6233), .A2(REIP_REG_26__SCAN_IN), .ZN(n5628) );
  AOI21_X1 U6628 ( .B1(n5565), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5628), 
        .ZN(n5466) );
  OAI21_X1 U6629 ( .B1(n6182), .B2(n5467), .A(n5466), .ZN(n5468) );
  AOI21_X1 U6630 ( .B1(n5469), .B2(n6177), .A(n5468), .ZN(n5470) );
  OAI21_X1 U6631 ( .B1(n5633), .B2(n6159), .A(n5470), .ZN(U2960) );
  OAI21_X1 U6632 ( .B1(n5473), .B2(n5471), .A(n5472), .ZN(n5474) );
  INV_X1 U6633 ( .A(n5474), .ZN(n5643) );
  AND2_X1 U6634 ( .A1(n6233), .A2(REIP_REG_25__SCAN_IN), .ZN(n5635) );
  AOI21_X1 U6635 ( .B1(n5565), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5635), 
        .ZN(n5475) );
  OAI21_X1 U6636 ( .B1(n6182), .B2(n5476), .A(n5475), .ZN(n5477) );
  AOI21_X1 U6637 ( .B1(n5478), .B2(n6177), .A(n5477), .ZN(n5479) );
  OAI21_X1 U6638 ( .B1(n5643), .B2(n6159), .A(n5479), .ZN(U2961) );
  AOI21_X1 U6639 ( .B1(n5565), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5480), 
        .ZN(n5481) );
  OAI21_X1 U6640 ( .B1(n6182), .B2(n5482), .A(n5481), .ZN(n5483) );
  AOI21_X1 U6641 ( .B1(n5484), .B2(n6177), .A(n5483), .ZN(n5485) );
  OAI21_X1 U6642 ( .B1(n5486), .B2(n6159), .A(n5485), .ZN(U2962) );
  NOR2_X1 U6643 ( .A1(n5533), .A2(n5731), .ZN(n5488) );
  OAI22_X2 U6644 ( .A1(n5487), .A2(n5488), .B1(n3933), .B2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U6645 ( .A1(n6146), .A2(n5721), .ZN(n5532) );
  NAND4_X1 U6646 ( .A1(n5532), .A2(n5490), .A3(n5489), .A4(n6146), .ZN(n5491)
         );
  XNOR2_X1 U6647 ( .A(n5492), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5652)
         );
  NAND2_X1 U6648 ( .A1(n6233), .A2(REIP_REG_23__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U6649 ( .A1(n5565), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5493)
         );
  OAI211_X1 U6650 ( .C1(n6182), .C2(n5494), .A(n5646), .B(n5493), .ZN(n5495)
         );
  AOI21_X1 U6651 ( .B1(n5496), .B2(n6177), .A(n5495), .ZN(n5497) );
  OAI21_X1 U6652 ( .B1(n5652), .B2(n6159), .A(n5497), .ZN(U2963) );
  AOI21_X1 U6653 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5533), .A(n5498), 
        .ZN(n5499) );
  XNOR2_X1 U6654 ( .A(n5500), .B(n5499), .ZN(n5662) );
  AND2_X1 U6655 ( .A1(n6233), .A2(REIP_REG_22__SCAN_IN), .ZN(n5656) );
  AOI21_X1 U6656 ( .B1(n5565), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5656), 
        .ZN(n5501) );
  OAI21_X1 U6657 ( .B1(n6182), .B2(n5502), .A(n5501), .ZN(n5503) );
  AOI21_X1 U6658 ( .B1(n5504), .B2(n6177), .A(n5503), .ZN(n5505) );
  OAI21_X1 U6659 ( .B1(n5662), .B2(n6159), .A(n5505), .ZN(U2964) );
  OAI21_X1 U6660 ( .B1(n5508), .B2(n5507), .A(n5506), .ZN(n5509) );
  INV_X1 U6661 ( .A(n5509), .ZN(n5670) );
  INV_X1 U6662 ( .A(n5510), .ZN(n5512) );
  AND2_X1 U6663 ( .A1(n6233), .A2(REIP_REG_21__SCAN_IN), .ZN(n5665) );
  AOI21_X1 U6664 ( .B1(n5565), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5665), 
        .ZN(n5511) );
  OAI21_X1 U6665 ( .B1(n6182), .B2(n5512), .A(n5511), .ZN(n5513) );
  AOI21_X1 U6666 ( .B1(n5514), .B2(n6177), .A(n5513), .ZN(n5515) );
  OAI21_X1 U6667 ( .B1(n5670), .B2(n6159), .A(n5515), .ZN(U2965) );
  NAND3_X1 U6668 ( .A1(n5535), .A2(n3933), .A3(n5721), .ZN(n5524) );
  NAND3_X1 U6669 ( .A1(n5532), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5533), .ZN(n5516) );
  OAI22_X1 U6670 ( .A1(n5524), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .B1(n5516), .B2(n5535), .ZN(n5517) );
  XNOR2_X1 U6671 ( .A(n5517), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5702)
         );
  INV_X1 U6672 ( .A(n5518), .ZN(n5522) );
  AND2_X1 U6673 ( .A1(n6233), .A2(REIP_REG_18__SCAN_IN), .ZN(n5697) );
  AOI21_X1 U6674 ( .B1(n5565), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5697), 
        .ZN(n5519) );
  OAI21_X1 U6675 ( .B1(n6182), .B2(n5520), .A(n5519), .ZN(n5521) );
  AOI21_X1 U6676 ( .B1(n5522), .B2(n6177), .A(n5521), .ZN(n5523) );
  OAI21_X1 U6677 ( .B1(n5702), .B2(n6159), .A(n5523), .ZN(U2968) );
  NAND2_X1 U6678 ( .A1(n5533), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5525) );
  OAI21_X1 U6679 ( .B1(n5535), .B2(n5525), .A(n5524), .ZN(n5526) );
  XNOR2_X1 U6680 ( .A(n5526), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5711)
         );
  INV_X1 U6681 ( .A(n5527), .ZN(n5529) );
  AND2_X1 U6682 ( .A1(n6233), .A2(REIP_REG_17__SCAN_IN), .ZN(n5704) );
  AOI21_X1 U6683 ( .B1(n5565), .B2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n5704), 
        .ZN(n5528) );
  OAI21_X1 U6684 ( .B1(n6182), .B2(n5529), .A(n5528), .ZN(n5530) );
  AOI21_X1 U6685 ( .B1(n6069), .B2(n6177), .A(n5530), .ZN(n5531) );
  OAI21_X1 U6686 ( .B1(n5711), .B2(n6159), .A(n5531), .ZN(U2969) );
  OAI21_X1 U6687 ( .B1(n5721), .B2(n5533), .A(n5532), .ZN(n5534) );
  XNOR2_X1 U6688 ( .A(n5535), .B(n5534), .ZN(n5725) );
  INV_X1 U6689 ( .A(n5955), .ZN(n5537) );
  AND2_X1 U6690 ( .A1(n6233), .A2(REIP_REG_16__SCAN_IN), .ZN(n5720) );
  AOI21_X1 U6691 ( .B1(n5565), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5720), 
        .ZN(n5536) );
  OAI21_X1 U6692 ( .B1(n6182), .B2(n5537), .A(n5536), .ZN(n5538) );
  AOI21_X1 U6693 ( .B1(n6074), .B2(n6177), .A(n5538), .ZN(n5539) );
  OAI21_X1 U6694 ( .B1(n6159), .B2(n5725), .A(n5539), .ZN(U2970) );
  XNOR2_X1 U6695 ( .A(n6146), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5540)
         );
  XNOR2_X1 U6696 ( .A(n5487), .B(n5540), .ZN(n5735) );
  AND2_X1 U6697 ( .A1(n6233), .A2(REIP_REG_15__SCAN_IN), .ZN(n5729) );
  AOI21_X1 U6698 ( .B1(n5565), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5729), 
        .ZN(n5541) );
  OAI21_X1 U6699 ( .B1(n6182), .B2(n5542), .A(n5541), .ZN(n5543) );
  AOI21_X1 U6700 ( .B1(n5544), .B2(n6177), .A(n5543), .ZN(n5545) );
  OAI21_X1 U6701 ( .B1(n5735), .B2(n6159), .A(n5545), .ZN(U2971) );
  XNOR2_X1 U6702 ( .A(n6146), .B(n5740), .ZN(n5547) );
  XNOR2_X1 U6703 ( .A(n5546), .B(n5547), .ZN(n5748) );
  INV_X1 U6704 ( .A(n5970), .ZN(n5549) );
  AND2_X1 U6705 ( .A1(n6233), .A2(REIP_REG_14__SCAN_IN), .ZN(n5742) );
  AOI21_X1 U6706 ( .B1(n5565), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5742), 
        .ZN(n5548) );
  OAI21_X1 U6707 ( .B1(n6182), .B2(n5549), .A(n5548), .ZN(n5550) );
  AOI21_X1 U6708 ( .B1(n5971), .B2(n6177), .A(n5550), .ZN(n5551) );
  OAI21_X1 U6709 ( .B1(n6159), .B2(n5748), .A(n5551), .ZN(U2972) );
  NAND2_X1 U6710 ( .A1(n5553), .A2(n5552), .ZN(n5556) );
  XOR2_X1 U6711 ( .A(n5556), .B(n5555), .Z(n5756) );
  INV_X1 U6712 ( .A(n5756), .ZN(n5561) );
  NAND2_X1 U6713 ( .A1(n6233), .A2(REIP_REG_12__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U6714 ( .A1(n5565), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5557)
         );
  OAI211_X1 U6715 ( .C1(n6182), .C2(n6777), .A(n5752), .B(n5557), .ZN(n5558)
         );
  AOI21_X1 U6716 ( .B1(n5559), .B2(n6177), .A(n5558), .ZN(n5560) );
  OAI21_X1 U6717 ( .B1(n5561), .B2(n6159), .A(n5560), .ZN(U2974) );
  NAND2_X1 U6718 ( .A1(n3933), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5574)
         );
  NOR2_X1 U6719 ( .A1(n3933), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6144)
         );
  NAND2_X1 U6720 ( .A1(n3933), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6143) );
  INV_X1 U6721 ( .A(n6143), .ZN(n5563) );
  NOR2_X1 U6722 ( .A1(n6144), .A2(n5563), .ZN(n5564) );
  XNOR2_X1 U6723 ( .A(n6145), .B(n5564), .ZN(n6199) );
  INV_X1 U6724 ( .A(n6199), .ZN(n5571) );
  AOI22_X1 U6725 ( .A1(n5565), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6233), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5566) );
  OAI21_X1 U6726 ( .B1(n6182), .B2(n5567), .A(n5566), .ZN(n5568) );
  AOI21_X1 U6727 ( .B1(n5569), .B2(n6177), .A(n5568), .ZN(n5570) );
  OAI21_X1 U6728 ( .B1(n5571), .B2(n6159), .A(n5570), .ZN(U2976) );
  NAND2_X1 U6729 ( .A1(n5574), .A2(n5573), .ZN(n5575) );
  XNOR2_X1 U6730 ( .A(n5572), .B(n5575), .ZN(n6209) );
  NAND2_X1 U6731 ( .A1(n6209), .A2(n3910), .ZN(n5579) );
  INV_X1 U6732 ( .A(n6182), .ZN(n6150) );
  NAND2_X1 U6733 ( .A1(n6233), .A2(REIP_REG_9__SCAN_IN), .ZN(n6205) );
  OAI21_X1 U6734 ( .B1(n5576), .B2(n6001), .A(n6205), .ZN(n5577) );
  AOI21_X1 U6735 ( .B1(n6150), .B2(n5996), .A(n5577), .ZN(n5578) );
  OAI211_X1 U6736 ( .C1(n6157), .C2(n5995), .A(n5579), .B(n5578), .ZN(U2977)
         );
  OAI21_X1 U6737 ( .B1(n5580), .B2(n5582), .A(n5581), .ZN(n5583) );
  INV_X1 U6738 ( .A(n5583), .ZN(n6216) );
  NAND2_X1 U6739 ( .A1(n6216), .A2(n3910), .ZN(n5587) );
  NOR2_X1 U6740 ( .A1(n6248), .A2(n6541), .ZN(n6214) );
  NOR2_X1 U6741 ( .A1(n6182), .A2(n5584), .ZN(n5585) );
  AOI211_X1 U6742 ( .C1(n5565), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6214), 
        .B(n5585), .ZN(n5586) );
  OAI211_X1 U6743 ( .C1(n6157), .C2(n5588), .A(n5587), .B(n5586), .ZN(U2978)
         );
  NOR3_X1 U6744 ( .A1(n5603), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5589), 
        .ZN(n5595) );
  INV_X1 U6745 ( .A(n5590), .ZN(n5591) );
  OAI21_X1 U6746 ( .B1(n5593), .B2(n5592), .A(n5591), .ZN(n5594) );
  AOI211_X1 U6747 ( .C1(n5596), .C2(n6262), .A(n5595), .B(n5594), .ZN(n5597)
         );
  OAI21_X1 U6748 ( .B1(n5598), .B2(n6184), .A(n5597), .ZN(U2988) );
  INV_X1 U6749 ( .A(n5599), .ZN(n5605) );
  AOI21_X1 U6750 ( .B1(n5601), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5600), 
        .ZN(n5602) );
  OAI21_X1 U6751 ( .B1(n5603), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5602), 
        .ZN(n5604) );
  AOI21_X1 U6752 ( .B1(n5605), .B2(n6262), .A(n5604), .ZN(n5606) );
  OAI21_X1 U6753 ( .B1(n5607), .B2(n6184), .A(n5606), .ZN(U2989) );
  INV_X1 U6754 ( .A(n5621), .ZN(n5615) );
  INV_X1 U6755 ( .A(n5608), .ZN(n5609) );
  OAI21_X1 U6756 ( .B1(n5610), .B2(n6250), .A(n5609), .ZN(n5614) );
  INV_X1 U6757 ( .A(n5623), .ZN(n5612) );
  NOR3_X1 U6758 ( .A1(n5612), .A2(n3001), .A3(n5611), .ZN(n5613) );
  AOI211_X1 U6759 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5615), .A(n5614), .B(n5613), .ZN(n5616) );
  OAI21_X1 U6760 ( .B1(n5617), .B2(n6184), .A(n5616), .ZN(U2990) );
  AOI21_X1 U6761 ( .B1(n5619), .B2(n6262), .A(n5618), .ZN(n5620) );
  OAI21_X1 U6762 ( .B1(n5621), .B2(n6756), .A(n5620), .ZN(n5622) );
  AOI21_X1 U6763 ( .B1(n5623), .B2(n6756), .A(n5622), .ZN(n5624) );
  OAI21_X1 U6764 ( .B1(n5625), .B2(n6184), .A(n5624), .ZN(U2991) );
  NOR2_X1 U6765 ( .A1(n5626), .A2(n6250), .ZN(n5627) );
  AOI211_X1 U6766 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5634), .A(n5628), .B(n5627), .ZN(n5632) );
  INV_X1 U6767 ( .A(n5629), .ZN(n5641) );
  OAI211_X1 U6768 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5641), .B(n5630), .ZN(n5631) );
  OAI211_X1 U6769 ( .C1(n5633), .C2(n6184), .A(n5632), .B(n5631), .ZN(U2992)
         );
  INV_X1 U6770 ( .A(n5634), .ZN(n5638) );
  AOI21_X1 U6771 ( .B1(n5636), .B2(n6262), .A(n5635), .ZN(n5637) );
  OAI21_X1 U6772 ( .B1(n5638), .B2(n5640), .A(n5637), .ZN(n5639) );
  AOI21_X1 U6773 ( .B1(n5641), .B2(n5640), .A(n5639), .ZN(n5642) );
  OAI21_X1 U6774 ( .B1(n5643), .B2(n6184), .A(n5642), .ZN(U2993) );
  INV_X1 U6775 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U6776 ( .A1(n5644), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5645) );
  OAI211_X1 U6777 ( .C1(n5647), .C2(n6250), .A(n5646), .B(n5645), .ZN(n5648)
         );
  AOI21_X1 U6778 ( .B1(n5650), .B2(n5649), .A(n5648), .ZN(n5651) );
  OAI21_X1 U6779 ( .B1(n5652), .B2(n6184), .A(n5651), .ZN(U2995) );
  INV_X1 U6780 ( .A(n5653), .ZN(n5666) );
  NOR2_X1 U6781 ( .A1(n5654), .A2(n6250), .ZN(n5655) );
  AOI211_X1 U6782 ( .C1(n5666), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5656), .B(n5655), .ZN(n5661) );
  INV_X1 U6783 ( .A(n5657), .ZN(n5658) );
  NAND3_X1 U6784 ( .A1(n5667), .A2(n5659), .A3(n5658), .ZN(n5660) );
  OAI211_X1 U6785 ( .C1(n5662), .C2(n6184), .A(n5661), .B(n5660), .ZN(U2996)
         );
  NOR2_X1 U6786 ( .A1(n5663), .A2(n6250), .ZN(n5664) );
  AOI211_X1 U6787 ( .C1(n5666), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5665), .B(n5664), .ZN(n5669) );
  INV_X1 U6788 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6707) );
  NAND2_X1 U6789 ( .A1(n5667), .A2(n6707), .ZN(n5668) );
  OAI211_X1 U6790 ( .C1(n5670), .C2(n6184), .A(n5669), .B(n5668), .ZN(U2997)
         );
  INV_X1 U6791 ( .A(n5671), .ZN(n5677) );
  INV_X1 U6792 ( .A(n5695), .ZN(n5706) );
  NAND2_X1 U6793 ( .A1(n5706), .A2(n5672), .ZN(n5689) );
  NOR3_X1 U6794 ( .A1(n5689), .A2(n5674), .A3(n5673), .ZN(n5675) );
  AOI211_X1 U6795 ( .C1(n6262), .C2(n5677), .A(n5676), .B(n5675), .ZN(n5683)
         );
  AOI21_X1 U6796 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5678), .A(n5712), 
        .ZN(n5679) );
  AOI21_X1 U6797 ( .B1(n6193), .B2(n5680), .A(n5679), .ZN(n5708) );
  OAI21_X1 U6798 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6268), .A(n5708), 
        .ZN(n5699) );
  INV_X1 U6799 ( .A(n5699), .ZN(n5681) );
  OAI21_X1 U6800 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5718), .A(n5681), 
        .ZN(n5691) );
  NAND2_X1 U6801 ( .A1(n5691), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5682) );
  OAI211_X1 U6802 ( .C1(n5684), .C2(n6184), .A(n5683), .B(n5682), .ZN(U2998)
         );
  INV_X1 U6803 ( .A(n5685), .ZN(n5687) );
  AOI21_X1 U6804 ( .B1(n5687), .B2(n6262), .A(n5686), .ZN(n5688) );
  OAI21_X1 U6805 ( .B1(n5689), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5688), 
        .ZN(n5690) );
  AOI21_X1 U6806 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5691), .A(n5690), 
        .ZN(n5692) );
  OAI21_X1 U6807 ( .B1(n5693), .B2(n6184), .A(n5692), .ZN(U2999) );
  INV_X1 U6808 ( .A(n5694), .ZN(n5698) );
  NOR3_X1 U6809 ( .A1(n5695), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n5707), 
        .ZN(n5696) );
  AOI211_X1 U6810 ( .C1(n6262), .C2(n5698), .A(n5697), .B(n5696), .ZN(n5701)
         );
  NAND2_X1 U6811 ( .A1(n5699), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5700) );
  OAI211_X1 U6812 ( .C1(n5702), .C2(n6184), .A(n5701), .B(n5700), .ZN(U3000)
         );
  NOR2_X1 U6813 ( .A1(n5703), .A2(n6250), .ZN(n5705) );
  AOI211_X1 U6814 ( .C1(n5706), .C2(n5707), .A(n5705), .B(n5704), .ZN(n5710)
         );
  OR2_X1 U6815 ( .A1(n5708), .A2(n5707), .ZN(n5709) );
  OAI211_X1 U6816 ( .C1(n5711), .C2(n6184), .A(n5710), .B(n5709), .ZN(U3001)
         );
  OR2_X1 U6817 ( .A1(n5713), .A2(n5712), .ZN(n5716) );
  NAND2_X1 U6818 ( .A1(n6193), .A2(n5714), .ZN(n5715) );
  NAND2_X1 U6819 ( .A1(n5716), .A2(n5715), .ZN(n6188) );
  INV_X1 U6820 ( .A(n6188), .ZN(n5750) );
  OAI21_X1 U6821 ( .B1(n5718), .B2(n5717), .A(n5750), .ZN(n5730) );
  NOR2_X1 U6822 ( .A1(n5957), .A2(n6250), .ZN(n5719) );
  AOI211_X1 U6823 ( .C1(n5730), .C2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5720), .B(n5719), .ZN(n5724) );
  XNOR2_X1 U6824 ( .A(n5721), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5722)
         );
  NAND2_X1 U6825 ( .A1(n5732), .A2(n5722), .ZN(n5723) );
  OAI211_X1 U6826 ( .C1(n5725), .C2(n6184), .A(n5724), .B(n5723), .ZN(U3002)
         );
  INV_X1 U6827 ( .A(n5726), .ZN(n5727) );
  NOR2_X1 U6828 ( .A1(n5727), .A2(n6250), .ZN(n5728) );
  AOI211_X1 U6829 ( .C1(n5730), .C2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5729), .B(n5728), .ZN(n5734) );
  NAND2_X1 U6830 ( .A1(n5732), .A2(n5731), .ZN(n5733) );
  OAI211_X1 U6831 ( .C1(n5735), .C2(n6184), .A(n5734), .B(n5733), .ZN(U3003)
         );
  NAND2_X1 U6832 ( .A1(n5924), .A2(n5736), .ZN(n5918) );
  OAI22_X1 U6833 ( .A1(n5738), .A2(n5741), .B1(n5737), .B2(n5736), .ZN(n5739)
         );
  NOR2_X1 U6834 ( .A1(n6188), .A2(n5739), .ZN(n5925) );
  OAI21_X1 U6835 ( .B1(n2974), .B2(n5918), .A(n5925), .ZN(n5746) );
  NAND3_X1 U6836 ( .A1(n5919), .A2(n5741), .A3(n5740), .ZN(n5744) );
  INV_X1 U6837 ( .A(n5742), .ZN(n5743) );
  OAI211_X1 U6838 ( .C1(n6250), .C2(n5967), .A(n5744), .B(n5743), .ZN(n5745)
         );
  AOI21_X1 U6839 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n5746), .A(n5745), 
        .ZN(n5747) );
  OAI21_X1 U6840 ( .B1(n5748), .B2(n6184), .A(n5747), .ZN(U3004) );
  INV_X1 U6841 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5749) );
  NAND2_X1 U6842 ( .A1(n5749), .A2(n5919), .ZN(n6189) );
  AOI21_X1 U6843 ( .B1(n5750), .B2(n6189), .A(n5751), .ZN(n5755) );
  NAND3_X1 U6844 ( .A1(n5919), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n5751), .ZN(n5753) );
  OAI211_X1 U6845 ( .C1(n6250), .C2(n6772), .A(n5753), .B(n5752), .ZN(n5754)
         );
  AOI211_X1 U6846 ( .C1(n5756), .C2(n6266), .A(n5755), .B(n5754), .ZN(n5757)
         );
  INV_X1 U6847 ( .A(n5757), .ZN(U3006) );
  INV_X1 U6848 ( .A(n6310), .ZN(n6402) );
  OAI211_X1 U6849 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n2964), .A(n6402), .B(
        n6401), .ZN(n5758) );
  OAI21_X1 U6850 ( .B1(n5761), .B2(n5759), .A(n5758), .ZN(n5760) );
  MUX2_X1 U6851 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5760), .S(n6274), 
        .Z(U3464) );
  XNOR2_X1 U6852 ( .A(n6402), .B(n4633), .ZN(n5762) );
  OAI22_X1 U6853 ( .A1(n5762), .A2(n6406), .B1(n4590), .B2(n5761), .ZN(n5763)
         );
  MUX2_X1 U6854 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5763), .S(n6274), 
        .Z(U3463) );
  OAI22_X1 U6855 ( .A1(n5765), .A2(n5926), .B1(n5764), .B2(n6502), .ZN(n5766)
         );
  MUX2_X1 U6856 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5766), .S(n5930), 
        .Z(U3456) );
  NAND3_X1 U6857 ( .A1(n4633), .A2(n5767), .A3(n2964), .ZN(n5768) );
  NOR2_X1 U6858 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5769), .ZN(n5782)
         );
  INV_X1 U6859 ( .A(n5782), .ZN(n5816) );
  INV_X1 U6860 ( .A(n5770), .ZN(n5772) );
  INV_X1 U6861 ( .A(n5869), .ZN(n5771) );
  OAI22_X1 U6862 ( .A1(n5774), .A2(n5773), .B1(n5772), .B2(n5771), .ZN(n5814)
         );
  AOI21_X1 U6863 ( .B1(n6339), .B2(n5775), .A(n6604), .ZN(n5776) );
  AOI211_X1 U6864 ( .C1(n5778), .C2(n5777), .A(n5776), .B(n6406), .ZN(n5780)
         );
  NOR3_X1 U6865 ( .A1(n6279), .A2(n5780), .A3(n5779), .ZN(n5781) );
  AOI22_X1 U6866 ( .A1(n5814), .A2(n6413), .B1(INSTQUEUE_REG_4__0__SCAN_IN), 
        .B2(n5813), .ZN(n5783) );
  OAI21_X1 U6867 ( .B1(n5784), .B2(n5816), .A(n5783), .ZN(n5785) );
  AOI21_X1 U6868 ( .B1(n6400), .B2(n5819), .A(n5785), .ZN(n5786) );
  OAI21_X1 U6869 ( .B1(n6416), .B2(n6339), .A(n5786), .ZN(U3052) );
  AOI22_X1 U6870 ( .A1(n5814), .A2(n6419), .B1(INSTQUEUE_REG_4__1__SCAN_IN), 
        .B2(n5813), .ZN(n5787) );
  OAI21_X1 U6871 ( .B1(n5788), .B2(n5816), .A(n5787), .ZN(n5789) );
  AOI21_X1 U6872 ( .B1(n6418), .B2(n5819), .A(n5789), .ZN(n5790) );
  OAI21_X1 U6873 ( .B1(n6422), .B2(n6339), .A(n5790), .ZN(U3053) );
  AOI22_X1 U6874 ( .A1(n5814), .A2(n6425), .B1(INSTQUEUE_REG_4__2__SCAN_IN), 
        .B2(n5813), .ZN(n5791) );
  OAI21_X1 U6875 ( .B1(n5792), .B2(n5816), .A(n5791), .ZN(n5793) );
  AOI21_X1 U6876 ( .B1(n6424), .B2(n5819), .A(n5793), .ZN(n5794) );
  OAI21_X1 U6877 ( .B1(n6428), .B2(n6339), .A(n5794), .ZN(U3054) );
  AOI22_X1 U6878 ( .A1(n5814), .A2(n6431), .B1(INSTQUEUE_REG_4__3__SCAN_IN), 
        .B2(n5813), .ZN(n5795) );
  OAI21_X1 U6879 ( .B1(n5796), .B2(n5816), .A(n5795), .ZN(n5797) );
  AOI21_X1 U6880 ( .B1(n5798), .B2(n5819), .A(n5797), .ZN(n5799) );
  OAI21_X1 U6881 ( .B1(n5842), .B2(n6339), .A(n5799), .ZN(U3055) );
  AOI22_X1 U6882 ( .A1(n5814), .A2(n6437), .B1(INSTQUEUE_REG_4__4__SCAN_IN), 
        .B2(n5813), .ZN(n5800) );
  OAI21_X1 U6883 ( .B1(n5801), .B2(n5816), .A(n5800), .ZN(n5802) );
  AOI21_X1 U6884 ( .B1(n6436), .B2(n5819), .A(n5802), .ZN(n5803) );
  OAI21_X1 U6885 ( .B1(n6440), .B2(n6339), .A(n5803), .ZN(U3056) );
  AOI22_X1 U6886 ( .A1(n5814), .A2(n6443), .B1(INSTQUEUE_REG_4__5__SCAN_IN), 
        .B2(n5813), .ZN(n5804) );
  OAI21_X1 U6887 ( .B1(n5805), .B2(n5816), .A(n5804), .ZN(n5806) );
  AOI21_X1 U6888 ( .B1(n5807), .B2(n5819), .A(n5806), .ZN(n5808) );
  OAI21_X1 U6889 ( .B1(n5849), .B2(n6339), .A(n5808), .ZN(U3057) );
  AOI22_X1 U6890 ( .A1(n5814), .A2(n6450), .B1(INSTQUEUE_REG_4__6__SCAN_IN), 
        .B2(n5813), .ZN(n5809) );
  OAI21_X1 U6891 ( .B1(n5810), .B2(n5816), .A(n5809), .ZN(n5811) );
  AOI21_X1 U6892 ( .B1(n6386), .B2(n5819), .A(n5811), .ZN(n5812) );
  OAI21_X1 U6893 ( .B1(n6389), .B2(n6339), .A(n5812), .ZN(U3058) );
  AOI22_X1 U6894 ( .A1(n5814), .A2(n6460), .B1(INSTQUEUE_REG_4__7__SCAN_IN), 
        .B2(n5813), .ZN(n5815) );
  OAI21_X1 U6895 ( .B1(n5817), .B2(n5816), .A(n5815), .ZN(n5818) );
  AOI21_X1 U6896 ( .B1(n6457), .B2(n5819), .A(n5818), .ZN(n5820) );
  OAI21_X1 U6897 ( .B1(n6465), .B2(n6339), .A(n5820), .ZN(U3059) );
  AOI21_X1 U6898 ( .B1(n5862), .B2(n6385), .A(n6604), .ZN(n5829) );
  OAI21_X1 U6899 ( .B1(n5823), .B2(n6278), .A(n6401), .ZN(n5828) );
  NOR2_X1 U6900 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5824), .ZN(n5859)
         );
  INV_X1 U6901 ( .A(n5859), .ZN(n5825) );
  AOI21_X1 U6902 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5825), .A(n5869), .ZN(
        n5826) );
  NAND2_X1 U6903 ( .A1(n5856), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5835) );
  AOI22_X1 U6904 ( .A1(n5832), .A2(n5831), .B1(n6279), .B2(n5830), .ZN(n5857)
         );
  OAI22_X1 U6905 ( .A1(n6385), .A2(n6416), .B1(n5857), .B2(n5878), .ZN(n5833)
         );
  AOI21_X1 U6906 ( .B1(n6399), .B2(n5859), .A(n5833), .ZN(n5834) );
  OAI211_X1 U6907 ( .C1(n6369), .C2(n5862), .A(n5835), .B(n5834), .ZN(U3084)
         );
  NAND2_X1 U6908 ( .A1(n5856), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5838) );
  OAI22_X1 U6909 ( .A1(n6385), .A2(n6422), .B1(n5857), .B2(n5882), .ZN(n5836)
         );
  AOI21_X1 U6910 ( .B1(n6417), .B2(n5859), .A(n5836), .ZN(n5837) );
  OAI211_X1 U6911 ( .C1(n6373), .C2(n5862), .A(n5838), .B(n5837), .ZN(U3085)
         );
  NAND2_X1 U6912 ( .A1(n5856), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5841) );
  OAI22_X1 U6913 ( .A1(n6385), .A2(n6428), .B1(n5857), .B2(n5886), .ZN(n5839)
         );
  AOI21_X1 U6914 ( .B1(n6423), .B2(n5859), .A(n5839), .ZN(n5840) );
  OAI211_X1 U6915 ( .C1(n6329), .C2(n5862), .A(n5841), .B(n5840), .ZN(U3086)
         );
  NAND2_X1 U6916 ( .A1(n5856), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5845) );
  OAI22_X1 U6917 ( .A1(n6385), .A2(n5842), .B1(n5857), .B2(n5890), .ZN(n5843)
         );
  AOI21_X1 U6918 ( .B1(n6429), .B2(n5859), .A(n5843), .ZN(n5844) );
  OAI211_X1 U6919 ( .C1(n6434), .C2(n5862), .A(n5845), .B(n5844), .ZN(U3087)
         );
  NAND2_X1 U6920 ( .A1(n5856), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5848) );
  OAI22_X1 U6921 ( .A1(n6385), .A2(n6440), .B1(n5857), .B2(n5894), .ZN(n5846)
         );
  AOI21_X1 U6922 ( .B1(n6435), .B2(n5859), .A(n5846), .ZN(n5847) );
  OAI211_X1 U6923 ( .C1(n6381), .C2(n5862), .A(n5848), .B(n5847), .ZN(U3088)
         );
  NAND2_X1 U6924 ( .A1(n5856), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5852) );
  OAI22_X1 U6925 ( .A1(n6385), .A2(n5849), .B1(n5857), .B2(n5898), .ZN(n5850)
         );
  AOI21_X1 U6926 ( .B1(n6441), .B2(n5859), .A(n5850), .ZN(n5851) );
  OAI211_X1 U6927 ( .C1(n6446), .C2(n5862), .A(n5852), .B(n5851), .ZN(U3089)
         );
  NAND2_X1 U6928 ( .A1(n5856), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5855) );
  OAI22_X1 U6929 ( .A1(n6385), .A2(n6389), .B1(n5857), .B2(n5902), .ZN(n5853)
         );
  AOI21_X1 U6930 ( .B1(n6447), .B2(n5859), .A(n5853), .ZN(n5854) );
  OAI211_X1 U6931 ( .C1(n6454), .C2(n5862), .A(n5855), .B(n5854), .ZN(U3090)
         );
  NAND2_X1 U6932 ( .A1(n5856), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5861) );
  OAI22_X1 U6933 ( .A1(n6385), .A2(n6465), .B1(n5857), .B2(n5909), .ZN(n5858)
         );
  AOI21_X1 U6934 ( .B1(n6456), .B2(n5859), .A(n5858), .ZN(n5860) );
  OAI211_X1 U6935 ( .C1(n6308), .C2(n5862), .A(n5861), .B(n5860), .ZN(U3091)
         );
  AND2_X1 U6936 ( .A1(n5865), .A2(n4590), .ZN(n6277) );
  NAND3_X1 U6937 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6474), .ZN(n6410) );
  NOR2_X1 U6938 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6410), .ZN(n5904)
         );
  NOR2_X1 U6939 ( .A1(n5869), .A2(n5868), .ZN(n6285) );
  INV_X1 U6940 ( .A(n6404), .ZN(n5871) );
  INV_X1 U6941 ( .A(n5904), .ZN(n5870) );
  AOI22_X1 U6942 ( .A1(n5872), .A2(n5871), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5870), .ZN(n5873) );
  AOI22_X1 U6943 ( .A1(n6399), .A2(n5904), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5903), .ZN(n5875) );
  OAI21_X1 U6944 ( .B1(n6369), .B2(n6464), .A(n5875), .ZN(n5876) );
  AOI21_X1 U6945 ( .B1(n6355), .B2(n5907), .A(n5876), .ZN(n5877) );
  OAI21_X1 U6946 ( .B1(n5910), .B2(n5878), .A(n5877), .ZN(U3100) );
  AOI22_X1 U6947 ( .A1(n6417), .A2(n5904), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5903), .ZN(n5879) );
  OAI21_X1 U6948 ( .B1(n6373), .B2(n6464), .A(n5879), .ZN(n5880) );
  AOI21_X1 U6949 ( .B1(n5907), .B2(n6370), .A(n5880), .ZN(n5881) );
  OAI21_X1 U6950 ( .B1(n5910), .B2(n5882), .A(n5881), .ZN(U3101) );
  AOI22_X1 U6951 ( .A1(n6423), .A2(n5904), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5903), .ZN(n5883) );
  OAI21_X1 U6952 ( .B1(n6329), .B2(n6464), .A(n5883), .ZN(n5884) );
  AOI21_X1 U6953 ( .B1(n5907), .B2(n6326), .A(n5884), .ZN(n5885) );
  OAI21_X1 U6954 ( .B1(n5910), .B2(n5886), .A(n5885), .ZN(U3102) );
  AOI22_X1 U6955 ( .A1(n6429), .A2(n5904), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5903), .ZN(n5887) );
  OAI21_X1 U6956 ( .B1(n6434), .B2(n6464), .A(n5887), .ZN(n5888) );
  AOI21_X1 U6957 ( .B1(n5907), .B2(n6430), .A(n5888), .ZN(n5889) );
  OAI21_X1 U6958 ( .B1(n5910), .B2(n5890), .A(n5889), .ZN(U3103) );
  AOI22_X1 U6959 ( .A1(n6435), .A2(n5904), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5903), .ZN(n5891) );
  OAI21_X1 U6960 ( .B1(n6381), .B2(n6464), .A(n5891), .ZN(n5892) );
  AOI21_X1 U6961 ( .B1(n5907), .B2(n6378), .A(n5892), .ZN(n5893) );
  OAI21_X1 U6962 ( .B1(n5910), .B2(n5894), .A(n5893), .ZN(U3104) );
  AOI22_X1 U6963 ( .A1(n6441), .A2(n5904), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5903), .ZN(n5895) );
  OAI21_X1 U6964 ( .B1(n6446), .B2(n6464), .A(n5895), .ZN(n5896) );
  AOI21_X1 U6965 ( .B1(n5907), .B2(n6442), .A(n5896), .ZN(n5897) );
  OAI21_X1 U6966 ( .B1(n5910), .B2(n5898), .A(n5897), .ZN(U3105) );
  AOI22_X1 U6967 ( .A1(n6447), .A2(n5904), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5903), .ZN(n5899) );
  OAI21_X1 U6968 ( .B1(n6454), .B2(n6464), .A(n5899), .ZN(n5900) );
  AOI21_X1 U6969 ( .B1(n5907), .B2(n6448), .A(n5900), .ZN(n5901) );
  OAI21_X1 U6970 ( .B1(n5910), .B2(n5902), .A(n5901), .ZN(U3106) );
  AOI22_X1 U6971 ( .A1(n6456), .A2(n5904), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5903), .ZN(n5905) );
  OAI21_X1 U6972 ( .B1(n6308), .B2(n6464), .A(n5905), .ZN(n5906) );
  AOI21_X1 U6973 ( .B1(n5907), .B2(n6304), .A(n5906), .ZN(n5908) );
  OAI21_X1 U6974 ( .B1(n5910), .B2(n5909), .A(n5908), .ZN(U3107) );
  AND2_X1 U6975 ( .A1(n6112), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6976 ( .A1(n6233), .A2(REIP_REG_13__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n5565), .ZN(n5915) );
  INV_X1 U6977 ( .A(n5911), .ZN(n6060) );
  XNOR2_X1 U6978 ( .A(n5912), .B(n5913), .ZN(n5921) );
  AOI22_X1 U6979 ( .A1(n6060), .A2(n6177), .B1(n3910), .B2(n5921), .ZN(n5914)
         );
  OAI211_X1 U6980 ( .C1(n6182), .C2(n5984), .A(n5915), .B(n5914), .ZN(U2973)
         );
  AOI21_X1 U6981 ( .B1(n5917), .B2(n5916), .A(n5359), .ZN(n6059) );
  AOI22_X1 U6982 ( .A1(n6059), .A2(n6262), .B1(n6233), .B2(
        REIP_REG_13__SCAN_IN), .ZN(n5923) );
  INV_X1 U6983 ( .A(n5918), .ZN(n5920) );
  AOI22_X1 U6984 ( .A1(n5921), .A2(n6266), .B1(n5920), .B2(n5919), .ZN(n5922)
         );
  OAI211_X1 U6985 ( .C1(n5925), .C2(n5924), .A(n5923), .B(n5922), .ZN(U3005)
         );
  OR4_X1 U6986 ( .A1(n6036), .A2(n5928), .A3(n5927), .A4(n5926), .ZN(n5929) );
  OAI21_X1 U6987 ( .B1(n5930), .B2(n3884), .A(n5929), .ZN(U3455) );
  INV_X1 U6988 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6752) );
  AOI21_X1 U6989 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6752), .A(n4196), .ZN(n5937) );
  INV_X1 U6990 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5931) );
  INV_X1 U6991 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6524) );
  AOI21_X1 U6992 ( .B1(n5937), .B2(n5931), .A(n6615), .ZN(U2789) );
  NAND2_X1 U6993 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6610), .ZN(n5935) );
  INV_X1 U6994 ( .A(n6511), .ZN(n5932) );
  OAI21_X1 U6995 ( .B1(n5933), .B2(n5932), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5934) );
  OAI21_X1 U6996 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5935), .A(n5934), .ZN(
        U2790) );
  NOR2_X1 U6997 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5938) );
  OAI21_X1 U6998 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5938), .A(n6579), .ZN(n5936)
         );
  OAI21_X1 U6999 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6598), .A(n5936), .ZN(
        U2791) );
  NOR2_X1 U7000 ( .A1(n6615), .A2(n5937), .ZN(n6585) );
  OAI21_X1 U7001 ( .B1(BS16_N), .B2(n5938), .A(n6585), .ZN(n6583) );
  OAI21_X1 U7002 ( .B1(n6585), .B2(n6604), .A(n6583), .ZN(U2792) );
  INV_X1 U7003 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5939) );
  OAI21_X1 U7004 ( .B1(n5940), .B2(n5939), .A(n6159), .ZN(U2793) );
  NOR4_X1 U7005 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n5944) );
  NOR4_X1 U7006 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n5943) );
  NOR4_X1 U7007 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5942) );
  NOR4_X1 U7008 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n5941) );
  NAND4_X1 U7009 ( .A1(n5944), .A2(n5943), .A3(n5942), .A4(n5941), .ZN(n5950)
         );
  NOR4_X1 U7010 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), 
        .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(DATAWIDTH_REG_5__SCAN_IN), .ZN(
        n5948) );
  AOI211_X1 U7011 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_20__SCAN_IN), .B(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n5947) );
  NOR4_X1 U7012 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(
        DATAWIDTH_REG_13__SCAN_IN), .ZN(n5946) );
  NOR4_X1 U7013 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(
        n5945) );
  NAND4_X1 U7014 ( .A1(n5948), .A2(n5947), .A3(n5946), .A4(n5945), .ZN(n5949)
         );
  NOR2_X1 U7015 ( .A1(n5950), .A2(n5949), .ZN(n6596) );
  INV_X1 U7016 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5952) );
  NOR3_X1 U7017 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5953) );
  OAI21_X1 U7018 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5953), .A(n6596), .ZN(n5951)
         );
  OAI21_X1 U7019 ( .B1(n6596), .B2(n5952), .A(n5951), .ZN(U2794) );
  INV_X1 U7020 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6584) );
  AOI21_X1 U7021 ( .B1(n6589), .B2(n6584), .A(n5953), .ZN(n5954) );
  INV_X1 U7022 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6683) );
  INV_X1 U7023 ( .A(n6596), .ZN(n6591) );
  AOI22_X1 U7024 ( .A1(n6596), .A2(n5954), .B1(n6683), .B2(n6591), .ZN(U2795)
         );
  AOI21_X1 U7025 ( .B1(n6779), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6033), 
        .ZN(n5964) );
  AOI22_X1 U7026 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6780), .B1(n5955), .B2(n6054), .ZN(n5963) );
  AOI22_X1 U7027 ( .A1(n5960), .A2(n6551), .B1(n5965), .B2(n6030), .ZN(n5956)
         );
  INV_X1 U7028 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5959) );
  OAI22_X1 U7029 ( .A1(n5957), .A2(n6044), .B1(n5956), .B2(n5959), .ZN(n5958)
         );
  AOI21_X1 U7030 ( .B1(n6074), .B2(n6025), .A(n5958), .ZN(n5962) );
  NAND3_X1 U7031 ( .A1(n5960), .A2(REIP_REG_15__SCAN_IN), .A3(n5959), .ZN(
        n5961) );
  NAND4_X1 U7032 ( .A1(n5964), .A2(n5963), .A3(n5962), .A4(n5961), .ZN(U2811)
         );
  NAND3_X1 U7033 ( .A1(n6030), .A2(REIP_REG_14__SCAN_IN), .A3(n5965), .ZN(
        n5966) );
  OAI21_X1 U7034 ( .B1(n5967), .B2(n6044), .A(n5966), .ZN(n5968) );
  INV_X1 U7035 ( .A(n5968), .ZN(n5975) );
  AOI22_X1 U7036 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6780), .B1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n6779), .ZN(n5974) );
  NOR2_X1 U7037 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5976), .ZN(n5969) );
  AOI21_X1 U7038 ( .B1(REIP_REG_13__SCAN_IN), .B2(n5969), .A(n6033), .ZN(n5973) );
  AOI22_X1 U7039 ( .A1(n5971), .A2(n6025), .B1(n5970), .B2(n6054), .ZN(n5972)
         );
  NAND4_X1 U7040 ( .A1(n5975), .A2(n5974), .A3(n5973), .A4(n5972), .ZN(U2813)
         );
  NOR2_X1 U7041 ( .A1(n5976), .A2(REIP_REG_13__SCAN_IN), .ZN(n5979) );
  INV_X1 U7042 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7043 ( .A1(n6779), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5977)
         );
  OAI211_X1 U7044 ( .C1(n6029), .C2(n6062), .A(n5977), .B(n6781), .ZN(n5978)
         );
  AOI211_X1 U7045 ( .C1(n6059), .C2(n6787), .A(n5979), .B(n5978), .ZN(n5983)
         );
  OAI21_X1 U7046 ( .B1(n3017), .B2(n6773), .A(n6030), .ZN(n6783) );
  OAI21_X1 U7047 ( .B1(REIP_REG_12__SCAN_IN), .B2(n5980), .A(n6783), .ZN(n5981) );
  AOI22_X1 U7048 ( .A1(n6060), .A2(n6025), .B1(REIP_REG_13__SCAN_IN), .B2(
        n5981), .ZN(n5982) );
  OAI211_X1 U7049 ( .C1(n5984), .C2(n6778), .A(n5983), .B(n5982), .ZN(U2814)
         );
  AOI21_X1 U7050 ( .B1(n5985), .B2(n6004), .A(REIP_REG_11__SCAN_IN), .ZN(n5994) );
  INV_X1 U7051 ( .A(n5276), .ZN(n5989) );
  INV_X1 U7052 ( .A(n5986), .ZN(n5988) );
  OAI21_X1 U7053 ( .B1(n5989), .B2(n5988), .A(n5987), .ZN(n6183) );
  INV_X1 U7054 ( .A(n6183), .ZN(n6063) );
  INV_X1 U7055 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6720) );
  NOR2_X1 U7056 ( .A1(n6029), .A2(n6720), .ZN(n5991) );
  OAI21_X1 U7057 ( .B1(n6047), .B2(n6673), .A(n6781), .ZN(n5990) );
  AOI211_X1 U7058 ( .C1(n6063), .C2(n6787), .A(n5991), .B(n5990), .ZN(n5993)
         );
  AOI22_X1 U7059 ( .A1(n6151), .A2(n6025), .B1(n6054), .B2(n6149), .ZN(n5992)
         );
  OAI211_X1 U7060 ( .C1(n5994), .C2(n6783), .A(n5993), .B(n5992), .ZN(U2816)
         );
  INV_X1 U7061 ( .A(n5995), .ZN(n5997) );
  AOI22_X1 U7062 ( .A1(n5997), .A2(n6025), .B1(n6054), .B2(n5996), .ZN(n6006)
         );
  OAI22_X1 U7063 ( .A1(n6029), .A2(n5998), .B1(n6044), .B2(n6204), .ZN(n5999)
         );
  INV_X1 U7064 ( .A(n5999), .ZN(n6000) );
  OAI211_X1 U7065 ( .C1(n6047), .C2(n6001), .A(n6000), .B(n6781), .ZN(n6002)
         );
  AOI221_X1 U7066 ( .B1(n6004), .B2(n6543), .C1(n6003), .C2(
        REIP_REG_9__SCAN_IN), .A(n6002), .ZN(n6005) );
  NAND2_X1 U7067 ( .A1(n6006), .A2(n6005), .ZN(U2818) );
  NAND2_X1 U7068 ( .A1(n6007), .A2(n6538), .ZN(n6021) );
  INV_X1 U7069 ( .A(n6008), .ZN(n6009) );
  AOI22_X1 U7070 ( .A1(n6787), .A2(n6222), .B1(n6009), .B2(n6054), .ZN(n6010)
         );
  OAI211_X1 U7071 ( .C1(n6047), .C2(n6011), .A(n6010), .B(n6781), .ZN(n6015)
         );
  OAI22_X1 U7072 ( .A1(n6013), .A2(n6790), .B1(REIP_REG_7__SCAN_IN), .B2(n6012), .ZN(n6014) );
  AOI211_X1 U7073 ( .C1(EBX_REG_7__SCAN_IN), .C2(n6780), .A(n6015), .B(n6014), 
        .ZN(n6016) );
  OAI221_X1 U7074 ( .B1(n6017), .B2(n6019), .C1(n6017), .C2(n6021), .A(n6016), 
        .ZN(U2820) );
  OAI22_X1 U7075 ( .A1(n6538), .A2(n6019), .B1(n6044), .B2(n6018), .ZN(n6020)
         );
  AOI211_X1 U7076 ( .C1(n6779), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6033), 
        .B(n6020), .ZN(n6022) );
  OAI211_X1 U7077 ( .C1(n6029), .C2(n6023), .A(n6022), .B(n6021), .ZN(n6024)
         );
  AOI21_X1 U7078 ( .B1(n6026), .B2(n6025), .A(n6024), .ZN(n6027) );
  OAI21_X1 U7079 ( .B1(n6163), .B2(n6778), .A(n6027), .ZN(U2821) );
  OR2_X1 U7080 ( .A1(n6029), .A2(n6028), .ZN(n6035) );
  OAI21_X1 U7081 ( .B1(n3017), .B2(n6031), .A(n6030), .ZN(n6058) );
  OAI22_X1 U7082 ( .A1(n6740), .A2(n6058), .B1(n6044), .B2(n6241), .ZN(n6032)
         );
  AOI211_X1 U7083 ( .C1(n6779), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6033), 
        .B(n6032), .ZN(n6034) );
  OAI211_X1 U7084 ( .C1(n6045), .C2(n6036), .A(n6035), .B(n6034), .ZN(n6039)
         );
  NOR2_X1 U7085 ( .A1(n6037), .A2(n6051), .ZN(n6038) );
  AOI211_X1 U7086 ( .C1(n6040), .C2(n6740), .A(n6039), .B(n6038), .ZN(n6041)
         );
  OAI21_X1 U7087 ( .B1(n6172), .B2(n6778), .A(n6041), .ZN(U2823) );
  INV_X1 U7088 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6658) );
  OR2_X1 U7089 ( .A1(n6043), .A2(n6042), .ZN(n6057) );
  NOR2_X1 U7090 ( .A1(n6044), .A2(n6249), .ZN(n6049) );
  OAI22_X1 U7091 ( .A1(n6047), .A2(n6046), .B1(n6045), .B2(n6278), .ZN(n6048)
         );
  AOI211_X1 U7092 ( .C1(n6780), .C2(EBX_REG_3__SCAN_IN), .A(n6049), .B(n6048), 
        .ZN(n6050) );
  OAI21_X1 U7093 ( .B1(n6052), .B2(n6051), .A(n6050), .ZN(n6053) );
  AOI21_X1 U7094 ( .B1(n6055), .B2(n6054), .A(n6053), .ZN(n6056) );
  OAI221_X1 U7095 ( .B1(n6058), .B2(n6658), .C1(n6058), .C2(n6057), .A(n6056), 
        .ZN(U2824) );
  AOI22_X1 U7096 ( .A1(n6060), .A2(n4264), .B1(n6065), .B2(n6059), .ZN(n6061)
         );
  OAI21_X1 U7097 ( .B1(n6062), .B2(n6067), .A(n6061), .ZN(U2846) );
  AOI22_X1 U7098 ( .A1(n6151), .A2(n4264), .B1(n6065), .B2(n6063), .ZN(n6064)
         );
  OAI21_X1 U7099 ( .B1(n6720), .B2(n6067), .A(n6064), .ZN(U2848) );
  AOI22_X1 U7100 ( .A1(n6178), .A2(n4264), .B1(n6065), .B2(n6261), .ZN(n6066)
         );
  OAI21_X1 U7101 ( .B1(n6068), .B2(n6067), .A(n6066), .ZN(U2857) );
  AOI22_X1 U7102 ( .A1(n6069), .A2(n6073), .B1(n6072), .B2(DATAI_17_), .ZN(
        n6071) );
  AOI22_X1 U7103 ( .A1(n6076), .A2(DATAI_1_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n6075), .ZN(n6070) );
  NAND2_X1 U7104 ( .A1(n6071), .A2(n6070), .ZN(U2874) );
  AOI22_X1 U7105 ( .A1(n6074), .A2(n6073), .B1(n6072), .B2(DATAI_16_), .ZN(
        n6078) );
  AOI22_X1 U7106 ( .A1(n6076), .A2(DATAI_0_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n6075), .ZN(n6077) );
  NAND2_X1 U7107 ( .A1(n6078), .A2(n6077), .ZN(U2875) );
  INV_X1 U7108 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n6637) );
  INV_X1 U7109 ( .A(n6079), .ZN(n6082) );
  AOI22_X1 U7110 ( .A1(n6112), .A2(DATAO_REG_24__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n6082), .ZN(n6080) );
  OAI21_X1 U7111 ( .B1(n6637), .B2(n6111), .A(n6080), .ZN(U2899) );
  INV_X1 U7112 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n6689) );
  AOI22_X1 U7113 ( .A1(n6082), .A2(EAX_REG_18__SCAN_IN), .B1(
        UWORD_REG_2__SCAN_IN), .B2(n6601), .ZN(n6081) );
  OAI21_X1 U7114 ( .B1(n6689), .B2(n6108), .A(n6081), .ZN(U2905) );
  INV_X1 U7115 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n6719) );
  AOI22_X1 U7116 ( .A1(n6112), .A2(DATAO_REG_16__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6082), .ZN(n6083) );
  OAI21_X1 U7117 ( .B1(n6719), .B2(n6111), .A(n6083), .ZN(U2907) );
  AOI22_X1 U7118 ( .A1(LWORD_REG_15__SCAN_IN), .A2(n6601), .B1(n6112), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6084) );
  OAI21_X1 U7119 ( .B1(n4458), .B2(n6114), .A(n6084), .ZN(U2908) );
  INV_X1 U7120 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n6739) );
  AOI22_X1 U7121 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6098), .B1(
        LWORD_REG_14__SCAN_IN), .B2(n6085), .ZN(n6086) );
  OAI21_X1 U7122 ( .B1(n6739), .B2(n6108), .A(n6086), .ZN(U2909) );
  AOI22_X1 U7123 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n6601), .B1(n6112), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6087) );
  OAI21_X1 U7124 ( .B1(n6641), .B2(n6114), .A(n6087), .ZN(U2910) );
  INV_X1 U7125 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6089) );
  AOI22_X1 U7126 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n6601), .B1(n6112), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6088) );
  OAI21_X1 U7127 ( .B1(n6089), .B2(n6114), .A(n6088), .ZN(U2911) );
  INV_X1 U7128 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6091) );
  AOI22_X1 U7129 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6601), .B1(n6112), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6090) );
  OAI21_X1 U7130 ( .B1(n6091), .B2(n6114), .A(n6090), .ZN(U2912) );
  INV_X1 U7131 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6093) );
  AOI22_X1 U7132 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n6601), .B1(n6112), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6092) );
  OAI21_X1 U7133 ( .B1(n6093), .B2(n6114), .A(n6092), .ZN(U2913) );
  INV_X1 U7134 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6095) );
  AOI22_X1 U7135 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n6601), .B1(n6112), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6094) );
  OAI21_X1 U7136 ( .B1(n6095), .B2(n6114), .A(n6094), .ZN(U2914) );
  INV_X1 U7137 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6129) );
  AOI22_X1 U7138 ( .A1(LWORD_REG_8__SCAN_IN), .A2(n6601), .B1(n6112), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6096) );
  OAI21_X1 U7139 ( .B1(n6129), .B2(n6114), .A(n6096), .ZN(U2915) );
  INV_X1 U7140 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n6661) );
  AOI22_X1 U7141 ( .A1(EAX_REG_7__SCAN_IN), .A2(n6098), .B1(n6112), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6097) );
  OAI21_X1 U7142 ( .B1(n6661), .B2(n6111), .A(n6097), .ZN(U2916) );
  INV_X1 U7143 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n6676) );
  AOI22_X1 U7144 ( .A1(EAX_REG_6__SCAN_IN), .A2(n6098), .B1(n6112), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6099) );
  OAI21_X1 U7145 ( .B1(n6676), .B2(n6111), .A(n6099), .ZN(U2917) );
  AOI22_X1 U7146 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n6601), .B1(n6112), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6100) );
  OAI21_X1 U7147 ( .B1(n6101), .B2(n6114), .A(n6100), .ZN(U2918) );
  AOI22_X1 U7148 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n6601), .B1(n6112), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6102) );
  OAI21_X1 U7149 ( .B1(n6103), .B2(n6114), .A(n6102), .ZN(U2919) );
  AOI22_X1 U7150 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n6601), .B1(n6112), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6104) );
  OAI21_X1 U7151 ( .B1(n6105), .B2(n6114), .A(n6104), .ZN(U2920) );
  AOI22_X1 U7152 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n6601), .B1(n6112), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6106) );
  OAI21_X1 U7153 ( .B1(n6107), .B2(n6114), .A(n6106), .ZN(U2921) );
  INV_X1 U7154 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n6110) );
  INV_X1 U7155 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n6725) );
  OAI222_X1 U7156 ( .A1(n6111), .A2(n6110), .B1(n6114), .B2(n6109), .C1(n6725), 
        .C2(n6108), .ZN(U2922) );
  AOI22_X1 U7157 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n6601), .B1(n6112), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6113) );
  OAI21_X1 U7158 ( .B1(n6115), .B2(n6114), .A(n6113), .ZN(U2923) );
  INV_X1 U7159 ( .A(n6140), .ZN(n6118) );
  INV_X1 U7160 ( .A(DATAI_8_), .ZN(n6116) );
  NOR2_X1 U7161 ( .A1(n6125), .A2(n6116), .ZN(n6127) );
  AOI21_X1 U7162 ( .B1(n6136), .B2(EAX_REG_24__SCAN_IN), .A(n6127), .ZN(n6117)
         );
  OAI21_X1 U7163 ( .B1(n6637), .B2(n6118), .A(n6117), .ZN(U2932) );
  AOI22_X1 U7164 ( .A1(EAX_REG_25__SCAN_IN), .A2(n6136), .B1(n6140), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7165 ( .A1(n6122), .A2(DATAI_9_), .ZN(n6130) );
  NAND2_X1 U7166 ( .A1(n6119), .A2(n6130), .ZN(U2933) );
  AOI22_X1 U7167 ( .A1(EAX_REG_26__SCAN_IN), .A2(n6136), .B1(n6140), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7168 ( .A1(n6122), .A2(DATAI_10_), .ZN(n6132) );
  NAND2_X1 U7169 ( .A1(n6120), .A2(n6132), .ZN(U2934) );
  AOI22_X1 U7170 ( .A1(EAX_REG_27__SCAN_IN), .A2(n6136), .B1(n6140), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7171 ( .A1(n6122), .A2(DATAI_11_), .ZN(n6134) );
  NAND2_X1 U7172 ( .A1(n6121), .A2(n6134), .ZN(U2935) );
  AOI22_X1 U7173 ( .A1(EAX_REG_28__SCAN_IN), .A2(n6136), .B1(n6140), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7174 ( .A1(n6122), .A2(DATAI_12_), .ZN(n6137) );
  NAND2_X1 U7175 ( .A1(n6123), .A2(n6137), .ZN(U2936) );
  NOR2_X1 U7176 ( .A1(n6125), .A2(n6124), .ZN(n6139) );
  AOI21_X1 U7177 ( .B1(n6140), .B2(UWORD_REG_13__SCAN_IN), .A(n6139), .ZN(
        n6126) );
  OAI21_X1 U7178 ( .B1(n6652), .B2(n6142), .A(n6126), .ZN(U2937) );
  AOI21_X1 U7179 ( .B1(n6140), .B2(LWORD_REG_8__SCAN_IN), .A(n6127), .ZN(n6128) );
  OAI21_X1 U7180 ( .B1(n6129), .B2(n6142), .A(n6128), .ZN(U2947) );
  AOI22_X1 U7181 ( .A1(EAX_REG_9__SCAN_IN), .A2(n6136), .B1(n6140), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7182 ( .A1(n6131), .A2(n6130), .ZN(U2948) );
  AOI22_X1 U7183 ( .A1(EAX_REG_10__SCAN_IN), .A2(n6136), .B1(n6140), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n6133) );
  NAND2_X1 U7184 ( .A1(n6133), .A2(n6132), .ZN(U2949) );
  AOI22_X1 U7185 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6136), .B1(n6140), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7186 ( .A1(n6135), .A2(n6134), .ZN(U2950) );
  AOI22_X1 U7187 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6136), .B1(n6140), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7188 ( .A1(n6138), .A2(n6137), .ZN(U2951) );
  AOI21_X1 U7189 ( .B1(n6140), .B2(LWORD_REG_13__SCAN_IN), .A(n6139), .ZN(
        n6141) );
  OAI21_X1 U7190 ( .B1(n6641), .B2(n6142), .A(n6141), .ZN(U2952) );
  OAI21_X1 U7191 ( .B1(n6145), .B2(n6144), .A(n6143), .ZN(n6148) );
  XNOR2_X1 U7192 ( .A(n6146), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6147)
         );
  XNOR2_X1 U7193 ( .A(n6148), .B(n6147), .ZN(n6185) );
  AOI22_X1 U7194 ( .A1(n6233), .A2(REIP_REG_11__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n5565), .ZN(n6153) );
  AOI22_X1 U7195 ( .A1(n6151), .A2(n6177), .B1(n6150), .B2(n6149), .ZN(n6152)
         );
  OAI211_X1 U7196 ( .C1(n6185), .C2(n6159), .A(n6153), .B(n6152), .ZN(U2975)
         );
  AOI22_X1 U7197 ( .A1(n6233), .A2(REIP_REG_6__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n5565), .ZN(n6162) );
  OAI21_X1 U7198 ( .B1(n6154), .B2(n6156), .A(n6155), .ZN(n6230) );
  OAI22_X1 U7199 ( .A1(n6230), .A2(n6159), .B1(n6158), .B2(n6157), .ZN(n6160)
         );
  INV_X1 U7200 ( .A(n6160), .ZN(n6161) );
  OAI211_X1 U7201 ( .C1(n6182), .C2(n6163), .A(n6162), .B(n6161), .ZN(U2980)
         );
  AOI22_X1 U7202 ( .A1(n6233), .A2(REIP_REG_4__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n5565), .ZN(n6171) );
  INV_X1 U7203 ( .A(n6164), .ZN(n6165) );
  NAND2_X1 U7204 ( .A1(n6246), .A2(n6165), .ZN(n6168) );
  XNOR2_X1 U7205 ( .A(n6166), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6167)
         );
  XNOR2_X1 U7206 ( .A(n6168), .B(n6167), .ZN(n6240) );
  AOI22_X1 U7207 ( .A1(n6169), .A2(n6177), .B1(n3910), .B2(n6240), .ZN(n6170)
         );
  OAI211_X1 U7208 ( .C1(n6182), .C2(n6172), .A(n6171), .B(n6170), .ZN(U2982)
         );
  AOI22_X1 U7209 ( .A1(n6233), .A2(REIP_REG_2__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n5565), .ZN(n6180) );
  XNOR2_X1 U7210 ( .A(n6174), .B(n6173), .ZN(n6176) );
  XNOR2_X1 U7211 ( .A(n6176), .B(n6175), .ZN(n6265) );
  AOI22_X1 U7212 ( .A1(n6178), .A2(n6177), .B1(n3910), .B2(n6265), .ZN(n6179)
         );
  OAI211_X1 U7213 ( .C1(n6182), .C2(n6181), .A(n6180), .B(n6179), .ZN(U2984)
         );
  INV_X1 U7214 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6674) );
  OAI22_X1 U7215 ( .A1(n6183), .A2(n6250), .B1(n6674), .B2(n6248), .ZN(n6187)
         );
  NOR2_X1 U7216 ( .A1(n6185), .A2(n6184), .ZN(n6186) );
  AOI211_X1 U7217 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n6188), .A(n6187), .B(n6186), .ZN(n6190) );
  NAND2_X1 U7218 ( .A1(n6190), .A2(n6189), .ZN(U3007) );
  AOI22_X1 U7219 ( .A1(n6194), .A2(n6193), .B1(n6192), .B2(n6191), .ZN(n6195)
         );
  INV_X1 U7220 ( .A(n6195), .ZN(n6225) );
  AOI21_X1 U7221 ( .B1(n6213), .B2(n6196), .A(n6225), .ZN(n6212) );
  OAI22_X1 U7222 ( .A1(n6197), .A2(n6250), .B1(n6542), .B2(n6248), .ZN(n6198)
         );
  AOI21_X1 U7223 ( .B1(n6199), .B2(n6266), .A(n6198), .ZN(n6203) );
  OAI21_X1 U7224 ( .B1(n6259), .B2(n6268), .A(n6200), .ZN(n6239) );
  NAND2_X1 U7225 ( .A1(n6201), .A2(n6239), .ZN(n6228) );
  NOR2_X1 U7226 ( .A1(n6213), .A2(n6228), .ZN(n6208) );
  OAI221_X1 U7227 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n6710), .C2(n6735), .A(n6208), 
        .ZN(n6202) );
  OAI211_X1 U7228 ( .C1(n6212), .C2(n6710), .A(n6203), .B(n6202), .ZN(U3008)
         );
  INV_X1 U7229 ( .A(n6204), .ZN(n6207) );
  INV_X1 U7230 ( .A(n6205), .ZN(n6206) );
  AOI21_X1 U7231 ( .B1(n6262), .B2(n6207), .A(n6206), .ZN(n6211) );
  AOI22_X1 U7232 ( .A1(n6209), .A2(n6266), .B1(n6208), .B2(n6735), .ZN(n6210)
         );
  OAI211_X1 U7233 ( .C1(n6212), .C2(n6735), .A(n6211), .B(n6210), .ZN(U3009)
         );
  OAI21_X1 U7234 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6213), .ZN(n6219) );
  AOI21_X1 U7235 ( .B1(n6262), .B2(n6215), .A(n6214), .ZN(n6218) );
  AOI22_X1 U7236 ( .A1(n6216), .A2(n6266), .B1(n6225), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6217) );
  OAI211_X1 U7237 ( .C1(n6228), .C2(n6219), .A(n6218), .B(n6217), .ZN(U3010)
         );
  INV_X1 U7238 ( .A(n6220), .ZN(n6221) );
  AOI21_X1 U7239 ( .B1(n6262), .B2(n6222), .A(n6221), .ZN(n6227) );
  INV_X1 U7240 ( .A(n6223), .ZN(n6224) );
  AOI22_X1 U7241 ( .A1(n6225), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .B1(n6266), 
        .B2(n6224), .ZN(n6226) );
  OAI211_X1 U7242 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6228), .A(n6227), 
        .B(n6226), .ZN(U3011) );
  NAND2_X1 U7243 ( .A1(n6239), .A2(n6229), .ZN(n6237) );
  INV_X1 U7244 ( .A(n6230), .ZN(n6231) );
  AOI222_X1 U7245 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6233), .B1(n6262), .B2(
        n6232), .C1(n6266), .C2(n6231), .ZN(n6234) );
  OAI221_X1 U7246 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6237), .C1(n6236), .C2(n6235), .A(n6234), .ZN(U3012) );
  INV_X1 U7247 ( .A(n6258), .ZN(n6238) );
  AOI21_X1 U7248 ( .B1(n6264), .B2(n6238), .A(n6267), .ZN(n6255) );
  NAND2_X1 U7249 ( .A1(n6239), .A2(n6258), .ZN(n6257) );
  AOI221_X1 U7250 ( .B1(INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .C1(n3762), .C2(n6256), .A(n6257), 
        .ZN(n6244) );
  AND2_X1 U7251 ( .A1(n6240), .A2(n6266), .ZN(n6243) );
  OAI22_X1 U7252 ( .A1(n6250), .A2(n6241), .B1(n6740), .B2(n6248), .ZN(n6242)
         );
  NOR3_X1 U7253 ( .A1(n6244), .A2(n6243), .A3(n6242), .ZN(n6245) );
  OAI21_X1 U7254 ( .B1(n6255), .B2(n3762), .A(n6245), .ZN(U3014) );
  NAND3_X1 U7255 ( .A1(n6247), .A2(n6266), .A3(n6246), .ZN(n6253) );
  OAI22_X1 U7256 ( .A1(n6250), .A2(n6249), .B1(n6658), .B2(n6248), .ZN(n6251)
         );
  INV_X1 U7257 ( .A(n6251), .ZN(n6252) );
  AND2_X1 U7258 ( .A1(n6253), .A2(n6252), .ZN(n6254) );
  OAI221_X1 U7259 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n6257), .C1(n6256), .C2(n6255), .A(n6254), .ZN(U3015) );
  OAI21_X1 U7260 ( .B1(n6260), .B2(n6259), .A(n6258), .ZN(n6263) );
  AOI22_X1 U7261 ( .A1(n6264), .A2(n6263), .B1(n6262), .B2(n6261), .ZN(n6273)
         );
  AOI22_X1 U7262 ( .A1(n6267), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6266), 
        .B2(n6265), .ZN(n6272) );
  NAND2_X1 U7263 ( .A1(n6233), .A2(REIP_REG_2__SCAN_IN), .ZN(n6271) );
  OR3_X1 U7264 ( .A1(n6269), .A2(n6268), .A3(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6270) );
  NAND4_X1 U7265 ( .A1(n6273), .A2(n6272), .A3(n6271), .A4(n6270), .ZN(U3016)
         );
  NOR2_X1 U7266 ( .A1(n6478), .A2(n6274), .ZN(U3019) );
  NAND3_X1 U7267 ( .A1(n4633), .A2(n6275), .A3(n2964), .ZN(n6276) );
  NAND3_X1 U7268 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6397), .A3(n6474), .ZN(n6319) );
  NOR2_X1 U7269 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6319), .ZN(n6302)
         );
  NAND2_X1 U7270 ( .A1(n6278), .A2(n6277), .ZN(n6314) );
  INV_X1 U7271 ( .A(n6279), .ZN(n6282) );
  INV_X1 U7272 ( .A(n6280), .ZN(n6281) );
  OAI22_X1 U7273 ( .A1(n6314), .A2(n6406), .B1(n6282), .B2(n6281), .ZN(n6301)
         );
  AOI22_X1 U7274 ( .A1(n6399), .A2(n6302), .B1(n6413), .B2(n6301), .ZN(n6288)
         );
  OAI21_X1 U7275 ( .B1(n6303), .B2(n6336), .A(n6283), .ZN(n6284) );
  AOI21_X1 U7276 ( .B1(n6284), .B2(n6314), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n6286) );
  AOI22_X1 U7277 ( .A1(n6305), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n6355), 
        .B2(n6303), .ZN(n6287) );
  OAI211_X1 U7278 ( .C1(n6369), .C2(n6346), .A(n6288), .B(n6287), .ZN(U3036)
         );
  AOI22_X1 U7279 ( .A1(n6417), .A2(n6302), .B1(n6419), .B2(n6301), .ZN(n6290)
         );
  AOI22_X1 U7280 ( .A1(n6305), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n6370), 
        .B2(n6303), .ZN(n6289) );
  OAI211_X1 U7281 ( .C1(n6346), .C2(n6373), .A(n6290), .B(n6289), .ZN(U3037)
         );
  AOI22_X1 U7282 ( .A1(n6423), .A2(n6302), .B1(n6425), .B2(n6301), .ZN(n6292)
         );
  AOI22_X1 U7283 ( .A1(n6305), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n6326), 
        .B2(n6303), .ZN(n6291) );
  OAI211_X1 U7284 ( .C1(n6346), .C2(n6329), .A(n6292), .B(n6291), .ZN(U3038)
         );
  AOI22_X1 U7285 ( .A1(n6429), .A2(n6302), .B1(n6431), .B2(n6301), .ZN(n6294)
         );
  AOI22_X1 U7286 ( .A1(n6305), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n6430), 
        .B2(n6303), .ZN(n6293) );
  OAI211_X1 U7287 ( .C1(n6346), .C2(n6434), .A(n6294), .B(n6293), .ZN(U3039)
         );
  AOI22_X1 U7288 ( .A1(n6435), .A2(n6302), .B1(n6437), .B2(n6301), .ZN(n6296)
         );
  AOI22_X1 U7289 ( .A1(n6305), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n6378), 
        .B2(n6303), .ZN(n6295) );
  OAI211_X1 U7290 ( .C1(n6346), .C2(n6381), .A(n6296), .B(n6295), .ZN(U3040)
         );
  AOI22_X1 U7291 ( .A1(n6441), .A2(n6302), .B1(n6443), .B2(n6301), .ZN(n6298)
         );
  AOI22_X1 U7292 ( .A1(n6305), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n6442), 
        .B2(n6303), .ZN(n6297) );
  OAI211_X1 U7293 ( .C1(n6346), .C2(n6446), .A(n6298), .B(n6297), .ZN(U3041)
         );
  AOI22_X1 U7294 ( .A1(n6447), .A2(n6302), .B1(n6450), .B2(n6301), .ZN(n6300)
         );
  AOI22_X1 U7295 ( .A1(n6305), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n6448), 
        .B2(n6303), .ZN(n6299) );
  OAI211_X1 U7296 ( .C1(n6346), .C2(n6454), .A(n6300), .B(n6299), .ZN(U3042)
         );
  AOI22_X1 U7297 ( .A1(n6456), .A2(n6302), .B1(n6460), .B2(n6301), .ZN(n6307)
         );
  AOI22_X1 U7298 ( .A1(n6305), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n6304), 
        .B2(n6303), .ZN(n6306) );
  OAI211_X1 U7299 ( .C1(n6346), .C2(n6308), .A(n6307), .B(n6306), .ZN(U3043)
         );
  INV_X1 U7300 ( .A(n6398), .ZN(n6309) );
  NAND2_X1 U7301 ( .A1(n6309), .A2(n6397), .ZN(n6315) );
  INV_X1 U7302 ( .A(n6315), .ZN(n6341) );
  INV_X1 U7303 ( .A(n6339), .ZN(n6340) );
  AOI22_X1 U7304 ( .A1(n6399), .A2(n6341), .B1(n6340), .B2(n6400), .ZN(n6323)
         );
  NAND2_X1 U7305 ( .A1(n6310), .A2(n4633), .ZN(n6311) );
  OAI21_X1 U7306 ( .B1(n6312), .B2(n6311), .A(n6401), .ZN(n6321) );
  OR2_X1 U7307 ( .A1(n6314), .A2(n6313), .ZN(n6316) );
  INV_X1 U7308 ( .A(n6320), .ZN(n6318) );
  AOI21_X1 U7309 ( .B1(n6406), .B2(n6319), .A(n6405), .ZN(n6317) );
  AOI22_X1 U7310 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6343), .B1(n6413), 
        .B2(n6342), .ZN(n6322) );
  OAI211_X1 U7311 ( .C1(n6416), .C2(n6346), .A(n6323), .B(n6322), .ZN(U3044)
         );
  AOI22_X1 U7312 ( .A1(n6417), .A2(n6341), .B1(n6340), .B2(n6418), .ZN(n6325)
         );
  AOI22_X1 U7313 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6343), .B1(n6419), 
        .B2(n6342), .ZN(n6324) );
  OAI211_X1 U7314 ( .C1(n6346), .C2(n6422), .A(n6325), .B(n6324), .ZN(U3045)
         );
  AOI22_X1 U7315 ( .A1(n6423), .A2(n6341), .B1(n6336), .B2(n6326), .ZN(n6328)
         );
  AOI22_X1 U7316 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6343), .B1(n6425), 
        .B2(n6342), .ZN(n6327) );
  OAI211_X1 U7317 ( .C1(n6329), .C2(n6339), .A(n6328), .B(n6327), .ZN(U3046)
         );
  AOI22_X1 U7318 ( .A1(n6429), .A2(n6341), .B1(n6336), .B2(n6430), .ZN(n6331)
         );
  AOI22_X1 U7319 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6343), .B1(n6431), 
        .B2(n6342), .ZN(n6330) );
  OAI211_X1 U7320 ( .C1(n6434), .C2(n6339), .A(n6331), .B(n6330), .ZN(U3047)
         );
  AOI22_X1 U7321 ( .A1(n6435), .A2(n6341), .B1(n6336), .B2(n6378), .ZN(n6333)
         );
  AOI22_X1 U7322 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6343), .B1(n6437), 
        .B2(n6342), .ZN(n6332) );
  OAI211_X1 U7323 ( .C1(n6381), .C2(n6339), .A(n6333), .B(n6332), .ZN(U3048)
         );
  AOI22_X1 U7324 ( .A1(n6441), .A2(n6341), .B1(n6336), .B2(n6442), .ZN(n6335)
         );
  AOI22_X1 U7325 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6343), .B1(n6443), 
        .B2(n6342), .ZN(n6334) );
  OAI211_X1 U7326 ( .C1(n6446), .C2(n6339), .A(n6335), .B(n6334), .ZN(U3049)
         );
  AOI22_X1 U7327 ( .A1(n6447), .A2(n6341), .B1(n6336), .B2(n6448), .ZN(n6338)
         );
  AOI22_X1 U7328 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6343), .B1(n6450), 
        .B2(n6342), .ZN(n6337) );
  OAI211_X1 U7329 ( .C1(n6454), .C2(n6339), .A(n6338), .B(n6337), .ZN(U3050)
         );
  AOI22_X1 U7330 ( .A1(n6456), .A2(n6341), .B1(n6340), .B2(n6457), .ZN(n6345)
         );
  AOI22_X1 U7331 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6343), .B1(n6460), 
        .B2(n6342), .ZN(n6344) );
  OAI211_X1 U7332 ( .C1(n6346), .C2(n6465), .A(n6345), .B(n6344), .ZN(U3051)
         );
  INV_X1 U7333 ( .A(n6347), .ZN(n6348) );
  AOI22_X1 U7334 ( .A1(n6399), .A2(n6349), .B1(n6413), .B2(n6348), .ZN(n6353)
         );
  AOI22_X1 U7335 ( .A1(n6351), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6355), 
        .B2(n6350), .ZN(n6352) );
  OAI211_X1 U7336 ( .C1(n6369), .C2(n6396), .A(n6353), .B(n6352), .ZN(U3068)
         );
  INV_X1 U7337 ( .A(n6354), .ZN(n6390) );
  AOI22_X1 U7338 ( .A1(n6355), .A2(n6382), .B1(n6399), .B2(n6390), .ZN(n6368)
         );
  NAND2_X1 U7339 ( .A1(n6356), .A2(n6401), .ZN(n6366) );
  INV_X1 U7340 ( .A(n6366), .ZN(n6360) );
  INV_X1 U7341 ( .A(n6357), .ZN(n6358) );
  AOI21_X1 U7342 ( .B1(n6359), .B2(n6358), .A(n6390), .ZN(n6365) );
  NAND2_X1 U7343 ( .A1(n6360), .A2(n6365), .ZN(n6362) );
  OAI211_X1 U7344 ( .C1(n6401), .C2(n6363), .A(n6362), .B(n6361), .ZN(n6393)
         );
  OAI22_X1 U7345 ( .A1(n6366), .A2(n6365), .B1(n6364), .B2(n6409), .ZN(n6392)
         );
  AOI22_X1 U7346 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6393), .B1(n6413), 
        .B2(n6392), .ZN(n6367) );
  OAI211_X1 U7347 ( .C1(n6369), .C2(n6385), .A(n6368), .B(n6367), .ZN(U3076)
         );
  AOI22_X1 U7348 ( .A1(n6370), .A2(n6382), .B1(n6417), .B2(n6390), .ZN(n6372)
         );
  AOI22_X1 U7349 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6393), .B1(n6419), 
        .B2(n6392), .ZN(n6371) );
  OAI211_X1 U7350 ( .C1(n6373), .C2(n6385), .A(n6372), .B(n6371), .ZN(U3077)
         );
  INV_X1 U7351 ( .A(n6385), .ZN(n6391) );
  AOI22_X1 U7352 ( .A1(n6424), .A2(n6391), .B1(n6423), .B2(n6390), .ZN(n6375)
         );
  AOI22_X1 U7353 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6393), .B1(n6425), 
        .B2(n6392), .ZN(n6374) );
  OAI211_X1 U7354 ( .C1(n6428), .C2(n6396), .A(n6375), .B(n6374), .ZN(U3078)
         );
  AOI22_X1 U7355 ( .A1(n6430), .A2(n6382), .B1(n6429), .B2(n6390), .ZN(n6377)
         );
  AOI22_X1 U7356 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6393), .B1(n6431), 
        .B2(n6392), .ZN(n6376) );
  OAI211_X1 U7357 ( .C1(n6434), .C2(n6385), .A(n6377), .B(n6376), .ZN(U3079)
         );
  AOI22_X1 U7358 ( .A1(n6378), .A2(n6382), .B1(n6435), .B2(n6390), .ZN(n6380)
         );
  AOI22_X1 U7359 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6393), .B1(n6437), 
        .B2(n6392), .ZN(n6379) );
  OAI211_X1 U7360 ( .C1(n6381), .C2(n6385), .A(n6380), .B(n6379), .ZN(U3080)
         );
  AOI22_X1 U7361 ( .A1(n6442), .A2(n6382), .B1(n6441), .B2(n6390), .ZN(n6384)
         );
  AOI22_X1 U7362 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6393), .B1(n6443), 
        .B2(n6392), .ZN(n6383) );
  OAI211_X1 U7363 ( .C1(n6446), .C2(n6385), .A(n6384), .B(n6383), .ZN(U3081)
         );
  AOI22_X1 U7364 ( .A1(n6386), .A2(n6391), .B1(n6447), .B2(n6390), .ZN(n6388)
         );
  AOI22_X1 U7365 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6393), .B1(n6450), 
        .B2(n6392), .ZN(n6387) );
  OAI211_X1 U7366 ( .C1(n6389), .C2(n6396), .A(n6388), .B(n6387), .ZN(U3082)
         );
  AOI22_X1 U7367 ( .A1(n6457), .A2(n6391), .B1(n6456), .B2(n6390), .ZN(n6395)
         );
  AOI22_X1 U7368 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6393), .B1(n6460), 
        .B2(n6392), .ZN(n6394) );
  OAI211_X1 U7369 ( .C1(n6465), .C2(n6396), .A(n6395), .B(n6394), .ZN(U3083)
         );
  NOR2_X1 U7370 ( .A1(n6398), .A2(n6397), .ZN(n6455) );
  AOI22_X1 U7371 ( .A1(n6458), .A2(n6400), .B1(n6399), .B2(n6455), .ZN(n6415)
         );
  OAI21_X1 U7372 ( .B1(n6403), .B2(n6402), .A(n6401), .ZN(n6412) );
  INV_X1 U7373 ( .A(n6411), .ZN(n6408) );
  AOI21_X1 U7374 ( .B1(n6406), .B2(n6410), .A(n6405), .ZN(n6407) );
  OAI22_X1 U7375 ( .A1(n6412), .A2(n6411), .B1(n6410), .B2(n6409), .ZN(n6459)
         );
  AOI22_X1 U7376 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6461), .B1(n6413), 
        .B2(n6459), .ZN(n6414) );
  OAI211_X1 U7377 ( .C1(n6416), .C2(n6464), .A(n6415), .B(n6414), .ZN(U3108)
         );
  AOI22_X1 U7378 ( .A1(n6458), .A2(n6418), .B1(n6417), .B2(n6455), .ZN(n6421)
         );
  AOI22_X1 U7379 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6461), .B1(n6419), 
        .B2(n6459), .ZN(n6420) );
  OAI211_X1 U7380 ( .C1(n6422), .C2(n6464), .A(n6421), .B(n6420), .ZN(U3109)
         );
  AOI22_X1 U7381 ( .A1(n6458), .A2(n6424), .B1(n6423), .B2(n6455), .ZN(n6427)
         );
  AOI22_X1 U7382 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6461), .B1(n6425), 
        .B2(n6459), .ZN(n6426) );
  OAI211_X1 U7383 ( .C1(n6428), .C2(n6464), .A(n6427), .B(n6426), .ZN(U3110)
         );
  AOI22_X1 U7384 ( .A1(n6449), .A2(n6430), .B1(n6429), .B2(n6455), .ZN(n6433)
         );
  AOI22_X1 U7385 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6461), .B1(n6431), 
        .B2(n6459), .ZN(n6432) );
  OAI211_X1 U7386 ( .C1(n6434), .C2(n6453), .A(n6433), .B(n6432), .ZN(U3111)
         );
  AOI22_X1 U7387 ( .A1(n6458), .A2(n6436), .B1(n6435), .B2(n6455), .ZN(n6439)
         );
  AOI22_X1 U7388 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6461), .B1(n6437), 
        .B2(n6459), .ZN(n6438) );
  OAI211_X1 U7389 ( .C1(n6440), .C2(n6464), .A(n6439), .B(n6438), .ZN(U3112)
         );
  AOI22_X1 U7390 ( .A1(n6449), .A2(n6442), .B1(n6441), .B2(n6455), .ZN(n6445)
         );
  AOI22_X1 U7391 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6461), .B1(n6443), 
        .B2(n6459), .ZN(n6444) );
  OAI211_X1 U7392 ( .C1(n6446), .C2(n6453), .A(n6445), .B(n6444), .ZN(U3113)
         );
  AOI22_X1 U7393 ( .A1(n6449), .A2(n6448), .B1(n6447), .B2(n6455), .ZN(n6452)
         );
  AOI22_X1 U7394 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6461), .B1(n6450), 
        .B2(n6459), .ZN(n6451) );
  OAI211_X1 U7395 ( .C1(n6454), .C2(n6453), .A(n6452), .B(n6451), .ZN(U3114)
         );
  AOI22_X1 U7396 ( .A1(n6458), .A2(n6457), .B1(n6456), .B2(n6455), .ZN(n6463)
         );
  AOI22_X1 U7397 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6461), .B1(n6460), 
        .B2(n6459), .ZN(n6462) );
  OAI211_X1 U7398 ( .C1(n6465), .C2(n6464), .A(n6463), .B(n6462), .ZN(U3115)
         );
  AND3_X1 U7399 ( .A1(n6467), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6466), 
        .ZN(n6471) );
  NAND2_X1 U7400 ( .A1(n6469), .A2(n6468), .ZN(n6470) );
  AOI222_X1 U7401 ( .A1(n6471), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n6471), .B2(n6470), .C1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n6470), 
        .ZN(n6472) );
  AOI222_X1 U7402 ( .A1(n6474), .A2(n6473), .B1(n6474), .B2(n6472), .C1(n6473), 
        .C2(n6472), .ZN(n6477) );
  OR2_X1 U7403 ( .A1(n6477), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6476)
         );
  NAND2_X1 U7404 ( .A1(n6476), .A2(n6475), .ZN(n6480) );
  NAND2_X1 U7405 ( .A1(n6477), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6479) );
  NAND3_X1 U7406 ( .A1(n6480), .A2(n6479), .A3(n6478), .ZN(n6490) );
  NOR2_X1 U7407 ( .A1(MORE_REG_SCAN_IN), .A2(FLUSH_REG_SCAN_IN), .ZN(n6482) );
  OAI21_X1 U7408 ( .B1(n6483), .B2(n6482), .A(n6481), .ZN(n6484) );
  OR3_X1 U7409 ( .A1(n6486), .A2(n6485), .A3(n6484), .ZN(n6487) );
  NOR2_X1 U7410 ( .A1(n6488), .A2(n6487), .ZN(n6489) );
  INV_X1 U7411 ( .A(n6497), .ZN(n6501) );
  NOR2_X1 U7412 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6606), .ZN(n6507) );
  NOR2_X1 U7413 ( .A1(n6507), .A2(n6491), .ZN(n6498) );
  INV_X1 U7414 ( .A(n6492), .ZN(n6496) );
  NAND3_X1 U7415 ( .A1(STATE2_REG_2__SCAN_IN), .A2(READY_N), .A3(n6509), .ZN(
        n6494) );
  AOI22_X1 U7416 ( .A1(n6496), .A2(n6495), .B1(n6494), .B2(n6493), .ZN(n6506)
         );
  OAI221_X1 U7417 ( .B1(STATE2_REG_1__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_1__SCAN_IN), .C2(n6497), .A(n6506), .ZN(n6587) );
  AOI21_X1 U7418 ( .B1(n6498), .B2(n6587), .A(n6509), .ZN(n6499) );
  AOI211_X1 U7419 ( .C1(n6511), .C2(n6501), .A(n6500), .B(n6499), .ZN(n6505)
         );
  OAI211_X1 U7420 ( .C1(n6503), .C2(n6502), .A(n6509), .B(n6587), .ZN(n6504)
         );
  NAND2_X1 U7421 ( .A1(n6505), .A2(n6504), .ZN(U3148) );
  AOI21_X1 U7422 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6507), .A(n6506), .ZN(
        n6514) );
  INV_X1 U7423 ( .A(n6508), .ZN(n6513) );
  NOR2_X1 U7424 ( .A1(READY_N), .A2(n6509), .ZN(n6515) );
  OAI221_X1 U7425 ( .B1(n6511), .B2(n6510), .C1(n6511), .C2(n6515), .A(n6587), 
        .ZN(n6512) );
  OAI211_X1 U7426 ( .C1(n6514), .C2(n6749), .A(n6513), .B(n6512), .ZN(U3149)
         );
  AOI21_X1 U7427 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n6515), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n6517) );
  OAI21_X1 U7428 ( .B1(n6518), .B2(n6517), .A(n6516), .ZN(U3150) );
  AND2_X1 U7429 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6581), .ZN(U3151) );
  INV_X1 U7430 ( .A(DATAWIDTH_REG_30__SCAN_IN), .ZN(n6737) );
  NOR2_X1 U7431 ( .A1(n6585), .A2(n6737), .ZN(U3152) );
  AND2_X1 U7432 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6581), .ZN(U3153) );
  AND2_X1 U7433 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6581), .ZN(U3154) );
  AND2_X1 U7434 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6581), .ZN(U3155) );
  AND2_X1 U7435 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6581), .ZN(U3156) );
  AND2_X1 U7436 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6581), .ZN(U3157) );
  AND2_X1 U7437 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6581), .ZN(U3158) );
  AND2_X1 U7438 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6581), .ZN(U3159) );
  AND2_X1 U7439 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6581), .ZN(U3160) );
  AND2_X1 U7440 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6581), .ZN(U3161) );
  INV_X1 U7441 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6684) );
  NOR2_X1 U7442 ( .A1(n6585), .A2(n6684), .ZN(U3162) );
  AND2_X1 U7443 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6581), .ZN(U3163) );
  AND2_X1 U7444 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6581), .ZN(U3164) );
  AND2_X1 U7445 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6581), .ZN(U3165) );
  AND2_X1 U7446 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6581), .ZN(U3166) );
  AND2_X1 U7447 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6581), .ZN(U3167) );
  AND2_X1 U7448 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6581), .ZN(U3168) );
  AND2_X1 U7449 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6581), .ZN(U3169) );
  AND2_X1 U7450 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6581), .ZN(U3170) );
  AND2_X1 U7451 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6581), .ZN(U3171) );
  AND2_X1 U7452 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6581), .ZN(U3172) );
  AND2_X1 U7453 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6581), .ZN(U3173) );
  AND2_X1 U7454 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6581), .ZN(U3174) );
  AND2_X1 U7455 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6581), .ZN(U3175) );
  AND2_X1 U7456 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6581), .ZN(U3176) );
  AND2_X1 U7457 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6581), .ZN(U3177) );
  AND2_X1 U7458 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6581), .ZN(U3178) );
  AND2_X1 U7459 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6581), .ZN(U3179) );
  AND2_X1 U7460 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6581), .ZN(U3180) );
  NOR2_X1 U7461 ( .A1(n6752), .A2(n6524), .ZN(n6520) );
  AOI22_X1 U7462 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6531) );
  AND2_X1 U7463 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6522) );
  INV_X1 U7464 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6614) );
  INV_X1 U7465 ( .A(NA_N), .ZN(n6525) );
  AOI221_X1 U7466 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6525), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6528) );
  AOI221_X1 U7467 ( .B1(n6522), .B2(n6579), .C1(n6614), .C2(n6579), .A(n6528), 
        .ZN(n6519) );
  OAI21_X1 U7468 ( .B1(n6520), .B2(n6531), .A(n6519), .ZN(U3181) );
  NOR2_X1 U7469 ( .A1(n4196), .A2(n6614), .ZN(n6526) );
  NAND2_X1 U7470 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6521) );
  OAI21_X1 U7471 ( .B1(n6526), .B2(n6522), .A(n6521), .ZN(n6523) );
  OAI211_X1 U7472 ( .C1(n6524), .C2(n6606), .A(n6603), .B(n6523), .ZN(U3182)
         );
  AOI22_X1 U7473 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .B1(
        n6526), .B2(n6525), .ZN(n6530) );
  AOI221_X1 U7474 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6606), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6527) );
  AOI221_X1 U7475 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6527), .C2(HOLD), .A(n4196), .ZN(n6529) );
  OAI22_X1 U7476 ( .A1(n6531), .A2(n6530), .B1(n6529), .B2(n6528), .ZN(U3183)
         );
  NAND2_X1 U7477 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6615), .ZN(n6573) );
  NOR2_X2 U7478 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6579), .ZN(n6567) );
  AOI22_X1 U7479 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6598), .ZN(n6532) );
  OAI21_X1 U7480 ( .B1(n6589), .B2(n6573), .A(n6532), .ZN(U3184) );
  AOI22_X1 U7481 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6575), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6598), .ZN(n6533) );
  OAI21_X1 U7482 ( .B1(n6658), .B2(n6577), .A(n6533), .ZN(U3185) );
  AOI22_X1 U7483 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6598), .ZN(n6534) );
  OAI21_X1 U7484 ( .B1(n6658), .B2(n6573), .A(n6534), .ZN(U3186) );
  AOI22_X1 U7485 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6598), .ZN(n6535) );
  OAI21_X1 U7486 ( .B1(n6740), .B2(n6573), .A(n6535), .ZN(U3187) );
  AOI22_X1 U7487 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6575), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6598), .ZN(n6536) );
  OAI21_X1 U7488 ( .B1(n6538), .B2(n6577), .A(n6536), .ZN(U3188) );
  AOI22_X1 U7489 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6598), .ZN(n6537) );
  OAI21_X1 U7490 ( .B1(n6538), .B2(n6573), .A(n6537), .ZN(U3189) );
  AOI22_X1 U7491 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6575), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6598), .ZN(n6539) );
  OAI21_X1 U7492 ( .B1(n6541), .B2(n6577), .A(n6539), .ZN(U3190) );
  AOI22_X1 U7493 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6598), .ZN(n6540) );
  OAI21_X1 U7494 ( .B1(n6541), .B2(n6573), .A(n6540), .ZN(U3191) );
  INV_X1 U7495 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6723) );
  OAI222_X1 U7496 ( .A1(n6573), .A2(n6543), .B1(n6723), .B2(n6615), .C1(n6542), 
        .C2(n6577), .ZN(U3192) );
  AOI22_X1 U7497 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6575), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6579), .ZN(n6544) );
  OAI21_X1 U7498 ( .B1(n6674), .B2(n6577), .A(n6544), .ZN(U3193) );
  AOI22_X1 U7499 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6598), .ZN(n6545) );
  OAI21_X1 U7500 ( .B1(n6674), .B2(n6573), .A(n6545), .ZN(U3194) );
  AOI22_X1 U7501 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6598), .ZN(n6546) );
  OAI21_X1 U7502 ( .B1(n6784), .B2(n6573), .A(n6546), .ZN(U3195) );
  INV_X1 U7503 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6548) );
  AOI22_X1 U7504 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6598), .ZN(n6547) );
  OAI21_X1 U7505 ( .B1(n6548), .B2(n6573), .A(n6547), .ZN(U3196) );
  AOI22_X1 U7506 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6575), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6598), .ZN(n6549) );
  OAI21_X1 U7507 ( .B1(n6551), .B2(n6577), .A(n6549), .ZN(U3197) );
  AOI22_X1 U7508 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6598), .ZN(n6550) );
  OAI21_X1 U7509 ( .B1(n6551), .B2(n6573), .A(n6550), .ZN(U3198) );
  AOI22_X1 U7510 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6575), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6598), .ZN(n6552) );
  OAI21_X1 U7511 ( .B1(n6554), .B2(n6577), .A(n6552), .ZN(U3199) );
  AOI22_X1 U7512 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6598), .ZN(n6553) );
  OAI21_X1 U7513 ( .B1(n6554), .B2(n6573), .A(n6553), .ZN(U3200) );
  INV_X1 U7514 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6557) );
  AOI22_X1 U7515 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6575), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6598), .ZN(n6555) );
  OAI21_X1 U7516 ( .B1(n6557), .B2(n6577), .A(n6555), .ZN(U3201) );
  AOI22_X1 U7517 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6598), .ZN(n6556) );
  OAI21_X1 U7518 ( .B1(n6557), .B2(n6573), .A(n6556), .ZN(U3202) );
  AOI22_X1 U7519 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6575), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6598), .ZN(n6558) );
  OAI21_X1 U7520 ( .B1(n6670), .B2(n6577), .A(n6558), .ZN(U3203) );
  INV_X1 U7521 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6561) );
  AOI22_X1 U7522 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6575), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6579), .ZN(n6559) );
  OAI21_X1 U7523 ( .B1(n6561), .B2(n6577), .A(n6559), .ZN(U3204) );
  AOI22_X1 U7524 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6579), .ZN(n6560) );
  OAI21_X1 U7525 ( .B1(n6561), .B2(n6573), .A(n6560), .ZN(U3205) );
  AOI22_X1 U7526 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6575), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6579), .ZN(n6562) );
  OAI21_X1 U7527 ( .B1(n6564), .B2(n6577), .A(n6562), .ZN(U3206) );
  AOI22_X1 U7528 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6598), .ZN(n6563) );
  OAI21_X1 U7529 ( .B1(n6564), .B2(n6573), .A(n6563), .ZN(U3207) );
  AOI22_X1 U7530 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6579), .ZN(n6565) );
  OAI21_X1 U7531 ( .B1(n6566), .B2(n6573), .A(n6565), .ZN(U3208) );
  AOI22_X1 U7532 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6579), .ZN(n6568) );
  OAI21_X1 U7533 ( .B1(n6569), .B2(n6573), .A(n6568), .ZN(U3209) );
  INV_X1 U7534 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6572) );
  AOI22_X1 U7535 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6575), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6579), .ZN(n6570) );
  OAI21_X1 U7536 ( .B1(n6572), .B2(n6577), .A(n6570), .ZN(U3210) );
  INV_X1 U7537 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6690) );
  OAI222_X1 U7538 ( .A1(n6573), .A2(n6572), .B1(n6690), .B2(n6615), .C1(n6571), 
        .C2(n6577), .ZN(U3211) );
  AOI22_X1 U7539 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6575), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6579), .ZN(n6574) );
  OAI21_X1 U7540 ( .B1(n6660), .B2(n6577), .A(n6574), .ZN(U3212) );
  INV_X1 U7541 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6578) );
  AOI22_X1 U7542 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6575), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6579), .ZN(n6576) );
  OAI21_X1 U7543 ( .B1(n6578), .B2(n6577), .A(n6576), .ZN(U3213) );
  INV_X1 U7544 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n6709) );
  AOI22_X1 U7545 ( .A1(n6615), .A2(n6683), .B1(n6709), .B2(n6579), .ZN(U3445)
         );
  MUX2_X1 U7546 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6615), .Z(U3446) );
  MUX2_X1 U7547 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6615), .Z(U3447) );
  MUX2_X1 U7548 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6615), .Z(U3448) );
  INV_X1 U7549 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6582) );
  INV_X1 U7550 ( .A(n6583), .ZN(n6580) );
  AOI21_X1 U7551 ( .B1(n6582), .B2(n6581), .A(n6580), .ZN(U3451) );
  OAI21_X1 U7552 ( .B1(n6585), .B2(n6584), .A(n6583), .ZN(U3452) );
  OAI221_X1 U7553 ( .B1(n6588), .B2(STATE2_REG_0__SCAN_IN), .C1(n6588), .C2(
        n6587), .A(n6586), .ZN(U3453) );
  AOI21_X1 U7554 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6590) );
  AOI22_X1 U7555 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6590), .B2(n6589), .ZN(n6593) );
  INV_X1 U7556 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6592) );
  AOI22_X1 U7557 ( .A1(n6596), .A2(n6593), .B1(n6592), .B2(n6591), .ZN(U3468)
         );
  INV_X1 U7558 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6595) );
  OAI21_X1 U7559 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6596), .ZN(n6594) );
  OAI21_X1 U7560 ( .B1(n6596), .B2(n6595), .A(n6594), .ZN(U3469) );
  NAND2_X1 U7561 ( .A1(n6598), .A2(W_R_N_REG_SCAN_IN), .ZN(n6597) );
  OAI21_X1 U7562 ( .B1(n6598), .B2(READREQUEST_REG_SCAN_IN), .A(n6597), .ZN(
        U3470) );
  AOI211_X1 U7563 ( .C1(n6601), .C2(n6606), .A(n6600), .B(n6599), .ZN(n6613)
         );
  INV_X1 U7564 ( .A(n6602), .ZN(n6608) );
  AOI21_X1 U7565 ( .B1(n6605), .B2(n6604), .A(n6603), .ZN(n6607) );
  OAI211_X1 U7566 ( .C1(n6608), .C2(n6607), .A(STATE2_REG_2__SCAN_IN), .B(
        n6606), .ZN(n6609) );
  NAND2_X1 U7567 ( .A1(n6609), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6612) );
  NOR2_X1 U7568 ( .A1(n6613), .A2(n6610), .ZN(n6611) );
  AOI22_X1 U7569 ( .A1(n6614), .A2(n6613), .B1(n6612), .B2(n6611), .ZN(U3472)
         );
  MUX2_X1 U7570 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6615), .Z(U3473) );
  NAND4_X1 U7571 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(
        INSTQUEUE_REG_12__0__SCAN_IN), .A3(PHYADDRPOINTER_REG_20__SCAN_IN), 
        .A4(DATAO_REG_1__SCAN_IN), .ZN(n6625) );
  NOR4_X1 U7572 ( .A1(EBX_REG_11__SCAN_IN), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .A3(ADDRESS_REG_8__SCAN_IN), .A4(UWORD_REG_0__SCAN_IN), .ZN(n6618) );
  NOR4_X1 U7573 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(EAX_REG_20__SCAN_IN), 
        .A3(n6707), .A4(n6703), .ZN(n6617) );
  INV_X1 U7574 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n6712) );
  NOR3_X1 U7575 ( .A1(BS16_N), .A2(n6710), .A3(n6712), .ZN(n6616) );
  NAND4_X1 U7576 ( .A1(n6618), .A2(n6617), .A3(BE_N_REG_3__SCAN_IN), .A4(n6616), .ZN(n6624) );
  NAND4_X1 U7577 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        DATAWIDTH_REG_30__SCAN_IN), .A3(n6735), .A4(n6734), .ZN(n6623) );
  NOR4_X1 U7578 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(REIP_REG_4__SCAN_IN), 
        .A3(DATAO_REG_14__SCAN_IN), .A4(n6743), .ZN(n6621) );
  NOR4_X1 U7579 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .A3(PHYADDRPOINTER_REG_19__SCAN_IN), 
        .A4(n6750), .ZN(n6619) );
  AND3_X1 U7580 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(DATAI_15_), .A3(n6619), 
        .ZN(n6620) );
  NAND4_X1 U7581 ( .A1(n6621), .A2(n6620), .A3(n6752), .A4(n6757), .ZN(n6622)
         );
  NOR4_X1 U7582 ( .A1(n6625), .A2(n6624), .A3(n6623), .A4(n6622), .ZN(n6771)
         );
  NAND4_X1 U7583 ( .A1(REIP_REG_3__SCAN_IN), .A2(REIP_REG_30__SCAN_IN), .A3(
        LWORD_REG_7__SCAN_IN), .A4(n6657), .ZN(n6635) );
  NOR4_X1 U7584 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n6640), .A4(n6641), .ZN(n6628) );
  NOR4_X1 U7585 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(
        INSTQUEUE_REG_13__0__SCAN_IN), .A3(UWORD_REG_8__SCAN_IN), .A4(n6638), 
        .ZN(n6627) );
  NOR3_X1 U7586 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(
        INSTQUEUE_REG_10__2__SCAN_IN), .A3(EBX_REG_19__SCAN_IN), .ZN(n6626) );
  NAND4_X1 U7587 ( .A1(EAX_REG_29__SCAN_IN), .A2(n6628), .A3(n6627), .A4(n6626), .ZN(n6634) );
  NAND4_X1 U7588 ( .A1(EBX_REG_7__SCAN_IN), .A2(ADDRESS_REG_27__SCAN_IN), .A3(
        DATAO_REG_18__SCAN_IN), .A4(n6692), .ZN(n6633) );
  NOR4_X1 U7589 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(DATAI_19_), .A3(
        n6670), .A4(n6667), .ZN(n6631) );
  NOR4_X1 U7590 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .A3(REIP_REG_11__SCAN_IN), .A4(
        LWORD_REG_6__SCAN_IN), .ZN(n6630) );
  NOR3_X1 U7591 ( .A1(DATAI_24_), .A2(BYTEENABLE_REG_3__SCAN_IN), .A3(n6684), 
        .ZN(n6629) );
  NAND4_X1 U7592 ( .A1(DATAI_29_), .A2(n6631), .A3(n6630), .A4(n6629), .ZN(
        n6632) );
  NOR4_X1 U7593 ( .A1(n6635), .A2(n6634), .A3(n6633), .A4(n6632), .ZN(n6770)
         );
  AOI22_X1 U7594 ( .A1(n6638), .A2(keyinput16), .B1(keyinput28), .B2(n6637), 
        .ZN(n6636) );
  OAI221_X1 U7595 ( .B1(n6638), .B2(keyinput16), .C1(n6637), .C2(keyinput28), 
        .A(n6636), .ZN(n6649) );
  AOI22_X1 U7596 ( .A1(n6641), .A2(keyinput42), .B1(n6640), .B2(keyinput47), 
        .ZN(n6639) );
  OAI221_X1 U7597 ( .B1(n6641), .B2(keyinput42), .C1(n6640), .C2(keyinput47), 
        .A(n6639), .ZN(n6648) );
  INV_X1 U7598 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n6642) );
  XOR2_X1 U7599 ( .A(n6642), .B(keyinput14), .Z(n6646) );
  XNOR2_X1 U7600 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .B(keyinput5), .ZN(n6645)
         );
  XNOR2_X1 U7601 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .B(keyinput22), .ZN(
        n6644) );
  XNOR2_X1 U7602 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .B(keyinput38), .ZN(n6643) );
  NAND4_X1 U7603 ( .A1(n6646), .A2(n6645), .A3(n6644), .A4(n6643), .ZN(n6647)
         );
  NOR3_X1 U7604 ( .A1(n6649), .A2(n6648), .A3(n6647), .ZN(n6701) );
  AOI22_X1 U7605 ( .A1(n6652), .A2(keyinput59), .B1(n6651), .B2(keyinput45), 
        .ZN(n6650) );
  OAI221_X1 U7606 ( .B1(n6652), .B2(keyinput59), .C1(n6651), .C2(keyinput45), 
        .A(n6650), .ZN(n6665) );
  INV_X1 U7607 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6654) );
  AOI22_X1 U7608 ( .A1(n6655), .A2(keyinput63), .B1(n6654), .B2(keyinput29), 
        .ZN(n6653) );
  OAI221_X1 U7609 ( .B1(n6655), .B2(keyinput63), .C1(n6654), .C2(keyinput29), 
        .A(n6653), .ZN(n6664) );
  AOI22_X1 U7610 ( .A1(n6658), .A2(keyinput7), .B1(keyinput19), .B2(n6657), 
        .ZN(n6656) );
  OAI221_X1 U7611 ( .B1(n6658), .B2(keyinput7), .C1(n6657), .C2(keyinput19), 
        .A(n6656), .ZN(n6663) );
  AOI22_X1 U7612 ( .A1(n6661), .A2(keyinput33), .B1(n6660), .B2(keyinput58), 
        .ZN(n6659) );
  OAI221_X1 U7613 ( .B1(n6661), .B2(keyinput33), .C1(n6660), .C2(keyinput58), 
        .A(n6659), .ZN(n6662) );
  NOR4_X1 U7614 ( .A1(n6665), .A2(n6664), .A3(n6663), .A4(n6662), .ZN(n6700)
         );
  AOI22_X1 U7615 ( .A1(n6668), .A2(keyinput55), .B1(keyinput12), .B2(n6667), 
        .ZN(n6666) );
  OAI221_X1 U7616 ( .B1(n6668), .B2(keyinput55), .C1(n6667), .C2(keyinput12), 
        .A(n6666), .ZN(n6681) );
  INV_X1 U7617 ( .A(DATAI_19_), .ZN(n6671) );
  AOI22_X1 U7618 ( .A1(n6671), .A2(keyinput31), .B1(n6670), .B2(keyinput1), 
        .ZN(n6669) );
  OAI221_X1 U7619 ( .B1(n6671), .B2(keyinput31), .C1(n6670), .C2(keyinput1), 
        .A(n6669), .ZN(n6680) );
  AOI22_X1 U7620 ( .A1(n6674), .A2(keyinput34), .B1(n6673), .B2(keyinput41), 
        .ZN(n6672) );
  OAI221_X1 U7621 ( .B1(n6674), .B2(keyinput34), .C1(n6673), .C2(keyinput41), 
        .A(n6672), .ZN(n6679) );
  INV_X1 U7622 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6677) );
  AOI22_X1 U7623 ( .A1(n6677), .A2(keyinput17), .B1(keyinput4), .B2(n6676), 
        .ZN(n6675) );
  OAI221_X1 U7624 ( .B1(n6677), .B2(keyinput17), .C1(n6676), .C2(keyinput4), 
        .A(n6675), .ZN(n6678) );
  NOR4_X1 U7625 ( .A1(n6681), .A2(n6680), .A3(n6679), .A4(n6678), .ZN(n6699)
         );
  AOI22_X1 U7626 ( .A1(n6684), .A2(keyinput54), .B1(keyinput6), .B2(n6683), 
        .ZN(n6682) );
  OAI221_X1 U7627 ( .B1(n6684), .B2(keyinput54), .C1(n6683), .C2(keyinput6), 
        .A(n6682), .ZN(n6697) );
  INV_X1 U7628 ( .A(DATAI_29_), .ZN(n6687) );
  INV_X1 U7629 ( .A(DATAI_24_), .ZN(n6686) );
  AOI22_X1 U7630 ( .A1(n6687), .A2(keyinput3), .B1(keyinput57), .B2(n6686), 
        .ZN(n6685) );
  OAI221_X1 U7631 ( .B1(n6687), .B2(keyinput3), .C1(n6686), .C2(keyinput57), 
        .A(n6685), .ZN(n6696) );
  AOI22_X1 U7632 ( .A1(n6690), .A2(keyinput11), .B1(keyinput49), .B2(n6689), 
        .ZN(n6688) );
  OAI221_X1 U7633 ( .B1(n6690), .B2(keyinput11), .C1(n6689), .C2(keyinput49), 
        .A(n6688), .ZN(n6695) );
  AOI22_X1 U7634 ( .A1(n6693), .A2(keyinput48), .B1(keyinput13), .B2(n6692), 
        .ZN(n6691) );
  OAI221_X1 U7635 ( .B1(n6693), .B2(keyinput48), .C1(n6692), .C2(keyinput13), 
        .A(n6691), .ZN(n6694) );
  NOR4_X1 U7636 ( .A1(n6697), .A2(n6696), .A3(n6695), .A4(n6694), .ZN(n6698)
         );
  NAND4_X1 U7637 ( .A1(n6701), .A2(n6700), .A3(n6699), .A4(n6698), .ZN(n6769)
         );
  AOI22_X1 U7638 ( .A1(n6704), .A2(keyinput40), .B1(n6703), .B2(keyinput53), 
        .ZN(n6702) );
  OAI221_X1 U7639 ( .B1(n6704), .B2(keyinput40), .C1(n6703), .C2(keyinput53), 
        .A(n6702), .ZN(n6717) );
  AOI22_X1 U7640 ( .A1(n6707), .A2(keyinput21), .B1(keyinput2), .B2(n6706), 
        .ZN(n6705) );
  OAI221_X1 U7641 ( .B1(n6707), .B2(keyinput21), .C1(n6706), .C2(keyinput2), 
        .A(n6705), .ZN(n6716) );
  AOI22_X1 U7642 ( .A1(n6710), .A2(keyinput51), .B1(keyinput39), .B2(n6709), 
        .ZN(n6708) );
  OAI221_X1 U7643 ( .B1(n6710), .B2(keyinput51), .C1(n6709), .C2(keyinput39), 
        .A(n6708), .ZN(n6715) );
  INV_X1 U7644 ( .A(BS16_N), .ZN(n6713) );
  AOI22_X1 U7645 ( .A1(n6713), .A2(keyinput52), .B1(n6712), .B2(keyinput56), 
        .ZN(n6711) );
  OAI221_X1 U7646 ( .B1(n6713), .B2(keyinput52), .C1(n6712), .C2(keyinput56), 
        .A(n6711), .ZN(n6714) );
  NOR4_X1 U7647 ( .A1(n6717), .A2(n6716), .A3(n6715), .A4(n6714), .ZN(n6767)
         );
  AOI22_X1 U7648 ( .A1(n6720), .A2(keyinput43), .B1(keyinput18), .B2(n6719), 
        .ZN(n6718) );
  OAI221_X1 U7649 ( .B1(n6720), .B2(keyinput43), .C1(n6719), .C2(keyinput18), 
        .A(n6718), .ZN(n6732) );
  INV_X1 U7650 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6722) );
  AOI22_X1 U7651 ( .A1(n6723), .A2(keyinput20), .B1(n6722), .B2(keyinput36), 
        .ZN(n6721) );
  OAI221_X1 U7652 ( .B1(n6723), .B2(keyinput20), .C1(n6722), .C2(keyinput36), 
        .A(n6721), .ZN(n6731) );
  INV_X1 U7653 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n6726) );
  AOI22_X1 U7654 ( .A1(n6726), .A2(keyinput46), .B1(keyinput27), .B2(n6725), 
        .ZN(n6724) );
  OAI221_X1 U7655 ( .B1(n6726), .B2(keyinput46), .C1(n6725), .C2(keyinput27), 
        .A(n6724), .ZN(n6730) );
  INV_X1 U7656 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n6728) );
  AOI22_X1 U7657 ( .A1(n5210), .A2(keyinput15), .B1(n6728), .B2(keyinput23), 
        .ZN(n6727) );
  OAI221_X1 U7658 ( .B1(n5210), .B2(keyinput15), .C1(n6728), .C2(keyinput23), 
        .A(n6727), .ZN(n6729) );
  NOR4_X1 U7659 ( .A1(n6732), .A2(n6731), .A3(n6730), .A4(n6729), .ZN(n6766)
         );
  AOI22_X1 U7660 ( .A1(n6735), .A2(keyinput60), .B1(keyinput9), .B2(n6734), 
        .ZN(n6733) );
  OAI221_X1 U7661 ( .B1(n6735), .B2(keyinput60), .C1(n6734), .C2(keyinput9), 
        .A(n6733), .ZN(n6747) );
  AOI22_X1 U7662 ( .A1(n6737), .A2(keyinput32), .B1(n3762), .B2(keyinput30), 
        .ZN(n6736) );
  OAI221_X1 U7663 ( .B1(n6737), .B2(keyinput32), .C1(n3762), .C2(keyinput30), 
        .A(n6736), .ZN(n6746) );
  AOI22_X1 U7664 ( .A1(n6740), .A2(keyinput0), .B1(keyinput35), .B2(n6739), 
        .ZN(n6738) );
  OAI221_X1 U7665 ( .B1(n6740), .B2(keyinput0), .C1(n6739), .C2(keyinput35), 
        .A(n6738), .ZN(n6745) );
  INV_X1 U7666 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6742) );
  AOI22_X1 U7667 ( .A1(n6743), .A2(keyinput37), .B1(n6742), .B2(keyinput26), 
        .ZN(n6741) );
  OAI221_X1 U7668 ( .B1(n6743), .B2(keyinput37), .C1(n6742), .C2(keyinput26), 
        .A(n6741), .ZN(n6744) );
  NOR4_X1 U7669 ( .A1(n6747), .A2(n6746), .A3(n6745), .A4(n6744), .ZN(n6765)
         );
  AOI22_X1 U7670 ( .A1(n6750), .A2(keyinput61), .B1(n6749), .B2(keyinput8), 
        .ZN(n6748) );
  OAI221_X1 U7671 ( .B1(n6750), .B2(keyinput61), .C1(n6749), .C2(keyinput8), 
        .A(n6748), .ZN(n6763) );
  AOI22_X1 U7672 ( .A1(n6753), .A2(keyinput10), .B1(n6752), .B2(keyinput44), 
        .ZN(n6751) );
  OAI221_X1 U7673 ( .B1(n6753), .B2(keyinput10), .C1(n6752), .C2(keyinput44), 
        .A(n6751), .ZN(n6762) );
  AOI22_X1 U7674 ( .A1(n6756), .A2(keyinput25), .B1(keyinput24), .B2(n6755), 
        .ZN(n6754) );
  OAI221_X1 U7675 ( .B1(n6756), .B2(keyinput25), .C1(n6755), .C2(keyinput24), 
        .A(n6754), .ZN(n6761) );
  XOR2_X1 U7676 ( .A(n6757), .B(keyinput62), .Z(n6759) );
  XNOR2_X1 U7677 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .B(keyinput50), .ZN(n6758)
         );
  NAND2_X1 U7678 ( .A1(n6759), .A2(n6758), .ZN(n6760) );
  NOR4_X1 U7679 ( .A1(n6763), .A2(n6762), .A3(n6761), .A4(n6760), .ZN(n6764)
         );
  NAND4_X1 U7680 ( .A1(n6767), .A2(n6766), .A3(n6765), .A4(n6764), .ZN(n6768)
         );
  AOI211_X1 U7681 ( .C1(n6771), .C2(n6770), .A(n6769), .B(n6768), .ZN(n6793)
         );
  INV_X1 U7682 ( .A(n6772), .ZN(n6788) );
  INV_X1 U7683 ( .A(n6773), .ZN(n6774) );
  NAND3_X1 U7684 ( .A1(n6775), .A2(n6784), .A3(n6774), .ZN(n6776) );
  OAI21_X1 U7685 ( .B1(n6778), .B2(n6777), .A(n6776), .ZN(n6786) );
  AOI22_X1 U7686 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6780), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6779), .ZN(n6782) );
  OAI211_X1 U7687 ( .C1(n6784), .C2(n6783), .A(n6782), .B(n6781), .ZN(n6785)
         );
  AOI211_X1 U7688 ( .C1(n6788), .C2(n6787), .A(n6786), .B(n6785), .ZN(n6789)
         );
  OAI21_X1 U7689 ( .B1(n6791), .B2(n6790), .A(n6789), .ZN(n6792) );
  XOR2_X1 U7690 ( .A(n6793), .B(n6792), .Z(U2815) );
  NAND2_X1 U3420 ( .A1(n4681), .A2(n3253), .ZN(n5297) );
  BUF_X2 U3932 ( .A(n3340), .Z(n4288) );
  NAND2_X1 U3707 ( .A1(n3452), .A2(n3451), .ZN(n3893) );
  CLKBUF_X1 U3441 ( .A(n3385), .Z(n3446) );
  CLKBUF_X1 U3533 ( .A(n3284), .Z(n4212) );
  CLKBUF_X1 U3583 ( .A(n3381), .Z(n3299) );
  CLKBUF_X1 U4357 ( .A(n3289), .Z(n3685) );
  OAI21_X1 U4429 ( .B1(n5188), .B2(n5187), .A(n3149), .ZN(n5190) );
endmodule

