

module b14_C_gen_AntiSAT_k_128_10 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, 
        U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, 
        U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, 
        U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, 
        U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, 
        U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, 
        U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, 
        U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, 
        U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, 
        U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, 
        U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, 
        U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, 
        U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, 
        U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, 
        U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, 
        U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, 
        U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, 
        U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, 
        U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, 
        U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, 
        U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, 
        U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, 
        U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, 
        U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, 
        U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737;

  INV_X1 U2285 ( .A(n3602), .ZN(n3591) );
  CLKBUF_X2 U2286 ( .A(n2433), .Z(n2471) );
  INV_X1 U2288 ( .A(n3601), .ZN(n2857) );
  INV_X2 U2289 ( .A(n2878), .ZN(n3600) );
  OAI21_X1 U2290 ( .B1(n3262), .B2(n2189), .A(n2186), .ZN(n3427) );
  INV_X1 U2291 ( .A(n2401), .ZN(n2455) );
  NAND2_X1 U2292 ( .A1(n2687), .A2(IR_REG_31__SCAN_IN), .ZN(n2689) );
  AND4_X1 U2293 ( .A1(n2438), .A2(n2437), .A3(n2436), .A4(n2435), .ZN(n2978)
         );
  NOR2_X2 U2294 ( .A1(n3470), .A2(n4344), .ZN(n3469) );
  NAND2_X1 U2295 ( .A1(n2329), .A2(IR_REG_31__SCAN_IN), .ZN(n2312) );
  NOR2_X1 U2296 ( .A1(n2250), .A2(n2249), .ZN(n4415) );
  OAI22_X2 U2297 ( .A1(n3227), .A2(n2520), .B1(n3388), .B2(n3309), .ZN(n3286)
         );
  OAI21_X2 U2298 ( .B1(n3185), .B2(n2509), .A(n2510), .ZN(n3227) );
  XNOR2_X2 U2299 ( .A(n2689), .B(n2688), .ZN(n2691) );
  XNOR2_X2 U2300 ( .A(n2312), .B(IR_REG_24__SCAN_IN), .ZN(n2729) );
  XNOR2_X2 U2301 ( .A(n2399), .B(IR_REG_29__SCAN_IN), .ZN(n3497) );
  OR2_X2 U2302 ( .A1(n2398), .A2(n3493), .ZN(n2399) );
  NAND2_X1 U2303 ( .A1(n2121), .A2(n2671), .ZN(n3615) );
  AND2_X1 U2304 ( .A1(n2206), .A2(n2062), .ZN(n3149) );
  INV_X1 U2306 ( .A(n2875), .ZN(n2856) );
  INV_X1 U2307 ( .A(n3962), .ZN(n3178) );
  NAND4_X1 U2308 ( .A1(n2475), .A2(n2474), .A3(n2473), .A4(n2472), .ZN(n4253)
         );
  NAND4_X1 U2309 ( .A1(n2462), .A2(n2461), .A3(n2460), .A4(n2459), .ZN(n3962)
         );
  CLKBUF_X2 U2310 ( .A(n2434), .Z(n2401) );
  INV_X1 U2311 ( .A(n4227), .ZN(n4011) );
  AND2_X1 U2312 ( .A1(n3726), .A2(n3648), .ZN(n3727) );
  OR2_X1 U2313 ( .A1(n3667), .A2(n3647), .ZN(n3726) );
  AOI21_X1 U2314 ( .B1(n3615), .B2(n3614), .A(n2214), .ZN(n2686) );
  INV_X1 U2315 ( .A(n2207), .ZN(n2205) );
  AND2_X1 U2316 ( .A1(n3117), .A2(n3116), .ZN(n3121) );
  AND2_X1 U2317 ( .A1(n3810), .A2(n3814), .ZN(n3893) );
  INV_X1 U2318 ( .A(n3895), .ZN(n2763) );
  NAND2_X2 U2319 ( .A1(n2856), .A2(n3107), .ZN(n3601) );
  AND2_X1 U2320 ( .A1(n3800), .A2(n3803), .ZN(n3895) );
  INV_X1 U2321 ( .A(n3961), .ZN(n3221) );
  NAND3_X1 U2322 ( .A1(n2450), .A2(n2449), .A3(n2448), .ZN(n3963) );
  INV_X1 U2323 ( .A(n3049), .ZN(n2043) );
  INV_X2 U2324 ( .A(n3049), .ZN(n2878) );
  NAND2_X1 U2325 ( .A1(n2871), .A2(n2858), .ZN(n2875) );
  NAND2_X1 U2326 ( .A1(n2469), .A2(n2050), .ZN(n3961) );
  NAND2_X1 U2327 ( .A1(n2847), .A2(n2858), .ZN(n3049) );
  AND2_X1 U2328 ( .A1(n2442), .A2(n2441), .ZN(n2450) );
  NAND3_X1 U2329 ( .A1(n2729), .A2(n2788), .A3(n4408), .ZN(n2858) );
  NAND2_X2 U2330 ( .A1(n2871), .A2(n2870), .ZN(n3602) );
  OAI21_X1 U2331 ( .B1(n2609), .B2(n2477), .A(n2476), .ZN(n2995) );
  INV_X1 U2332 ( .A(n3218), .ZN(n3101) );
  AND2_X1 U2333 ( .A1(n2321), .A2(n2323), .ZN(n2788) );
  NAND2_X1 U2334 ( .A1(n2609), .A2(n4414), .ZN(n2476) );
  AND2_X1 U2335 ( .A1(n2608), .A2(n2687), .ZN(n4227) );
  AND2_X1 U2336 ( .A1(n2325), .A2(n2324), .ZN(n4408) );
  NAND2_X1 U2337 ( .A1(n2342), .A2(n2340), .ZN(n2345) );
  OR2_X1 U2338 ( .A1(n2323), .A2(n2210), .ZN(n2342) );
  AND4_X1 U2339 ( .A1(n2307), .A2(n2306), .A3(n2305), .A4(n2304), .ZN(n2308)
         );
  NAND2_X1 U2340 ( .A1(n2338), .A2(n2211), .ZN(n2210) );
  NAND3_X1 U2341 ( .A1(n2079), .A2(n2259), .A3(n2222), .ZN(n2239) );
  INV_X1 U2342 ( .A(IR_REG_3__SCAN_IN), .ZN(n2259) );
  NOR2_X1 U2343 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2225)
         );
  NOR2_X1 U2344 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_2__SCAN_IN), .ZN(n2222)
         );
  NOR2_X1 U2345 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2226)
         );
  NOR2_X1 U2346 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2224)
         );
  NOR2_X1 U2347 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2223)
         );
  NOR2_X2 U2348 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2079)
         );
  INV_X1 U2349 ( .A(IR_REG_14__SCAN_IN), .ZN(n2236) );
  INV_X1 U2350 ( .A(IR_REG_15__SCAN_IN), .ZN(n2297) );
  AND3_X2 U2351 ( .A1(n2582), .A2(n2581), .A3(n2580), .ZN(n4338) );
  NOR2_X2 U2352 ( .A1(n2239), .A2(n2078), .ZN(n2309) );
  AOI21_X4 U2353 ( .B1(n3175), .B2(n3174), .A(n2064), .ZN(n3262) );
  INV_X2 U2354 ( .A(n3779), .ZN(n2609) );
  AND3_X1 U2355 ( .A1(n2318), .A2(n2317), .A3(n2316), .ZN(n2319) );
  NOR2_X1 U2356 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2317)
         );
  INV_X1 U2357 ( .A(n2124), .ZN(n2123) );
  OAI22_X1 U2358 ( .A1(n2063), .A2(n2647), .B1(n4132), .B2(n4112), .ZN(n2124)
         );
  INV_X1 U2359 ( .A(n3499), .ZN(n2202) );
  NAND2_X1 U2360 ( .A1(n3501), .A2(n2202), .ZN(n2200) );
  AND2_X1 U2361 ( .A1(n4411), .A2(n4510), .ZN(n2119) );
  INV_X1 U2362 ( .A(n3779), .ZN(n3780) );
  INV_X1 U2363 ( .A(n2079), .ZN(n2252) );
  NAND2_X1 U2364 ( .A1(n2392), .A2(REG3_REG_23__SCAN_IN), .ZN(n2649) );
  INV_X1 U2365 ( .A(n2639), .ZN(n2392) );
  OAI22_X1 U2366 ( .A1(n2880), .A2(n3049), .B1(n2876), .B2(n2875), .ZN(n2877)
         );
  OR2_X1 U2367 ( .A1(n4411), .A2(n4510), .ZN(n2120) );
  NOR2_X1 U2368 ( .A1(n2117), .A2(n2119), .ZN(n2116) );
  INV_X1 U2369 ( .A(n4432), .ZN(n2117) );
  XNOR2_X1 U2370 ( .A(n2285), .B(n2284), .ZN(n4445) );
  NAND2_X1 U2371 ( .A1(n4454), .A2(n4455), .ZN(n4453) );
  XNOR2_X1 U2372 ( .A(n2289), .B(n2288), .ZN(n4467) );
  AND2_X1 U2373 ( .A1(n2380), .A2(n2375), .ZN(n2156) );
  OR2_X1 U2374 ( .A1(n2661), .A2(n3751), .ZN(n2663) );
  OAI21_X1 U2375 ( .B1(n4158), .B2(n2628), .A(n2627), .ZN(n4147) );
  INV_X1 U2376 ( .A(n2139), .ZN(n2138) );
  AOI21_X1 U2377 ( .B1(n2139), .B2(n2137), .A(n2059), .ZN(n2136) );
  AOI21_X1 U2378 ( .B1(n3894), .B2(n2530), .A(n2052), .ZN(n2139) );
  NAND2_X1 U2379 ( .A1(n2691), .A2(n3006), .ZN(n3107) );
  INV_X2 U2380 ( .A(n2439), .ZN(n3779) );
  NAND2_X1 U2381 ( .A1(n2402), .A2(n3497), .ZN(n2433) );
  NOR2_X1 U2382 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2306)
         );
  NOR2_X1 U2383 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2305)
         );
  NOR2_X1 U2384 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2304)
         );
  INV_X1 U2385 ( .A(n2210), .ZN(n2209) );
  INV_X1 U2386 ( .A(n2555), .ZN(n2131) );
  INV_X1 U2387 ( .A(n3306), .ZN(n2190) );
  INV_X1 U2388 ( .A(n3261), .ZN(n2195) );
  INV_X1 U2389 ( .A(n3381), .ZN(n3382) );
  NOR2_X1 U2390 ( .A1(n3533), .A2(n2169), .ZN(n2168) );
  INV_X1 U2391 ( .A(n3525), .ZN(n2169) );
  NOR2_X1 U2392 ( .A1(n3532), .A2(n3531), .ZN(n2166) );
  OAI21_X1 U2393 ( .B1(n3500), .B2(n2199), .A(n2198), .ZN(n3685) );
  AOI21_X1 U2394 ( .B1(n2200), .B2(n2201), .A(n2070), .ZN(n2198) );
  NAND2_X1 U2395 ( .A1(n2111), .A2(n2110), .ZN(n2109) );
  NAND2_X1 U2396 ( .A1(n4415), .A2(REG2_REG_2__SCAN_IN), .ZN(n2110) );
  AND2_X1 U2397 ( .A1(n2700), .A2(n2048), .ZN(n2088) );
  NAND2_X1 U2398 ( .A1(n2556), .A2(REG3_REG_16__SCAN_IN), .ZN(n2583) );
  OAI21_X1 U2399 ( .B1(n2695), .B2(n2097), .A(n3819), .ZN(n2096) );
  NOR2_X1 U2400 ( .A1(n2142), .A2(n2141), .ZN(n2140) );
  INV_X1 U2401 ( .A(n3015), .ZN(n2141) );
  INV_X1 U2402 ( .A(n3016), .ZN(n2142) );
  NAND2_X1 U2403 ( .A1(n2480), .A2(n3893), .ZN(n2479) );
  NAND2_X1 U2404 ( .A1(n2320), .A2(n2316), .ZN(n2335) );
  INV_X1 U2405 ( .A(IR_REG_19__SCAN_IN), .ZN(n2606) );
  NOR2_X1 U2406 ( .A1(n3501), .A2(n2202), .ZN(n2201) );
  INV_X1 U2407 ( .A(n2200), .ZN(n2199) );
  INV_X1 U2408 ( .A(n2193), .ZN(n2192) );
  OAI22_X1 U2409 ( .A1(n3300), .A2(n2194), .B1(n3298), .B2(n3299), .ZN(n2193)
         );
  NAND2_X1 U2410 ( .A1(n3262), .A2(n2049), .ZN(n2191) );
  NOR2_X1 U2411 ( .A1(n2163), .A2(n2159), .ZN(n2158) );
  INV_X1 U2412 ( .A(n2165), .ZN(n2163) );
  INV_X1 U2413 ( .A(n3688), .ZN(n2159) );
  INV_X1 U2414 ( .A(n2168), .ZN(n2162) );
  NOR2_X1 U2415 ( .A1(n3737), .A2(n2166), .ZN(n2165) );
  INV_X1 U2416 ( .A(n3606), .ZN(n2176) );
  AOI21_X1 U2417 ( .B1(n2181), .B2(n2179), .A(n2071), .ZN(n2178) );
  INV_X1 U2418 ( .A(n2184), .ZN(n2179) );
  NAND2_X1 U2419 ( .A1(n2204), .A2(n2203), .ZN(n2206) );
  AOI21_X1 U2420 ( .B1(n2205), .B2(n3058), .A(n3087), .ZN(n2203) );
  NOR2_X1 U2421 ( .A1(n3057), .A2(n3058), .ZN(n3080) );
  NAND2_X1 U2422 ( .A1(n3546), .A2(n3545), .ZN(n3547) );
  NAND2_X1 U2423 ( .A1(n4011), .A2(n4409), .ZN(n2870) );
  AND3_X1 U2424 ( .A1(n2257), .A2(n2256), .A3(n2255), .ZN(n3972) );
  OR2_X1 U2425 ( .A1(n3971), .A2(n2254), .ZN(n2257) );
  XNOR2_X1 U2426 ( .A(n2109), .B(n4414), .ZN(n3982) );
  OAI22_X1 U2427 ( .A1(n3982), .A2(n3238), .B1(n2355), .B2(n2108), .ZN(n2263)
         );
  INV_X1 U2428 ( .A(n2109), .ZN(n2108) );
  NOR2_X1 U2429 ( .A1(n2802), .A2(n2268), .ZN(n2271) );
  NOR2_X1 U2430 ( .A1(n2806), .A2(n2267), .ZN(n2268) );
  AOI21_X1 U2431 ( .B1(n2116), .B2(n2113), .A(n2065), .ZN(n2112) );
  INV_X1 U2432 ( .A(n2116), .ZN(n2114) );
  INV_X1 U2433 ( .A(n2120), .ZN(n2113) );
  NAND2_X1 U2434 ( .A1(n4445), .A2(REG2_REG_10__SCAN_IN), .ZN(n4444) );
  NAND2_X1 U2435 ( .A1(n4449), .A2(n2365), .ZN(n4454) );
  NAND2_X1 U2436 ( .A1(n4471), .A2(n2368), .ZN(n3255) );
  NAND2_X1 U2437 ( .A1(n3255), .A2(n3254), .ZN(n3253) );
  NAND2_X1 U2438 ( .A1(n4456), .A2(n2287), .ZN(n2289) );
  NAND2_X1 U2439 ( .A1(n4467), .A2(REG2_REG_12__SCAN_IN), .ZN(n4465) );
  NAND2_X1 U2440 ( .A1(n2153), .A2(n2154), .ZN(n2155) );
  NOR2_X1 U2441 ( .A1(n2670), .A2(n2669), .ZN(n4052) );
  AND2_X1 U2442 ( .A1(n4286), .A2(n4076), .ZN(n2669) );
  NOR2_X1 U2443 ( .A1(n3866), .A2(n4103), .ZN(n4067) );
  OR2_X1 U2444 ( .A1(n2629), .A2(n2391), .ZN(n2639) );
  OAI22_X1 U2445 ( .A1(n4172), .A2(n2621), .B1(n3668), .B2(n4188), .ZN(n4158)
         );
  AND2_X1 U2446 ( .A1(n3913), .A2(n3788), .ZN(n3881) );
  NAND2_X1 U2447 ( .A1(n2135), .A2(n2134), .ZN(n3332) );
  INV_X1 U2448 ( .A(n3889), .ZN(n2134) );
  INV_X1 U2449 ( .A(n3334), .ZN(n2135) );
  OR2_X1 U2450 ( .A1(n3286), .A2(n3894), .ZN(n3284) );
  AND2_X1 U2451 ( .A1(n3796), .A2(n3834), .ZN(n3894) );
  NAND2_X1 U2452 ( .A1(n2144), .A2(n2500), .ZN(n3185) );
  NAND2_X1 U2453 ( .A1(n3128), .A2(n2499), .ZN(n2144) );
  NAND2_X1 U2454 ( .A1(n2957), .A2(n3804), .ZN(n2991) );
  NAND2_X1 U2455 ( .A1(n2991), .A2(n3877), .ZN(n2990) );
  AND2_X1 U2456 ( .A1(n2725), .A2(n2771), .ZN(n3006) );
  NOR2_X1 U2457 ( .A1(n4264), .A2(n4267), .ZN(n4263) );
  NAND2_X1 U2458 ( .A1(n3612), .A2(n4024), .ZN(n4264) );
  INV_X1 U2459 ( .A(n3503), .ZN(n3639) );
  AND4_X1 U2460 ( .A1(n2528), .A2(n2527), .A3(n2526), .A4(n2525), .ZN(n3439)
         );
  NAND2_X1 U2461 ( .A1(n3047), .A2(n3026), .ZN(n3038) );
  NAND2_X1 U2462 ( .A1(n4185), .A2(n4530), .ZN(n4340) );
  AND2_X1 U2463 ( .A1(n2858), .A2(n4522), .ZN(n2864) );
  NOR2_X1 U2464 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2318)
         );
  NOR2_X1 U2465 ( .A1(n2283), .A2(n2282), .ZN(n2791) );
  AND2_X1 U2466 ( .A1(n2613), .A2(n2598), .ZN(n4211) );
  NAND2_X1 U2467 ( .A1(n2057), .A2(n3591), .ZN(n2873) );
  OR2_X1 U2468 ( .A1(n2433), .A2(n2416), .ZN(n2423) );
  INV_X1 U2469 ( .A(n3287), .ZN(n3387) );
  INV_X1 U2470 ( .A(n3958), .ZN(n3388) );
  INV_X1 U2471 ( .A(n3776), .ZN(n3757) );
  AND2_X1 U2472 ( .A1(n2663), .A2(n2662), .ZN(n4077) );
  NAND2_X1 U2473 ( .A1(n2656), .A2(n2655), .ZN(n4283) );
  INV_X1 U2474 ( .A(n3700), .ZN(n4334) );
  NAND4_X1 U2475 ( .A1(n2429), .A2(n2428), .A3(n2427), .A4(n2426), .ZN(n3966)
         );
  NAND2_X1 U2476 ( .A1(n2579), .A2(REG1_REG_0__SCAN_IN), .ZN(n2429) );
  NOR2_X1 U2477 ( .A1(n2804), .A2(n2803), .ZN(n2802) );
  NAND2_X1 U2478 ( .A1(n4457), .A2(n4458), .ZN(n4456) );
  INV_X1 U2479 ( .A(n2155), .ZN(n3990) );
  NOR2_X1 U2480 ( .A1(n2346), .A2(n2347), .ZN(n4002) );
  INV_X1 U2481 ( .A(n4466), .ZN(n4495) );
  AND2_X1 U2482 ( .A1(n4426), .A2(n2378), .ZN(n4502) );
  OR2_X1 U2483 ( .A1(n4002), .A2(n2102), .ZN(n2101) );
  AND2_X1 U2484 ( .A1(n4003), .A2(REG2_REG_18__SCAN_IN), .ZN(n2102) );
  OAI21_X1 U2485 ( .B1(n2153), .B2(n2152), .A(n2151), .ZN(n4008) );
  AOI21_X1 U2486 ( .B1(n2156), .B2(n3988), .A(n2073), .ZN(n2151) );
  XNOR2_X1 U2487 ( .A(n2686), .B(n3862), .ZN(n4022) );
  NAND2_X1 U2488 ( .A1(n2724), .A2(n2723), .ZN(n4029) );
  NAND2_X1 U2489 ( .A1(n2722), .A2(n2212), .ZN(n2723) );
  NAND2_X1 U2490 ( .A1(n4215), .A2(n2775), .ZN(n4213) );
  INV_X1 U2491 ( .A(n4213), .ZN(n4514) );
  INV_X1 U2492 ( .A(IR_REG_29__SCAN_IN), .ZN(n2396) );
  INV_X1 U2493 ( .A(n3543), .ZN(n3546) );
  AND2_X1 U2494 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2443) );
  NOR2_X1 U2495 ( .A1(n2557), .A2(n3766), .ZN(n2556) );
  INV_X1 U2496 ( .A(IR_REG_6__SCAN_IN), .ZN(n2240) );
  NAND2_X1 U2497 ( .A1(n2128), .A2(n2127), .ZN(n2126) );
  INV_X1 U2498 ( .A(n2647), .ZN(n2127) );
  AND2_X1 U2499 ( .A1(n2576), .A2(REG3_REG_19__SCAN_IN), .ZN(n2595) );
  NOR2_X1 U2500 ( .A1(n2585), .A2(n2577), .ZN(n2576) );
  INV_X1 U2501 ( .A(n2133), .ZN(n2132) );
  AOI21_X1 U2502 ( .B1(n2133), .B2(n2131), .A(n2058), .ZN(n2130) );
  AOI21_X1 U2503 ( .B1(n3889), .B2(n2555), .A(n2053), .ZN(n2133) );
  NAND2_X1 U2504 ( .A1(n2083), .A2(n2086), .ZN(n2082) );
  AND2_X1 U2505 ( .A1(n3343), .A2(n3318), .ZN(n3835) );
  INV_X1 U2506 ( .A(n2530), .ZN(n2137) );
  INV_X1 U2507 ( .A(n3834), .ZN(n2086) );
  AOI21_X1 U2508 ( .B1(n2085), .B2(n3834), .A(n2084), .ZN(n2083) );
  INV_X1 U2509 ( .A(n3796), .ZN(n2084) );
  INV_X1 U2510 ( .A(n3828), .ZN(n2085) );
  AND2_X1 U2511 ( .A1(n2512), .A2(REG3_REG_11__SCAN_IN), .ZN(n2521) );
  NOR2_X1 U2512 ( .A1(n3780), .A2(n2620), .ZN(n4178) );
  NOR2_X1 U2513 ( .A1(n3229), .A2(n3287), .ZN(n2076) );
  INV_X1 U2514 ( .A(n3050), .ZN(n3047) );
  AND2_X1 U2515 ( .A1(n3937), .A2(n4409), .ZN(n2841) );
  INV_X1 U2516 ( .A(IR_REG_26__SCAN_IN), .ZN(n2211) );
  NAND2_X1 U2517 ( .A1(n2314), .A2(IR_REG_31__SCAN_IN), .ZN(n2327) );
  INV_X1 U2518 ( .A(IR_REG_23__SCAN_IN), .ZN(n2326) );
  INV_X1 U2519 ( .A(IR_REG_17__SCAN_IN), .ZN(n2229) );
  OR3_X1 U2520 ( .A1(n2248), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2279) );
  INV_X1 U2521 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4639) );
  OR2_X1 U2522 ( .A1(n3649), .A2(n3650), .ZN(n3570) );
  INV_X1 U2523 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4658) );
  OAI22_X1 U2524 ( .A1(n3640), .A2(n3601), .B1(n3600), .B2(n3486), .ZN(n3499)
         );
  AOI21_X1 U2525 ( .B1(n2188), .B2(n2187), .A(n2068), .ZN(n2186) );
  INV_X1 U2526 ( .A(n2049), .ZN(n2187) );
  NAND2_X1 U2527 ( .A1(n2170), .A2(n2168), .ZN(n2167) );
  INV_X1 U2528 ( .A(n2166), .ZN(n2164) );
  AND2_X1 U2529 ( .A1(n2443), .A2(REG3_REG_5__SCAN_IN), .ZN(n2458) );
  OR2_X1 U2530 ( .A1(n2548), .A2(n4639), .ZN(n2557) );
  INV_X1 U2531 ( .A(n2888), .ZN(n2867) );
  AND3_X1 U2532 ( .A1(n2574), .A2(n2573), .A3(n2572), .ZN(n3700) );
  OR2_X1 U2533 ( .A1(n2912), .A2(n2911), .ZN(n2111) );
  NAND2_X1 U2534 ( .A1(n2809), .A2(n2145), .ZN(n2360) );
  NAND2_X1 U2535 ( .A1(n2143), .A2(REG1_REG_5__SCAN_IN), .ZN(n2145) );
  INV_X1 U2536 ( .A(IR_REG_7__SCAN_IN), .ZN(n2273) );
  INV_X1 U2537 ( .A(n2119), .ZN(n2115) );
  NAND2_X1 U2538 ( .A1(n4453), .A2(n2366), .ZN(n2367) );
  AND2_X1 U2539 ( .A1(n2309), .A2(n2227), .ZN(n2292) );
  INV_X1 U2540 ( .A(IR_REG_13__SCAN_IN), .ZN(n2227) );
  NAND2_X1 U2541 ( .A1(n3253), .A2(n2369), .ZN(n2370) );
  XNOR2_X1 U2542 ( .A(n2104), .B(n2554), .ZN(n4477) );
  NOR2_X1 U2543 ( .A1(n4477), .A2(n4478), .ZN(n4476) );
  INV_X1 U2544 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3766) );
  NAND2_X1 U2545 ( .A1(n4498), .A2(n4496), .ZN(n4497) );
  INV_X1 U2546 ( .A(n2156), .ZN(n2152) );
  AOI21_X1 U2547 ( .B1(n3616), .B2(n3783), .A(n2711), .ZN(n2712) );
  NAND2_X1 U2548 ( .A1(n4052), .A2(n2122), .ZN(n2121) );
  NAND2_X1 U2549 ( .A1(n3849), .A2(n4057), .ZN(n2122) );
  AOI21_X1 U2550 ( .B1(n4067), .B2(n2710), .A(n2709), .ZN(n4049) );
  INV_X1 U2551 ( .A(n3848), .ZN(n2709) );
  NAND2_X1 U2552 ( .A1(n4283), .A2(n4291), .ZN(n2657) );
  NAND2_X1 U2553 ( .A1(n2090), .A2(n3915), .ZN(n4121) );
  NAND2_X1 U2554 ( .A1(n3474), .A2(n2087), .ZN(n2090) );
  AND2_X1 U2555 ( .A1(n2088), .A2(n3787), .ZN(n2087) );
  NAND2_X1 U2556 ( .A1(n3474), .A2(n2088), .ZN(n4175) );
  AND2_X1 U2557 ( .A1(n4198), .A2(n4199), .ZN(n4238) );
  OR2_X1 U2558 ( .A1(n2583), .A2(n4646), .ZN(n2585) );
  INV_X1 U2559 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2577) );
  NAND2_X1 U2560 ( .A1(n2080), .A2(n3791), .ZN(n3367) );
  NAND2_X1 U2561 ( .A1(n3335), .A2(n3889), .ZN(n2080) );
  OR2_X1 U2562 ( .A1(n3367), .A2(n3875), .ZN(n3368) );
  AND2_X1 U2563 ( .A1(n3791), .A2(n3789), .ZN(n3889) );
  NAND2_X1 U2564 ( .A1(n2521), .A2(REG3_REG_12__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U2565 ( .A1(n2696), .A2(n3828), .ZN(n3288) );
  AOI21_X1 U2566 ( .B1(n2095), .B2(n2097), .A(n2093), .ZN(n2092) );
  INV_X1 U2567 ( .A(n2096), .ZN(n2095) );
  NAND2_X1 U2568 ( .A1(n2493), .A2(REG3_REG_8__SCAN_IN), .ZN(n2502) );
  NAND2_X1 U2569 ( .A1(n2094), .A2(n3821), .ZN(n3129) );
  NAND2_X1 U2570 ( .A1(n3109), .A2(n2695), .ZN(n2094) );
  NOR2_X1 U2571 ( .A1(n2051), .A2(n3121), .ZN(n2489) );
  NAND2_X1 U2572 ( .A1(n2479), .A2(n2140), .ZN(n2491) );
  AOI21_X1 U2573 ( .B1(n3068), .B2(n3812), .A(n3798), .ZN(n3109) );
  OAI21_X1 U2574 ( .B1(n3034), .B2(n3032), .A(n3823), .ZN(n3068) );
  NAND2_X1 U2575 ( .A1(n2694), .A2(n3204), .ZN(n2457) );
  NAND2_X1 U2576 ( .A1(n2693), .A2(n3814), .ZN(n3034) );
  NAND2_X1 U2577 ( .A1(n2990), .A2(n2098), .ZN(n2693) );
  AND2_X1 U2578 ( .A1(n3810), .A2(n3809), .ZN(n2098) );
  NAND2_X1 U2579 ( .A1(n2759), .A2(n3803), .ZN(n2958) );
  NAND2_X1 U2580 ( .A1(n3895), .A2(n2692), .ZN(n2759) );
  NAND2_X1 U2581 ( .A1(n4088), .A2(n4076), .ZN(n4075) );
  INV_X1 U2582 ( .A(n3864), .ZN(n4076) );
  NOR2_X1 U2583 ( .A1(n4106), .A2(n4282), .ZN(n4088) );
  INV_X1 U2584 ( .A(n4291), .ZN(n4107) );
  OR2_X1 U2585 ( .A1(n4131), .A2(n4291), .ZN(n4106) );
  OR2_X1 U2586 ( .A1(n4148), .A2(n3558), .ZN(n4131) );
  NAND2_X1 U2587 ( .A1(n4161), .A2(n4149), .ZN(n4148) );
  INV_X1 U2588 ( .A(n2638), .ZN(n4149) );
  AND2_X1 U2589 ( .A1(n4186), .A2(n4167), .ZN(n4161) );
  NOR2_X2 U2590 ( .A1(n4208), .A2(n4178), .ZN(n4186) );
  NAND2_X1 U2591 ( .A1(n3469), .A2(n2066), .ZN(n4218) );
  AND2_X1 U2592 ( .A1(n3469), .A2(n3699), .ZN(n4220) );
  INV_X1 U2593 ( .A(n3953), .ZN(n4350) );
  OR2_X1 U2594 ( .A1(n3371), .A2(n3512), .ZN(n3470) );
  NAND2_X1 U2595 ( .A1(n3336), .A2(n3639), .ZN(n3371) );
  INV_X1 U2596 ( .A(n3955), .ZN(n3640) );
  NOR2_X1 U2597 ( .A1(n3349), .A2(n3326), .ZN(n3336) );
  NAND2_X1 U2598 ( .A1(n2076), .A2(n3438), .ZN(n3349) );
  INV_X1 U2599 ( .A(n2076), .ZN(n3347) );
  INV_X1 U2600 ( .A(n3302), .ZN(n3309) );
  AND2_X1 U2601 ( .A1(n3190), .A2(n3268), .ZN(n3228) );
  NAND2_X1 U2602 ( .A1(n3072), .A2(n2054), .ZN(n3136) );
  INV_X1 U2603 ( .A(n3168), .ZN(n3159) );
  NOR2_X2 U2604 ( .A1(n3136), .A2(n3159), .ZN(n3190) );
  NAND2_X1 U2605 ( .A1(n3072), .A2(n3101), .ZN(n3108) );
  INV_X1 U2606 ( .A(n4349), .ZN(n4333) );
  NOR2_X1 U2607 ( .A1(n2995), .A2(n4251), .ZN(n2074) );
  INV_X1 U2608 ( .A(n2996), .ZN(n2075) );
  INV_X1 U2609 ( .A(n2995), .ZN(n3239) );
  INV_X1 U2610 ( .A(n4346), .ZN(n4337) );
  INV_X1 U2611 ( .A(n3107), .ZN(n4352) );
  INV_X1 U2612 ( .A(n4203), .ZN(n4345) );
  AND2_X1 U2613 ( .A1(n4418), .A2(n2841), .ZN(n4346) );
  INV_X1 U2614 ( .A(n2838), .ZN(n2770) );
  AND3_X1 U2615 ( .A1(n2745), .A2(n2744), .A3(n2765), .ZN(n2754) );
  AND2_X1 U2616 ( .A1(n2731), .A2(n4408), .ZN(n2766) );
  NAND2_X1 U2617 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2213) );
  NAND2_X1 U2618 ( .A1(n2327), .A2(n2326), .ZN(n2329) );
  XNOR2_X1 U2619 ( .A(n2336), .B(n2310), .ZN(n2725) );
  INV_X1 U2620 ( .A(IR_REG_20__SCAN_IN), .ZN(n2688) );
  XNOR2_X1 U2621 ( .A(n2246), .B(IR_REG_11__SCAN_IN), .ZN(n2529) );
  NOR2_X1 U2622 ( .A1(n2239), .A2(IR_REG_5__SCAN_IN), .ZN(n2269) );
  INV_X1 U2623 ( .A(IR_REG_5__SCAN_IN), .ZN(n2265) );
  NAND2_X1 U2624 ( .A1(n2253), .A2(n2252), .ZN(n3971) );
  MUX2_X1 U2625 ( .A(IR_REG_31__SCAN_IN), .B(n2251), .S(IR_REG_1__SCAN_IN), 
        .Z(n2253) );
  INV_X1 U2626 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4646) );
  INV_X1 U2627 ( .A(n2201), .ZN(n2197) );
  NAND2_X1 U2628 ( .A1(n2191), .A2(n2192), .ZN(n3307) );
  AOI21_X1 U2629 ( .B1(n2165), .B2(n2162), .A(n2161), .ZN(n2160) );
  INV_X1 U2630 ( .A(n3738), .ZN(n2161) );
  AND2_X1 U2631 ( .A1(n2178), .A2(n2176), .ZN(n2172) );
  OAI21_X1 U2632 ( .B1(n2178), .B2(n3606), .A(n2174), .ZN(n2173) );
  NAND2_X1 U2633 ( .A1(n2178), .A2(n2175), .ZN(n2174) );
  NAND2_X1 U2634 ( .A1(n2180), .A2(n2176), .ZN(n2175) );
  NAND2_X1 U2635 ( .A1(n2181), .A2(n3606), .ZN(n2177) );
  AND2_X1 U2636 ( .A1(n2636), .A2(n2635), .ZN(n4315) );
  INV_X1 U2637 ( .A(n3204), .ZN(n3090) );
  NOR2_X1 U2638 ( .A1(n3080), .A2(n2207), .ZN(n3088) );
  AND4_X1 U2639 ( .A1(n2498), .A2(n2497), .A3(n2496), .A4(n2495), .ZN(n3269)
         );
  INV_X1 U2640 ( .A(n3263), .ZN(n3268) );
  AOI21_X1 U2641 ( .B1(n3262), .B2(n3261), .A(n2045), .ZN(n3301) );
  NAND2_X1 U2642 ( .A1(n2882), .A2(n2881), .ZN(n2884) );
  INV_X1 U2643 ( .A(n4222), .ZN(n4219) );
  AND2_X1 U2644 ( .A1(n2983), .A2(n2982), .ZN(n3776) );
  INV_X1 U2645 ( .A(n3512), .ZN(n3767) );
  INV_X1 U2646 ( .A(n3753), .ZN(n3770) );
  INV_X1 U2647 ( .A(n3755), .ZN(n3772) );
  INV_X1 U2648 ( .A(n3759), .ZN(n3764) );
  NAND2_X1 U2649 ( .A1(n2668), .A2(n2667), .ZN(n4270) );
  NAND2_X1 U2650 ( .A1(n2645), .A2(n2644), .ZN(n4292) );
  INV_X1 U2651 ( .A(n4315), .ZN(n4162) );
  NAND2_X1 U2652 ( .A1(n2626), .A2(n2625), .ZN(n4141) );
  NAND2_X1 U2653 ( .A1(n2619), .A2(n2618), .ZN(n4312) );
  NAND2_X1 U2654 ( .A1(n2604), .A2(n2603), .ZN(n4179) );
  INV_X1 U2655 ( .A(n2111), .ZN(n2910) );
  NAND2_X1 U2656 ( .A1(n2935), .A2(n2055), .ZN(n2810) );
  NAND2_X1 U2657 ( .A1(n2810), .A2(n2811), .ZN(n2809) );
  AOI21_X1 U2658 ( .B1(n2934), .B2(REG2_REG_4__SCAN_IN), .A(n2264), .ZN(n2804)
         );
  XNOR2_X1 U2659 ( .A(n2360), .B(n4412), .ZN(n2818) );
  AOI22_X1 U2660 ( .A1(n2814), .A2(REG2_REG_6__SCAN_IN), .B1(n4412), .B2(n2272), .ZN(n2832) );
  AOI21_X1 U2661 ( .B1(n4412), .B2(n2360), .A(n2815), .ZN(n2827) );
  XNOR2_X1 U2662 ( .A(n2362), .B(n2148), .ZN(n2945) );
  XNOR2_X1 U2663 ( .A(n2278), .B(n4411), .ZN(n2947) );
  OAI21_X1 U2664 ( .B1(n2945), .B2(n2492), .A(n2147), .ZN(n4436) );
  NAND2_X1 U2665 ( .A1(n2362), .A2(n2148), .ZN(n2147) );
  NAND2_X1 U2666 ( .A1(n2118), .A2(n2116), .ZN(n4431) );
  AND2_X1 U2667 ( .A1(n2118), .A2(n2115), .ZN(n4433) );
  NAND2_X1 U2668 ( .A1(n2278), .A2(n2120), .ZN(n2118) );
  NAND2_X1 U2669 ( .A1(n4444), .A2(n2286), .ZN(n4457) );
  XNOR2_X1 U2670 ( .A(n2367), .B(n2288), .ZN(n4472) );
  AND2_X1 U2671 ( .A1(n4426), .A2(n3943), .ZN(n4466) );
  NAND2_X1 U2672 ( .A1(n2290), .A2(n4465), .ZN(n3251) );
  XNOR2_X1 U2673 ( .A(n2370), .B(n2146), .ZN(n4482) );
  OAI21_X1 U2674 ( .B1(n4477), .B2(n2106), .A(n2105), .ZN(n4485) );
  NAND2_X1 U2675 ( .A1(n2107), .A2(REG2_REG_14__SCAN_IN), .ZN(n2106) );
  NAND2_X1 U2676 ( .A1(n2295), .A2(n2107), .ZN(n2105) );
  INV_X1 U2677 ( .A(n4486), .ZN(n2107) );
  AND2_X1 U2678 ( .A1(n2383), .A2(n2382), .ZN(n4501) );
  NAND2_X1 U2679 ( .A1(n3993), .A2(n2103), .ZN(n2346) );
  NAND2_X1 U2680 ( .A1(n4001), .A2(n2586), .ZN(n2103) );
  NAND2_X1 U2681 ( .A1(n2155), .A2(n2156), .ZN(n4005) );
  NOR2_X1 U2682 ( .A1(n3990), .A2(n2377), .ZN(n2379) );
  INV_X1 U2683 ( .A(n4067), .ZN(n4083) );
  NAND2_X1 U2684 ( .A1(n3474), .A2(n3788), .ZN(n3455) );
  NAND2_X1 U2685 ( .A1(n3332), .A2(n2555), .ZN(n3370) );
  NAND2_X1 U2686 ( .A1(n3284), .A2(n2530), .ZN(n3346) );
  NAND4_X1 U2687 ( .A1(n2519), .A2(n2518), .A3(n2517), .A4(n2516), .ZN(n3958)
         );
  INV_X1 U2688 ( .A(n3959), .ZN(n3310) );
  INV_X1 U2689 ( .A(n4113), .ZN(n4254) );
  NAND2_X1 U2690 ( .A1(n2990), .A2(n3809), .ZN(n3021) );
  AND2_X1 U2691 ( .A1(n4511), .A2(n4333), .ZN(n4248) );
  NAND2_X1 U2692 ( .A1(n4536), .A2(n2772), .ZN(n4508) );
  INV_X1 U2693 ( .A(n4419), .ZN(n4215) );
  AND2_X2 U2694 ( .A1(n2754), .A2(n2838), .ZN(n4552) );
  NOR2_X1 U2695 ( .A1(n4029), .A2(n2099), .ZN(n2755) );
  NAND2_X1 U2696 ( .A1(n2100), .A2(n2727), .ZN(n2099) );
  NAND2_X1 U2697 ( .A1(n4022), .A2(n4340), .ZN(n2100) );
  NAND2_X1 U2698 ( .A1(n4264), .A2(n2751), .ZN(n4027) );
  OR2_X1 U2699 ( .A1(n3612), .A2(n4024), .ZN(n2751) );
  AND2_X2 U2700 ( .A1(n2754), .A2(n2770), .ZN(n4546) );
  NAND2_X1 U2701 ( .A1(n3494), .A2(IR_REG_31__SCAN_IN), .ZN(n2397) );
  AND2_X1 U2702 ( .A1(n2320), .A2(n2046), .ZN(n2398) );
  MUX2_X1 U2703 ( .A(IR_REG_31__SCAN_IN), .B(n2315), .S(IR_REG_25__SCAN_IN), 
        .Z(n2321) );
  AND2_X1 U2704 ( .A1(n2337), .A2(STATE_REG_SCAN_IN), .ZN(n4522) );
  INV_X1 U2705 ( .A(n2771), .ZN(n3937) );
  XNOR2_X1 U2706 ( .A(n2101), .B(n4004), .ZN(n4015) );
  AOI22_X1 U2707 ( .A1(n4420), .A2(n4514), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4419), .ZN(n4421) );
  NAND2_X1 U2708 ( .A1(n2056), .A2(n3520), .ZN(n2170) );
  AND2_X1 U2709 ( .A1(n3162), .A2(n3163), .ZN(n2045) );
  AND2_X1 U2710 ( .A1(n2061), .A2(n2319), .ZN(n2046) );
  OAI21_X1 U2711 ( .B1(n2827), .B2(n2361), .A(n2069), .ZN(n2362) );
  NOR2_X1 U2712 ( .A1(n4233), .A2(n2593), .ZN(n2047) );
  INV_X1 U2713 ( .A(n2189), .ZN(n2188) );
  NAND2_X1 U2714 ( .A1(n2192), .A2(n2190), .ZN(n2189) );
  INV_X1 U2715 ( .A(n3822), .ZN(n2093) );
  NOR2_X1 U2716 ( .A1(n3454), .A2(n2089), .ZN(n2048) );
  INV_X1 U2717 ( .A(n2554), .ZN(n2146) );
  INV_X1 U2718 ( .A(n3988), .ZN(n2154) );
  NOR2_X1 U2719 ( .A1(n3300), .A2(n2195), .ZN(n2049) );
  AND3_X1 U2720 ( .A1(n2468), .A2(n2467), .A3(n2466), .ZN(n2050) );
  AND2_X1 U2721 ( .A1(n3961), .A2(n3152), .ZN(n2051) );
  XNOR2_X1 U2722 ( .A(n2877), .B(n3602), .ZN(n2882) );
  INV_X1 U2723 ( .A(n4414), .ZN(n2355) );
  AND2_X1 U2724 ( .A1(n2308), .A2(n2309), .ZN(n2320) );
  NAND2_X1 U2725 ( .A1(n2707), .A2(n3869), .ZN(n4103) );
  NAND2_X1 U2726 ( .A1(n2183), .A2(n3748), .ZN(n3627) );
  NAND2_X1 U2727 ( .A1(n2170), .A2(n3525), .ZN(n3695) );
  NAND2_X1 U2728 ( .A1(n2167), .A2(n2164), .ZN(n3736) );
  AND4_X1 U2729 ( .A1(n2423), .A2(n2422), .A3(n2421), .A4(n2420), .ZN(n2880)
         );
  XNOR2_X1 U2730 ( .A(n2397), .B(IR_REG_30__SCAN_IN), .ZN(n4407) );
  AND2_X1 U2731 ( .A1(n3956), .A2(n3433), .ZN(n2052) );
  NOR2_X1 U2732 ( .A1(n2323), .A2(IR_REG_26__SCAN_IN), .ZN(n2339) );
  AND2_X1 U2733 ( .A1(n3953), .A2(n3512), .ZN(n2053) );
  AND2_X1 U2734 ( .A1(n3101), .A2(n3177), .ZN(n2054) );
  INV_X1 U2735 ( .A(n4251), .ZN(n2962) );
  INV_X1 U2736 ( .A(n2077), .ZN(n4056) );
  OR2_X1 U2737 ( .A1(n2359), .A2(n2940), .ZN(n2055) );
  AND2_X1 U2738 ( .A1(n3683), .A2(n3688), .ZN(n2056) );
  AND2_X1 U2739 ( .A1(n2854), .A2(n2853), .ZN(n2057) );
  AND2_X1 U2740 ( .A1(n4350), .A2(n3767), .ZN(n2058) );
  AND2_X1 U2741 ( .A1(n3487), .A2(n3438), .ZN(n2059) );
  INV_X1 U2742 ( .A(IR_REG_2__SCAN_IN), .ZN(n4585) );
  NAND2_X1 U2743 ( .A1(n3474), .A2(n2048), .ZN(n2060) );
  AND2_X1 U2744 ( .A1(n2209), .A2(n2208), .ZN(n2061) );
  NAND2_X1 U2745 ( .A1(n3096), .A2(n3095), .ZN(n2062) );
  INV_X1 U2746 ( .A(IR_REG_31__SCAN_IN), .ZN(n3493) );
  NAND2_X1 U2747 ( .A1(n4162), .A2(n2638), .ZN(n2063) );
  OAI21_X1 U2748 ( .B1(n2696), .B2(n2086), .A(n2083), .ZN(n3316) );
  AND2_X1 U2749 ( .A1(n4125), .A2(n2704), .ZN(n4146) );
  INV_X1 U2750 ( .A(n4146), .ZN(n2128) );
  AND2_X1 U2751 ( .A1(n3157), .A2(n3156), .ZN(n2064) );
  AND2_X1 U2752 ( .A1(n3429), .A2(n3428), .ZN(n3480) );
  INV_X1 U2753 ( .A(n2196), .ZN(n3634) );
  AND2_X1 U2754 ( .A1(n2129), .A2(n2063), .ZN(n4120) );
  INV_X1 U2755 ( .A(n3748), .ZN(n2182) );
  NAND2_X1 U2756 ( .A1(n3961), .A2(n3177), .ZN(n3821) );
  INV_X1 U2757 ( .A(n3821), .ZN(n2097) );
  NAND2_X1 U2758 ( .A1(n2407), .A2(n2406), .ZN(n4072) );
  AND2_X1 U2759 ( .A1(n2791), .A2(REG2_REG_9__SCAN_IN), .ZN(n2065) );
  AND2_X1 U2760 ( .A1(n3699), .A2(n4219), .ZN(n2066) );
  NOR2_X1 U2761 ( .A1(n4476), .A2(n2295), .ZN(n2067) );
  AND2_X1 U2762 ( .A1(n3380), .A2(n3382), .ZN(n2068) );
  XOR2_X1 U2763 ( .A(n3602), .B(n3483), .Z(n3501) );
  OR2_X1 U2764 ( .A1(n2829), .A2(n4550), .ZN(n2069) );
  INV_X1 U2765 ( .A(n2181), .ZN(n2180) );
  NOR2_X1 U2766 ( .A1(n3628), .A2(n2182), .ZN(n2181) );
  NAND2_X1 U2767 ( .A1(n3636), .A2(n3507), .ZN(n2070) );
  OR2_X1 U2768 ( .A1(n4147), .A2(n4146), .ZN(n2129) );
  AND2_X1 U2769 ( .A1(n3598), .A2(n3597), .ZN(n2071) );
  AND2_X1 U2770 ( .A1(n3835), .A2(n2082), .ZN(n2072) );
  BUF_X1 U2771 ( .A(n2432), .Z(n2680) );
  INV_X1 U2772 ( .A(n3788), .ZN(n2089) );
  NAND2_X1 U2773 ( .A1(n2191), .A2(n2188), .ZN(n3383) );
  AND4_X1 U2774 ( .A1(n2484), .A2(n2483), .A3(n2482), .A4(n2481), .ZN(n3084)
         );
  NAND2_X1 U2775 ( .A1(n2691), .A2(n3937), .ZN(n2871) );
  INV_X1 U2776 ( .A(IR_REG_28__SCAN_IN), .ZN(n2208) );
  INV_X1 U2777 ( .A(n2045), .ZN(n2194) );
  NOR2_X1 U2778 ( .A1(n4523), .A2(n4006), .ZN(n2073) );
  INV_X1 U2779 ( .A(n2806), .ZN(n2143) );
  INV_X1 U2780 ( .A(n4411), .ZN(n2148) );
  NOR2_X1 U2781 ( .A1(n4075), .A2(n4269), .ZN(n2077) );
  NOR3_X1 U2782 ( .A1(n4075), .A2(n4269), .A3(n3618), .ZN(n3612) );
  AND2_X2 U2783 ( .A1(n2075), .A2(n2074), .ZN(n3026) );
  OR2_X2 U2784 ( .A1(n4218), .A2(n3539), .ZN(n4208) );
  NAND4_X1 U2785 ( .A1(n2224), .A2(n2225), .A3(n2226), .A4(n2223), .ZN(n2078)
         );
  NAND3_X1 U2786 ( .A1(n2308), .A2(n2309), .A3(n2319), .ZN(n2323) );
  NAND2_X1 U2787 ( .A1(n2079), .A2(n4585), .ZN(n2258) );
  NAND2_X1 U2788 ( .A1(n2696), .A2(n2083), .ZN(n2081) );
  NAND2_X1 U2789 ( .A1(n2081), .A2(n2072), .ZN(n2698) );
  NAND2_X1 U2790 ( .A1(n3109), .A2(n2095), .ZN(n2091) );
  NAND2_X1 U2791 ( .A1(n2091), .A2(n2092), .ZN(n3186) );
  NAND4_X1 U2792 ( .A1(n2046), .A2(n2308), .A3(n2309), .A4(n2396), .ZN(n3494)
         );
  OAI21_X1 U2793 ( .B1(n3186), .B2(n3831), .A(n3820), .ZN(n3226) );
  OAI21_X1 U2794 ( .B1(n4121), .B2(n2706), .A(n3917), .ZN(n2707) );
  INV_X1 U2795 ( .A(n2294), .ZN(n2104) );
  OAI21_X1 U2796 ( .B1(n2278), .B2(n2114), .A(n2112), .ZN(n2285) );
  NAND2_X2 U2797 ( .A1(n2125), .A2(n2123), .ZN(n4101) );
  OR2_X2 U2798 ( .A1(n4147), .A2(n2126), .ZN(n2125) );
  INV_X1 U2799 ( .A(n2129), .ZN(n4306) );
  INV_X1 U2800 ( .A(n4101), .ZN(n2658) );
  OAI21_X1 U2801 ( .B1(n3334), .B2(n2132), .A(n2130), .ZN(n3457) );
  OAI21_X1 U2802 ( .B1(n3286), .B2(n2138), .A(n2136), .ZN(n3325) );
  NOR2_X1 U2803 ( .A1(n3113), .A2(n2051), .ZN(n2480) );
  MUX2_X1 U2804 ( .A(n2143), .B(DATAI_5_), .S(n3779), .Z(n3204) );
  NAND2_X1 U2805 ( .A1(n4436), .A2(n4435), .ZN(n4434) );
  NAND2_X1 U2806 ( .A1(n2150), .A2(n2149), .ZN(n2250) );
  NAND2_X1 U2807 ( .A1(n4585), .A2(n3493), .ZN(n2149) );
  NAND3_X1 U2808 ( .A1(n2252), .A2(IR_REG_2__SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n2150) );
  INV_X1 U2809 ( .A(n3989), .ZN(n2153) );
  NAND3_X1 U2810 ( .A1(n3520), .A2(n2158), .A3(n3683), .ZN(n2157) );
  NAND2_X1 U2811 ( .A1(n2157), .A2(n2160), .ZN(n3658) );
  NAND2_X1 U2812 ( .A1(n3588), .A2(n2172), .ZN(n2171) );
  NAND2_X1 U2813 ( .A1(n3588), .A2(n2184), .ZN(n2183) );
  OAI211_X1 U2814 ( .C1(n3588), .C2(n2177), .A(n2173), .B(n2171), .ZN(n3611)
         );
  NAND2_X1 U2815 ( .A1(n3588), .A2(n3675), .ZN(n3747) );
  NOR2_X1 U2816 ( .A1(n3749), .A2(n2185), .ZN(n2184) );
  INV_X1 U2817 ( .A(n3675), .ZN(n2185) );
  AOI21_X1 U2818 ( .B1(n3500), .B2(n2197), .A(n2199), .ZN(n2196) );
  NAND2_X1 U2819 ( .A1(n3057), .A2(n2205), .ZN(n2204) );
  INV_X1 U2820 ( .A(n2206), .ZN(n3097) );
  AND2_X1 U2821 ( .A1(n3081), .A2(n3082), .ZN(n2207) );
  OR2_X1 U2822 ( .A1(n3019), .A2(n3893), .ZN(n3115) );
  OAI211_X1 U2823 ( .C1(n3461), .C2(n2680), .A(n2588), .B(n2587), .ZN(n4347)
         );
  NAND2_X1 U2824 ( .A1(n2862), .A2(n2861), .ZN(n2874) );
  NAND2_X1 U2825 ( .A1(n3963), .A2(n3050), .ZN(n3031) );
  NAND2_X1 U2826 ( .A1(n2402), .A2(n2400), .ZN(n2425) );
  INV_X1 U2827 ( .A(n2871), .ZN(n2847) );
  OR2_X1 U2828 ( .A1(n2425), .A2(n2431), .ZN(n2438) );
  AOI21_X1 U2829 ( .B1(n2658), .B2(n2657), .A(n2215), .ZN(n4086) );
  OR2_X1 U2830 ( .A1(n2432), .A2(n3010), .ZN(n2427) );
  NAND2_X1 U2831 ( .A1(n4407), .A2(n2400), .ZN(n2434) );
  INV_X1 U2832 ( .A(n2881), .ZN(n2883) );
  NAND2_X1 U2833 ( .A1(n4407), .A2(n3497), .ZN(n2432) );
  AOI21_X2 U2834 ( .B1(n3646), .B2(n3572), .A(n3571), .ZN(n3651) );
  AND2_X1 U2835 ( .A1(n2714), .A2(n2713), .ZN(n4206) );
  INV_X1 U2836 ( .A(n4206), .ZN(n2715) );
  AND2_X1 U2837 ( .A1(n4346), .A2(n2721), .ZN(n2212) );
  INV_X1 U2838 ( .A(n3785), .ZN(n2700) );
  INV_X1 U2839 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2501) );
  INV_X1 U2840 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2254) );
  INV_X1 U2841 ( .A(IR_REG_27__SCAN_IN), .ZN(n2338) );
  AND2_X1 U2842 ( .A1(n4061), .A2(n3618), .ZN(n2214) );
  AND2_X1 U2843 ( .A1(n3653), .A2(n4107), .ZN(n2215) );
  OR2_X1 U2844 ( .A1(n2858), .A2(n2855), .ZN(n2216) );
  INV_X1 U2845 ( .A(U4043), .ZN(n3965) );
  NOR2_X1 U2846 ( .A1(n3780), .A2(n2408), .ZN(n4282) );
  NOR2_X1 U2847 ( .A1(n3780), .A2(n2390), .ZN(n4269) );
  XNOR2_X1 U2848 ( .A(n2882), .B(n2883), .ZN(n2924) );
  INV_X1 U2849 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2539) );
  NAND2_X1 U2850 ( .A1(n2415), .A2(n2414), .ZN(n3950) );
  INV_X1 U2851 ( .A(DATAI_3_), .ZN(n2477) );
  INV_X1 U2852 ( .A(n4404), .ZN(n3362) );
  NAND2_X1 U2853 ( .A1(n3017), .A2(n2480), .ZN(n2217) );
  NAND2_X1 U2854 ( .A1(n4552), .A2(n4352), .ZN(n4343) );
  NOR2_X1 U2855 ( .A1(n2593), .A2(n4234), .ZN(n2218) );
  AND2_X1 U2856 ( .A1(n4270), .A2(n3864), .ZN(n2219) );
  INV_X1 U2857 ( .A(n3923), .ZN(n2710) );
  INV_X1 U2858 ( .A(n3875), .ZN(n2699) );
  XNOR2_X1 U2859 ( .A(n2247), .B(IR_REG_10__SCAN_IN), .ZN(n4443) );
  INV_X1 U2860 ( .A(n4464), .ZN(n2288) );
  AND2_X1 U2861 ( .A1(n3577), .A2(n3578), .ZN(n2220) );
  INV_X1 U2862 ( .A(n3799), .ZN(n2692) );
  OR2_X1 U2863 ( .A1(n3149), .A2(n3148), .ZN(n2221) );
  INV_X1 U2864 ( .A(n3544), .ZN(n3545) );
  INV_X1 U2865 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2267) );
  NAND2_X1 U2866 ( .A1(n3962), .A2(n3218), .ZN(n2486) );
  INV_X1 U2867 ( .A(n2649), .ZN(n2393) );
  INV_X1 U2868 ( .A(n4443), .ZN(n2284) );
  AND2_X1 U2869 ( .A1(n2697), .A2(n3319), .ZN(n3794) );
  NAND2_X1 U2870 ( .A1(n3063), .A2(n2486), .ZN(n3113) );
  INV_X1 U2871 ( .A(IR_REG_21__SCAN_IN), .ZN(n2316) );
  OR2_X1 U2872 ( .A1(n2651), .A2(n2409), .ZN(n2661) );
  NAND2_X1 U2873 ( .A1(n2393), .A2(REG3_REG_24__SCAN_IN), .ZN(n2651) );
  INV_X1 U2874 ( .A(n3497), .ZN(n2400) );
  NAND2_X1 U2875 ( .A1(n4072), .A2(n4269), .ZN(n2671) );
  NAND2_X1 U2876 ( .A1(n3950), .A2(n4282), .ZN(n2659) );
  INV_X1 U2877 ( .A(n3950), .ZN(n4295) );
  INV_X1 U2878 ( .A(n3113), .ZN(n3114) );
  AND2_X1 U2879 ( .A1(n3804), .A2(n3807), .ZN(n3892) );
  NOR2_X1 U2880 ( .A1(n2279), .A2(IR_REG_9__SCAN_IN), .ZN(n2282) );
  INV_X1 U2881 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2463) );
  NOR2_X1 U2882 ( .A1(n2513), .A2(n4658), .ZN(n2512) );
  NAND2_X1 U2883 ( .A1(n2595), .A2(REG3_REG_20__SCAN_IN), .ZN(n2629) );
  NAND2_X1 U2884 ( .A1(n3651), .A2(n2220), .ZN(n3707) );
  INV_X1 U2885 ( .A(n4179), .ZN(n4224) );
  INV_X1 U2886 ( .A(n4072), .ZN(n3849) );
  NOR2_X1 U2887 ( .A1(n3600), .A2(n2849), .ZN(n3944) );
  OAI21_X1 U2888 ( .B1(n4507), .B2(n4523), .A(n2384), .ZN(n2385) );
  INV_X1 U2889 ( .A(n3614), .ZN(n3908) );
  INV_X1 U2890 ( .A(n4270), .ZN(n4286) );
  NOR2_X1 U2891 ( .A1(n3780), .A2(n4588), .ZN(n4291) );
  NAND2_X1 U2892 ( .A1(n3228), .A2(n3309), .ZN(n3229) );
  NAND2_X1 U2893 ( .A1(n3009), .A2(n2725), .ZN(n4530) );
  NOR2_X1 U2894 ( .A1(n2464), .A2(n2463), .ZN(n2493) );
  OR2_X1 U2895 ( .A1(n2502), .A2(n2501), .ZN(n2513) );
  OR2_X1 U2896 ( .A1(n2540), .A2(n2539), .ZN(n2548) );
  NAND2_X1 U2897 ( .A1(n2458), .A2(REG3_REG_6__SCAN_IN), .ZN(n2464) );
  AND2_X1 U2898 ( .A1(n2679), .A2(n2678), .ZN(n4273) );
  AND4_X1 U2899 ( .A1(n2553), .A2(n2552), .A3(n2551), .A4(n2550), .ZN(n3769)
         );
  AND2_X1 U2900 ( .A1(n2383), .A2(n2381), .ZN(n4426) );
  OR2_X1 U2901 ( .A1(n3457), .A2(n3881), .ZN(n4230) );
  INV_X1 U2902 ( .A(n4239), .ZN(n4159) );
  NAND2_X1 U2903 ( .A1(n2773), .A2(n4508), .ZN(n4511) );
  AND2_X1 U2904 ( .A1(n2749), .A2(n2748), .ZN(n2838) );
  INV_X1 U2905 ( .A(n4332), .ZN(n3699) );
  AND2_X1 U2906 ( .A1(n3115), .A2(n3020), .ZN(n4537) );
  INV_X1 U2907 ( .A(n4530), .ZN(n4536) );
  XNOR2_X1 U2908 ( .A(n2245), .B(IR_REG_12__SCAN_IN), .ZN(n4464) );
  NAND2_X1 U2909 ( .A1(n2867), .A2(n2866), .ZN(n3759) );
  INV_X1 U2910 ( .A(n4273), .ZN(n4061) );
  INV_X1 U2911 ( .A(n3965), .ZN(n3951) );
  INV_X1 U2912 ( .A(n3439), .ZN(n3957) );
  NAND2_X1 U2913 ( .A1(n2387), .A2(n2386), .ZN(n2388) );
  NAND2_X1 U2914 ( .A1(n4215), .A2(n3120), .ZN(n4239) );
  INV_X1 U2915 ( .A(n4511), .ZN(n4520) );
  OR2_X1 U2916 ( .A1(n4027), .A2(n4343), .ZN(n2752) );
  INV_X1 U2917 ( .A(n4552), .ZN(n4549) );
  OR2_X1 U2918 ( .A1(n4027), .A2(n4404), .ZN(n2757) );
  NAND2_X1 U2919 ( .A1(n4546), .A2(n4352), .ZN(n4404) );
  INV_X1 U2920 ( .A(n4546), .ZN(n4544) );
  INV_X1 U2921 ( .A(n2725), .ZN(n4409) );
  NAND2_X1 U2922 ( .A1(n2236), .A2(n2297), .ZN(n2303) );
  NOR2_X1 U2923 ( .A1(n2303), .A2(IR_REG_16__SCAN_IN), .ZN(n2228) );
  NAND2_X1 U2924 ( .A1(n2292), .A2(n2228), .ZN(n2233) );
  INV_X1 U2925 ( .A(n2233), .ZN(n2230) );
  NAND2_X1 U2926 ( .A1(n2230), .A2(n2229), .ZN(n2605) );
  NAND2_X1 U2927 ( .A1(n2605), .A2(IR_REG_31__SCAN_IN), .ZN(n2231) );
  XNOR2_X1 U2928 ( .A(n2231), .B(IR_REG_18__SCAN_IN), .ZN(n4003) );
  INV_X1 U2929 ( .A(n4003), .ZN(n4523) );
  INV_X1 U2930 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2232) );
  AOI22_X1 U2931 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4523), .B1(n4003), .B2(
        n2232), .ZN(n2347) );
  NAND2_X1 U2932 ( .A1(n2233), .A2(IR_REG_31__SCAN_IN), .ZN(n2234) );
  MUX2_X1 U2933 ( .A(IR_REG_31__SCAN_IN), .B(n2234), .S(IR_REG_17__SCAN_IN), 
        .Z(n2235) );
  AND2_X1 U2934 ( .A1(n2605), .A2(n2235), .ZN(n2784) );
  NAND2_X1 U2935 ( .A1(n2292), .A2(n2236), .ZN(n2237) );
  NAND2_X1 U2936 ( .A1(n2237), .A2(IR_REG_31__SCAN_IN), .ZN(n2298) );
  XNOR2_X1 U2937 ( .A(n2298), .B(IR_REG_15__SCAN_IN), .ZN(n2564) );
  INV_X1 U2938 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4478) );
  OR2_X1 U2939 ( .A1(n2292), .A2(n3493), .ZN(n2238) );
  XNOR2_X1 U2940 ( .A(n2238), .B(IR_REG_14__SCAN_IN), .ZN(n2554) );
  NAND2_X1 U2941 ( .A1(n2269), .A2(n2240), .ZN(n2248) );
  INV_X1 U2942 ( .A(IR_REG_10__SCAN_IN), .ZN(n2241) );
  NAND2_X1 U2943 ( .A1(n2282), .A2(n2241), .ZN(n2242) );
  NAND2_X1 U2944 ( .A1(n2242), .A2(IR_REG_31__SCAN_IN), .ZN(n2246) );
  INV_X1 U2945 ( .A(IR_REG_11__SCAN_IN), .ZN(n2243) );
  NAND2_X1 U2946 ( .A1(n2246), .A2(n2243), .ZN(n2244) );
  NAND2_X1 U2947 ( .A1(n2244), .A2(IR_REG_31__SCAN_IN), .ZN(n2245) );
  NAND2_X1 U2948 ( .A1(REG2_REG_11__SCAN_IN), .A2(n2529), .ZN(n2287) );
  INV_X1 U2949 ( .A(n2529), .ZN(n4527) );
  INV_X1 U2950 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U2951 ( .A1(REG2_REG_11__SCAN_IN), .A2(n2529), .B1(n4527), .B2(
        n3292), .ZN(n4458) );
  OR2_X1 U2952 ( .A1(n2282), .A2(n3493), .ZN(n2247) );
  NAND2_X1 U2953 ( .A1(n2248), .A2(IR_REG_31__SCAN_IN), .ZN(n2274) );
  XNOR2_X1 U2954 ( .A(n2274), .B(IR_REG_7__SCAN_IN), .ZN(n2825) );
  INV_X1 U2955 ( .A(n2258), .ZN(n2249) );
  NAND2_X1 U2956 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2251)
         );
  INV_X1 U2957 ( .A(n3971), .ZN(n4416) );
  NAND2_X1 U2958 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3970) );
  INV_X1 U2959 ( .A(n3970), .ZN(n2256) );
  NAND2_X1 U2960 ( .A1(n3971), .A2(n2254), .ZN(n2255) );
  AOI21_X1 U2961 ( .B1(n4416), .B2(REG2_REG_1__SCAN_IN), .A(n3972), .ZN(n2912)
         );
  MUX2_X1 U2962 ( .A(n4245), .B(REG2_REG_2__SCAN_IN), .S(n4415), .Z(n2911) );
  NAND2_X1 U2963 ( .A1(n2258), .A2(IR_REG_31__SCAN_IN), .ZN(n2260) );
  XNOR2_X1 U2964 ( .A(n2260), .B(IR_REG_3__SCAN_IN), .ZN(n4414) );
  INV_X1 U2965 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3238) );
  NAND2_X1 U2966 ( .A1(n2260), .A2(n2259), .ZN(n2261) );
  NAND2_X1 U2967 ( .A1(n2261), .A2(IR_REG_31__SCAN_IN), .ZN(n2262) );
  XNOR2_X1 U2968 ( .A(n2262), .B(IR_REG_4__SCAN_IN), .ZN(n4413) );
  INV_X1 U2969 ( .A(n4413), .ZN(n2940) );
  XNOR2_X1 U2970 ( .A(n2263), .B(n2940), .ZN(n2934) );
  AND2_X1 U2971 ( .A1(n2263), .A2(n4413), .ZN(n2264) );
  NAND2_X1 U2972 ( .A1(n2239), .A2(IR_REG_31__SCAN_IN), .ZN(n2266) );
  XNOR2_X1 U2973 ( .A(n2266), .B(n2265), .ZN(n2806) );
  MUX2_X1 U2974 ( .A(REG2_REG_5__SCAN_IN), .B(n2267), .S(n2806), .Z(n2803) );
  OR2_X1 U2975 ( .A1(n2269), .A2(n3493), .ZN(n2270) );
  XNOR2_X1 U2976 ( .A(n2270), .B(IR_REG_6__SCAN_IN), .ZN(n4412) );
  XNOR2_X1 U2977 ( .A(n2271), .B(n4412), .ZN(n2814) );
  INV_X1 U2978 ( .A(n2271), .ZN(n2272) );
  INV_X1 U2979 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3123) );
  MUX2_X1 U2980 ( .A(n3123), .B(REG2_REG_7__SCAN_IN), .S(n2825), .Z(n2831) );
  NOR2_X1 U2981 ( .A1(n2832), .A2(n2831), .ZN(n2830) );
  AOI21_X1 U2982 ( .B1(n2825), .B2(REG2_REG_7__SCAN_IN), .A(n2830), .ZN(n2278)
         );
  NAND2_X1 U2983 ( .A1(n2274), .A2(n2273), .ZN(n2275) );
  NAND2_X1 U2984 ( .A1(n2275), .A2(IR_REG_31__SCAN_IN), .ZN(n2277) );
  INV_X1 U2985 ( .A(IR_REG_8__SCAN_IN), .ZN(n2276) );
  XNOR2_X1 U2986 ( .A(n2277), .B(n2276), .ZN(n4411) );
  INV_X1 U2987 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4510) );
  INV_X1 U2988 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2504) );
  NAND2_X1 U2989 ( .A1(n2279), .A2(IR_REG_31__SCAN_IN), .ZN(n2280) );
  MUX2_X1 U2990 ( .A(IR_REG_31__SCAN_IN), .B(n2280), .S(IR_REG_9__SCAN_IN), 
        .Z(n2281) );
  INV_X1 U2991 ( .A(n2281), .ZN(n2283) );
  MUX2_X1 U2992 ( .A(REG2_REG_9__SCAN_IN), .B(n2504), .S(n2791), .Z(n4432) );
  NAND2_X1 U2993 ( .A1(n4443), .A2(n2285), .ZN(n2286) );
  NAND2_X1 U2994 ( .A1(n4464), .A2(n2289), .ZN(n2290) );
  NOR2_X1 U2995 ( .A1(n2309), .A2(n3493), .ZN(n2291) );
  MUX2_X1 U2996 ( .A(n3493), .B(n2291), .S(IR_REG_13__SCAN_IN), .Z(n2293) );
  OR2_X1 U2997 ( .A1(n2293), .A2(n2292), .ZN(n3258) );
  INV_X1 U2998 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3249) );
  NOR2_X1 U2999 ( .A1(n3258), .A2(n3249), .ZN(n3248) );
  INV_X1 U3000 ( .A(n3258), .ZN(n2781) );
  OAI22_X1 U3001 ( .A1(n3251), .A2(n3248), .B1(REG2_REG_13__SCAN_IN), .B2(
        n2781), .ZN(n2294) );
  NOR2_X1 U3002 ( .A1(n2146), .A2(n2294), .ZN(n2295) );
  NAND2_X1 U3003 ( .A1(REG2_REG_15__SCAN_IN), .A2(n2564), .ZN(n2296) );
  OAI21_X1 U3004 ( .B1(REG2_REG_15__SCAN_IN), .B2(n2564), .A(n2296), .ZN(n4486) );
  AOI21_X1 U3005 ( .B1(n2564), .B2(REG2_REG_15__SCAN_IN), .A(n4485), .ZN(n2301) );
  NAND2_X1 U3006 ( .A1(n2298), .A2(n2297), .ZN(n2299) );
  NAND2_X1 U3007 ( .A1(n2299), .A2(IR_REG_31__SCAN_IN), .ZN(n2300) );
  XNOR2_X1 U3008 ( .A(n2300), .B(IR_REG_16__SCAN_IN), .ZN(n2575) );
  INV_X1 U3009 ( .A(n2575), .ZN(n4524) );
  NAND2_X1 U3010 ( .A1(n2301), .A2(n4524), .ZN(n2302) );
  XNOR2_X1 U3011 ( .A(n2301), .B(n2575), .ZN(n4498) );
  INV_X1 U3012 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4496) );
  NAND2_X1 U3013 ( .A1(n2302), .A2(n4497), .ZN(n3992) );
  INV_X1 U3014 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2586) );
  XNOR2_X1 U3015 ( .A(n2784), .B(n2586), .ZN(n3994) );
  NAND2_X1 U3016 ( .A1(n3992), .A2(n3994), .ZN(n3993) );
  INV_X1 U3017 ( .A(n2303), .ZN(n2307) );
  INV_X1 U3018 ( .A(n2335), .ZN(n2311) );
  INV_X1 U3019 ( .A(IR_REG_22__SCAN_IN), .ZN(n2310) );
  NAND2_X1 U3020 ( .A1(n2311), .A2(n2310), .ZN(n2314) );
  INV_X1 U3021 ( .A(n2318), .ZN(n2313) );
  OAI21_X1 U3022 ( .B1(n2314), .B2(n2313), .A(IR_REG_31__SCAN_IN), .ZN(n2315)
         );
  NAND2_X1 U3023 ( .A1(n2323), .A2(IR_REG_31__SCAN_IN), .ZN(n2322) );
  MUX2_X1 U3024 ( .A(IR_REG_31__SCAN_IN), .B(n2322), .S(IR_REG_26__SCAN_IN), 
        .Z(n2325) );
  INV_X1 U3025 ( .A(n2339), .ZN(n2324) );
  OR2_X1 U3026 ( .A1(n2327), .A2(n2326), .ZN(n2328) );
  NAND2_X1 U3027 ( .A1(n2329), .A2(n2328), .ZN(n2337) );
  INV_X1 U3028 ( .A(n2864), .ZN(n2331) );
  INV_X1 U3029 ( .A(n2337), .ZN(n2330) );
  NAND2_X1 U3030 ( .A1(n2330), .A2(STATE_REG_SCAN_IN), .ZN(n3947) );
  NAND2_X1 U3031 ( .A1(n2331), .A2(n3947), .ZN(n2383) );
  INV_X1 U3032 ( .A(n2320), .ZN(n2332) );
  NAND2_X1 U3033 ( .A1(n2332), .A2(IR_REG_31__SCAN_IN), .ZN(n2333) );
  MUX2_X1 U3034 ( .A(IR_REG_31__SCAN_IN), .B(n2333), .S(IR_REG_21__SCAN_IN), 
        .Z(n2334) );
  NAND2_X1 U3035 ( .A1(n2334), .A2(n2335), .ZN(n2771) );
  NAND2_X1 U3036 ( .A1(n2335), .A2(IR_REG_31__SCAN_IN), .ZN(n2336) );
  AND2_X1 U3037 ( .A1(n2841), .A2(n2337), .ZN(n2341) );
  NAND2_X1 U3038 ( .A1(n2338), .A2(n3493), .ZN(n2340) );
  NOR2_X1 U3039 ( .A1(n2339), .A2(n2213), .ZN(n2344) );
  MUX2_X2 U3040 ( .A(n2345), .B(n2344), .S(IR_REG_28__SCAN_IN), .Z(n2439) );
  NOR2_X1 U3041 ( .A1(n2341), .A2(n3780), .ZN(n2381) );
  NAND2_X1 U3042 ( .A1(n2342), .A2(IR_REG_31__SCAN_IN), .ZN(n2343) );
  XNOR2_X1 U3043 ( .A(n2343), .B(n2208), .ZN(n4418) );
  INV_X1 U3044 ( .A(n4418), .ZN(n2906) );
  NOR2_X1 U3045 ( .A1(n2345), .A2(n2344), .ZN(n4424) );
  AND2_X1 U3046 ( .A1(n2906), .A2(n4424), .ZN(n3943) );
  AOI211_X1 U3047 ( .C1(n2347), .C2(n2346), .A(n4002), .B(n4495), .ZN(n2389)
         );
  INV_X1 U3048 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U3049 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4003), .B1(n4523), .B2(
        n4006), .ZN(n2380) );
  NOR2_X1 U3050 ( .A1(n2784), .A2(REG1_REG_17__SCAN_IN), .ZN(n2377) );
  NAND2_X1 U3051 ( .A1(REG1_REG_15__SCAN_IN), .A2(n2564), .ZN(n2372) );
  INV_X1 U3052 ( .A(n2564), .ZN(n4525) );
  INV_X1 U3053 ( .A(REG1_REG_15__SCAN_IN), .ZN(n2348) );
  AOI22_X1 U3054 ( .A1(REG1_REG_15__SCAN_IN), .A2(n2564), .B1(n4525), .B2(
        n2348), .ZN(n4491) );
  INV_X1 U3055 ( .A(REG1_REG_13__SCAN_IN), .ZN(n2542) );
  NOR2_X1 U3056 ( .A1(n3258), .A2(n2542), .ZN(n2349) );
  INV_X1 U3057 ( .A(n2349), .ZN(n2369) );
  AOI21_X1 U3058 ( .B1(n2542), .B2(n3258), .A(n2349), .ZN(n3254) );
  NAND2_X1 U3059 ( .A1(REG1_REG_11__SCAN_IN), .A2(n2529), .ZN(n2366) );
  INV_X1 U3060 ( .A(REG1_REG_11__SCAN_IN), .ZN(n2350) );
  AOI22_X1 U3061 ( .A1(REG1_REG_11__SCAN_IN), .A2(n2529), .B1(n4527), .B2(
        n2350), .ZN(n4455) );
  NAND2_X1 U3062 ( .A1(n2791), .A2(REG1_REG_9__SCAN_IN), .ZN(n2363) );
  INV_X1 U3063 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2351) );
  MUX2_X1 U3064 ( .A(n2351), .B(REG1_REG_9__SCAN_IN), .S(n2791), .Z(n2352) );
  INV_X1 U3065 ( .A(n2352), .ZN(n4435) );
  INV_X1 U3066 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2451) );
  INV_X1 U3067 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2964) );
  XNOR2_X1 U3068 ( .A(n4415), .B(n2964), .ZN(n2915) );
  XNOR2_X1 U3069 ( .A(n3971), .B(REG1_REG_1__SCAN_IN), .ZN(n3969) );
  AND2_X1 U3070 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3968)
         );
  NAND2_X1 U3071 ( .A1(n3969), .A2(n3968), .ZN(n3967) );
  NAND2_X1 U3072 ( .A1(n4416), .A2(REG1_REG_1__SCAN_IN), .ZN(n2353) );
  NAND2_X1 U3073 ( .A1(n3967), .A2(n2353), .ZN(n2914) );
  NAND2_X1 U3074 ( .A1(n2915), .A2(n2914), .ZN(n2913) );
  NAND2_X1 U3075 ( .A1(n4415), .A2(REG1_REG_2__SCAN_IN), .ZN(n2354) );
  NAND2_X1 U3076 ( .A1(n2913), .A2(n2354), .ZN(n2356) );
  XNOR2_X1 U3077 ( .A(n2356), .B(n2355), .ZN(n3981) );
  NAND2_X1 U3078 ( .A1(n3981), .A2(REG1_REG_3__SCAN_IN), .ZN(n3980) );
  NAND2_X1 U3079 ( .A1(n2356), .A2(n4414), .ZN(n2357) );
  NAND2_X1 U3080 ( .A1(n3980), .A2(n2357), .ZN(n2358) );
  INV_X1 U3081 ( .A(n2358), .ZN(n2359) );
  XNOR2_X1 U3082 ( .A(n2358), .B(n2940), .ZN(n2936) );
  NAND2_X1 U3083 ( .A1(n2936), .A2(REG1_REG_4__SCAN_IN), .ZN(n2935) );
  XNOR2_X1 U3084 ( .A(n2806), .B(REG1_REG_5__SCAN_IN), .ZN(n2811) );
  INV_X1 U3085 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2817) );
  NOR2_X1 U3086 ( .A1(n2818), .A2(n2817), .ZN(n2815) );
  NOR2_X1 U3087 ( .A1(n2825), .A2(REG1_REG_7__SCAN_IN), .ZN(n2361) );
  INV_X1 U3088 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4550) );
  INV_X1 U3089 ( .A(n2825), .ZN(n2829) );
  INV_X1 U3090 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2492) );
  NAND2_X1 U3091 ( .A1(n2363), .A2(n4434), .ZN(n2364) );
  NAND2_X1 U3092 ( .A1(n4443), .A2(n2364), .ZN(n2365) );
  XOR2_X1 U3093 ( .A(n2364), .B(n4443), .Z(n4450) );
  NAND2_X1 U3094 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4450), .ZN(n4449) );
  NAND2_X1 U3095 ( .A1(n4464), .A2(n2367), .ZN(n2368) );
  NAND2_X1 U3096 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4472), .ZN(n4471) );
  NAND2_X1 U3097 ( .A1(n2554), .A2(n2370), .ZN(n2371) );
  NAND2_X1 U3098 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4482), .ZN(n4481) );
  NAND2_X1 U3099 ( .A1(n2371), .A2(n4481), .ZN(n4490) );
  NAND2_X1 U3100 ( .A1(n4491), .A2(n4490), .ZN(n4489) );
  NAND2_X1 U3101 ( .A1(n2372), .A2(n4489), .ZN(n2373) );
  NOR2_X1 U3102 ( .A1(n2575), .A2(n2373), .ZN(n2374) );
  XNOR2_X1 U3103 ( .A(n2373), .B(n2575), .ZN(n4503) );
  NOR2_X1 U3104 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4503), .ZN(n4504) );
  NOR2_X1 U3105 ( .A1(n2374), .A2(n4504), .ZN(n3989) );
  INV_X1 U3106 ( .A(REG1_REG_17__SCAN_IN), .ZN(n2376) );
  INV_X1 U3107 ( .A(n2784), .ZN(n4001) );
  INV_X1 U3108 ( .A(n2377), .ZN(n2375) );
  OAI21_X1 U3109 ( .B1(n2376), .B2(n4001), .A(n2375), .ZN(n3988) );
  INV_X1 U3110 ( .A(n4424), .ZN(n2378) );
  OAI211_X1 U3111 ( .C1(n2380), .C2(n2379), .A(n4502), .B(n4005), .ZN(n2387)
         );
  NAND2_X1 U3112 ( .A1(n4426), .A2(n4418), .ZN(n4507) );
  INV_X1 U3113 ( .A(n2381), .ZN(n2382) );
  NOR2_X1 U3114 ( .A1(n2577), .A2(STATE_REG_SCAN_IN), .ZN(n3744) );
  AOI21_X1 U3115 ( .B1(n4501), .B2(ADDR_REG_18__SCAN_IN), .A(n3744), .ZN(n2384) );
  INV_X1 U3116 ( .A(n2385), .ZN(n2386) );
  OR2_X1 U3117 ( .A1(n2389), .A2(n2388), .ZN(U3258) );
  INV_X1 U3118 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2750) );
  INV_X1 U3119 ( .A(DATAI_27_), .ZN(n2390) );
  NAND2_X1 U3120 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2391) );
  INV_X1 U3121 ( .A(REG3_REG_25__SCAN_IN), .ZN(n2409) );
  INV_X1 U3122 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3751) );
  INV_X1 U3123 ( .A(n2663), .ZN(n2394) );
  NAND2_X1 U3124 ( .A1(n2394), .A2(REG3_REG_27__SCAN_IN), .ZN(n2673) );
  INV_X1 U3125 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4640) );
  NAND2_X1 U3126 ( .A1(n2663), .A2(n4640), .ZN(n2395) );
  NAND2_X1 U3127 ( .A1(n2673), .A2(n2395), .ZN(n4055) );
  OR2_X1 U3128 ( .A1(n4055), .A2(n2680), .ZN(n2407) );
  INV_X1 U3129 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4276) );
  NAND2_X1 U3130 ( .A1(n2455), .A2(REG2_REG_27__SCAN_IN), .ZN(n2404) );
  INV_X1 U3131 ( .A(n4407), .ZN(n2402) );
  INV_X2 U3132 ( .A(n2425), .ZN(n2470) );
  NAND2_X1 U3133 ( .A1(n2470), .A2(REG0_REG_27__SCAN_IN), .ZN(n2403) );
  OAI211_X1 U3134 ( .C1(n4276), .C2(n2471), .A(n2404), .B(n2403), .ZN(n2405)
         );
  INV_X1 U3135 ( .A(n2405), .ZN(n2406) );
  INV_X1 U3136 ( .A(DATAI_25_), .ZN(n2408) );
  NAND2_X1 U3137 ( .A1(n2651), .A2(n2409), .ZN(n2410) );
  NAND2_X1 U3138 ( .A1(n2661), .A2(n2410), .ZN(n4093) );
  OR2_X1 U3139 ( .A1(n4093), .A2(n2680), .ZN(n2415) );
  INV_X1 U3140 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4289) );
  NAND2_X1 U3141 ( .A1(n2470), .A2(REG0_REG_25__SCAN_IN), .ZN(n2412) );
  NAND2_X1 U3142 ( .A1(n2455), .A2(REG2_REG_25__SCAN_IN), .ZN(n2411) );
  OAI211_X1 U3143 ( .C1(n4289), .C2(n2471), .A(n2412), .B(n2411), .ZN(n2413)
         );
  INV_X1 U3144 ( .A(n2413), .ZN(n2414) );
  INV_X1 U3145 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2416) );
  INV_X1 U3146 ( .A(n2434), .ZN(n2417) );
  NAND2_X1 U3147 ( .A1(n2417), .A2(REG2_REG_1__SCAN_IN), .ZN(n2422) );
  INV_X1 U31480 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2418) );
  OR2_X1 U31490 ( .A1(n2425), .A2(n2418), .ZN(n2421) );
  INV_X1 U3150 ( .A(n2432), .ZN(n2419) );
  NAND2_X1 U3151 ( .A1(n2419), .A2(REG3_REG_1__SCAN_IN), .ZN(n2420) );
  INV_X1 U3152 ( .A(n2880), .ZN(n4247) );
  MUX2_X1 U3153 ( .A(DATAI_1_), .B(n4416), .S(n2439), .Z(n2929) );
  INV_X1 U3154 ( .A(n2929), .ZN(n2876) );
  NAND2_X1 U3155 ( .A1(n4247), .A2(n2876), .ZN(n3800) );
  NAND2_X1 U3156 ( .A1(n2880), .A2(n2929), .ZN(n3803) );
  INV_X1 U3157 ( .A(n2433), .ZN(n2579) );
  INV_X1 U3158 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3011) );
  OR2_X1 U3159 ( .A1(n2434), .A2(n3011), .ZN(n2428) );
  INV_X1 U3160 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3010) );
  INV_X1 U3161 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2424) );
  OR2_X1 U3162 ( .A1(n2425), .A2(n2424), .ZN(n2426) );
  MUX2_X1 U3163 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(n2439), .Z(n3007) );
  AND2_X1 U3164 ( .A1(n3966), .A2(n3007), .ZN(n2762) );
  NAND2_X1 U3165 ( .A1(n2763), .A2(n2762), .ZN(n2761) );
  NAND2_X1 U3166 ( .A1(n4247), .A2(n2929), .ZN(n2430) );
  NAND2_X1 U3167 ( .A1(n2761), .A2(n2430), .ZN(n2953) );
  INV_X1 U3168 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2431) );
  INV_X1 U3169 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2917) );
  OR2_X1 U3170 ( .A1(n2432), .A2(n2917), .ZN(n2437) );
  OR2_X1 U3171 ( .A1(n2433), .A2(n2964), .ZN(n2436) );
  INV_X1 U3172 ( .A(REG2_REG_2__SCAN_IN), .ZN(n4245) );
  OR2_X1 U3173 ( .A1(n2434), .A2(n4245), .ZN(n2435) );
  MUX2_X1 U3174 ( .A(DATAI_2_), .B(n4415), .S(n2439), .Z(n4251) );
  NAND2_X1 U3175 ( .A1(n2978), .A2(n4251), .ZN(n3804) );
  INV_X1 U3176 ( .A(n2978), .ZN(n3964) );
  NAND2_X1 U3177 ( .A1(n3964), .A2(n2962), .ZN(n3807) );
  OR2_X2 U3178 ( .A1(n2953), .A2(n3892), .ZN(n3016) );
  INV_X1 U3179 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2440) );
  OR2_X1 U3180 ( .A1(n2471), .A2(n2440), .ZN(n2442) );
  NAND2_X1 U3181 ( .A1(n2455), .A2(REG2_REG_4__SCAN_IN), .ZN(n2441) );
  INV_X1 U3182 ( .A(n2443), .ZN(n2452) );
  INV_X1 U3183 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2445) );
  INV_X1 U3184 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2444) );
  NAND2_X1 U3185 ( .A1(n2445), .A2(n2444), .ZN(n2446) );
  NAND2_X1 U3186 ( .A1(n2452), .A2(n2446), .ZN(n3043) );
  OR2_X1 U3187 ( .A1(n2680), .A2(n3043), .ZN(n2449) );
  INV_X1 U3188 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2447) );
  OR2_X1 U3189 ( .A1(n2425), .A2(n2447), .ZN(n2448) );
  MUX2_X1 U3190 ( .A(DATAI_4_), .B(n4413), .S(n2609), .Z(n3050) );
  OR2_X1 U3191 ( .A1(n2471), .A2(n2451), .ZN(n2484) );
  NAND2_X1 U3192 ( .A1(n2470), .A2(REG0_REG_5__SCAN_IN), .ZN(n2483) );
  INV_X1 U3193 ( .A(n2458), .ZN(n2454) );
  NAND2_X1 U3194 ( .A1(n2452), .A2(n4656), .ZN(n2453) );
  NAND2_X1 U3195 ( .A1(n2454), .A2(n2453), .ZN(n3205) );
  OR2_X1 U3196 ( .A1(n2680), .A2(n3205), .ZN(n2482) );
  OR2_X1 U3197 ( .A1(n2401), .A2(n2267), .ZN(n2481) );
  NAND4_X1 U3198 ( .A1(n2484), .A2(n2483), .A3(n2482), .A4(n2481), .ZN(n2694)
         );
  INV_X1 U3199 ( .A(DATAI_5_), .ZN(n2456) );
  AND2_X1 U3200 ( .A1(n3031), .A2(n2457), .ZN(n3063) );
  NAND2_X1 U3201 ( .A1(n2470), .A2(REG0_REG_6__SCAN_IN), .ZN(n2462) );
  INV_X1 U3202 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3215) );
  OR2_X1 U3203 ( .A1(n2401), .A2(n3215), .ZN(n2461) );
  OAI21_X1 U3204 ( .B1(n2458), .B2(REG3_REG_6__SCAN_IN), .A(n2464), .ZN(n3214)
         );
  OR2_X1 U3205 ( .A1(n2680), .A2(n3214), .ZN(n2460) );
  OR2_X1 U3206 ( .A1(n2471), .A2(n2817), .ZN(n2459) );
  MUX2_X1 U3207 ( .A(DATAI_6_), .B(n4412), .S(n2609), .Z(n3218) );
  OR2_X1 U3208 ( .A1(n2471), .A2(n4550), .ZN(n2469) );
  NAND2_X1 U3209 ( .A1(n2470), .A2(REG0_REG_7__SCAN_IN), .ZN(n2468) );
  AND2_X1 U32100 ( .A1(n2464), .A2(n2463), .ZN(n2465) );
  OR2_X1 U32110 ( .A1(n2465), .A2(n2493), .ZN(n3183) );
  OR2_X1 U32120 ( .A1(n2680), .A2(n3183), .ZN(n2467) );
  OR2_X1 U32130 ( .A1(n2401), .A2(n3123), .ZN(n2466) );
  MUX2_X1 U32140 ( .A(DATAI_7_), .B(n2825), .S(n2609), .Z(n3152) );
  INV_X2 U32150 ( .A(n3963), .ZN(n3240) );
  NAND2_X1 U32160 ( .A1(n3240), .A2(n3050), .ZN(n3810) );
  NAND2_X1 U32170 ( .A1(n3963), .A2(n3047), .ZN(n3814) );
  NAND2_X1 U32180 ( .A1(n2978), .A2(n2962), .ZN(n2988) );
  NAND2_X1 U32190 ( .A1(n2470), .A2(REG0_REG_3__SCAN_IN), .ZN(n2475) );
  OR2_X1 U32200 ( .A1(n2680), .A2(REG3_REG_3__SCAN_IN), .ZN(n2474) );
  INV_X1 U32210 ( .A(REG1_REG_3__SCAN_IN), .ZN(n3000) );
  OR2_X1 U32220 ( .A1(n2471), .A2(n3000), .ZN(n2473) );
  OR2_X1 U32230 ( .A1(n2401), .A2(n3238), .ZN(n2472) );
  INV_X1 U32240 ( .A(n4253), .ZN(n2977) );
  NAND2_X1 U32250 ( .A1(n2977), .A2(n3239), .ZN(n2478) );
  AND2_X1 U32260 ( .A1(n2988), .A2(n2478), .ZN(n3015) );
  NAND2_X1 U32270 ( .A1(n4253), .A2(n2995), .ZN(n3017) );
  NAND2_X1 U32280 ( .A1(n2479), .A2(n2217), .ZN(n2490) );
  NAND2_X1 U32290 ( .A1(n3221), .A2(n3152), .ZN(n2695) );
  INV_X1 U32300 ( .A(n3152), .ZN(n3177) );
  NAND2_X1 U32310 ( .A1(n2695), .A2(n3821), .ZN(n3117) );
  NAND2_X1 U32320 ( .A1(n3084), .A2(n3090), .ZN(n3064) );
  INV_X1 U32330 ( .A(n3064), .ZN(n2485) );
  NAND2_X1 U32340 ( .A1(n2486), .A2(n2485), .ZN(n2488) );
  NAND2_X1 U32350 ( .A1(n3178), .A2(n3101), .ZN(n2487) );
  AND2_X1 U32360 ( .A1(n2488), .A2(n2487), .ZN(n3116) );
  AOI21_X2 U32370 ( .B1(n2491), .B2(n2490), .A(n2489), .ZN(n3128) );
  NAND2_X1 U32380 ( .A1(n2470), .A2(REG0_REG_8__SCAN_IN), .ZN(n2498) );
  OR2_X1 U32390 ( .A1(n2471), .A2(n2492), .ZN(n2497) );
  OR2_X1 U32400 ( .A1(n2493), .A2(REG3_REG_8__SCAN_IN), .ZN(n2494) );
  NAND2_X1 U32410 ( .A1(n2502), .A2(n2494), .ZN(n4509) );
  OR2_X1 U32420 ( .A1(n2680), .A2(n4509), .ZN(n2496) );
  OR2_X1 U32430 ( .A1(n2401), .A2(n4510), .ZN(n2495) );
  INV_X1 U32440 ( .A(DATAI_8_), .ZN(n4670) );
  MUX2_X1 U32450 ( .A(n4670), .B(n4411), .S(n2609), .Z(n3168) );
  NAND2_X1 U32460 ( .A1(n3269), .A2(n3168), .ZN(n2499) );
  INV_X1 U32470 ( .A(n3269), .ZN(n3960) );
  NAND2_X1 U32480 ( .A1(n3960), .A2(n3159), .ZN(n2500) );
  NAND2_X1 U32490 ( .A1(n2470), .A2(REG0_REG_9__SCAN_IN), .ZN(n2508) );
  NAND2_X1 U32500 ( .A1(n2502), .A2(n2501), .ZN(n2503) );
  NAND2_X1 U32510 ( .A1(n2513), .A2(n2503), .ZN(n3273) );
  OR2_X1 U32520 ( .A1(n2680), .A2(n3273), .ZN(n2507) );
  OR2_X1 U32530 ( .A1(n2471), .A2(n2351), .ZN(n2506) );
  OR2_X1 U32540 ( .A1(n2401), .A2(n2504), .ZN(n2505) );
  NAND4_X1 U32550 ( .A1(n2508), .A2(n2507), .A3(n2506), .A4(n2505), .ZN(n3959)
         );
  MUX2_X1 U32560 ( .A(DATAI_9_), .B(n2791), .S(n2609), .Z(n3263) );
  AND2_X1 U32570 ( .A1(n3959), .A2(n3263), .ZN(n2509) );
  NAND2_X1 U32580 ( .A1(n3310), .A2(n3268), .ZN(n2510) );
  NAND2_X1 U32590 ( .A1(n2470), .A2(REG0_REG_10__SCAN_IN), .ZN(n2519) );
  INV_X1 U32600 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2511) );
  OR2_X1 U32610 ( .A1(n2471), .A2(n2511), .ZN(n2518) );
  INV_X1 U32620 ( .A(n2512), .ZN(n2523) );
  NAND2_X1 U32630 ( .A1(n2513), .A2(n4658), .ZN(n2514) );
  NAND2_X1 U32640 ( .A1(n2523), .A2(n2514), .ZN(n3315) );
  OR2_X1 U32650 ( .A1(n2680), .A2(n3315), .ZN(n2517) );
  INV_X1 U32660 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2515) );
  OR2_X1 U32670 ( .A1(n2401), .A2(n2515), .ZN(n2516) );
  MUX2_X1 U32680 ( .A(DATAI_10_), .B(n4443), .S(n2609), .Z(n3302) );
  NOR2_X1 U32690 ( .A1(n3958), .A2(n3302), .ZN(n2520) );
  NAND2_X1 U32700 ( .A1(n2470), .A2(REG0_REG_11__SCAN_IN), .ZN(n2528) );
  OR2_X1 U32710 ( .A1(n2471), .A2(n2350), .ZN(n2527) );
  INV_X1 U32720 ( .A(n2521), .ZN(n2532) );
  INV_X1 U32730 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U32740 ( .A1(n2523), .A2(n2522), .ZN(n2524) );
  NAND2_X1 U32750 ( .A1(n2532), .A2(n2524), .ZN(n3392) );
  OR2_X1 U32760 ( .A1(n2680), .A2(n3392), .ZN(n2526) );
  OR2_X1 U32770 ( .A1(n2401), .A2(n3292), .ZN(n2525) );
  MUX2_X1 U32780 ( .A(DATAI_11_), .B(n2529), .S(n3780), .Z(n3287) );
  NAND2_X1 U32790 ( .A1(n3439), .A2(n3287), .ZN(n3796) );
  NAND2_X1 U32800 ( .A1(n3957), .A2(n3387), .ZN(n3834) );
  NAND2_X1 U32810 ( .A1(n3439), .A2(n3387), .ZN(n2530) );
  NAND2_X1 U32820 ( .A1(n2470), .A2(REG0_REG_12__SCAN_IN), .ZN(n2538) );
  INV_X1 U32830 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3350) );
  OR2_X1 U32840 ( .A1(n2401), .A2(n3350), .ZN(n2537) );
  INV_X1 U32850 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U32860 ( .A1(n2532), .A2(n2531), .ZN(n2533) );
  NAND2_X1 U32870 ( .A1(n2540), .A2(n2533), .ZN(n3437) );
  OR2_X1 U32880 ( .A1(n2680), .A2(n3437), .ZN(n2536) );
  INV_X1 U32890 ( .A(REG1_REG_12__SCAN_IN), .ZN(n2534) );
  OR2_X1 U32900 ( .A1(n2471), .A2(n2534), .ZN(n2535) );
  NAND4_X1 U32910 ( .A1(n2538), .A2(n2537), .A3(n2536), .A4(n2535), .ZN(n3956)
         );
  MUX2_X1 U32920 ( .A(DATAI_12_), .B(n4464), .S(n3780), .Z(n3433) );
  INV_X1 U32930 ( .A(n3956), .ZN(n3487) );
  INV_X1 U32940 ( .A(n3433), .ZN(n3438) );
  NAND2_X1 U32950 ( .A1(n2470), .A2(REG0_REG_13__SCAN_IN), .ZN(n2546) );
  OR2_X1 U32960 ( .A1(n2401), .A2(n3249), .ZN(n2545) );
  NAND2_X1 U32970 ( .A1(n2540), .A2(n2539), .ZN(n2541) );
  NAND2_X1 U32980 ( .A1(n2548), .A2(n2541), .ZN(n3492) );
  OR2_X1 U32990 ( .A1(n2680), .A2(n3492), .ZN(n2544) );
  OR2_X1 U33000 ( .A1(n2471), .A2(n2542), .ZN(n2543) );
  NAND4_X1 U33010 ( .A1(n2546), .A2(n2545), .A3(n2544), .A4(n2543), .ZN(n3955)
         );
  MUX2_X1 U33020 ( .A(DATAI_13_), .B(n2781), .S(n2609), .Z(n3326) );
  NOR2_X1 U33030 ( .A1(n3955), .A2(n3326), .ZN(n2547) );
  INV_X1 U33040 ( .A(n3326), .ZN(n3486) );
  OAI22_X2 U33050 ( .A1(n3325), .A2(n2547), .B1(n3640), .B2(n3486), .ZN(n3334)
         );
  NAND2_X1 U33060 ( .A1(n2470), .A2(REG0_REG_14__SCAN_IN), .ZN(n2553) );
  INV_X1 U33070 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3413) );
  OR2_X1 U33080 ( .A1(n2471), .A2(n3413), .ZN(n2552) );
  NAND2_X1 U33090 ( .A1(n2548), .A2(n4639), .ZN(n2549) );
  NAND2_X1 U33100 ( .A1(n2557), .A2(n2549), .ZN(n3638) );
  OR2_X1 U33110 ( .A1(n2680), .A2(n3638), .ZN(n2551) );
  OR2_X1 U33120 ( .A1(n2401), .A2(n4478), .ZN(n2550) );
  MUX2_X1 U33130 ( .A(DATAI_14_), .B(n2554), .S(n2609), .Z(n3503) );
  NAND2_X1 U33140 ( .A1(n3769), .A2(n3503), .ZN(n3791) );
  INV_X1 U33150 ( .A(n3769), .ZN(n3954) );
  NAND2_X1 U33160 ( .A1(n3954), .A2(n3639), .ZN(n3789) );
  NAND2_X1 U33170 ( .A1(n3769), .A2(n3639), .ZN(n2555) );
  INV_X1 U33180 ( .A(n2556), .ZN(n2569) );
  NAND2_X1 U33190 ( .A1(n2557), .A2(n3766), .ZN(n2558) );
  NAND2_X1 U33200 ( .A1(n2569), .A2(n2558), .ZN(n3775) );
  OR2_X1 U33210 ( .A1(n2680), .A2(n3775), .ZN(n2563) );
  INV_X1 U33220 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2559) );
  OR2_X1 U33230 ( .A1(n2401), .A2(n2559), .ZN(n2562) );
  INV_X1 U33240 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3449) );
  OR2_X1 U33250 ( .A1(n2425), .A2(n3449), .ZN(n2561) );
  OR2_X1 U33260 ( .A1(n2471), .A2(n2348), .ZN(n2560) );
  NAND4_X1 U33270 ( .A1(n2563), .A2(n2562), .A3(n2561), .A4(n2560), .ZN(n3953)
         );
  MUX2_X1 U33280 ( .A(DATAI_15_), .B(n2564), .S(n2609), .Z(n3512) );
  INV_X1 U33290 ( .A(n3457), .ZN(n2594) );
  OR2_X1 U33300 ( .A1(n2401), .A2(n4496), .ZN(n2567) );
  INV_X1 U33310 ( .A(REG0_REG_16__SCAN_IN), .ZN(n2565) );
  OR2_X1 U33320 ( .A1(n2425), .A2(n2565), .ZN(n2566) );
  AND2_X1 U33330 ( .A1(n2567), .A2(n2566), .ZN(n2574) );
  INV_X1 U33340 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2568) );
  NAND2_X1 U33350 ( .A1(n2569), .A2(n2568), .ZN(n2570) );
  NAND2_X1 U33360 ( .A1(n2583), .A2(n2570), .ZN(n3471) );
  OR2_X1 U33370 ( .A1(n3471), .A2(n2680), .ZN(n2573) );
  INV_X1 U33380 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2571) );
  OR2_X1 U33390 ( .A1(n2471), .A2(n2571), .ZN(n2572) );
  MUX2_X1 U33400 ( .A(DATAI_16_), .B(n2575), .S(n3780), .Z(n4344) );
  NAND2_X1 U33410 ( .A1(n3700), .A2(n4344), .ZN(n3913) );
  INV_X1 U33420 ( .A(n4344), .ZN(n3689) );
  NAND2_X1 U33430 ( .A1(n4334), .A2(n3689), .ZN(n3788) );
  INV_X1 U33440 ( .A(n2576), .ZN(n2597) );
  NAND2_X1 U33450 ( .A1(n2585), .A2(n2577), .ZN(n2578) );
  NAND2_X1 U33460 ( .A1(n2597), .A2(n2578), .ZN(n4228) );
  OR2_X1 U33470 ( .A1(n4228), .A2(n2680), .ZN(n2582) );
  AOI22_X1 U33480 ( .A1(n2579), .A2(REG1_REG_18__SCAN_IN), .B1(n2470), .B2(
        REG0_REG_18__SCAN_IN), .ZN(n2581) );
  NAND2_X1 U33490 ( .A1(n2455), .A2(REG2_REG_18__SCAN_IN), .ZN(n2580) );
  MUX2_X1 U33500 ( .A(DATAI_18_), .B(n4003), .S(n3780), .Z(n4222) );
  NAND2_X1 U33510 ( .A1(n4338), .A2(n4222), .ZN(n4198) );
  INV_X1 U33520 ( .A(n4338), .ZN(n3952) );
  NAND2_X1 U3353 ( .A1(n3952), .A2(n4219), .ZN(n4199) );
  NAND2_X1 U33540 ( .A1(n2583), .A2(n4646), .ZN(n2584) );
  NAND2_X1 U3355 ( .A1(n2585), .A2(n2584), .ZN(n3461) );
  AOI22_X1 U3356 ( .A1(n2579), .A2(REG1_REG_17__SCAN_IN), .B1(n2470), .B2(
        REG0_REG_17__SCAN_IN), .ZN(n2588) );
  OR2_X1 U3357 ( .A1(n2401), .A2(n2586), .ZN(n2587) );
  MUX2_X1 U3358 ( .A(DATAI_17_), .B(n2784), .S(n3780), .Z(n4332) );
  OR2_X1 U3359 ( .A1(n4347), .A2(n4332), .ZN(n4231) );
  NOR2_X1 U3360 ( .A1(n4238), .A2(n4231), .ZN(n2592) );
  OR2_X1 U3361 ( .A1(n3881), .A2(n2592), .ZN(n4233) );
  AND2_X1 U3362 ( .A1(n4338), .A2(n4219), .ZN(n2593) );
  NAND2_X1 U3363 ( .A1(n4334), .A2(n4344), .ZN(n3458) );
  NAND2_X1 U3364 ( .A1(n4347), .A2(n4332), .ZN(n2589) );
  AND2_X1 U3365 ( .A1(n3458), .A2(n2589), .ZN(n4229) );
  INV_X1 U3366 ( .A(n4238), .ZN(n2590) );
  AND2_X1 U3367 ( .A1(n4229), .A2(n2590), .ZN(n2591) );
  OR2_X1 U3368 ( .A1(n2592), .A2(n2591), .ZN(n4234) );
  AOI21_X1 U3369 ( .B1(n2594), .B2(n2047), .A(n2218), .ZN(n4196) );
  INV_X1 U3370 ( .A(n2595), .ZN(n2613) );
  INV_X1 U3371 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2596) );
  NAND2_X1 U3372 ( .A1(n2597), .A2(n2596), .ZN(n2598) );
  NAND2_X1 U3373 ( .A1(n4211), .A2(n2419), .ZN(n2604) );
  INV_X1 U3374 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4327) );
  NAND2_X1 U3375 ( .A1(n2470), .A2(REG0_REG_19__SCAN_IN), .ZN(n2601) );
  INV_X1 U3376 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2599) );
  OR2_X1 U3377 ( .A1(n2401), .A2(n2599), .ZN(n2600) );
  OAI211_X1 U3378 ( .C1(n4327), .C2(n2471), .A(n2601), .B(n2600), .ZN(n2602)
         );
  INV_X1 U3379 ( .A(n2602), .ZN(n2603) );
  OAI21_X2 U3380 ( .B1(n2605), .B2(IR_REG_18__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2607) );
  OR2_X1 U3381 ( .A1(n2607), .A2(n2606), .ZN(n2608) );
  NAND2_X1 U3382 ( .A1(n2607), .A2(n2606), .ZN(n2687) );
  MUX2_X1 U3383 ( .A(DATAI_19_), .B(n4227), .S(n2609), .Z(n3539) );
  NAND2_X1 U3384 ( .A1(n4179), .A2(n3539), .ZN(n2610) );
  NAND2_X1 U3385 ( .A1(n4196), .A2(n2610), .ZN(n2612) );
  INV_X1 U3386 ( .A(n3539), .ZN(n4209) );
  NAND2_X1 U3387 ( .A1(n4224), .A2(n4209), .ZN(n2611) );
  NAND2_X1 U3388 ( .A1(n2612), .A2(n2611), .ZN(n4172) );
  INV_X1 U3389 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4574) );
  NAND2_X1 U3390 ( .A1(n2613), .A2(n4574), .ZN(n2614) );
  NAND2_X1 U3391 ( .A1(n2629), .A2(n2614), .ZN(n4191) );
  OR2_X1 U3392 ( .A1(n4191), .A2(n2680), .ZN(n2619) );
  INV_X1 U3393 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4323) );
  NAND2_X1 U3394 ( .A1(n2455), .A2(REG2_REG_20__SCAN_IN), .ZN(n2616) );
  NAND2_X1 U3395 ( .A1(n2470), .A2(REG0_REG_20__SCAN_IN), .ZN(n2615) );
  OAI211_X1 U3396 ( .C1(n4323), .C2(n2471), .A(n2616), .B(n2615), .ZN(n2617)
         );
  INV_X1 U3397 ( .A(n2617), .ZN(n2618) );
  INV_X1 U3398 ( .A(DATAI_20_), .ZN(n2620) );
  NOR2_X1 U3399 ( .A1(n4312), .A2(n4178), .ZN(n2621) );
  INV_X1 U3400 ( .A(n4312), .ZN(n3668) );
  INV_X1 U3401 ( .A(n4178), .ZN(n4188) );
  XNOR2_X1 U3402 ( .A(n2629), .B(REG3_REG_21__SCAN_IN), .ZN(n4163) );
  NAND2_X1 U3403 ( .A1(n4163), .A2(n2419), .ZN(n2626) );
  INV_X1 U3404 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4318) );
  NAND2_X1 U3405 ( .A1(n2470), .A2(REG0_REG_21__SCAN_IN), .ZN(n2623) );
  NAND2_X1 U3406 ( .A1(n2455), .A2(REG2_REG_21__SCAN_IN), .ZN(n2622) );
  OAI211_X1 U3407 ( .C1(n2471), .C2(n4318), .A(n2623), .B(n2622), .ZN(n2624)
         );
  INV_X1 U3408 ( .A(n2624), .ZN(n2625) );
  NAND2_X1 U3409 ( .A1(n3779), .A2(DATAI_21_), .ZN(n4167) );
  INV_X1 U3410 ( .A(n4167), .ZN(n4311) );
  AND2_X1 U3411 ( .A1(n4141), .A2(n4311), .ZN(n2628) );
  OR2_X1 U3412 ( .A1(n4141), .A2(n4311), .ZN(n2627) );
  INV_X1 U3413 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3669) );
  INV_X1 U3414 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3730) );
  OAI21_X1 U3415 ( .B1(n2629), .B2(n3669), .A(n3730), .ZN(n2630) );
  NAND2_X1 U3416 ( .A1(n2630), .A2(n2639), .ZN(n4151) );
  OR2_X1 U3417 ( .A1(n4151), .A2(n2680), .ZN(n2636) );
  INV_X1 U3418 ( .A(REG1_REG_22__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U3419 ( .A1(n2470), .A2(REG0_REG_22__SCAN_IN), .ZN(n2632) );
  NAND2_X1 U3420 ( .A1(n2455), .A2(REG2_REG_22__SCAN_IN), .ZN(n2631) );
  OAI211_X1 U3421 ( .C1(n2471), .C2(n2633), .A(n2632), .B(n2631), .ZN(n2634)
         );
  INV_X1 U3422 ( .A(n2634), .ZN(n2635) );
  INV_X1 U3423 ( .A(DATAI_22_), .ZN(n2637) );
  NOR2_X1 U3424 ( .A1(n3780), .A2(n2637), .ZN(n2638) );
  NAND2_X1 U3425 ( .A1(n4315), .A2(n2638), .ZN(n4125) );
  NAND2_X1 U3426 ( .A1(n4162), .A2(n4149), .ZN(n2704) );
  INV_X1 U3427 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4611) );
  NAND2_X1 U3428 ( .A1(n2639), .A2(n4611), .ZN(n2640) );
  NAND2_X1 U3429 ( .A1(n2649), .A2(n2640), .ZN(n4134) );
  OR2_X1 U3430 ( .A1(n4134), .A2(n2680), .ZN(n2645) );
  INV_X1 U3431 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4302) );
  NAND2_X1 U3432 ( .A1(n2455), .A2(REG2_REG_23__SCAN_IN), .ZN(n2642) );
  NAND2_X1 U3433 ( .A1(n2470), .A2(REG0_REG_23__SCAN_IN), .ZN(n2641) );
  OAI211_X1 U3434 ( .C1(n4302), .C2(n2471), .A(n2642), .B(n2641), .ZN(n2643)
         );
  INV_X1 U3435 ( .A(n2643), .ZN(n2644) );
  INV_X1 U3436 ( .A(DATAI_23_), .ZN(n2646) );
  NOR2_X1 U3437 ( .A1(n3780), .A2(n2646), .ZN(n3558) );
  NOR2_X1 U3438 ( .A1(n4292), .A2(n3558), .ZN(n2647) );
  INV_X1 U3439 ( .A(n4292), .ZN(n4112) );
  INV_X1 U3440 ( .A(n3558), .ZN(n4132) );
  INV_X1 U3441 ( .A(REG3_REG_24__SCAN_IN), .ZN(n2648) );
  NAND2_X1 U3442 ( .A1(n2649), .A2(n2648), .ZN(n2650) );
  NAND2_X1 U3443 ( .A1(n2651), .A2(n2650), .ZN(n4110) );
  OR2_X1 U3444 ( .A1(n4110), .A2(n2680), .ZN(n2656) );
  INV_X1 U3445 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4298) );
  NAND2_X1 U3446 ( .A1(n2455), .A2(REG2_REG_24__SCAN_IN), .ZN(n2653) );
  NAND2_X1 U3447 ( .A1(n2470), .A2(REG0_REG_24__SCAN_IN), .ZN(n2652) );
  OAI211_X1 U3448 ( .C1(n4298), .C2(n2471), .A(n2653), .B(n2652), .ZN(n2654)
         );
  INV_X1 U3449 ( .A(n2654), .ZN(n2655) );
  INV_X1 U3450 ( .A(DATAI_24_), .ZN(n4588) );
  INV_X1 U3451 ( .A(n4283), .ZN(n3653) );
  OAI21_X1 U3452 ( .B1(n4282), .B2(n3950), .A(n4086), .ZN(n2660) );
  INV_X1 U3453 ( .A(n4282), .ZN(n4091) );
  NAND2_X1 U3454 ( .A1(n2660), .A2(n2659), .ZN(n4064) );
  NAND2_X1 U3455 ( .A1(n2661), .A2(n3751), .ZN(n2662) );
  NAND2_X1 U3456 ( .A1(n4077), .A2(n2419), .ZN(n2668) );
  INV_X1 U3457 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4280) );
  NAND2_X1 U34580 ( .A1(n2455), .A2(REG2_REG_26__SCAN_IN), .ZN(n2665) );
  NAND2_X1 U34590 ( .A1(n2470), .A2(REG0_REG_26__SCAN_IN), .ZN(n2664) );
  OAI211_X1 U3460 ( .C1(n4280), .C2(n2471), .A(n2665), .B(n2664), .ZN(n2666)
         );
  INV_X1 U3461 ( .A(n2666), .ZN(n2667) );
  INV_X1 U3462 ( .A(DATAI_26_), .ZN(n4642) );
  NOR2_X1 U3463 ( .A1(n3780), .A2(n4642), .ZN(n3864) );
  NOR2_X1 U3464 ( .A1(n4064), .A2(n2219), .ZN(n2670) );
  INV_X1 U3465 ( .A(n4269), .ZN(n4057) );
  INV_X1 U3466 ( .A(n2673), .ZN(n2672) );
  NAND2_X1 U34670 ( .A1(n2672), .A2(REG3_REG_28__SCAN_IN), .ZN(n4026) );
  INV_X1 U3468 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3607) );
  NAND2_X1 U34690 ( .A1(n2673), .A2(n3607), .ZN(n2674) );
  NAND2_X1 U3470 ( .A1(n4026), .A2(n2674), .ZN(n4035) );
  OR2_X1 U34710 ( .A1(n4035), .A2(n2680), .ZN(n2679) );
  INV_X1 U3472 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3625) );
  NAND2_X1 U34730 ( .A1(n2455), .A2(REG2_REG_28__SCAN_IN), .ZN(n2676) );
  NAND2_X1 U3474 ( .A1(n2470), .A2(REG0_REG_28__SCAN_IN), .ZN(n2675) );
  OAI211_X1 U34750 ( .C1(n3625), .C2(n2471), .A(n2676), .B(n2675), .ZN(n2677)
         );
  INV_X1 U3476 ( .A(n2677), .ZN(n2678) );
  INV_X1 U34770 ( .A(DATAI_28_), .ZN(n4417) );
  NOR2_X1 U3478 ( .A1(n3780), .A2(n4417), .ZN(n3618) );
  NAND2_X1 U34790 ( .A1(n4273), .A2(n3618), .ZN(n3851) );
  INV_X1 U3480 ( .A(n3618), .ZN(n4037) );
  NAND2_X1 U34810 ( .A1(n4061), .A2(n4037), .ZN(n3783) );
  NAND2_X1 U3482 ( .A1(n3851), .A2(n3783), .ZN(n3614) );
  OR2_X1 U34830 ( .A1(n4026), .A2(n2680), .ZN(n2685) );
  NAND2_X1 U3484 ( .A1(n2455), .A2(REG2_REG_29__SCAN_IN), .ZN(n2682) );
  NAND2_X1 U34850 ( .A1(n2470), .A2(REG0_REG_29__SCAN_IN), .ZN(n2681) );
  OAI211_X1 U3486 ( .C1(n2750), .C2(n2471), .A(n2682), .B(n2681), .ZN(n2683)
         );
  INV_X1 U34870 ( .A(n2683), .ZN(n2684) );
  NAND2_X1 U3488 ( .A1(n2685), .A2(n2684), .ZN(n3949) );
  NAND2_X1 U34890 ( .A1(n3779), .A2(DATAI_29_), .ZN(n4024) );
  XNOR2_X1 U3490 ( .A(n3949), .B(n4024), .ZN(n3862) );
  XNOR2_X1 U34910 ( .A(n2871), .B(n4409), .ZN(n2690) );
  NAND2_X1 U3492 ( .A1(n2690), .A2(n4011), .ZN(n4185) );
  AND2_X1 U34930 ( .A1(n2691), .A2(n4227), .ZN(n3009) );
  INV_X1 U3494 ( .A(n3966), .ZN(n2927) );
  NAND2_X1 U34950 ( .A1(n2927), .A2(n3007), .ZN(n3799) );
  NAND2_X1 U3496 ( .A1(n2958), .A2(n3892), .ZN(n2957) );
  NAND2_X1 U34970 ( .A1(n2977), .A2(n2995), .ZN(n3809) );
  NAND2_X1 U3498 ( .A1(n4253), .A2(n3239), .ZN(n3806) );
  AND2_X1 U34990 ( .A1(n3809), .A2(n3806), .ZN(n3877) );
  AND2_X1 U3500 ( .A1(n2694), .A2(n3090), .ZN(n3032) );
  NAND2_X1 U35010 ( .A1(n3084), .A2(n3204), .ZN(n3823) );
  NAND2_X1 U3502 ( .A1(n3962), .A2(n3101), .ZN(n3812) );
  NOR2_X1 U35030 ( .A1(n3962), .A2(n3101), .ZN(n3798) );
  NAND2_X1 U3504 ( .A1(n3269), .A2(n3159), .ZN(n3819) );
  NAND2_X1 U35050 ( .A1(n3960), .A2(n3168), .ZN(n3822) );
  AND2_X1 U35060 ( .A1(n3959), .A2(n3268), .ZN(n3831) );
  NAND2_X1 U35070 ( .A1(n3310), .A2(n3263), .ZN(n3820) );
  NAND2_X1 U35080 ( .A1(n3958), .A2(n3309), .ZN(n3833) );
  NAND2_X1 U35090 ( .A1(n3226), .A2(n3833), .ZN(n2696) );
  NAND2_X1 U35100 ( .A1(n3388), .A2(n3302), .ZN(n3828) );
  NAND2_X1 U35110 ( .A1(n3956), .A2(n3438), .ZN(n3343) );
  NAND2_X1 U35120 ( .A1(n3955), .A2(n3486), .ZN(n3318) );
  INV_X1 U35130 ( .A(n3835), .ZN(n3795) );
  NAND2_X1 U35140 ( .A1(n3487), .A2(n3433), .ZN(n3344) );
  OR2_X1 U35150 ( .A1(n3795), .A2(n3344), .ZN(n2697) );
  NAND2_X1 U35160 ( .A1(n3640), .A2(n3326), .ZN(n3319) );
  NAND2_X1 U35170 ( .A1(n2698), .A2(n3794), .ZN(n3335) );
  NAND2_X1 U35180 ( .A1(n4350), .A2(n3512), .ZN(n3792) );
  NAND2_X1 U35190 ( .A1(n3953), .A2(n3767), .ZN(n3790) );
  NAND2_X1 U35200 ( .A1(n3792), .A2(n3790), .ZN(n3875) );
  NAND2_X1 U35210 ( .A1(n3368), .A2(n3790), .ZN(n3475) );
  NAND2_X1 U35220 ( .A1(n3475), .A2(n3881), .ZN(n3474) );
  AND2_X1 U35230 ( .A1(n4347), .A2(n3699), .ZN(n3454) );
  NAND2_X1 U35240 ( .A1(n4179), .A2(n4209), .ZN(n3870) );
  NAND2_X1 U35250 ( .A1(n3870), .A2(n4199), .ZN(n3785) );
  NAND2_X1 U35260 ( .A1(n4312), .A2(n4188), .ZN(n3787) );
  OR2_X1 U35270 ( .A1(n4347), .A2(n3699), .ZN(n4197) );
  AND2_X1 U35280 ( .A1(n4198), .A2(n4197), .ZN(n2701) );
  NAND2_X1 U35290 ( .A1(n4224), .A2(n3539), .ZN(n3871) );
  OAI21_X1 U35300 ( .B1(n3785), .B2(n2701), .A(n3871), .ZN(n4173) );
  NOR2_X1 U35310 ( .A1(n4312), .A2(n4188), .ZN(n2702) );
  OR2_X1 U35320 ( .A1(n4173), .A2(n2702), .ZN(n2703) );
  NAND2_X1 U35330 ( .A1(n2703), .A2(n3787), .ZN(n3915) );
  OR2_X1 U35340 ( .A1(n4141), .A2(n4167), .ZN(n3867) );
  AND2_X1 U35350 ( .A1(n4125), .A2(n3867), .ZN(n3916) );
  INV_X1 U35360 ( .A(n3916), .ZN(n2706) );
  NAND2_X1 U35370 ( .A1(n4292), .A2(n4132), .ZN(n3868) );
  NAND2_X1 U35380 ( .A1(n3868), .A2(n2704), .ZN(n3845) );
  AND2_X1 U35390 ( .A1(n4141), .A2(n4167), .ZN(n4122) );
  AND2_X1 U35400 ( .A1(n4125), .A2(n4122), .ZN(n2705) );
  NOR2_X1 U35410 ( .A1(n3845), .A2(n2705), .ZN(n3917) );
  OR2_X1 U35420 ( .A1(n4292), .A2(n4132), .ZN(n3869) );
  NOR2_X1 U35430 ( .A1(n4283), .A2(n4107), .ZN(n3866) );
  NAND2_X1 U35440 ( .A1(n4286), .A2(n3864), .ZN(n2708) );
  NAND2_X1 U35450 ( .A1(n4295), .A2(n4282), .ZN(n4065) );
  NAND2_X1 U35460 ( .A1(n2708), .A2(n4065), .ZN(n3923) );
  NAND2_X1 U35470 ( .A1(n3950), .A2(n4091), .ZN(n3905) );
  NAND2_X1 U35480 ( .A1(n4283), .A2(n4107), .ZN(n4082) );
  NAND2_X1 U35490 ( .A1(n3905), .A2(n4082), .ZN(n4066) );
  AND2_X1 U35500 ( .A1(n4270), .A2(n4076), .ZN(n3926) );
  AOI21_X1 U35510 ( .B1(n2710), .B2(n4066), .A(n3926), .ZN(n3848) );
  XNOR2_X1 U35520 ( .A(n4072), .B(n4269), .ZN(n4051) );
  NAND2_X1 U35530 ( .A1(n4049), .A2(n4051), .ZN(n4048) );
  NAND2_X1 U35540 ( .A1(n3849), .A2(n4269), .ZN(n3850) );
  NAND2_X1 U35550 ( .A1(n4048), .A2(n3850), .ZN(n3616) );
  INV_X1 U35560 ( .A(n3851), .ZN(n2711) );
  XNOR2_X1 U35570 ( .A(n2712), .B(n3862), .ZN(n2716) );
  INV_X1 U35580 ( .A(n2691), .ZN(n4410) );
  NAND2_X1 U35590 ( .A1(n4410), .A2(n3937), .ZN(n2714) );
  NAND2_X1 U35600 ( .A1(n4227), .A2(n4409), .ZN(n2713) );
  NAND2_X1 U35610 ( .A1(n2716), .A2(n2715), .ZN(n2724) );
  NAND2_X1 U35620 ( .A1(n2455), .A2(REG2_REG_30__SCAN_IN), .ZN(n2720) );
  NAND2_X1 U35630 ( .A1(n2470), .A2(REG0_REG_30__SCAN_IN), .ZN(n2719) );
  INV_X1 U35640 ( .A(REG1_REG_30__SCAN_IN), .ZN(n2717) );
  OR2_X1 U35650 ( .A1(n2471), .A2(n2717), .ZN(n2718) );
  AND3_X1 U35660 ( .A1(n2720), .A2(n2719), .A3(n2718), .ZN(n3852) );
  INV_X1 U35670 ( .A(n3852), .ZN(n2722) );
  NAND2_X1 U35680 ( .A1(n4424), .A2(B_REG_SCAN_IN), .ZN(n2721) );
  NAND2_X1 U35690 ( .A1(n2906), .A2(n2841), .ZN(n4349) );
  NAND2_X1 U35700 ( .A1(n4410), .A2(n3006), .ZN(n4203) );
  OAI22_X1 U35710 ( .A1(n4273), .A2(n4349), .B1(n4024), .B2(n4203), .ZN(n2726)
         );
  INV_X1 U35720 ( .A(n2726), .ZN(n2727) );
  NAND2_X1 U35730 ( .A1(n2691), .A2(n4011), .ZN(n2840) );
  NAND2_X1 U35740 ( .A1(n2840), .A2(n2841), .ZN(n2845) );
  OAI211_X1 U35750 ( .C1(n4530), .C2(n3937), .A(n2864), .B(n2845), .ZN(n2728)
         );
  INV_X1 U35760 ( .A(n2728), .ZN(n2745) );
  INV_X1 U35770 ( .A(n2788), .ZN(n2733) );
  NAND2_X1 U35780 ( .A1(n2733), .A2(B_REG_SCAN_IN), .ZN(n2730) );
  MUX2_X1 U35790 ( .A(n2730), .B(B_REG_SCAN_IN), .S(n2729), .Z(n2731) );
  INV_X1 U35800 ( .A(D_REG_1__SCAN_IN), .ZN(n2732) );
  NAND2_X1 U35810 ( .A1(n2766), .A2(n2732), .ZN(n2837) );
  INV_X1 U3582 ( .A(n4408), .ZN(n2746) );
  NAND2_X1 U3583 ( .A1(n2733), .A2(n2746), .ZN(n2799) );
  NAND2_X1 U3584 ( .A1(n2837), .A2(n2799), .ZN(n2744) );
  NOR4_X1 U3585 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2737) );
  NOR4_X1 U3586 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2736) );
  NOR4_X1 U3587 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2735) );
  NOR4_X1 U3588 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2734) );
  NAND4_X1 U3589 ( .A1(n2737), .A2(n2736), .A3(n2735), .A4(n2734), .ZN(n2743)
         );
  NOR2_X1 U3590 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_3__SCAN_IN), .ZN(n2741) );
  NOR4_X1 U3591 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2740) );
  NOR4_X1 U3592 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2739) );
  NOR4_X1 U3593 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2738) );
  NAND4_X1 U3594 ( .A1(n2741), .A2(n2740), .A3(n2739), .A4(n2738), .ZN(n2742)
         );
  OAI21_X1 U3595 ( .B1(n2743), .B2(n2742), .A(n2766), .ZN(n2765) );
  INV_X1 U3596 ( .A(D_REG_0__SCAN_IN), .ZN(n2798) );
  NAND2_X1 U3597 ( .A1(n2766), .A2(n2798), .ZN(n2749) );
  INV_X1 U3598 ( .A(n2729), .ZN(n2747) );
  NAND2_X1 U3599 ( .A1(n2747), .A2(n2746), .ZN(n2748) );
  MUX2_X1 U3600 ( .A(n2750), .B(n2755), .S(n4552), .Z(n2753) );
  INV_X1 U3601 ( .A(n3007), .ZN(n3005) );
  NAND2_X1 U3602 ( .A1(n2876), .A2(n3005), .ZN(n2996) );
  NOR2_X2 U3603 ( .A1(n3038), .A2(n3204), .ZN(n3072) );
  NAND2_X1 U3604 ( .A1(n2753), .A2(n2752), .ZN(U3547) );
  INV_X1 U3605 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2756) );
  MUX2_X1 U3606 ( .A(n2756), .B(n2755), .S(n4546), .Z(n2758) );
  NAND2_X1 U3607 ( .A1(n2758), .A2(n2757), .ZN(U3515) );
  INV_X1 U3608 ( .A(n4522), .ZN(n2796) );
  NOR2_X1 U3609 ( .A1(n2858), .A2(n2796), .ZN(U4043) );
  INV_X1 U3610 ( .A(n2759), .ZN(n2760) );
  AOI21_X1 U3611 ( .B1(n2763), .B2(n3799), .A(n2760), .ZN(n2764) );
  OAI21_X1 U3612 ( .B1(n2763), .B2(n2762), .A(n2761), .ZN(n2894) );
  OAI22_X1 U3613 ( .A1(n2764), .A2(n4206), .B1(n4185), .B2(n2894), .ZN(n2896)
         );
  AND2_X1 U3614 ( .A1(n2765), .A2(n2799), .ZN(n2839) );
  INV_X1 U3615 ( .A(n2766), .ZN(n2767) );
  NAND2_X2 U3616 ( .A1(n2767), .A2(n2864), .ZN(n4521) );
  NAND2_X1 U3617 ( .A1(n2864), .A2(D_REG_1__SCAN_IN), .ZN(n2768) );
  NAND2_X1 U3618 ( .A1(n4521), .A2(n2768), .ZN(n2769) );
  NAND4_X1 U3619 ( .A1(n2770), .A2(n2839), .A3(n2845), .A4(n2769), .ZN(n2773)
         );
  AND2_X1 U3620 ( .A1(n2864), .A2(n2771), .ZN(n2772) );
  MUX2_X1 U3621 ( .A(REG2_REG_1__SCAN_IN), .B(n2896), .S(n4511), .Z(n2780) );
  INV_X1 U3622 ( .A(n4248), .ZN(n4111) );
  NAND2_X1 U3623 ( .A1(n4215), .A2(n4346), .ZN(n4113) );
  OAI22_X1 U3624 ( .A1(n4111), .A2(n2927), .B1(n2978), .B2(n4113), .ZN(n2779)
         );
  OR2_X1 U3625 ( .A1(n2871), .A2(n4011), .ZN(n3119) );
  INV_X1 U3626 ( .A(n3119), .ZN(n2774) );
  NAND2_X1 U3627 ( .A1(n4511), .A2(n2774), .ZN(n4246) );
  INV_X1 U3628 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2932) );
  OAI22_X1 U3629 ( .A1(n2894), .A2(n4246), .B1(n2932), .B2(n4508), .ZN(n2778)
         );
  NAND2_X1 U3630 ( .A1(n4215), .A2(n4345), .ZN(n4166) );
  AND2_X1 U3631 ( .A1(n4352), .A2(n4011), .ZN(n2775) );
  NAND2_X1 U3632 ( .A1(n2929), .A2(n3007), .ZN(n2776) );
  NAND2_X1 U3633 ( .A1(n2996), .A2(n2776), .ZN(n2901) );
  OAI22_X1 U3634 ( .A1(n2876), .A2(n4166), .B1(n4213), .B2(n2901), .ZN(n2777)
         );
  OR4_X1 U3635 ( .A1(n2780), .A2(n2779), .A3(n2778), .A4(n2777), .ZN(U3289) );
  INV_X2 U3636 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3637 ( .A(DATAI_13_), .ZN(n4587) );
  NAND2_X1 U3638 ( .A1(n2781), .A2(STATE_REG_SCAN_IN), .ZN(n2782) );
  OAI21_X1 U3639 ( .B1(STATE_REG_SCAN_IN), .B2(n4587), .A(n2782), .ZN(U3339)
         );
  INV_X1 U3640 ( .A(DATAI_21_), .ZN(n4669) );
  NAND2_X1 U3641 ( .A1(n3937), .A2(STATE_REG_SCAN_IN), .ZN(n2783) );
  OAI21_X1 U3642 ( .B1(STATE_REG_SCAN_IN), .B2(n4669), .A(n2783), .ZN(U3331)
         );
  INV_X1 U3643 ( .A(DATAI_17_), .ZN(n4680) );
  NAND2_X1 U3644 ( .A1(n2784), .A2(STATE_REG_SCAN_IN), .ZN(n2785) );
  OAI21_X1 U3645 ( .B1(STATE_REG_SCAN_IN), .B2(n4680), .A(n2785), .ZN(U3335)
         );
  INV_X1 U3646 ( .A(DATAI_7_), .ZN(n2786) );
  MUX2_X1 U3647 ( .A(n2786), .B(n2829), .S(STATE_REG_SCAN_IN), .Z(n2787) );
  INV_X1 U3648 ( .A(n2787), .ZN(U3345) );
  NAND2_X1 U3649 ( .A1(n2788), .A2(STATE_REG_SCAN_IN), .ZN(n2789) );
  OAI21_X1 U3650 ( .B1(STATE_REG_SCAN_IN), .B2(n2408), .A(n2789), .ZN(U3327)
         );
  NAND2_X1 U3651 ( .A1(n4424), .A2(STATE_REG_SCAN_IN), .ZN(n2790) );
  OAI21_X1 U3652 ( .B1(STATE_REG_SCAN_IN), .B2(n2390), .A(n2790), .ZN(U3325)
         );
  INV_X1 U3653 ( .A(n2791), .ZN(n4439) );
  INV_X1 U3654 ( .A(DATAI_9_), .ZN(n2792) );
  MUX2_X1 U3655 ( .A(n4439), .B(n2792), .S(U3149), .Z(n2793) );
  INV_X1 U3656 ( .A(n2793), .ZN(U3343) );
  INV_X1 U3657 ( .A(DATAI_19_), .ZN(n2794) );
  MUX2_X1 U3658 ( .A(n4011), .B(n2794), .S(U3149), .Z(n2795) );
  INV_X1 U3659 ( .A(n2795), .ZN(U3333) );
  NOR3_X1 U3660 ( .A1(n2796), .A2(n2729), .A3(n4408), .ZN(n2797) );
  AOI21_X1 U3661 ( .B1(n4521), .B2(n2798), .A(n2797), .ZN(U3458) );
  INV_X1 U3662 ( .A(n2799), .ZN(n2800) );
  AOI22_X1 U3663 ( .A1(n4521), .A2(n2732), .B1(n2800), .B2(n4522), .ZN(U3459)
         );
  NAND2_X1 U3664 ( .A1(n3965), .A2(DATAO_REG_30__SCAN_IN), .ZN(n2801) );
  OAI21_X1 U3665 ( .B1(n3852), .B2(n3965), .A(n2801), .ZN(U3580) );
  NOR2_X1 U3666 ( .A1(n4501), .A2(n3951), .ZN(U3148) );
  AOI211_X1 U3667 ( .C1(n2804), .C2(n2803), .A(n4495), .B(n2802), .ZN(n2808)
         );
  INV_X1 U3668 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4656) );
  NOR2_X1 U3669 ( .A1(STATE_REG_SCAN_IN), .A2(n4656), .ZN(n3092) );
  AOI21_X1 U3670 ( .B1(n4501), .B2(ADDR_REG_5__SCAN_IN), .A(n3092), .ZN(n2805)
         );
  OAI21_X1 U3671 ( .B1(n4507), .B2(n2806), .A(n2805), .ZN(n2807) );
  NOR2_X1 U3672 ( .A1(n2808), .A2(n2807), .ZN(n2813) );
  OAI211_X1 U3673 ( .C1(n2811), .C2(n2810), .A(n4502), .B(n2809), .ZN(n2812)
         );
  NAND2_X1 U3674 ( .A1(n2813), .A2(n2812), .ZN(U3245) );
  XOR2_X1 U3675 ( .A(REG2_REG_6__SCAN_IN), .B(n2814), .Z(n2823) );
  INV_X1 U3676 ( .A(n4502), .ZN(n2816) );
  AOI211_X1 U3677 ( .C1(n2818), .C2(n2817), .A(n2816), .B(n2815), .ZN(n2822)
         );
  INV_X1 U3678 ( .A(n4412), .ZN(n2820) );
  AND2_X1 U3679 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3103) );
  AOI21_X1 U3680 ( .B1(n4501), .B2(ADDR_REG_6__SCAN_IN), .A(n3103), .ZN(n2819)
         );
  OAI21_X1 U3681 ( .B1(n4507), .B2(n2820), .A(n2819), .ZN(n2821) );
  AOI211_X1 U3682 ( .C1(n2823), .C2(n4466), .A(n2822), .B(n2821), .ZN(n2824)
         );
  INV_X1 U3683 ( .A(n2824), .ZN(U3246) );
  MUX2_X1 U3684 ( .A(REG1_REG_7__SCAN_IN), .B(n4550), .S(n2825), .Z(n2826) );
  XNOR2_X1 U3685 ( .A(n2827), .B(n2826), .ZN(n2835) );
  NOR2_X1 U3686 ( .A1(STATE_REG_SCAN_IN), .A2(n2463), .ZN(n3180) );
  AOI21_X1 U3687 ( .B1(n4501), .B2(ADDR_REG_7__SCAN_IN), .A(n3180), .ZN(n2828)
         );
  OAI21_X1 U3688 ( .B1(n4507), .B2(n2829), .A(n2828), .ZN(n2834) );
  AOI211_X1 U3689 ( .C1(n2832), .C2(n2831), .A(n4495), .B(n2830), .ZN(n2833)
         );
  AOI211_X1 U3690 ( .C1(n4502), .C2(n2835), .A(n2834), .B(n2833), .ZN(n2836)
         );
  INV_X1 U3691 ( .A(n2836), .ZN(U3247) );
  NAND3_X1 U3692 ( .A1(n2839), .A2(n2838), .A3(n2837), .ZN(n2888) );
  NAND2_X1 U3693 ( .A1(n2840), .A2(n3006), .ZN(n2843) );
  INV_X1 U3694 ( .A(n2841), .ZN(n2842) );
  NAND2_X1 U3695 ( .A1(n2843), .A2(n2842), .ZN(n2863) );
  NAND2_X1 U3696 ( .A1(n2863), .A2(n4203), .ZN(n2844) );
  NAND2_X1 U3697 ( .A1(n2888), .A2(n2844), .ZN(n2846) );
  NAND2_X1 U3698 ( .A1(n2846), .A2(n2845), .ZN(n2980) );
  INV_X1 U3699 ( .A(n2980), .ZN(n2850) );
  INV_X1 U3700 ( .A(n2870), .ZN(n2848) );
  NAND2_X1 U3701 ( .A1(n2848), .A2(n4522), .ZN(n2849) );
  NAND2_X1 U3702 ( .A1(n2888), .A2(n3944), .ZN(n2981) );
  NAND3_X1 U3703 ( .A1(n2850), .A2(n2864), .A3(n2981), .ZN(n2891) );
  INV_X1 U3704 ( .A(n2891), .ZN(n2933) );
  AND2_X1 U3705 ( .A1(n2864), .A2(n4345), .ZN(n2851) );
  NAND2_X1 U3706 ( .A1(n2867), .A2(n2851), .ZN(n2852) );
  AND2_X2 U3707 ( .A1(n2852), .A2(n4508), .ZN(n3768) );
  INV_X1 U3708 ( .A(n3768), .ZN(n3044) );
  NAND2_X1 U3709 ( .A1(n3966), .A2(n2043), .ZN(n2854) );
  NAND2_X1 U3710 ( .A1(n3007), .A2(n2044), .ZN(n2853) );
  INV_X1 U3711 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2855) );
  NAND2_X1 U3712 ( .A1(n2057), .A2(n2216), .ZN(n2862) );
  NAND2_X1 U3713 ( .A1(n3966), .A2(n2857), .ZN(n2860) );
  INV_X1 U3714 ( .A(n2858), .ZN(n2979) );
  AOI22_X1 U3715 ( .A1(n2878), .A2(n3007), .B1(n2979), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2859) );
  NAND2_X1 U3716 ( .A1(n2860), .A2(n2859), .ZN(n2861) );
  OAI21_X1 U3717 ( .B1(n2862), .B2(n2861), .A(n2874), .ZN(n2907) );
  INV_X1 U3718 ( .A(n2863), .ZN(n2865) );
  AND2_X1 U3719 ( .A1(n2865), .A2(n2864), .ZN(n2866) );
  NAND3_X1 U3720 ( .A1(n2867), .A2(n3944), .A3(n4418), .ZN(n3755) );
  OAI22_X1 U3721 ( .A1(n2907), .A2(n3759), .B1(n3755), .B2(n2880), .ZN(n2868)
         );
  AOI21_X1 U3722 ( .B1(n3007), .B2(n3044), .A(n2868), .ZN(n2869) );
  OAI21_X1 U3723 ( .B1(n2933), .B2(n3010), .A(n2869), .ZN(U3229) );
  OAI22_X1 U3724 ( .A1(n2978), .A2(n3049), .B1(n3599), .B2(n2962), .ZN(n2872)
         );
  XNOR2_X1 U3725 ( .A(n2872), .B(n3602), .ZN(n2970) );
  OAI22_X1 U3726 ( .A1(n2978), .A2(n3601), .B1(n3049), .B2(n2962), .ZN(n2969)
         );
  XNOR2_X1 U3727 ( .A(n2970), .B(n2969), .ZN(n2886) );
  NAND2_X1 U3728 ( .A1(n2874), .A2(n2873), .ZN(n2926) );
  NAND2_X1 U3729 ( .A1(n2929), .A2(n2043), .ZN(n2879) );
  OAI21_X1 U3730 ( .B1(n3601), .B2(n2880), .A(n2879), .ZN(n2881) );
  NAND2_X1 U3731 ( .A1(n2926), .A2(n2924), .ZN(n2925) );
  NAND2_X1 U3732 ( .A1(n2925), .A2(n2884), .ZN(n2885) );
  NOR2_X1 U3733 ( .A1(n2885), .A2(n2886), .ZN(n2971) );
  AOI21_X1 U3734 ( .B1(n2886), .B2(n2885), .A(n2971), .ZN(n2893) );
  INV_X1 U3735 ( .A(n3944), .ZN(n2887) );
  NOR3_X2 U3736 ( .A1(n2888), .A2(n2887), .A3(n4418), .ZN(n3753) );
  AOI22_X1 U3737 ( .A1(n3753), .A2(n4247), .B1(n3772), .B2(n4253), .ZN(n2889)
         );
  OAI21_X1 U3738 ( .B1(n3768), .B2(n2962), .A(n2889), .ZN(n2890) );
  AOI21_X1 U3739 ( .B1(REG3_REG_2__SCAN_IN), .B2(n2891), .A(n2890), .ZN(n2892)
         );
  OAI21_X1 U3740 ( .B1(n2893), .B2(n3759), .A(n2892), .ZN(U3234) );
  INV_X1 U3741 ( .A(n2894), .ZN(n2898) );
  AOI22_X1 U3742 ( .A1(n3964), .A2(n4346), .B1(n4345), .B2(n2929), .ZN(n2895)
         );
  OAI21_X1 U3743 ( .B1(n2927), .B2(n4349), .A(n2895), .ZN(n2897) );
  AOI211_X1 U3744 ( .C1(n4536), .C2(n2898), .A(n2897), .B(n2896), .ZN(n2904)
         );
  OAI22_X1 U3745 ( .A1(n4343), .A2(n2901), .B1(n4552), .B2(n2416), .ZN(n2899)
         );
  INV_X1 U3746 ( .A(n2899), .ZN(n2900) );
  OAI21_X1 U3747 ( .B1(n2904), .B2(n4549), .A(n2900), .ZN(U3519) );
  OAI22_X1 U3748 ( .A1(n4404), .A2(n2901), .B1(n4546), .B2(n2418), .ZN(n2902)
         );
  INV_X1 U3749 ( .A(n2902), .ZN(n2903) );
  OAI21_X1 U3750 ( .B1(n2904), .B2(n4544), .A(n2903), .ZN(U3469) );
  INV_X1 U3751 ( .A(IR_REG_0__SCAN_IN), .ZN(n4429) );
  NAND2_X1 U3752 ( .A1(n4424), .A2(n3011), .ZN(n2905) );
  NAND2_X1 U3753 ( .A1(n2906), .A2(n2905), .ZN(n4425) );
  NOR2_X1 U3754 ( .A1(n2907), .A2(n4424), .ZN(n2908) );
  AOI211_X1 U3755 ( .C1(n4424), .C2(n3970), .A(n4418), .B(n2908), .ZN(n2909)
         );
  AOI211_X1 U3756 ( .C1(n4429), .C2(n4425), .A(n3965), .B(n2909), .ZN(n2941)
         );
  AOI211_X1 U3757 ( .C1(n2912), .C2(n2911), .A(n2910), .B(n4495), .ZN(n2923)
         );
  OAI211_X1 U3758 ( .C1(n2915), .C2(n2914), .A(n4502), .B(n2913), .ZN(n2916)
         );
  INV_X1 U3759 ( .A(n2916), .ZN(n2922) );
  INV_X1 U3760 ( .A(n4415), .ZN(n2920) );
  NOR2_X1 U3761 ( .A1(n2917), .A2(STATE_REG_SCAN_IN), .ZN(n2918) );
  AOI21_X1 U3762 ( .B1(n4501), .B2(ADDR_REG_2__SCAN_IN), .A(n2918), .ZN(n2919)
         );
  OAI21_X1 U3763 ( .B1(n4507), .B2(n2920), .A(n2919), .ZN(n2921) );
  OR4_X1 U3764 ( .A1(n2941), .A2(n2923), .A3(n2922), .A4(n2921), .ZN(U3242) );
  OAI211_X1 U3765 ( .C1(n2924), .C2(n2926), .A(n2925), .B(n3764), .ZN(n2931)
         );
  OAI22_X1 U3766 ( .A1(n3770), .A2(n2927), .B1(n2978), .B2(n3755), .ZN(n2928)
         );
  AOI21_X1 U3767 ( .B1(n2929), .B2(n3044), .A(n2928), .ZN(n2930) );
  OAI211_X1 U3768 ( .C1(n2933), .C2(n2932), .A(n2931), .B(n2930), .ZN(U3219)
         );
  XOR2_X1 U3769 ( .A(REG2_REG_4__SCAN_IN), .B(n2934), .Z(n2943) );
  OAI211_X1 U3770 ( .C1(REG1_REG_4__SCAN_IN), .C2(n2936), .A(n4502), .B(n2935), 
        .ZN(n2939) );
  NAND2_X1 U3771 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3045) );
  INV_X1 U3772 ( .A(n3045), .ZN(n2937) );
  AOI21_X1 U3773 ( .B1(n4501), .B2(ADDR_REG_4__SCAN_IN), .A(n2937), .ZN(n2938)
         );
  OAI211_X1 U3774 ( .C1(n4507), .C2(n2940), .A(n2939), .B(n2938), .ZN(n2942)
         );
  AOI211_X1 U3775 ( .C1(n4466), .C2(n2943), .A(n2942), .B(n2941), .ZN(n2944)
         );
  INV_X1 U3776 ( .A(n2944), .ZN(U3244) );
  XNOR2_X1 U3777 ( .A(n2945), .B(REG1_REG_8__SCAN_IN), .ZN(n2946) );
  NAND2_X1 U3778 ( .A1(n2946), .A2(n4502), .ZN(n2952) );
  XNOR2_X1 U3779 ( .A(REG2_REG_8__SCAN_IN), .B(n2947), .ZN(n2948) );
  NAND2_X1 U3780 ( .A1(n4466), .A2(n2948), .ZN(n2949) );
  NAND2_X1 U3781 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3167) );
  NAND2_X1 U3782 ( .A1(n2949), .A2(n3167), .ZN(n2950) );
  AOI21_X1 U3783 ( .B1(n4501), .B2(ADDR_REG_8__SCAN_IN), .A(n2950), .ZN(n2951)
         );
  OAI211_X1 U3784 ( .C1(n4507), .C2(n4411), .A(n2952), .B(n2951), .ZN(U3248)
         );
  INV_X1 U3785 ( .A(n2953), .ZN(n2955) );
  INV_X1 U3786 ( .A(n3892), .ZN(n2954) );
  OAI21_X1 U3787 ( .B1(n2955), .B2(n2954), .A(n3016), .ZN(n4249) );
  AOI22_X1 U3788 ( .A1(n4253), .A2(n4346), .B1(n4251), .B2(n4345), .ZN(n2956)
         );
  OAI21_X1 U3789 ( .B1(n2880), .B2(n4349), .A(n2956), .ZN(n2961) );
  INV_X1 U3790 ( .A(n4185), .ZN(n3134) );
  OAI21_X1 U3791 ( .B1(n3892), .B2(n2958), .A(n2957), .ZN(n2959) );
  AOI22_X1 U3792 ( .A1(n4249), .A2(n3134), .B1(n2715), .B2(n2959), .ZN(n4244)
         );
  INV_X1 U3793 ( .A(n4244), .ZN(n2960) );
  AOI211_X1 U3794 ( .C1(n4536), .C2(n4249), .A(n2961), .B(n2960), .ZN(n2968)
         );
  XNOR2_X1 U3795 ( .A(n2996), .B(n2962), .ZN(n4255) );
  AOI22_X1 U3796 ( .A1(n3362), .A2(n4255), .B1(REG0_REG_2__SCAN_IN), .B2(n4544), .ZN(n2963) );
  OAI21_X1 U3797 ( .B1(n2968), .B2(n4544), .A(n2963), .ZN(U3471) );
  INV_X1 U3798 ( .A(n4255), .ZN(n2965) );
  OAI22_X1 U3799 ( .A1(n4343), .A2(n2965), .B1(n4552), .B2(n2964), .ZN(n2966)
         );
  INV_X1 U3800 ( .A(n2966), .ZN(n2967) );
  OAI21_X1 U3801 ( .B1(n2968), .B2(n4549), .A(n2967), .ZN(U3520) );
  INV_X1 U3802 ( .A(n2969), .ZN(n2973) );
  INV_X1 U3803 ( .A(n2970), .ZN(n2972) );
  AOI21_X1 U3804 ( .B1(n2973), .B2(n2972), .A(n2971), .ZN(n3056) );
  NAND2_X1 U3805 ( .A1(n4253), .A2(n2878), .ZN(n2975) );
  NAND2_X1 U3806 ( .A1(n2995), .A2(n2044), .ZN(n2974) );
  NAND2_X1 U3807 ( .A1(n2975), .A2(n2974), .ZN(n2976) );
  XNOR2_X1 U3808 ( .A(n2976), .B(n3602), .ZN(n3054) );
  OAI22_X1 U3809 ( .A1(n2977), .A2(n3601), .B1(n3600), .B2(n3239), .ZN(n3053)
         );
  XNOR2_X1 U3810 ( .A(n3054), .B(n3053), .ZN(n3055) );
  XOR2_X1 U3811 ( .A(n3056), .B(n3055), .Z(n2987) );
  OAI22_X1 U3812 ( .A1(n3770), .A2(n2978), .B1(n3240), .B2(n3755), .ZN(n2985)
         );
  OAI21_X1 U3813 ( .B1(n2980), .B2(n2979), .A(STATE_REG_SCAN_IN), .ZN(n2983)
         );
  AND2_X1 U3814 ( .A1(n2981), .A2(n3947), .ZN(n2982) );
  MUX2_X1 U3815 ( .A(n3757), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n2984) );
  AOI211_X1 U3816 ( .C1(n2995), .C2(n3044), .A(n2985), .B(n2984), .ZN(n2986)
         );
  OAI21_X1 U3817 ( .B1(n2987), .B2(n3759), .A(n2986), .ZN(U3215) );
  NAND2_X1 U3818 ( .A1(n3016), .A2(n2988), .ZN(n2989) );
  XOR2_X1 U3819 ( .A(n3877), .B(n2989), .Z(n3244) );
  OAI22_X1 U3820 ( .A1(n3240), .A2(n4337), .B1(n4203), .B2(n3239), .ZN(n2994)
         );
  OAI21_X1 U3821 ( .B1(n3877), .B2(n2991), .A(n2990), .ZN(n2992) );
  AOI22_X1 U3822 ( .A1(n2992), .A2(n2715), .B1(n4333), .B2(n3964), .ZN(n3247)
         );
  INV_X1 U3823 ( .A(n3247), .ZN(n2993) );
  AOI211_X1 U3824 ( .C1(n4340), .C2(n3244), .A(n2994), .B(n2993), .ZN(n3004)
         );
  OAI21_X1 U3825 ( .B1(n2996), .B2(n4251), .A(n2995), .ZN(n2997) );
  INV_X1 U3826 ( .A(n2997), .ZN(n2998) );
  NOR2_X1 U3827 ( .A1(n2998), .A2(n3026), .ZN(n3243) );
  AOI22_X1 U3828 ( .A1(n3362), .A2(n3243), .B1(REG0_REG_3__SCAN_IN), .B2(n4544), .ZN(n2999) );
  OAI21_X1 U3829 ( .B1(n3004), .B2(n4544), .A(n2999), .ZN(U3473) );
  INV_X1 U3830 ( .A(n3243), .ZN(n3001) );
  OAI22_X1 U3831 ( .A1(n4343), .A2(n3001), .B1(n4552), .B2(n3000), .ZN(n3002)
         );
  INV_X1 U3832 ( .A(n3002), .ZN(n3003) );
  OAI21_X1 U3833 ( .B1(n3004), .B2(n4549), .A(n3003), .ZN(U3521) );
  NAND2_X1 U3834 ( .A1(n3966), .A2(n3005), .ZN(n3801) );
  AND2_X1 U3835 ( .A1(n3799), .A2(n3801), .ZN(n4531) );
  NAND2_X1 U3836 ( .A1(n3007), .A2(n3006), .ZN(n4528) );
  AOI21_X1 U3837 ( .B1(n4206), .B2(n4185), .A(n4531), .ZN(n3008) );
  AOI21_X1 U3838 ( .B1(n4346), .B2(n4247), .A(n3008), .ZN(n4529) );
  OAI21_X1 U3839 ( .B1(n3009), .B2(n4528), .A(n4529), .ZN(n3013) );
  OAI22_X1 U3840 ( .A1(n4511), .A2(n3011), .B1(n3010), .B2(n4508), .ZN(n3012)
         );
  AOI21_X1 U3841 ( .B1(n3013), .B2(n4215), .A(n3012), .ZN(n3014) );
  OAI21_X1 U3842 ( .B1(n4531), .B2(n4246), .A(n3014), .ZN(U3290) );
  NAND2_X1 U3843 ( .A1(n3016), .A2(n3015), .ZN(n3018) );
  AND2_X1 U3844 ( .A1(n3018), .A2(n3017), .ZN(n3019) );
  NAND2_X1 U3845 ( .A1(n3019), .A2(n3893), .ZN(n3020) );
  INV_X1 U3846 ( .A(n4537), .ZN(n3030) );
  XOR2_X1 U3847 ( .A(n3893), .B(n3021), .Z(n3025) );
  AOI22_X1 U3848 ( .A1(n4253), .A2(n4333), .B1(n3050), .B2(n4345), .ZN(n3022)
         );
  OAI21_X1 U3849 ( .B1(n3084), .B2(n4337), .A(n3022), .ZN(n3023) );
  AOI21_X1 U3850 ( .B1(n4537), .B2(n3134), .A(n3023), .ZN(n3024) );
  OAI21_X1 U3851 ( .B1(n3025), .B2(n4206), .A(n3024), .ZN(n4534) );
  OAI211_X1 U3852 ( .C1(n3026), .C2(n3047), .A(n3038), .B(n4352), .ZN(n4533)
         );
  OAI22_X1 U3853 ( .A1(n4533), .A2(n4227), .B1(n4508), .B2(n3043), .ZN(n3027)
         );
  OAI21_X1 U3854 ( .B1(n4534), .B2(n3027), .A(n4215), .ZN(n3029) );
  NAND2_X1 U3855 ( .A1(n4520), .A2(REG2_REG_4__SCAN_IN), .ZN(n3028) );
  OAI211_X1 U3856 ( .C1(n3030), .C2(n4246), .A(n3029), .B(n3028), .ZN(U3286)
         );
  NAND2_X1 U3857 ( .A1(n3115), .A2(n3031), .ZN(n3033) );
  INV_X1 U3858 ( .A(n3032), .ZN(n3813) );
  AND2_X1 U3859 ( .A1(n3813), .A2(n3823), .ZN(n3890) );
  XNOR2_X1 U3860 ( .A(n3033), .B(n3890), .ZN(n3211) );
  XOR2_X1 U3861 ( .A(n3890), .B(n3034), .Z(n3035) );
  NAND2_X1 U3862 ( .A1(n3035), .A2(n2715), .ZN(n3213) );
  AOI22_X1 U3863 ( .A1(n3962), .A2(n4346), .B1(n4345), .B2(n3204), .ZN(n3036)
         );
  OAI211_X1 U3864 ( .C1(n3240), .C2(n4349), .A(n3213), .B(n3036), .ZN(n3037)
         );
  AOI21_X1 U3865 ( .B1(n3211), .B2(n4340), .A(n3037), .ZN(n3042) );
  INV_X1 U3866 ( .A(n4343), .ZN(n3279) );
  AND2_X1 U3867 ( .A1(n3038), .A2(n3204), .ZN(n3039) );
  NOR2_X1 U3868 ( .A1(n3072), .A2(n3039), .ZN(n3207) );
  AOI22_X1 U3869 ( .A1(n3279), .A2(n3207), .B1(REG1_REG_5__SCAN_IN), .B2(n4549), .ZN(n3040) );
  OAI21_X1 U3870 ( .B1(n3042), .B2(n4549), .A(n3040), .ZN(U3523) );
  AOI22_X1 U3871 ( .A1(n3362), .A2(n3207), .B1(REG0_REG_5__SCAN_IN), .B2(n4544), .ZN(n3041) );
  OAI21_X1 U3872 ( .B1(n3042), .B2(n4544), .A(n3041), .ZN(U3477) );
  INV_X1 U3873 ( .A(n3043), .ZN(n3061) );
  AOI22_X1 U3874 ( .A1(n3050), .A2(n3044), .B1(n3753), .B2(n4253), .ZN(n3046)
         );
  OAI211_X1 U3875 ( .C1(n3084), .C2(n3755), .A(n3046), .B(n3045), .ZN(n3060)
         );
  OAI22_X1 U3876 ( .A1(n3240), .A2(n3600), .B1(n3599), .B2(n3047), .ZN(n3048)
         );
  XNOR2_X1 U3877 ( .A(n3048), .B(n3602), .ZN(n3081) );
  OR2_X1 U3878 ( .A1(n3240), .A2(n3601), .ZN(n3052) );
  NAND2_X1 U3879 ( .A1(n3050), .A2(n2878), .ZN(n3051) );
  NAND2_X1 U3880 ( .A1(n3052), .A2(n3051), .ZN(n3082) );
  XNOR2_X1 U3881 ( .A(n3081), .B(n3082), .ZN(n3058) );
  OAI22_X1 U3882 ( .A1(n3056), .A2(n3055), .B1(n3054), .B2(n3053), .ZN(n3057)
         );
  AOI211_X1 U3883 ( .C1(n3058), .C2(n3057), .A(n3759), .B(n3080), .ZN(n3059)
         );
  AOI211_X1 U3884 ( .C1(n3061), .C2(n3757), .A(n3060), .B(n3059), .ZN(n3062)
         );
  INV_X1 U3885 ( .A(n3062), .ZN(U3227) );
  NAND2_X1 U3886 ( .A1(n3115), .A2(n3063), .ZN(n3065) );
  AND2_X1 U3887 ( .A1(n3065), .A2(n3064), .ZN(n3066) );
  INV_X1 U3888 ( .A(n3812), .ZN(n3824) );
  OR2_X1 U3889 ( .A1(n3824), .A2(n3798), .ZN(n3067) );
  INV_X1 U3890 ( .A(n3067), .ZN(n3878) );
  XNOR2_X1 U3891 ( .A(n3066), .B(n3878), .ZN(n3223) );
  XNOR2_X1 U3892 ( .A(n3068), .B(n3067), .ZN(n3225) );
  OAI22_X1 U3893 ( .A1(n3221), .A2(n4337), .B1(n3101), .B2(n4203), .ZN(n3069)
         );
  AOI21_X1 U3894 ( .B1(n4333), .B2(n2694), .A(n3069), .ZN(n3070) );
  OAI21_X1 U3895 ( .B1(n3225), .B2(n4206), .A(n3070), .ZN(n3071) );
  AOI21_X1 U3896 ( .B1(n3223), .B2(n4340), .A(n3071), .ZN(n3079) );
  INV_X1 U3897 ( .A(n3072), .ZN(n3074) );
  INV_X1 U3898 ( .A(n3108), .ZN(n3073) );
  AOI21_X1 U3899 ( .B1(n3218), .B2(n3074), .A(n3073), .ZN(n3217) );
  INV_X1 U3900 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3075) );
  NOR2_X1 U3901 ( .A1(n4546), .A2(n3075), .ZN(n3076) );
  AOI21_X1 U3902 ( .B1(n3217), .B2(n3362), .A(n3076), .ZN(n3077) );
  OAI21_X1 U3903 ( .B1(n3079), .B2(n4544), .A(n3077), .ZN(U3479) );
  AOI22_X1 U3904 ( .A1(n3217), .A2(n3279), .B1(n4549), .B2(REG1_REG_6__SCAN_IN), .ZN(n3078) );
  OAI21_X1 U3905 ( .B1(n3079), .B2(n4549), .A(n3078), .ZN(U3524) );
  OAI22_X1 U3906 ( .A1(n3084), .A2(n3600), .B1(n3599), .B2(n3090), .ZN(n3083)
         );
  XNOR2_X1 U3907 ( .A(n3083), .B(n3602), .ZN(n3096) );
  OR2_X1 U3908 ( .A1(n3084), .A2(n3601), .ZN(n3086) );
  NAND2_X1 U3909 ( .A1(n3204), .A2(n2878), .ZN(n3085) );
  NAND2_X1 U3910 ( .A1(n3086), .A2(n3085), .ZN(n3095) );
  XNOR2_X1 U3911 ( .A(n3096), .B(n3095), .ZN(n3087) );
  AOI211_X1 U3912 ( .C1(n3088), .C2(n3087), .A(n3759), .B(n3097), .ZN(n3089)
         );
  INV_X1 U3913 ( .A(n3089), .ZN(n3094) );
  OAI22_X1 U3914 ( .A1(n3770), .A2(n3240), .B1(n3768), .B2(n3090), .ZN(n3091)
         );
  AOI211_X1 U3915 ( .C1(n3772), .C2(n3962), .A(n3092), .B(n3091), .ZN(n3093)
         );
  OAI211_X1 U3916 ( .C1(n3776), .C2(n3205), .A(n3094), .B(n3093), .ZN(U3224)
         );
  OAI22_X1 U3917 ( .A1(n3178), .A2(n3600), .B1(n3599), .B2(n3101), .ZN(n3098)
         );
  XNOR2_X1 U3918 ( .A(n3098), .B(n3602), .ZN(n3145) );
  OAI22_X1 U3919 ( .A1(n3178), .A2(n3601), .B1(n3600), .B2(n3101), .ZN(n3144)
         );
  INV_X1 U3920 ( .A(n3144), .ZN(n3148) );
  XNOR2_X1 U3921 ( .A(n3145), .B(n3148), .ZN(n3099) );
  XNOR2_X1 U3922 ( .A(n3149), .B(n3099), .ZN(n3100) );
  NAND2_X1 U3923 ( .A1(n3100), .A2(n3764), .ZN(n3105) );
  OAI22_X1 U3924 ( .A1(n3770), .A2(n3084), .B1(n3768), .B2(n3101), .ZN(n3102)
         );
  AOI211_X1 U3925 ( .C1(n3772), .C2(n3961), .A(n3103), .B(n3102), .ZN(n3104)
         );
  OAI211_X1 U3926 ( .C1(n3776), .C2(n3214), .A(n3105), .B(n3104), .ZN(U3236)
         );
  INV_X1 U3927 ( .A(n3136), .ZN(n3106) );
  AOI211_X1 U3928 ( .C1(n3152), .C2(n3108), .A(n3107), .B(n3106), .ZN(n4541)
         );
  INV_X1 U3929 ( .A(n3117), .ZN(n3880) );
  XNOR2_X1 U3930 ( .A(n3109), .B(n3880), .ZN(n3112) );
  OAI22_X1 U3931 ( .A1(n3269), .A2(n4337), .B1(n4203), .B2(n3177), .ZN(n3110)
         );
  AOI21_X1 U3932 ( .B1(n4333), .B2(n3962), .A(n3110), .ZN(n3111) );
  OAI21_X1 U3933 ( .B1(n3112), .B2(n4206), .A(n3111), .ZN(n4540) );
  AOI21_X1 U3934 ( .B1(n4541), .B2(n4011), .A(n4540), .ZN(n3127) );
  INV_X1 U3935 ( .A(n4511), .ZN(n4419) );
  NAND2_X1 U3936 ( .A1(n3115), .A2(n3114), .ZN(n3122) );
  AND2_X1 U3937 ( .A1(n3122), .A2(n3116), .ZN(n3118) );
  NOR2_X1 U3938 ( .A1(n3118), .A2(n3117), .ZN(n4539) );
  NAND2_X1 U3939 ( .A1(n4185), .A2(n3119), .ZN(n3120) );
  NOR2_X1 U3940 ( .A1(n4539), .A2(n4239), .ZN(n3125) );
  NAND2_X1 U3941 ( .A1(n3122), .A2(n3121), .ZN(n4542) );
  OAI22_X1 U3942 ( .A1(n4511), .A2(n3123), .B1(n3183), .B2(n4508), .ZN(n3124)
         );
  AOI21_X1 U3943 ( .B1(n3125), .B2(n4542), .A(n3124), .ZN(n3126) );
  OAI21_X1 U3944 ( .B1(n3127), .B2(n4419), .A(n3126), .ZN(U3283) );
  AND2_X1 U3945 ( .A1(n3819), .A2(n3822), .ZN(n3876) );
  XNOR2_X1 U3946 ( .A(n3128), .B(n3876), .ZN(n4516) );
  INV_X1 U3947 ( .A(n4516), .ZN(n3135) );
  XNOR2_X1 U3948 ( .A(n3129), .B(n3876), .ZN(n3132) );
  OAI22_X1 U3949 ( .A1(n3221), .A2(n4349), .B1(n3168), .B2(n4203), .ZN(n3130)
         );
  AOI21_X1 U3950 ( .B1(n4346), .B2(n3959), .A(n3130), .ZN(n3131) );
  OAI21_X1 U3951 ( .B1(n3132), .B2(n4206), .A(n3131), .ZN(n3133) );
  AOI21_X1 U3952 ( .B1(n3134), .B2(n4516), .A(n3133), .ZN(n4519) );
  OAI21_X1 U3953 ( .B1(n4530), .B2(n3135), .A(n4519), .ZN(n3140) );
  NAND2_X1 U3954 ( .A1(n3140), .A2(n4552), .ZN(n3139) );
  AND2_X1 U3955 ( .A1(n3136), .A2(n3159), .ZN(n3137) );
  NOR2_X1 U3956 ( .A1(n3190), .A2(n3137), .ZN(n4513) );
  NAND2_X1 U3957 ( .A1(n4513), .A2(n3279), .ZN(n3138) );
  OAI211_X1 U3958 ( .C1(n4552), .C2(n2492), .A(n3139), .B(n3138), .ZN(U3526)
         );
  INV_X1 U3959 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3143) );
  NAND2_X1 U3960 ( .A1(n3140), .A2(n4546), .ZN(n3142) );
  NAND2_X1 U3961 ( .A1(n4513), .A2(n3362), .ZN(n3141) );
  OAI211_X1 U3962 ( .C1(n4546), .C2(n3143), .A(n3142), .B(n3141), .ZN(U3483)
         );
  INV_X1 U3963 ( .A(n3145), .ZN(n3146) );
  AOI21_X1 U3964 ( .B1(n3149), .B2(n3148), .A(n3146), .ZN(n3147) );
  INV_X1 U3965 ( .A(n3147), .ZN(n3150) );
  NAND2_X1 U3966 ( .A1(n3150), .A2(n2221), .ZN(n3175) );
  OAI22_X1 U3967 ( .A1(n3221), .A2(n3600), .B1(n3599), .B2(n3177), .ZN(n3151)
         );
  XNOR2_X1 U3968 ( .A(n3151), .B(n3591), .ZN(n3155) );
  OR2_X1 U3969 ( .A1(n3221), .A2(n3601), .ZN(n3154) );
  NAND2_X1 U3970 ( .A1(n3152), .A2(n2878), .ZN(n3153) );
  NAND2_X1 U3971 ( .A1(n3154), .A2(n3153), .ZN(n3156) );
  XNOR2_X1 U3972 ( .A(n3155), .B(n3156), .ZN(n3174) );
  INV_X1 U3973 ( .A(n3155), .ZN(n3157) );
  OAI22_X1 U3974 ( .A1(n3269), .A2(n3600), .B1(n3599), .B2(n3168), .ZN(n3158)
         );
  XNOR2_X1 U3975 ( .A(n3158), .B(n3591), .ZN(n3162) );
  OR2_X1 U3976 ( .A1(n3269), .A2(n3601), .ZN(n3161) );
  NAND2_X1 U3977 ( .A1(n3159), .A2(n2878), .ZN(n3160) );
  AND2_X1 U3978 ( .A1(n3161), .A2(n3160), .ZN(n3163) );
  INV_X1 U3979 ( .A(n3162), .ZN(n3165) );
  INV_X1 U3980 ( .A(n3163), .ZN(n3164) );
  NAND2_X1 U3981 ( .A1(n3165), .A2(n3164), .ZN(n3261) );
  NAND2_X1 U3982 ( .A1(n2194), .A2(n3261), .ZN(n3166) );
  XNOR2_X1 U3983 ( .A(n3262), .B(n3166), .ZN(n3173) );
  INV_X1 U3984 ( .A(n4509), .ZN(n3171) );
  OAI21_X1 U3985 ( .B1(n3755), .B2(n3310), .A(n3167), .ZN(n3170) );
  OAI22_X1 U3986 ( .A1(n3770), .A2(n3221), .B1(n3768), .B2(n3168), .ZN(n3169)
         );
  AOI211_X1 U3987 ( .C1(n3171), .C2(n3757), .A(n3170), .B(n3169), .ZN(n3172)
         );
  OAI21_X1 U3988 ( .B1(n3173), .B2(n3759), .A(n3172), .ZN(U3218) );
  XOR2_X1 U3989 ( .A(n3175), .B(n3174), .Z(n3176) );
  NAND2_X1 U3990 ( .A1(n3176), .A2(n3764), .ZN(n3182) );
  OAI22_X1 U3991 ( .A1(n3770), .A2(n3178), .B1(n3768), .B2(n3177), .ZN(n3179)
         );
  AOI211_X1 U3992 ( .C1(n3772), .C2(n3960), .A(n3180), .B(n3179), .ZN(n3181)
         );
  OAI211_X1 U3993 ( .C1(n3776), .C2(n3183), .A(n3182), .B(n3181), .ZN(U3210)
         );
  INV_X1 U3994 ( .A(n3831), .ZN(n3184) );
  AND2_X1 U3995 ( .A1(n3184), .A2(n3820), .ZN(n3891) );
  XNOR2_X1 U3996 ( .A(n3185), .B(n3891), .ZN(n3202) );
  XOR2_X1 U3997 ( .A(n3891), .B(n3186), .Z(n3187) );
  NAND2_X1 U3998 ( .A1(n3187), .A2(n2715), .ZN(n3200) );
  AOI22_X1 U3999 ( .A1(n3958), .A2(n4346), .B1(n4345), .B2(n3263), .ZN(n3188)
         );
  OAI211_X1 U4000 ( .C1(n3269), .C2(n4349), .A(n3200), .B(n3188), .ZN(n3189)
         );
  AOI21_X1 U4001 ( .B1(n3202), .B2(n4340), .A(n3189), .ZN(n3194) );
  INV_X1 U4002 ( .A(n3190), .ZN(n3191) );
  AOI21_X1 U4003 ( .B1(n3263), .B2(n3191), .A(n3228), .ZN(n3197) );
  AOI22_X1 U4004 ( .A1(n3197), .A2(n3279), .B1(REG1_REG_9__SCAN_IN), .B2(n4549), .ZN(n3192) );
  OAI21_X1 U4005 ( .B1(n3194), .B2(n4549), .A(n3192), .ZN(U3527) );
  AOI22_X1 U4006 ( .A1(n3197), .A2(n3362), .B1(REG0_REG_9__SCAN_IN), .B2(n4544), .ZN(n3193) );
  OAI21_X1 U4007 ( .B1(n3194), .B2(n4544), .A(n3193), .ZN(U3485) );
  INV_X1 U4008 ( .A(n4166), .ZN(n4252) );
  OAI22_X1 U4009 ( .A1(n3273), .A2(n4508), .B1(n2504), .B2(n4511), .ZN(n3196)
         );
  OAI22_X1 U4010 ( .A1(n4111), .A2(n3269), .B1(n3388), .B2(n4113), .ZN(n3195)
         );
  AOI211_X1 U4011 ( .C1(n4252), .C2(n3263), .A(n3196), .B(n3195), .ZN(n3199)
         );
  NAND2_X1 U4012 ( .A1(n3197), .A2(n4514), .ZN(n3198) );
  OAI211_X1 U4013 ( .C1(n3200), .C2(n4520), .A(n3199), .B(n3198), .ZN(n3201)
         );
  AOI21_X1 U4014 ( .B1(n4159), .B2(n3202), .A(n3201), .ZN(n3203) );
  INV_X1 U4015 ( .A(n3203), .ZN(U3281) );
  AOI22_X1 U4016 ( .A1(n4252), .A2(n3204), .B1(n4254), .B2(n3962), .ZN(n3209)
         );
  OAI22_X1 U4017 ( .A1(n4511), .A2(n2267), .B1(n3205), .B2(n4508), .ZN(n3206)
         );
  AOI21_X1 U4018 ( .B1(n4514), .B2(n3207), .A(n3206), .ZN(n3208) );
  OAI211_X1 U4019 ( .C1(n3240), .C2(n4111), .A(n3209), .B(n3208), .ZN(n3210)
         );
  AOI21_X1 U4020 ( .B1(n3211), .B2(n4159), .A(n3210), .ZN(n3212) );
  OAI21_X1 U4021 ( .B1(n3213), .B2(n4419), .A(n3212), .ZN(U3285) );
  NOR2_X1 U4022 ( .A1(n4520), .A2(n4206), .ZN(n3341) );
  INV_X1 U4023 ( .A(n3341), .ZN(n3237) );
  OAI22_X1 U4024 ( .A1(n4511), .A2(n3215), .B1(n3214), .B2(n4508), .ZN(n3216)
         );
  AOI21_X1 U4025 ( .B1(n3217), .B2(n4514), .A(n3216), .ZN(n3220) );
  AOI22_X1 U4026 ( .A1(n4252), .A2(n3218), .B1(n4248), .B2(n2694), .ZN(n3219)
         );
  OAI211_X1 U4027 ( .C1(n3221), .C2(n4113), .A(n3220), .B(n3219), .ZN(n3222)
         );
  AOI21_X1 U4028 ( .B1(n3223), .B2(n4159), .A(n3222), .ZN(n3224) );
  OAI21_X1 U4029 ( .B1(n3237), .B2(n3225), .A(n3224), .ZN(U3284) );
  AND2_X1 U4030 ( .A1(n3828), .A2(n3833), .ZN(n3888) );
  XOR2_X1 U4031 ( .A(n3888), .B(n3226), .Z(n3276) );
  XOR2_X1 U4032 ( .A(n3227), .B(n3888), .Z(n3278) );
  NAND2_X1 U4033 ( .A1(n3278), .A2(n4159), .ZN(n3236) );
  INV_X1 U4034 ( .A(n3228), .ZN(n3230) );
  INV_X1 U4035 ( .A(n3229), .ZN(n3293) );
  AOI21_X1 U4036 ( .B1(n3302), .B2(n3230), .A(n3293), .ZN(n3281) );
  AOI22_X1 U4037 ( .A1(n4252), .A2(n3302), .B1(n4254), .B2(n3957), .ZN(n3233)
         );
  INV_X1 U4038 ( .A(n3315), .ZN(n3231) );
  INV_X1 U4039 ( .A(n4508), .ZN(n4250) );
  AOI22_X1 U4040 ( .A1(n4520), .A2(REG2_REG_10__SCAN_IN), .B1(n3231), .B2(
        n4250), .ZN(n3232) );
  OAI211_X1 U4041 ( .C1(n3310), .C2(n4111), .A(n3233), .B(n3232), .ZN(n3234)
         );
  AOI21_X1 U4042 ( .B1(n3281), .B2(n4514), .A(n3234), .ZN(n3235) );
  OAI211_X1 U40430 ( .C1(n3276), .C2(n3237), .A(n3236), .B(n3235), .ZN(U3280)
         );
  OAI22_X1 U4044 ( .A1(n4511), .A2(n3238), .B1(REG3_REG_3__SCAN_IN), .B2(n4508), .ZN(n3242) );
  OAI22_X1 U4045 ( .A1(n3240), .A2(n4113), .B1(n4166), .B2(n3239), .ZN(n3241)
         );
  AOI211_X1 U4046 ( .C1(n4514), .C2(n3243), .A(n3242), .B(n3241), .ZN(n3246)
         );
  NAND2_X1 U4047 ( .A1(n3244), .A2(n4159), .ZN(n3245) );
  OAI211_X1 U4048 ( .C1(n3247), .C2(n4520), .A(n3246), .B(n3245), .ZN(U3287)
         );
  AOI21_X1 U4049 ( .B1(n3249), .B2(n3258), .A(n3248), .ZN(n3252) );
  OAI21_X1 U4050 ( .B1(n3252), .B2(n3251), .A(n4466), .ZN(n3250) );
  AOI21_X1 U4051 ( .B1(n3252), .B2(n3251), .A(n3250), .ZN(n3260) );
  OAI211_X1 U4052 ( .C1(n3255), .C2(n3254), .A(n4502), .B(n3253), .ZN(n3257)
         );
  NOR2_X1 U4053 ( .A1(STATE_REG_SCAN_IN), .A2(n2539), .ZN(n3489) );
  AOI21_X1 U4054 ( .B1(n4501), .B2(ADDR_REG_13__SCAN_IN), .A(n3489), .ZN(n3256) );
  OAI211_X1 U4055 ( .C1(n4507), .C2(n3258), .A(n3257), .B(n3256), .ZN(n3259)
         );
  OR2_X1 U4056 ( .A1(n3260), .A2(n3259), .ZN(U3253) );
  NAND2_X1 U4057 ( .A1(n3959), .A2(n2878), .ZN(n3265) );
  NAND2_X1 U4058 ( .A1(n3263), .A2(n2044), .ZN(n3264) );
  NAND2_X1 U4059 ( .A1(n3265), .A2(n3264), .ZN(n3266) );
  XNOR2_X1 U4060 ( .A(n3266), .B(n3602), .ZN(n3299) );
  OAI22_X1 U4061 ( .A1(n3310), .A2(n3601), .B1(n3600), .B2(n3268), .ZN(n3298)
         );
  XNOR2_X1 U4062 ( .A(n3299), .B(n3298), .ZN(n3300) );
  XNOR2_X1 U4063 ( .A(n3301), .B(n3300), .ZN(n3267) );
  NAND2_X1 U4064 ( .A1(n3267), .A2(n3764), .ZN(n3272) );
  NOR2_X1 U4065 ( .A1(STATE_REG_SCAN_IN), .A2(n2501), .ZN(n4441) );
  OAI22_X1 U4066 ( .A1(n3770), .A2(n3269), .B1(n3768), .B2(n3268), .ZN(n3270)
         );
  AOI211_X1 U4067 ( .C1(n3772), .C2(n3958), .A(n4441), .B(n3270), .ZN(n3271)
         );
  OAI211_X1 U4068 ( .C1(n3776), .C2(n3273), .A(n3272), .B(n3271), .ZN(U3228)
         );
  OAI22_X1 U4069 ( .A1(n3439), .A2(n4337), .B1(n4203), .B2(n3309), .ZN(n3274)
         );
  AOI21_X1 U4070 ( .B1(n4333), .B2(n3959), .A(n3274), .ZN(n3275) );
  OAI21_X1 U4071 ( .B1(n3276), .B2(n4206), .A(n3275), .ZN(n3277) );
  AOI21_X1 U4072 ( .B1(n4340), .B2(n3278), .A(n3277), .ZN(n3283) );
  AOI22_X1 U4073 ( .A1(n3281), .A2(n3279), .B1(REG1_REG_10__SCAN_IN), .B2(
        n4549), .ZN(n3280) );
  OAI21_X1 U4074 ( .B1(n3283), .B2(n4549), .A(n3280), .ZN(U3528) );
  AOI22_X1 U4075 ( .A1(n3281), .A2(n3362), .B1(REG0_REG_10__SCAN_IN), .B2(
        n4544), .ZN(n3282) );
  OAI21_X1 U4076 ( .B1(n3283), .B2(n4544), .A(n3282), .ZN(U3487) );
  INV_X1 U4077 ( .A(n3284), .ZN(n3285) );
  AOI21_X1 U4078 ( .B1(n3894), .B2(n3286), .A(n3285), .ZN(n3358) );
  AOI22_X1 U4079 ( .A1(n3956), .A2(n4346), .B1(n4345), .B2(n3287), .ZN(n3291)
         );
  XNOR2_X1 U4080 ( .A(n3288), .B(n3894), .ZN(n3289) );
  NAND2_X1 U4081 ( .A1(n3289), .A2(n2715), .ZN(n3290) );
  OAI211_X1 U4082 ( .C1(n3358), .C2(n4185), .A(n3291), .B(n3290), .ZN(n3360)
         );
  NAND2_X1 U4083 ( .A1(n3360), .A2(n4215), .ZN(n3297) );
  OAI22_X1 U4084 ( .A1(n4511), .A2(n3292), .B1(n3392), .B2(n4508), .ZN(n3295)
         );
  OAI21_X1 U4085 ( .B1(n3293), .B2(n3387), .A(n3347), .ZN(n3366) );
  NOR2_X1 U4086 ( .A1(n3366), .A2(n4213), .ZN(n3294) );
  AOI211_X1 U4087 ( .C1(n4248), .C2(n3958), .A(n3295), .B(n3294), .ZN(n3296)
         );
  OAI211_X1 U4088 ( .C1(n3358), .C2(n4246), .A(n3297), .B(n3296), .ZN(U3279)
         );
  AOI22_X1 U4089 ( .A1(n3958), .A2(n2857), .B1(n2043), .B2(n3302), .ZN(n3381)
         );
  NAND2_X1 U4090 ( .A1(n3958), .A2(n2043), .ZN(n3304) );
  NAND2_X1 U4091 ( .A1(n3302), .A2(n2044), .ZN(n3303) );
  NAND2_X1 U4092 ( .A1(n3304), .A2(n3303), .ZN(n3305) );
  XNOR2_X1 U4093 ( .A(n3305), .B(n3602), .ZN(n3380) );
  XOR2_X1 U4094 ( .A(n3381), .B(n3380), .Z(n3306) );
  AOI21_X1 U4095 ( .B1(n3307), .B2(n3306), .A(n3759), .ZN(n3308) );
  NAND2_X1 U4096 ( .A1(n3308), .A2(n3383), .ZN(n3314) );
  NAND2_X1 U4097 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4446) );
  INV_X1 U4098 ( .A(n4446), .ZN(n3312) );
  OAI22_X1 U4099 ( .A1(n3770), .A2(n3310), .B1(n3768), .B2(n3309), .ZN(n3311)
         );
  AOI211_X1 U4100 ( .C1(n3772), .C2(n3957), .A(n3312), .B(n3311), .ZN(n3313)
         );
  OAI211_X1 U4101 ( .C1(n3776), .C2(n3315), .A(n3314), .B(n3313), .ZN(U3214)
         );
  INV_X1 U4102 ( .A(n3344), .ZN(n3317) );
  OAI21_X1 U4103 ( .B1(n3316), .B2(n3317), .A(n3343), .ZN(n3320) );
  NAND2_X1 U4104 ( .A1(n3319), .A2(n3318), .ZN(n3872) );
  XNOR2_X1 U4105 ( .A(n3320), .B(n3872), .ZN(n3324) );
  NAND2_X1 U4106 ( .A1(n3326), .A2(n4345), .ZN(n3322) );
  NAND2_X1 U4107 ( .A1(n3956), .A2(n4333), .ZN(n3321) );
  OAI211_X1 U4108 ( .C1(n3769), .C2(n4337), .A(n3322), .B(n3321), .ZN(n3323)
         );
  AOI21_X1 U4109 ( .B1(n3324), .B2(n2715), .A(n3323), .ZN(n3417) );
  XNOR2_X1 U4110 ( .A(n3325), .B(n3872), .ZN(n3416) );
  INV_X1 U4111 ( .A(n3336), .ZN(n3328) );
  NAND2_X1 U4112 ( .A1(n3349), .A2(n3326), .ZN(n3327) );
  NAND2_X1 U4113 ( .A1(n3328), .A2(n3327), .ZN(n3424) );
  NOR2_X1 U4114 ( .A1(n3424), .A2(n4213), .ZN(n3330) );
  OAI22_X1 U4115 ( .A1(n4511), .A2(n3249), .B1(n3492), .B2(n4508), .ZN(n3329)
         );
  AOI211_X1 U4116 ( .C1(n3416), .C2(n4159), .A(n3330), .B(n3329), .ZN(n3331)
         );
  OAI21_X1 U4117 ( .B1(n4520), .B2(n3417), .A(n3331), .ZN(U3277) );
  INV_X1 U4118 ( .A(n3332), .ZN(n3333) );
  AOI21_X1 U4119 ( .B1(n3889), .B2(n3334), .A(n3333), .ZN(n3406) );
  XNOR2_X1 U4120 ( .A(n3335), .B(n3889), .ZN(n3409) );
  OAI21_X1 U4121 ( .B1(n3336), .B2(n3639), .A(n3371), .ZN(n3415) );
  OAI22_X1 U4122 ( .A1(n4511), .A2(n4478), .B1(n3638), .B2(n4508), .ZN(n3338)
         );
  OAI22_X1 U4123 ( .A1(n4350), .A2(n4113), .B1(n4166), .B2(n3639), .ZN(n3337)
         );
  AOI211_X1 U4124 ( .C1(n4248), .C2(n3955), .A(n3338), .B(n3337), .ZN(n3339)
         );
  OAI21_X1 U4125 ( .B1(n3415), .B2(n4213), .A(n3339), .ZN(n3340) );
  AOI21_X1 U4126 ( .B1(n3409), .B2(n3341), .A(n3340), .ZN(n3342) );
  OAI21_X1 U4127 ( .B1(n3406), .B2(n4239), .A(n3342), .ZN(U3276) );
  AND2_X1 U4128 ( .A1(n3344), .A2(n3343), .ZN(n3879) );
  INV_X1 U4129 ( .A(n3879), .ZN(n3345) );
  XNOR2_X1 U4130 ( .A(n3346), .B(n3345), .ZN(n3396) );
  NAND2_X1 U4131 ( .A1(n3347), .A2(n3433), .ZN(n3348) );
  NAND2_X1 U4132 ( .A1(n3349), .A2(n3348), .ZN(n3404) );
  OAI22_X1 U4133 ( .A1(n4511), .A2(n3350), .B1(n3437), .B2(n4508), .ZN(n3351)
         );
  AOI21_X1 U4134 ( .B1(n3433), .B2(n4252), .A(n3351), .ZN(n3353) );
  AOI22_X1 U4135 ( .A1(n4254), .A2(n3955), .B1(n4248), .B2(n3957), .ZN(n3352)
         );
  OAI211_X1 U4136 ( .C1(n3404), .C2(n4213), .A(n3353), .B(n3352), .ZN(n3356)
         );
  XNOR2_X1 U4137 ( .A(n3316), .B(n3879), .ZN(n3354) );
  NAND2_X1 U4138 ( .A1(n3354), .A2(n2715), .ZN(n3394) );
  NOR2_X1 U4139 ( .A1(n3394), .A2(n4419), .ZN(n3355) );
  AOI211_X1 U4140 ( .C1(n4159), .C2(n3396), .A(n3356), .B(n3355), .ZN(n3357)
         );
  INV_X1 U4141 ( .A(n3357), .ZN(U3278) );
  OAI22_X1 U4142 ( .A1(n3358), .A2(n4530), .B1(n3388), .B2(n4349), .ZN(n3359)
         );
  NOR2_X1 U4143 ( .A1(n3360), .A2(n3359), .ZN(n3363) );
  MUX2_X1 U4144 ( .A(n2350), .B(n3363), .S(n4552), .Z(n3361) );
  OAI21_X1 U4145 ( .B1(n4343), .B2(n3366), .A(n3361), .ZN(U3529) );
  INV_X1 U4146 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3364) );
  MUX2_X1 U4147 ( .A(n3364), .B(n3363), .S(n4546), .Z(n3365) );
  OAI21_X1 U4148 ( .B1(n3366), .B2(n4404), .A(n3365), .ZN(U3489) );
  AOI21_X1 U4149 ( .B1(n3367), .B2(n3875), .A(n4206), .ZN(n3369) );
  NAND2_X1 U4150 ( .A1(n3369), .A2(n3368), .ZN(n3446) );
  XNOR2_X1 U4151 ( .A(n3370), .B(n3875), .ZN(n3448) );
  NAND2_X1 U4152 ( .A1(n3448), .A2(n4159), .ZN(n3379) );
  INV_X1 U4153 ( .A(n3371), .ZN(n3372) );
  OAI21_X1 U4154 ( .B1(n3372), .B2(n3767), .A(n3470), .ZN(n3453) );
  INV_X1 U4155 ( .A(n3453), .ZN(n3377) );
  AOI22_X1 U4156 ( .A1(n4254), .A2(n4334), .B1(n4248), .B2(n3954), .ZN(n3375)
         );
  INV_X1 U4157 ( .A(n3775), .ZN(n3373) );
  AOI22_X1 U4158 ( .A1(n4520), .A2(REG2_REG_15__SCAN_IN), .B1(n3373), .B2(
        n4250), .ZN(n3374) );
  OAI211_X1 U4159 ( .C1(n3767), .C2(n4166), .A(n3375), .B(n3374), .ZN(n3376)
         );
  AOI21_X1 U4160 ( .B1(n3377), .B2(n4514), .A(n3376), .ZN(n3378) );
  OAI211_X1 U4161 ( .C1(n4520), .C2(n3446), .A(n3379), .B(n3378), .ZN(U3275)
         );
  OAI22_X1 U4162 ( .A1(n3439), .A2(n3600), .B1(n3599), .B2(n3387), .ZN(n3384)
         );
  XNOR2_X1 U4163 ( .A(n3384), .B(n3602), .ZN(n3425) );
  OAI22_X1 U4164 ( .A1(n3439), .A2(n3601), .B1(n3600), .B2(n3387), .ZN(n3426)
         );
  XNOR2_X1 U4165 ( .A(n3425), .B(n3426), .ZN(n3385) );
  XNOR2_X1 U4166 ( .A(n3427), .B(n3385), .ZN(n3386) );
  NAND2_X1 U4167 ( .A1(n3386), .A2(n3764), .ZN(n3391) );
  AND2_X1 U4168 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4462) );
  OAI22_X1 U4169 ( .A1(n3770), .A2(n3388), .B1(n3768), .B2(n3387), .ZN(n3389)
         );
  AOI211_X1 U4170 ( .C1(n3772), .C2(n3956), .A(n4462), .B(n3389), .ZN(n3390)
         );
  OAI211_X1 U4171 ( .C1(n3776), .C2(n3392), .A(n3391), .B(n3390), .ZN(U3233)
         );
  AOI22_X1 U4172 ( .A1(n3957), .A2(n4333), .B1(n4346), .B2(n3955), .ZN(n3393)
         );
  OAI211_X1 U4173 ( .C1(n4203), .C2(n3438), .A(n3394), .B(n3393), .ZN(n3395)
         );
  INV_X1 U4174 ( .A(n3395), .ZN(n3398) );
  NAND2_X1 U4175 ( .A1(n3396), .A2(n4340), .ZN(n3397) );
  NAND2_X1 U4176 ( .A1(n3398), .A2(n3397), .ZN(n3401) );
  MUX2_X1 U4177 ( .A(n3401), .B(REG1_REG_12__SCAN_IN), .S(n4549), .Z(n3399) );
  INV_X1 U4178 ( .A(n3399), .ZN(n3400) );
  OAI21_X1 U4179 ( .B1(n4343), .B2(n3404), .A(n3400), .ZN(U3530) );
  MUX2_X1 U4180 ( .A(REG0_REG_12__SCAN_IN), .B(n3401), .S(n4546), .Z(n3402) );
  INV_X1 U4181 ( .A(n3402), .ZN(n3403) );
  OAI21_X1 U4182 ( .B1(n3404), .B2(n4404), .A(n3403), .ZN(U3491) );
  INV_X1 U4183 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4184 ( .A1(n3953), .A2(n4346), .B1(n4345), .B2(n3503), .ZN(n3405)
         );
  OAI21_X1 U4185 ( .B1(n3640), .B2(n4349), .A(n3405), .ZN(n3408) );
  INV_X1 U4186 ( .A(n4340), .ZN(n4538) );
  NOR2_X1 U4187 ( .A1(n3406), .A2(n4538), .ZN(n3407) );
  AOI211_X1 U4188 ( .C1(n3409), .C2(n2715), .A(n3408), .B(n3407), .ZN(n3412)
         );
  MUX2_X1 U4189 ( .A(n3410), .B(n3412), .S(n4546), .Z(n3411) );
  OAI21_X1 U4190 ( .B1(n3415), .B2(n4404), .A(n3411), .ZN(U3495) );
  MUX2_X1 U4191 ( .A(n3413), .B(n3412), .S(n4552), .Z(n3414) );
  OAI21_X1 U4192 ( .B1(n4343), .B2(n3415), .A(n3414), .ZN(U3532) );
  NAND2_X1 U4193 ( .A1(n3416), .A2(n4340), .ZN(n3418) );
  NAND2_X1 U4194 ( .A1(n3418), .A2(n3417), .ZN(n3421) );
  MUX2_X1 U4195 ( .A(REG1_REG_13__SCAN_IN), .B(n3421), .S(n4552), .Z(n3419) );
  INV_X1 U4196 ( .A(n3419), .ZN(n3420) );
  OAI21_X1 U4197 ( .B1(n4343), .B2(n3424), .A(n3420), .ZN(U3531) );
  MUX2_X1 U4198 ( .A(REG0_REG_13__SCAN_IN), .B(n3421), .S(n4546), .Z(n3422) );
  INV_X1 U4199 ( .A(n3422), .ZN(n3423) );
  OAI21_X1 U4200 ( .B1(n3424), .B2(n4404), .A(n3423), .ZN(U3493) );
  OAI21_X1 U4201 ( .B1(n3427), .B2(n3426), .A(n3425), .ZN(n3429) );
  NAND2_X1 U4202 ( .A1(n3427), .A2(n3426), .ZN(n3428) );
  NAND2_X1 U4203 ( .A1(n3956), .A2(n2878), .ZN(n3431) );
  NAND2_X1 U4204 ( .A1(n3433), .A2(n2044), .ZN(n3430) );
  NAND2_X1 U4205 ( .A1(n3431), .A2(n3430), .ZN(n3432) );
  XNOR2_X1 U4206 ( .A(n3432), .B(n3591), .ZN(n3435) );
  AOI22_X1 U4207 ( .A1(n3956), .A2(n2857), .B1(n2043), .B2(n3433), .ZN(n3434)
         );
  OR2_X1 U4208 ( .A1(n3435), .A2(n3434), .ZN(n3479) );
  NAND2_X1 U4209 ( .A1(n3435), .A2(n3434), .ZN(n3481) );
  NAND2_X1 U4210 ( .A1(n3479), .A2(n3481), .ZN(n3436) );
  XNOR2_X1 U4211 ( .A(n3480), .B(n3436), .ZN(n3444) );
  INV_X1 U4212 ( .A(n3437), .ZN(n3442) );
  NAND2_X1 U4213 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4468) );
  OAI21_X1 U4214 ( .B1(n3755), .B2(n3640), .A(n4468), .ZN(n3441) );
  OAI22_X1 U4215 ( .A1(n3770), .A2(n3439), .B1(n3768), .B2(n3438), .ZN(n3440)
         );
  AOI211_X1 U4216 ( .C1(n3442), .C2(n3757), .A(n3441), .B(n3440), .ZN(n3443)
         );
  OAI21_X1 U4217 ( .B1(n3444), .B2(n3759), .A(n3443), .ZN(U3221) );
  AOI22_X1 U4218 ( .A1(n4334), .A2(n4346), .B1(n3512), .B2(n4345), .ZN(n3445)
         );
  OAI211_X1 U4219 ( .C1(n3769), .C2(n4349), .A(n3446), .B(n3445), .ZN(n3447)
         );
  AOI21_X1 U4220 ( .B1(n3448), .B2(n4340), .A(n3447), .ZN(n3451) );
  MUX2_X1 U4221 ( .A(n3449), .B(n3451), .S(n4546), .Z(n3450) );
  OAI21_X1 U4222 ( .B1(n3453), .B2(n4404), .A(n3450), .ZN(U3497) );
  MUX2_X1 U4223 ( .A(n2348), .B(n3451), .S(n4552), .Z(n3452) );
  OAI21_X1 U4224 ( .B1(n4343), .B2(n3453), .A(n3452), .ZN(U3533) );
  INV_X1 U4225 ( .A(n3454), .ZN(n3786) );
  NAND2_X1 U4226 ( .A1(n3786), .A2(n4197), .ZN(n3873) );
  XNOR2_X1 U4227 ( .A(n3455), .B(n3873), .ZN(n3456) );
  NAND2_X1 U4228 ( .A1(n3456), .A2(n2715), .ZN(n4336) );
  NAND2_X1 U4229 ( .A1(n4230), .A2(n3458), .ZN(n3459) );
  XOR2_X1 U4230 ( .A(n3873), .B(n3459), .Z(n4341) );
  NAND2_X1 U4231 ( .A1(n4341), .A2(n4159), .ZN(n3467) );
  INV_X1 U4232 ( .A(n4220), .ZN(n3460) );
  OAI21_X1 U4233 ( .B1(n3469), .B2(n3699), .A(n3460), .ZN(n4405) );
  INV_X1 U4234 ( .A(n4405), .ZN(n3465) );
  AOI22_X1 U4235 ( .A1(n4254), .A2(n3952), .B1(n4248), .B2(n4334), .ZN(n3463)
         );
  INV_X1 U4236 ( .A(n3461), .ZN(n3703) );
  AOI22_X1 U4237 ( .A1(n4520), .A2(REG2_REG_17__SCAN_IN), .B1(n3703), .B2(
        n4250), .ZN(n3462) );
  OAI211_X1 U4238 ( .C1(n3699), .C2(n4166), .A(n3463), .B(n3462), .ZN(n3464)
         );
  AOI21_X1 U4239 ( .B1(n3465), .B2(n4514), .A(n3464), .ZN(n3466) );
  OAI211_X1 U4240 ( .C1(n4520), .C2(n4336), .A(n3467), .B(n3466), .ZN(U3273)
         );
  INV_X1 U4241 ( .A(n3881), .ZN(n3468) );
  OAI21_X1 U4242 ( .B1(n2594), .B2(n3468), .A(n4230), .ZN(n4356) );
  AOI21_X1 U4243 ( .B1(n4344), .B2(n3470), .A(n3469), .ZN(n4353) );
  AOI22_X1 U4244 ( .A1(n4254), .A2(n4347), .B1(n4248), .B2(n3953), .ZN(n3473)
         );
  INV_X1 U4245 ( .A(n3471), .ZN(n3692) );
  AOI22_X1 U4246 ( .A1(n4520), .A2(REG2_REG_16__SCAN_IN), .B1(n3692), .B2(
        n4250), .ZN(n3472) );
  OAI211_X1 U4247 ( .C1(n3689), .C2(n4166), .A(n3473), .B(n3472), .ZN(n3477)
         );
  OAI211_X1 U4248 ( .C1(n3475), .C2(n3881), .A(n3474), .B(n2715), .ZN(n4354)
         );
  NOR2_X1 U4249 ( .A1(n4354), .A2(n4520), .ZN(n3476) );
  AOI211_X1 U4250 ( .C1(n4353), .C2(n4514), .A(n3477), .B(n3476), .ZN(n3478)
         );
  OAI21_X1 U4251 ( .B1(n4239), .B2(n4356), .A(n3478), .ZN(U3274) );
  NAND2_X1 U4252 ( .A1(n3480), .A2(n3479), .ZN(n3482) );
  NAND2_X1 U4253 ( .A1(n3482), .A2(n3481), .ZN(n3500) );
  OAI22_X1 U4254 ( .A1(n3640), .A2(n3600), .B1(n3599), .B2(n3486), .ZN(n3483)
         );
  XNOR2_X1 U4255 ( .A(n3501), .B(n3499), .ZN(n3484) );
  XNOR2_X1 U4256 ( .A(n3500), .B(n3484), .ZN(n3485) );
  NAND2_X1 U4257 ( .A1(n3485), .A2(n3764), .ZN(n3491) );
  OAI22_X1 U4258 ( .A1(n3770), .A2(n3487), .B1(n3768), .B2(n3486), .ZN(n3488)
         );
  AOI211_X1 U4259 ( .C1(n3772), .C2(n3954), .A(n3489), .B(n3488), .ZN(n3490)
         );
  OAI211_X1 U4260 ( .C1(n3776), .C2(n3492), .A(n3491), .B(n3490), .ZN(U3231)
         );
  INV_X1 U4261 ( .A(DATAI_31_), .ZN(n3496) );
  OR4_X1 U4262 ( .A1(n3494), .A2(IR_REG_30__SCAN_IN), .A3(n3493), .A4(U3149), 
        .ZN(n3495) );
  OAI21_X1 U4263 ( .B1(STATE_REG_SCAN_IN), .B2(n3496), .A(n3495), .ZN(U3321)
         );
  INV_X1 U4264 ( .A(DATAI_29_), .ZN(n4591) );
  NAND2_X1 U4265 ( .A1(n3497), .A2(STATE_REG_SCAN_IN), .ZN(n3498) );
  OAI21_X1 U4266 ( .B1(STATE_REG_SCAN_IN), .B2(n4591), .A(n3498), .ZN(U3323)
         );
  OAI22_X1 U4267 ( .A1(n3769), .A2(n3600), .B1(n3599), .B2(n3639), .ZN(n3502)
         );
  XNOR2_X1 U4268 ( .A(n3502), .B(n3602), .ZN(n3508) );
  OR2_X1 U4269 ( .A1(n3769), .A2(n3601), .ZN(n3505) );
  NAND2_X1 U4270 ( .A1(n3503), .A2(n2878), .ZN(n3504) );
  NAND2_X1 U4271 ( .A1(n3505), .A2(n3504), .ZN(n3509) );
  NAND2_X1 U4272 ( .A1(n3508), .A2(n3509), .ZN(n3636) );
  OAI22_X1 U4273 ( .A1(n4350), .A2(n3600), .B1(n3599), .B2(n3767), .ZN(n3506)
         );
  XOR2_X1 U4274 ( .A(n3602), .B(n3506), .Z(n3507) );
  INV_X1 U4275 ( .A(n3507), .ZN(n3516) );
  INV_X1 U4276 ( .A(n3508), .ZN(n3511) );
  INV_X1 U4277 ( .A(n3509), .ZN(n3510) );
  NAND2_X1 U4278 ( .A1(n3511), .A2(n3510), .ZN(n3635) );
  OR2_X1 U4279 ( .A1(n3516), .A2(n3635), .ZN(n3684) );
  NAND2_X1 U4280 ( .A1(n3953), .A2(n2857), .ZN(n3514) );
  NAND2_X1 U4281 ( .A1(n3512), .A2(n2878), .ZN(n3513) );
  NAND2_X1 U4282 ( .A1(n3514), .A2(n3513), .ZN(n3762) );
  AND2_X1 U4283 ( .A1(n3684), .A2(n3762), .ZN(n3515) );
  NAND2_X1 U4284 ( .A1(n3685), .A2(n3515), .ZN(n3520) );
  NAND2_X1 U4285 ( .A1(n3634), .A2(n3636), .ZN(n3518) );
  AND2_X1 U4286 ( .A1(n3635), .A2(n3516), .ZN(n3517) );
  NAND2_X1 U4287 ( .A1(n3518), .A2(n3517), .ZN(n3683) );
  OAI22_X1 U4288 ( .A1(n3700), .A2(n3601), .B1(n3600), .B2(n3689), .ZN(n3522)
         );
  OAI22_X1 U4289 ( .A1(n3700), .A2(n3600), .B1(n3599), .B2(n3689), .ZN(n3519)
         );
  XNOR2_X1 U4290 ( .A(n3519), .B(n3602), .ZN(n3521) );
  XOR2_X1 U4291 ( .A(n3522), .B(n3521), .Z(n3688) );
  INV_X1 U4292 ( .A(n3521), .ZN(n3524) );
  INV_X1 U4293 ( .A(n3522), .ZN(n3523) );
  NAND2_X1 U4294 ( .A1(n3524), .A2(n3523), .ZN(n3525) );
  NAND2_X1 U4295 ( .A1(n4347), .A2(n2878), .ZN(n3527) );
  NAND2_X1 U4296 ( .A1(n4332), .A2(n2044), .ZN(n3526) );
  NAND2_X1 U4297 ( .A1(n3527), .A2(n3526), .ZN(n3528) );
  XNOR2_X1 U4298 ( .A(n3528), .B(n3602), .ZN(n3697) );
  NAND2_X1 U4299 ( .A1(n4347), .A2(n2857), .ZN(n3530) );
  NAND2_X1 U4300 ( .A1(n4332), .A2(n2043), .ZN(n3529) );
  NAND2_X1 U4301 ( .A1(n3530), .A2(n3529), .ZN(n3696) );
  NOR2_X1 U4302 ( .A1(n3697), .A2(n3696), .ZN(n3533) );
  INV_X1 U4303 ( .A(n3697), .ZN(n3532) );
  INV_X1 U4304 ( .A(n3696), .ZN(n3531) );
  OAI22_X1 U4305 ( .A1(n4338), .A2(n3600), .B1(n3599), .B2(n4219), .ZN(n3534)
         );
  XNOR2_X1 U4306 ( .A(n3534), .B(n3602), .ZN(n3535) );
  OAI22_X1 U4307 ( .A1(n4338), .A2(n3601), .B1(n3600), .B2(n4219), .ZN(n3536)
         );
  AND2_X1 U4308 ( .A1(n3535), .A2(n3536), .ZN(n3737) );
  INV_X1 U4309 ( .A(n3535), .ZN(n3538) );
  INV_X1 U4310 ( .A(n3536), .ZN(n3537) );
  NAND2_X1 U4311 ( .A1(n3538), .A2(n3537), .ZN(n3738) );
  OAI22_X1 U4312 ( .A1(n4224), .A2(n3601), .B1(n3600), .B2(n4209), .ZN(n3544)
         );
  NAND2_X1 U4313 ( .A1(n4179), .A2(n2878), .ZN(n3541) );
  NAND2_X1 U4314 ( .A1(n3539), .A2(n2044), .ZN(n3540) );
  NAND2_X1 U4315 ( .A1(n3541), .A2(n3540), .ZN(n3542) );
  XNOR2_X1 U4316 ( .A(n3542), .B(n3602), .ZN(n3543) );
  XOR2_X1 U4317 ( .A(n3544), .B(n3543), .Z(n3659) );
  NAND2_X1 U4318 ( .A1(n3658), .A2(n3659), .ZN(n3548) );
  NAND2_X1 U4319 ( .A1(n3548), .A2(n3547), .ZN(n3715) );
  NAND2_X1 U4320 ( .A1(n4312), .A2(n2878), .ZN(n3550) );
  NAND2_X1 U4321 ( .A1(n2044), .A2(n4178), .ZN(n3549) );
  NAND2_X1 U4322 ( .A1(n3550), .A2(n3549), .ZN(n3551) );
  XNOR2_X1 U4323 ( .A(n3551), .B(n3591), .ZN(n3565) );
  NOR2_X1 U4324 ( .A1(n3600), .A2(n4188), .ZN(n3552) );
  AOI21_X1 U4325 ( .B1(n4312), .B2(n2857), .A(n3552), .ZN(n3564) );
  OR2_X1 U4326 ( .A1(n3565), .A2(n3564), .ZN(n3716) );
  NAND2_X1 U4327 ( .A1(n3715), .A2(n3716), .ZN(n3646) );
  NAND2_X1 U4328 ( .A1(n4141), .A2(n2878), .ZN(n3554) );
  NAND2_X1 U4329 ( .A1(n2044), .A2(n4311), .ZN(n3553) );
  NAND2_X1 U4330 ( .A1(n3554), .A2(n3553), .ZN(n3555) );
  XNOR2_X1 U4331 ( .A(n3555), .B(n3602), .ZN(n3665) );
  NAND2_X1 U4332 ( .A1(n4141), .A2(n2857), .ZN(n3557) );
  OR2_X1 U4333 ( .A1(n4167), .A2(n3600), .ZN(n3556) );
  NAND2_X1 U4334 ( .A1(n3557), .A2(n3556), .ZN(n3664) );
  NOR2_X1 U4335 ( .A1(n3665), .A2(n3664), .ZN(n3647) );
  NAND2_X1 U4336 ( .A1(n4292), .A2(n2043), .ZN(n3560) );
  NAND2_X1 U4337 ( .A1(n2044), .A2(n3558), .ZN(n3559) );
  NAND2_X1 U4338 ( .A1(n3560), .A2(n3559), .ZN(n3561) );
  XNOR2_X1 U4339 ( .A(n3561), .B(n3591), .ZN(n3574) );
  NOR2_X1 U4340 ( .A1(n3600), .A2(n4132), .ZN(n3562) );
  AOI21_X1 U4341 ( .B1(n4292), .B2(n2857), .A(n3562), .ZN(n3573) );
  XNOR2_X1 U4342 ( .A(n3574), .B(n3573), .ZN(n3649) );
  OAI22_X1 U4343 ( .A1(n4315), .A2(n3600), .B1(n3599), .B2(n4149), .ZN(n3563)
         );
  XNOR2_X1 U4344 ( .A(n3563), .B(n3602), .ZN(n3568) );
  OAI22_X1 U4345 ( .A1(n4315), .A2(n3601), .B1(n3600), .B2(n4149), .ZN(n3567)
         );
  NOR2_X1 U4346 ( .A1(n3568), .A2(n3567), .ZN(n3650) );
  NOR2_X1 U4347 ( .A1(n3647), .A2(n3570), .ZN(n3566) );
  NAND2_X1 U4348 ( .A1(n3565), .A2(n3564), .ZN(n3718) );
  AND2_X1 U4349 ( .A1(n3566), .A2(n3718), .ZN(n3572) );
  NAND2_X1 U4350 ( .A1(n3665), .A2(n3664), .ZN(n3725) );
  XNOR2_X1 U4351 ( .A(n3568), .B(n3567), .ZN(n3729) );
  INV_X1 U4352 ( .A(n3729), .ZN(n3569) );
  AND2_X1 U4353 ( .A1(n3725), .A2(n3569), .ZN(n3648) );
  NOR2_X1 U4354 ( .A1(n3570), .A2(n3648), .ZN(n3571) );
  OR2_X1 U4355 ( .A1(n3574), .A2(n3573), .ZN(n3577) );
  NOR2_X1 U4356 ( .A1(n3600), .A2(n4107), .ZN(n3575) );
  AOI21_X1 U4357 ( .B1(n4283), .B2(n2857), .A(n3575), .ZN(n3578) );
  OAI22_X1 U4358 ( .A1(n3653), .A2(n3600), .B1(n3599), .B2(n4107), .ZN(n3576)
         );
  XNOR2_X1 U4359 ( .A(n3576), .B(n3602), .ZN(n3709) );
  NAND2_X1 U4360 ( .A1(n3707), .A2(n3709), .ZN(n3581) );
  NAND2_X1 U4361 ( .A1(n3651), .A2(n3577), .ZN(n3580) );
  INV_X1 U4362 ( .A(n3578), .ZN(n3579) );
  NAND2_X1 U4363 ( .A1(n3580), .A2(n3579), .ZN(n3706) );
  NAND2_X1 U4364 ( .A1(n3581), .A2(n3706), .ZN(n3676) );
  NAND2_X1 U4365 ( .A1(n3950), .A2(n2043), .ZN(n3583) );
  NAND2_X1 U4366 ( .A1(n2044), .A2(n4282), .ZN(n3582) );
  NAND2_X1 U4367 ( .A1(n3583), .A2(n3582), .ZN(n3584) );
  XNOR2_X1 U4368 ( .A(n3584), .B(n3591), .ZN(n3587) );
  NOR2_X1 U4369 ( .A1(n3600), .A2(n4091), .ZN(n3585) );
  AOI21_X1 U4370 ( .B1(n3950), .B2(n2857), .A(n3585), .ZN(n3586) );
  NAND2_X1 U4371 ( .A1(n3587), .A2(n3586), .ZN(n3674) );
  NAND2_X1 U4372 ( .A1(n3676), .A2(n3674), .ZN(n3588) );
  OR2_X1 U4373 ( .A1(n3587), .A2(n3586), .ZN(n3675) );
  NAND2_X1 U4374 ( .A1(n4270), .A2(n2878), .ZN(n3590) );
  NAND2_X1 U4375 ( .A1(n2044), .A2(n3864), .ZN(n3589) );
  NAND2_X1 U4376 ( .A1(n3590), .A2(n3589), .ZN(n3592) );
  XNOR2_X1 U4377 ( .A(n3592), .B(n3591), .ZN(n3595) );
  NOR2_X1 U4378 ( .A1(n3600), .A2(n4076), .ZN(n3593) );
  AOI21_X1 U4379 ( .B1(n4270), .B2(n2857), .A(n3593), .ZN(n3594) );
  NOR2_X1 U4380 ( .A1(n3595), .A2(n3594), .ZN(n3749) );
  NAND2_X1 U4381 ( .A1(n3595), .A2(n3594), .ZN(n3748) );
  OAI22_X1 U4382 ( .A1(n3849), .A2(n3600), .B1(n4057), .B2(n3599), .ZN(n3596)
         );
  XNOR2_X1 U4383 ( .A(n3596), .B(n3602), .ZN(n3598) );
  OAI22_X1 U4384 ( .A1(n3849), .A2(n3601), .B1(n4057), .B2(n3600), .ZN(n3597)
         );
  XNOR2_X1 U4385 ( .A(n3598), .B(n3597), .ZN(n3628) );
  OAI22_X1 U4386 ( .A1(n4273), .A2(n3049), .B1(n3599), .B2(n4037), .ZN(n3605)
         );
  OAI22_X1 U4387 ( .A1(n4273), .A2(n3601), .B1(n3600), .B2(n4037), .ZN(n3603)
         );
  XNOR2_X1 U4388 ( .A(n3603), .B(n3602), .ZN(n3604) );
  XOR2_X1 U4389 ( .A(n3605), .B(n3604), .Z(n3606) );
  OAI22_X1 U4390 ( .A1(n3768), .A2(n4037), .B1(STATE_REG_SCAN_IN), .B2(n3607), 
        .ZN(n3609) );
  INV_X1 U4391 ( .A(n3949), .ZN(n4042) );
  OAI22_X1 U4392 ( .A1(n4042), .A2(n3755), .B1(n3776), .B2(n4035), .ZN(n3608)
         );
  AOI211_X1 U4393 ( .C1(n3753), .C2(n4072), .A(n3609), .B(n3608), .ZN(n3610)
         );
  OAI21_X1 U4394 ( .B1(n3611), .B2(n3759), .A(n3610), .ZN(U3217) );
  INV_X1 U4395 ( .A(n3612), .ZN(n3613) );
  OAI21_X1 U4396 ( .B1(n2077), .B2(n4037), .A(n3613), .ZN(n4034) );
  OR2_X1 U4397 ( .A1(n4034), .A2(n4404), .ZN(n3623) );
  INV_X1 U4398 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3621) );
  XNOR2_X1 U4399 ( .A(n3908), .B(n3615), .ZN(n4033) );
  XNOR2_X1 U4400 ( .A(n3616), .B(n3908), .ZN(n3617) );
  NAND2_X1 U4401 ( .A1(n3617), .A2(n2715), .ZN(n4047) );
  AOI22_X1 U4402 ( .A1(n4072), .A2(n4333), .B1(n4345), .B2(n3618), .ZN(n3619)
         );
  OAI211_X1 U4403 ( .C1(n4042), .C2(n4337), .A(n4047), .B(n3619), .ZN(n3620)
         );
  AOI21_X1 U4404 ( .B1(n4033), .B2(n4340), .A(n3620), .ZN(n3624) );
  MUX2_X1 U4405 ( .A(n3621), .B(n3624), .S(n4546), .Z(n3622) );
  NAND2_X1 U4406 ( .A1(n3623), .A2(n3622), .ZN(U3514) );
  MUX2_X1 U4407 ( .A(n3625), .B(n3624), .S(n4552), .Z(n3626) );
  OAI21_X1 U4408 ( .B1(n4343), .B2(n4034), .A(n3626), .ZN(U3546) );
  XNOR2_X1 U4409 ( .A(n3627), .B(n3628), .ZN(n3633) );
  OAI22_X1 U4410 ( .A1(n3768), .A2(n4057), .B1(STATE_REG_SCAN_IN), .B2(n4640), 
        .ZN(n3629) );
  AOI21_X1 U4411 ( .B1(n4270), .B2(n3753), .A(n3629), .ZN(n3630) );
  OAI21_X1 U4412 ( .B1(n3776), .B2(n4055), .A(n3630), .ZN(n3631) );
  AOI21_X1 U4413 ( .B1(n4061), .B2(n3772), .A(n3631), .ZN(n3632) );
  OAI21_X1 U4414 ( .B1(n3633), .B2(n3759), .A(n3632), .ZN(U3211) );
  NAND2_X1 U4415 ( .A1(n3636), .A2(n3635), .ZN(n3637) );
  XNOR2_X1 U4416 ( .A(n3634), .B(n3637), .ZN(n3645) );
  INV_X1 U4417 ( .A(n3638), .ZN(n3643) );
  NAND2_X1 U4418 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4475) );
  OAI21_X1 U4419 ( .B1(n3755), .B2(n4350), .A(n4475), .ZN(n3642) );
  OAI22_X1 U4420 ( .A1(n3770), .A2(n3640), .B1(n3768), .B2(n3639), .ZN(n3641)
         );
  AOI211_X1 U4421 ( .C1(n3643), .C2(n3757), .A(n3642), .B(n3641), .ZN(n3644)
         );
  OAI21_X1 U4422 ( .B1(n3645), .B2(n3759), .A(n3644), .ZN(U3212) );
  NAND2_X1 U4423 ( .A1(n3646), .A2(n3718), .ZN(n3667) );
  OAI21_X1 U4424 ( .B1(n3727), .B2(n3650), .A(n3649), .ZN(n3652) );
  NAND3_X1 U4425 ( .A1(n3652), .A2(n3764), .A3(n3651), .ZN(n3657) );
  NOR2_X1 U4426 ( .A1(n4611), .A2(STATE_REG_SCAN_IN), .ZN(n3655) );
  OAI22_X1 U4427 ( .A1(n3653), .A2(n3755), .B1(n3768), .B2(n4132), .ZN(n3654)
         );
  AOI211_X1 U4428 ( .C1(n3753), .C2(n4162), .A(n3655), .B(n3654), .ZN(n3656)
         );
  OAI211_X1 U4429 ( .C1(n3776), .C2(n4134), .A(n3657), .B(n3656), .ZN(U3213)
         );
  XOR2_X1 U4430 ( .A(n3659), .B(n3658), .Z(n3663) );
  NAND2_X1 U4431 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4010) );
  OAI21_X1 U4432 ( .B1(n3668), .B2(n3755), .A(n4010), .ZN(n3661) );
  OAI22_X1 U4433 ( .A1(n3770), .A2(n4338), .B1(n3768), .B2(n4209), .ZN(n3660)
         );
  AOI211_X1 U4434 ( .C1(n4211), .C2(n3757), .A(n3661), .B(n3660), .ZN(n3662)
         );
  OAI21_X1 U4435 ( .B1(n3663), .B2(n3759), .A(n3662), .ZN(U3216) );
  XNOR2_X1 U4436 ( .A(n3665), .B(n3664), .ZN(n3666) );
  XNOR2_X1 U4437 ( .A(n3667), .B(n3666), .ZN(n3673) );
  OAI22_X1 U4438 ( .A1(n3770), .A2(n3668), .B1(n3768), .B2(n4167), .ZN(n3671)
         );
  OAI22_X1 U4439 ( .A1(n4315), .A2(n3755), .B1(STATE_REG_SCAN_IN), .B2(n3669), 
        .ZN(n3670) );
  AOI211_X1 U4440 ( .C1(n4163), .C2(n3757), .A(n3671), .B(n3670), .ZN(n3672)
         );
  OAI21_X1 U4441 ( .B1(n3673), .B2(n3759), .A(n3672), .ZN(U3220) );
  NAND2_X1 U4442 ( .A1(n3675), .A2(n3674), .ZN(n3677) );
  XOR2_X1 U4443 ( .A(n3677), .B(n3676), .Z(n3682) );
  NOR2_X1 U4444 ( .A1(n4093), .A2(n3776), .ZN(n3680) );
  AOI22_X1 U4445 ( .A1(n4283), .A2(n3753), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3678) );
  OAI21_X1 U4446 ( .B1(n3768), .B2(n4091), .A(n3678), .ZN(n3679) );
  AOI211_X1 U4447 ( .C1(n3772), .C2(n4270), .A(n3680), .B(n3679), .ZN(n3681)
         );
  OAI21_X1 U4448 ( .B1(n3682), .B2(n3759), .A(n3681), .ZN(U3222) );
  INV_X1 U4449 ( .A(n3683), .ZN(n3686) );
  AND2_X1 U4450 ( .A1(n3685), .A2(n3684), .ZN(n3761) );
  OAI21_X1 U4451 ( .B1(n3686), .B2(n3762), .A(n3761), .ZN(n3687) );
  XOR2_X1 U4452 ( .A(n3688), .B(n3687), .Z(n3694) );
  INV_X1 U4453 ( .A(n4347), .ZN(n3742) );
  NAND2_X1 U4454 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4494) );
  OAI21_X1 U4455 ( .B1(n3755), .B2(n3742), .A(n4494), .ZN(n3691) );
  OAI22_X1 U4456 ( .A1(n3770), .A2(n4350), .B1(n3768), .B2(n3689), .ZN(n3690)
         );
  AOI211_X1 U4457 ( .C1(n3692), .C2(n3757), .A(n3691), .B(n3690), .ZN(n3693)
         );
  OAI21_X1 U4458 ( .B1(n3694), .B2(n3759), .A(n3693), .ZN(U3223) );
  XNOR2_X1 U4459 ( .A(n3697), .B(n3696), .ZN(n3698) );
  XNOR2_X1 U4460 ( .A(n3695), .B(n3698), .ZN(n3705) );
  NAND2_X1 U4461 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n3997) );
  OAI21_X1 U4462 ( .B1(n3755), .B2(n4338), .A(n3997), .ZN(n3702) );
  OAI22_X1 U4463 ( .A1(n3770), .A2(n3700), .B1(n3768), .B2(n3699), .ZN(n3701)
         );
  AOI211_X1 U4464 ( .C1(n3703), .C2(n3757), .A(n3702), .B(n3701), .ZN(n3704)
         );
  OAI21_X1 U4465 ( .B1(n3705), .B2(n3759), .A(n3704), .ZN(U3225) );
  NAND2_X1 U4466 ( .A1(n3706), .A2(n3707), .ZN(n3708) );
  XOR2_X1 U4467 ( .A(n3709), .B(n3708), .Z(n3714) );
  NOR2_X1 U4468 ( .A1(n4110), .A2(n3776), .ZN(n3712) );
  AOI22_X1 U4469 ( .A1(n4292), .A2(n3753), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3710) );
  OAI21_X1 U4470 ( .B1(n3768), .B2(n4107), .A(n3710), .ZN(n3711) );
  AOI211_X1 U4471 ( .C1(n3772), .C2(n3950), .A(n3712), .B(n3711), .ZN(n3713)
         );
  OAI21_X1 U4472 ( .B1(n3714), .B2(n3759), .A(n3713), .ZN(U3226) );
  INV_X1 U4473 ( .A(n3646), .ZN(n3719) );
  AOI21_X1 U4474 ( .B1(n3718), .B2(n3716), .A(n3715), .ZN(n3717) );
  AOI21_X1 U4475 ( .B1(n3719), .B2(n3718), .A(n3717), .ZN(n3724) );
  INV_X1 U4476 ( .A(n4191), .ZN(n3722) );
  OAI22_X1 U4477 ( .A1(n3770), .A2(n4224), .B1(STATE_REG_SCAN_IN), .B2(n4574), 
        .ZN(n3721) );
  INV_X1 U4478 ( .A(n4141), .ZN(n4181) );
  OAI22_X1 U4479 ( .A1(n4181), .A2(n3755), .B1(n3768), .B2(n4188), .ZN(n3720)
         );
  AOI211_X1 U4480 ( .C1(n3722), .C2(n3757), .A(n3721), .B(n3720), .ZN(n3723)
         );
  OAI21_X1 U4481 ( .B1(n3724), .B2(n3759), .A(n3723), .ZN(U3230) );
  NAND2_X1 U4482 ( .A1(n3726), .A2(n3725), .ZN(n3728) );
  AOI21_X1 U4483 ( .B1(n3729), .B2(n3728), .A(n3727), .ZN(n3735) );
  INV_X1 U4484 ( .A(n4151), .ZN(n3733) );
  OAI22_X1 U4485 ( .A1(n4181), .A2(n3770), .B1(n3768), .B2(n4149), .ZN(n3732)
         );
  OAI22_X1 U4486 ( .A1(n4112), .A2(n3755), .B1(STATE_REG_SCAN_IN), .B2(n3730), 
        .ZN(n3731) );
  AOI211_X1 U4487 ( .C1(n3733), .C2(n3757), .A(n3732), .B(n3731), .ZN(n3734)
         );
  OAI21_X1 U4488 ( .B1(n3735), .B2(n3759), .A(n3734), .ZN(U3232) );
  INV_X1 U4489 ( .A(n3737), .ZN(n3739) );
  NAND2_X1 U4490 ( .A1(n3739), .A2(n3738), .ZN(n3740) );
  XNOR2_X1 U4491 ( .A(n3736), .B(n3740), .ZN(n3741) );
  NAND2_X1 U4492 ( .A1(n3741), .A2(n3764), .ZN(n3746) );
  OAI22_X1 U4493 ( .A1(n3770), .A2(n3742), .B1(n3768), .B2(n4219), .ZN(n3743)
         );
  AOI211_X1 U4494 ( .C1(n3772), .C2(n4179), .A(n3744), .B(n3743), .ZN(n3745)
         );
  OAI211_X1 U4495 ( .C1(n3776), .C2(n4228), .A(n3746), .B(n3745), .ZN(U3235)
         );
  NOR2_X1 U4496 ( .A1(n3749), .A2(n2182), .ZN(n3750) );
  XNOR2_X1 U4497 ( .A(n3747), .B(n3750), .ZN(n3760) );
  OAI22_X1 U4498 ( .A1(n3768), .A2(n4076), .B1(STATE_REG_SCAN_IN), .B2(n3751), 
        .ZN(n3752) );
  AOI21_X1 U4499 ( .B1(n3950), .B2(n3753), .A(n3752), .ZN(n3754) );
  OAI21_X1 U4500 ( .B1(n3849), .B2(n3755), .A(n3754), .ZN(n3756) );
  AOI21_X1 U4501 ( .B1(n4077), .B2(n3757), .A(n3756), .ZN(n3758) );
  OAI21_X1 U4502 ( .B1(n3760), .B2(n3759), .A(n3758), .ZN(U3237) );
  NAND2_X1 U4503 ( .A1(n3683), .A2(n3761), .ZN(n3763) );
  XNOR2_X1 U4504 ( .A(n3763), .B(n3762), .ZN(n3765) );
  NAND2_X1 U4505 ( .A1(n3765), .A2(n3764), .ZN(n3774) );
  NOR2_X1 U4506 ( .A1(n3766), .A2(STATE_REG_SCAN_IN), .ZN(n4488) );
  OAI22_X1 U4507 ( .A1(n3770), .A2(n3769), .B1(n3768), .B2(n3767), .ZN(n3771)
         );
  AOI211_X1 U4508 ( .C1(n3772), .C2(n4334), .A(n4488), .B(n3771), .ZN(n3773)
         );
  OAI211_X1 U4509 ( .C1(n3776), .C2(n3775), .A(n3774), .B(n3773), .ZN(U3238)
         );
  INV_X1 U4510 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4260) );
  NAND2_X1 U4511 ( .A1(n2455), .A2(REG2_REG_31__SCAN_IN), .ZN(n3778) );
  NAND2_X1 U4512 ( .A1(n2470), .A2(REG0_REG_31__SCAN_IN), .ZN(n3777) );
  OAI211_X1 U4513 ( .C1(n2471), .C2(n4260), .A(n3778), .B(n3777), .ZN(n4017)
         );
  NAND2_X1 U4514 ( .A1(n3779), .A2(DATAI_31_), .ZN(n4016) );
  NAND2_X1 U4515 ( .A1(n4017), .A2(n4016), .ZN(n3853) );
  INV_X1 U4516 ( .A(n3853), .ZN(n3861) );
  INV_X1 U4517 ( .A(DATAI_30_), .ZN(n4555) );
  NOR2_X1 U4518 ( .A1(n3780), .A2(n4555), .ZN(n4267) );
  NOR2_X1 U4519 ( .A1(n3852), .A2(n4267), .ZN(n3934) );
  INV_X1 U4520 ( .A(n3934), .ZN(n3782) );
  OR2_X1 U4521 ( .A1(n4017), .A2(n4016), .ZN(n3781) );
  NAND2_X1 U4522 ( .A1(n3782), .A2(n3781), .ZN(n3886) );
  INV_X1 U4523 ( .A(n3886), .ZN(n3860) );
  INV_X1 U4524 ( .A(n4024), .ZN(n3784) );
  OAI21_X1 U4525 ( .B1(n4042), .B2(n3784), .A(n3783), .ZN(n3927) );
  NAND3_X1 U4526 ( .A1(n3787), .A2(n2700), .A3(n3786), .ZN(n3912) );
  INV_X1 U4527 ( .A(n3912), .ZN(n3841) );
  NAND2_X1 U4528 ( .A1(n3790), .A2(n3789), .ZN(n3797) );
  NAND2_X1 U4529 ( .A1(n3797), .A2(n3792), .ZN(n3910) );
  NAND2_X1 U4530 ( .A1(n3792), .A2(n3791), .ZN(n3911) );
  INV_X1 U4531 ( .A(n3911), .ZN(n3793) );
  OAI211_X1 U4532 ( .C1(n3796), .C2(n3795), .A(n3794), .B(n3793), .ZN(n3837)
         );
  INV_X1 U4533 ( .A(n3797), .ZN(n3827) );
  INV_X1 U4534 ( .A(n3798), .ZN(n3816) );
  OAI211_X1 U4535 ( .C1(n3937), .C2(n2692), .A(n3801), .B(n3800), .ZN(n3802)
         );
  NAND3_X1 U4536 ( .A1(n3804), .A2(n3803), .A3(n3802), .ZN(n3805) );
  NAND3_X1 U4537 ( .A1(n3807), .A2(n3806), .A3(n3805), .ZN(n3808) );
  NAND3_X1 U4538 ( .A1(n3810), .A2(n3809), .A3(n3808), .ZN(n3811) );
  NAND4_X1 U4539 ( .A1(n3814), .A2(n3813), .A3(n3812), .A4(n3811), .ZN(n3815)
         );
  NAND3_X1 U4540 ( .A1(n3880), .A2(n3816), .A3(n3815), .ZN(n3817) );
  NAND3_X1 U4541 ( .A1(n3821), .A2(n3822), .A3(n3817), .ZN(n3818) );
  NAND3_X1 U4542 ( .A1(n3820), .A2(n3819), .A3(n3818), .ZN(n3826) );
  NOR4_X1 U4543 ( .A1(n2097), .A2(n2093), .A3(n3824), .A4(n3823), .ZN(n3825)
         );
  AOI22_X1 U4544 ( .A1(n3827), .A2(n3826), .B1(n3825), .B2(n3910), .ZN(n3830)
         );
  INV_X1 U4545 ( .A(n3910), .ZN(n3829) );
  OAI22_X1 U4546 ( .A1(n3831), .A2(n3830), .B1(n3829), .B2(n3828), .ZN(n3832)
         );
  AND4_X1 U4547 ( .A1(n3835), .A2(n3834), .A3(n3833), .A4(n3832), .ZN(n3836)
         );
  AOI21_X1 U4548 ( .B1(n3910), .B2(n3837), .A(n3836), .ZN(n3838) );
  OAI21_X1 U4549 ( .B1(n2089), .B2(n3838), .A(n3913), .ZN(n3840) );
  INV_X1 U4550 ( .A(n3915), .ZN(n3839) );
  AOI21_X1 U4551 ( .B1(n3841), .B2(n3840), .A(n3839), .ZN(n3842) );
  OAI21_X1 U4552 ( .B1(n4122), .B2(n3842), .A(n3916), .ZN(n3843) );
  INV_X1 U4553 ( .A(n3843), .ZN(n3846) );
  INV_X1 U4554 ( .A(n3869), .ZN(n3844) );
  NOR2_X1 U4555 ( .A1(n3844), .A2(n3866), .ZN(n3920) );
  OAI211_X1 U4556 ( .C1(n3846), .C2(n3845), .A(n2710), .B(n3920), .ZN(n3847)
         );
  OAI211_X1 U4557 ( .C1(n3849), .C2(n4269), .A(n3848), .B(n3847), .ZN(n3858)
         );
  NAND2_X1 U4558 ( .A1(n3851), .A2(n3850), .ZN(n3924) );
  INV_X1 U4559 ( .A(n3924), .ZN(n3856) );
  NAND2_X1 U4560 ( .A1(n3852), .A2(n4267), .ZN(n3854) );
  AND2_X1 U4561 ( .A1(n3854), .A2(n3853), .ZN(n3884) );
  OAI21_X1 U4562 ( .B1(n3949), .B2(n4024), .A(n3884), .ZN(n3922) );
  INV_X1 U4563 ( .A(n3922), .ZN(n3855) );
  OAI21_X1 U4564 ( .B1(n3856), .B2(n3927), .A(n3855), .ZN(n3928) );
  INV_X1 U4565 ( .A(n3928), .ZN(n3857) );
  OAI21_X1 U4566 ( .B1(n3927), .B2(n3858), .A(n3857), .ZN(n3859) );
  OAI21_X1 U4567 ( .B1(n3861), .B2(n3860), .A(n3859), .ZN(n3941) );
  INV_X1 U4568 ( .A(n4051), .ZN(n3863) );
  NOR2_X1 U4569 ( .A1(n3863), .A2(n3862), .ZN(n3909) );
  XNOR2_X1 U4570 ( .A(n4270), .B(n3864), .ZN(n4068) );
  INV_X1 U4571 ( .A(n4082), .ZN(n3865) );
  OR2_X1 U4572 ( .A1(n3866), .A2(n3865), .ZN(n4102) );
  INV_X1 U4573 ( .A(n4102), .ZN(n4104) );
  INV_X1 U4574 ( .A(n3867), .ZN(n4123) );
  NOR2_X1 U4575 ( .A1(n4123), .A2(n4122), .ZN(n4157) );
  XNOR2_X1 U4576 ( .A(n4312), .B(n4178), .ZN(n4176) );
  AND2_X1 U4577 ( .A1(n4146), .A2(n4176), .ZN(n3904) );
  NAND2_X1 U4578 ( .A1(n3869), .A2(n3868), .ZN(n4126) );
  NAND2_X1 U4579 ( .A1(n3871), .A2(n3870), .ZN(n4202) );
  OR2_X1 U4580 ( .A1(n3873), .A2(n3872), .ZN(n3874) );
  NOR2_X1 U4581 ( .A1(n4202), .A2(n3874), .ZN(n3901) );
  NAND4_X1 U4582 ( .A1(n3878), .A2(n2699), .A3(n3877), .A4(n3876), .ZN(n3883)
         );
  NAND4_X1 U4583 ( .A1(n3881), .A2(n3880), .A3(n3879), .A4(n4531), .ZN(n3882)
         );
  NOR2_X1 U4584 ( .A1(n3883), .A2(n3882), .ZN(n3900) );
  INV_X1 U4585 ( .A(n3884), .ZN(n3885) );
  NOR2_X1 U4586 ( .A1(n3886), .A2(n3885), .ZN(n3887) );
  AND2_X1 U4587 ( .A1(n4238), .A2(n3887), .ZN(n3899) );
  NAND4_X1 U4588 ( .A1(n3891), .A2(n3890), .A3(n3889), .A4(n3888), .ZN(n3897)
         );
  NAND4_X1 U4589 ( .A1(n3895), .A2(n3894), .A3(n3893), .A4(n3892), .ZN(n3896)
         );
  NOR2_X1 U4590 ( .A1(n3897), .A2(n3896), .ZN(n3898) );
  NAND4_X1 U4591 ( .A1(n3901), .A2(n3900), .A3(n3899), .A4(n3898), .ZN(n3902)
         );
  NOR2_X1 U4592 ( .A1(n4126), .A2(n3902), .ZN(n3903) );
  NAND4_X1 U4593 ( .A1(n4104), .A2(n4157), .A3(n3904), .A4(n3903), .ZN(n3906)
         );
  NAND2_X1 U4594 ( .A1(n4065), .A2(n3905), .ZN(n4087) );
  NOR2_X1 U4595 ( .A1(n3906), .A2(n4087), .ZN(n3907) );
  NAND4_X1 U4596 ( .A1(n3909), .A2(n3908), .A3(n4068), .A4(n3907), .ZN(n3939)
         );
  OAI21_X1 U4597 ( .B1(n3335), .B2(n3911), .A(n3910), .ZN(n3914) );
  AOI211_X1 U4598 ( .C1(n3914), .C2(n3913), .A(n2089), .B(n3912), .ZN(n3919)
         );
  NAND2_X1 U4599 ( .A1(n3916), .A2(n3915), .ZN(n3918) );
  OAI21_X1 U4600 ( .B1(n3919), .B2(n3918), .A(n3917), .ZN(n3921) );
  AOI21_X1 U4601 ( .B1(n3921), .B2(n3920), .A(n4066), .ZN(n3925) );
  NOR4_X1 U4602 ( .A1(n3925), .A2(n3924), .A3(n3923), .A4(n3922), .ZN(n3932)
         );
  NOR2_X1 U4603 ( .A1(n3927), .A2(n3926), .ZN(n3929) );
  AOI21_X1 U4604 ( .B1(n4051), .B2(n3929), .A(n3928), .ZN(n3931) );
  INV_X1 U4605 ( .A(n4267), .ZN(n3930) );
  OAI22_X1 U4606 ( .A1(n3932), .A2(n3931), .B1(n3930), .B2(n4017), .ZN(n3936)
         );
  INV_X1 U4607 ( .A(n4017), .ZN(n3933) );
  INV_X1 U4608 ( .A(n4016), .ZN(n4018) );
  OAI21_X1 U4609 ( .B1(n3934), .B2(n3933), .A(n4018), .ZN(n3935) );
  NAND2_X1 U4610 ( .A1(n3936), .A2(n3935), .ZN(n3938) );
  MUX2_X1 U4611 ( .A(n3939), .B(n3938), .S(n3937), .Z(n3940) );
  MUX2_X1 U4612 ( .A(n3941), .B(n3940), .S(n4410), .Z(n3942) );
  XNOR2_X1 U4613 ( .A(n3942), .B(n4011), .ZN(n3948) );
  NAND2_X1 U4614 ( .A1(n3944), .A2(n3943), .ZN(n3945) );
  OAI211_X1 U4615 ( .C1(n4409), .C2(n3947), .A(n3945), .B(B_REG_SCAN_IN), .ZN(
        n3946) );
  OAI21_X1 U4616 ( .B1(n3948), .B2(n3947), .A(n3946), .ZN(U3239) );
  MUX2_X1 U4617 ( .A(DATAO_REG_31__SCAN_IN), .B(n4017), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4618 ( .A(DATAO_REG_29__SCAN_IN), .B(n3949), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4619 ( .A(DATAO_REG_28__SCAN_IN), .B(n4061), .S(n3951), .Z(U3578)
         );
  MUX2_X1 U4620 ( .A(DATAO_REG_27__SCAN_IN), .B(n4072), .S(n3951), .Z(U3577)
         );
  MUX2_X1 U4621 ( .A(DATAO_REG_26__SCAN_IN), .B(n4270), .S(n3951), .Z(U3576)
         );
  MUX2_X1 U4622 ( .A(DATAO_REG_25__SCAN_IN), .B(n3950), .S(n3951), .Z(U3575)
         );
  MUX2_X1 U4623 ( .A(DATAO_REG_24__SCAN_IN), .B(n4283), .S(n3951), .Z(U3574)
         );
  MUX2_X1 U4624 ( .A(DATAO_REG_23__SCAN_IN), .B(n4292), .S(n3951), .Z(U3573)
         );
  MUX2_X1 U4625 ( .A(DATAO_REG_22__SCAN_IN), .B(n4162), .S(n3951), .Z(U3572)
         );
  MUX2_X1 U4626 ( .A(DATAO_REG_21__SCAN_IN), .B(n4141), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4627 ( .A(n4312), .B(DATAO_REG_20__SCAN_IN), .S(n3965), .Z(U3570)
         );
  MUX2_X1 U4628 ( .A(n4179), .B(DATAO_REG_19__SCAN_IN), .S(n3965), .Z(U3569)
         );
  MUX2_X1 U4629 ( .A(DATAO_REG_18__SCAN_IN), .B(n3952), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4630 ( .A(n4347), .B(DATAO_REG_17__SCAN_IN), .S(n3965), .Z(U3567)
         );
  MUX2_X1 U4631 ( .A(DATAO_REG_16__SCAN_IN), .B(n4334), .S(n3951), .Z(U3566)
         );
  MUX2_X1 U4632 ( .A(n3953), .B(DATAO_REG_15__SCAN_IN), .S(n3965), .Z(U3565)
         );
  MUX2_X1 U4633 ( .A(DATAO_REG_14__SCAN_IN), .B(n3954), .S(n3951), .Z(U3564)
         );
  MUX2_X1 U4634 ( .A(n3955), .B(DATAO_REG_13__SCAN_IN), .S(n3965), .Z(U3563)
         );
  MUX2_X1 U4635 ( .A(n3956), .B(DATAO_REG_12__SCAN_IN), .S(n3965), .Z(U3562)
         );
  MUX2_X1 U4636 ( .A(DATAO_REG_11__SCAN_IN), .B(n3957), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4637 ( .A(n3958), .B(DATAO_REG_10__SCAN_IN), .S(n3965), .Z(U3560)
         );
  MUX2_X1 U4638 ( .A(n3959), .B(DATAO_REG_9__SCAN_IN), .S(n3965), .Z(U3559) );
  MUX2_X1 U4639 ( .A(DATAO_REG_8__SCAN_IN), .B(n3960), .S(n3951), .Z(U3558) );
  MUX2_X1 U4640 ( .A(DATAO_REG_7__SCAN_IN), .B(n3961), .S(n3951), .Z(U3557) );
  MUX2_X1 U4641 ( .A(n3962), .B(DATAO_REG_6__SCAN_IN), .S(n3965), .Z(U3556) );
  MUX2_X1 U4642 ( .A(DATAO_REG_5__SCAN_IN), .B(n2694), .S(n3951), .Z(U3555) );
  MUX2_X1 U4643 ( .A(DATAO_REG_4__SCAN_IN), .B(n3963), .S(U4043), .Z(U3554) );
  MUX2_X1 U4644 ( .A(n4253), .B(DATAO_REG_3__SCAN_IN), .S(n3965), .Z(U3553) );
  MUX2_X1 U4645 ( .A(DATAO_REG_2__SCAN_IN), .B(n3964), .S(U4043), .Z(U3552) );
  MUX2_X1 U4646 ( .A(DATAO_REG_1__SCAN_IN), .B(n4247), .S(U4043), .Z(U3551) );
  MUX2_X1 U4647 ( .A(n3966), .B(DATAO_REG_0__SCAN_IN), .S(n3965), .Z(U3550) );
  INV_X1 U4648 ( .A(n4507), .ZN(n3979) );
  NAND2_X1 U4649 ( .A1(n3979), .A2(n4416), .ZN(n3978) );
  OAI211_X1 U4650 ( .C1(n3969), .C2(n3968), .A(n4502), .B(n3967), .ZN(n3977)
         );
  MUX2_X1 U4651 ( .A(n2254), .B(REG2_REG_1__SCAN_IN), .S(n3971), .Z(n3974) );
  INV_X1 U4652 ( .A(n3972), .ZN(n3973) );
  OAI211_X1 U4653 ( .C1(n2256), .C2(n3974), .A(n4466), .B(n3973), .ZN(n3976)
         );
  AOI22_X1 U4654 ( .A1(n4501), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3975) );
  NAND4_X1 U4655 ( .A1(n3978), .A2(n3977), .A3(n3976), .A4(n3975), .ZN(U3241)
         );
  NAND2_X1 U4656 ( .A1(n3979), .A2(n4414), .ZN(n3987) );
  OAI211_X1 U4657 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3981), .A(n4502), .B(n3980), 
        .ZN(n3986) );
  AOI22_X1 U4658 ( .A1(n4501), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3985) );
  XNOR2_X1 U4659 ( .A(n3982), .B(REG2_REG_3__SCAN_IN), .ZN(n3983) );
  NAND2_X1 U4660 ( .A1(n4466), .A2(n3983), .ZN(n3984) );
  NAND4_X1 U4661 ( .A1(n3987), .A2(n3986), .A3(n3985), .A4(n3984), .ZN(U3243)
         );
  AND2_X1 U4662 ( .A1(n3989), .A2(n3988), .ZN(n3991) );
  OAI21_X1 U4663 ( .B1(n3991), .B2(n3990), .A(n4502), .ZN(n4000) );
  AOI221_X1 U4664 ( .B1(n3994), .B2(n3993), .C1(n3992), .C2(n3993), .A(n4495), 
        .ZN(n3995) );
  INV_X1 U4665 ( .A(n3995), .ZN(n3996) );
  NAND2_X1 U4666 ( .A1(n3997), .A2(n3996), .ZN(n3998) );
  AOI21_X1 U4667 ( .B1(n4501), .B2(ADDR_REG_17__SCAN_IN), .A(n3998), .ZN(n3999) );
  OAI211_X1 U4668 ( .C1(n4507), .C2(n4001), .A(n4000), .B(n3999), .ZN(U3257)
         );
  MUX2_X1 U4669 ( .A(REG2_REG_19__SCAN_IN), .B(n2599), .S(n4227), .Z(n4004) );
  MUX2_X1 U4670 ( .A(n4327), .B(REG1_REG_19__SCAN_IN), .S(n4227), .Z(n4007) );
  XNOR2_X1 U4671 ( .A(n4008), .B(n4007), .ZN(n4013) );
  NAND2_X1 U4672 ( .A1(n4501), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4009) );
  OAI211_X1 U4673 ( .C1(n4507), .C2(n4011), .A(n4010), .B(n4009), .ZN(n4012)
         );
  AOI21_X1 U4674 ( .B1(n4013), .B2(n4502), .A(n4012), .ZN(n4014) );
  OAI21_X1 U4675 ( .B1(n4015), .B2(n4495), .A(n4014), .ZN(U3259) );
  XNOR2_X1 U4676 ( .A(n4263), .B(n4016), .ZN(n4360) );
  NAND2_X1 U4677 ( .A1(n4017), .A2(n2212), .ZN(n4265) );
  NAND2_X1 U4678 ( .A1(n4345), .A2(n4018), .ZN(n4019) );
  NAND2_X1 U4679 ( .A1(n4265), .A2(n4019), .ZN(n4357) );
  NAND2_X1 U4680 ( .A1(n4215), .A2(n4357), .ZN(n4021) );
  NAND2_X1 U4681 ( .A1(n4520), .A2(REG2_REG_31__SCAN_IN), .ZN(n4020) );
  OAI211_X1 U4682 ( .C1(n4360), .C2(n4213), .A(n4021), .B(n4020), .ZN(U3260)
         );
  INV_X1 U4683 ( .A(n4022), .ZN(n4032) );
  INV_X1 U4684 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4023) );
  OAI22_X1 U4685 ( .A1(n4166), .A2(n4024), .B1(n4023), .B2(n4215), .ZN(n4025)
         );
  AOI21_X1 U4686 ( .B1(n4061), .B2(n4248), .A(n4025), .ZN(n4031) );
  OAI22_X1 U4687 ( .A1(n4027), .A2(n4213), .B1(n4026), .B2(n4508), .ZN(n4028)
         );
  OAI21_X1 U4688 ( .B1(n4029), .B2(n4028), .A(n4215), .ZN(n4030) );
  OAI211_X1 U4689 ( .C1(n4032), .C2(n4239), .A(n4031), .B(n4030), .ZN(U3354)
         );
  NAND2_X1 U4690 ( .A1(n4033), .A2(n4159), .ZN(n4046) );
  INV_X1 U4691 ( .A(n4034), .ZN(n4044) );
  INV_X1 U4692 ( .A(n4035), .ZN(n4039) );
  INV_X1 U4693 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4036) );
  OAI22_X1 U4694 ( .A1(n4166), .A2(n4037), .B1(n4036), .B2(n4511), .ZN(n4038)
         );
  AOI21_X1 U4695 ( .B1(n4039), .B2(n4250), .A(n4038), .ZN(n4041) );
  NAND2_X1 U4696 ( .A1(n4072), .A2(n4248), .ZN(n4040) );
  OAI211_X1 U4697 ( .C1(n4042), .C2(n4113), .A(n4041), .B(n4040), .ZN(n4043)
         );
  AOI21_X1 U4698 ( .B1(n4044), .B2(n4514), .A(n4043), .ZN(n4045) );
  OAI211_X1 U4699 ( .C1(n4520), .C2(n4047), .A(n4046), .B(n4045), .ZN(U3262)
         );
  OAI21_X1 U4700 ( .B1(n4051), .B2(n4049), .A(n4048), .ZN(n4050) );
  NAND2_X1 U4701 ( .A1(n4050), .A2(n2715), .ZN(n4272) );
  XNOR2_X1 U4702 ( .A(n4052), .B(n4051), .ZN(n4275) );
  NAND2_X1 U4703 ( .A1(n4275), .A2(n4159), .ZN(n4063) );
  NAND2_X1 U4704 ( .A1(n4270), .A2(n4248), .ZN(n4054) );
  AOI22_X1 U4705 ( .A1(n4252), .A2(n4269), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4419), .ZN(n4053) );
  OAI211_X1 U4706 ( .C1(n4508), .C2(n4055), .A(n4054), .B(n4053), .ZN(n4060)
         );
  INV_X1 U4707 ( .A(n4075), .ZN(n4058) );
  OAI21_X1 U4708 ( .B1(n4058), .B2(n4057), .A(n4056), .ZN(n4367) );
  NOR2_X1 U4709 ( .A1(n4367), .A2(n4213), .ZN(n4059) );
  AOI211_X1 U4710 ( .C1(n4254), .C2(n4061), .A(n4060), .B(n4059), .ZN(n4062)
         );
  OAI211_X1 U4711 ( .C1(n4520), .C2(n4272), .A(n4063), .B(n4062), .ZN(U3263)
         );
  XNOR2_X1 U4712 ( .A(n4064), .B(n4068), .ZN(n4279) );
  INV_X1 U4713 ( .A(n4279), .ZN(n4081) );
  OAI21_X1 U4714 ( .B1(n4067), .B2(n4066), .A(n4065), .ZN(n4070) );
  INV_X1 U4715 ( .A(n4068), .ZN(n4069) );
  XNOR2_X1 U4716 ( .A(n4070), .B(n4069), .ZN(n4074) );
  OAI22_X1 U4717 ( .A1(n4295), .A2(n4349), .B1(n4076), .B2(n4203), .ZN(n4071)
         );
  AOI21_X1 U4718 ( .B1(n4072), .B2(n4346), .A(n4071), .ZN(n4073) );
  OAI21_X1 U4719 ( .B1(n4074), .B2(n4206), .A(n4073), .ZN(n4278) );
  OAI21_X1 U4720 ( .B1(n4088), .B2(n4076), .A(n4075), .ZN(n4371) );
  AOI22_X1 U4721 ( .A1(n4077), .A2(n4250), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4419), .ZN(n4078) );
  OAI21_X1 U4722 ( .B1(n4371), .B2(n4213), .A(n4078), .ZN(n4079) );
  AOI21_X1 U4723 ( .B1(n4278), .B2(n4215), .A(n4079), .ZN(n4080) );
  OAI21_X1 U4724 ( .B1(n4081), .B2(n4239), .A(n4080), .ZN(U3264) );
  NAND2_X1 U4725 ( .A1(n4083), .A2(n4082), .ZN(n4084) );
  XNOR2_X1 U4726 ( .A(n4084), .B(n4087), .ZN(n4085) );
  NAND2_X1 U4727 ( .A1(n4085), .A2(n2715), .ZN(n4285) );
  XOR2_X1 U4728 ( .A(n4087), .B(n4086), .Z(n4288) );
  NAND2_X1 U4729 ( .A1(n4288), .A2(n4159), .ZN(n4100) );
  INV_X1 U4730 ( .A(n4088), .ZN(n4090) );
  NAND2_X1 U4731 ( .A1(n4106), .A2(n4282), .ZN(n4089) );
  NAND2_X1 U4732 ( .A1(n4090), .A2(n4089), .ZN(n4375) );
  INV_X1 U4733 ( .A(n4375), .ZN(n4098) );
  NOR2_X1 U4734 ( .A1(n4166), .A2(n4091), .ZN(n4095) );
  INV_X1 U4735 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4092) );
  OAI22_X1 U4736 ( .A1(n4093), .A2(n4508), .B1(n4092), .B2(n4215), .ZN(n4094)
         );
  AOI211_X1 U4737 ( .C1(n4248), .C2(n4283), .A(n4095), .B(n4094), .ZN(n4096)
         );
  OAI21_X1 U4738 ( .B1(n4286), .B2(n4113), .A(n4096), .ZN(n4097) );
  AOI21_X1 U4739 ( .B1(n4098), .B2(n4514), .A(n4097), .ZN(n4099) );
  OAI211_X1 U4740 ( .C1(n4520), .C2(n4285), .A(n4100), .B(n4099), .ZN(U3265)
         );
  XOR2_X1 U4741 ( .A(n4102), .B(n4101), .Z(n4297) );
  XNOR2_X1 U4742 ( .A(n4103), .B(n4104), .ZN(n4105) );
  NAND2_X1 U4743 ( .A1(n4105), .A2(n2715), .ZN(n4294) );
  NOR2_X1 U4744 ( .A1(n4294), .A2(n4419), .ZN(n4118) );
  INV_X1 U4745 ( .A(n4131), .ZN(n4108) );
  OAI21_X1 U4746 ( .B1(n4108), .B2(n4107), .A(n4106), .ZN(n4379) );
  INV_X1 U4747 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4109) );
  OAI22_X1 U4748 ( .A1(n4110), .A2(n4508), .B1(n4109), .B2(n4215), .ZN(n4115)
         );
  OAI22_X1 U4749 ( .A1(n4295), .A2(n4113), .B1(n4112), .B2(n4111), .ZN(n4114)
         );
  AOI211_X1 U4750 ( .C1(n4291), .C2(n4252), .A(n4115), .B(n4114), .ZN(n4116)
         );
  OAI21_X1 U4751 ( .B1(n4379), .B2(n4213), .A(n4116), .ZN(n4117) );
  AOI211_X1 U4752 ( .C1(n4297), .C2(n4159), .A(n4118), .B(n4117), .ZN(n4119)
         );
  INV_X1 U4753 ( .A(n4119), .ZN(U3266) );
  XNOR2_X1 U4754 ( .A(n4120), .B(n4126), .ZN(n4301) );
  INV_X1 U4755 ( .A(n4301), .ZN(n4139) );
  INV_X1 U4756 ( .A(n4122), .ZN(n4124) );
  AOI21_X1 U4757 ( .B1(n4121), .B2(n4124), .A(n4123), .ZN(n4140) );
  OAI21_X1 U4758 ( .B1(n4140), .B2(n2128), .A(n4125), .ZN(n4127) );
  XNOR2_X1 U4759 ( .A(n4127), .B(n4126), .ZN(n4130) );
  OAI22_X1 U4760 ( .A1(n4315), .A2(n4349), .B1(n4203), .B2(n4132), .ZN(n4128)
         );
  AOI21_X1 U4761 ( .B1(n4346), .B2(n4283), .A(n4128), .ZN(n4129) );
  OAI21_X1 U4762 ( .B1(n4130), .B2(n4206), .A(n4129), .ZN(n4300) );
  INV_X1 U4763 ( .A(n4148), .ZN(n4133) );
  OAI21_X1 U4764 ( .B1(n4133), .B2(n4132), .A(n4131), .ZN(n4383) );
  INV_X1 U4765 ( .A(n4134), .ZN(n4135) );
  AOI22_X1 U4766 ( .A1(n4135), .A2(n4250), .B1(REG2_REG_23__SCAN_IN), .B2(
        n4419), .ZN(n4136) );
  OAI21_X1 U4767 ( .B1(n4383), .B2(n4213), .A(n4136), .ZN(n4137) );
  AOI21_X1 U4768 ( .B1(n4300), .B2(n4215), .A(n4137), .ZN(n4138) );
  OAI21_X1 U4769 ( .B1(n4139), .B2(n4239), .A(n4138), .ZN(U3267) );
  XNOR2_X1 U4770 ( .A(n4140), .B(n2128), .ZN(n4145) );
  NAND2_X1 U4771 ( .A1(n4292), .A2(n4346), .ZN(n4143) );
  NAND2_X1 U4772 ( .A1(n4141), .A2(n4333), .ZN(n4142) );
  OAI211_X1 U4773 ( .C1(n4203), .C2(n4149), .A(n4143), .B(n4142), .ZN(n4144)
         );
  AOI21_X1 U4774 ( .B1(n4145), .B2(n2715), .A(n4144), .ZN(n4307) );
  NAND2_X1 U4775 ( .A1(n4147), .A2(n4146), .ZN(n4304) );
  NAND3_X1 U4776 ( .A1(n2129), .A2(n4159), .A3(n4304), .ZN(n4155) );
  OAI21_X1 U4777 ( .B1(n4161), .B2(n4149), .A(n4148), .ZN(n4387) );
  INV_X1 U4778 ( .A(n4387), .ZN(n4153) );
  INV_X1 U4779 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4150) );
  OAI22_X1 U4780 ( .A1(n4151), .A2(n4508), .B1(n4150), .B2(n4511), .ZN(n4152)
         );
  AOI21_X1 U4781 ( .B1(n4153), .B2(n4514), .A(n4152), .ZN(n4154) );
  OAI211_X1 U4782 ( .C1(n4520), .C2(n4307), .A(n4155), .B(n4154), .ZN(U3268)
         );
  XNOR2_X1 U4783 ( .A(n4121), .B(n4157), .ZN(n4156) );
  NAND2_X1 U4784 ( .A1(n4156), .A2(n2715), .ZN(n4314) );
  XNOR2_X1 U4785 ( .A(n4158), .B(n4157), .ZN(n4317) );
  NAND2_X1 U4786 ( .A1(n4317), .A2(n4159), .ZN(n4171) );
  NOR2_X1 U4787 ( .A1(n4186), .A2(n4167), .ZN(n4160) );
  OR2_X1 U4788 ( .A1(n4161), .A2(n4160), .ZN(n4391) );
  INV_X1 U4789 ( .A(n4391), .ZN(n4169) );
  AOI22_X1 U4790 ( .A1(n4162), .A2(n4254), .B1(n4248), .B2(n4312), .ZN(n4165)
         );
  AOI22_X1 U4791 ( .A1(n4163), .A2(n4250), .B1(n4520), .B2(
        REG2_REG_21__SCAN_IN), .ZN(n4164) );
  OAI211_X1 U4792 ( .C1(n4167), .C2(n4166), .A(n4165), .B(n4164), .ZN(n4168)
         );
  AOI21_X1 U4793 ( .B1(n4169), .B2(n4514), .A(n4168), .ZN(n4170) );
  OAI211_X1 U4794 ( .C1(n4520), .C2(n4314), .A(n4171), .B(n4170), .ZN(U3269)
         );
  XNOR2_X1 U4795 ( .A(n4172), .B(n4176), .ZN(n4320) );
  INV_X1 U4796 ( .A(n4173), .ZN(n4174) );
  NAND2_X1 U4797 ( .A1(n4175), .A2(n4174), .ZN(n4177) );
  XNOR2_X1 U4798 ( .A(n4177), .B(n4176), .ZN(n4183) );
  AOI22_X1 U4799 ( .A1(n4179), .A2(n4333), .B1(n4178), .B2(n4345), .ZN(n4180)
         );
  OAI21_X1 U4800 ( .B1(n4181), .B2(n4337), .A(n4180), .ZN(n4182) );
  AOI21_X1 U4801 ( .B1(n4183), .B2(n2715), .A(n4182), .ZN(n4184) );
  OAI21_X1 U4802 ( .B1(n4320), .B2(n4185), .A(n4184), .ZN(n4321) );
  NAND2_X1 U4803 ( .A1(n4321), .A2(n4215), .ZN(n4195) );
  INV_X1 U4804 ( .A(n4208), .ZN(n4189) );
  INV_X1 U4805 ( .A(n4186), .ZN(n4187) );
  OAI21_X1 U4806 ( .B1(n4189), .B2(n4188), .A(n4187), .ZN(n4395) );
  INV_X1 U4807 ( .A(n4395), .ZN(n4193) );
  INV_X1 U4808 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4190) );
  OAI22_X1 U4809 ( .A1(n4191), .A2(n4508), .B1(n4511), .B2(n4190), .ZN(n4192)
         );
  AOI21_X1 U4810 ( .B1(n4193), .B2(n4514), .A(n4192), .ZN(n4194) );
  OAI211_X1 U4811 ( .C1(n4320), .C2(n4246), .A(n4195), .B(n4194), .ZN(U3270)
         );
  XNOR2_X1 U4812 ( .A(n4196), .B(n4202), .ZN(n4326) );
  INV_X1 U4813 ( .A(n4326), .ZN(n4217) );
  NAND2_X1 U4814 ( .A1(n2060), .A2(n4197), .ZN(n4221) );
  INV_X1 U4815 ( .A(n4198), .ZN(n4200) );
  OAI21_X1 U4816 ( .B1(n4221), .B2(n4200), .A(n4199), .ZN(n4201) );
  XOR2_X1 U4817 ( .A(n4202), .B(n4201), .Z(n4207) );
  OAI22_X1 U4818 ( .A1(n4338), .A2(n4349), .B1(n4203), .B2(n4209), .ZN(n4204)
         );
  AOI21_X1 U4819 ( .B1(n4346), .B2(n4312), .A(n4204), .ZN(n4205) );
  OAI21_X1 U4820 ( .B1(n4207), .B2(n4206), .A(n4205), .ZN(n4325) );
  INV_X1 U4821 ( .A(n4218), .ZN(n4210) );
  OAI21_X1 U4822 ( .B1(n4210), .B2(n4209), .A(n4208), .ZN(n4399) );
  AOI22_X1 U4823 ( .A1(n4520), .A2(REG2_REG_19__SCAN_IN), .B1(n4211), .B2(
        n4250), .ZN(n4212) );
  OAI21_X1 U4824 ( .B1(n4399), .B2(n4213), .A(n4212), .ZN(n4214) );
  AOI21_X1 U4825 ( .B1(n4325), .B2(n4215), .A(n4214), .ZN(n4216) );
  OAI21_X1 U4826 ( .B1(n4217), .B2(n4239), .A(n4216), .ZN(U3271) );
  OAI211_X1 U4827 ( .C1(n4220), .C2(n4219), .A(n4352), .B(n4218), .ZN(n4329)
         );
  XNOR2_X1 U4828 ( .A(n4221), .B(n4238), .ZN(n4226) );
  AOI22_X1 U4829 ( .A1(n4347), .A2(n4333), .B1(n4222), .B2(n4345), .ZN(n4223)
         );
  OAI21_X1 U4830 ( .B1(n4224), .B2(n4337), .A(n4223), .ZN(n4225) );
  AOI21_X1 U4831 ( .B1(n4226), .B2(n2715), .A(n4225), .ZN(n4330) );
  OAI21_X1 U4832 ( .B1(n4227), .B2(n4329), .A(n4330), .ZN(n4242) );
  OAI22_X1 U4833 ( .A1(n4511), .A2(n2232), .B1(n4228), .B2(n4508), .ZN(n4241)
         );
  NAND2_X1 U4834 ( .A1(n4230), .A2(n4229), .ZN(n4232) );
  AND2_X1 U4835 ( .A1(n4232), .A2(n4231), .ZN(n4237) );
  OR2_X1 U4836 ( .A1(n3457), .A2(n4233), .ZN(n4235) );
  AND2_X1 U4837 ( .A1(n4235), .A2(n4234), .ZN(n4236) );
  AOI21_X1 U4838 ( .B1(n4238), .B2(n4237), .A(n4236), .ZN(n4331) );
  NOR2_X1 U4839 ( .A1(n4331), .A2(n4239), .ZN(n4240) );
  AOI211_X1 U4840 ( .C1(n4511), .C2(n4242), .A(n4241), .B(n4240), .ZN(n4243)
         );
  INV_X1 U4841 ( .A(n4243), .ZN(U3272) );
  MUX2_X1 U4842 ( .A(n4245), .B(n4244), .S(n4511), .Z(n4259) );
  INV_X1 U4843 ( .A(n4246), .ZN(n4515) );
  AOI22_X1 U4844 ( .A1(n4249), .A2(n4515), .B1(n4248), .B2(n4247), .ZN(n4258)
         );
  AOI22_X1 U4845 ( .A1(n4252), .A2(n4251), .B1(REG3_REG_2__SCAN_IN), .B2(n4250), .ZN(n4257) );
  AOI22_X1 U4846 ( .A1(n4514), .A2(n4255), .B1(n4254), .B2(n4253), .ZN(n4256)
         );
  NAND4_X1 U4847 ( .A1(n4259), .A2(n4258), .A3(n4257), .A4(n4256), .ZN(U3288)
         );
  NOR2_X1 U4848 ( .A1(n4552), .A2(n4260), .ZN(n4261) );
  AOI21_X1 U4849 ( .B1(n4552), .B2(n4357), .A(n4261), .ZN(n4262) );
  OAI21_X1 U4850 ( .B1(n4360), .B2(n4343), .A(n4262), .ZN(U3549) );
  AOI21_X1 U4851 ( .B1(n4267), .B2(n4264), .A(n4263), .ZN(n4420) );
  INV_X1 U4852 ( .A(n4420), .ZN(n4363) );
  INV_X1 U4853 ( .A(n4265), .ZN(n4266) );
  AOI21_X1 U4854 ( .B1(n4267), .B2(n4345), .A(n4266), .ZN(n4422) );
  MUX2_X1 U4855 ( .A(n2717), .B(n4422), .S(n4552), .Z(n4268) );
  OAI21_X1 U4856 ( .B1(n4363), .B2(n4343), .A(n4268), .ZN(U3548) );
  AOI22_X1 U4857 ( .A1(n4270), .A2(n4333), .B1(n4269), .B2(n4345), .ZN(n4271)
         );
  OAI211_X1 U4858 ( .C1(n4273), .C2(n4337), .A(n4272), .B(n4271), .ZN(n4274)
         );
  AOI21_X1 U4859 ( .B1(n4275), .B2(n4340), .A(n4274), .ZN(n4364) );
  MUX2_X1 U4860 ( .A(n4276), .B(n4364), .S(n4552), .Z(n4277) );
  OAI21_X1 U4861 ( .B1(n4343), .B2(n4367), .A(n4277), .ZN(U3545) );
  AOI21_X1 U4862 ( .B1(n4279), .B2(n4340), .A(n4278), .ZN(n4368) );
  MUX2_X1 U4863 ( .A(n4280), .B(n4368), .S(n4552), .Z(n4281) );
  OAI21_X1 U4864 ( .B1(n4343), .B2(n4371), .A(n4281), .ZN(U3544) );
  AOI22_X1 U4865 ( .A1(n4283), .A2(n4333), .B1(n4282), .B2(n4345), .ZN(n4284)
         );
  OAI211_X1 U4866 ( .C1(n4286), .C2(n4337), .A(n4285), .B(n4284), .ZN(n4287)
         );
  AOI21_X1 U4867 ( .B1(n4288), .B2(n4340), .A(n4287), .ZN(n4372) );
  MUX2_X1 U4868 ( .A(n4289), .B(n4372), .S(n4552), .Z(n4290) );
  OAI21_X1 U4869 ( .B1(n4343), .B2(n4375), .A(n4290), .ZN(U3543) );
  AOI22_X1 U4870 ( .A1(n4292), .A2(n4333), .B1(n4345), .B2(n4291), .ZN(n4293)
         );
  OAI211_X1 U4871 ( .C1(n4295), .C2(n4337), .A(n4294), .B(n4293), .ZN(n4296)
         );
  AOI21_X1 U4872 ( .B1(n4297), .B2(n4340), .A(n4296), .ZN(n4376) );
  MUX2_X1 U4873 ( .A(n4298), .B(n4376), .S(n4552), .Z(n4299) );
  OAI21_X1 U4874 ( .B1(n4343), .B2(n4379), .A(n4299), .ZN(U3542) );
  AOI21_X1 U4875 ( .B1(n4301), .B2(n4340), .A(n4300), .ZN(n4380) );
  MUX2_X1 U4876 ( .A(n4302), .B(n4380), .S(n4552), .Z(n4303) );
  OAI21_X1 U4877 ( .B1(n4343), .B2(n4383), .A(n4303), .ZN(U3541) );
  NAND2_X1 U4878 ( .A1(n4304), .A2(n4340), .ZN(n4305) );
  OR2_X1 U4879 ( .A1(n4306), .A2(n4305), .ZN(n4308) );
  NAND2_X1 U4880 ( .A1(n4308), .A2(n4307), .ZN(n4384) );
  MUX2_X1 U4881 ( .A(n4384), .B(REG1_REG_22__SCAN_IN), .S(n4549), .Z(n4309) );
  INV_X1 U4882 ( .A(n4309), .ZN(n4310) );
  OAI21_X1 U4883 ( .B1(n4343), .B2(n4387), .A(n4310), .ZN(U3540) );
  AOI22_X1 U4884 ( .A1(n4312), .A2(n4333), .B1(n4311), .B2(n4345), .ZN(n4313)
         );
  OAI211_X1 U4885 ( .C1(n4315), .C2(n4337), .A(n4314), .B(n4313), .ZN(n4316)
         );
  AOI21_X1 U4886 ( .B1(n4317), .B2(n4340), .A(n4316), .ZN(n4388) );
  MUX2_X1 U4887 ( .A(n4318), .B(n4388), .S(n4552), .Z(n4319) );
  OAI21_X1 U4888 ( .B1(n4343), .B2(n4391), .A(n4319), .ZN(U3539) );
  INV_X1 U4889 ( .A(n4320), .ZN(n4322) );
  AOI21_X1 U4890 ( .B1(n4536), .B2(n4322), .A(n4321), .ZN(n4392) );
  MUX2_X1 U4891 ( .A(n4323), .B(n4392), .S(n4552), .Z(n4324) );
  OAI21_X1 U4892 ( .B1(n4343), .B2(n4395), .A(n4324), .ZN(U3538) );
  AOI21_X1 U4893 ( .B1(n4326), .B2(n4340), .A(n4325), .ZN(n4397) );
  MUX2_X1 U4894 ( .A(n4397), .B(n4327), .S(n4549), .Z(n4328) );
  OAI21_X1 U4895 ( .B1(n4343), .B2(n4399), .A(n4328), .ZN(U3537) );
  OAI211_X1 U4896 ( .C1(n4331), .C2(n4538), .A(n4330), .B(n4329), .ZN(n4400)
         );
  MUX2_X1 U4897 ( .A(REG1_REG_18__SCAN_IN), .B(n4400), .S(n4552), .Z(U3536) );
  AOI22_X1 U4898 ( .A1(n4334), .A2(n4333), .B1(n4332), .B2(n4345), .ZN(n4335)
         );
  OAI211_X1 U4899 ( .C1(n4338), .C2(n4337), .A(n4336), .B(n4335), .ZN(n4339)
         );
  AOI21_X1 U4900 ( .B1(n4341), .B2(n4340), .A(n4339), .ZN(n4402) );
  MUX2_X1 U4901 ( .A(n4402), .B(n2376), .S(n4549), .Z(n4342) );
  OAI21_X1 U4902 ( .B1(n4343), .B2(n4405), .A(n4342), .ZN(U3535) );
  AOI22_X1 U4903 ( .A1(n4347), .A2(n4346), .B1(n4345), .B2(n4344), .ZN(n4348)
         );
  OAI21_X1 U4904 ( .B1(n4350), .B2(n4349), .A(n4348), .ZN(n4351) );
  AOI21_X1 U4905 ( .B1(n4353), .B2(n4352), .A(n4351), .ZN(n4355) );
  OAI211_X1 U4906 ( .C1(n4356), .C2(n4538), .A(n4355), .B(n4354), .ZN(n4406)
         );
  MUX2_X1 U4907 ( .A(REG1_REG_16__SCAN_IN), .B(n4406), .S(n4552), .Z(U3534) );
  NAND2_X1 U4908 ( .A1(n4546), .A2(n4357), .ZN(n4359) );
  NAND2_X1 U4909 ( .A1(n4544), .A2(REG0_REG_31__SCAN_IN), .ZN(n4358) );
  OAI211_X1 U4910 ( .C1(n4360), .C2(n4404), .A(n4359), .B(n4358), .ZN(U3517)
         );
  INV_X1 U4911 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4361) );
  MUX2_X1 U4912 ( .A(n4361), .B(n4422), .S(n4546), .Z(n4362) );
  OAI21_X1 U4913 ( .B1(n4363), .B2(n4404), .A(n4362), .ZN(U3516) );
  INV_X1 U4914 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4365) );
  MUX2_X1 U4915 ( .A(n4365), .B(n4364), .S(n4546), .Z(n4366) );
  OAI21_X1 U4916 ( .B1(n4367), .B2(n4404), .A(n4366), .ZN(U3513) );
  INV_X1 U4917 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4369) );
  MUX2_X1 U4918 ( .A(n4369), .B(n4368), .S(n4546), .Z(n4370) );
  OAI21_X1 U4919 ( .B1(n4371), .B2(n4404), .A(n4370), .ZN(U3512) );
  INV_X1 U4920 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4373) );
  MUX2_X1 U4921 ( .A(n4373), .B(n4372), .S(n4546), .Z(n4374) );
  OAI21_X1 U4922 ( .B1(n4375), .B2(n4404), .A(n4374), .ZN(U3511) );
  INV_X1 U4923 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4377) );
  MUX2_X1 U4924 ( .A(n4377), .B(n4376), .S(n4546), .Z(n4378) );
  OAI21_X1 U4925 ( .B1(n4379), .B2(n4404), .A(n4378), .ZN(U3510) );
  INV_X1 U4926 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4381) );
  MUX2_X1 U4927 ( .A(n4381), .B(n4380), .S(n4546), .Z(n4382) );
  OAI21_X1 U4928 ( .B1(n4383), .B2(n4404), .A(n4382), .ZN(U3509) );
  MUX2_X1 U4929 ( .A(REG0_REG_22__SCAN_IN), .B(n4384), .S(n4546), .Z(n4385) );
  INV_X1 U4930 ( .A(n4385), .ZN(n4386) );
  OAI21_X1 U4931 ( .B1(n4387), .B2(n4404), .A(n4386), .ZN(U3508) );
  INV_X1 U4932 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4389) );
  MUX2_X1 U4933 ( .A(n4389), .B(n4388), .S(n4546), .Z(n4390) );
  OAI21_X1 U4934 ( .B1(n4391), .B2(n4404), .A(n4390), .ZN(U3507) );
  INV_X1 U4935 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4393) );
  MUX2_X1 U4936 ( .A(n4393), .B(n4392), .S(n4546), .Z(n4394) );
  OAI21_X1 U4937 ( .B1(n4395), .B2(n4404), .A(n4394), .ZN(U3506) );
  INV_X1 U4938 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4396) );
  MUX2_X1 U4939 ( .A(n4397), .B(n4396), .S(n4544), .Z(n4398) );
  OAI21_X1 U4940 ( .B1(n4399), .B2(n4404), .A(n4398), .ZN(U3505) );
  MUX2_X1 U4941 ( .A(REG0_REG_18__SCAN_IN), .B(n4400), .S(n4546), .Z(U3503) );
  INV_X1 U4942 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4401) );
  MUX2_X1 U4943 ( .A(n4402), .B(n4401), .S(n4544), .Z(n4403) );
  OAI21_X1 U4944 ( .B1(n4405), .B2(n4404), .A(n4403), .ZN(U3501) );
  MUX2_X1 U4945 ( .A(REG0_REG_16__SCAN_IN), .B(n4406), .S(n4546), .Z(U3499) );
  MUX2_X1 U4946 ( .A(DATAI_30_), .B(n4407), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4947 ( .A(n4408), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4948 ( .A(n2729), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U4949 ( .A(DATAI_22_), .B(n4409), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4950 ( .A(DATAI_20_), .B(n4410), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4951 ( .A(DATAI_8_), .B(n2148), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U4952 ( .A(n4412), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4953 ( .A(DATAI_5_), .B(n2143), .S(STATE_REG_SCAN_IN), .Z(U3347) );
  MUX2_X1 U4954 ( .A(DATAI_4_), .B(n4413), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4955 ( .A(DATAI_3_), .B(n4414), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U4956 ( .A(DATAI_2_), .B(n4415), .S(STATE_REG_SCAN_IN), .Z(U3350) );
  MUX2_X1 U4957 ( .A(n4416), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U4958 ( .A1(STATE_REG_SCAN_IN), .A2(n4418), .B1(n4417), .B2(U3149), 
        .ZN(U3324) );
  OAI21_X1 U4959 ( .B1(n4520), .B2(n4422), .A(n4421), .ZN(U3261) );
  INV_X1 U4960 ( .A(n4425), .ZN(n4423) );
  OAI211_X1 U4961 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4424), .A(n4426), .B(n4423), 
        .ZN(n4430) );
  AOI22_X1 U4962 ( .A1(n4426), .A2(n4425), .B1(n4502), .B2(n2855), .ZN(n4428)
         );
  AOI22_X1 U4963 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4501), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4427) );
  OAI221_X1 U4964 ( .B1(IR_REG_0__SCAN_IN), .B2(n4430), .C1(n4429), .C2(n4428), 
        .A(n4427), .ZN(U3240) );
  OAI211_X1 U4965 ( .C1(n4433), .C2(n4432), .A(n4466), .B(n4431), .ZN(n4438)
         );
  OAI211_X1 U4966 ( .C1(n4436), .C2(n4435), .A(n4502), .B(n4434), .ZN(n4437)
         );
  OAI211_X1 U4967 ( .C1(n4507), .C2(n4439), .A(n4438), .B(n4437), .ZN(n4440)
         );
  AOI211_X1 U4968 ( .C1(n4501), .C2(ADDR_REG_9__SCAN_IN), .A(n4441), .B(n4440), 
        .ZN(n4442) );
  INV_X1 U4969 ( .A(n4442), .ZN(U3249) );
  OAI211_X1 U4970 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4445), .A(n4466), .B(n4444), .ZN(n4447) );
  NAND2_X1 U4971 ( .A1(n4447), .A2(n4446), .ZN(n4448) );
  AOI21_X1 U4972 ( .B1(n4501), .B2(ADDR_REG_10__SCAN_IN), .A(n4448), .ZN(n4452) );
  OAI211_X1 U4973 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4450), .A(n4502), .B(n4449), .ZN(n4451) );
  OAI211_X1 U4974 ( .C1(n4507), .C2(n2284), .A(n4452), .B(n4451), .ZN(U3250)
         );
  OAI211_X1 U4975 ( .C1(n4455), .C2(n4454), .A(n4502), .B(n4453), .ZN(n4460)
         );
  OAI211_X1 U4976 ( .C1(n4458), .C2(n4457), .A(n4466), .B(n4456), .ZN(n4459)
         );
  OAI211_X1 U4977 ( .C1(n4507), .C2(n4527), .A(n4460), .B(n4459), .ZN(n4461)
         );
  AOI211_X1 U4978 ( .C1(n4501), .C2(ADDR_REG_11__SCAN_IN), .A(n4462), .B(n4461), .ZN(n4463) );
  INV_X1 U4979 ( .A(n4463), .ZN(U3251) );
  OAI211_X1 U4980 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4467), .A(n4466), .B(n4465), .ZN(n4469) );
  NAND2_X1 U4981 ( .A1(n4469), .A2(n4468), .ZN(n4470) );
  AOI21_X1 U4982 ( .B1(n4501), .B2(ADDR_REG_12__SCAN_IN), .A(n4470), .ZN(n4474) );
  OAI211_X1 U4983 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4472), .A(n4502), .B(n4471), .ZN(n4473) );
  OAI211_X1 U4984 ( .C1(n4507), .C2(n2288), .A(n4474), .B(n4473), .ZN(U3252)
         );
  INV_X1 U4985 ( .A(n4475), .ZN(n4480) );
  AOI211_X1 U4986 ( .C1(n4478), .C2(n4477), .A(n4476), .B(n4495), .ZN(n4479)
         );
  AOI211_X1 U4987 ( .C1(n4501), .C2(ADDR_REG_14__SCAN_IN), .A(n4480), .B(n4479), .ZN(n4484) );
  OAI211_X1 U4988 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4482), .A(n4502), .B(n4481), .ZN(n4483) );
  OAI211_X1 U4989 ( .C1(n4507), .C2(n2146), .A(n4484), .B(n4483), .ZN(U3254)
         );
  AOI211_X1 U4990 ( .C1(n2067), .C2(n4486), .A(n4485), .B(n4495), .ZN(n4487)
         );
  AOI211_X1 U4991 ( .C1(n4501), .C2(ADDR_REG_15__SCAN_IN), .A(n4488), .B(n4487), .ZN(n4493) );
  OAI211_X1 U4992 ( .C1(n4491), .C2(n4490), .A(n4502), .B(n4489), .ZN(n4492)
         );
  OAI211_X1 U4993 ( .C1(n4507), .C2(n4525), .A(n4493), .B(n4492), .ZN(U3255)
         );
  INV_X1 U4994 ( .A(n4494), .ZN(n4500) );
  AOI221_X1 U4995 ( .B1(n4498), .B2(n4497), .C1(n4496), .C2(n4497), .A(n4495), 
        .ZN(n4499) );
  AOI211_X1 U4996 ( .C1(n4501), .C2(ADDR_REG_16__SCAN_IN), .A(n4500), .B(n4499), .ZN(n4506) );
  OAI221_X1 U4997 ( .B1(n4504), .B2(REG1_REG_16__SCAN_IN), .C1(n4504), .C2(
        n4503), .A(n4502), .ZN(n4505) );
  OAI211_X1 U4998 ( .C1(n4507), .C2(n4524), .A(n4506), .B(n4505), .ZN(U3256)
         );
  OAI22_X1 U4999 ( .A1(n4511), .A2(n4510), .B1(n4509), .B2(n4508), .ZN(n4512)
         );
  INV_X1 U5000 ( .A(n4512), .ZN(n4518) );
  AOI22_X1 U5001 ( .A1(n4516), .A2(n4515), .B1(n4514), .B2(n4513), .ZN(n4517)
         );
  OAI211_X1 U5002 ( .C1(n4520), .C2(n4519), .A(n4518), .B(n4517), .ZN(U3282)
         );
  AND2_X1 U5003 ( .A1(D_REG_31__SCAN_IN), .A2(n4521), .ZN(U3291) );
  AND2_X1 U5004 ( .A1(D_REG_30__SCAN_IN), .A2(n4521), .ZN(U3292) );
  AND2_X1 U5005 ( .A1(D_REG_29__SCAN_IN), .A2(n4521), .ZN(U3293) );
  AND2_X1 U5006 ( .A1(D_REG_28__SCAN_IN), .A2(n4521), .ZN(U3294) );
  AND2_X1 U5007 ( .A1(D_REG_27__SCAN_IN), .A2(n4521), .ZN(U3295) );
  AND2_X1 U5008 ( .A1(D_REG_26__SCAN_IN), .A2(n4521), .ZN(U3296) );
  AND2_X1 U5009 ( .A1(D_REG_25__SCAN_IN), .A2(n4521), .ZN(U3297) );
  AND2_X1 U5010 ( .A1(D_REG_24__SCAN_IN), .A2(n4521), .ZN(U3298) );
  AND2_X1 U5011 ( .A1(D_REG_23__SCAN_IN), .A2(n4521), .ZN(U3299) );
  AND2_X1 U5012 ( .A1(D_REG_22__SCAN_IN), .A2(n4521), .ZN(U3300) );
  AND2_X1 U5013 ( .A1(D_REG_21__SCAN_IN), .A2(n4521), .ZN(U3301) );
  AND2_X1 U5014 ( .A1(D_REG_20__SCAN_IN), .A2(n4521), .ZN(U3302) );
  AND2_X1 U5015 ( .A1(D_REG_19__SCAN_IN), .A2(n4521), .ZN(U3303) );
  AND2_X1 U5016 ( .A1(D_REG_18__SCAN_IN), .A2(n4521), .ZN(U3304) );
  AND2_X1 U5017 ( .A1(D_REG_17__SCAN_IN), .A2(n4521), .ZN(U3305) );
  AND2_X1 U5018 ( .A1(D_REG_16__SCAN_IN), .A2(n4521), .ZN(U3306) );
  AND2_X1 U5019 ( .A1(D_REG_15__SCAN_IN), .A2(n4521), .ZN(U3307) );
  AND2_X1 U5020 ( .A1(D_REG_14__SCAN_IN), .A2(n4521), .ZN(U3308) );
  AND2_X1 U5021 ( .A1(D_REG_13__SCAN_IN), .A2(n4521), .ZN(U3309) );
  AND2_X1 U5022 ( .A1(D_REG_12__SCAN_IN), .A2(n4521), .ZN(U3310) );
  AND2_X1 U5023 ( .A1(D_REG_11__SCAN_IN), .A2(n4521), .ZN(U3311) );
  AND2_X1 U5024 ( .A1(D_REG_10__SCAN_IN), .A2(n4521), .ZN(U3312) );
  AND2_X1 U5025 ( .A1(D_REG_9__SCAN_IN), .A2(n4521), .ZN(U3313) );
  AND2_X1 U5026 ( .A1(D_REG_8__SCAN_IN), .A2(n4521), .ZN(U3314) );
  AND2_X1 U5027 ( .A1(D_REG_7__SCAN_IN), .A2(n4521), .ZN(U3315) );
  AND2_X1 U5028 ( .A1(D_REG_6__SCAN_IN), .A2(n4521), .ZN(U3316) );
  AND2_X1 U5029 ( .A1(D_REG_5__SCAN_IN), .A2(n4521), .ZN(U3317) );
  AND2_X1 U5030 ( .A1(D_REG_4__SCAN_IN), .A2(n4521), .ZN(U3318) );
  AND2_X1 U5031 ( .A1(D_REG_3__SCAN_IN), .A2(n4521), .ZN(U3319) );
  AND2_X1 U5032 ( .A1(D_REG_2__SCAN_IN), .A2(n4521), .ZN(U3320) );
  AOI21_X1 U5033 ( .B1(U3149), .B2(n2646), .A(n4522), .ZN(U3329) );
  INV_X1 U5034 ( .A(DATAI_18_), .ZN(n4576) );
  AOI22_X1 U5035 ( .A1(STATE_REG_SCAN_IN), .A2(n4523), .B1(n4576), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5036 ( .A(DATAI_16_), .ZN(n4590) );
  AOI22_X1 U5037 ( .A1(STATE_REG_SCAN_IN), .A2(n4524), .B1(n4590), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5038 ( .A(DATAI_15_), .ZN(n4666) );
  AOI22_X1 U5039 ( .A1(STATE_REG_SCAN_IN), .A2(n4525), .B1(n4666), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5040 ( .A(DATAI_14_), .ZN(n4645) );
  AOI22_X1 U5041 ( .A1(STATE_REG_SCAN_IN), .A2(n2146), .B1(n4645), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5042 ( .A(DATAI_12_), .ZN(n4526) );
  AOI22_X1 U5043 ( .A1(STATE_REG_SCAN_IN), .A2(n2288), .B1(n4526), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5044 ( .A(DATAI_11_), .ZN(n4643) );
  AOI22_X1 U5045 ( .A1(STATE_REG_SCAN_IN), .A2(n4527), .B1(n4643), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5046 ( .A(DATAI_10_), .ZN(n4667) );
  AOI22_X1 U5047 ( .A1(STATE_REG_SCAN_IN), .A2(n2284), .B1(n4667), .B2(U3149), 
        .ZN(U3342) );
  OAI211_X1 U5048 ( .C1(n4531), .C2(n4530), .A(n4529), .B(n4528), .ZN(n4532)
         );
  INV_X1 U5049 ( .A(n4532), .ZN(n4547) );
  AOI22_X1 U5050 ( .A1(n4546), .A2(n4547), .B1(n2424), .B2(n4544), .ZN(U3467)
         );
  INV_X1 U5051 ( .A(n4533), .ZN(n4535) );
  AOI211_X1 U5052 ( .C1(n4537), .C2(n4536), .A(n4535), .B(n4534), .ZN(n4548)
         );
  AOI22_X1 U5053 ( .A1(n4546), .A2(n4548), .B1(n2447), .B2(n4544), .ZN(U3475)
         );
  NOR2_X1 U5054 ( .A1(n4539), .A2(n4538), .ZN(n4543) );
  AOI211_X1 U5055 ( .C1(n4543), .C2(n4542), .A(n4541), .B(n4540), .ZN(n4551)
         );
  INV_X1 U5056 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4545) );
  AOI22_X1 U5057 ( .A1(n4546), .A2(n4551), .B1(n4545), .B2(n4544), .ZN(U3481)
         );
  AOI22_X1 U5058 ( .A1(n4552), .A2(n4547), .B1(n2855), .B2(n4549), .ZN(U3518)
         );
  AOI22_X1 U5059 ( .A1(n4552), .A2(n4548), .B1(n2440), .B2(n4549), .ZN(U3522)
         );
  AOI22_X1 U5060 ( .A1(n4552), .A2(n4551), .B1(n4550), .B2(n4549), .ZN(U3525)
         );
  AOI22_X1 U5061 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n4737) );
  AOI22_X1 U5062 ( .A1(n4646), .A2(keyinput_g48), .B1(keyinput_g6), .B2(n2408), 
        .ZN(n4553) );
  OAI221_X1 U5063 ( .B1(n4646), .B2(keyinput_g48), .C1(n2408), .C2(keyinput_g6), .A(n4553), .ZN(n4562) );
  AOI22_X1 U5064 ( .A1(n4555), .A2(keyinput_g1), .B1(n4645), .B2(keyinput_g17), 
        .ZN(n4554) );
  OAI221_X1 U5065 ( .B1(n4555), .B2(keyinput_g1), .C1(n4645), .C2(keyinput_g17), .A(n4554), .ZN(n4561) );
  XOR2_X1 U5066 ( .A(n2501), .B(keyinput_g51), .Z(n4559) );
  XNOR2_X1 U5067 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_g59), .ZN(n4558) );
  XNOR2_X1 U5068 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_g35), .ZN(n4557) );
  XNOR2_X1 U5069 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_g61), .ZN(n4556) );
  NAND4_X1 U5070 ( .A1(n4559), .A2(n4558), .A3(n4557), .A4(n4556), .ZN(n4560)
         );
  NOR3_X1 U5071 ( .A1(n4562), .A2(n4561), .A3(n4560), .ZN(n4601) );
  AOI22_X1 U5072 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput_g34), .B1(n2390), 
        .B2(keyinput_g4), .ZN(n4563) );
  OAI221_X1 U5073 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput_g34), .C1(n2390), 
        .C2(keyinput_g4), .A(n4563), .ZN(n4571) );
  AOI22_X1 U5074 ( .A1(DATAI_9_), .A2(keyinput_g22), .B1(DATAI_11_), .B2(
        keyinput_g20), .ZN(n4564) );
  OAI221_X1 U5075 ( .B1(DATAI_9_), .B2(keyinput_g22), .C1(DATAI_11_), .C2(
        keyinput_g20), .A(n4564), .ZN(n4570) );
  AOI22_X1 U5076 ( .A1(REG3_REG_10__SCAN_IN), .A2(keyinput_g37), .B1(
        REG3_REG_16__SCAN_IN), .B2(keyinput_g46), .ZN(n4565) );
  OAI221_X1 U5077 ( .B1(REG3_REG_10__SCAN_IN), .B2(keyinput_g37), .C1(
        REG3_REG_16__SCAN_IN), .C2(keyinput_g46), .A(n4565), .ZN(n4569) );
  XNOR2_X1 U5078 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_g58), .ZN(n4567) );
  XNOR2_X1 U5079 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_g39), .ZN(n4566) );
  NAND2_X1 U5080 ( .A1(n4567), .A2(n4566), .ZN(n4568) );
  NOR4_X1 U5081 ( .A1(n4571), .A2(n4570), .A3(n4569), .A4(n4568), .ZN(n4600)
         );
  INV_X1 U5082 ( .A(DATAI_1_), .ZN(n4573) );
  AOI22_X1 U5083 ( .A1(n4574), .A2(keyinput_g53), .B1(keyinput_g30), .B2(n4573), .ZN(n4572) );
  OAI221_X1 U5084 ( .B1(n4574), .B2(keyinput_g53), .C1(n4573), .C2(
        keyinput_g30), .A(n4572), .ZN(n4583) );
  AOI22_X1 U5085 ( .A1(n3607), .A2(keyinput_g40), .B1(keyinput_g13), .B2(n4576), .ZN(n4575) );
  OAI221_X1 U5086 ( .B1(n3607), .B2(keyinput_g40), .C1(n4576), .C2(
        keyinput_g13), .A(n4575), .ZN(n4582) );
  XOR2_X1 U5087 ( .A(n4666), .B(keyinput_g16), .Z(n4580) );
  XOR2_X1 U5088 ( .A(n2273), .B(keyinput_g62), .Z(n4579) );
  XNOR2_X1 U5089 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_g38), .ZN(n4578) );
  XNOR2_X1 U5090 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_g42), .ZN(n4577) );
  NAND4_X1 U5091 ( .A1(n4580), .A2(n4579), .A3(n4578), .A4(n4577), .ZN(n4581)
         );
  NOR3_X1 U5092 ( .A1(n4583), .A2(n4582), .A3(n4581), .ZN(n4599) );
  AOI22_X1 U5093 ( .A1(n2463), .A2(keyinput_g33), .B1(n4585), .B2(keyinput_g57), .ZN(n4584) );
  OAI221_X1 U5094 ( .B1(n2463), .B2(keyinput_g33), .C1(n4585), .C2(
        keyinput_g57), .A(n4584), .ZN(n4597) );
  AOI22_X1 U5095 ( .A1(n4588), .A2(keyinput_g7), .B1(n4587), .B2(keyinput_g18), 
        .ZN(n4586) );
  OAI221_X1 U5096 ( .B1(n4588), .B2(keyinput_g7), .C1(n4587), .C2(keyinput_g18), .A(n4586), .ZN(n4596) );
  INV_X1 U5097 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4681) );
  AOI22_X1 U5098 ( .A1(n4681), .A2(keyinput_g41), .B1(keyinput_g15), .B2(n4590), .ZN(n4589) );
  OAI221_X1 U5099 ( .B1(n4681), .B2(keyinput_g41), .C1(n4590), .C2(
        keyinput_g15), .A(n4589), .ZN(n4595) );
  XOR2_X1 U5100 ( .A(n4591), .B(keyinput_g2), .Z(n4593) );
  XNOR2_X1 U5101 ( .A(DATAI_2_), .B(keyinput_g29), .ZN(n4592) );
  NAND2_X1 U5102 ( .A1(n4593), .A2(n4592), .ZN(n4594) );
  NOR4_X1 U5103 ( .A1(n4597), .A2(n4596), .A3(n4595), .A4(n4594), .ZN(n4598)
         );
  NAND4_X1 U5104 ( .A1(n4601), .A2(n4600), .A3(n4599), .A4(n4598), .ZN(n4735)
         );
  AOI22_X1 U5105 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput_g52), .B1(DATAI_19_), 
        .B2(keyinput_g12), .ZN(n4602) );
  OAI221_X1 U5106 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput_g52), .C1(DATAI_19_), .C2(keyinput_g12), .A(n4602), .ZN(n4609) );
  AOI22_X1 U5107 ( .A1(DATAI_4_), .A2(keyinput_g27), .B1(DATAI_28_), .B2(
        keyinput_g3), .ZN(n4603) );
  OAI221_X1 U5108 ( .B1(DATAI_4_), .B2(keyinput_g27), .C1(DATAI_28_), .C2(
        keyinput_g3), .A(n4603), .ZN(n4608) );
  AOI22_X1 U5109 ( .A1(DATAI_23_), .A2(keyinput_g8), .B1(DATAI_26_), .B2(
        keyinput_g5), .ZN(n4604) );
  OAI221_X1 U5110 ( .B1(DATAI_23_), .B2(keyinput_g8), .C1(DATAI_26_), .C2(
        keyinput_g5), .A(n4604), .ZN(n4607) );
  AOI22_X1 U5111 ( .A1(DATAI_31_), .A2(keyinput_g0), .B1(REG3_REG_24__SCAN_IN), 
        .B2(keyinput_g49), .ZN(n4605) );
  OAI221_X1 U5112 ( .B1(DATAI_31_), .B2(keyinput_g0), .C1(REG3_REG_24__SCAN_IN), .C2(keyinput_g49), .A(n4605), .ZN(n4606) );
  NOR4_X1 U5113 ( .A1(n4609), .A2(n4608), .A3(n4607), .A4(n4606), .ZN(n4637)
         );
  XNOR2_X1 U5114 ( .A(DATAI_22_), .B(keyinput_g9), .ZN(n4617) );
  AOI22_X1 U5115 ( .A1(DATAI_10_), .A2(keyinput_g21), .B1(n4611), .B2(
        keyinput_g36), .ZN(n4610) );
  OAI221_X1 U5116 ( .B1(DATAI_10_), .B2(keyinput_g21), .C1(n4611), .C2(
        keyinput_g36), .A(n4610), .ZN(n4616) );
  AOI22_X1 U5117 ( .A1(REG3_REG_25__SCAN_IN), .A2(keyinput_g45), .B1(
        STATE_REG_SCAN_IN), .B2(keyinput_g32), .ZN(n4612) );
  OAI221_X1 U5118 ( .B1(REG3_REG_25__SCAN_IN), .B2(keyinput_g45), .C1(
        STATE_REG_SCAN_IN), .C2(keyinput_g32), .A(n4612), .ZN(n4615) );
  AOI22_X1 U5119 ( .A1(DATAI_21_), .A2(keyinput_g10), .B1(REG3_REG_21__SCAN_IN), .B2(keyinput_g43), .ZN(n4613) );
  OAI221_X1 U5120 ( .B1(DATAI_21_), .B2(keyinput_g10), .C1(
        REG3_REG_21__SCAN_IN), .C2(keyinput_g43), .A(n4613), .ZN(n4614) );
  NOR4_X1 U5121 ( .A1(n4617), .A2(n4616), .A3(n4615), .A4(n4614), .ZN(n4636)
         );
  AOI22_X1 U5122 ( .A1(DATAI_3_), .A2(keyinput_g28), .B1(REG3_REG_4__SCAN_IN), 
        .B2(keyinput_g50), .ZN(n4618) );
  OAI221_X1 U5123 ( .B1(DATAI_3_), .B2(keyinput_g28), .C1(REG3_REG_4__SCAN_IN), 
        .C2(keyinput_g50), .A(n4618), .ZN(n4625) );
  AOI22_X1 U5124 ( .A1(DATAI_0_), .A2(keyinput_g31), .B1(IR_REG_1__SCAN_IN), 
        .B2(keyinput_g56), .ZN(n4619) );
  OAI221_X1 U5125 ( .B1(DATAI_0_), .B2(keyinput_g31), .C1(IR_REG_1__SCAN_IN), 
        .C2(keyinput_g56), .A(n4619), .ZN(n4624) );
  AOI22_X1 U5126 ( .A1(DATAI_8_), .A2(keyinput_g23), .B1(IR_REG_8__SCAN_IN), 
        .B2(keyinput_g63), .ZN(n4620) );
  OAI221_X1 U5127 ( .B1(DATAI_8_), .B2(keyinput_g23), .C1(IR_REG_8__SCAN_IN), 
        .C2(keyinput_g63), .A(n4620), .ZN(n4623) );
  AOI22_X1 U5128 ( .A1(REG3_REG_5__SCAN_IN), .A2(keyinput_g47), .B1(
        IR_REG_5__SCAN_IN), .B2(keyinput_g60), .ZN(n4621) );
  OAI221_X1 U5129 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput_g47), .C1(
        IR_REG_5__SCAN_IN), .C2(keyinput_g60), .A(n4621), .ZN(n4622) );
  NOR4_X1 U5130 ( .A1(n4625), .A2(n4624), .A3(n4623), .A4(n4622), .ZN(n4635)
         );
  AOI22_X1 U5131 ( .A1(REG3_REG_12__SCAN_IN), .A2(keyinput_g44), .B1(
        IR_REG_0__SCAN_IN), .B2(keyinput_g55), .ZN(n4626) );
  OAI221_X1 U5132 ( .B1(REG3_REG_12__SCAN_IN), .B2(keyinput_g44), .C1(
        IR_REG_0__SCAN_IN), .C2(keyinput_g55), .A(n4626), .ZN(n4633) );
  AOI22_X1 U5133 ( .A1(DATAI_17_), .A2(keyinput_g14), .B1(DATAI_20_), .B2(
        keyinput_g11), .ZN(n4627) );
  OAI221_X1 U5134 ( .B1(DATAI_17_), .B2(keyinput_g14), .C1(DATAI_20_), .C2(
        keyinput_g11), .A(n4627), .ZN(n4632) );
  AOI22_X1 U5135 ( .A1(DATAI_6_), .A2(keyinput_g25), .B1(DATAI_12_), .B2(
        keyinput_g19), .ZN(n4628) );
  OAI221_X1 U5136 ( .B1(DATAI_6_), .B2(keyinput_g25), .C1(DATAI_12_), .C2(
        keyinput_g19), .A(n4628), .ZN(n4631) );
  AOI22_X1 U5137 ( .A1(DATAI_7_), .A2(keyinput_g24), .B1(REG3_REG_13__SCAN_IN), 
        .B2(keyinput_g54), .ZN(n4629) );
  OAI221_X1 U5138 ( .B1(DATAI_7_), .B2(keyinput_g24), .C1(REG3_REG_13__SCAN_IN), .C2(keyinput_g54), .A(n4629), .ZN(n4630) );
  NOR4_X1 U5139 ( .A1(n4633), .A2(n4632), .A3(n4631), .A4(n4630), .ZN(n4634)
         );
  NAND4_X1 U5140 ( .A1(n4637), .A2(n4636), .A3(n4635), .A4(n4634), .ZN(n4734)
         );
  AOI22_X1 U5141 ( .A1(n4640), .A2(keyinput_f34), .B1(keyinput_f35), .B2(n4639), .ZN(n4638) );
  OAI221_X1 U5142 ( .B1(n4640), .B2(keyinput_f34), .C1(n4639), .C2(
        keyinput_f35), .A(n4638), .ZN(n4652) );
  AOI22_X1 U5143 ( .A1(n4643), .A2(keyinput_f20), .B1(n4642), .B2(keyinput_f5), 
        .ZN(n4641) );
  OAI221_X1 U5144 ( .B1(n4643), .B2(keyinput_f20), .C1(n4642), .C2(keyinput_f5), .A(n4641), .ZN(n4651) );
  AOI22_X1 U5145 ( .A1(n4646), .A2(keyinput_f48), .B1(keyinput_f17), .B2(n4645), .ZN(n4644) );
  OAI221_X1 U5146 ( .B1(n4646), .B2(keyinput_f48), .C1(n4645), .C2(
        keyinput_f17), .A(n4644), .ZN(n4650) );
  XNOR2_X1 U5147 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_f59), .ZN(n4648) );
  XNOR2_X1 U5148 ( .A(DATAI_12_), .B(keyinput_f19), .ZN(n4647) );
  NAND2_X1 U5149 ( .A1(n4648), .A2(n4647), .ZN(n4649) );
  NOR4_X1 U5150 ( .A1(n4652), .A2(n4651), .A3(n4650), .A4(n4649), .ZN(n4692)
         );
  AOI22_X1 U5151 ( .A1(DATAI_22_), .A2(keyinput_f9), .B1(REG3_REG_20__SCAN_IN), 
        .B2(keyinput_f53), .ZN(n4653) );
  OAI221_X1 U5152 ( .B1(DATAI_22_), .B2(keyinput_f9), .C1(REG3_REG_20__SCAN_IN), .C2(keyinput_f53), .A(n4653), .ZN(n4662) );
  AOI22_X1 U5153 ( .A1(DATAI_18_), .A2(keyinput_f13), .B1(STATE_REG_SCAN_IN), 
        .B2(keyinput_f32), .ZN(n4654) );
  OAI221_X1 U5154 ( .B1(DATAI_18_), .B2(keyinput_f13), .C1(STATE_REG_SCAN_IN), 
        .C2(keyinput_f32), .A(n4654), .ZN(n4661) );
  AOI22_X1 U5155 ( .A1(n4656), .A2(keyinput_f47), .B1(n2539), .B2(keyinput_f54), .ZN(n4655) );
  OAI221_X1 U5156 ( .B1(n4656), .B2(keyinput_f47), .C1(n2539), .C2(
        keyinput_f54), .A(n4655), .ZN(n4660) );
  AOI22_X1 U5157 ( .A1(n4658), .A2(keyinput_f37), .B1(keyinput_f28), .B2(n2477), .ZN(n4657) );
  OAI221_X1 U5158 ( .B1(n4658), .B2(keyinput_f37), .C1(n2477), .C2(
        keyinput_f28), .A(n4657), .ZN(n4659) );
  NOR4_X1 U5159 ( .A1(n4662), .A2(n4661), .A3(n4660), .A4(n4659), .ZN(n4691)
         );
  INV_X1 U5160 ( .A(DATAI_0_), .ZN(n4664) );
  AOI22_X1 U5161 ( .A1(n2273), .A2(keyinput_f62), .B1(keyinput_f31), .B2(n4664), .ZN(n4663) );
  OAI221_X1 U5162 ( .B1(n2273), .B2(keyinput_f62), .C1(n4664), .C2(
        keyinput_f31), .A(n4663), .ZN(n4677) );
  AOI22_X1 U5163 ( .A1(n4667), .A2(keyinput_f21), .B1(n4666), .B2(keyinput_f16), .ZN(n4665) );
  OAI221_X1 U5164 ( .B1(n4667), .B2(keyinput_f21), .C1(n4666), .C2(
        keyinput_f16), .A(n4665), .ZN(n4676) );
  AOI22_X1 U5165 ( .A1(n4670), .A2(keyinput_f23), .B1(n4669), .B2(keyinput_f10), .ZN(n4668) );
  OAI221_X1 U5166 ( .B1(n4670), .B2(keyinput_f23), .C1(n4669), .C2(
        keyinput_f10), .A(n4668), .ZN(n4675) );
  INV_X1 U5167 ( .A(IR_REG_1__SCAN_IN), .ZN(n4671) );
  XOR2_X1 U5168 ( .A(n4671), .B(keyinput_f56), .Z(n4673) );
  XNOR2_X1 U5169 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_f42), .ZN(n4672) );
  NAND2_X1 U5170 ( .A1(n4673), .A2(n4672), .ZN(n4674) );
  NOR4_X1 U5171 ( .A1(n4677), .A2(n4676), .A3(n4675), .A4(n4674), .ZN(n4690)
         );
  AOI22_X1 U5172 ( .A1(n2646), .A2(keyinput_f8), .B1(n2463), .B2(keyinput_f33), 
        .ZN(n4678) );
  OAI221_X1 U5173 ( .B1(n2646), .B2(keyinput_f8), .C1(n2463), .C2(keyinput_f33), .A(n4678), .ZN(n4688) );
  AOI22_X1 U5174 ( .A1(n4681), .A2(keyinput_f41), .B1(keyinput_f14), .B2(n4680), .ZN(n4679) );
  OAI221_X1 U5175 ( .B1(n4681), .B2(keyinput_f41), .C1(n4680), .C2(
        keyinput_f14), .A(n4679), .ZN(n4687) );
  XNOR2_X1 U5176 ( .A(REG3_REG_25__SCAN_IN), .B(keyinput_f45), .ZN(n4685) );
  XNOR2_X1 U5177 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_f50), .ZN(n4684) );
  XNOR2_X1 U5178 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_f61), .ZN(n4683) );
  XNOR2_X1 U5179 ( .A(DATAI_2_), .B(keyinput_f29), .ZN(n4682) );
  NAND4_X1 U5180 ( .A1(n4685), .A2(n4684), .A3(n4683), .A4(n4682), .ZN(n4686)
         );
  NOR3_X1 U5181 ( .A1(n4688), .A2(n4687), .A3(n4686), .ZN(n4689) );
  NAND4_X1 U5182 ( .A1(n4692), .A2(n4691), .A3(n4690), .A4(n4689), .ZN(n4729)
         );
  AOI22_X1 U5183 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(DATAI_25_), .B2(
        keyinput_f6), .ZN(n4693) );
  OAI221_X1 U5184 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(DATAI_25_), .C2(
        keyinput_f6), .A(n4693), .ZN(n4700) );
  AOI22_X1 U5185 ( .A1(DATAI_31_), .A2(keyinput_f0), .B1(DATAI_27_), .B2(
        keyinput_f4), .ZN(n4694) );
  OAI221_X1 U5186 ( .B1(DATAI_31_), .B2(keyinput_f0), .C1(DATAI_27_), .C2(
        keyinput_f4), .A(n4694), .ZN(n4699) );
  AOI22_X1 U5187 ( .A1(REG3_REG_12__SCAN_IN), .A2(keyinput_f44), .B1(
        IR_REG_0__SCAN_IN), .B2(keyinput_f55), .ZN(n4695) );
  OAI221_X1 U5188 ( .B1(REG3_REG_12__SCAN_IN), .B2(keyinput_f44), .C1(
        IR_REG_0__SCAN_IN), .C2(keyinput_f55), .A(n4695), .ZN(n4698) );
  AOI22_X1 U5189 ( .A1(DATAI_20_), .A2(keyinput_f11), .B1(REG3_REG_3__SCAN_IN), 
        .B2(keyinput_f38), .ZN(n4696) );
  OAI221_X1 U5190 ( .B1(DATAI_20_), .B2(keyinput_f11), .C1(REG3_REG_3__SCAN_IN), .C2(keyinput_f38), .A(n4696), .ZN(n4697) );
  NOR4_X1 U5191 ( .A1(n4700), .A2(n4699), .A3(n4698), .A4(n4697), .ZN(n4727)
         );
  XNOR2_X1 U5192 ( .A(DATAI_4_), .B(keyinput_f27), .ZN(n4707) );
  AOI22_X1 U5193 ( .A1(DATAI_28_), .A2(keyinput_f3), .B1(n3669), .B2(
        keyinput_f43), .ZN(n4701) );
  OAI221_X1 U5194 ( .B1(DATAI_28_), .B2(keyinput_f3), .C1(n3669), .C2(
        keyinput_f43), .A(n4701), .ZN(n4706) );
  AOI22_X1 U5195 ( .A1(REG3_REG_24__SCAN_IN), .A2(keyinput_f49), .B1(
        REG3_REG_28__SCAN_IN), .B2(keyinput_f40), .ZN(n4702) );
  OAI221_X1 U5196 ( .B1(REG3_REG_24__SCAN_IN), .B2(keyinput_f49), .C1(
        REG3_REG_28__SCAN_IN), .C2(keyinput_f40), .A(n4702), .ZN(n4705) );
  AOI22_X1 U5197 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput_f52), .B1(DATAI_19_), 
        .B2(keyinput_f12), .ZN(n4703) );
  OAI221_X1 U5198 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput_f52), .C1(DATAI_19_), .C2(keyinput_f12), .A(n4703), .ZN(n4704) );
  NOR4_X1 U5199 ( .A1(n4707), .A2(n4706), .A3(n4705), .A4(n4704), .ZN(n4726)
         );
  AOI22_X1 U5200 ( .A1(DATAI_16_), .A2(keyinput_f15), .B1(REG3_REG_23__SCAN_IN), .B2(keyinput_f36), .ZN(n4708) );
  OAI221_X1 U5201 ( .B1(DATAI_16_), .B2(keyinput_f15), .C1(
        REG3_REG_23__SCAN_IN), .C2(keyinput_f36), .A(n4708), .ZN(n4715) );
  AOI22_X1 U5202 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput_f51), .B1(
        REG3_REG_16__SCAN_IN), .B2(keyinput_f46), .ZN(n4709) );
  OAI221_X1 U5203 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput_f51), .C1(
        REG3_REG_16__SCAN_IN), .C2(keyinput_f46), .A(n4709), .ZN(n4714) );
  AOI22_X1 U5204 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(REG3_REG_19__SCAN_IN), 
        .B2(keyinput_f39), .ZN(n4710) );
  OAI221_X1 U5205 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(REG3_REG_19__SCAN_IN), .C2(keyinput_f39), .A(n4710), .ZN(n4713) );
  AOI22_X1 U5206 ( .A1(DATAI_13_), .A2(keyinput_f18), .B1(DATAI_29_), .B2(
        keyinput_f2), .ZN(n4711) );
  OAI221_X1 U5207 ( .B1(DATAI_13_), .B2(keyinput_f18), .C1(DATAI_29_), .C2(
        keyinput_f2), .A(n4711), .ZN(n4712) );
  NOR4_X1 U5208 ( .A1(n4715), .A2(n4714), .A3(n4713), .A4(n4712), .ZN(n4725)
         );
  AOI22_X1 U5209 ( .A1(DATAI_1_), .A2(keyinput_f30), .B1(IR_REG_2__SCAN_IN), 
        .B2(keyinput_f57), .ZN(n4716) );
  OAI221_X1 U5210 ( .B1(DATAI_1_), .B2(keyinput_f30), .C1(IR_REG_2__SCAN_IN), 
        .C2(keyinput_f57), .A(n4716), .ZN(n4723) );
  AOI22_X1 U5211 ( .A1(DATAI_7_), .A2(keyinput_f24), .B1(DATAI_6_), .B2(
        keyinput_f25), .ZN(n4717) );
  OAI221_X1 U5212 ( .B1(DATAI_7_), .B2(keyinput_f24), .C1(DATAI_6_), .C2(
        keyinput_f25), .A(n4717), .ZN(n4722) );
  AOI22_X1 U5213 ( .A1(DATAI_9_), .A2(keyinput_f22), .B1(IR_REG_8__SCAN_IN), 
        .B2(keyinput_f63), .ZN(n4718) );
  OAI221_X1 U5214 ( .B1(DATAI_9_), .B2(keyinput_f22), .C1(IR_REG_8__SCAN_IN), 
        .C2(keyinput_f63), .A(n4718), .ZN(n4721) );
  AOI22_X1 U5215 ( .A1(IR_REG_3__SCAN_IN), .A2(keyinput_f58), .B1(
        IR_REG_5__SCAN_IN), .B2(keyinput_f60), .ZN(n4719) );
  OAI221_X1 U5216 ( .B1(IR_REG_3__SCAN_IN), .B2(keyinput_f58), .C1(
        IR_REG_5__SCAN_IN), .C2(keyinput_f60), .A(n4719), .ZN(n4720) );
  NOR4_X1 U5217 ( .A1(n4723), .A2(n4722), .A3(n4721), .A4(n4720), .ZN(n4724)
         );
  NAND4_X1 U5218 ( .A1(n4727), .A2(n4726), .A3(n4725), .A4(n4724), .ZN(n4728)
         );
  OAI22_X1 U5219 ( .A1(keyinput_f26), .A2(n2456), .B1(n4729), .B2(n4728), .ZN(
        n4730) );
  OAI21_X1 U5220 ( .B1(n4730), .B2(keyinput_f26), .A(n2456), .ZN(n4732) );
  NAND3_X1 U5221 ( .A1(n4730), .A2(keyinput_g26), .A3(DATAI_5_), .ZN(n4731) );
  OAI21_X1 U5222 ( .B1(keyinput_g26), .B2(n4732), .A(n4731), .ZN(n4733) );
  OAI21_X1 U5223 ( .B1(n4735), .B2(n4734), .A(n4733), .ZN(n4736) );
  XOR2_X1 U5224 ( .A(n4737), .B(n4736), .Z(U3352) );
  CLKBUF_X1 U2287 ( .A(n2856), .Z(n2044) );
  CLKBUF_X1 U2305 ( .A(n2875), .Z(n3599) );
endmodule

