

module b15_C_gen_AntiSAT_k_128_5 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, 
        U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, 
        U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, 
        U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, 
        U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, 
        U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, 
        U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, 
        U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, 
        U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, 
        U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, 
        U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, 
        U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, 
        U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, 
        U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, 
        U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, 
        U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, 
        U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, 
        U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, 
        U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, 
        U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, 
        U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, 
        U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, 
        U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, 
        U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, 
        U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, 
        U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, 
        U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, 
        U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, 
        U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, 
        U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, 
        U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, 
        U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, 
        U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, 
        U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, 
        U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, 
        U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, 
        U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, 
        U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, 
        U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, 
        U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, 
        U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, 
        U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, 
        U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, 
        U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, 
        U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, 
        U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838;

  CLKBUF_X2 U3433 ( .A(n3565), .Z(n3796) );
  CLKBUF_X2 U3434 ( .A(n3795), .Z(n3881) );
  CLKBUF_X2 U3435 ( .A(n3283), .Z(n3879) );
  CLKBUF_X2 U3436 ( .A(n3148), .Z(n3819) );
  CLKBUF_X2 U3437 ( .A(n3168), .Z(n3840) );
  CLKBUF_X2 U3438 ( .A(n3107), .Z(n3769) );
  INV_X1 U3440 ( .A(n5391), .ZN(n4295) );
  INV_X1 U3441 ( .A(n4222), .ZN(n3207) );
  CLKBUF_X2 U3442 ( .A(n3158), .Z(n5392) );
  CLKBUF_X2 U3443 ( .A(n3566), .Z(n3775) );
  INV_X1 U3444 ( .A(n6210), .ZN(n6156) );
  INV_X1 U34450 ( .A(n4442), .ZN(n4285) );
  AND2_X2 U34470 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4484) );
  INV_X1 U34480 ( .A(n4398), .ZN(n2986) );
  INV_X1 U3449 ( .A(n4117), .ZN(n4442) );
  INV_X1 U34510 ( .A(n6338), .ZN(n6376) );
  NAND2_X1 U34520 ( .A1(n3973), .A2(n3976), .ZN(n4003) );
  AND2_X1 U34530 ( .A1(n3389), .A2(n3412), .ZN(n4637) );
  NAND2_X2 U34550 ( .A1(n5626), .A2(n5613), .ZN(n5644) );
  NAND2_X2 U34560 ( .A1(n3236), .A2(n3264), .ZN(n3365) );
  OR2_X1 U3457 ( .A1(n3222), .A2(n4650), .ZN(n2985) );
  OR2_X1 U3458 ( .A1(n3222), .A2(n4650), .ZN(n4118) );
  AND2_X4 U34590 ( .A1(n4424), .A2(n4489), .ZN(n3862) );
  AND2_X4 U34600 ( .A1(n4489), .A2(n4484), .ZN(n3251) );
  AND2_X4 U34610 ( .A1(n3070), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4489) );
  XNOR2_X2 U34620 ( .A(n3942), .B(n4133), .ZN(n4618) );
  NAND2_X2 U34630 ( .A1(n3941), .A2(n3940), .ZN(n3942) );
  NAND2_X1 U34640 ( .A1(n5690), .A2(n5689), .ZN(n5669) );
  INV_X1 U34650 ( .A(n4003), .ZN(n2998) );
  NOR2_X2 U3466 ( .A1(n4563), .A2(n4686), .ZN(n4685) );
  OAI21_X1 U3467 ( .B1(n3950), .B2(n3975), .A(n3949), .ZN(n3952) );
  NAND2_X1 U34680 ( .A1(n4628), .A2(n3364), .ZN(n4564) );
  CLKBUF_X1 U34690 ( .A(n4637), .Z(n4638) );
  BUF_X2 U34700 ( .A(n3184), .Z(n3195) );
  AND2_X1 U34710 ( .A1(n4081), .A2(n4080), .ZN(n4082) );
  XNOR2_X1 U34720 ( .A(n4269), .B(n3905), .ZN(n5369) );
  OR2_X1 U34730 ( .A1(n5712), .A2(n6297), .ZN(n4081) );
  AOI21_X1 U34740 ( .B1(n5495), .B2(n5494), .A(n4364), .ZN(n6007) );
  AOI22_X1 U3475 ( .A1(n5597), .A2(n5596), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5595), .ZN(n5599) );
  NAND2_X1 U3476 ( .A1(n4088), .A2(n4087), .ZN(n5596) );
  NAND2_X1 U3477 ( .A1(n5669), .A2(n3015), .ZN(n5610) );
  NAND2_X1 U3478 ( .A1(n3036), .A2(n3038), .ZN(n5309) );
  OR2_X1 U3479 ( .A1(n2990), .A2(n3048), .ZN(n2989) );
  NAND2_X1 U3480 ( .A1(n4003), .A2(n3980), .ZN(n3981) );
  INV_X4 U3481 ( .A(n2998), .ZN(n2999) );
  OAI21_X1 U3482 ( .B1(n3957), .B2(n3975), .A(n3956), .ZN(n3959) );
  XNOR2_X1 U3483 ( .A(n3973), .B(n3472), .ZN(n3962) );
  OAI21_X1 U3484 ( .B1(n3950), .B2(n3552), .A(n3445), .ZN(n4713) );
  NAND2_X1 U3485 ( .A1(n3458), .A2(n3459), .ZN(n3973) );
  XNOR2_X1 U3486 ( .A(n3934), .B(n3912), .ZN(n4555) );
  NAND2_X1 U3487 ( .A1(n3911), .A2(n3910), .ZN(n3934) );
  NAND2_X1 U3488 ( .A1(n4314), .A2(n4313), .ZN(n6210) );
  NAND2_X1 U3489 ( .A1(n3386), .A2(n3385), .ZN(n4663) );
  CLKBUF_X1 U3490 ( .A(n4639), .Z(n5821) );
  CLKBUF_X1 U3491 ( .A(n4482), .Z(n6399) );
  CLKBUF_X1 U3492 ( .A(n3341), .Z(n3342) );
  NOR2_X1 U3493 ( .A1(n6715), .A2(n4806), .ZN(n6481) );
  NAND2_X2 U3494 ( .A1(n3354), .A2(n3353), .ZN(n5052) );
  NOR2_X1 U3495 ( .A1(n6712), .A2(n4806), .ZN(n6475) );
  NOR2_X1 U3496 ( .A1(n6662), .A2(n4806), .ZN(n6496) );
  NOR2_X1 U3497 ( .A1(n4676), .A2(n4806), .ZN(n6469) );
  NAND2_X1 U3498 ( .A1(n3320), .A2(n3319), .ZN(n3340) );
  NAND2_X1 U3499 ( .A1(n3281), .A2(n3280), .ZN(n3341) );
  NOR2_X1 U3500 ( .A1(n6284), .A2(n4471), .ZN(n6283) );
  NAND2_X1 U3501 ( .A1(n4395), .A2(n4393), .ZN(n6638) );
  OAI21_X1 U3502 ( .B1(n3232), .B2(n3231), .A(n4650), .ZN(n4220) );
  NAND2_X1 U3503 ( .A1(n3052), .A2(n4398), .ZN(n3051) );
  AND3_X1 U3504 ( .A1(n3211), .A2(n3210), .A3(n2997), .ZN(n4216) );
  AND3_X1 U3505 ( .A1(n5100), .A2(n3208), .A3(n3207), .ZN(n3214) );
  AND2_X2 U3506 ( .A1(n4277), .A2(n3373), .ZN(n4057) );
  INV_X1 U3507 ( .A(n3221), .ZN(n4544) );
  NAND2_X1 U3508 ( .A1(n3313), .A2(n3195), .ZN(n4069) );
  CLKBUF_X1 U3509 ( .A(n3908), .Z(n6634) );
  CLKBUF_X1 U3510 ( .A(n3183), .Z(n3155) );
  OR2_X1 U3511 ( .A1(n3212), .A2(n6636), .ZN(n4277) );
  INV_X1 U3512 ( .A(n3187), .ZN(n3194) );
  NAND4_X1 U3513 ( .A1(n3180), .A2(n3179), .A3(n3178), .A4(n3177), .ZN(n3187)
         );
  INV_X2 U3514 ( .A(n4650), .ZN(n2987) );
  NAND2_X1 U3515 ( .A1(n3113), .A2(n3112), .ZN(n3184) );
  AND4_X1 U3516 ( .A1(n3117), .A2(n3116), .A3(n3115), .A4(n3114), .ZN(n3122)
         );
  AND4_X1 U3517 ( .A1(n3090), .A2(n3089), .A3(n3088), .A4(n3087), .ZN(n3101)
         );
  AND4_X1 U3518 ( .A1(n3094), .A2(n3093), .A3(n3092), .A4(n3091), .ZN(n3100)
         );
  AND4_X1 U3519 ( .A1(n3098), .A2(n3097), .A3(n3096), .A4(n3095), .ZN(n3099)
         );
  AND4_X1 U3520 ( .A1(n3111), .A2(n3110), .A3(n3109), .A4(n3108), .ZN(n3112)
         );
  AND4_X1 U3521 ( .A1(n3167), .A2(n3166), .A3(n3165), .A4(n3164), .ZN(n3179)
         );
  AND4_X1 U3522 ( .A1(n3162), .A2(n3161), .A3(n3160), .A4(n3159), .ZN(n3180)
         );
  AND4_X1 U3523 ( .A1(n3135), .A2(n3134), .A3(n3133), .A4(n3132), .ZN(n3140)
         );
  INV_X1 U3524 ( .A(n3378), .ZN(n2996) );
  AND4_X1 U3525 ( .A1(n3106), .A2(n3105), .A3(n3104), .A4(n3103), .ZN(n3113)
         );
  BUF_X2 U3526 ( .A(n3887), .Z(n3768) );
  AND2_X1 U3527 ( .A1(n3147), .A2(n3146), .ZN(n3152) );
  AND4_X1 U3528 ( .A1(n3176), .A2(n3175), .A3(n3174), .A4(n3173), .ZN(n3177)
         );
  AND4_X1 U3529 ( .A1(n3086), .A2(n3085), .A3(n3084), .A4(n3083), .ZN(n3102)
         );
  AND4_X1 U3530 ( .A1(n3172), .A2(n3171), .A3(n3170), .A4(n3169), .ZN(n3178)
         );
  AND4_X1 U3531 ( .A1(n3145), .A2(n3144), .A3(n3143), .A4(n3142), .ZN(n3154)
         );
  BUF_X2 U3532 ( .A(n3862), .Z(n3813) );
  INV_X2 U3533 ( .A(n3250), .ZN(n3774) );
  BUF_X2 U3534 ( .A(n3273), .Z(n3880) );
  NAND2_X1 U3535 ( .A1(n3906), .A2(n6408), .ZN(n6335) );
  BUF_X2 U3536 ( .A(n3282), .Z(n3877) );
  BUF_X2 U3537 ( .A(n3878), .Z(n3818) );
  AND2_X2 U3538 ( .A1(n4425), .A2(n4485), .ZN(n3283) );
  AND2_X2 U3539 ( .A1(n4488), .A2(n4484), .ZN(n3245) );
  AND2_X2 U3540 ( .A1(n4489), .A2(n4425), .ZN(n3273) );
  AND2_X4 U3541 ( .A1(n4520), .A2(n4485), .ZN(n3565) );
  AND2_X2 U3542 ( .A1(n3069), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4425)
         );
  INV_X1 U3543 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3396) );
  NAND2_X2 U3544 ( .A1(n3972), .A2(n3971), .ZN(n5160) );
  AND2_X2 U3545 ( .A1(n5005), .A2(n5177), .ZN(n5156) );
  NAND2_X1 U3546 ( .A1(n5160), .A2(n2991), .ZN(n2988) );
  AND2_X2 U3547 ( .A1(n2988), .A2(n2989), .ZN(n5269) );
  INV_X1 U3548 ( .A(n3983), .ZN(n2990) );
  AND2_X1 U3549 ( .A1(n5161), .A2(n3983), .ZN(n2991) );
  NOR2_X2 U3550 ( .A1(n5530), .A2(n5532), .ZN(n5460) );
  NAND2_X1 U3551 ( .A1(n5810), .A2(n2995), .ZN(n2992) );
  AND2_X2 U3552 ( .A1(n2992), .A2(n2993), .ZN(n5690) );
  OR2_X1 U3553 ( .A1(n2994), .A2(n3987), .ZN(n2993) );
  INV_X1 U3554 ( .A(n3988), .ZN(n2994) );
  AND2_X1 U3555 ( .A1(n3986), .A2(n3988), .ZN(n2995) );
  NAND2_X1 U3556 ( .A1(n3158), .A2(n3183), .ZN(n2997) );
  NAND2_X1 U3557 ( .A1(n3158), .A2(n3183), .ZN(n3209) );
  NAND2_X2 U3558 ( .A1(n5610), .A2(n3995), .ZN(n5659) );
  NOR2_X2 U3559 ( .A1(n5512), .A2(n5514), .ZN(n5447) );
  BUF_X4 U3560 ( .A(n3845), .Z(n3888) );
  NAND2_X1 U3561 ( .A1(n4022), .A2(n4020), .ZN(n4052) );
  NOR2_X1 U3562 ( .A1(n5500), .A2(n5491), .ZN(n3032) );
  NAND2_X1 U3563 ( .A1(n3182), .A2(n2987), .ZN(n4300) );
  OR2_X1 U3564 ( .A1(n4306), .A2(n5535), .ZN(n4307) );
  OR2_X1 U3565 ( .A1(n4053), .A2(n6394), .ZN(n4055) );
  INV_X1 U3566 ( .A(n4098), .ZN(n4060) );
  NOR2_X1 U3567 ( .A1(n5414), .A2(n3062), .ZN(n3061) );
  INV_X1 U3568 ( .A(n5422), .ZN(n3062) );
  INV_X1 U3569 ( .A(n5495), .ZN(n3058) );
  NAND2_X1 U3570 ( .A1(n5156), .A2(n3017), .ZN(n3559) );
  OR2_X1 U3571 ( .A1(n4117), .A2(n5467), .ZN(n4305) );
  AND2_X1 U3572 ( .A1(n3195), .A2(n4398), .ZN(n4020) );
  AND2_X2 U3573 ( .A1(n3225), .A2(n3195), .ZN(n3221) );
  AND2_X1 U3574 ( .A1(n3260), .A2(n3212), .ZN(n4022) );
  XNOR2_X1 U3575 ( .A(n4522), .B(n4873), .ZN(n4482) );
  AND3_X1 U3576 ( .A1(n3207), .A2(n5392), .A3(n3222), .ZN(n3181) );
  NOR2_X1 U3577 ( .A1(n5500), .A2(n3022), .ZN(n5426) );
  AND2_X1 U3578 ( .A1(n3032), .A2(n3033), .ZN(n4306) );
  NOR3_X1 U3579 ( .A1(n4209), .A2(n3034), .A3(n3035), .ZN(n3033) );
  NOR2_X2 U3580 ( .A1(n5478), .A2(n5477), .ZN(n5563) );
  OR2_X1 U3581 ( .A1(n4534), .A2(n4108), .ZN(n4109) );
  OR2_X1 U3582 ( .A1(n4104), .A2(n4211), .ZN(n6531) );
  INV_X1 U3583 ( .A(n3938), .ZN(n3945) );
  AOI22_X1 U3584 ( .A1(n3251), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3163), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3111) );
  CLKBUF_X1 U3585 ( .A(n3888), .Z(n3857) );
  OAI21_X1 U3586 ( .B1(n4057), .B2(n3435), .A(n3434), .ZN(n3438) );
  OAI21_X1 U3587 ( .B1(n4057), .B2(n3457), .A(n3456), .ZN(n3459) );
  OR2_X1 U3588 ( .A1(n3257), .A2(n3256), .ZN(n3907) );
  NAND2_X1 U3589 ( .A1(n3251), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3146)
         );
  INV_X1 U3590 ( .A(n5498), .ZN(n3788) );
  INV_X1 U3591 ( .A(n5542), .ZN(n3657) );
  INV_X1 U3592 ( .A(n3872), .ZN(n3900) );
  NOR2_X1 U3593 ( .A1(n3056), .A2(n3055), .ZN(n3054) );
  INV_X1 U3594 ( .A(n5560), .ZN(n3055) );
  NAND2_X1 U3595 ( .A1(n3057), .A2(n5344), .ZN(n3056) );
  INV_X1 U3596 ( .A(n5475), .ZN(n3057) );
  INV_X1 U3597 ( .A(n5264), .ZN(n3537) );
  AND2_X1 U3598 ( .A1(n3156), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3356) );
  INV_X1 U3599 ( .A(n4199), .ZN(n4205) );
  INV_X1 U3600 ( .A(n5296), .ZN(n3040) );
  NOR2_X1 U3601 ( .A1(n3040), .A2(n5271), .ZN(n3037) );
  INV_X1 U3602 ( .A(n5008), .ZN(n3031) );
  INV_X1 U3603 ( .A(n4305), .ZN(n4200) );
  OR2_X1 U3604 ( .A1(n4285), .A2(n5535), .ZN(n4199) );
  OAI21_X1 U3605 ( .B1(n4305), .B2(EBX_REG_1__SCAN_IN), .A(n4120), .ZN(n4123)
         );
  OR2_X1 U3606 ( .A1(n3293), .A2(n3292), .ZN(n3977) );
  OR2_X1 U3607 ( .A1(n3310), .A2(n3309), .ZN(n3917) );
  OAI211_X1 U3608 ( .C1(n3296), .C2(n3373), .A(n3295), .B(n3300), .ZN(n3339)
         );
  AND2_X1 U3609 ( .A1(n4224), .A2(n4223), .ZN(n4420) );
  AND2_X1 U3610 ( .A1(n4216), .A2(n4068), .ZN(n4113) );
  INV_X1 U3611 ( .A(n4740), .ZN(n4143) );
  INV_X1 U3612 ( .A(n4741), .ZN(n4144) );
  NAND2_X1 U3613 ( .A1(n4118), .A2(n5467), .ZN(n4409) );
  AND2_X1 U3614 ( .A1(n4113), .A2(n4112), .ZN(n4540) );
  OR2_X2 U3615 ( .A1(n3082), .A2(n3081), .ZN(n4398) );
  NOR2_X1 U3616 ( .A1(n4534), .A2(n4396), .ZN(n4399) );
  XNOR2_X1 U3617 ( .A(n4076), .B(n4323), .ZN(n4350) );
  NAND2_X1 U3618 ( .A1(n4363), .A2(n3016), .ZN(n4269) );
  NAND2_X1 U3619 ( .A1(n3834), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3875)
         );
  NOR2_X1 U3620 ( .A1(n3807), .A2(n5606), .ZN(n3808) );
  CLKBUF_X1 U3621 ( .A(n5530), .Z(n5531) );
  NOR2_X1 U3622 ( .A1(n3506), .A2(n6128), .ZN(n3521) );
  INV_X1 U3623 ( .A(n3442), .ZN(n3443) );
  INV_X1 U3624 ( .A(n4565), .ZN(n3398) );
  AND2_X1 U3625 ( .A1(n4177), .A2(n3029), .ZN(n3028) );
  INV_X1 U3626 ( .A(n5538), .ZN(n3029) );
  NAND2_X1 U3627 ( .A1(n5303), .A2(n3014), .ZN(n5478) );
  INV_X1 U3628 ( .A(n5346), .ZN(n3024) );
  AND2_X1 U3629 ( .A1(n3007), .A2(n3982), .ZN(n3048) );
  CLKBUF_X1 U3630 ( .A(n4426), .Z(n4427) );
  CLKBUF_X1 U3631 ( .A(n4503), .Z(n4504) );
  AOI21_X1 U3632 ( .B1(n4872), .B2(STATEBS16_REG_SCAN_IN), .A(n5896), .ZN(
        n5047) );
  NAND2_X1 U3633 ( .A1(n5107), .A2(n4770), .ZN(n4967) );
  NAND2_X1 U3634 ( .A1(n6636), .A2(n4648), .ZN(n4806) );
  NAND2_X1 U3635 ( .A1(n4482), .A2(n6636), .ZN(n3386) );
  INV_X1 U3636 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6517) );
  AND2_X2 U3637 ( .A1(n4066), .A2(n4065), .ZN(n5406) );
  NAND2_X1 U3638 ( .A1(n4064), .A2(n4063), .ZN(n4065) );
  INV_X1 U3639 ( .A(n4100), .ZN(n4063) );
  INV_X1 U3640 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6822) );
  INV_X1 U3641 ( .A(n5380), .ZN(n5397) );
  AND2_X1 U3642 ( .A1(n5394), .A2(n3156), .ZN(n6247) );
  AND2_X1 U3643 ( .A1(n5394), .A2(n4546), .ZN(n5583) );
  AOI21_X1 U3644 ( .B1(n6310), .B2(n5435), .A(n4369), .ZN(n4370) );
  NOR2_X1 U3645 ( .A1(n4084), .A2(n4089), .ZN(n4090) );
  INV_X1 U3646 ( .A(n5596), .ZN(n4089) );
  NAND2_X1 U3647 ( .A1(n4374), .A2(n4383), .ZN(n4262) );
  NAND2_X1 U3648 ( .A1(n4294), .A2(n4293), .ZN(n5381) );
  NOR2_X1 U3649 ( .A1(n4384), .A2(n4383), .ZN(n4386) );
  INV_X1 U3650 ( .A(n6035), .ZN(n6383) );
  AND2_X1 U3651 ( .A1(n4235), .A2(n4213), .ZN(n6382) );
  INV_X1 U3652 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6401) );
  OR2_X1 U3653 ( .A1(n3352), .A2(n3351), .ZN(n3353) );
  AND2_X1 U3654 ( .A1(n4067), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6539) );
  INV_X1 U3655 ( .A(n6539), .ZN(n6545) );
  OAI21_X1 U3656 ( .B1(n4057), .B2(n3945), .A(n3410), .ZN(n3413) );
  OR2_X1 U3657 ( .A1(n3455), .A2(n3454), .ZN(n3964) );
  OR2_X1 U3658 ( .A1(n3433), .A2(n3432), .ZN(n3947) );
  OR2_X1 U3659 ( .A1(n3409), .A2(n3408), .ZN(n3938) );
  NAND2_X1 U3660 ( .A1(n3878), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3172) );
  OR2_X1 U3661 ( .A1(n3279), .A2(n3278), .ZN(n3916) );
  NAND2_X1 U3662 ( .A1(n2987), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4010) );
  NAND2_X1 U3663 ( .A1(n3221), .A2(n3313), .ZN(n3211) );
  AOI22_X1 U3664 ( .A1(n3163), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3148), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3080) );
  AND2_X1 U3665 ( .A1(n5622), .A2(n3829), .ZN(n3764) );
  AND2_X1 U3666 ( .A1(n5374), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3872) );
  AND2_X1 U3667 ( .A1(n3557), .A2(n3556), .ZN(n3558) );
  NOR2_X1 U3668 ( .A1(n3060), .A2(n5242), .ZN(n3059) );
  INV_X1 U3669 ( .A(n5158), .ZN(n3060) );
  INV_X1 U3670 ( .A(n5604), .ZN(n4002) );
  NOR2_X1 U3671 ( .A1(n3991), .A2(n3047), .ZN(n3046) );
  INV_X1 U3672 ( .A(n5677), .ZN(n3991) );
  INV_X1 U3673 ( .A(n3990), .ZN(n3047) );
  NOR2_X1 U3674 ( .A1(n5365), .A2(n3026), .ZN(n3025) );
  INV_X1 U3675 ( .A(n5281), .ZN(n3026) );
  XNOR2_X1 U3676 ( .A(n3263), .B(n3262), .ZN(n3328) );
  AOI22_X1 U3677 ( .A1(n4022), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3261), 
        .B2(n3907), .ZN(n3262) );
  NAND2_X1 U3678 ( .A1(n3259), .A2(n3258), .ZN(n3263) );
  NAND2_X1 U3679 ( .A1(n3328), .A2(n3327), .ZN(n3387) );
  INV_X1 U3680 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3070) );
  NAND2_X1 U3681 ( .A1(n3244), .A2(n3243), .ZN(n3366) );
  NAND2_X2 U3682 ( .A1(n3122), .A2(n3004), .ZN(n4222) );
  INV_X1 U3683 ( .A(n3184), .ZN(n3158) );
  AOI22_X1 U3684 ( .A1(n3283), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3107), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3145) );
  OAI21_X1 U3685 ( .B1(n6535), .B2(n4529), .A(n5838), .ZN(n4648) );
  INV_X1 U3686 ( .A(n4057), .ZN(n4035) );
  INV_X1 U3687 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5018) );
  INV_X1 U3688 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6512) );
  OR2_X1 U3689 ( .A1(n4057), .A2(n4100), .ZN(n4058) );
  INV_X1 U3690 ( .A(n4052), .ZN(n4064) );
  CLKBUF_X1 U3691 ( .A(n4300), .Z(n5398) );
  NOR2_X1 U3692 ( .A1(n4650), .A2(n4398), .ZN(n3908) );
  CLKBUF_X1 U3693 ( .A(n4093), .Z(n5402) );
  NOR2_X1 U3694 ( .A1(n6083), .A2(n4326), .ZN(n5965) );
  INV_X1 U3695 ( .A(n3577), .ZN(n3591) );
  NOR2_X1 U3696 ( .A1(n6582), .A2(n6140), .ZN(n5249) );
  NAND2_X1 U3697 ( .A1(n6156), .A2(n4324), .ZN(n6140) );
  INV_X1 U3698 ( .A(n3297), .ZN(n3298) );
  NOR2_X1 U3699 ( .A1(n5493), .A2(n4209), .ZN(n5424) );
  AND2_X1 U3700 ( .A1(n4204), .A2(n4203), .ZN(n5491) );
  INV_X1 U3701 ( .A(n3032), .ZN(n5493) );
  AOI21_X1 U3702 ( .B1(n3536), .B2(n3829), .A(n3535), .ZN(n5264) );
  INV_X1 U3703 ( .A(n6286), .ZN(n4471) );
  AND2_X1 U3704 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n3833), .ZN(n3834)
         );
  MUX2_X1 U3705 ( .A(n5592), .B(n3854), .S(n4301), .Z(n5422) );
  NAND2_X1 U3706 ( .A1(n3810), .A2(n3809), .ZN(n5495) );
  NAND2_X1 U3707 ( .A1(n3767), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3807)
         );
  AND2_X1 U3708 ( .A1(n3761), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3767)
         );
  CLKBUF_X1 U3709 ( .A(n4353), .Z(n5448) );
  INV_X1 U3710 ( .A(n3704), .ZN(n3705) );
  CLKBUF_X1 U3711 ( .A(n5512), .Z(n5513) );
  NOR2_X1 U3712 ( .A1(n3673), .A2(n5982), .ZN(n3674) );
  NAND2_X1 U3713 ( .A1(n3674), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3704)
         );
  NOR2_X1 U3714 ( .A1(n3653), .A2(n6084), .ZN(n3654) );
  NAND2_X1 U3715 ( .A1(n3654), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3673)
         );
  NAND2_X1 U3716 ( .A1(n3620), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3653)
         );
  NOR2_X1 U3717 ( .A1(n3607), .A2(n5686), .ZN(n3620) );
  CLKBUF_X1 U3718 ( .A(n5549), .Z(n5550) );
  NAND2_X1 U3719 ( .A1(n3591), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3607)
         );
  INV_X1 U3720 ( .A(n5342), .ZN(n3053) );
  AND2_X1 U3721 ( .A1(n3554), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3555)
         );
  NAND2_X1 U3722 ( .A1(n3555), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3577)
         );
  INV_X1 U3723 ( .A(n5358), .ZN(n3574) );
  OAI211_X1 U3724 ( .C1(n3553), .C2(n3552), .A(n3551), .B(n3550), .ZN(n5280)
         );
  NAND2_X1 U3725 ( .A1(n3521), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3549)
         );
  INV_X1 U3726 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3548) );
  INV_X1 U3727 ( .A(n3491), .ZN(n3492) );
  INV_X1 U3728 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U3729 ( .A1(n3473), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3491)
         );
  CLKBUF_X1 U3730 ( .A(n5005), .Z(n5006) );
  INV_X1 U3731 ( .A(n3467), .ZN(n3468) );
  INV_X1 U3732 ( .A(n3441), .ZN(n3444) );
  AOI21_X1 U3733 ( .B1(n3937), .B2(n3600), .A(n3423), .ZN(n4686) );
  INV_X1 U3734 ( .A(n3422), .ZN(n3423) );
  NOR2_X1 U3735 ( .A1(n3391), .A2(n3390), .ZN(n3417) );
  INV_X1 U3736 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3390) );
  NAND2_X1 U3737 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3391) );
  AND2_X1 U3738 ( .A1(n3362), .A2(n3361), .ZN(n4440) );
  OR2_X1 U3739 ( .A1(n4411), .A2(n3829), .ZN(n3361) );
  INV_X1 U3740 ( .A(n5703), .ZN(n3043) );
  NOR2_X1 U3741 ( .A1(n2999), .A2(n4086), .ZN(n4087) );
  INV_X1 U3742 ( .A(n4085), .ZN(n4088) );
  OR2_X1 U3743 ( .A1(n5503), .A2(n5502), .ZN(n5500) );
  NOR2_X1 U3744 ( .A1(n5519), .A2(n5452), .ZN(n5453) );
  OR2_X1 U3745 ( .A1(n5516), .A2(n5517), .ZN(n5519) );
  INV_X1 U3746 ( .A(n4185), .ZN(n3027) );
  AND2_X1 U3747 ( .A1(n4180), .A2(n4179), .ZN(n5538) );
  AND2_X1 U3748 ( .A1(n4173), .A2(n4172), .ZN(n5553) );
  NAND2_X1 U3749 ( .A1(n5303), .A2(n3025), .ZN(n5362) );
  NAND2_X1 U3750 ( .A1(n5303), .A2(n5281), .ZN(n5364) );
  INV_X1 U3751 ( .A(n3039), .ZN(n3038) );
  OAI21_X1 U3752 ( .B1(n5270), .B2(n3040), .A(n5297), .ZN(n3039) );
  NOR2_X1 U3753 ( .A1(n5301), .A2(n5300), .ZN(n5303) );
  NAND2_X1 U3754 ( .A1(n4144), .A2(n3030), .ZN(n5245) );
  AND2_X1 U3755 ( .A1(n3013), .A2(n5182), .ZN(n3030) );
  NAND2_X1 U3756 ( .A1(n4158), .A2(n4157), .ZN(n5301) );
  INV_X1 U3757 ( .A(n5244), .ZN(n4157) );
  INV_X1 U3758 ( .A(n5245), .ZN(n4158) );
  AND2_X1 U3759 ( .A1(n4144), .A2(n3013), .ZN(n5183) );
  NOR2_X1 U3760 ( .A1(n4622), .A2(n4621), .ZN(n4705) );
  NAND2_X1 U3761 ( .A1(n4130), .A2(n4129), .ZN(n4633) );
  INV_X1 U3762 ( .A(n4631), .ZN(n4130) );
  OR2_X1 U3763 ( .A1(n4633), .A2(n4558), .ZN(n4622) );
  INV_X1 U3764 ( .A(n4300), .ZN(n3052) );
  NAND2_X1 U3765 ( .A1(n3157), .A2(n3156), .ZN(n4212) );
  OAI21_X1 U3766 ( .B1(n5052), .B2(n3975), .A(n3915), .ZN(n6325) );
  NAND2_X1 U3767 ( .A1(n3317), .A2(n3316), .ZN(n3350) );
  AND3_X1 U3768 ( .A1(n3315), .A2(n3314), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3316) );
  INV_X1 U3769 ( .A(n3312), .ZN(n3351) );
  XNOR2_X1 U3770 ( .A(n3343), .B(n3342), .ZN(n4639) );
  CLKBUF_X1 U3771 ( .A(n4489), .Z(n4491) );
  AND3_X1 U3772 ( .A1(n4423), .A2(n4422), .A3(n4421), .ZN(n6507) );
  OAI21_X1 U3773 ( .B1(n5850), .B2(n5852), .A(n5849), .ZN(n5886) );
  NOR2_X1 U3774 ( .A1(n4638), .A2(n5015), .ZN(n5024) );
  OR2_X1 U3775 ( .A1(n5821), .A2(n5107), .ZN(n5015) );
  NAND2_X1 U3776 ( .A1(n5107), .A2(n4769), .ZN(n4871) );
  OR2_X1 U3777 ( .A1(n5895), .A2(n5939), .ZN(n5897) );
  AND2_X1 U3778 ( .A1(n4640), .A2(n6399), .ZN(n5901) );
  NAND2_X1 U3779 ( .A1(n3372), .A2(n3371), .ZN(n4873) );
  NAND2_X1 U3780 ( .A1(n4649), .A2(n4648), .ZN(n4719) );
  INV_X1 U3781 ( .A(n4663), .ZN(n4769) );
  AND2_X1 U3782 ( .A1(n6542), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4067) );
  AND2_X1 U3783 ( .A1(n5247), .A2(n4304), .ZN(n6145) );
  INV_X1 U3784 ( .A(n6218), .ZN(n6205) );
  INV_X1 U3785 ( .A(n6200), .ZN(n6177) );
  NOR2_X1 U3786 ( .A1(n5099), .A2(n4312), .ZN(n4313) );
  INV_X1 U3787 ( .A(n6220), .ZN(n6216) );
  INV_X1 U3788 ( .A(n5247), .ZN(n6217) );
  AND2_X1 U3789 ( .A1(n5247), .A2(n4351), .ZN(n6225) );
  AND2_X1 U3790 ( .A1(n5247), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6218) );
  INV_X1 U3791 ( .A(n6209), .ZN(n6227) );
  OAI21_X1 U3792 ( .B1(n4379), .B2(n4308), .A(n4307), .ZN(n4310) );
  OR2_X1 U3793 ( .A1(n5381), .A2(n5557), .ZN(n4297) );
  NAND2_X1 U3794 ( .A1(n4144), .A2(n4143), .ZN(n5009) );
  INV_X1 U3795 ( .A(n5988), .ZN(n6248) );
  NAND2_X1 U3796 ( .A1(n4543), .A2(n4542), .ZN(n5394) );
  AOI21_X1 U3797 ( .B1(n4541), .B2(n4540), .A(n4539), .ZN(n4542) );
  OR2_X1 U3799 ( .A1(n5413), .A2(n4267), .ZN(n4268) );
  OAI21_X1 U3800 ( .B1(n4363), .B2(n5422), .A(n5412), .ZN(n5602) );
  AND2_X1 U3801 ( .A1(n5494), .A2(n5499), .ZN(n5991) );
  INV_X1 U3802 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5982) );
  AND2_X1 U3803 ( .A1(n5531), .A2(n5543), .ZN(n6241) );
  INV_X1 U3804 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6084) );
  INV_X1 U3805 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U3806 ( .A1(n6314), .A2(n6329), .ZN(n6324) );
  INV_X1 U3807 ( .A(n6335), .ZN(n6319) );
  INV_X1 U3808 ( .A(n6314), .ZN(n6330) );
  AND2_X1 U3809 ( .A1(n5740), .A2(n4249), .ZN(n6027) );
  AND2_X1 U3810 ( .A1(n4232), .A2(n4243), .ZN(n5760) );
  NAND2_X1 U3811 ( .A1(n5563), .A2(n3028), .ZN(n5466) );
  NAND2_X1 U3812 ( .A1(n3985), .A2(n3984), .ZN(n3041) );
  CLKBUF_X1 U3813 ( .A(n4619), .Z(n4620) );
  OR2_X1 U3814 ( .A1(n4242), .A2(n6372), .ZN(n6369) );
  CLKBUF_X1 U3815 ( .A(n3924), .Z(n5826) );
  INV_X1 U3816 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6394) );
  OR2_X1 U3817 ( .A1(n4528), .A2(n4867), .ZN(n6393) );
  NOR2_X1 U3818 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6052) );
  AND2_X1 U3819 ( .A1(n5024), .A2(n5052), .ZN(n5889) );
  INV_X1 U3820 ( .A(n5194), .ZN(n5222) );
  OAI21_X1 U3821 ( .B1(n5051), .B2(n5050), .A(n5049), .ZN(n5082) );
  INV_X1 U3822 ( .A(n6460), .ZN(n6404) );
  NOR2_X1 U3823 ( .A1(n6818), .A2(n4806), .ZN(n6403) );
  NOR2_X1 U3824 ( .A1(n6777), .A2(n4806), .ZN(n6437) );
  NOR2_X2 U3825 ( .A1(n4967), .A2(n5016), .ZN(n4997) );
  OAI211_X1 U3826 ( .C1(n4776), .C2(n4775), .A(n6410), .B(n4774), .ZN(n4799)
         );
  INV_X1 U3827 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6636) );
  NOR2_X1 U3828 ( .A1(n6623), .A2(n5406), .ZN(n6534) );
  INV_X1 U3829 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6542) );
  INV_X1 U3830 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6623) );
  AND2_X1 U3831 ( .A1(n6533), .A2(n6532), .ZN(n6619) );
  INV_X1 U3832 ( .A(n4372), .ZN(n4373) );
  OAI21_X1 U3833 ( .B1(n4371), .B2(n6297), .A(n4370), .ZN(n4372) );
  AOI21_X1 U3834 ( .B1(n5707), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n4340), 
        .ZN(n4341) );
  AOI211_X1 U3835 ( .C1(n5486), .C2(n6382), .A(n4386), .B(n4385), .ZN(n4387)
         );
  NAND2_X1 U3836 ( .A1(n4001), .A2(n3009), .ZN(n4005) );
  NOR2_X1 U3837 ( .A1(n3053), .A2(n3056), .ZN(n5474) );
  NAND2_X1 U3838 ( .A1(n4353), .A2(n3011), .ZN(n5494) );
  INV_X2 U3839 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6633) );
  INV_X1 U3840 ( .A(n2999), .ZN(n5670) );
  AND2_X1 U3841 ( .A1(n5156), .A2(n3012), .ZN(n5266) );
  NAND2_X1 U3842 ( .A1(n5156), .A2(n5158), .ZN(n5157) );
  NAND2_X1 U3843 ( .A1(n3222), .A2(n4398), .ZN(n4124) );
  INV_X1 U3844 ( .A(n4124), .ZN(n5535) );
  AND2_X1 U3845 ( .A1(n3028), .A2(n3027), .ZN(n3000) );
  AND2_X1 U3846 ( .A1(n4143), .A2(n3031), .ZN(n3001) );
  AND2_X2 U3847 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4485) );
  AND4_X1 U3848 ( .A1(n3139), .A2(n3138), .A3(n3137), .A4(n3136), .ZN(n3002)
         );
  AND2_X1 U3849 ( .A1(n3045), .A2(n3046), .ZN(n5668) );
  NAND2_X1 U3850 ( .A1(n4353), .A2(n4355), .ZN(n4354) );
  AND4_X1 U3851 ( .A1(n3131), .A2(n3130), .A3(n3129), .A4(n3128), .ZN(n3003)
         );
  AND4_X1 U3852 ( .A1(n3121), .A2(n3120), .A3(n3119), .A4(n3118), .ZN(n3004)
         );
  OR2_X1 U3853 ( .A1(n5434), .A2(n6335), .ZN(n3005) );
  AND4_X1 U3854 ( .A1(n3229), .A2(n3228), .A3(n4512), .A4(n3227), .ZN(n3006)
         );
  AND2_X2 U3855 ( .A1(n3076), .A2(n4425), .ZN(n3148) );
  OR2_X1 U3856 ( .A1(n2999), .A2(n6355), .ZN(n3007) );
  AND2_X1 U3857 ( .A1(n3045), .A2(n3990), .ZN(n3008) );
  AND2_X1 U3858 ( .A1(n4002), .A2(n4000), .ZN(n3009) );
  OR2_X1 U3859 ( .A1(n4300), .A2(n4095), .ZN(n3010) );
  NOR2_X1 U3860 ( .A1(n4260), .A2(n3065), .ZN(n4084) );
  AND2_X2 U3861 ( .A1(n4488), .A2(n4425), .ZN(n3282) );
  INV_X1 U3862 ( .A(n3632), .ZN(n3870) );
  INV_X1 U3863 ( .A(n3870), .ZN(n4278) );
  NAND2_X1 U3864 ( .A1(n5563), .A2(n4177), .ZN(n5534) );
  NOR2_X2 U3865 ( .A1(n3155), .A2(n6633), .ZN(n3600) );
  INV_X1 U3866 ( .A(n3600), .ZN(n3552) );
  NAND2_X1 U3867 ( .A1(n5342), .A2(n5344), .ZN(n5343) );
  AND2_X1 U3868 ( .A1(n5156), .A2(n3059), .ZN(n5241) );
  INV_X1 U3869 ( .A(n4105), .ZN(n3156) );
  AND2_X1 U3870 ( .A1(n3788), .A2(n4355), .ZN(n3011) );
  NAND2_X1 U3871 ( .A1(n3041), .A2(n5270), .ZN(n5298) );
  INV_X2 U3872 ( .A(n5535), .ZN(n5467) );
  NAND2_X1 U3873 ( .A1(n3049), .A2(n3982), .ZN(n5257) );
  AND2_X1 U3874 ( .A1(n3059), .A2(n3537), .ZN(n3012) );
  AOI21_X1 U3875 ( .B1(n3962), .B2(n3600), .A(n3476), .ZN(n5004) );
  AND2_X1 U3876 ( .A1(n3001), .A2(n5163), .ZN(n3013) );
  NOR2_X1 U3877 ( .A1(n3471), .A2(n4277), .ZN(n3974) );
  AND2_X1 U3878 ( .A1(n3025), .A2(n3024), .ZN(n3014) );
  NAND2_X1 U3879 ( .A1(n5360), .A2(n3576), .ZN(n5342) );
  AND2_X1 U3880 ( .A1(n3046), .A2(n3993), .ZN(n3015) );
  AND2_X1 U3881 ( .A1(n3061), .A2(n4267), .ZN(n3016) );
  AND2_X1 U3882 ( .A1(n3012), .A2(n5280), .ZN(n3017) );
  OAI21_X1 U3883 ( .B1(n3957), .B2(n3552), .A(n3468), .ZN(n4725) );
  AND2_X1 U3884 ( .A1(n3000), .A2(n5525), .ZN(n3018) );
  NAND2_X1 U3885 ( .A1(n5563), .A2(n3018), .ZN(n5516) );
  AND2_X1 U3886 ( .A1(n5563), .A2(n3000), .ZN(n3019) );
  AND2_X1 U3887 ( .A1(n3011), .A2(n3058), .ZN(n3020) );
  NAND2_X1 U3888 ( .A1(n6633), .A2(n6822), .ZN(n4301) );
  INV_X1 U3889 ( .A(n4301), .ZN(n3829) );
  AND2_X1 U3890 ( .A1(n4144), .A2(n3001), .ZN(n3021) );
  AND2_X1 U3891 ( .A1(n6633), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3903) );
  AND2_X1 U3892 ( .A1(n2986), .A2(n4650), .ZN(n4112) );
  OR3_X1 U3893 ( .A1(n4209), .A2(n5491), .A3(n3035), .ZN(n3022) );
  AND2_X2 U3894 ( .A1(n3396), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4488)
         );
  AND2_X1 U3895 ( .A1(n4417), .A2(n3051), .ZN(n4111) );
  INV_X1 U3896 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6164) );
  AND2_X1 U3897 ( .A1(n4335), .A2(n3043), .ZN(n3023) );
  INV_X1 U3898 ( .A(n4378), .ZN(n3034) );
  INV_X1 U3899 ( .A(n5423), .ZN(n3035) );
  NAND2_X1 U3900 ( .A1(n3985), .A2(n3037), .ZN(n3036) );
  NAND2_X1 U3901 ( .A1(n4084), .A2(n4335), .ZN(n4259) );
  NAND2_X1 U3902 ( .A1(n3042), .A2(n4007), .ZN(n3044) );
  NAND2_X1 U3903 ( .A1(n4084), .A2(n3023), .ZN(n3042) );
  XNOR2_X1 U3904 ( .A(n3044), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5712)
         );
  CLKBUF_X1 U3905 ( .A(n5669), .Z(n3045) );
  NAND2_X1 U3906 ( .A1(n4001), .A2(n4000), .ZN(n4085) );
  NAND2_X1 U3907 ( .A1(n4005), .A2(n4004), .ZN(n4260) );
  NAND2_X1 U3908 ( .A1(n5160), .A2(n5161), .ZN(n3049) );
  NOR2_X2 U3909 ( .A1(n4724), .A2(n5004), .ZN(n5005) );
  NAND2_X1 U3910 ( .A1(n3469), .A2(n4725), .ZN(n4724) );
  NAND2_X1 U3911 ( .A1(n3399), .A2(n3398), .ZN(n4563) );
  NAND2_X2 U3912 ( .A1(n3050), .A2(n2986), .ZN(n4417) );
  INV_X1 U3913 ( .A(n4093), .ZN(n3050) );
  NAND4_X1 U3914 ( .A1(n3010), .A2(n4212), .A3(n3051), .A4(n4417), .ZN(n3197)
         );
  NAND2_X1 U3915 ( .A1(n5342), .A2(n3054), .ZN(n5549) );
  INV_X1 U3916 ( .A(n5549), .ZN(n3638) );
  AND2_X2 U3917 ( .A1(n4353), .A2(n3020), .ZN(n4364) );
  AND2_X1 U3918 ( .A1(n4363), .A2(n3061), .ZN(n5413) );
  NAND2_X1 U3919 ( .A1(n4363), .A2(n5422), .ZN(n5412) );
  NOR2_X2 U3920 ( .A1(n5644), .A2(n5645), .ZN(n5643) );
  NAND2_X1 U3921 ( .A1(n5380), .A2(n6319), .ZN(n4274) );
  NAND2_X1 U3922 ( .A1(n3237), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3218) );
  NAND2_X1 U3923 ( .A1(n3218), .A2(n3217), .ZN(n3299) );
  XNOR2_X1 U3924 ( .A(n3299), .B(n3298), .ZN(n3357) );
  NAND2_X1 U3925 ( .A1(n3299), .A2(n3297), .ZN(n3266) );
  NAND2_X1 U3926 ( .A1(n3201), .A2(n3200), .ZN(n3265) );
  CLKBUF_X1 U3927 ( .A(n3412), .Z(n3415) );
  NAND2_X1 U3928 ( .A1(n3795), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3147) );
  AND2_X1 U3929 ( .A1(n6306), .A2(n3829), .ZN(n3063) );
  AND2_X1 U3930 ( .A1(n4282), .A2(n4281), .ZN(n5504) );
  AOI21_X1 U3931 ( .B1(n6401), .B2(STATE2_REG_3__SCAN_IN), .A(n4806), .ZN(
        n5020) );
  OR2_X1 U3932 ( .A1(n5567), .A2(n4296), .ZN(n3064) );
  OR2_X1 U3933 ( .A1(n5670), .A2(n5595), .ZN(n3065) );
  INV_X1 U3934 ( .A(n5241), .ZN(n5265) );
  AND2_X1 U3935 ( .A1(n5567), .A2(n4295), .ZN(n5569) );
  AND4_X1 U3936 ( .A1(n3126), .A2(n3125), .A3(n3124), .A4(n3123), .ZN(n3066)
         );
  INV_X1 U3937 ( .A(n6236), .ZN(n4283) );
  OR2_X1 U3938 ( .A1(n4409), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3067)
         );
  NAND2_X1 U3939 ( .A1(n5812), .A2(n5811), .ZN(n5810) );
  AND2_X1 U3940 ( .A1(n3225), .A2(n5391), .ZN(n3068) );
  OR2_X1 U3941 ( .A1(n4534), .A2(n6521), .ZN(n6297) );
  NAND2_X1 U3942 ( .A1(n3187), .A2(n3225), .ZN(n3189) );
  INV_X1 U3943 ( .A(n3947), .ZN(n3435) );
  AND2_X1 U3944 ( .A1(n3862), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3127) );
  AOI22_X1 U3945 ( .A1(n3163), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3148), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3151) );
  INV_X1 U3946 ( .A(n4010), .ZN(n3260) );
  NAND2_X1 U3947 ( .A1(n3209), .A2(n3194), .ZN(n3185) );
  INV_X1 U3948 ( .A(n3964), .ZN(n3457) );
  INV_X1 U3949 ( .A(n3378), .ZN(n4486) );
  AOI21_X1 U3950 ( .B1(n3565), .B2(INSTQUEUE_REG_12__3__SCAN_IN), .A(n3127), 
        .ZN(n3130) );
  AND2_X1 U3951 ( .A1(n6401), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4024)
         );
  OR2_X1 U3952 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n4055), .ZN(n4047)
         );
  INV_X1 U3953 ( .A(n5523), .ZN(n3702) );
  OR2_X1 U3954 ( .A1(n2999), .A2(n3994), .ZN(n3995) );
  OR2_X1 U3955 ( .A1(n3384), .A2(n3383), .ZN(n3909) );
  AND2_X1 U3956 ( .A1(n4048), .A2(n4047), .ZN(n4098) );
  INV_X1 U3957 ( .A(n5551), .ZN(n3637) );
  INV_X1 U3958 ( .A(n4630), .ZN(n4129) );
  INV_X1 U3959 ( .A(n3831), .ZN(n4365) );
  NOR2_X1 U3960 ( .A1(n3444), .A2(n3063), .ZN(n3445) );
  INV_X1 U3961 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4506) );
  NAND2_X1 U3962 ( .A1(n4056), .A2(n4055), .ZN(n4100) );
  AND2_X1 U3963 ( .A1(n5553), .A2(n5562), .ZN(n4177) );
  AND2_X1 U3964 ( .A1(n4181), .A2(n5536), .ZN(n5465) );
  AND2_X1 U3965 ( .A1(n4168), .A2(n4167), .ZN(n5346) );
  AOI22_X1 U3966 ( .A1(n3107), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        INSTQUEUE_REG_13__1__SCAN_IN), .B2(n3283), .ZN(n3075) );
  AND2_X1 U3967 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3705), .ZN(n3706)
         );
  INV_X1 U3968 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5614) );
  AND2_X1 U3969 ( .A1(n4839), .A2(n6408), .ZN(n4842) );
  NAND2_X1 U3970 ( .A1(n3367), .A2(n3366), .ZN(n4522) );
  AND2_X1 U3971 ( .A1(n4191), .A2(n4190), .ZN(n5517) );
  NOR2_X1 U3972 ( .A1(n3549), .A2(n3548), .ZN(n3554) );
  NAND2_X1 U3973 ( .A1(n3417), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3442)
         );
  AND2_X1 U3974 ( .A1(n4156), .A2(n4155), .ZN(n5244) );
  INV_X1 U3975 ( .A(n6284), .ZN(n6529) );
  AND2_X1 U3976 ( .A1(n3706), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3761)
         );
  NAND2_X1 U3977 ( .A1(n3492), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3506)
         );
  NOR2_X1 U3978 ( .A1(n3464), .A2(n6164), .ZN(n3473) );
  AND2_X1 U3979 ( .A1(n2999), .A2(n5759), .ZN(n5616) );
  AND2_X1 U3980 ( .A1(n4142), .A2(n4141), .ZN(n4740) );
  INV_X1 U3981 ( .A(n6382), .ZN(n6339) );
  NAND2_X1 U3982 ( .A1(n4235), .A2(n4226), .ZN(n5796) );
  INV_X1 U3983 ( .A(n5826), .ZN(n5107) );
  OR2_X1 U3984 ( .A1(n4871), .A2(n5821), .ZN(n5053) );
  OR2_X1 U3985 ( .A1(n4871), .A2(n4869), .ZN(n6450) );
  OR2_X1 U3986 ( .A1(n5105), .A2(n5821), .ZN(n4845) );
  INV_X1 U3987 ( .A(n5887), .ZN(n4731) );
  OR3_X1 U3988 ( .A1(n5402), .A2(n6545), .A3(n5400), .ZN(n4393) );
  NOR2_X1 U3989 ( .A1(n6592), .A2(n5352), .ZN(n6104) );
  OR2_X1 U3990 ( .A1(n6638), .A2(n4303), .ZN(n5247) );
  NAND2_X1 U3991 ( .A1(n3443), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3464)
         );
  NAND2_X1 U3992 ( .A1(n4347), .A2(n4346), .ZN(n6220) );
  NAND2_X1 U3993 ( .A1(n4368), .A2(n4367), .ZN(n5434) );
  AND2_X1 U3994 ( .A1(n5394), .A2(n5393), .ZN(n6251) );
  INV_X1 U3995 ( .A(n4543), .ZN(n6288) );
  NAND2_X1 U3996 ( .A1(n3808), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3832)
         );
  AND2_X1 U3997 ( .A1(n5513), .A2(n5524), .ZN(n5997) );
  INV_X1 U3998 ( .A(n6324), .ZN(n6310) );
  OR2_X1 U3999 ( .A1(n5406), .A2(n6545), .ZN(n4534) );
  INV_X1 U4000 ( .A(n6297), .ZN(n6332) );
  BUF_X1 U4001 ( .A(n5626), .Z(n5653) );
  NAND2_X1 U4002 ( .A1(n4110), .A2(n4109), .ZN(n4235) );
  INV_X1 U4003 ( .A(n5796), .ZN(n6372) );
  INV_X1 U4004 ( .A(n4806), .ZN(n4867) );
  INV_X1 U4005 ( .A(n6534), .ZN(n5838) );
  AND2_X1 U4006 ( .A1(n5107), .A2(n4665), .ZN(n5887) );
  INV_X1 U4007 ( .A(n5052), .ZN(n5016) );
  INV_X1 U4008 ( .A(n5193), .ZN(n5220) );
  INV_X1 U4009 ( .A(n4877), .ZN(n5149) );
  NOR2_X1 U4010 ( .A1(n5053), .A2(n5052), .ZN(n6445) );
  AND2_X1 U4011 ( .A1(n5821), .A2(n5052), .ZN(n5117) );
  OR2_X1 U4012 ( .A1(n4922), .A2(n4921), .ZN(n4956) );
  NOR2_X2 U4013 ( .A1(n4845), .A2(n5052), .ZN(n5939) );
  NAND2_X1 U4014 ( .A1(n4638), .A2(n5826), .ZN(n5105) );
  INV_X1 U4015 ( .A(n6408), .ZN(n5896) );
  INV_X1 U4016 ( .A(n4777), .ZN(n4998) );
  OR4_X1 U4017 ( .A1(n6528), .A2(n6527), .A3(n6526), .A4(n6525), .ZN(n6538) );
  NOR2_X1 U4018 ( .A1(n6542), .A2(n6633), .ZN(n4529) );
  INV_X1 U4019 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6564) );
  INV_X1 U4020 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6569) );
  OR2_X1 U4021 ( .A1(n4534), .A2(n5398), .ZN(n4395) );
  AND2_X1 U4022 ( .A1(n6564), .A2(STATE_REG_1__SCAN_IN), .ZN(n6836) );
  INV_X1 U4023 ( .A(n6145), .ZN(n6167) );
  INV_X1 U4024 ( .A(n6225), .ZN(n6206) );
  OR2_X1 U4025 ( .A1(n4117), .A2(n6232), .ZN(n6200) );
  AND2_X1 U4026 ( .A1(n4297), .A2(n3064), .ZN(n4298) );
  NAND2_X1 U4027 ( .A1(n5394), .A2(n4545), .ZN(n5988) );
  OR2_X1 U4028 ( .A1(n4534), .A2(n4470), .ZN(n6286) );
  OR2_X1 U4029 ( .A1(n4534), .A2(n6531), .ZN(n6291) );
  NAND2_X1 U4030 ( .A1(n6297), .A2(n4071), .ZN(n6314) );
  AOI21_X1 U4031 ( .B1(n4256), .B2(n6382), .A(n4255), .ZN(n4257) );
  NAND2_X1 U4032 ( .A1(n4235), .A2(n4115), .ZN(n6035) );
  INV_X1 U4033 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U4034 ( .A1(n5024), .A2(n5016), .ZN(n5194) );
  AOI21_X1 U4035 ( .B1(n5192), .B2(n5191), .A(n5190), .ZN(n5226) );
  AOI211_X2 U4036 ( .C1(n5114), .C2(n5115), .A(n5113), .B(n5112), .ZN(n5155)
         );
  AND2_X1 U4037 ( .A1(n4876), .A2(n4875), .ZN(n4906) );
  NAND2_X1 U4038 ( .A1(n4748), .A2(n5117), .ZN(n6460) );
  NAND2_X1 U4039 ( .A1(n4837), .A2(n5052), .ZN(n4963) );
  AOI22_X1 U4040 ( .A1(n5904), .A2(n5901), .B1(n6396), .B2(n5899), .ZN(n5942)
         );
  OR2_X1 U4041 ( .A1(n5105), .A2(n4646), .ZN(n6500) );
  AOI21_X1 U4042 ( .B1(n4809), .B2(n4808), .A(n4807), .ZN(n4836) );
  INV_X1 U4043 ( .A(n6403), .ZN(n5910) );
  INV_X1 U4044 ( .A(n6437), .ZN(n5934) );
  INV_X1 U4045 ( .A(n6618), .ZN(n6552) );
  INV_X1 U4046 ( .A(n6609), .ZN(n6614) );
  NAND2_X1 U4047 ( .A1(n3005), .A2(n4373), .ZN(U2959) );
  NAND2_X1 U4048 ( .A1(n4388), .A2(n4387), .ZN(U2989) );
  NAND2_X1 U4049 ( .A1(n4258), .A2(n4257), .ZN(U2991) );
  NOR2_X4 U4050 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3076) );
  NOR2_X4 U4051 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4520) );
  AND2_X2 U4052 ( .A1(n3076), .A2(n4520), .ZN(n3107) );
  INV_X1 U4053 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3069) );
  AND2_X2 U4054 ( .A1(n4488), .A2(n4520), .ZN(n3141) );
  AOI22_X1 U4055 ( .A1(n3245), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3141), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3074) );
  AND2_X2 U4056 ( .A1(n3076), .A2(n4484), .ZN(n3168) );
  AOI22_X1 U4057 ( .A1(n3273), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3168), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3073) );
  INV_X1 U4058 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3071) );
  AND2_X4 U4059 ( .A1(n3071), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4424)
         );
  AND2_X4 U4060 ( .A1(n4424), .A2(n4488), .ZN(n3878) );
  AOI22_X1 U4061 ( .A1(n3878), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3072) );
  NAND4_X1 U4062 ( .A1(n3075), .A2(n3074), .A3(n3073), .A4(n3072), .ZN(n3082)
         );
  NAND2_X2 U4063 ( .A1(n4424), .A2(n4485), .ZN(n3250) );
  INV_X2 U4064 ( .A(n3250), .ZN(n3163) );
  AND2_X4 U4065 ( .A1(n3076), .A2(n4424), .ZN(n3795) );
  AOI22_X1 U4066 ( .A1(n3251), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3079) );
  AOI22_X1 U4067 ( .A1(n3862), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3565), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3078) );
  AND2_X4 U4068 ( .A1(n4520), .A2(n4489), .ZN(n3845) );
  AND2_X2 U4069 ( .A1(n4484), .A2(n4485), .ZN(n3566) );
  AOI22_X1 U4070 ( .A1(n3845), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3566), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3077) );
  NAND4_X1 U4071 ( .A1(n3080), .A2(n3079), .A3(n3078), .A4(n3077), .ZN(n3081)
         );
  NAND2_X1 U4072 ( .A1(n3282), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3086) );
  NAND2_X1 U4073 ( .A1(n3878), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3085) );
  NAND2_X1 U4074 ( .A1(n3273), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3084) );
  NAND2_X1 U4075 ( .A1(n3168), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3083) );
  NAND2_X1 U4076 ( .A1(n3245), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3090) );
  BUF_X4 U4077 ( .A(n3141), .Z(n3887) );
  NAND2_X1 U4078 ( .A1(n3887), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3089) );
  NAND2_X1 U4079 ( .A1(n3283), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3088)
         );
  NAND2_X1 U4080 ( .A1(n3107), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3087) );
  NAND2_X1 U4081 ( .A1(n3148), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3094) );
  NAND2_X1 U4082 ( .A1(n3862), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3093)
         );
  NAND2_X1 U4083 ( .A1(n3163), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3092)
         );
  NAND2_X1 U4084 ( .A1(n3565), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3091)
         );
  NAND2_X1 U4085 ( .A1(n3251), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3098)
         );
  NAND2_X1 U4086 ( .A1(n3795), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3097) );
  NAND2_X1 U4087 ( .A1(n3888), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3096) );
  NAND2_X1 U4088 ( .A1(n3566), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3095)
         );
  AND4_X4 U4089 ( .A1(n3102), .A2(n3101), .A3(n3100), .A4(n3099), .ZN(n4650)
         );
  AOI22_X1 U4090 ( .A1(n3862), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3106) );
  AOI22_X1 U4091 ( .A1(n3565), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3148), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3105) );
  AOI22_X1 U4092 ( .A1(n3282), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3168), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3104) );
  AOI22_X1 U4093 ( .A1(n3245), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3103) );
  AOI22_X1 U4094 ( .A1(n3283), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3107), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3110) );
  AOI22_X1 U4095 ( .A1(n3878), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3141), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3109) );
  AOI22_X1 U4096 ( .A1(n3845), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3566), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3108) );
  AOI22_X1 U4097 ( .A1(n3878), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3141), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3117) );
  AOI22_X1 U4098 ( .A1(n3148), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3107), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3116) );
  AOI22_X1 U4099 ( .A1(n3251), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3565), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3115) );
  AOI22_X1 U4100 ( .A1(n3845), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3566), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3114) );
  AOI22_X1 U4101 ( .A1(n3245), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3121) );
  AOI22_X1 U4102 ( .A1(n3283), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3163), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3120) );
  AOI22_X1 U4103 ( .A1(n3862), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3119) );
  AOI22_X1 U4104 ( .A1(n3282), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3168), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3118) );
  AOI22_X1 U4105 ( .A1(n3878), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3126) );
  AOI22_X1 U4106 ( .A1(n3245), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3887), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3125) );
  AOI22_X1 U4107 ( .A1(n3273), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3168), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3124) );
  AOI22_X1 U4108 ( .A1(n3283), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3107), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3123) );
  AOI22_X1 U4109 ( .A1(n3251), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3131) );
  AOI22_X1 U4110 ( .A1(n3163), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3148), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3129) );
  AOI22_X1 U4111 ( .A1(n3845), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3566), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3128) );
  NAND2_X2 U4112 ( .A1(n3066), .A2(n3003), .ZN(n3222) );
  NOR2_X1 U4113 ( .A1(n4222), .A2(n3222), .ZN(n4279) );
  NAND3_X1 U4114 ( .A1(n4112), .A2(n5392), .A3(n4279), .ZN(n4428) );
  INV_X1 U4115 ( .A(n4428), .ZN(n3157) );
  AOI22_X1 U4116 ( .A1(n3163), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3148), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3135) );
  AOI22_X1 U4117 ( .A1(n3251), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3134) );
  AOI22_X1 U4118 ( .A1(n3862), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3565), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3133) );
  AOI22_X1 U4119 ( .A1(n3845), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3566), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3132) );
  AOI22_X1 U4120 ( .A1(n3245), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3141), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3139) );
  AOI22_X1 U4121 ( .A1(n3283), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3107), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3138) );
  AOI22_X1 U4122 ( .A1(n3273), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3168), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3137) );
  AOI22_X1 U4123 ( .A1(n3878), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3136) );
  NAND2_X4 U4124 ( .A1(n3140), .A2(n3002), .ZN(n5391) );
  AOI22_X1 U4125 ( .A1(n3878), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3144) );
  AOI22_X1 U4126 ( .A1(n3845), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3566), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3143) );
  AOI22_X1 U4127 ( .A1(n3245), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3141), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3142) );
  AOI22_X1 U4128 ( .A1(n3282), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3168), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3150) );
  AOI22_X1 U4129 ( .A1(n3862), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3565), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3149) );
  NAND2_X2 U4130 ( .A1(n3154), .A2(n3153), .ZN(n3183) );
  NAND2_X1 U4131 ( .A1(n5391), .A2(n3155), .ZN(n4105) );
  NAND2_X1 U4132 ( .A1(n3148), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3162) );
  NAND2_X1 U4133 ( .A1(n3845), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3161) );
  NAND2_X1 U4134 ( .A1(n3565), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3160)
         );
  NAND2_X1 U4135 ( .A1(n3566), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3159)
         );
  NAND2_X1 U4136 ( .A1(n3141), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3167) );
  NAND2_X1 U4137 ( .A1(n3282), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3166) );
  NAND2_X1 U4138 ( .A1(n3163), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3165)
         );
  NAND2_X1 U4139 ( .A1(n3107), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3164) );
  NAND2_X1 U4140 ( .A1(n3245), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3171) );
  NAND2_X1 U4141 ( .A1(n3273), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3170) );
  NAND2_X1 U4142 ( .A1(n3168), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3169) );
  NAND2_X1 U4143 ( .A1(n3862), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3176)
         );
  NAND2_X1 U4144 ( .A1(n3283), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3175)
         );
  NAND2_X1 U4145 ( .A1(n3251), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3174)
         );
  NAND2_X1 U4146 ( .A1(n3795), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3173) );
  NOR2_X2 U4147 ( .A1(n3185), .A2(n4295), .ZN(n4091) );
  NAND2_X1 U4148 ( .A1(n3181), .A2(n4091), .ZN(n4104) );
  INV_X1 U4149 ( .A(n4104), .ZN(n3182) );
  NAND2_X1 U4150 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .ZN(
        n6567) );
  OAI21_X1 U4151 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_1__SCAN_IN), .A(
        n6567), .ZN(n4095) );
  INV_X2 U4152 ( .A(n3183), .ZN(n3225) );
  INV_X1 U4153 ( .A(n3222), .ZN(n4672) );
  NAND2_X1 U4154 ( .A1(n3185), .A2(n4222), .ZN(n3186) );
  OAI211_X1 U4155 ( .C1(n3221), .C2(n4672), .A(n3186), .B(n5391), .ZN(n3193)
         );
  INV_X1 U4156 ( .A(n2997), .ZN(n3191) );
  NAND2_X1 U4157 ( .A1(n4222), .A2(n3183), .ZN(n3188) );
  NAND2_X1 U4158 ( .A1(n3189), .A2(n3188), .ZN(n3190) );
  NOR2_X1 U4159 ( .A1(n3191), .A2(n3190), .ZN(n3192) );
  NOR2_X1 U4160 ( .A1(n3193), .A2(n3192), .ZN(n3202) );
  NOR2_X1 U4161 ( .A1(n4069), .A2(n2987), .ZN(n3196) );
  NAND2_X1 U4162 ( .A1(n3202), .A2(n3196), .ZN(n4093) );
  NAND2_X1 U4163 ( .A1(n3197), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3235) );
  INV_X1 U4164 ( .A(n3235), .ZN(n3201) );
  NAND2_X1 U4165 ( .A1(n6052), .A2(n6636), .ZN(n4077) );
  INV_X1 U4166 ( .A(n4077), .ZN(n3242) );
  XNOR2_X1 U4167 ( .A(n6401), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6396)
         );
  NAND2_X1 U4168 ( .A1(n3242), .A2(n6396), .ZN(n3199) );
  INV_X1 U4169 ( .A(n4067), .ZN(n3241) );
  NAND2_X1 U4170 ( .A1(n3241), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3198) );
  NAND2_X1 U4171 ( .A1(n3199), .A2(n3198), .ZN(n3233) );
  OR2_X1 U4172 ( .A1(n3233), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3200)
         );
  INV_X1 U4173 ( .A(n3202), .ZN(n3230) );
  NAND2_X1 U4174 ( .A1(n3230), .A2(n4650), .ZN(n3215) );
  INV_X1 U4175 ( .A(n4091), .ZN(n3203) );
  NAND2_X1 U4176 ( .A1(n3203), .A2(n3908), .ZN(n3205) );
  AND2_X2 U4178 ( .A1(n3205), .A2(n3204), .ZN(n3227) );
  NAND2_X1 U4179 ( .A1(n4650), .A2(n4398), .ZN(n5100) );
  INV_X1 U4180 ( .A(n4095), .ZN(n3206) );
  OAI21_X1 U4181 ( .B1(n4398), .B2(n3206), .A(n5392), .ZN(n3208) );
  AND2_X1 U4182 ( .A1(n5391), .A2(n3222), .ZN(n3210) );
  NAND2_X1 U4184 ( .A1(n4544), .A2(n3212), .ZN(n3213) );
  AND2_X2 U4185 ( .A1(n4216), .A2(n3213), .ZN(n3219) );
  NAND4_X1 U4186 ( .A1(n3215), .A2(n3227), .A3(n3214), .A4(n3219), .ZN(n3216)
         );
  AND2_X2 U4187 ( .A1(n3216), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3237) );
  MUX2_X1 U4188 ( .A(n4067), .B(n4077), .S(n6401), .Z(n3217) );
  INV_X1 U4189 ( .A(n3219), .ZN(n3220) );
  NAND2_X1 U4190 ( .A1(n3220), .A2(n4398), .ZN(n3229) );
  NAND2_X1 U4191 ( .A1(n3908), .A2(n5374), .ZN(n3224) );
  NAND2_X1 U4192 ( .A1(n6052), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6544) );
  INV_X1 U4193 ( .A(n6544), .ZN(n3223) );
  NAND2_X1 U4194 ( .A1(n2987), .A2(n4222), .ZN(n4215) );
  AND4_X1 U4195 ( .A1(n3224), .A2(n3223), .A3(n2985), .A4(n4215), .ZN(n3228)
         );
  AND3_X1 U4196 ( .A1(n3225), .A2(n3212), .A3(n5391), .ZN(n3226) );
  NAND2_X1 U4197 ( .A1(n4279), .A2(n3226), .ZN(n4512) );
  AND2_X1 U4199 ( .A1(n4069), .A2(n4398), .ZN(n3231) );
  NAND2_X1 U4200 ( .A1(n3006), .A2(n4220), .ZN(n3297) );
  NAND2_X1 U4201 ( .A1(n3265), .A2(n3266), .ZN(n3236) );
  AOI21_X1 U4202 ( .B1(n3237), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3233), 
        .ZN(n3234) );
  NAND2_X1 U4203 ( .A1(n3235), .A2(n3234), .ZN(n3264) );
  NAND2_X1 U4204 ( .A1(n3237), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3244) );
  AND2_X1 U4205 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3238) );
  NAND2_X1 U4206 ( .A1(n3238), .A2(n6512), .ZN(n5110) );
  INV_X1 U4207 ( .A(n3238), .ZN(n3239) );
  NAND2_X1 U4208 ( .A1(n3239), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3240) );
  NAND2_X1 U4209 ( .A1(n5110), .A2(n3240), .ZN(n4772) );
  AOI22_X1 U4210 ( .A1(n3242), .A2(n4772), .B1(n3241), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3243) );
  XNOR2_X1 U4211 ( .A(n3365), .B(n3366), .ZN(n4503) );
  NAND2_X1 U4212 ( .A1(n4503), .A2(n6636), .ZN(n3259) );
  INV_X1 U4213 ( .A(n4277), .ZN(n3294) );
  AOI22_X1 U4214 ( .A1(n3818), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3249) );
  INV_X1 U4215 ( .A(n3245), .ZN(n4493) );
  AOI22_X1 U4216 ( .A1(n3886), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3248) );
  AOI22_X1 U4217 ( .A1(n3880), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3247) );
  AOI22_X1 U4218 ( .A1(n3879), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3246) );
  NAND4_X1 U4219 ( .A1(n3249), .A2(n3248), .A3(n3247), .A4(n3246), .ZN(n3257)
         );
  AOI22_X1 U4220 ( .A1(n3774), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3255) );
  INV_X1 U4221 ( .A(n3251), .ZN(n3378) );
  AOI22_X1 U4222 ( .A1(n4486), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3254) );
  AOI22_X1 U4223 ( .A1(n3813), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4224 ( .A1(n3888), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3252) );
  NAND4_X1 U4225 ( .A1(n3255), .A2(n3254), .A3(n3253), .A4(n3252), .ZN(n3256)
         );
  NAND2_X1 U4226 ( .A1(n3294), .A2(n3907), .ZN(n3258) );
  NAND2_X1 U4227 ( .A1(n4650), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3373) );
  INV_X1 U4228 ( .A(n3373), .ZN(n3261) );
  NAND2_X1 U4229 ( .A1(n3265), .A2(n3264), .ZN(n3268) );
  INV_X1 U4230 ( .A(n3266), .ZN(n3267) );
  XNOR2_X1 U4231 ( .A(n3268), .B(n3267), .ZN(n4426) );
  NAND2_X1 U4232 ( .A1(n4426), .A2(n6636), .ZN(n3281) );
  AOI22_X1 U4233 ( .A1(n3818), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3272) );
  AOI22_X1 U4234 ( .A1(n3886), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3271) );
  AOI22_X1 U4235 ( .A1(n2996), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3888), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3270) );
  AOI22_X1 U4236 ( .A1(n3819), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3269) );
  NAND4_X1 U4237 ( .A1(n3272), .A2(n3271), .A3(n3270), .A4(n3269), .ZN(n3279)
         );
  AOI22_X1 U4238 ( .A1(n3879), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U4239 ( .A1(n3880), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3276) );
  AOI22_X1 U4240 ( .A1(n3813), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3275) );
  AOI22_X1 U4241 ( .A1(n3881), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3274) );
  NAND4_X1 U4242 ( .A1(n3277), .A2(n3276), .A3(n3275), .A4(n3274), .ZN(n3278)
         );
  NAND2_X1 U4243 ( .A1(n3294), .A2(n3916), .ZN(n3280) );
  INV_X1 U4244 ( .A(n3916), .ZN(n3296) );
  NAND2_X1 U4245 ( .A1(n4022), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3295) );
  AOI22_X1 U4246 ( .A1(n3818), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4247 ( .A1(n3886), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4248 ( .A1(n3273), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4249 ( .A1(n3879), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3284) );
  NAND4_X1 U4250 ( .A1(n3287), .A2(n3286), .A3(n3285), .A4(n3284), .ZN(n3293)
         );
  AOI22_X1 U4251 ( .A1(n3774), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4252 ( .A1(n3251), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3290) );
  AOI22_X1 U4253 ( .A1(n3813), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3289) );
  AOI22_X1 U4254 ( .A1(n3845), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3288) );
  NAND4_X1 U4255 ( .A1(n3291), .A2(n3290), .A3(n3289), .A4(n3288), .ZN(n3292)
         );
  INV_X1 U4256 ( .A(n3977), .ZN(n3471) );
  NAND2_X1 U4257 ( .A1(n3294), .A2(n3471), .ZN(n3300) );
  NAND2_X1 U4258 ( .A1(n3341), .A2(n3339), .ZN(n3322) );
  NAND2_X1 U4259 ( .A1(n3357), .A2(n6636), .ZN(n3348) );
  INV_X1 U4260 ( .A(n3300), .ZN(n3311) );
  AOI22_X1 U4261 ( .A1(n3886), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3304) );
  AOI22_X1 U4262 ( .A1(n3813), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U4263 ( .A1(n3774), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4264 ( .A1(n2996), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3301) );
  NAND4_X1 U4265 ( .A1(n3304), .A2(n3303), .A3(n3302), .A4(n3301), .ZN(n3310)
         );
  AOI22_X1 U4266 ( .A1(n3818), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4267 ( .A1(n3819), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3888), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U4268 ( .A1(n3879), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4269 ( .A1(n3273), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3305) );
  NAND4_X1 U4270 ( .A1(n3308), .A2(n3307), .A3(n3306), .A4(n3305), .ZN(n3309)
         );
  MUX2_X1 U4271 ( .A(n3974), .B(n3311), .S(n3917), .Z(n3312) );
  NAND2_X1 U4272 ( .A1(n3348), .A2(n3351), .ZN(n3318) );
  NAND2_X1 U4273 ( .A1(n4022), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3317) );
  NAND2_X1 U4274 ( .A1(n4650), .A2(n3917), .ZN(n3315) );
  NAND2_X1 U4275 ( .A1(n3313), .A2(n3977), .ZN(n3314) );
  NAND2_X1 U4276 ( .A1(n3318), .A2(n3350), .ZN(n3320) );
  INV_X1 U4277 ( .A(n3974), .ZN(n3319) );
  INV_X1 U4278 ( .A(n3340), .ZN(n3321) );
  NAND2_X1 U4279 ( .A1(n3322), .A2(n3321), .ZN(n3326) );
  INV_X1 U4280 ( .A(n3341), .ZN(n3324) );
  INV_X1 U4281 ( .A(n3339), .ZN(n3323) );
  NAND2_X1 U4282 ( .A1(n3324), .A2(n3323), .ZN(n3325) );
  AND2_X2 U4283 ( .A1(n3326), .A2(n3325), .ZN(n3327) );
  OAI21_X1 U4284 ( .B1(n3328), .B2(n3327), .A(n3387), .ZN(n3924) );
  INV_X1 U4285 ( .A(n3924), .ZN(n3329) );
  NAND2_X1 U4286 ( .A1(n3329), .A2(n3600), .ZN(n3330) );
  NAND2_X1 U4287 ( .A1(n3330), .A2(n3762), .ZN(n3338) );
  INV_X1 U4288 ( .A(n3338), .ZN(n3335) );
  NAND2_X1 U4289 ( .A1(n3356), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3334) );
  NOR2_X2 U4290 ( .A1(n5391), .A2(n6633), .ZN(n3632) );
  OAI21_X1 U4291 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3391), .ZN(n6323) );
  INV_X1 U4292 ( .A(n6323), .ZN(n3331) );
  INV_X1 U4293 ( .A(n3903), .ZN(n3762) );
  INV_X1 U4294 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6204) );
  OAI22_X1 U4295 ( .A1(n4301), .A2(n3331), .B1(n3762), .B2(n6204), .ZN(n3332)
         );
  AOI21_X1 U4296 ( .B1(n4278), .B2(EAX_REG_2__SCAN_IN), .A(n3332), .ZN(n3333)
         );
  AND2_X1 U4297 ( .A1(n3334), .A2(n3333), .ZN(n3336) );
  NAND2_X1 U4298 ( .A1(n3335), .A2(n3336), .ZN(n4628) );
  INV_X1 U4299 ( .A(n3336), .ZN(n3337) );
  NAND2_X1 U4300 ( .A1(n3338), .A2(n3337), .ZN(n3363) );
  XNOR2_X1 U4301 ( .A(n3340), .B(n3339), .ZN(n3343) );
  NAND2_X1 U4302 ( .A1(n4639), .A2(n3600), .ZN(n3347) );
  AOI22_X1 U4303 ( .A1(n4278), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6633), .ZN(n3345) );
  NAND2_X1 U4304 ( .A1(n3356), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3344) );
  AND2_X1 U4305 ( .A1(n3345), .A2(n3344), .ZN(n3346) );
  NAND2_X1 U4306 ( .A1(n3347), .A2(n3346), .ZN(n4441) );
  NAND2_X1 U4307 ( .A1(n3348), .A2(n3350), .ZN(n3349) );
  NAND2_X1 U4308 ( .A1(n3349), .A2(n3351), .ZN(n3354) );
  INV_X1 U4309 ( .A(n3350), .ZN(n3352) );
  NAND2_X1 U4310 ( .A1(n5052), .A2(n3068), .ZN(n3355) );
  NAND2_X1 U4311 ( .A1(n3355), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4410) );
  INV_X1 U4312 ( .A(n3356), .ZN(n3420) );
  INV_X1 U4313 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U4314 ( .A1(n3358), .A2(n3600), .ZN(n3360) );
  AOI22_X1 U4315 ( .A1(n3632), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6633), .ZN(n3359) );
  OAI211_X1 U4316 ( .C1(n3420), .C2(n6503), .A(n3360), .B(n3359), .ZN(n4411)
         );
  NAND2_X1 U4317 ( .A1(n4410), .A2(n4411), .ZN(n3362) );
  NAND2_X1 U4318 ( .A1(n4441), .A2(n4440), .ZN(n4439) );
  NAND2_X1 U4319 ( .A1(n3363), .A2(n4439), .ZN(n3364) );
  INV_X1 U4320 ( .A(n4564), .ZN(n3399) );
  INV_X1 U4321 ( .A(n3365), .ZN(n3367) );
  NAND2_X1 U4322 ( .A1(n3237), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3372) );
  NAND3_X1 U4323 ( .A1(n6517), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4745) );
  INV_X1 U4324 ( .A(n4745), .ZN(n3368) );
  NAND2_X1 U4325 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3368), .ZN(n6451) );
  NAND2_X1 U4326 ( .A1(n6517), .A2(n6451), .ZN(n3369) );
  NOR3_X1 U4327 ( .A1(n6517), .A2(n6512), .A3(n5018), .ZN(n4773) );
  NAND2_X1 U4328 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4773), .ZN(n4732) );
  NAND2_X1 U4329 ( .A1(n3369), .A2(n4732), .ZN(n4865) );
  OAI22_X1 U4330 ( .A1(n4077), .A2(n4865), .B1(n4067), .B2(n6517), .ZN(n3370)
         );
  INV_X1 U4331 ( .A(n3370), .ZN(n3371) );
  AOI22_X1 U4332 ( .A1(n3818), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3377) );
  INV_X2 U4333 ( .A(n4493), .ZN(n3886) );
  AOI22_X1 U4334 ( .A1(n3886), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4335 ( .A1(n3880), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U4336 ( .A1(n3879), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3374) );
  NAND4_X1 U4337 ( .A1(n3377), .A2(n3376), .A3(n3375), .A4(n3374), .ZN(n3384)
         );
  AOI22_X1 U4338 ( .A1(n3774), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4339 ( .A1(n4486), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4340 ( .A1(n3813), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3380) );
  AOI22_X1 U4341 ( .A1(n3857), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3379) );
  NAND4_X1 U4342 ( .A1(n3382), .A2(n3381), .A3(n3380), .A4(n3379), .ZN(n3383)
         );
  AOI22_X1 U4343 ( .A1(n4035), .A2(n3909), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n4022), .ZN(n3385) );
  NAND2_X1 U4344 ( .A1(n3387), .A2(n4769), .ZN(n3389) );
  INV_X1 U4345 ( .A(n3387), .ZN(n3388) );
  NAND2_X1 U4346 ( .A1(n3388), .A2(n4663), .ZN(n3412) );
  INV_X1 U4347 ( .A(n3391), .ZN(n3393) );
  INV_X1 U4348 ( .A(n3417), .ZN(n3392) );
  OAI21_X1 U4349 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3393), .A(n3392), 
        .ZN(n5236) );
  AOI22_X1 U4350 ( .A1(n3829), .A2(n5236), .B1(n3903), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3395) );
  NAND2_X1 U4351 ( .A1(n4278), .A2(EAX_REG_3__SCAN_IN), .ZN(n3394) );
  OAI211_X1 U4352 ( .C1(n3420), .C2(n3396), .A(n3395), .B(n3394), .ZN(n3397)
         );
  AOI21_X1 U4353 ( .B1(n4637), .B2(n3600), .A(n3397), .ZN(n4565) );
  INV_X1 U4354 ( .A(n3412), .ZN(n3411) );
  AOI22_X1 U4355 ( .A1(n3818), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4356 ( .A1(n3886), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3402) );
  AOI22_X1 U4357 ( .A1(n3880), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3401) );
  AOI22_X1 U4358 ( .A1(n3879), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3400) );
  NAND4_X1 U4359 ( .A1(n3403), .A2(n3402), .A3(n3401), .A4(n3400), .ZN(n3409)
         );
  AOI22_X1 U4360 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n3819), .B1(n3774), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3407) );
  AOI22_X1 U4361 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n3881), .B1(n4486), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3406) );
  AOI22_X1 U4362 ( .A1(n3813), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4363 ( .A1(n3857), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3404) );
  NAND4_X1 U4364 ( .A1(n3407), .A2(n3406), .A3(n3405), .A4(n3404), .ZN(n3408)
         );
  NAND2_X1 U4365 ( .A1(n4022), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3410) );
  NAND2_X1 U4366 ( .A1(n3411), .A2(n3413), .ZN(n3437) );
  INV_X1 U4367 ( .A(n3413), .ZN(n3414) );
  NAND2_X1 U4368 ( .A1(n3415), .A2(n3414), .ZN(n3416) );
  AND2_X2 U4369 ( .A1(n3437), .A2(n3416), .ZN(n3937) );
  OAI21_X1 U4370 ( .B1(n3417), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3442), 
        .ZN(n6193) );
  INV_X1 U4371 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6057) );
  OAI21_X1 U4372 ( .B1(n6822), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6633), 
        .ZN(n3419) );
  NAND2_X1 U4373 ( .A1(n4278), .A2(EAX_REG_4__SCAN_IN), .ZN(n3418) );
  OAI211_X1 U4374 ( .C1(n3420), .C2(n6057), .A(n3419), .B(n3418), .ZN(n3421)
         );
  OAI21_X1 U4375 ( .B1(n6193), .B2(n4301), .A(n3421), .ZN(n3422) );
  AOI22_X1 U4376 ( .A1(n3877), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4377 ( .A1(n3774), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3426) );
  AOI22_X1 U4378 ( .A1(n3813), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4486), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U4379 ( .A1(n3857), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3424) );
  NAND4_X1 U4380 ( .A1(n3427), .A2(n3426), .A3(n3425), .A4(n3424), .ZN(n3433)
         );
  AOI22_X1 U4381 ( .A1(n3887), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4382 ( .A1(n3818), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4383 ( .A1(n3886), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4384 ( .A1(n3881), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3428) );
  NAND4_X1 U4385 ( .A1(n3431), .A2(n3430), .A3(n3429), .A4(n3428), .ZN(n3432)
         );
  NAND2_X1 U4386 ( .A1(n4022), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3434) );
  INV_X1 U4387 ( .A(n3438), .ZN(n3436) );
  NAND2_X1 U4388 ( .A1(n3437), .A2(n3436), .ZN(n3440) );
  INV_X1 U4389 ( .A(n3437), .ZN(n3439) );
  NAND2_X1 U4390 ( .A1(n3439), .A2(n3438), .ZN(n3461) );
  NAND2_X1 U4391 ( .A1(n3440), .A2(n3461), .ZN(n3950) );
  AOI22_X1 U4392 ( .A1(n4278), .A2(EAX_REG_5__SCAN_IN), .B1(n3903), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3441) );
  OAI21_X1 U4393 ( .B1(n3443), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3464), 
        .ZN(n6306) );
  NAND2_X1 U4394 ( .A1(n4685), .A2(n4713), .ZN(n4714) );
  INV_X1 U4395 ( .A(n4714), .ZN(n3469) );
  INV_X1 U4396 ( .A(n3461), .ZN(n3458) );
  AOI22_X1 U4397 ( .A1(n3818), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4398 ( .A1(n3886), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3448) );
  AOI22_X1 U4399 ( .A1(n3880), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3447) );
  AOI22_X1 U4400 ( .A1(n3879), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3446) );
  NAND4_X1 U4401 ( .A1(n3449), .A2(n3448), .A3(n3447), .A4(n3446), .ZN(n3455)
         );
  AOI22_X1 U4402 ( .A1(n3774), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4403 ( .A1(n4486), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3452) );
  AOI22_X1 U4404 ( .A1(n3813), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4405 ( .A1(n3857), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3450) );
  NAND4_X1 U4406 ( .A1(n3453), .A2(n3452), .A3(n3451), .A4(n3450), .ZN(n3454)
         );
  NAND2_X1 U4407 ( .A1(n4022), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3456) );
  INV_X1 U4408 ( .A(n3459), .ZN(n3460) );
  NAND2_X1 U4409 ( .A1(n3461), .A2(n3460), .ZN(n3462) );
  NAND2_X1 U4410 ( .A1(n3973), .A2(n3462), .ZN(n3957) );
  NAND2_X1 U4411 ( .A1(n3632), .A2(EAX_REG_6__SCAN_IN), .ZN(n3466) );
  AOI21_X1 U4412 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n6164), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3463) );
  INV_X1 U4413 ( .A(n3463), .ZN(n3465) );
  AOI21_X1 U4414 ( .B1(n3464), .B2(n6164), .A(n3473), .ZN(n6165) );
  AOI22_X1 U4415 ( .A1(n3466), .A2(n3465), .B1(n3829), .B2(n6165), .ZN(n3467)
         );
  NAND2_X1 U4416 ( .A1(n4022), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3470) );
  OAI21_X1 U4417 ( .B1(n4057), .B2(n3471), .A(n3470), .ZN(n3472) );
  OAI21_X1 U4418 ( .B1(n3473), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3491), 
        .ZN(n6299) );
  NAND2_X1 U4419 ( .A1(n6299), .A2(n3829), .ZN(n3475) );
  AOI22_X1 U4420 ( .A1(n3632), .A2(EAX_REG_7__SCAN_IN), .B1(n3903), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3474) );
  NAND2_X1 U4421 ( .A1(n3475), .A2(n3474), .ZN(n3476) );
  AOI22_X1 U4422 ( .A1(n3879), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3480) );
  AOI22_X1 U4423 ( .A1(n4486), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4424 ( .A1(n3880), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4425 ( .A1(n3877), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3477) );
  NAND4_X1 U4426 ( .A1(n3480), .A2(n3479), .A3(n3478), .A4(n3477), .ZN(n3486)
         );
  AOI22_X1 U4427 ( .A1(n3818), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3484) );
  AOI22_X1 U4428 ( .A1(n3886), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4429 ( .A1(n3813), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4430 ( .A1(n3857), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3481) );
  NAND4_X1 U4431 ( .A1(n3484), .A2(n3483), .A3(n3482), .A4(n3481), .ZN(n3485)
         );
  NOR2_X1 U4432 ( .A1(n3486), .A2(n3485), .ZN(n3490) );
  INV_X1 U4433 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3487) );
  XNOR2_X1 U4434 ( .A(n3491), .B(n3487), .ZN(n6143) );
  NAND2_X1 U4435 ( .A1(n6143), .A2(n3829), .ZN(n3489) );
  AOI22_X1 U4436 ( .A1(n3632), .A2(EAX_REG_8__SCAN_IN), .B1(n3903), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3488) );
  OAI211_X1 U4437 ( .C1(n3490), .C2(n3552), .A(n3489), .B(n3488), .ZN(n5177)
         );
  XOR2_X1 U4438 ( .A(n6128), .B(n3506), .Z(n6132) );
  AOI22_X1 U4439 ( .A1(n3887), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3496) );
  AOI22_X1 U4440 ( .A1(n3813), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4441 ( .A1(n3881), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3888), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U4442 ( .A1(n3879), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3493) );
  NAND4_X1 U4443 ( .A1(n3496), .A2(n3495), .A3(n3494), .A4(n3493), .ZN(n3502)
         );
  AOI22_X1 U4444 ( .A1(n3818), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U4445 ( .A1(n3886), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3499) );
  AOI22_X1 U4446 ( .A1(n3819), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3498) );
  AOI22_X1 U4447 ( .A1(n4486), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3497) );
  NAND4_X1 U4448 ( .A1(n3500), .A2(n3499), .A3(n3498), .A4(n3497), .ZN(n3501)
         );
  OR2_X1 U4449 ( .A1(n3502), .A2(n3501), .ZN(n3503) );
  AOI22_X1 U4450 ( .A1(n3600), .A2(n3503), .B1(n3903), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3505) );
  NAND2_X1 U4451 ( .A1(n3632), .A2(EAX_REG_9__SCAN_IN), .ZN(n3504) );
  OAI211_X1 U4452 ( .C1(n6132), .C2(n4301), .A(n3505), .B(n3504), .ZN(n5158)
         );
  XNOR2_X1 U4453 ( .A(n3521), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5275)
         );
  AOI22_X1 U4454 ( .A1(n3886), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3510) );
  AOI22_X1 U4455 ( .A1(n4486), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3509) );
  AOI22_X1 U4456 ( .A1(n3774), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3508) );
  AOI22_X1 U4457 ( .A1(n3877), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3507) );
  NAND4_X1 U4458 ( .A1(n3510), .A2(n3509), .A3(n3508), .A4(n3507), .ZN(n3516)
         );
  AOI22_X1 U4459 ( .A1(n3818), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3887), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4460 ( .A1(n3879), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4461 ( .A1(n3813), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4462 ( .A1(n3857), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3511) );
  NAND4_X1 U4463 ( .A1(n3514), .A2(n3513), .A3(n3512), .A4(n3511), .ZN(n3515)
         );
  OAI21_X1 U4464 ( .B1(n3516), .B2(n3515), .A(n3600), .ZN(n3519) );
  NAND2_X1 U4465 ( .A1(n3632), .A2(EAX_REG_10__SCAN_IN), .ZN(n3518) );
  NAND2_X1 U4466 ( .A1(n3903), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3517)
         );
  NAND3_X1 U4467 ( .A1(n3519), .A2(n3518), .A3(n3517), .ZN(n3520) );
  AOI21_X1 U4468 ( .B1(n5275), .B2(n3829), .A(n3520), .ZN(n5242) );
  XOR2_X1 U4469 ( .A(n3548), .B(n3549), .Z(n6293) );
  INV_X1 U4470 ( .A(n6293), .ZN(n3536) );
  AOI22_X1 U4471 ( .A1(n3818), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3525) );
  AOI22_X1 U4472 ( .A1(n3813), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3524) );
  AOI22_X1 U4473 ( .A1(n3886), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3523) );
  AOI22_X1 U4474 ( .A1(n4486), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3522) );
  NAND4_X1 U4475 ( .A1(n3525), .A2(n3524), .A3(n3523), .A4(n3522), .ZN(n3531)
         );
  AOI22_X1 U4476 ( .A1(n3879), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U4477 ( .A1(n3819), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3888), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3528) );
  AOI22_X1 U4478 ( .A1(n3887), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U4479 ( .A1(n3880), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3526) );
  NAND4_X1 U4480 ( .A1(n3529), .A2(n3528), .A3(n3527), .A4(n3526), .ZN(n3530)
         );
  OAI21_X1 U4481 ( .B1(n3531), .B2(n3530), .A(n3600), .ZN(n3534) );
  NAND2_X1 U4482 ( .A1(n3632), .A2(EAX_REG_11__SCAN_IN), .ZN(n3533) );
  NAND2_X1 U4483 ( .A1(n3903), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3532)
         );
  NAND3_X1 U4484 ( .A1(n3534), .A2(n3533), .A3(n3532), .ZN(n3535) );
  AOI22_X1 U4485 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3768), .B1(n3886), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4486 ( .A1(n3813), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4487 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4486), .B1(n3881), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4488 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3877), .B1(n3840), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3538) );
  NAND4_X1 U4489 ( .A1(n3541), .A2(n3540), .A3(n3539), .A4(n3538), .ZN(n3547)
         );
  AOI22_X1 U4490 ( .A1(n3818), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3545) );
  AOI22_X1 U4491 ( .A1(n3774), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4492 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n3819), .B1(n3796), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3543) );
  AOI22_X1 U4493 ( .A1(n3845), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3542) );
  NAND4_X1 U4494 ( .A1(n3545), .A2(n3544), .A3(n3543), .A4(n3542), .ZN(n3546)
         );
  NOR2_X1 U4495 ( .A1(n3547), .A2(n3546), .ZN(n3553) );
  XNOR2_X1 U4496 ( .A(n3554), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5326)
         );
  NAND2_X1 U4497 ( .A1(n5326), .A2(n3829), .ZN(n3551) );
  AOI22_X1 U4498 ( .A1(n3632), .A2(EAX_REG_12__SCAN_IN), .B1(n3903), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3550) );
  NAND2_X1 U4499 ( .A1(n4278), .A2(EAX_REG_13__SCAN_IN), .ZN(n3557) );
  OAI21_X1 U4500 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3555), .A(n3577), 
        .ZN(n6118) );
  AOI22_X1 U4501 ( .A1(n3829), .A2(n6118), .B1(n3903), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3556) );
  OR2_X2 U4502 ( .A1(n3559), .A2(n3558), .ZN(n3576) );
  NAND2_X1 U4503 ( .A1(n3559), .A2(n3558), .ZN(n3560) );
  NAND2_X1 U4504 ( .A1(n3576), .A2(n3560), .ZN(n5357) );
  INV_X1 U4505 ( .A(n5357), .ZN(n3575) );
  AOI22_X1 U4506 ( .A1(n3886), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4507 ( .A1(n3813), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4508 ( .A1(n4486), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3888), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4509 ( .A1(n3818), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3561) );
  NAND4_X1 U4510 ( .A1(n3564), .A2(n3563), .A3(n3562), .A4(n3561), .ZN(n3572)
         );
  AOI22_X1 U4511 ( .A1(n3877), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4512 ( .A1(n3768), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4513 ( .A1(n3774), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4514 ( .A1(n3881), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3567) );
  NAND4_X1 U4515 ( .A1(n3570), .A2(n3569), .A3(n3568), .A4(n3567), .ZN(n3571)
         );
  OR2_X1 U4516 ( .A1(n3572), .A2(n3571), .ZN(n3573) );
  NAND2_X1 U4517 ( .A1(n3600), .A2(n3573), .ZN(n5358) );
  NAND2_X1 U4518 ( .A1(n3575), .A2(n3574), .ZN(n5360) );
  XOR2_X1 U4519 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3591), .Z(n5697) );
  AOI22_X1 U4520 ( .A1(n3877), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4521 ( .A1(n4486), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4522 ( .A1(n3813), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4523 ( .A1(n3857), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3578) );
  NAND4_X1 U4524 ( .A1(n3581), .A2(n3580), .A3(n3579), .A4(n3578), .ZN(n3587)
         );
  AOI22_X1 U4525 ( .A1(n3887), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4526 ( .A1(n3879), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4527 ( .A1(n3886), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4528 ( .A1(n3818), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3582) );
  NAND4_X1 U4529 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(n3586)
         );
  OR2_X1 U4530 ( .A1(n3587), .A2(n3586), .ZN(n3588) );
  AOI22_X1 U4531 ( .A1(n3600), .A2(n3588), .B1(n3903), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3590) );
  NAND2_X1 U4532 ( .A1(n3632), .A2(EAX_REG_14__SCAN_IN), .ZN(n3589) );
  OAI211_X1 U4533 ( .C1(n5697), .C2(n4301), .A(n3590), .B(n3589), .ZN(n5344)
         );
  XNOR2_X1 U4534 ( .A(n3607), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5688)
         );
  INV_X1 U4535 ( .A(n5688), .ZN(n3606) );
  AOI22_X1 U4536 ( .A1(n3818), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4537 ( .A1(n3774), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4538 ( .A1(n3886), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4539 ( .A1(n3857), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3592) );
  NAND4_X1 U4540 ( .A1(n3595), .A2(n3594), .A3(n3593), .A4(n3592), .ZN(n3602)
         );
  AOI22_X1 U4541 ( .A1(n3768), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3599) );
  AOI22_X1 U4542 ( .A1(n3813), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4543 ( .A1(n3877), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4544 ( .A1(n4486), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3596) );
  NAND4_X1 U4545 ( .A1(n3599), .A2(n3598), .A3(n3597), .A4(n3596), .ZN(n3601)
         );
  OAI21_X1 U4546 ( .B1(n3602), .B2(n3601), .A(n3600), .ZN(n3604) );
  NAND2_X1 U4547 ( .A1(n4278), .A2(EAX_REG_15__SCAN_IN), .ZN(n3603) );
  OAI211_X1 U4548 ( .C1(n3762), .C2(n5686), .A(n3604), .B(n3603), .ZN(n3605)
         );
  AOI21_X1 U4549 ( .B1(n3606), .B2(n3829), .A(n3605), .ZN(n5475) );
  XOR2_X1 U4550 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3620), .Z(n6098) );
  AOI22_X1 U4551 ( .A1(n3632), .A2(EAX_REG_16__SCAN_IN), .B1(n3903), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4552 ( .A1(n3877), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4553 ( .A1(n3886), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4554 ( .A1(n3879), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4555 ( .A1(n3813), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3608) );
  NAND4_X1 U4556 ( .A1(n3611), .A2(n3610), .A3(n3609), .A4(n3608), .ZN(n3617)
         );
  AOI22_X1 U4557 ( .A1(n3768), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4558 ( .A1(n3881), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4559 ( .A1(n4486), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3888), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4560 ( .A1(n3818), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3612) );
  NAND4_X1 U4561 ( .A1(n3615), .A2(n3614), .A3(n3613), .A4(n3612), .ZN(n3616)
         );
  OAI21_X1 U4562 ( .B1(n3617), .B2(n3616), .A(n3872), .ZN(n3618) );
  OAI211_X1 U4563 ( .C1(n6098), .C2(n4301), .A(n3619), .B(n3618), .ZN(n5560)
         );
  XNOR2_X1 U4564 ( .A(n3653), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6087)
         );
  NAND2_X1 U4565 ( .A1(n6087), .A2(n3829), .ZN(n3636) );
  AOI22_X1 U4566 ( .A1(n3818), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4567 ( .A1(n3886), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3887), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4568 ( .A1(n3880), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4569 ( .A1(n3879), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3621) );
  NAND4_X1 U4570 ( .A1(n3624), .A2(n3623), .A3(n3622), .A4(n3621), .ZN(n3630)
         );
  AOI22_X1 U4571 ( .A1(n3774), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4572 ( .A1(n4486), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3627) );
  AOI22_X1 U4573 ( .A1(n3813), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4574 ( .A1(n3857), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3625) );
  NAND4_X1 U4575 ( .A1(n3628), .A2(n3627), .A3(n3626), .A4(n3625), .ZN(n3629)
         );
  NOR2_X1 U4576 ( .A1(n3630), .A2(n3629), .ZN(n3634) );
  AOI21_X1 U4577 ( .B1(n6084), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3631) );
  AOI21_X1 U4578 ( .B1(n3632), .B2(EAX_REG_17__SCAN_IN), .A(n3631), .ZN(n3633)
         );
  OAI21_X1 U4579 ( .B1(n3900), .B2(n3634), .A(n3633), .ZN(n3635) );
  NAND2_X1 U4580 ( .A1(n3636), .A2(n3635), .ZN(n5551) );
  NAND2_X1 U4581 ( .A1(n3638), .A2(n3637), .ZN(n5541) );
  INV_X1 U4582 ( .A(n5541), .ZN(n3658) );
  AOI22_X1 U4583 ( .A1(n3818), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4584 ( .A1(n3813), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4486), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4585 ( .A1(n3886), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4586 ( .A1(n3857), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3639) );
  NAND4_X1 U4587 ( .A1(n3642), .A2(n3641), .A3(n3640), .A4(n3639), .ZN(n3648)
         );
  AOI22_X1 U4588 ( .A1(n3879), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4589 ( .A1(n3881), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4590 ( .A1(n3768), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4591 ( .A1(n3877), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3643) );
  NAND4_X1 U4592 ( .A1(n3646), .A2(n3645), .A3(n3644), .A4(n3643), .ZN(n3647)
         );
  NOR2_X1 U4593 ( .A1(n3648), .A2(n3647), .ZN(n3652) );
  OAI21_X1 U4594 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6822), .A(n6633), 
        .ZN(n3649) );
  INV_X1 U4595 ( .A(n3649), .ZN(n3650) );
  AOI21_X1 U4596 ( .B1(n4278), .B2(EAX_REG_18__SCAN_IN), .A(n3650), .ZN(n3651)
         );
  OAI21_X1 U4597 ( .B1(n3900), .B2(n3652), .A(n3651), .ZN(n3656) );
  OAI21_X1 U4598 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n3654), .A(n3673), 
        .ZN(n6077) );
  OR2_X1 U4599 ( .A1(n4301), .A2(n6077), .ZN(n3655) );
  NAND2_X1 U4600 ( .A1(n3656), .A2(n3655), .ZN(n5542) );
  NAND2_X1 U4601 ( .A1(n3658), .A2(n3657), .ZN(n5530) );
  XNOR2_X1 U4602 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n3673), .ZN(n5980)
         );
  AOI22_X1 U4603 ( .A1(n3877), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4604 ( .A1(n3813), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U4605 ( .A1(n3819), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4606 ( .A1(n4486), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3659) );
  NAND4_X1 U4607 ( .A1(n3662), .A2(n3661), .A3(n3660), .A4(n3659), .ZN(n3668)
         );
  AOI22_X1 U4608 ( .A1(n3886), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3887), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3666) );
  AOI22_X1 U4609 ( .A1(n3774), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3857), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4610 ( .A1(n3879), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4611 ( .A1(n3818), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3663) );
  NAND4_X1 U4612 ( .A1(n3666), .A2(n3665), .A3(n3664), .A4(n3663), .ZN(n3667)
         );
  NOR2_X1 U4613 ( .A1(n3668), .A2(n3667), .ZN(n3670) );
  AOI22_X1 U4614 ( .A1(n3632), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6633), .ZN(n3669) );
  OAI21_X1 U4615 ( .B1(n3900), .B2(n3670), .A(n3669), .ZN(n3671) );
  INV_X1 U4616 ( .A(n3671), .ZN(n3672) );
  MUX2_X1 U4617 ( .A(n5980), .B(n3672), .S(n4301), .Z(n5532) );
  OAI21_X1 U4618 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n3674), .A(n3704), 
        .ZN(n5656) );
  AOI22_X1 U4619 ( .A1(n3818), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3678) );
  AOI22_X1 U4620 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n3819), .B1(n3774), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3677) );
  AOI22_X1 U4621 ( .A1(n4486), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4622 ( .A1(n3886), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3675) );
  NAND4_X1 U4623 ( .A1(n3678), .A2(n3677), .A3(n3676), .A4(n3675), .ZN(n3684)
         );
  AOI22_X1 U4624 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3768), .B1(n3879), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4625 ( .A1(n3880), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4626 ( .A1(n3813), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4627 ( .A1(n3857), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3679) );
  NAND4_X1 U4628 ( .A1(n3682), .A2(n3681), .A3(n3680), .A4(n3679), .ZN(n3683)
         );
  NOR2_X1 U4629 ( .A1(n3684), .A2(n3683), .ZN(n3686) );
  AOI22_X1 U4630 ( .A1(n3632), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6633), .ZN(n3685) );
  OAI21_X1 U4631 ( .B1(n3900), .B2(n3686), .A(n3685), .ZN(n3687) );
  MUX2_X1 U4632 ( .A(n5656), .B(n3687), .S(n4301), .Z(n5462) );
  NAND2_X1 U4633 ( .A1(n5460), .A2(n5462), .ZN(n5461) );
  INV_X1 U4634 ( .A(n5461), .ZN(n3703) );
  XNOR2_X1 U4635 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n3704), .ZN(n5970)
         );
  AOI22_X1 U4636 ( .A1(n3768), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4637 ( .A1(n3879), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4638 ( .A1(n3886), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4639 ( .A1(n4486), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3688) );
  NAND4_X1 U4640 ( .A1(n3691), .A2(n3690), .A3(n3689), .A4(n3688), .ZN(n3697)
         );
  AOI22_X1 U4641 ( .A1(n3880), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4642 ( .A1(n3881), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3857), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4643 ( .A1(n3818), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3693) );
  AOI22_X1 U4644 ( .A1(n3813), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3692) );
  NAND4_X1 U4645 ( .A1(n3695), .A2(n3694), .A3(n3693), .A4(n3692), .ZN(n3696)
         );
  NOR2_X1 U4646 ( .A1(n3697), .A2(n3696), .ZN(n3699) );
  AOI22_X1 U4647 ( .A1(n3632), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6633), .ZN(n3698) );
  OAI21_X1 U4648 ( .B1(n3900), .B2(n3699), .A(n3698), .ZN(n3700) );
  INV_X1 U4649 ( .A(n3700), .ZN(n3701) );
  MUX2_X1 U4650 ( .A(n5970), .B(n3701), .S(n4301), .Z(n5523) );
  NAND2_X1 U4651 ( .A1(n3703), .A2(n3702), .ZN(n5512) );
  NOR2_X1 U4652 ( .A1(n3706), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3707)
         );
  NOR2_X1 U4653 ( .A1(n3761), .A2(n3707), .ZN(n5960) );
  AOI22_X1 U4654 ( .A1(n3768), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3711) );
  AOI22_X1 U4655 ( .A1(n3879), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4656 ( .A1(n4486), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3857), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3709) );
  AOI22_X1 U4657 ( .A1(n3877), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3708) );
  NAND4_X1 U4658 ( .A1(n3711), .A2(n3710), .A3(n3709), .A4(n3708), .ZN(n3717)
         );
  AOI22_X1 U4659 ( .A1(n3818), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3886), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4660 ( .A1(n3774), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4661 ( .A1(n3819), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3713) );
  AOI22_X1 U4662 ( .A1(n3813), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3712) );
  NAND4_X1 U4663 ( .A1(n3715), .A2(n3714), .A3(n3713), .A4(n3712), .ZN(n3716)
         );
  NOR2_X1 U4664 ( .A1(n3717), .A2(n3716), .ZN(n3719) );
  AOI22_X1 U4665 ( .A1(n3632), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6633), .ZN(n3718) );
  OAI21_X1 U4666 ( .B1(n3900), .B2(n3719), .A(n3718), .ZN(n3720) );
  INV_X1 U4667 ( .A(n3720), .ZN(n3721) );
  MUX2_X1 U4668 ( .A(n5960), .B(n3721), .S(n4301), .Z(n5514) );
  AOI22_X1 U4669 ( .A1(n3818), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4670 ( .A1(n3880), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4671 ( .A1(n3774), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4672 ( .A1(n3888), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3722) );
  NAND4_X1 U4673 ( .A1(n3725), .A2(n3724), .A3(n3723), .A4(n3722), .ZN(n3731)
         );
  AOI22_X1 U4674 ( .A1(n3886), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3729) );
  AOI22_X1 U4675 ( .A1(n3879), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3728) );
  AOI22_X1 U4676 ( .A1(n3813), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4677 ( .A1(n4486), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3726) );
  NAND4_X1 U4678 ( .A1(n3729), .A2(n3728), .A3(n3727), .A4(n3726), .ZN(n3730)
         );
  NOR2_X1 U4679 ( .A1(n3731), .A2(n3730), .ZN(n3747) );
  AOI22_X1 U4680 ( .A1(n3818), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4681 ( .A1(n3768), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4682 ( .A1(n3862), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4683 ( .A1(n3845), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3732) );
  NAND4_X1 U4684 ( .A1(n3735), .A2(n3734), .A3(n3733), .A4(n3732), .ZN(n3741)
         );
  AOI22_X1 U4685 ( .A1(n3879), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4686 ( .A1(n3880), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4687 ( .A1(n3886), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4688 ( .A1(n4486), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3736) );
  NAND4_X1 U4689 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3740)
         );
  NOR2_X1 U4690 ( .A1(n3741), .A2(n3740), .ZN(n3748) );
  XOR2_X1 U4691 ( .A(n3747), .B(n3748), .Z(n3744) );
  INV_X1 U4692 ( .A(EAX_REG_23__SCAN_IN), .ZN(n3742) );
  INV_X1 U4693 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5632) );
  OAI22_X1 U4694 ( .A1(n3870), .A2(n3742), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5632), .ZN(n3743) );
  AOI21_X1 U4695 ( .B1(n3744), .B2(n3872), .A(n3743), .ZN(n3745) );
  XNOR2_X1 U4696 ( .A(n3761), .B(n5632), .ZN(n5630) );
  MUX2_X1 U4697 ( .A(n3745), .B(n5630), .S(n3829), .Z(n5450) );
  INV_X1 U4698 ( .A(n5450), .ZN(n3746) );
  AND2_X2 U4699 ( .A1(n5447), .A2(n3746), .ZN(n4353) );
  NOR2_X1 U4700 ( .A1(n3748), .A2(n3747), .ZN(n3783) );
  AOI22_X1 U4701 ( .A1(n3818), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4702 ( .A1(n3886), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4703 ( .A1(n3880), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4704 ( .A1(n3879), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3749) );
  NAND4_X1 U4705 ( .A1(n3752), .A2(n3751), .A3(n3750), .A4(n3749), .ZN(n3758)
         );
  AOI22_X1 U4706 ( .A1(n3774), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4707 ( .A1(n4486), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4708 ( .A1(n3862), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3754) );
  AOI22_X1 U4709 ( .A1(n3888), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3753) );
  NAND4_X1 U4710 ( .A1(n3756), .A2(n3755), .A3(n3754), .A4(n3753), .ZN(n3757)
         );
  OR2_X1 U4711 ( .A1(n3758), .A2(n3757), .ZN(n3782) );
  INV_X1 U4712 ( .A(n3782), .ZN(n3759) );
  XNOR2_X1 U4713 ( .A(n3783), .B(n3759), .ZN(n3760) );
  NAND2_X1 U4714 ( .A1(n3760), .A2(n3872), .ZN(n3766) );
  XNOR2_X1 U4715 ( .A(n3767), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5622)
         );
  INV_X1 U4716 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4348) );
  NOR2_X1 U4717 ( .A1(n3762), .A2(n4348), .ZN(n3763) );
  AOI211_X1 U4718 ( .C1(n4278), .C2(EAX_REG_24__SCAN_IN), .A(n3764), .B(n3763), 
        .ZN(n3765) );
  NAND2_X1 U4719 ( .A1(n3766), .A2(n3765), .ZN(n4355) );
  XNOR2_X1 U4720 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .B(n3807), .ZN(n5952)
         );
  AOI22_X1 U4721 ( .A1(n3818), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4722 ( .A1(n3886), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4723 ( .A1(n3880), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4724 ( .A1(n3879), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3770) );
  NAND4_X1 U4725 ( .A1(n3773), .A2(n3772), .A3(n3771), .A4(n3770), .ZN(n3781)
         );
  AOI22_X1 U4726 ( .A1(n3774), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4727 ( .A1(n4486), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4728 ( .A1(n3813), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4729 ( .A1(n3857), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3776) );
  NAND4_X1 U4730 ( .A1(n3779), .A2(n3778), .A3(n3777), .A4(n3776), .ZN(n3780)
         );
  NOR2_X1 U4731 ( .A1(n3781), .A2(n3780), .ZN(n3790) );
  NAND2_X1 U4732 ( .A1(n3783), .A2(n3782), .ZN(n3789) );
  XOR2_X1 U4733 ( .A(n3790), .B(n3789), .Z(n3786) );
  INV_X1 U4734 ( .A(EAX_REG_25__SCAN_IN), .ZN(n3784) );
  INV_X1 U4735 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5606) );
  OAI22_X1 U4736 ( .A1(n3870), .A2(n3784), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5606), .ZN(n3785) );
  AOI21_X1 U4737 ( .B1(n3786), .B2(n3872), .A(n3785), .ZN(n3787) );
  MUX2_X1 U4738 ( .A(n5952), .B(n3787), .S(n4301), .Z(n5498) );
  NOR2_X1 U4739 ( .A1(n3790), .A2(n3789), .ZN(n3812) );
  AOI22_X1 U4740 ( .A1(n3818), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4741 ( .A1(n3886), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4742 ( .A1(n3880), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4743 ( .A1(n3879), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3791) );
  NAND4_X1 U4744 ( .A1(n3794), .A2(n3793), .A3(n3792), .A4(n3791), .ZN(n3802)
         );
  AOI22_X1 U4745 ( .A1(n3774), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4746 ( .A1(n2996), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4747 ( .A1(n3813), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4748 ( .A1(n3888), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3797) );
  NAND4_X1 U4749 ( .A1(n3800), .A2(n3799), .A3(n3798), .A4(n3797), .ZN(n3801)
         );
  OR2_X1 U4750 ( .A1(n3802), .A2(n3801), .ZN(n3811) );
  XNOR2_X1 U4751 ( .A(n3812), .B(n3811), .ZN(n3806) );
  INV_X1 U4752 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3803) );
  AOI21_X1 U4753 ( .B1(n3803), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3804) );
  AOI21_X1 U4754 ( .B1(n4278), .B2(EAX_REG_26__SCAN_IN), .A(n3804), .ZN(n3805)
         );
  OAI21_X1 U4755 ( .B1(n3806), .B2(n3900), .A(n3805), .ZN(n3810) );
  OAI21_X1 U4756 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n3808), .A(n3832), 
        .ZN(n6010) );
  OR2_X1 U4757 ( .A1(n4301), .A2(n6010), .ZN(n3809) );
  NAND2_X1 U4758 ( .A1(n3812), .A2(n3811), .ZN(n3838) );
  AOI22_X1 U4759 ( .A1(n3768), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4760 ( .A1(n3813), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4761 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n3774), .B1(n3565), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4762 ( .A1(n3888), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3814) );
  NAND4_X1 U4763 ( .A1(n3817), .A2(n3816), .A3(n3815), .A4(n3814), .ZN(n3825)
         );
  AOI22_X1 U4764 ( .A1(n3818), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4765 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3881), .B1(n3819), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4766 ( .A1(n3879), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4767 ( .A1(n3886), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3820) );
  NAND4_X1 U4768 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3824)
         );
  NOR2_X1 U4769 ( .A1(n3825), .A2(n3824), .ZN(n3839) );
  XOR2_X1 U4770 ( .A(n3838), .B(n3839), .Z(n3828) );
  INV_X1 U4771 ( .A(EAX_REG_27__SCAN_IN), .ZN(n3826) );
  INV_X1 U4772 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5437) );
  OAI22_X1 U4773 ( .A1(n3870), .A2(n3826), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5437), .ZN(n3827) );
  AOI21_X1 U4774 ( .B1(n3828), .B2(n3872), .A(n3827), .ZN(n3830) );
  XNOR2_X1 U4775 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .B(n3832), .ZN(n5435)
         );
  MUX2_X1 U4776 ( .A(n3830), .B(n5435), .S(n3829), .Z(n3831) );
  AND2_X2 U4777 ( .A1(n4364), .A2(n4365), .ZN(n4363) );
  INV_X1 U4778 ( .A(n3832), .ZN(n3833) );
  INV_X1 U4779 ( .A(n3834), .ZN(n3836) );
  INV_X1 U4780 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3835) );
  NAND2_X1 U4781 ( .A1(n3836), .A2(n3835), .ZN(n3837) );
  NAND2_X1 U4782 ( .A1(n3875), .A2(n3837), .ZN(n5592) );
  NOR2_X1 U4783 ( .A1(n3839), .A2(n3838), .ZN(n3856) );
  AOI22_X1 U4784 ( .A1(n3878), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4785 ( .A1(n3886), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4786 ( .A1(n3880), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4787 ( .A1(n3879), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3841) );
  NAND4_X1 U4788 ( .A1(n3844), .A2(n3843), .A3(n3842), .A4(n3841), .ZN(n3851)
         );
  AOI22_X1 U4789 ( .A1(n3774), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4790 ( .A1(n2996), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4791 ( .A1(n3862), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3565), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4792 ( .A1(n3845), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3846) );
  NAND4_X1 U4793 ( .A1(n3849), .A2(n3848), .A3(n3847), .A4(n3846), .ZN(n3850)
         );
  OR2_X1 U4794 ( .A1(n3851), .A2(n3850), .ZN(n3855) );
  XNOR2_X1 U4795 ( .A(n3856), .B(n3855), .ZN(n3853) );
  AOI22_X1 U4796 ( .A1(n3632), .A2(EAX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6633), .ZN(n3852) );
  OAI21_X1 U4797 ( .B1(n3853), .B2(n3900), .A(n3852), .ZN(n3854) );
  XNOR2_X1 U4798 ( .A(n3875), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5588)
         );
  NAND2_X1 U4799 ( .A1(n3856), .A2(n3855), .ZN(n3895) );
  AOI22_X1 U4800 ( .A1(n3774), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4801 ( .A1(n2996), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3857), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4802 ( .A1(n3877), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4803 ( .A1(n3881), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3565), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3858) );
  NAND4_X1 U4804 ( .A1(n3861), .A2(n3860), .A3(n3859), .A4(n3858), .ZN(n3868)
         );
  AOI22_X1 U4805 ( .A1(n3886), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4806 ( .A1(n3878), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4807 ( .A1(n3879), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4808 ( .A1(n3862), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3863) );
  NAND4_X1 U4809 ( .A1(n3866), .A2(n3865), .A3(n3864), .A4(n3863), .ZN(n3867)
         );
  NOR2_X1 U4810 ( .A1(n3868), .A2(n3867), .ZN(n3896) );
  XOR2_X1 U4811 ( .A(n3895), .B(n3896), .Z(n3873) );
  INV_X1 U4812 ( .A(EAX_REG_29__SCAN_IN), .ZN(n3869) );
  INV_X1 U4813 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5586) );
  OAI22_X1 U4814 ( .A1(n3870), .A2(n3869), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5586), .ZN(n3871) );
  AOI21_X1 U4815 ( .B1(n3873), .B2(n3872), .A(n3871), .ZN(n3874) );
  MUX2_X1 U4816 ( .A(n5588), .B(n3874), .S(n4301), .Z(n5414) );
  INV_X1 U4817 ( .A(n3875), .ZN(n3876) );
  NAND2_X1 U4818 ( .A1(n3876), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4074)
         );
  INV_X1 U4819 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4270) );
  XNOR2_X1 U4820 ( .A(n4074), .B(n4270), .ZN(n5386) );
  AOI22_X1 U4821 ( .A1(n3878), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4822 ( .A1(n3880), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4823 ( .A1(n2996), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4824 ( .A1(n3774), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3565), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3882) );
  NAND4_X1 U4825 ( .A1(n3885), .A2(n3884), .A3(n3883), .A4(n3882), .ZN(n3894)
         );
  AOI22_X1 U4826 ( .A1(n3862), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4827 ( .A1(n3886), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4828 ( .A1(n3887), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4829 ( .A1(n3888), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3889) );
  NAND4_X1 U4830 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(n3893)
         );
  NOR2_X1 U4831 ( .A1(n3894), .A2(n3893), .ZN(n3898) );
  NOR2_X1 U4832 ( .A1(n3896), .A2(n3895), .ZN(n3897) );
  XOR2_X1 U4833 ( .A(n3898), .B(n3897), .Z(n3901) );
  AOI22_X1 U4834 ( .A1(n3632), .A2(EAX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6633), .ZN(n3899) );
  OAI21_X1 U4835 ( .B1(n3901), .B2(n3900), .A(n3899), .ZN(n3902) );
  MUX2_X1 U4836 ( .A(n5386), .B(n3902), .S(n4301), .Z(n4267) );
  AOI22_X1 U4837 ( .A1(n3632), .A2(EAX_REG_31__SCAN_IN), .B1(n3903), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3904) );
  INV_X1 U4838 ( .A(n3904), .ZN(n3905) );
  NAND3_X1 U4839 ( .A1(n6636), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6549) );
  INV_X1 U4840 ( .A(n6549), .ZN(n3906) );
  NOR2_X2 U4841 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6408) );
  NAND2_X1 U4842 ( .A1(n5369), .A2(n6319), .ZN(n4083) );
  NAND2_X1 U4843 ( .A1(n4637), .A2(n4020), .ZN(n3911) );
  NAND2_X1 U4844 ( .A1(n3916), .A2(n3917), .ZN(n3926) );
  INV_X1 U4845 ( .A(n3907), .ZN(n3927) );
  NAND2_X1 U4846 ( .A1(n3926), .A2(n3927), .ZN(n3925) );
  NAND2_X1 U4847 ( .A1(n3925), .A2(n3909), .ZN(n3946) );
  OAI211_X1 U4848 ( .C1(n3909), .C2(n3925), .A(n3946), .B(n6634), .ZN(n3910)
         );
  INV_X1 U4849 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3912) );
  INV_X1 U4850 ( .A(n4020), .ZN(n3975) );
  INV_X1 U4851 ( .A(n6634), .ZN(n4211) );
  AND2_X1 U4852 ( .A1(n4650), .A2(n3222), .ZN(n3928) );
  INV_X1 U4853 ( .A(n3928), .ZN(n3913) );
  OAI21_X1 U4854 ( .B1(n4211), .B2(n3917), .A(n3913), .ZN(n3914) );
  INV_X1 U4855 ( .A(n3914), .ZN(n3915) );
  NAND2_X1 U4856 ( .A1(n6325), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6326)
         );
  XNOR2_X1 U4857 ( .A(n6326), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4549)
         );
  NAND2_X1 U4858 ( .A1(n4639), .A2(n4020), .ZN(n3922) );
  OAI21_X1 U4859 ( .B1(n3917), .B2(n3916), .A(n3926), .ZN(n3918) );
  INV_X1 U4860 ( .A(n3918), .ZN(n3920) );
  NAND3_X1 U4861 ( .A1(n3207), .A2(n3195), .A3(n3222), .ZN(n3919) );
  AOI21_X1 U4862 ( .B1(n6634), .B2(n3920), .A(n3919), .ZN(n3921) );
  NAND2_X1 U4863 ( .A1(n3922), .A2(n3921), .ZN(n4548) );
  NAND2_X1 U4864 ( .A1(n4549), .A2(n4548), .ZN(n4547) );
  INV_X1 U4865 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6378) );
  OR2_X1 U4866 ( .A1(n6326), .A2(n6378), .ZN(n3923) );
  NAND2_X1 U4867 ( .A1(n4547), .A2(n3923), .ZN(n6317) );
  OR2_X1 U4868 ( .A1(n3924), .A2(n3975), .ZN(n3931) );
  OAI21_X1 U4869 ( .B1(n3927), .B2(n3926), .A(n3925), .ZN(n3929) );
  AOI21_X1 U4870 ( .B1(n3929), .B2(n6634), .A(n3928), .ZN(n3930) );
  NAND2_X1 U4871 ( .A1(n3931), .A2(n3930), .ZN(n6316) );
  OAI21_X1 U4872 ( .B1(n6317), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(n6316), 
        .ZN(n3933) );
  NAND2_X1 U4873 ( .A1(n6317), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3932)
         );
  NAND2_X1 U4874 ( .A1(n3933), .A2(n3932), .ZN(n4556) );
  NAND2_X1 U4875 ( .A1(n4555), .A2(n4556), .ZN(n3936) );
  NAND2_X1 U4876 ( .A1(n3934), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3935)
         );
  NAND2_X1 U4877 ( .A1(n3936), .A2(n3935), .ZN(n4619) );
  NAND2_X1 U4878 ( .A1(n3937), .A2(n4020), .ZN(n3941) );
  XNOR2_X1 U4879 ( .A(n3946), .B(n3938), .ZN(n3939) );
  NAND2_X1 U4880 ( .A1(n3939), .A2(n6634), .ZN(n3940) );
  INV_X1 U4881 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4133) );
  NAND2_X1 U4882 ( .A1(n4619), .A2(n4618), .ZN(n3944) );
  NAND2_X1 U4883 ( .A1(n3942), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3943)
         );
  NAND2_X1 U4884 ( .A1(n3944), .A2(n3943), .ZN(n4703) );
  NOR2_X1 U4885 ( .A1(n3946), .A2(n3945), .ZN(n3948) );
  NAND2_X1 U4886 ( .A1(n3948), .A2(n3947), .ZN(n3963) );
  OAI211_X1 U4887 ( .C1(n3948), .C2(n3947), .A(n3963), .B(n6634), .ZN(n3949)
         );
  INV_X1 U4888 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3951) );
  XNOR2_X1 U4889 ( .A(n3952), .B(n3951), .ZN(n4702) );
  NAND2_X1 U4890 ( .A1(n4703), .A2(n4702), .ZN(n3954) );
  NAND2_X1 U4891 ( .A1(n3952), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3953)
         );
  NAND2_X1 U4892 ( .A1(n3954), .A2(n3953), .ZN(n4907) );
  XNOR2_X1 U4893 ( .A(n3963), .B(n3964), .ZN(n3955) );
  NAND2_X1 U4894 ( .A1(n3955), .A2(n6634), .ZN(n3956) );
  INV_X1 U4895 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3958) );
  XNOR2_X1 U4896 ( .A(n3959), .B(n3958), .ZN(n4908) );
  NAND2_X1 U4897 ( .A1(n4907), .A2(n4908), .ZN(n3961) );
  NAND2_X1 U4898 ( .A1(n3959), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3960)
         );
  NAND2_X1 U4899 ( .A1(n3961), .A2(n3960), .ZN(n5171) );
  NAND2_X1 U4900 ( .A1(n3962), .A2(n4020), .ZN(n3968) );
  INV_X1 U4901 ( .A(n3963), .ZN(n3965) );
  NAND2_X1 U4902 ( .A1(n3965), .A2(n3964), .ZN(n3979) );
  XNOR2_X1 U4903 ( .A(n3979), .B(n3977), .ZN(n3966) );
  NAND2_X1 U4904 ( .A1(n3966), .A2(n6634), .ZN(n3967) );
  NAND2_X1 U4905 ( .A1(n3968), .A2(n3967), .ZN(n3970) );
  INV_X1 U4906 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3969) );
  XNOR2_X1 U4907 ( .A(n3970), .B(n3969), .ZN(n5172) );
  NAND2_X1 U4908 ( .A1(n5171), .A2(n5172), .ZN(n3972) );
  NAND2_X1 U4909 ( .A1(n3970), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3971)
         );
  NOR2_X1 U4910 ( .A1(n3319), .A2(n3975), .ZN(n3976) );
  NAND2_X1 U4911 ( .A1(n6634), .A2(n3977), .ZN(n3978) );
  OR2_X1 U4912 ( .A1(n3979), .A2(n3978), .ZN(n3980) );
  INV_X1 U4913 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4147) );
  XNOR2_X1 U4914 ( .A(n3981), .B(n4147), .ZN(n5161) );
  NAND2_X1 U4915 ( .A1(n3981), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3982)
         );
  INV_X1 U4916 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U4917 ( .A1(n2999), .A2(n6355), .ZN(n3983) );
  INV_X1 U4918 ( .A(n5269), .ZN(n3985) );
  INV_X1 U4919 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6348) );
  AND2_X1 U4920 ( .A1(n2999), .A2(n6348), .ZN(n5271) );
  INV_X1 U4921 ( .A(n5271), .ZN(n3984) );
  OR2_X1 U4922 ( .A1(n2999), .A2(n6348), .ZN(n5270) );
  INV_X1 U4923 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5318) );
  NAND2_X1 U4924 ( .A1(n2999), .A2(n5318), .ZN(n5296) );
  OR2_X1 U4925 ( .A1(n2999), .A2(n5318), .ZN(n5297) );
  INV_X1 U4926 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4161) );
  NOR2_X1 U4927 ( .A1(n2999), .A2(n4161), .ZN(n5312) );
  NAND2_X1 U4928 ( .A1(n2999), .A2(n4161), .ZN(n5310) );
  OAI21_X1 U4929 ( .B1(n5309), .B2(n5312), .A(n5310), .ZN(n5812) );
  XNOR2_X1 U4930 ( .A(n2999), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5811)
         );
  INV_X1 U4931 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4214) );
  NAND2_X1 U4932 ( .A1(n2999), .A2(n4214), .ZN(n3986) );
  NAND2_X1 U4933 ( .A1(n5810), .A2(n3986), .ZN(n5694) );
  INV_X1 U4934 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5803) );
  OR2_X1 U4935 ( .A1(n2999), .A2(n5803), .ZN(n3987) );
  NAND2_X1 U4936 ( .A1(n2999), .A2(n5803), .ZN(n3988) );
  XNOR2_X1 U4937 ( .A(n2999), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5689)
         );
  INV_X1 U4938 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3989) );
  NAND2_X1 U4939 ( .A1(n2999), .A2(n3989), .ZN(n3990) );
  NAND2_X1 U4940 ( .A1(n2999), .A2(n6042), .ZN(n5677) );
  AND2_X1 U4941 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5767) );
  INV_X1 U4942 ( .A(n5767), .ZN(n3992) );
  NAND2_X1 U4943 ( .A1(n2999), .A2(n3992), .ZN(n3993) );
  INV_X1 U4944 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5765) );
  INV_X1 U4945 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5792) );
  AND3_X1 U4946 ( .A1(n6042), .A2(n5765), .A3(n5792), .ZN(n3994) );
  NAND2_X1 U4947 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5774) );
  AND2_X1 U4948 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5741) );
  AND2_X1 U4949 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4246) );
  AND2_X1 U4950 ( .A1(n5741), .A2(n4246), .ZN(n4233) );
  INV_X1 U4951 ( .A(n4233), .ZN(n3996) );
  OAI21_X1 U4952 ( .B1(n5774), .B2(n3996), .A(n2999), .ZN(n3997) );
  NAND2_X1 U4953 ( .A1(n5659), .A2(n3997), .ZN(n4001) );
  NOR2_X1 U4954 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3998) );
  NOR2_X1 U4955 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5764) );
  INV_X1 U4956 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5734) );
  INV_X1 U4957 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5759) );
  NAND4_X1 U4958 ( .A1(n3998), .A2(n5764), .A3(n5734), .A4(n5759), .ZN(n3999)
         );
  NAND2_X1 U4959 ( .A1(n5670), .A2(n3999), .ZN(n4000) );
  XNOR2_X1 U4960 ( .A(n2999), .B(n6026), .ZN(n5604) );
  NAND2_X1 U4961 ( .A1(n2999), .A2(n6026), .ZN(n4004) );
  INV_X1 U4962 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U4963 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5717) );
  INV_X1 U4964 ( .A(n5717), .ZN(n4335) );
  NAND2_X1 U4965 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5703) );
  INV_X1 U4966 ( .A(n4005), .ZN(n5603) );
  INV_X1 U4967 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4253) );
  INV_X1 U4968 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5598) );
  NAND3_X1 U4969 ( .A1(n5595), .A2(n4253), .A3(n5598), .ZN(n4006) );
  NOR2_X1 U4970 ( .A1(n2999), .A2(n4006), .ZN(n4261) );
  INV_X1 U4971 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4264) );
  INV_X1 U4972 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4383) );
  NAND4_X1 U4973 ( .A1(n5603), .A2(n4261), .A3(n4264), .A4(n4383), .ZN(n4007)
         );
  OR2_X1 U4974 ( .A1(n3195), .A2(n4650), .ZN(n4008) );
  NAND2_X1 U4975 ( .A1(n4008), .A2(n2986), .ZN(n4028) );
  INV_X1 U4976 ( .A(n4028), .ZN(n4034) );
  AND2_X1 U4977 ( .A1(n6503), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4009)
         );
  NOR2_X1 U4978 ( .A1(n4024), .A2(n4009), .ZN(n4014) );
  AOI21_X1 U4979 ( .B1(n4069), .B2(n4014), .A(n4010), .ZN(n4013) );
  OAI21_X1 U4980 ( .B1(n4057), .B2(n2986), .A(n3195), .ZN(n4015) );
  XNOR2_X1 U4981 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4023) );
  INV_X1 U4982 ( .A(n4023), .ZN(n4011) );
  XNOR2_X1 U4983 ( .A(n4011), .B(n4024), .ZN(n4096) );
  AND2_X1 U4984 ( .A1(n4096), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4016) );
  OR2_X1 U4985 ( .A1(n4015), .A2(n4016), .ZN(n4012) );
  OAI21_X1 U4986 ( .B1(n4034), .B2(n4013), .A(n4012), .ZN(n4021) );
  NAND2_X1 U4987 ( .A1(n4035), .A2(n4014), .ZN(n4019) );
  INV_X1 U4988 ( .A(n4015), .ZN(n4018) );
  INV_X1 U4989 ( .A(n4016), .ZN(n4017) );
  OAI22_X1 U4990 ( .A1(n4021), .A2(n4019), .B1(n4018), .B2(n4017), .ZN(n4033)
         );
  AOI21_X1 U4991 ( .B1(n4021), .B2(n4096), .A(n4052), .ZN(n4032) );
  INV_X1 U4992 ( .A(n4022), .ZN(n4049) );
  NAND2_X1 U4993 ( .A1(n4024), .A2(n4023), .ZN(n4026) );
  NAND2_X1 U4994 ( .A1(n5018), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4025) );
  NAND2_X1 U4995 ( .A1(n4026), .A2(n4025), .ZN(n4039) );
  XNOR2_X1 U4996 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4038) );
  INV_X1 U4997 ( .A(n4038), .ZN(n4027) );
  XNOR2_X1 U4998 ( .A(n4039), .B(n4027), .ZN(n4097) );
  NOR2_X1 U4999 ( .A1(n4049), .A2(n4097), .ZN(n4031) );
  INV_X1 U5000 ( .A(n4097), .ZN(n4029) );
  OAI21_X1 U5001 ( .B1(n4057), .B2(n4029), .A(n4028), .ZN(n4030) );
  OAI22_X1 U5002 ( .A1(n4033), .A2(n4032), .B1(n4031), .B2(n4030), .ZN(n4037)
         );
  NAND3_X1 U5003 ( .A1(n4035), .A2(n4097), .A3(n4034), .ZN(n4036) );
  NAND2_X1 U5004 ( .A1(n4037), .A2(n4036), .ZN(n4051) );
  NAND2_X1 U5005 ( .A1(n4039), .A2(n4038), .ZN(n4041) );
  NAND2_X1 U5006 ( .A1(n6512), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4040) );
  NAND2_X1 U5007 ( .A1(n4041), .A2(n4040), .ZN(n4044) );
  XNOR2_X1 U5008 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4043) );
  INV_X1 U5009 ( .A(n4043), .ZN(n4042) );
  XNOR2_X1 U5010 ( .A(n4044), .B(n4042), .ZN(n4048) );
  NAND2_X1 U5011 ( .A1(n4044), .A2(n4043), .ZN(n4046) );
  NAND2_X1 U5012 ( .A1(n6517), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4045) );
  NAND2_X1 U5013 ( .A1(n4046), .A2(n4045), .ZN(n4053) );
  NAND2_X1 U5014 ( .A1(n4049), .A2(n4060), .ZN(n4050) );
  NAND2_X1 U5015 ( .A1(n4051), .A2(n4050), .ZN(n4062) );
  NAND2_X1 U5016 ( .A1(n4053), .A2(n6394), .ZN(n4054) );
  NAND2_X1 U5017 ( .A1(n4054), .A2(n6057), .ZN(n4056) );
  OAI21_X1 U5018 ( .B1(n6057), .B2(STATE2_REG_0__SCAN_IN), .A(n4058), .ZN(
        n4059) );
  AOI21_X1 U5019 ( .B1(n4064), .B2(n4060), .A(n4059), .ZN(n4061) );
  NAND2_X1 U5020 ( .A1(n4062), .A2(n4061), .ZN(n4066) );
  AOI21_X1 U5021 ( .B1(n4544), .B2(n4650), .A(n4222), .ZN(n4068) );
  INV_X1 U5022 ( .A(n4069), .ZN(n4070) );
  NAND2_X1 U5023 ( .A1(n4113), .A2(n4070), .ZN(n6521) );
  NAND2_X1 U5024 ( .A1(n5896), .A2(n4077), .ZN(n6639) );
  NAND2_X1 U5025 ( .A1(n6639), .A2(n6636), .ZN(n4071) );
  NAND2_X1 U5026 ( .A1(n6636), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4073) );
  NAND2_X1 U5027 ( .A1(n6822), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4072) );
  NAND2_X1 U5028 ( .A1(n4073), .A2(n4072), .ZN(n6329) );
  INV_X1 U5029 ( .A(n4074), .ZN(n4075) );
  NAND2_X1 U5030 ( .A1(n4075), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4076)
         );
  INV_X1 U5031 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4323) );
  OR2_X2 U5032 ( .A1(n4077), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6338) );
  INV_X1 U5033 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6792) );
  NOR2_X1 U5034 ( .A1(n6338), .A2(n6792), .ZN(n5705) );
  AOI21_X1 U5035 ( .B1(n6330), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5705), 
        .ZN(n4078) );
  OAI21_X1 U5036 ( .B1(n6324), .B2(n4350), .A(n4078), .ZN(n4079) );
  INV_X1 U5037 ( .A(n4079), .ZN(n4080) );
  NAND2_X1 U5038 ( .A1(n4083), .A2(n4082), .ZN(U2955) );
  INV_X1 U5039 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U5040 ( .A1(n6026), .A2(n5595), .ZN(n4086) );
  XNOR2_X1 U5041 ( .A(n4090), .B(n4253), .ZN(n4371) );
  INV_X1 U5042 ( .A(n4371), .ZN(n4116) );
  AND2_X1 U5043 ( .A1(n5374), .A2(n4398), .ZN(n4225) );
  NAND2_X1 U5044 ( .A1(n5406), .A2(n4225), .ZN(n4423) );
  OR2_X1 U5045 ( .A1(n4091), .A2(n4650), .ZN(n4092) );
  MUX2_X1 U5046 ( .A(n4092), .B(n4211), .S(n5374), .Z(n4218) );
  NAND2_X1 U5047 ( .A1(n4218), .A2(n4113), .ZN(n4094) );
  NAND2_X1 U5048 ( .A1(n4094), .A2(n5402), .ZN(n4224) );
  OR2_X1 U5049 ( .A1(n4095), .A2(STATE_REG_0__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U5050 ( .A1(n4398), .A2(n6558), .ZN(n4101) );
  NAND3_X1 U5051 ( .A1(n4098), .A2(n4097), .A3(n4096), .ZN(n4099) );
  NAND2_X1 U5052 ( .A1(n4100), .A2(n4099), .ZN(n5400) );
  NOR2_X1 U5053 ( .A1(READY_N), .A2(n5400), .ZN(n4535) );
  NAND3_X1 U5054 ( .A1(n4101), .A2(n4535), .A3(n4222), .ZN(n4102) );
  NAND3_X1 U5055 ( .A1(n4423), .A2(n4224), .A3(n4102), .ZN(n4103) );
  NAND2_X1 U5056 ( .A1(n4103), .A2(n6539), .ZN(n4110) );
  NAND2_X1 U5057 ( .A1(n2986), .A2(n6558), .ZN(n4413) );
  INV_X1 U5058 ( .A(READY_N), .ZN(n6768) );
  NAND2_X1 U5059 ( .A1(n4413), .A2(n6768), .ZN(n4106) );
  OAI211_X1 U5060 ( .C1(n4104), .C2(n4106), .A(n2987), .B(n4105), .ZN(n4107)
         );
  NAND2_X1 U5061 ( .A1(n4107), .A2(n3207), .ZN(n4108) );
  INV_X1 U5062 ( .A(n6521), .ZN(n4114) );
  NOR2_X1 U5063 ( .A1(n4114), .A2(n4540), .ZN(n5399) );
  OAI211_X1 U5064 ( .C1(n3313), .C2(n4212), .A(n4111), .B(n5399), .ZN(n4115)
         );
  NAND2_X1 U5065 ( .A1(n4116), .A2(n6383), .ZN(n4258) );
  NAND2_X1 U5066 ( .A1(n2987), .A2(n4398), .ZN(n4117) );
  NAND2_X1 U5067 ( .A1(n4118), .A2(n6378), .ZN(n4119) );
  OAI211_X1 U5068 ( .C1(n4285), .C2(EBX_REG_1__SCAN_IN), .A(n5467), .B(n4119), 
        .ZN(n4120) );
  NAND2_X1 U5069 ( .A1(n4118), .A2(EBX_REG_0__SCAN_IN), .ZN(n4122) );
  INV_X1 U5070 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4412) );
  NAND2_X1 U5071 ( .A1(n5467), .A2(n4412), .ZN(n4121) );
  NAND2_X1 U5072 ( .A1(n4122), .A2(n4121), .ZN(n4408) );
  XNOR2_X1 U5073 ( .A(n4123), .B(n4408), .ZN(n4443) );
  NAND2_X1 U5074 ( .A1(n4443), .A2(n4442), .ZN(n6233) );
  NAND2_X1 U5075 ( .A1(n6233), .A2(n4123), .ZN(n4631) );
  INV_X1 U5076 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U5077 ( .A1(n4200), .A2(n6215), .ZN(n4128) );
  INV_X1 U5078 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4125) );
  NAND2_X1 U5079 ( .A1(n4118), .A2(n4125), .ZN(n4126) );
  OAI211_X1 U5080 ( .C1(n4285), .C2(EBX_REG_2__SCAN_IN), .A(n5467), .B(n4126), 
        .ZN(n4127) );
  AND2_X1 U5081 ( .A1(n4128), .A2(n4127), .ZN(n4630) );
  NAND2_X1 U5082 ( .A1(n5467), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4131)
         );
  OAI211_X1 U5083 ( .C1(n4285), .C2(EBX_REG_3__SCAN_IN), .A(n4118), .B(n4131), 
        .ZN(n4132) );
  OAI21_X1 U5084 ( .B1(n4199), .B2(EBX_REG_3__SCAN_IN), .A(n4132), .ZN(n4558)
         );
  INV_X1 U5085 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U5086 ( .A1(n4200), .A2(n6191), .ZN(n4136) );
  NAND2_X1 U5087 ( .A1(n4118), .A2(n4133), .ZN(n4134) );
  OAI211_X1 U5088 ( .C1(n4117), .C2(EBX_REG_4__SCAN_IN), .A(n5467), .B(n4134), 
        .ZN(n4135) );
  AND2_X1 U5089 ( .A1(n4136), .A2(n4135), .ZN(n4621) );
  INV_X1 U5090 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4717) );
  MUX2_X1 U5091 ( .A(n5535), .B(n4205), .S(n4717), .Z(n4138) );
  NOR2_X1 U5092 ( .A1(n4409), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4137)
         );
  NOR2_X1 U5093 ( .A1(n4138), .A2(n4137), .ZN(n4704) );
  NAND2_X1 U5094 ( .A1(n4705), .A2(n4704), .ZN(n4741) );
  INV_X1 U5095 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4742) );
  NAND2_X1 U5096 ( .A1(n4200), .A2(n4742), .ZN(n4142) );
  NAND2_X1 U5097 ( .A1(n5467), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4139)
         );
  NAND2_X1 U5098 ( .A1(n4118), .A2(n4139), .ZN(n4140) );
  OAI21_X1 U5099 ( .B1(n4285), .B2(EBX_REG_6__SCAN_IN), .A(n4140), .ZN(n4141)
         );
  OR2_X1 U5100 ( .A1(n4285), .A2(EBX_REG_7__SCAN_IN), .ZN(n4145) );
  OAI211_X1 U5101 ( .C1(n5535), .C2(n3969), .A(n4145), .B(n4118), .ZN(n4146)
         );
  OAI21_X1 U5102 ( .B1(n4199), .B2(EBX_REG_7__SCAN_IN), .A(n4146), .ZN(n5008)
         );
  NAND2_X1 U5103 ( .A1(n4118), .A2(n4147), .ZN(n4148) );
  OAI211_X1 U5104 ( .C1(n4117), .C2(EBX_REG_8__SCAN_IN), .A(n5467), .B(n4148), 
        .ZN(n4149) );
  OAI21_X1 U5105 ( .B1(n4305), .B2(EBX_REG_8__SCAN_IN), .A(n4149), .ZN(n5163)
         );
  INV_X1 U5106 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5184) );
  MUX2_X1 U5107 ( .A(n5535), .B(n4205), .S(n5184), .Z(n4151) );
  NOR2_X1 U5108 ( .A1(n4409), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4150)
         );
  NOR2_X1 U5109 ( .A1(n4151), .A2(n4150), .ZN(n5182) );
  INV_X1 U5110 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4152) );
  NAND2_X1 U5111 ( .A1(n4200), .A2(n4152), .ZN(n4156) );
  NAND2_X1 U5112 ( .A1(n5467), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4153) );
  NAND2_X1 U5113 ( .A1(n4118), .A2(n4153), .ZN(n4154) );
  OAI21_X1 U5114 ( .B1(n4117), .B2(EBX_REG_10__SCAN_IN), .A(n4154), .ZN(n4155)
         );
  NAND2_X1 U5115 ( .A1(n5467), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4159) );
  OAI211_X1 U5116 ( .C1(n4285), .C2(EBX_REG_11__SCAN_IN), .A(n4118), .B(n4159), 
        .ZN(n4160) );
  OAI21_X1 U5117 ( .B1(n4199), .B2(EBX_REG_11__SCAN_IN), .A(n4160), .ZN(n5300)
         );
  NAND2_X1 U5118 ( .A1(n4118), .A2(n4161), .ZN(n4162) );
  OAI211_X1 U5119 ( .C1(n4117), .C2(EBX_REG_12__SCAN_IN), .A(n5467), .B(n4162), 
        .ZN(n4163) );
  OAI21_X1 U5120 ( .B1(n4305), .B2(EBX_REG_12__SCAN_IN), .A(n4163), .ZN(n5281)
         );
  MUX2_X1 U5121 ( .A(n4205), .B(n5535), .S(EBX_REG_13__SCAN_IN), .Z(n4164) );
  INV_X1 U5122 ( .A(n4164), .ZN(n4165) );
  NAND2_X1 U5123 ( .A1(n4165), .A2(n3067), .ZN(n5365) );
  INV_X1 U5124 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U5125 ( .A1(n4200), .A2(n5348), .ZN(n4168) );
  NAND2_X1 U5126 ( .A1(n4118), .A2(n5803), .ZN(n4166) );
  OAI211_X1 U5127 ( .C1(n4285), .C2(EBX_REG_14__SCAN_IN), .A(n5467), .B(n4166), 
        .ZN(n4167) );
  NAND2_X1 U5128 ( .A1(n5467), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4169) );
  OAI211_X1 U5129 ( .C1(n4285), .C2(EBX_REG_15__SCAN_IN), .A(n4118), .B(n4169), 
        .ZN(n4170) );
  OAI21_X1 U5130 ( .B1(n4199), .B2(EBX_REG_15__SCAN_IN), .A(n4170), .ZN(n5477)
         );
  INV_X1 U5131 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U5132 ( .A1(n4205), .A2(n6085), .ZN(n4173) );
  NAND2_X1 U5133 ( .A1(n5467), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4171) );
  OAI211_X1 U5134 ( .C1(n4285), .C2(EBX_REG_17__SCAN_IN), .A(n4118), .B(n4171), 
        .ZN(n4172) );
  NAND2_X1 U5135 ( .A1(n5467), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4174) );
  NAND2_X1 U5136 ( .A1(n4118), .A2(n4174), .ZN(n4175) );
  OAI21_X1 U5137 ( .B1(n4117), .B2(EBX_REG_16__SCAN_IN), .A(n4175), .ZN(n4176)
         );
  OAI21_X1 U5138 ( .B1(n4305), .B2(EBX_REG_16__SCAN_IN), .A(n4176), .ZN(n5562)
         );
  INV_X1 U5139 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U5140 ( .A1(n4200), .A2(n5539), .ZN(n4180) );
  INV_X1 U5141 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U5142 ( .A1(n4118), .A2(n5661), .ZN(n4178) );
  OAI211_X1 U5143 ( .C1(n4285), .C2(EBX_REG_19__SCAN_IN), .A(n5467), .B(n4178), 
        .ZN(n4179) );
  INV_X1 U5144 ( .A(n4409), .ZN(n4288) );
  NAND2_X1 U5145 ( .A1(n4288), .A2(n5765), .ZN(n4181) );
  OR2_X1 U5146 ( .A1(n4117), .A2(EBX_REG_18__SCAN_IN), .ZN(n5536) );
  OR2_X1 U5147 ( .A1(n4117), .A2(EBX_REG_20__SCAN_IN), .ZN(n4182) );
  OAI21_X1 U5148 ( .B1(n4409), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n4182), 
        .ZN(n5468) );
  NAND2_X1 U5149 ( .A1(n5465), .A2(n5468), .ZN(n4184) );
  NAND2_X1 U5150 ( .A1(n5535), .A2(EBX_REG_20__SCAN_IN), .ZN(n4183) );
  OAI211_X1 U5151 ( .C1(n5465), .C2(n5535), .A(n4184), .B(n4183), .ZN(n4185)
         );
  INV_X1 U5152 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5527) );
  MUX2_X1 U5153 ( .A(n5535), .B(n4205), .S(n5527), .Z(n4187) );
  NOR2_X1 U5154 ( .A1(n4409), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4186)
         );
  NOR2_X1 U5155 ( .A1(n4187), .A2(n4186), .ZN(n5525) );
  INV_X1 U5156 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U5157 ( .A1(n4200), .A2(n5520), .ZN(n4191) );
  INV_X1 U5158 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4188) );
  NAND2_X1 U5159 ( .A1(n4118), .A2(n4188), .ZN(n4189) );
  OAI211_X1 U5160 ( .C1(n4285), .C2(EBX_REG_22__SCAN_IN), .A(n5467), .B(n4189), 
        .ZN(n4190) );
  NAND2_X1 U5161 ( .A1(n5467), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4192) );
  OAI211_X1 U5162 ( .C1(n4285), .C2(EBX_REG_23__SCAN_IN), .A(n4118), .B(n4192), 
        .ZN(n4193) );
  OAI21_X1 U5163 ( .B1(n4199), .B2(EBX_REG_23__SCAN_IN), .A(n4193), .ZN(n5452)
         );
  NAND2_X1 U5164 ( .A1(n5467), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4194) );
  NAND2_X1 U5165 ( .A1(n4118), .A2(n4194), .ZN(n4195) );
  OAI21_X1 U5166 ( .B1(n4117), .B2(EBX_REG_24__SCAN_IN), .A(n4195), .ZN(n4196)
         );
  OAI21_X1 U5167 ( .B1(n4305), .B2(EBX_REG_24__SCAN_IN), .A(n4196), .ZN(n4356)
         );
  NAND2_X1 U5168 ( .A1(n5453), .A2(n4356), .ZN(n5503) );
  NAND2_X1 U5169 ( .A1(n5467), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4197) );
  OAI211_X1 U5170 ( .C1(n4285), .C2(EBX_REG_25__SCAN_IN), .A(n4118), .B(n4197), 
        .ZN(n4198) );
  OAI21_X1 U5171 ( .B1(n4199), .B2(EBX_REG_25__SCAN_IN), .A(n4198), .ZN(n5502)
         );
  INV_X1 U5172 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U5173 ( .A1(n4200), .A2(n5497), .ZN(n4204) );
  NAND2_X1 U5174 ( .A1(n5467), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4201) );
  NAND2_X1 U5175 ( .A1(n4118), .A2(n4201), .ZN(n4202) );
  OAI21_X1 U5176 ( .B1(n4117), .B2(EBX_REG_26__SCAN_IN), .A(n4202), .ZN(n4203)
         );
  MUX2_X1 U5177 ( .A(n4205), .B(n5535), .S(EBX_REG_27__SCAN_IN), .Z(n4206) );
  INV_X1 U5178 ( .A(n4206), .ZN(n4208) );
  NAND2_X1 U5179 ( .A1(n4288), .A2(n4253), .ZN(n4207) );
  NAND2_X1 U5180 ( .A1(n4208), .A2(n4207), .ZN(n4209) );
  AND2_X1 U5181 ( .A1(n5493), .A2(n4209), .ZN(n4210) );
  OR2_X1 U5182 ( .A1(n4210), .A2(n5424), .ZN(n5489) );
  INV_X1 U5183 ( .A(n5489), .ZN(n4256) );
  OAI21_X1 U5184 ( .B1(n4212), .B2(n3212), .A(n6531), .ZN(n4213) );
  NOR2_X1 U5185 ( .A1(n5595), .A2(n6026), .ZN(n5726) );
  INV_X1 U5186 ( .A(n5726), .ZN(n4250) );
  NAND2_X1 U5187 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5815) );
  NOR2_X1 U5188 ( .A1(n4214), .A2(n5815), .ZN(n5804) );
  NAND2_X1 U5189 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5804), .ZN(n6045) );
  NAND2_X1 U5190 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6038) );
  NOR2_X1 U5191 ( .A1(n6045), .A2(n6038), .ZN(n4236) );
  NOR2_X1 U5192 ( .A1(n4125), .A2(n6378), .ZN(n6359) );
  NAND3_X1 U5193 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n4910) );
  NOR2_X1 U5194 ( .A1(n3958), .A2(n4910), .ZN(n5162) );
  NAND2_X1 U5195 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6344) );
  NAND2_X1 U5196 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6345) );
  NOR2_X1 U5197 ( .A1(n6344), .A2(n6345), .ZN(n4227) );
  NAND3_X1 U5198 ( .A1(n6359), .A2(n5162), .A3(n4227), .ZN(n5816) );
  OR2_X1 U5199 ( .A1(n5402), .A2(n2986), .ZN(n6504) );
  INV_X1 U5200 ( .A(n6504), .ZN(n5372) );
  NAND2_X1 U5201 ( .A1(n4235), .A2(n5372), .ZN(n6385) );
  OAI21_X1 U5202 ( .B1(n4216), .B2(n4288), .A(n4215), .ZN(n4217) );
  INV_X1 U5203 ( .A(n4217), .ZN(n4219) );
  AND3_X1 U5204 ( .A1(n4220), .A2(n4219), .A3(n4218), .ZN(n4430) );
  NAND2_X1 U5205 ( .A1(n4430), .A2(n4512), .ZN(n4221) );
  NAND2_X1 U5206 ( .A1(n4235), .A2(n4221), .ZN(n5798) );
  NAND2_X1 U5207 ( .A1(n6385), .A2(n5798), .ZN(n4242) );
  INV_X1 U5208 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6371) );
  NAND2_X1 U5209 ( .A1(n6385), .A2(n6371), .ZN(n6368) );
  NAND2_X1 U5210 ( .A1(n4242), .A2(n6368), .ZN(n4557) );
  NOR2_X1 U5211 ( .A1(n5816), .A2(n4557), .ZN(n5304) );
  NAND2_X1 U5212 ( .A1(n4236), .A2(n5304), .ZN(n5780) );
  OR2_X1 U5213 ( .A1(n5100), .A2(n4222), .ZN(n4223) );
  NAND2_X1 U5214 ( .A1(n4420), .A2(n4225), .ZN(n5405) );
  INV_X1 U5215 ( .A(n5405), .ZN(n4226) );
  INV_X1 U5216 ( .A(n4227), .ZN(n4229) );
  AOI21_X1 U5217 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n4708) );
  INV_X1 U5218 ( .A(n4708), .ZN(n4228) );
  NAND2_X1 U5219 ( .A1(n5162), .A2(n4228), .ZN(n5165) );
  NOR2_X1 U5220 ( .A1(n4229), .A2(n5165), .ZN(n5797) );
  INV_X1 U5221 ( .A(n4236), .ZN(n5763) );
  NOR2_X1 U5222 ( .A1(n5792), .A2(n5763), .ZN(n5783) );
  NAND2_X1 U5223 ( .A1(n5797), .A2(n5783), .ZN(n4238) );
  OR2_X1 U5224 ( .A1(n5796), .A2(n4238), .ZN(n4230) );
  NAND2_X1 U5225 ( .A1(n5780), .A2(n4230), .ZN(n4232) );
  AND2_X1 U5226 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4231) );
  AND2_X1 U5227 ( .A1(n5767), .A2(n4231), .ZN(n4243) );
  NAND2_X1 U5228 ( .A1(n5760), .A2(n4233), .ZN(n6019) );
  NOR2_X1 U5229 ( .A1(n4250), .A2(n6019), .ZN(n5719) );
  INV_X1 U5230 ( .A(n5741), .ZN(n4234) );
  NAND2_X1 U5231 ( .A1(n5760), .A2(n4234), .ZN(n5748) );
  INV_X1 U5232 ( .A(n4242), .ZN(n5768) );
  OAI22_X1 U5233 ( .A1(n4235), .A2(n6376), .B1(n5798), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6370) );
  AOI21_X1 U5234 ( .B1(n4242), .B2(n5816), .A(n6370), .ZN(n5305) );
  OAI21_X1 U5235 ( .B1(n5768), .B2(n4236), .A(n5305), .ZN(n4237) );
  INV_X1 U5236 ( .A(n4237), .ZN(n4241) );
  INV_X1 U5237 ( .A(n4238), .ZN(n4239) );
  OR2_X1 U5238 ( .A1(n5796), .A2(n4239), .ZN(n4240) );
  NAND2_X1 U5239 ( .A1(n4241), .A2(n4240), .ZN(n5788) );
  INV_X1 U5240 ( .A(n4243), .ZN(n4244) );
  AND2_X1 U5241 ( .A1(n6369), .A2(n4244), .ZN(n4245) );
  NOR2_X1 U5242 ( .A1(n5788), .A2(n4245), .ZN(n5756) );
  AND2_X1 U5243 ( .A1(n5748), .A2(n5756), .ZN(n5740) );
  NAND2_X1 U5244 ( .A1(n4557), .A2(n5796), .ZN(n4248) );
  INV_X1 U5245 ( .A(n4246), .ZN(n4247) );
  NAND2_X1 U5246 ( .A1(n4248), .A2(n4247), .ZN(n4249) );
  NAND2_X1 U5247 ( .A1(n6369), .A2(n4250), .ZN(n4251) );
  NAND2_X1 U5248 ( .A1(n6027), .A2(n4251), .ZN(n5721) );
  INV_X1 U5249 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6748) );
  NOR2_X1 U5250 ( .A1(n6338), .A2(n6748), .ZN(n4252) );
  AOI221_X1 U5251 ( .B1(n5719), .B2(n4253), .C1(n5721), .C2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .A(n4252), .ZN(n4254) );
  INV_X1 U5252 ( .A(n4254), .ZN(n4255) );
  NAND2_X1 U5253 ( .A1(n4259), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4263) );
  NAND2_X1 U5254 ( .A1(n4260), .A2(n4261), .ZN(n4374) );
  NAND2_X1 U5255 ( .A1(n4263), .A2(n4262), .ZN(n4265) );
  XNOR2_X1 U5256 ( .A(n4265), .B(n4264), .ZN(n4342) );
  INV_X1 U5257 ( .A(n4342), .ZN(n4266) );
  NAND2_X1 U5258 ( .A1(n4266), .A2(n6332), .ZN(n4275) );
  AND2_X2 U5259 ( .A1(n4269), .A2(n4268), .ZN(n5380) );
  NOR2_X1 U5260 ( .A1(n6324), .A2(n5386), .ZN(n4272) );
  INV_X1 U5261 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6787) );
  OR2_X1 U5262 ( .A1(n6338), .A2(n6787), .ZN(n4336) );
  OAI21_X1 U5263 ( .B1(n6314), .B2(n4270), .A(n4336), .ZN(n4271) );
  NOR2_X1 U5264 ( .A1(n4272), .A2(n4271), .ZN(n4273) );
  NAND3_X1 U5265 ( .A1(n4275), .A2(n4274), .A3(n4273), .ZN(U2956) );
  NOR2_X1 U5266 ( .A1(n5405), .A2(n6545), .ZN(n4276) );
  NAND2_X1 U5267 ( .A1(n5406), .A2(n4276), .ZN(n4282) );
  NOR2_X1 U5268 ( .A1(n2997), .A2(n4277), .ZN(n4280) );
  NAND4_X1 U5269 ( .A1(n4280), .A2(n4279), .A3(n4278), .A4(n6542), .ZN(n4536)
         );
  OR2_X1 U5270 ( .A1(n4536), .A2(n4285), .ZN(n4281) );
  NAND2_X2 U5271 ( .A1(n5391), .A2(n5567), .ZN(n6236) );
  NAND2_X1 U5272 ( .A1(n5380), .A2(n4283), .ZN(n4299) );
  NAND2_X1 U5273 ( .A1(n4118), .A2(n5598), .ZN(n4284) );
  OAI211_X1 U5274 ( .C1(n4285), .C2(EBX_REG_28__SCAN_IN), .A(n5467), .B(n4284), 
        .ZN(n4286) );
  OAI21_X1 U5275 ( .B1(n4305), .B2(EBX_REG_28__SCAN_IN), .A(n4286), .ZN(n5423)
         );
  INV_X1 U5276 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4287) );
  AOI22_X1 U5277 ( .A1(n4288), .A2(n4383), .B1(n4442), .B2(n4287), .ZN(n4378)
         );
  INV_X1 U5278 ( .A(n5426), .ZN(n4381) );
  NAND2_X1 U5279 ( .A1(n4409), .A2(EBX_REG_30__SCAN_IN), .ZN(n4290) );
  NAND2_X1 U5280 ( .A1(n4117), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4289) );
  NAND2_X1 U5281 ( .A1(n4290), .A2(n4289), .ZN(n4308) );
  OAI211_X1 U5282 ( .C1(n4306), .C2(n4381), .A(n4307), .B(n4308), .ZN(n4294)
         );
  INV_X1 U5283 ( .A(n4308), .ZN(n4291) );
  OAI21_X1 U5284 ( .B1(n5426), .B2(n5467), .A(n4291), .ZN(n4292) );
  OR2_X1 U5285 ( .A1(n4306), .A2(n4292), .ZN(n4293) );
  INV_X2 U5286 ( .A(n5504), .ZN(n5567) );
  INV_X1 U5287 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4296) );
  NAND2_X1 U5288 ( .A1(n4299), .A2(n4298), .ZN(U2829) );
  NOR2_X1 U5289 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6535) );
  INV_X1 U5290 ( .A(n6535), .ZN(n6635) );
  NOR3_X1 U5291 ( .A1(n6636), .A2(n6623), .A3(n6635), .ZN(n6537) );
  NOR3_X1 U5292 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6542), .A3(n4301), .ZN(
        n6548) );
  NOR2_X1 U5293 ( .A1(n6537), .A2(n6548), .ZN(n4302) );
  NAND2_X1 U5294 ( .A1(n6338), .A2(n4302), .ZN(n4303) );
  NOR2_X1 U5295 ( .A1(n4350), .A2(n6542), .ZN(n4304) );
  NAND2_X1 U5296 ( .A1(n5369), .A2(n6145), .ZN(n4333) );
  NOR2_X1 U5297 ( .A1(n4305), .A2(EBX_REG_29__SCAN_IN), .ZN(n4377) );
  AOI22_X1 U5298 ( .A1(n4306), .A2(n5467), .B1(n4377), .B2(n5426), .ZN(n4379)
         );
  OAI22_X1 U5299 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n4409), .B1(n4117), .B2(EBX_REG_31__SCAN_IN), .ZN(n4309) );
  XNOR2_X1 U5300 ( .A(n4310), .B(n4309), .ZN(n5708) );
  NAND2_X1 U5301 ( .A1(n6768), .A2(n6822), .ZN(n4312) );
  NOR2_X2 U5302 ( .A1(n6633), .A2(n6217), .ZN(n5097) );
  AND2_X1 U5303 ( .A1(n4312), .A2(n5097), .ZN(n4344) );
  NAND2_X1 U5304 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4344), .ZN(n6232) );
  OR2_X1 U5305 ( .A1(n4650), .A2(n6558), .ZN(n4311) );
  NAND2_X1 U5306 ( .A1(n4117), .A2(n4311), .ZN(n4314) );
  INV_X1 U5307 ( .A(n5097), .ZN(n5099) );
  INV_X1 U5308 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6793) );
  NAND2_X1 U5309 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4321) );
  NAND3_X1 U5310 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n4315) );
  INV_X1 U5311 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6590) );
  INV_X1 U5312 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6587) );
  NAND2_X1 U5313 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n6119) );
  NOR2_X1 U5314 ( .A1(n6587), .A2(n6119), .ZN(n5290) );
  NAND2_X1 U5315 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5290), .ZN(n6108) );
  NOR2_X1 U5316 ( .A1(n6590), .A2(n6108), .ZN(n4325) );
  INV_X1 U5317 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6580) );
  NAND3_X1 U5318 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U5319 ( .A1(REIP_REG_5__SCAN_IN), .A2(REIP_REG_4__SCAN_IN), .ZN(
        n6153) );
  NOR2_X1 U5320 ( .A1(n6174), .A2(n6153), .ZN(n6155) );
  NAND2_X1 U5321 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6155), .ZN(n6150) );
  NOR2_X1 U5322 ( .A1(n6580), .A2(n6150), .ZN(n4324) );
  AND3_X1 U5323 ( .A1(n5247), .A2(REIP_REG_8__SCAN_IN), .A3(n4324), .ZN(n5289)
         );
  NAND3_X1 U5324 ( .A1(REIP_REG_14__SCAN_IN), .A2(n4325), .A3(n5289), .ZN(
        n5351) );
  NOR2_X1 U5325 ( .A1(n4315), .A2(n5351), .ZN(n4316) );
  NAND2_X1 U5326 ( .A1(n5247), .A2(n6210), .ZN(n6152) );
  INV_X1 U5327 ( .A(n6152), .ZN(n5288) );
  OR2_X1 U5328 ( .A1(n4316), .A2(n5288), .ZN(n5979) );
  NAND3_X1 U5329 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n4326) );
  NAND2_X1 U5330 ( .A1(n6152), .A2(n4326), .ZN(n4317) );
  NAND2_X1 U5331 ( .A1(n5979), .A2(n4317), .ZN(n5971) );
  AND3_X1 U5332 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4318) );
  NOR2_X1 U5333 ( .A1(n6210), .A2(n4318), .ZN(n4319) );
  NOR2_X1 U5334 ( .A1(n5971), .A2(n4319), .ZN(n5451) );
  NAND3_X1 U5335 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U5336 ( .A1(n6152), .A2(n5440), .ZN(n4320) );
  NAND2_X1 U5337 ( .A1(n5451), .A2(n4320), .ZN(n5944) );
  AOI21_X1 U5338 ( .B1(n6156), .B2(n4321), .A(n5944), .ZN(n5418) );
  INV_X1 U5339 ( .A(n5418), .ZN(n5429) );
  AOI21_X1 U5340 ( .B1(n6156), .B2(n6793), .A(n5429), .ZN(n5382) );
  OAI21_X1 U5341 ( .B1(REIP_REG_30__SCAN_IN), .B2(n6210), .A(n5382), .ZN(n4329) );
  OR3_X1 U5342 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .A3(n6558), .ZN(
        n6530) );
  AND2_X1 U5343 ( .A1(n6530), .A2(n5097), .ZN(n4343) );
  NAND3_X1 U5344 ( .A1(n6634), .A2(EBX_REG_31__SCAN_IN), .A3(n4343), .ZN(n4322) );
  OAI21_X1 U5345 ( .B1(n6205), .B2(n4323), .A(n4322), .ZN(n4328) );
  INV_X1 U5346 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6592) );
  INV_X1 U5347 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6582) );
  NAND2_X1 U5348 ( .A1(n5249), .A2(n4325), .ZN(n5352) );
  NAND4_X1 U5349 ( .A1(n6104), .A2(REIP_REG_17__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .A4(REIP_REG_15__SCAN_IN), .ZN(n6083) );
  NAND4_X1 U5350 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5965), .ZN(n5943) );
  NOR3_X1 U5351 ( .A1(n5943), .A2(n5440), .A3(n6748), .ZN(n5432) );
  NAND2_X1 U5352 ( .A1(n5432), .A2(REIP_REG_28__SCAN_IN), .ZN(n5415) );
  NOR4_X1 U5353 ( .A1(n5415), .A2(REIP_REG_31__SCAN_IN), .A3(n6787), .A4(n6793), .ZN(n4327) );
  AOI211_X1 U5354 ( .C1(REIP_REG_31__SCAN_IN), .C2(n4329), .A(n4328), .B(n4327), .ZN(n4330) );
  OAI21_X1 U5355 ( .B1(n5708), .B2(n6200), .A(n4330), .ZN(n4331) );
  INV_X1 U5356 ( .A(n4331), .ZN(n4332) );
  NAND2_X1 U5357 ( .A1(n4333), .A2(n4332), .ZN(U2796) );
  AOI21_X1 U5358 ( .B1(n6369), .B2(n5717), .A(n5721), .ZN(n4384) );
  NAND2_X1 U5359 ( .A1(n6369), .A2(n5703), .ZN(n4334) );
  NAND2_X1 U5360 ( .A1(n4384), .A2(n4334), .ZN(n5707) );
  NAND2_X1 U5361 ( .A1(n4335), .A2(n5719), .ZN(n5704) );
  NOR2_X1 U5362 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n5704), .ZN(n4338)
         );
  INV_X1 U5363 ( .A(n4336), .ZN(n4337) );
  AOI21_X1 U5364 ( .B1(n4338), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n4337), 
        .ZN(n4339) );
  OAI21_X1 U5365 ( .B1(n5381), .B2(n6339), .A(n4339), .ZN(n4340) );
  OAI21_X1 U5366 ( .B1(n4342), .B2(n6035), .A(n4341), .ZN(U2988) );
  NOR2_X1 U5367 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5943), .ZN(n5954) );
  INV_X1 U5368 ( .A(n5954), .ZN(n4362) );
  NAND2_X1 U5369 ( .A1(n6634), .A2(n4343), .ZN(n4347) );
  INV_X1 U5370 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U5371 ( .A1(n5485), .A2(n4344), .ZN(n4345) );
  OR2_X1 U5372 ( .A1(n4650), .A2(n4345), .ZN(n4346) );
  INV_X1 U5373 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5508) );
  OAI22_X1 U5374 ( .A1(n6216), .A2(n5508), .B1(n4348), .B2(n6205), .ZN(n4349)
         );
  INV_X1 U5375 ( .A(n4349), .ZN(n4361) );
  INV_X1 U5376 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6771) );
  AND2_X1 U5377 ( .A1(n4350), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4351) );
  OAI22_X1 U5378 ( .A1(n5451), .A2(n6771), .B1(n5622), .B2(n6206), .ZN(n4352)
         );
  INV_X1 U5379 ( .A(n4352), .ZN(n4360) );
  OAI21_X1 U5380 ( .B1(n5448), .B2(n4355), .A(n4354), .ZN(n5620) );
  OR2_X1 U5381 ( .A1(n5453), .A2(n4356), .ZN(n4357) );
  AND2_X1 U5382 ( .A1(n5503), .A2(n4357), .ZN(n5737) );
  INV_X1 U5383 ( .A(n5737), .ZN(n5507) );
  OAI22_X1 U5384 ( .A1(n5620), .A2(n6167), .B1(n5507), .B2(n6200), .ZN(n4358)
         );
  INV_X1 U5385 ( .A(n4358), .ZN(n4359) );
  NAND4_X1 U5386 ( .A1(n4362), .A2(n4361), .A3(n4360), .A4(n4359), .ZN(U2803)
         );
  INV_X1 U5387 ( .A(n4363), .ZN(n4368) );
  INV_X1 U5388 ( .A(n4364), .ZN(n4366) );
  NAND2_X1 U5389 ( .A1(n4366), .A2(n3831), .ZN(n4367) );
  OAI22_X1 U5390 ( .A1(n6314), .A2(n5437), .B1(n6338), .B2(n6748), .ZN(n4369)
         );
  NAND2_X1 U5391 ( .A1(n4259), .A2(n4374), .ZN(n4375) );
  XNOR2_X1 U5392 ( .A(n4375), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5591)
         );
  INV_X1 U5393 ( .A(n5591), .ZN(n4376) );
  NAND2_X1 U5394 ( .A1(n4376), .A2(n6383), .ZN(n4388) );
  AOI21_X1 U5395 ( .B1(n4378), .B2(n5467), .A(n4377), .ZN(n4382) );
  INV_X1 U5396 ( .A(n4379), .ZN(n4380) );
  AOI21_X1 U5397 ( .B1(n4382), .B2(n4381), .A(n4380), .ZN(n5486) );
  OAI22_X1 U5398 ( .A1(n6793), .A2(n6338), .B1(n5704), .B2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4385) );
  INV_X1 U5399 ( .A(n4112), .ZN(n4537) );
  NAND2_X1 U5400 ( .A1(n5406), .A2(n4537), .ZN(n4390) );
  OAI21_X1 U5401 ( .B1(n5402), .B2(n5400), .A(n5398), .ZN(n4389) );
  NAND2_X1 U5402 ( .A1(n4390), .A2(n4389), .ZN(n5410) );
  NOR2_X1 U5403 ( .A1(n5410), .A2(n6545), .ZN(n4392) );
  INV_X1 U5404 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6804) );
  NOR2_X1 U5405 ( .A1(n5896), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U5406 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5248), .ZN(n4391) );
  OAI21_X1 U5407 ( .B1(n4392), .B2(n6804), .A(n4391), .ZN(U2790) );
  AOI21_X1 U5408 ( .B1(n4393), .B2(MEMORYFETCH_REG_SCAN_IN), .A(n5248), .ZN(
        n4394) );
  NAND2_X1 U5409 ( .A1(n4395), .A2(n4394), .ZN(U2788) );
  INV_X1 U5410 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4401) );
  OR2_X1 U5411 ( .A1(n5398), .A2(READY_N), .ZN(n4396) );
  INV_X1 U5412 ( .A(n4399), .ZN(n4397) );
  NAND2_X1 U5413 ( .A1(n4397), .A2(n6291), .ZN(n4449) );
  NAND2_X1 U5414 ( .A1(n4399), .A2(n4398), .ZN(n4543) );
  INV_X1 U5415 ( .A(DATAI_15_), .ZN(n6774) );
  INV_X1 U5416 ( .A(EAX_REG_15__SCAN_IN), .ZN(n4400) );
  OAI222_X1 U5417 ( .A1(n4401), .A2(n4449), .B1(n4543), .B2(n6774), .C1(n4400), 
        .C2(n6291), .ZN(U2954) );
  INV_X1 U5418 ( .A(LWORD_REG_10__SCAN_IN), .ZN(n4404) );
  INV_X1 U5419 ( .A(DATAI_10_), .ZN(n4403) );
  INV_X1 U5420 ( .A(EAX_REG_10__SCAN_IN), .ZN(n4402) );
  OAI222_X1 U5421 ( .A1(n4404), .A2(n4449), .B1(n4543), .B2(n4403), .C1(n4402), 
        .C2(n6291), .ZN(U2949) );
  INV_X1 U5422 ( .A(n6638), .ZN(n4407) );
  INV_X1 U5423 ( .A(n5100), .ZN(n4405) );
  OR2_X1 U5424 ( .A1(n6634), .A2(n4405), .ZN(n5409) );
  OAI21_X1 U5425 ( .B1(n5248), .B2(READREQUEST_REG_SCAN_IN), .A(n4407), .ZN(
        n4406) );
  OAI21_X1 U5426 ( .B1(n4407), .B2(n5409), .A(n4406), .ZN(U3474) );
  OAI21_X1 U5427 ( .B1(n4409), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4408), 
        .ZN(n6380) );
  XOR2_X1 U5428 ( .A(n4411), .B(n4410), .Z(n6336) );
  OAI222_X1 U5429 ( .A1(n6380), .A2(n5557), .B1(n5567), .B2(n4412), .C1(n6236), 
        .C2(n6336), .ZN(U2859) );
  NAND2_X1 U5430 ( .A1(n6636), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6621) );
  INV_X1 U5431 ( .A(n6621), .ZN(n4649) );
  INV_X1 U5432 ( .A(n4413), .ZN(n4414) );
  OAI22_X1 U5433 ( .A1(n6504), .A2(n6558), .B1(n4414), .B2(n5398), .ZN(n4415)
         );
  AOI21_X1 U5434 ( .B1(n4415), .B2(n6768), .A(n4540), .ZN(n4416) );
  OR2_X1 U5435 ( .A1(n5406), .A2(n4416), .ZN(n4422) );
  INV_X1 U5436 ( .A(n4535), .ZN(n4418) );
  OR2_X1 U5437 ( .A1(n4417), .A2(n4418), .ZN(n4419) );
  AND2_X1 U5438 ( .A1(n4420), .A2(n4419), .ZN(n4421) );
  NAND2_X1 U5439 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4529), .ZN(n6620) );
  INV_X1 U5440 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6802) );
  OAI22_X1 U5441 ( .A1(n6507), .A2(n6545), .B1(n6620), .B2(n6802), .ZN(n6053)
         );
  NOR2_X1 U5442 ( .A1(n4649), .A2(n6053), .ZN(n5842) );
  NOR2_X1 U5443 ( .A1(n4424), .A2(n4425), .ZN(n4435) );
  AND2_X1 U5444 ( .A1(n4428), .A2(n4104), .ZN(n4429) );
  AND2_X1 U5445 ( .A1(n4417), .A2(n4429), .ZN(n4431) );
  NAND2_X1 U5446 ( .A1(n4431), .A2(n4430), .ZN(n5373) );
  NAND2_X1 U5447 ( .A1(n4427), .A2(n5373), .ZN(n4433) );
  NOR2_X1 U5448 ( .A1(n6504), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4507)
         );
  INV_X1 U5449 ( .A(n4507), .ZN(n4432) );
  OAI211_X1 U5450 ( .C1(n4435), .C2(n4544), .A(n4433), .B(n4432), .ZN(n6502)
         );
  INV_X1 U5451 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4434) );
  AOI22_X1 U5452 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4434), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6378), .ZN(n5335) );
  NOR2_X1 U5453 ( .A1(n6542), .A2(n6371), .ZN(n5333) );
  INV_X1 U5454 ( .A(n4435), .ZN(n4436) );
  AOI222_X1 U5455 ( .A1(n6502), .A2(n6052), .B1(n5335), .B2(n5333), .C1(n4436), 
        .C2(n6534), .ZN(n4438) );
  NAND2_X1 U5456 ( .A1(n5842), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4437) );
  OAI21_X1 U5457 ( .B1(n5842), .B2(n4438), .A(n4437), .ZN(U3460) );
  OAI21_X1 U5458 ( .B1(n4441), .B2(n4440), .A(n4439), .ZN(n6228) );
  OR2_X1 U5459 ( .A1(n4443), .A2(n4442), .ZN(n4444) );
  NAND2_X1 U5460 ( .A1(n6233), .A2(n4444), .ZN(n6374) );
  INV_X1 U5461 ( .A(n6374), .ZN(n4446) );
  INV_X1 U5462 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4445) );
  OAI22_X1 U5463 ( .A1(n5557), .A2(n4446), .B1(n4445), .B2(n5567), .ZN(n4447)
         );
  INV_X1 U5464 ( .A(n4447), .ZN(n4448) );
  OAI21_X1 U5465 ( .B1(n6228), .B2(n6236), .A(n4448), .ZN(U2858) );
  INV_X2 U5466 ( .A(n4449), .ZN(n6289) );
  INV_X2 U5467 ( .A(n6291), .ZN(n4575) );
  AOI22_X1 U5468 ( .A1(n6289), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n4575), .ZN(n4451) );
  INV_X1 U5469 ( .A(DATAI_14_), .ZN(n4450) );
  OR2_X1 U5470 ( .A1(n4543), .A2(n4450), .ZN(n4459) );
  NAND2_X1 U5471 ( .A1(n4451), .A2(n4459), .ZN(U2953) );
  AOI22_X1 U5472 ( .A1(n6289), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n4575), .ZN(n4452) );
  NAND2_X1 U5473 ( .A1(n6288), .A2(DATAI_0_), .ZN(n4576) );
  NAND2_X1 U5474 ( .A1(n4452), .A2(n4576), .ZN(U2939) );
  AOI22_X1 U5475 ( .A1(n6289), .A2(LWORD_REG_4__SCAN_IN), .B1(n4575), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n4453) );
  NAND2_X1 U5476 ( .A1(n6288), .A2(DATAI_4_), .ZN(n4465) );
  NAND2_X1 U5477 ( .A1(n4453), .A2(n4465), .ZN(U2943) );
  AOI22_X1 U5478 ( .A1(n6289), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n4575), .ZN(n4454) );
  NAND2_X1 U5479 ( .A1(n6288), .A2(DATAI_8_), .ZN(n4585) );
  NAND2_X1 U5480 ( .A1(n4454), .A2(n4585), .ZN(U2932) );
  AOI22_X1 U5481 ( .A1(n6289), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n4575), .ZN(n4456) );
  INV_X1 U5482 ( .A(DATAI_13_), .ZN(n4455) );
  OR2_X1 U5483 ( .A1(n4543), .A2(n4455), .ZN(n4591) );
  NAND2_X1 U5484 ( .A1(n4456), .A2(n4591), .ZN(U2937) );
  AOI22_X1 U5485 ( .A1(n6289), .A2(UWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_27__SCAN_IN), .B2(n4575), .ZN(n4457) );
  NAND2_X1 U5486 ( .A1(n6288), .A2(DATAI_11_), .ZN(n4587) );
  NAND2_X1 U5487 ( .A1(n4457), .A2(n4587), .ZN(U2935) );
  AOI22_X1 U5488 ( .A1(n6289), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n4575), .ZN(n4458) );
  NAND2_X1 U5489 ( .A1(n6288), .A2(DATAI_5_), .ZN(n4578) );
  NAND2_X1 U5490 ( .A1(n4458), .A2(n4578), .ZN(U2929) );
  AOI22_X1 U5491 ( .A1(n6289), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n4575), .ZN(n4460) );
  NAND2_X1 U5492 ( .A1(n4460), .A2(n4459), .ZN(U2938) );
  AOI22_X1 U5493 ( .A1(n6289), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n4575), .ZN(n4461) );
  NAND2_X1 U5494 ( .A1(n6288), .A2(DATAI_2_), .ZN(n4593) );
  NAND2_X1 U5495 ( .A1(n4461), .A2(n4593), .ZN(U2926) );
  AOI22_X1 U5496 ( .A1(n6289), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n4575), .ZN(n4462) );
  NAND2_X1 U5497 ( .A1(n6288), .A2(DATAI_7_), .ZN(n4595) );
  NAND2_X1 U5498 ( .A1(n4462), .A2(n4595), .ZN(U2931) );
  AOI22_X1 U5499 ( .A1(n6289), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n4575), .ZN(n4463) );
  NAND2_X1 U5500 ( .A1(n6288), .A2(DATAI_6_), .ZN(n4589) );
  NAND2_X1 U5501 ( .A1(n4463), .A2(n4589), .ZN(U2930) );
  AOI22_X1 U5502 ( .A1(n6289), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n4575), .ZN(n4464) );
  NAND2_X1 U5503 ( .A1(n6288), .A2(DATAI_9_), .ZN(n4583) );
  NAND2_X1 U5504 ( .A1(n4464), .A2(n4583), .ZN(U2933) );
  AOI22_X1 U5505 ( .A1(n6289), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n4575), .ZN(n4466) );
  NAND2_X1 U5506 ( .A1(n4466), .A2(n4465), .ZN(U2928) );
  AOI22_X1 U5507 ( .A1(n6289), .A2(UWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_28__SCAN_IN), .B2(n4575), .ZN(n4467) );
  NAND2_X1 U5508 ( .A1(n6288), .A2(DATAI_12_), .ZN(n4597) );
  NAND2_X1 U5509 ( .A1(n4467), .A2(n4597), .ZN(U2936) );
  INV_X1 U5510 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4473) );
  NAND2_X1 U5511 ( .A1(n6504), .A2(n6531), .ZN(n4469) );
  INV_X1 U5512 ( .A(n6558), .ZN(n4468) );
  NAND2_X1 U5513 ( .A1(n4469), .A2(n4468), .ZN(n4470) );
  NAND2_X1 U5514 ( .A1(n4471), .A2(n2987), .ZN(n4616) );
  AND2_X2 U5515 ( .A1(n6636), .A2(n4529), .ZN(n6284) );
  AOI22_X1 U5516 ( .A1(n6284), .A2(UWORD_REG_8__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4472) );
  OAI21_X1 U5517 ( .B1(n4473), .B2(n4616), .A(n4472), .ZN(U2899) );
  AOI22_X1 U5518 ( .A1(n6284), .A2(UWORD_REG_9__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4474) );
  OAI21_X1 U5519 ( .B1(n3784), .B2(n4616), .A(n4474), .ZN(U2898) );
  INV_X1 U5520 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6292) );
  AOI22_X1 U5521 ( .A1(n6284), .A2(UWORD_REG_10__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4475) );
  OAI21_X1 U5522 ( .B1(n6292), .B2(n4616), .A(n4475), .ZN(U2897) );
  INV_X1 U5523 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4477) );
  AOI22_X1 U5524 ( .A1(n6284), .A2(UWORD_REG_14__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4476) );
  OAI21_X1 U5525 ( .B1(n4477), .B2(n4616), .A(n4476), .ZN(U2893) );
  AOI22_X1 U5526 ( .A1(n6284), .A2(UWORD_REG_11__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4478) );
  OAI21_X1 U5527 ( .B1(n3826), .B2(n4616), .A(n4478), .ZN(U2896) );
  INV_X1 U5528 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4480) );
  AOI22_X1 U5529 ( .A1(n6284), .A2(UWORD_REG_12__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4479) );
  OAI21_X1 U5530 ( .B1(n4480), .B2(n4616), .A(n4479), .ZN(U2895) );
  AOI22_X1 U5531 ( .A1(n6284), .A2(UWORD_REG_13__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4481) );
  OAI21_X1 U5532 ( .B1(n3869), .B2(n4616), .A(n4481), .ZN(U2894) );
  NAND2_X1 U5533 ( .A1(n6399), .A2(n5373), .ZN(n4499) );
  INV_X1 U5534 ( .A(n4540), .ZN(n4483) );
  NAND2_X1 U5535 ( .A1(n5405), .A2(n4483), .ZN(n4505) );
  INV_X1 U5536 ( .A(n4484), .ZN(n5331) );
  AOI21_X1 U5537 ( .B1(n5331), .B2(n3076), .A(n4485), .ZN(n4487) );
  NAND3_X1 U5538 ( .A1(n4505), .A2(n4487), .A3(n3378), .ZN(n4497) );
  AOI21_X1 U5539 ( .B1(n4488), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n4491), 
        .ZN(n4494) );
  AND2_X1 U5540 ( .A1(n4506), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4490)
         );
  NOR2_X1 U5541 ( .A1(n4491), .A2(n4490), .ZN(n4492) );
  AND3_X1 U5542 ( .A1(n4493), .A2(n3250), .A3(n4492), .ZN(n5839) );
  OAI22_X1 U5543 ( .A1(n6504), .A2(n4494), .B1(n5839), .B2(n4512), .ZN(n4495)
         );
  AOI21_X1 U5544 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n4507), .A(n4495), 
        .ZN(n4496) );
  AND2_X1 U5545 ( .A1(n4497), .A2(n4496), .ZN(n4498) );
  NAND2_X1 U5546 ( .A1(n4499), .A2(n4498), .ZN(n5837) );
  INV_X1 U5547 ( .A(n6507), .ZN(n4500) );
  NAND2_X1 U5548 ( .A1(n5837), .A2(n4500), .ZN(n4502) );
  NAND2_X1 U5549 ( .A1(n6507), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4501) );
  NAND2_X1 U5550 ( .A1(n4502), .A2(n4501), .ZN(n6518) );
  XNOR2_X1 U5551 ( .A(n4484), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4513)
         );
  NAND2_X1 U5552 ( .A1(n4505), .A2(n4513), .ZN(n4511) );
  NOR2_X1 U5553 ( .A1(n6504), .A2(n4506), .ZN(n4508) );
  MUX2_X1 U5554 ( .A(n4508), .B(n4507), .S(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .Z(n4509) );
  INV_X1 U5555 ( .A(n4509), .ZN(n4510) );
  OAI211_X1 U5556 ( .C1(n4513), .C2(n4512), .A(n4511), .B(n4510), .ZN(n4514)
         );
  AOI21_X1 U5557 ( .B1(n4504), .B2(n5373), .A(n4514), .ZN(n5332) );
  OR2_X1 U5558 ( .A1(n5332), .A2(n6507), .ZN(n4516) );
  NAND2_X1 U5559 ( .A1(n6507), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4515) );
  NAND2_X1 U5560 ( .A1(n4516), .A2(n4515), .ZN(n6513) );
  NAND3_X1 U5561 ( .A1(n6518), .A2(n6542), .A3(n6513), .ZN(n4519) );
  NOR2_X1 U5562 ( .A1(FLUSH_REG_SCAN_IN), .A2(n6542), .ZN(n4517) );
  NAND2_X1 U5563 ( .A1(n4485), .A2(n4517), .ZN(n4518) );
  NAND2_X1 U5564 ( .A1(n4519), .A2(n4518), .ZN(n6527) );
  INV_X1 U5565 ( .A(n4520), .ZN(n4527) );
  INV_X1 U5566 ( .A(n4873), .ZN(n4521) );
  OR2_X1 U5567 ( .A1(n4522), .A2(n4521), .ZN(n4523) );
  XNOR2_X1 U5568 ( .A(n4523), .B(n6057), .ZN(n6186) );
  OR2_X1 U5569 ( .A1(n4417), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4526) );
  MUX2_X1 U5570 ( .A(n6802), .B(n6507), .S(n6542), .Z(n4524) );
  NAND2_X1 U5571 ( .A1(n4524), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4525) );
  OAI21_X1 U5572 ( .B1(n6186), .B2(n4526), .A(n4525), .ZN(n6526) );
  AOI21_X1 U5573 ( .B1(n6527), .B2(n4527), .A(n6526), .ZN(n4530) );
  AOI21_X1 U5574 ( .B1(n4530), .B2(n6802), .A(n6620), .ZN(n4528) );
  NAND2_X1 U5575 ( .A1(n4530), .A2(n4529), .ZN(n6541) );
  INV_X1 U5576 ( .A(n6541), .ZN(n4532) );
  INV_X1 U5577 ( .A(n3358), .ZN(n5044) );
  AND2_X1 U5578 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6623), .ZN(n5833) );
  OAI22_X1 U5579 ( .A1(n5052), .A2(n5896), .B1(n5044), .B2(n5833), .ZN(n4531)
         );
  OAI21_X1 U5580 ( .B1(n4532), .B2(n4531), .A(n6393), .ZN(n4533) );
  OAI21_X1 U5581 ( .B1(n6393), .B2(n6401), .A(n4533), .ZN(U3465) );
  INV_X1 U5582 ( .A(n4534), .ZN(n4541) );
  NAND2_X1 U5583 ( .A1(n6539), .A2(n4535), .ZN(n4538) );
  OAI22_X1 U5584 ( .A1(n4417), .A2(n4538), .B1(n4537), .B2(n4536), .ZN(n4539)
         );
  NAND2_X1 U5585 ( .A1(n4544), .A2(n5391), .ZN(n4545) );
  INV_X1 U5586 ( .A(n4545), .ZN(n4546) );
  INV_X1 U5587 ( .A(n5583), .ZN(n4739) );
  INV_X1 U5588 ( .A(DATAI_0_), .ZN(n6818) );
  INV_X1 U5589 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6287) );
  OAI222_X1 U5590 ( .A1(n5988), .A2(n6336), .B1(n4739), .B2(n6818), .C1(n5394), 
        .C2(n6287), .ZN(U2891) );
  INV_X1 U5591 ( .A(DATAI_1_), .ZN(n4656) );
  INV_X1 U5592 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6282) );
  OAI222_X1 U5593 ( .A1(n6228), .A2(n5988), .B1(n4739), .B2(n4656), .C1(n5394), 
        .C2(n6282), .ZN(U2890) );
  OAI21_X1 U5594 ( .B1(n4549), .B2(n4548), .A(n4547), .ZN(n6373) );
  AOI22_X1 U5595 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6376), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4552) );
  INV_X1 U5596 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4550) );
  NAND2_X1 U5597 ( .A1(n6310), .A2(n4550), .ZN(n4551) );
  OAI211_X1 U5598 ( .C1(n6373), .C2(n6297), .A(n4552), .B(n4551), .ZN(n4553)
         );
  INV_X1 U5599 ( .A(n4553), .ZN(n4554) );
  OAI21_X1 U5600 ( .B1(n6335), .B2(n6228), .A(n4554), .ZN(U2985) );
  XNOR2_X1 U5601 ( .A(n4555), .B(n4556), .ZN(n4573) );
  INV_X1 U5602 ( .A(n4557), .ZN(n6357) );
  AOI21_X1 U5603 ( .B1(n6359), .B2(n6357), .A(n6372), .ZN(n5166) );
  NOR2_X1 U5604 ( .A1(n4708), .A2(n5166), .ZN(n4706) );
  NAND2_X1 U5605 ( .A1(n4706), .A2(n3912), .ZN(n4562) );
  INV_X1 U5606 ( .A(n6370), .ZN(n5315) );
  OAI21_X1 U5607 ( .B1(n5768), .B2(n6359), .A(n5315), .ZN(n4707) );
  INV_X1 U5608 ( .A(n4707), .ZN(n6366) );
  NAND2_X1 U5609 ( .A1(n6372), .A2(n4708), .ZN(n6361) );
  NAND2_X1 U5610 ( .A1(n6366), .A2(n6361), .ZN(n4625) );
  NAND2_X1 U5611 ( .A1(n4633), .A2(n4558), .ZN(n4559) );
  NAND2_X1 U5612 ( .A1(n4622), .A2(n4559), .ZN(n5235) );
  INV_X1 U5613 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6573) );
  OAI22_X1 U5614 ( .A1(n6339), .A2(n5235), .B1(n6573), .B2(n6338), .ZN(n4560)
         );
  AOI21_X1 U5615 ( .B1(n4625), .B2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n4560), 
        .ZN(n4561) );
  OAI211_X1 U5616 ( .C1(n4573), .C2(n6035), .A(n4562), .B(n4561), .ZN(U3015)
         );
  NAND2_X1 U5617 ( .A1(n4564), .A2(n4565), .ZN(n4566) );
  AND2_X1 U5618 ( .A1(n4563), .A2(n4566), .ZN(n4574) );
  INV_X1 U5619 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4567) );
  OAI22_X1 U5620 ( .A1(n5557), .A2(n5235), .B1(n4567), .B2(n5567), .ZN(n4568)
         );
  AOI21_X1 U5621 ( .B1(n4574), .B2(n4283), .A(n4568), .ZN(n4569) );
  INV_X1 U5622 ( .A(n4569), .ZN(U2856) );
  AOI22_X1 U5623 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n6376), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n4570) );
  OAI21_X1 U5624 ( .B1(n5236), .B2(n6324), .A(n4570), .ZN(n4571) );
  AOI21_X1 U5625 ( .B1(n4574), .B2(n6319), .A(n4571), .ZN(n4572) );
  OAI21_X1 U5626 ( .B1(n4573), .B2(n6297), .A(n4572), .ZN(U2983) );
  INV_X1 U5627 ( .A(n4574), .ZN(n5240) );
  INV_X1 U5628 ( .A(DATAI_3_), .ZN(n6712) );
  INV_X1 U5629 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6278) );
  OAI222_X1 U5630 ( .A1(n5240), .A2(n5988), .B1(n4739), .B2(n6712), .C1(n5394), 
        .C2(n6278), .ZN(U2888) );
  AOI22_X1 U5631 ( .A1(n6289), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n4575), .ZN(n4577) );
  NAND2_X1 U5632 ( .A1(n4577), .A2(n4576), .ZN(U2924) );
  AOI22_X1 U5633 ( .A1(n6289), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n4575), .ZN(n4579) );
  NAND2_X1 U5634 ( .A1(n4579), .A2(n4578), .ZN(U2944) );
  AOI22_X1 U5635 ( .A1(n6289), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n4575), .ZN(n4580) );
  NAND2_X1 U5636 ( .A1(n6288), .A2(DATAI_3_), .ZN(n4581) );
  NAND2_X1 U5637 ( .A1(n4580), .A2(n4581), .ZN(U2927) );
  AOI22_X1 U5638 ( .A1(n6289), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n4575), .ZN(n4582) );
  NAND2_X1 U5639 ( .A1(n4582), .A2(n4581), .ZN(U2942) );
  AOI22_X1 U5640 ( .A1(n6289), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n4575), .ZN(n4584) );
  NAND2_X1 U5641 ( .A1(n4584), .A2(n4583), .ZN(U2948) );
  AOI22_X1 U5642 ( .A1(n6289), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n4575), .ZN(n4586) );
  NAND2_X1 U5643 ( .A1(n4586), .A2(n4585), .ZN(U2947) );
  AOI22_X1 U5644 ( .A1(n6289), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n4575), .ZN(n4588) );
  NAND2_X1 U5645 ( .A1(n4588), .A2(n4587), .ZN(U2950) );
  AOI22_X1 U5646 ( .A1(n6289), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n4575), .ZN(n4590) );
  NAND2_X1 U5647 ( .A1(n4590), .A2(n4589), .ZN(U2945) );
  AOI22_X1 U5648 ( .A1(n6289), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n4575), .ZN(n4592) );
  NAND2_X1 U5649 ( .A1(n4592), .A2(n4591), .ZN(U2952) );
  AOI22_X1 U5650 ( .A1(n6289), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n4575), .ZN(n4594) );
  NAND2_X1 U5651 ( .A1(n4594), .A2(n4593), .ZN(U2941) );
  AOI22_X1 U5652 ( .A1(n6289), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n4575), .ZN(n4596) );
  NAND2_X1 U5653 ( .A1(n4596), .A2(n4595), .ZN(U2946) );
  AOI22_X1 U5654 ( .A1(n6289), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n4575), .ZN(n4598) );
  NAND2_X1 U5655 ( .A1(n4598), .A2(n4597), .ZN(U2951) );
  AOI22_X1 U5656 ( .A1(n6289), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n4575), .ZN(n4599) );
  NAND2_X1 U5657 ( .A1(n6288), .A2(DATAI_1_), .ZN(n4600) );
  NAND2_X1 U5658 ( .A1(n4599), .A2(n4600), .ZN(U2940) );
  AOI22_X1 U5659 ( .A1(n6289), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n4575), .ZN(n4601) );
  NAND2_X1 U5660 ( .A1(n4601), .A2(n4600), .ZN(U2925) );
  AOI22_X1 U5661 ( .A1(n6284), .A2(UWORD_REG_7__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4602) );
  OAI21_X1 U5662 ( .B1(n3742), .B2(n4616), .A(n4602), .ZN(U2900) );
  INV_X1 U5663 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4604) );
  AOI22_X1 U5664 ( .A1(n6284), .A2(UWORD_REG_6__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4603) );
  OAI21_X1 U5665 ( .B1(n4604), .B2(n4616), .A(n4603), .ZN(U2901) );
  INV_X1 U5666 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4606) );
  AOI22_X1 U5667 ( .A1(n6284), .A2(UWORD_REG_2__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4605) );
  OAI21_X1 U5668 ( .B1(n4606), .B2(n4616), .A(n4605), .ZN(U2905) );
  INV_X1 U5669 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4608) );
  AOI22_X1 U5670 ( .A1(n6284), .A2(UWORD_REG_1__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4607) );
  OAI21_X1 U5671 ( .B1(n4608), .B2(n4616), .A(n4607), .ZN(U2906) );
  INV_X1 U5672 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4610) );
  AOI22_X1 U5673 ( .A1(n6284), .A2(UWORD_REG_5__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4609) );
  OAI21_X1 U5674 ( .B1(n4610), .B2(n4616), .A(n4609), .ZN(U2902) );
  INV_X1 U5675 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4612) );
  AOI22_X1 U5676 ( .A1(n6284), .A2(UWORD_REG_3__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4611) );
  OAI21_X1 U5677 ( .B1(n4612), .B2(n4616), .A(n4611), .ZN(U2904) );
  INV_X1 U5678 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4614) );
  AOI22_X1 U5679 ( .A1(n6284), .A2(UWORD_REG_0__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4613) );
  OAI21_X1 U5680 ( .B1(n4614), .B2(n4616), .A(n4613), .ZN(U2907) );
  INV_X1 U5681 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4617) );
  AOI22_X1 U5682 ( .A1(n6284), .A2(UWORD_REG_4__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4615) );
  OAI21_X1 U5683 ( .B1(n4617), .B2(n4616), .A(n4615), .ZN(U2903) );
  XNOR2_X1 U5684 ( .A(n4618), .B(n4620), .ZN(n4701) );
  NAND2_X1 U5685 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4709) );
  OAI211_X1 U5686 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4706), .B(n4709), .ZN(n4627) );
  INV_X1 U5687 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6188) );
  NOR2_X1 U5688 ( .A1(n6338), .A2(n6188), .ZN(n4697) );
  AND2_X1 U5689 ( .A1(n4622), .A2(n4621), .ZN(n4623) );
  OR2_X1 U5690 ( .A1(n4623), .A2(n4705), .ZN(n6199) );
  NOR2_X1 U5691 ( .A1(n6339), .A2(n6199), .ZN(n4624) );
  AOI211_X1 U5692 ( .C1(n4625), .C2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4697), 
        .B(n4624), .ZN(n4626) );
  OAI211_X1 U5693 ( .C1(n6035), .C2(n4701), .A(n4627), .B(n4626), .ZN(U3014)
         );
  INV_X1 U5694 ( .A(n4628), .ZN(n4629) );
  AOI21_X1 U5695 ( .B1(n4629), .B2(n4439), .A(n3399), .ZN(n6320) );
  NAND2_X1 U5696 ( .A1(n4631), .A2(n4630), .ZN(n4632) );
  AND2_X1 U5697 ( .A1(n4633), .A2(n4632), .ZN(n6358) );
  INV_X1 U5698 ( .A(n6358), .ZN(n6201) );
  OAI22_X1 U5699 ( .A1(n5557), .A2(n6201), .B1(n6215), .B2(n5567), .ZN(n4634)
         );
  AOI21_X1 U5700 ( .B1(n6320), .B2(n4283), .A(n4634), .ZN(n4635) );
  INV_X1 U5701 ( .A(n4635), .ZN(U2857) );
  INV_X1 U5702 ( .A(n6320), .ZN(n4636) );
  INV_X1 U5703 ( .A(DATAI_2_), .ZN(n4676) );
  INV_X1 U5704 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6280) );
  OAI222_X1 U5705 ( .A1(n4636), .A2(n5988), .B1(n4739), .B2(n4676), .C1(n5394), 
        .C2(n6280), .ZN(U2889) );
  NAND2_X1 U5706 ( .A1(n5821), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5825) );
  OAI21_X1 U5707 ( .B1(n5105), .B2(n5825), .A(n6408), .ZN(n4644) );
  INV_X1 U5708 ( .A(n4427), .ZN(n5823) );
  OR2_X1 U5709 ( .A1(n4504), .A2(n5823), .ZN(n5109) );
  INV_X1 U5710 ( .A(n5109), .ZN(n4640) );
  NOR2_X1 U5711 ( .A1(n5110), .A2(n6517), .ZN(n6491) );
  AOI21_X1 U5712 ( .B1(n5901), .B2(n3358), .A(n6491), .ZN(n4641) );
  NAND3_X1 U5713 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6512), .ZN(n5900) );
  OAI22_X1 U5714 ( .A1(n4644), .A2(n4641), .B1(n5900), .B2(n6633), .ZN(n6495)
         );
  INV_X1 U5715 ( .A(n6495), .ZN(n4693) );
  INV_X1 U5716 ( .A(n4641), .ZN(n4643) );
  INV_X1 U5717 ( .A(n5020), .ZN(n5112) );
  AOI21_X1 U5718 ( .B1(n5896), .B2(n5900), .A(n5112), .ZN(n4642) );
  OAI21_X1 U5719 ( .B1(n4644), .B2(n4643), .A(n4642), .ZN(n6497) );
  INV_X1 U5720 ( .A(DATAI_24_), .ZN(n4645) );
  OR2_X1 U5721 ( .A1(n6335), .A2(n4645), .ZN(n5123) );
  INV_X1 U5722 ( .A(n5117), .ZN(n4646) );
  NAND2_X1 U5723 ( .A1(n5821), .A2(n5016), .ZN(n4869) );
  NOR2_X2 U5724 ( .A1(n5105), .A2(n4869), .ZN(n6494) );
  INV_X1 U5725 ( .A(DATAI_16_), .ZN(n4647) );
  OR2_X1 U5726 ( .A1(n6335), .A2(n4647), .ZN(n6415) );
  INV_X1 U5727 ( .A(n6415), .ZN(n5851) );
  NOR2_X2 U5728 ( .A1(n4719), .A2(n4650), .ZN(n6402) );
  AOI22_X1 U5729 ( .A1(n6494), .A2(n5851), .B1(n6402), .B2(n6491), .ZN(n4651)
         );
  OAI21_X1 U5730 ( .B1(n5123), .B2(n6500), .A(n4651), .ZN(n4652) );
  AOI21_X1 U5731 ( .B1(INSTQUEUE_REG_11__0__SCAN_IN), .B2(n6497), .A(n4652), 
        .ZN(n4653) );
  OAI21_X1 U5732 ( .B1(n4693), .B2(n5910), .A(n4653), .ZN(U3108) );
  NAND2_X1 U5733 ( .A1(n6399), .A2(n3358), .ZN(n4840) );
  NAND2_X1 U5734 ( .A1(n4504), .A2(n4427), .ZN(n4771) );
  OR2_X1 U5735 ( .A1(n4840), .A2(n4771), .ZN(n4654) );
  AND2_X1 U5736 ( .A1(n4654), .A2(n4732), .ZN(n4659) );
  INV_X1 U5737 ( .A(n4659), .ZN(n4655) );
  AOI22_X1 U5738 ( .A1(n4655), .A2(n6408), .B1(n4773), .B2(
        STATE2_REG_2__SCAN_IN), .ZN(n4737) );
  NOR2_X2 U5739 ( .A1(n4656), .A2(n4806), .ZN(n6463) );
  INV_X1 U5740 ( .A(n6463), .ZN(n5914) );
  INV_X1 U5741 ( .A(n5821), .ZN(n4657) );
  NOR3_X1 U5742 ( .A1(n5826), .A2(n4769), .A3(n4657), .ZN(n4658) );
  AND2_X1 U5743 ( .A1(n6408), .A2(n6822), .ZN(n5844) );
  INV_X1 U5744 ( .A(n5844), .ZN(n5834) );
  OAI21_X1 U5745 ( .B1(n4658), .B2(n6335), .A(n5834), .ZN(n4660) );
  NAND2_X1 U5746 ( .A1(n4660), .A2(n4659), .ZN(n4661) );
  OAI211_X1 U5747 ( .C1(n4773), .C2(n6408), .A(n5020), .B(n4661), .ZN(n4730)
         );
  NAND2_X1 U5748 ( .A1(n4730), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4668)
         );
  INV_X1 U5749 ( .A(DATAI_25_), .ZN(n4662) );
  OR2_X1 U5750 ( .A1(n6335), .A2(n4662), .ZN(n6466) );
  INV_X1 U5751 ( .A(n6466), .ZN(n6416) );
  NAND3_X1 U5752 ( .A1(n5107), .A2(n5117), .A3(n4663), .ZN(n4800) );
  INV_X1 U5753 ( .A(n4800), .ZN(n4734) );
  NOR2_X2 U5754 ( .A1(n4719), .A2(n2986), .ZN(n6461) );
  INV_X1 U5755 ( .A(n6461), .ZN(n5062) );
  INV_X1 U5756 ( .A(DATAI_17_), .ZN(n4664) );
  OR2_X1 U5757 ( .A1(n6335), .A2(n4664), .ZN(n6419) );
  AND3_X1 U5758 ( .A1(n5821), .A2(n5016), .A3(n4663), .ZN(n4665) );
  OAI22_X1 U5759 ( .A1(n5062), .A2(n4732), .B1(n6419), .B2(n4731), .ZN(n4666)
         );
  AOI21_X1 U5760 ( .B1(n6416), .B2(n4734), .A(n4666), .ZN(n4667) );
  OAI211_X1 U5761 ( .C1(n4737), .C2(n5914), .A(n4668), .B(n4667), .ZN(U3141)
         );
  NAND2_X1 U5762 ( .A1(n4730), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4671)
         );
  INV_X1 U5763 ( .A(n5123), .ZN(n6412) );
  INV_X1 U5764 ( .A(n6402), .ZN(n5054) );
  OAI22_X1 U5765 ( .A1(n5054), .A2(n4732), .B1(n6415), .B2(n4731), .ZN(n4669)
         );
  AOI21_X1 U5766 ( .B1(n6412), .B2(n4734), .A(n4669), .ZN(n4670) );
  OAI211_X1 U5767 ( .C1(n4737), .C2(n5910), .A(n4671), .B(n4670), .ZN(U3140)
         );
  INV_X1 U5768 ( .A(n6475), .ZN(n5922) );
  NAND2_X1 U5769 ( .A1(n4730), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4675)
         );
  INV_X1 U5770 ( .A(DATAI_27_), .ZN(n6799) );
  OR2_X1 U5771 ( .A1(n6335), .A2(n6799), .ZN(n6478) );
  INV_X1 U5772 ( .A(n6478), .ZN(n6424) );
  NOR2_X2 U5773 ( .A1(n4719), .A2(n4672), .ZN(n6473) );
  INV_X1 U5774 ( .A(n6473), .ZN(n5066) );
  OR2_X1 U5775 ( .A1(n6335), .A2(n6680), .ZN(n6427) );
  OAI22_X1 U5776 ( .A1(n5066), .A2(n4732), .B1(n6427), .B2(n4731), .ZN(n4673)
         );
  AOI21_X1 U5777 ( .B1(n6424), .B2(n4734), .A(n4673), .ZN(n4674) );
  OAI211_X1 U5778 ( .C1(n4737), .C2(n5922), .A(n4675), .B(n4674), .ZN(U3143)
         );
  INV_X1 U5779 ( .A(n6469), .ZN(n5918) );
  NAND2_X1 U5780 ( .A1(n4730), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4680)
         );
  INV_X1 U5781 ( .A(DATAI_26_), .ZN(n6807) );
  OR2_X1 U5782 ( .A1(n6335), .A2(n6807), .ZN(n6472) );
  INV_X1 U5783 ( .A(n6472), .ZN(n6420) );
  NOR2_X2 U5784 ( .A1(n4719), .A2(n3207), .ZN(n6467) );
  INV_X1 U5785 ( .A(n6467), .ZN(n5084) );
  INV_X1 U5786 ( .A(DATAI_18_), .ZN(n4677) );
  OR2_X1 U5787 ( .A1(n6335), .A2(n4677), .ZN(n6423) );
  OAI22_X1 U5788 ( .A1(n5084), .A2(n4732), .B1(n6423), .B2(n4731), .ZN(n4678)
         );
  AOI21_X1 U5789 ( .B1(n6420), .B2(n4734), .A(n4678), .ZN(n4679) );
  OAI211_X1 U5790 ( .C1(n4737), .C2(n5918), .A(n4680), .B(n4679), .ZN(U3142)
         );
  INV_X1 U5791 ( .A(DATAI_7_), .ZN(n6662) );
  INV_X1 U5792 ( .A(n6496), .ZN(n5941) );
  NAND2_X1 U5793 ( .A1(n4730), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4684)
         );
  INV_X1 U5794 ( .A(DATAI_31_), .ZN(n6801) );
  OR2_X1 U5795 ( .A1(n6335), .A2(n6801), .ZN(n6501) );
  INV_X1 U5796 ( .A(n6501), .ZN(n6444) );
  NOR2_X2 U5797 ( .A1(n4719), .A2(n4295), .ZN(n6492) );
  INV_X1 U5798 ( .A(n6492), .ZN(n5058) );
  INV_X1 U5799 ( .A(DATAI_23_), .ZN(n4681) );
  OR2_X1 U5800 ( .A1(n6335), .A2(n4681), .ZN(n6449) );
  OAI22_X1 U5801 ( .A1(n5058), .A2(n4732), .B1(n6449), .B2(n4731), .ZN(n4682)
         );
  AOI21_X1 U5802 ( .B1(n6444), .B2(n4734), .A(n4682), .ZN(n4683) );
  OAI211_X1 U5803 ( .C1(n4737), .C2(n5941), .A(n4684), .B(n4683), .ZN(U3147)
         );
  AOI21_X1 U5804 ( .B1(n4686), .B2(n4563), .A(n4685), .ZN(n4738) );
  OAI22_X1 U5805 ( .A1(n5557), .A2(n6199), .B1(n6191), .B2(n5567), .ZN(n4687)
         );
  AOI21_X1 U5806 ( .B1(n4738), .B2(n4283), .A(n4687), .ZN(n4688) );
  INV_X1 U5807 ( .A(n4688), .ZN(U2855) );
  INV_X1 U5808 ( .A(DATAI_6_), .ZN(n6777) );
  INV_X1 U5809 ( .A(DATAI_30_), .ZN(n6769) );
  OR2_X1 U5810 ( .A1(n6335), .A2(n6769), .ZN(n5132) );
  INV_X1 U5811 ( .A(DATAI_22_), .ZN(n4689) );
  OR2_X1 U5812 ( .A1(n6335), .A2(n4689), .ZN(n6441) );
  INV_X1 U5813 ( .A(n6441), .ZN(n5881) );
  NOR2_X2 U5814 ( .A1(n4719), .A2(n3225), .ZN(n6436) );
  AOI22_X1 U5815 ( .A1(n6494), .A2(n5881), .B1(n6436), .B2(n6491), .ZN(n4690)
         );
  OAI21_X1 U5816 ( .B1(n5132), .B2(n6500), .A(n4690), .ZN(n4691) );
  AOI21_X1 U5817 ( .B1(INSTQUEUE_REG_11__6__SCAN_IN), .B2(n6497), .A(n4691), 
        .ZN(n4692) );
  OAI21_X1 U5818 ( .B1(n4693), .B2(n5934), .A(n4692), .ZN(U3114) );
  INV_X1 U5819 ( .A(DATAI_4_), .ZN(n6715) );
  INV_X1 U5820 ( .A(n6481), .ZN(n5926) );
  NAND2_X1 U5821 ( .A1(n4730), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4696)
         );
  INV_X1 U5822 ( .A(DATAI_28_), .ZN(n6682) );
  OR2_X1 U5823 ( .A1(n6335), .A2(n6682), .ZN(n6484) );
  INV_X1 U5824 ( .A(n6484), .ZN(n6428) );
  NOR2_X2 U5825 ( .A1(n4719), .A2(n3313), .ZN(n6479) );
  INV_X1 U5826 ( .A(n6479), .ZN(n5074) );
  OR2_X1 U5827 ( .A1(n6335), .A2(n6789), .ZN(n6431) );
  OAI22_X1 U5828 ( .A1(n5074), .A2(n4732), .B1(n6431), .B2(n4731), .ZN(n4694)
         );
  AOI21_X1 U5829 ( .B1(n6428), .B2(n4734), .A(n4694), .ZN(n4695) );
  OAI211_X1 U5830 ( .C1(n4737), .C2(n5926), .A(n4696), .B(n4695), .ZN(U3144)
         );
  AOI21_X1 U5831 ( .B1(n6330), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n4697), 
        .ZN(n4698) );
  OAI21_X1 U5832 ( .B1(n6193), .B2(n6324), .A(n4698), .ZN(n4699) );
  AOI21_X1 U5833 ( .B1(n4738), .B2(n6319), .A(n4699), .ZN(n4700) );
  OAI21_X1 U5834 ( .B1(n6297), .B2(n4701), .A(n4700), .ZN(U2982) );
  XNOR2_X1 U5835 ( .A(n4702), .B(n4703), .ZN(n6307) );
  OAI21_X1 U5836 ( .B1(n4705), .B2(n4704), .A(n4741), .ZN(n4716) );
  INV_X1 U5837 ( .A(n4716), .ZN(n6176) );
  NAND2_X1 U5838 ( .A1(n6376), .A2(REIP_REG_5__SCAN_IN), .ZN(n6312) );
  INV_X1 U5839 ( .A(n6312), .ZN(n4711) );
  INV_X1 U5840 ( .A(n4706), .ZN(n4909) );
  AOI221_X1 U5841 ( .B1(n4708), .B2(n6369), .C1(n4910), .C2(n6369), .A(n4707), 
        .ZN(n4911) );
  AOI221_X1 U5842 ( .B1(n4709), .B2(n3951), .C1(n4909), .C2(n3951), .A(n4911), 
        .ZN(n4710) );
  AOI211_X1 U5843 ( .C1(n6382), .C2(n6176), .A(n4711), .B(n4710), .ZN(n4712)
         );
  OAI21_X1 U5844 ( .B1(n6035), .B2(n6307), .A(n4712), .ZN(U3013) );
  OR2_X1 U5845 ( .A1(n4685), .A2(n4713), .ZN(n4715) );
  CLKBUF_X1 U5846 ( .A(n4714), .Z(n4727) );
  AND2_X1 U5847 ( .A1(n4715), .A2(n4727), .ZN(n6309) );
  INV_X1 U5848 ( .A(n6309), .ZN(n4718) );
  INV_X2 U5849 ( .A(n5569), .ZN(n5557) );
  OAI222_X1 U5850 ( .A1(n4718), .A2(n6236), .B1(n5567), .B2(n4717), .C1(n5557), 
        .C2(n4716), .ZN(U2854) );
  INV_X1 U5851 ( .A(DATAI_5_), .ZN(n6785) );
  INV_X1 U5852 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6273) );
  OAI222_X1 U5853 ( .A1(n4718), .A2(n5988), .B1(n4739), .B2(n6785), .C1(n5394), 
        .C2(n6273), .ZN(U2886) );
  NOR2_X2 U5854 ( .A1(n6785), .A2(n4806), .ZN(n6487) );
  INV_X1 U5855 ( .A(n6487), .ZN(n5930) );
  NAND2_X1 U5856 ( .A1(n4730), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4723)
         );
  INV_X1 U5857 ( .A(DATAI_29_), .ZN(n6772) );
  OR2_X1 U5858 ( .A1(n6335), .A2(n6772), .ZN(n6490) );
  INV_X1 U5859 ( .A(n6490), .ZN(n6432) );
  NOR2_X2 U5860 ( .A1(n4719), .A2(n5392), .ZN(n6485) );
  INV_X1 U5861 ( .A(n6485), .ZN(n5078) );
  INV_X1 U5862 ( .A(DATAI_21_), .ZN(n4720) );
  OR2_X1 U5863 ( .A1(n6335), .A2(n4720), .ZN(n6435) );
  OAI22_X1 U5864 ( .A1(n5078), .A2(n4732), .B1(n6435), .B2(n4731), .ZN(n4721)
         );
  AOI21_X1 U5865 ( .B1(n6432), .B2(n4734), .A(n4721), .ZN(n4722) );
  OAI211_X1 U5866 ( .C1(n4737), .C2(n5930), .A(n4723), .B(n4722), .ZN(U3145)
         );
  CLKBUF_X1 U5867 ( .A(n4724), .Z(n5007) );
  INV_X1 U5868 ( .A(n4725), .ZN(n4726) );
  NAND2_X1 U5869 ( .A1(n4727), .A2(n4726), .ZN(n4728) );
  NAND2_X1 U5870 ( .A1(n5007), .A2(n4728), .ZN(n6168) );
  INV_X2 U5871 ( .A(n5394), .ZN(n6250) );
  AOI22_X1 U5872 ( .A1(n5583), .A2(DATAI_6_), .B1(n6250), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n4729) );
  OAI21_X1 U5873 ( .B1(n6168), .B2(n5988), .A(n4729), .ZN(U2885) );
  NAND2_X1 U5874 ( .A1(n4730), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4736)
         );
  INV_X1 U5875 ( .A(n5132), .ZN(n6438) );
  INV_X1 U5876 ( .A(n6436), .ZN(n5070) );
  OAI22_X1 U5877 ( .A1(n5070), .A2(n4732), .B1(n6441), .B2(n4731), .ZN(n4733)
         );
  AOI21_X1 U5878 ( .B1(n6438), .B2(n4734), .A(n4733), .ZN(n4735) );
  OAI211_X1 U5879 ( .C1(n4737), .C2(n5934), .A(n4736), .B(n4735), .ZN(U3146)
         );
  INV_X1 U5880 ( .A(n4738), .ZN(n6194) );
  INV_X1 U5881 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6276) );
  OAI222_X1 U5882 ( .A1(n5988), .A2(n6194), .B1(n5394), .B2(n6276), .C1(n4739), 
        .C2(n6715), .ZN(U2887) );
  XOR2_X1 U5883 ( .A(n4741), .B(n4740), .Z(n6171) );
  INV_X1 U5884 ( .A(n6171), .ZN(n4743) );
  OAI222_X1 U5885 ( .A1(n6168), .A2(n6236), .B1(n5557), .B2(n4743), .C1(n4742), 
        .C2(n5567), .ZN(U2853) );
  OR2_X1 U5886 ( .A1(n4771), .A2(n4873), .ZN(n6405) );
  OAI21_X1 U5887 ( .B1(n6405), .B2(n5044), .A(n6451), .ZN(n4746) );
  NAND2_X1 U5888 ( .A1(n4746), .A2(n6408), .ZN(n4744) );
  OAI21_X1 U5889 ( .B1(n4745), .B2(n6633), .A(n4744), .ZN(n6456) );
  INV_X1 U5890 ( .A(n6456), .ZN(n4767) );
  NOR2_X1 U5891 ( .A1(n4871), .A2(n5825), .ZN(n5829) );
  OR3_X1 U5892 ( .A1(n5829), .A2(n5896), .A3(n4746), .ZN(n4747) );
  OAI211_X1 U5893 ( .C1(n3368), .C2(n6408), .A(n5020), .B(n4747), .ZN(n6457)
         );
  NAND2_X1 U5894 ( .A1(n6457), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4751) );
  INV_X1 U5895 ( .A(n4871), .ZN(n4748) );
  OAI22_X1 U5896 ( .A1(n5084), .A2(n6451), .B1(n6423), .B2(n6450), .ZN(n4749)
         );
  AOI21_X1 U5897 ( .B1(n6420), .B2(n6404), .A(n4749), .ZN(n4750) );
  OAI211_X1 U5898 ( .C1(n4767), .C2(n5918), .A(n4751), .B(n4750), .ZN(U3078)
         );
  NAND2_X1 U5899 ( .A1(n6457), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4754) );
  OAI22_X1 U5900 ( .A1(n5074), .A2(n6451), .B1(n6431), .B2(n6450), .ZN(n4752)
         );
  AOI21_X1 U5901 ( .B1(n6428), .B2(n6404), .A(n4752), .ZN(n4753) );
  OAI211_X1 U5902 ( .C1(n4767), .C2(n5926), .A(n4754), .B(n4753), .ZN(U3080)
         );
  NAND2_X1 U5903 ( .A1(n6457), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4757) );
  OAI22_X1 U5904 ( .A1(n5070), .A2(n6451), .B1(n6441), .B2(n6450), .ZN(n4755)
         );
  AOI21_X1 U5905 ( .B1(n6438), .B2(n6404), .A(n4755), .ZN(n4756) );
  OAI211_X1 U5906 ( .C1(n4767), .C2(n5934), .A(n4757), .B(n4756), .ZN(U3082)
         );
  NAND2_X1 U5907 ( .A1(n6457), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4760) );
  OAI22_X1 U5908 ( .A1(n5066), .A2(n6451), .B1(n6427), .B2(n6450), .ZN(n4758)
         );
  AOI21_X1 U5909 ( .B1(n6424), .B2(n6404), .A(n4758), .ZN(n4759) );
  OAI211_X1 U5910 ( .C1(n4767), .C2(n5922), .A(n4760), .B(n4759), .ZN(U3079)
         );
  NAND2_X1 U5911 ( .A1(n6457), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4763) );
  OAI22_X1 U5912 ( .A1(n5054), .A2(n6451), .B1(n6415), .B2(n6450), .ZN(n4761)
         );
  AOI21_X1 U5913 ( .B1(n6412), .B2(n6404), .A(n4761), .ZN(n4762) );
  OAI211_X1 U5914 ( .C1(n4767), .C2(n5910), .A(n4763), .B(n4762), .ZN(U3076)
         );
  NAND2_X1 U5915 ( .A1(n6457), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4766) );
  OAI22_X1 U5916 ( .A1(n5058), .A2(n6451), .B1(n6449), .B2(n6450), .ZN(n4764)
         );
  AOI21_X1 U5917 ( .B1(n6444), .B2(n6404), .A(n4764), .ZN(n4765) );
  OAI211_X1 U5918 ( .C1(n4767), .C2(n5941), .A(n4766), .B(n4765), .ZN(U3083)
         );
  NOR2_X1 U5919 ( .A1(n4771), .A2(n5896), .ZN(n6395) );
  AND2_X1 U5920 ( .A1(n4772), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6397) );
  INV_X1 U5921 ( .A(n6397), .ZN(n4920) );
  NOR2_X1 U5922 ( .A1(n4920), .A2(n6517), .ZN(n4768) );
  AOI22_X1 U5923 ( .A1(n6395), .A2(n6399), .B1(n6396), .B2(n4768), .ZN(n4805)
         );
  NOR2_X1 U5924 ( .A1(n4769), .A2(n5821), .ZN(n4770) );
  OR2_X1 U5925 ( .A1(n4967), .A2(n5052), .ZN(n4777) );
  AOI21_X1 U5926 ( .B1(n4777), .B2(n4800), .A(n6822), .ZN(n4776) );
  NAND2_X1 U5927 ( .A1(n6408), .A2(n4771), .ZN(n4775) );
  NOR2_X1 U5928 ( .A1(n4772), .A2(n6633), .ZN(n5854) );
  OAI21_X1 U5929 ( .B1(n6396), .B2(n6633), .A(n4867), .ZN(n5189) );
  NOR2_X1 U5930 ( .A1(n5854), .A2(n5189), .ZN(n6410) );
  NAND2_X1 U5931 ( .A1(n6401), .A2(n4773), .ZN(n4801) );
  AOI21_X1 U5932 ( .B1(n4801), .B2(STATE2_REG_3__SCAN_IN), .A(n6517), .ZN(
        n4774) );
  NAND2_X1 U5933 ( .A1(n4799), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4780)
         );
  OAI22_X1 U5934 ( .A1(n5078), .A2(n4801), .B1(n6435), .B2(n4800), .ZN(n4778)
         );
  AOI21_X1 U5935 ( .B1(n6432), .B2(n4998), .A(n4778), .ZN(n4779) );
  OAI211_X1 U5936 ( .C1(n4805), .C2(n5930), .A(n4780), .B(n4779), .ZN(U3137)
         );
  NAND2_X1 U5937 ( .A1(n4799), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4783)
         );
  OAI22_X1 U5938 ( .A1(n5062), .A2(n4801), .B1(n6419), .B2(n4800), .ZN(n4781)
         );
  AOI21_X1 U5939 ( .B1(n6416), .B2(n4998), .A(n4781), .ZN(n4782) );
  OAI211_X1 U5940 ( .C1(n4805), .C2(n5914), .A(n4783), .B(n4782), .ZN(U3133)
         );
  NAND2_X1 U5941 ( .A1(n4799), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4786)
         );
  OAI22_X1 U5942 ( .A1(n5074), .A2(n4801), .B1(n6431), .B2(n4800), .ZN(n4784)
         );
  AOI21_X1 U5943 ( .B1(n6428), .B2(n4998), .A(n4784), .ZN(n4785) );
  OAI211_X1 U5944 ( .C1(n4805), .C2(n5926), .A(n4786), .B(n4785), .ZN(U3136)
         );
  NAND2_X1 U5945 ( .A1(n4799), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4789)
         );
  OAI22_X1 U5946 ( .A1(n5066), .A2(n4801), .B1(n6427), .B2(n4800), .ZN(n4787)
         );
  AOI21_X1 U5947 ( .B1(n6424), .B2(n4998), .A(n4787), .ZN(n4788) );
  OAI211_X1 U5948 ( .C1(n4805), .C2(n5922), .A(n4789), .B(n4788), .ZN(U3135)
         );
  NAND2_X1 U5949 ( .A1(n4799), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4792)
         );
  OAI22_X1 U5950 ( .A1(n5058), .A2(n4801), .B1(n6449), .B2(n4800), .ZN(n4790)
         );
  AOI21_X1 U5951 ( .B1(n6444), .B2(n4998), .A(n4790), .ZN(n4791) );
  OAI211_X1 U5952 ( .C1(n4805), .C2(n5941), .A(n4792), .B(n4791), .ZN(U3139)
         );
  NAND2_X1 U5953 ( .A1(n4799), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4795)
         );
  OAI22_X1 U5954 ( .A1(n5070), .A2(n4801), .B1(n6441), .B2(n4800), .ZN(n4793)
         );
  AOI21_X1 U5955 ( .B1(n6438), .B2(n4998), .A(n4793), .ZN(n4794) );
  OAI211_X1 U5956 ( .C1(n4805), .C2(n5934), .A(n4795), .B(n4794), .ZN(U3138)
         );
  NAND2_X1 U5957 ( .A1(n4799), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4798)
         );
  OAI22_X1 U5958 ( .A1(n5084), .A2(n4801), .B1(n6423), .B2(n4800), .ZN(n4796)
         );
  AOI21_X1 U5959 ( .B1(n6420), .B2(n4998), .A(n4796), .ZN(n4797) );
  OAI211_X1 U5960 ( .C1(n4805), .C2(n5918), .A(n4798), .B(n4797), .ZN(U3134)
         );
  NAND2_X1 U5961 ( .A1(n4799), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4804)
         );
  OAI22_X1 U5962 ( .A1(n5054), .A2(n4801), .B1(n6415), .B2(n4800), .ZN(n4802)
         );
  AOI21_X1 U5963 ( .B1(n6412), .B2(n4998), .A(n4802), .ZN(n4803) );
  OAI211_X1 U5964 ( .C1(n4805), .C2(n5910), .A(n4804), .B(n4803), .ZN(U3132)
         );
  OAI21_X1 U5965 ( .B1(n6494), .B2(n4997), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4809) );
  NAND2_X1 U5966 ( .A1(n4504), .A2(n5823), .ZN(n4874) );
  INV_X1 U5967 ( .A(n4874), .ZN(n4965) );
  AOI21_X1 U5968 ( .B1(n4965), .B2(n4873), .A(n5896), .ZN(n4808) );
  NAND2_X1 U5969 ( .A1(n5018), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4972) );
  NOR2_X1 U5970 ( .A1(n6517), .A2(n4972), .ZN(n4964) );
  AND2_X1 U5971 ( .A1(n6401), .A2(n4964), .ZN(n4831) );
  INV_X1 U5972 ( .A(n5854), .ZN(n5898) );
  OR2_X1 U5973 ( .A1(n6396), .A2(n4865), .ZN(n4924) );
  AOI21_X1 U5974 ( .B1(n4924), .B2(STATE2_REG_2__SCAN_IN), .A(n4806), .ZN(
        n4919) );
  OAI211_X1 U5975 ( .C1(n6623), .C2(n4831), .A(n5898), .B(n4919), .ZN(n4807)
         );
  INV_X1 U5976 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4812) );
  INV_X1 U5977 ( .A(n6419), .ZN(n6462) );
  AOI22_X1 U5978 ( .A1(n4997), .A2(n6462), .B1(n6461), .B2(n4831), .ZN(n4811)
         );
  NAND2_X1 U5979 ( .A1(n4965), .A2(n6408), .ZN(n4879) );
  INV_X1 U5980 ( .A(n6399), .ZN(n5832) );
  OAI22_X1 U5981 ( .A1(n4879), .A2(n5832), .B1(n4920), .B2(n4924), .ZN(n4832)
         );
  AOI22_X1 U5982 ( .A1(n6463), .A2(n4832), .B1(n6494), .B2(n6416), .ZN(n4810)
         );
  OAI211_X1 U5983 ( .C1(n4836), .C2(n4812), .A(n4811), .B(n4810), .ZN(U3117)
         );
  INV_X1 U5984 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4815) );
  INV_X1 U5985 ( .A(n6423), .ZN(n6468) );
  AOI22_X1 U5986 ( .A1(n4997), .A2(n6468), .B1(n6467), .B2(n4831), .ZN(n4814)
         );
  AOI22_X1 U5987 ( .A1(n6469), .A2(n4832), .B1(n6494), .B2(n6420), .ZN(n4813)
         );
  OAI211_X1 U5988 ( .C1(n4836), .C2(n4815), .A(n4814), .B(n4813), .ZN(U3118)
         );
  INV_X1 U5989 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4818) );
  AOI22_X1 U5990 ( .A1(n4997), .A2(n5881), .B1(n6436), .B2(n4831), .ZN(n4817)
         );
  AOI22_X1 U5991 ( .A1(n6437), .A2(n4832), .B1(n6494), .B2(n6438), .ZN(n4816)
         );
  OAI211_X1 U5992 ( .C1(n4836), .C2(n4818), .A(n4817), .B(n4816), .ZN(U3122)
         );
  INV_X1 U5993 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4821) );
  AOI22_X1 U5994 ( .A1(n4997), .A2(n5851), .B1(n6402), .B2(n4831), .ZN(n4820)
         );
  AOI22_X1 U5995 ( .A1(n6403), .A2(n4832), .B1(n6494), .B2(n6412), .ZN(n4819)
         );
  OAI211_X1 U5996 ( .C1(n4836), .C2(n4821), .A(n4820), .B(n4819), .ZN(U3116)
         );
  INV_X1 U5997 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4824) );
  INV_X1 U5998 ( .A(n6435), .ZN(n6486) );
  AOI22_X1 U5999 ( .A1(n4997), .A2(n6486), .B1(n6485), .B2(n4831), .ZN(n4823)
         );
  AOI22_X1 U6000 ( .A1(n6487), .A2(n4832), .B1(n6494), .B2(n6432), .ZN(n4822)
         );
  OAI211_X1 U6001 ( .C1(n4836), .C2(n4824), .A(n4823), .B(n4822), .ZN(U3121)
         );
  INV_X1 U6002 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4827) );
  INV_X1 U6003 ( .A(n6427), .ZN(n6474) );
  AOI22_X1 U6004 ( .A1(n4997), .A2(n6474), .B1(n6473), .B2(n4831), .ZN(n4826)
         );
  AOI22_X1 U6005 ( .A1(n6475), .A2(n4832), .B1(n6494), .B2(n6424), .ZN(n4825)
         );
  OAI211_X1 U6006 ( .C1(n4836), .C2(n4827), .A(n4826), .B(n4825), .ZN(U3119)
         );
  INV_X1 U6007 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4830) );
  INV_X1 U6008 ( .A(n6449), .ZN(n6493) );
  AOI22_X1 U6009 ( .A1(n4997), .A2(n6493), .B1(n6492), .B2(n4831), .ZN(n4829)
         );
  AOI22_X1 U6010 ( .A1(n6496), .A2(n4832), .B1(n6494), .B2(n6444), .ZN(n4828)
         );
  OAI211_X1 U6011 ( .C1(n4836), .C2(n4830), .A(n4829), .B(n4828), .ZN(U3123)
         );
  INV_X1 U6012 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4835) );
  INV_X1 U6013 ( .A(n6431), .ZN(n6480) );
  AOI22_X1 U6014 ( .A1(n4997), .A2(n6480), .B1(n6479), .B2(n4831), .ZN(n4834)
         );
  AOI22_X1 U6015 ( .A1(n6481), .A2(n4832), .B1(n6494), .B2(n6428), .ZN(n4833)
         );
  OAI211_X1 U6016 ( .C1(n4836), .C2(n4835), .A(n4834), .B(n4833), .ZN(U3120)
         );
  INV_X1 U6017 ( .A(n4845), .ZN(n4837) );
  OR2_X1 U6018 ( .A1(n5821), .A2(n6822), .ZN(n4838) );
  OR2_X1 U6019 ( .A1(n5105), .A2(n4838), .ZN(n4839) );
  INV_X1 U6020 ( .A(n4840), .ZN(n4966) );
  OR2_X1 U6021 ( .A1(n4504), .A2(n4427), .ZN(n5017) );
  INV_X1 U6022 ( .A(n5017), .ZN(n4916) );
  NAND3_X1 U6023 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6512), .A3(n5018), .ZN(n4918) );
  NOR2_X1 U6024 ( .A1(n6401), .A2(n4918), .ZN(n4862) );
  AOI21_X1 U6025 ( .B1(n4966), .B2(n4916), .A(n4862), .ZN(n4844) );
  AOI22_X1 U6026 ( .A1(n4842), .A2(n4844), .B1(n5896), .B2(n4918), .ZN(n4841)
         );
  NAND2_X1 U6027 ( .A1(n5020), .A2(n4841), .ZN(n4861) );
  INV_X1 U6028 ( .A(n4842), .ZN(n4843) );
  OAI22_X1 U6029 ( .A1(n4844), .A2(n4843), .B1(n6633), .B2(n4918), .ZN(n4860)
         );
  AOI22_X1 U6030 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4861), .B1(n6475), 
        .B2(n4860), .ZN(n4847) );
  AOI22_X1 U6031 ( .A1(n5939), .A2(n6474), .B1(n4862), .B2(n6473), .ZN(n4846)
         );
  OAI211_X1 U6032 ( .C1(n6478), .C2(n4963), .A(n4847), .B(n4846), .ZN(U3095)
         );
  AOI22_X1 U6033 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4861), .B1(n6487), 
        .B2(n4860), .ZN(n4849) );
  AOI22_X1 U6034 ( .A1(n5939), .A2(n6486), .B1(n4862), .B2(n6485), .ZN(n4848)
         );
  OAI211_X1 U6035 ( .C1(n6490), .C2(n4963), .A(n4849), .B(n4848), .ZN(U3097)
         );
  AOI22_X1 U6036 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4861), .B1(n6469), 
        .B2(n4860), .ZN(n4851) );
  AOI22_X1 U6037 ( .A1(n5939), .A2(n6468), .B1(n4862), .B2(n6467), .ZN(n4850)
         );
  OAI211_X1 U6038 ( .C1(n6472), .C2(n4963), .A(n4851), .B(n4850), .ZN(U3094)
         );
  AOI22_X1 U6039 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4861), .B1(n6496), 
        .B2(n4860), .ZN(n4853) );
  AOI22_X1 U6040 ( .A1(n5939), .A2(n6493), .B1(n4862), .B2(n6492), .ZN(n4852)
         );
  OAI211_X1 U6041 ( .C1(n6501), .C2(n4963), .A(n4853), .B(n4852), .ZN(U3099)
         );
  AOI22_X1 U6042 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4861), .B1(n6481), 
        .B2(n4860), .ZN(n4855) );
  AOI22_X1 U6043 ( .A1(n5939), .A2(n6480), .B1(n4862), .B2(n6479), .ZN(n4854)
         );
  OAI211_X1 U6044 ( .C1(n6484), .C2(n4963), .A(n4855), .B(n4854), .ZN(U3096)
         );
  AOI22_X1 U6045 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4861), .B1(n6437), 
        .B2(n4860), .ZN(n4857) );
  AOI22_X1 U6046 ( .A1(n5939), .A2(n5881), .B1(n4862), .B2(n6436), .ZN(n4856)
         );
  OAI211_X1 U6047 ( .C1(n5132), .C2(n4963), .A(n4857), .B(n4856), .ZN(U3098)
         );
  AOI22_X1 U6048 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4861), .B1(n6463), 
        .B2(n4860), .ZN(n4859) );
  AOI22_X1 U6049 ( .A1(n5939), .A2(n6462), .B1(n4862), .B2(n6461), .ZN(n4858)
         );
  OAI211_X1 U6050 ( .C1(n6466), .C2(n4963), .A(n4859), .B(n4858), .ZN(U3093)
         );
  AOI22_X1 U6051 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4861), .B1(n6403), 
        .B2(n4860), .ZN(n4864) );
  AOI22_X1 U6052 ( .A1(n5939), .A2(n5851), .B1(n6402), .B2(n4862), .ZN(n4863)
         );
  OAI211_X1 U6053 ( .C1(n5123), .C2(n4963), .A(n4864), .B(n4863), .ZN(U3092)
         );
  OR2_X1 U6054 ( .A1(n4972), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5048)
         );
  NOR2_X1 U6055 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5048), .ZN(n4901)
         );
  INV_X1 U6056 ( .A(n4901), .ZN(n4868) );
  INV_X1 U6057 ( .A(n4865), .ZN(n4866) );
  OR2_X1 U6058 ( .A1(n6396), .A2(n4866), .ZN(n4878) );
  INV_X1 U6059 ( .A(n4878), .ZN(n5853) );
  OAI21_X1 U6060 ( .B1(n5853), .B2(n6633), .A(n4867), .ZN(n5847) );
  AOI211_X1 U6061 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4868), .A(n5854), .B(
        n5847), .ZN(n4876) );
  INV_X1 U6062 ( .A(n4638), .ZN(n5835) );
  INV_X1 U6063 ( .A(n4869), .ZN(n4870) );
  NAND3_X1 U6064 ( .A1(n5835), .A2(n4870), .A3(n5826), .ZN(n4877) );
  INV_X1 U6065 ( .A(n5053), .ZN(n4872) );
  OR2_X1 U6066 ( .A1(n4874), .A2(n4873), .ZN(n5045) );
  OAI211_X1 U6067 ( .C1(n5844), .C2(n4877), .A(n5047), .B(n5045), .ZN(n4875)
         );
  INV_X1 U6068 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4882) );
  AOI22_X1 U6069 ( .A1(n5149), .A2(n6412), .B1(n6402), .B2(n4901), .ZN(n4881)
         );
  OAI22_X1 U6070 ( .A1(n4879), .A2(n6399), .B1(n4878), .B2(n4920), .ZN(n4902)
         );
  NOR2_X2 U6071 ( .A1(n5053), .A2(n5016), .ZN(n5087) );
  AOI22_X1 U6072 ( .A1(n6403), .A2(n4902), .B1(n5087), .B2(n5851), .ZN(n4880)
         );
  OAI211_X1 U6073 ( .C1(n4906), .C2(n4882), .A(n4881), .B(n4880), .ZN(U3052)
         );
  INV_X1 U6074 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4885) );
  AOI22_X1 U6075 ( .A1(n5149), .A2(n6416), .B1(n6461), .B2(n4901), .ZN(n4884)
         );
  AOI22_X1 U6076 ( .A1(n6463), .A2(n4902), .B1(n5087), .B2(n6462), .ZN(n4883)
         );
  OAI211_X1 U6077 ( .C1(n4906), .C2(n4885), .A(n4884), .B(n4883), .ZN(U3053)
         );
  INV_X1 U6078 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4888) );
  AOI22_X1 U6079 ( .A1(n5149), .A2(n6420), .B1(n6467), .B2(n4901), .ZN(n4887)
         );
  AOI22_X1 U6080 ( .A1(n6469), .A2(n4902), .B1(n5087), .B2(n6468), .ZN(n4886)
         );
  OAI211_X1 U6081 ( .C1(n4906), .C2(n4888), .A(n4887), .B(n4886), .ZN(U3054)
         );
  INV_X1 U6082 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4891) );
  AOI22_X1 U6083 ( .A1(n5149), .A2(n6424), .B1(n6473), .B2(n4901), .ZN(n4890)
         );
  AOI22_X1 U6084 ( .A1(n6475), .A2(n4902), .B1(n5087), .B2(n6474), .ZN(n4889)
         );
  OAI211_X1 U6085 ( .C1(n4906), .C2(n4891), .A(n4890), .B(n4889), .ZN(U3055)
         );
  INV_X1 U6086 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4894) );
  AOI22_X1 U6087 ( .A1(n5149), .A2(n6428), .B1(n6479), .B2(n4901), .ZN(n4893)
         );
  AOI22_X1 U6088 ( .A1(n6481), .A2(n4902), .B1(n5087), .B2(n6480), .ZN(n4892)
         );
  OAI211_X1 U6089 ( .C1(n4906), .C2(n4894), .A(n4893), .B(n4892), .ZN(U3056)
         );
  INV_X1 U6090 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4897) );
  AOI22_X1 U6091 ( .A1(n5149), .A2(n6432), .B1(n6485), .B2(n4901), .ZN(n4896)
         );
  AOI22_X1 U6092 ( .A1(n6487), .A2(n4902), .B1(n5087), .B2(n6486), .ZN(n4895)
         );
  OAI211_X1 U6093 ( .C1(n4906), .C2(n4897), .A(n4896), .B(n4895), .ZN(U3057)
         );
  INV_X1 U6094 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4900) );
  AOI22_X1 U6095 ( .A1(n5149), .A2(n6438), .B1(n6436), .B2(n4901), .ZN(n4899)
         );
  AOI22_X1 U6096 ( .A1(n6437), .A2(n4902), .B1(n5087), .B2(n5881), .ZN(n4898)
         );
  OAI211_X1 U6097 ( .C1(n4906), .C2(n4900), .A(n4899), .B(n4898), .ZN(U3058)
         );
  INV_X1 U6098 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4905) );
  AOI22_X1 U6099 ( .A1(n5149), .A2(n6444), .B1(n6492), .B2(n4901), .ZN(n4904)
         );
  AOI22_X1 U6100 ( .A1(n6496), .A2(n4902), .B1(n5087), .B2(n6493), .ZN(n4903)
         );
  OAI211_X1 U6101 ( .C1(n4906), .C2(n4905), .A(n4904), .B(n4903), .ZN(U3059)
         );
  XNOR2_X1 U6102 ( .A(n4908), .B(n4907), .ZN(n5096) );
  INV_X1 U6103 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6578) );
  NOR2_X1 U6104 ( .A1(n6338), .A2(n6578), .ZN(n5091) );
  NOR2_X1 U6105 ( .A1(n4910), .A2(n4909), .ZN(n4913) );
  INV_X1 U6106 ( .A(n4911), .ZN(n4912) );
  MUX2_X1 U6107 ( .A(n4913), .B(n4912), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4914) );
  AOI211_X1 U6108 ( .C1(n6382), .C2(n6171), .A(n5091), .B(n4914), .ZN(n4915)
         );
  OAI21_X1 U6109 ( .B1(n6035), .B2(n5096), .A(n4915), .ZN(U3012) );
  NAND3_X1 U6110 ( .A1(n4963), .A2(n6408), .A3(n6450), .ZN(n4917) );
  AND2_X1 U6111 ( .A1(n4916), .A2(n6399), .ZN(n4923) );
  AOI21_X1 U6112 ( .B1(n4917), .B2(n5834), .A(n4923), .ZN(n4922) );
  NOR2_X1 U6113 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4918), .ZN(n4957)
         );
  OAI211_X1 U6114 ( .C1(n6623), .C2(n4957), .A(n4920), .B(n4919), .ZN(n4921)
         );
  NAND2_X1 U6115 ( .A1(n4956), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4931) );
  NAND2_X1 U6116 ( .A1(n4923), .A2(n6408), .ZN(n4927) );
  INV_X1 U6117 ( .A(n4924), .ZN(n4925) );
  NAND2_X1 U6118 ( .A1(n5854), .A2(n4925), .ZN(n4926) );
  NAND2_X1 U6119 ( .A1(n4927), .A2(n4926), .ZN(n4960) );
  NAND2_X1 U6120 ( .A1(n6467), .A2(n4957), .ZN(n4928) );
  OAI21_X1 U6121 ( .B1(n6450), .B2(n6472), .A(n4928), .ZN(n4929) );
  AOI21_X1 U6122 ( .B1(n6469), .B2(n4960), .A(n4929), .ZN(n4930) );
  OAI211_X1 U6123 ( .C1(n6423), .C2(n4963), .A(n4931), .B(n4930), .ZN(U3086)
         );
  NAND2_X1 U6124 ( .A1(n4956), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4935) );
  NAND2_X1 U6125 ( .A1(n6473), .A2(n4957), .ZN(n4932) );
  OAI21_X1 U6126 ( .B1(n6450), .B2(n6478), .A(n4932), .ZN(n4933) );
  AOI21_X1 U6127 ( .B1(n6475), .B2(n4960), .A(n4933), .ZN(n4934) );
  OAI211_X1 U6128 ( .C1(n6427), .C2(n4963), .A(n4935), .B(n4934), .ZN(U3087)
         );
  NAND2_X1 U6129 ( .A1(n4956), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4939) );
  NAND2_X1 U6130 ( .A1(n6479), .A2(n4957), .ZN(n4936) );
  OAI21_X1 U6131 ( .B1(n6450), .B2(n6484), .A(n4936), .ZN(n4937) );
  AOI21_X1 U6132 ( .B1(n6481), .B2(n4960), .A(n4937), .ZN(n4938) );
  OAI211_X1 U6133 ( .C1(n6431), .C2(n4963), .A(n4939), .B(n4938), .ZN(U3088)
         );
  NAND2_X1 U6134 ( .A1(n4956), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4943) );
  NAND2_X1 U6135 ( .A1(n6485), .A2(n4957), .ZN(n4940) );
  OAI21_X1 U6136 ( .B1(n6450), .B2(n6490), .A(n4940), .ZN(n4941) );
  AOI21_X1 U6137 ( .B1(n6487), .B2(n4960), .A(n4941), .ZN(n4942) );
  OAI211_X1 U6138 ( .C1(n6435), .C2(n4963), .A(n4943), .B(n4942), .ZN(U3089)
         );
  NAND2_X1 U6139 ( .A1(n4956), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4947) );
  NAND2_X1 U6140 ( .A1(n6436), .A2(n4957), .ZN(n4944) );
  OAI21_X1 U6141 ( .B1(n6450), .B2(n5132), .A(n4944), .ZN(n4945) );
  AOI21_X1 U6142 ( .B1(n6437), .B2(n4960), .A(n4945), .ZN(n4946) );
  OAI211_X1 U6143 ( .C1(n6441), .C2(n4963), .A(n4947), .B(n4946), .ZN(U3090)
         );
  NAND2_X1 U6144 ( .A1(n4956), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4951) );
  NAND2_X1 U6145 ( .A1(n6402), .A2(n4957), .ZN(n4948) );
  OAI21_X1 U6146 ( .B1(n6450), .B2(n5123), .A(n4948), .ZN(n4949) );
  AOI21_X1 U6147 ( .B1(n6403), .B2(n4960), .A(n4949), .ZN(n4950) );
  OAI211_X1 U6148 ( .C1(n6415), .C2(n4963), .A(n4951), .B(n4950), .ZN(U3084)
         );
  NAND2_X1 U6149 ( .A1(n4956), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4955) );
  NAND2_X1 U6150 ( .A1(n6492), .A2(n4957), .ZN(n4952) );
  OAI21_X1 U6151 ( .B1(n6450), .B2(n6501), .A(n4952), .ZN(n4953) );
  AOI21_X1 U6152 ( .B1(n6496), .B2(n4960), .A(n4953), .ZN(n4954) );
  OAI211_X1 U6153 ( .C1(n6449), .C2(n4963), .A(n4955), .B(n4954), .ZN(U3091)
         );
  NAND2_X1 U6154 ( .A1(n4956), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4962) );
  NAND2_X1 U6155 ( .A1(n6461), .A2(n4957), .ZN(n4958) );
  OAI21_X1 U6156 ( .B1(n6450), .B2(n6466), .A(n4958), .ZN(n4959) );
  AOI21_X1 U6157 ( .B1(n6463), .B2(n4960), .A(n4959), .ZN(n4961) );
  OAI211_X1 U6158 ( .C1(n6419), .C2(n4963), .A(n4962), .B(n4961), .ZN(U3085)
         );
  INV_X1 U6159 ( .A(n4964), .ZN(n4971) );
  AND2_X1 U6160 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4964), .ZN(n4996)
         );
  AOI21_X1 U6161 ( .B1(n4966), .B2(n4965), .A(n4996), .ZN(n4974) );
  INV_X1 U6162 ( .A(n4967), .ZN(n4968) );
  NAND2_X1 U6163 ( .A1(n4968), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5106) );
  NAND2_X1 U6164 ( .A1(n4974), .A2(n5106), .ZN(n4969) );
  NOR2_X1 U6165 ( .A1(n5896), .A2(n4969), .ZN(n4970) );
  AOI211_X2 U6166 ( .C1(n5896), .C2(n4971), .A(n4970), .B(n5112), .ZN(n5003)
         );
  INV_X1 U6167 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4977) );
  AOI22_X1 U6168 ( .A1(n4997), .A2(n6444), .B1(n6492), .B2(n4996), .ZN(n4976)
         );
  NAND2_X1 U6169 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4973) );
  OAI22_X1 U6170 ( .A1(n4974), .A2(n5896), .B1(n4973), .B2(n4972), .ZN(n4999)
         );
  AOI22_X1 U6171 ( .A1(n6496), .A2(n4999), .B1(n6493), .B2(n4998), .ZN(n4975)
         );
  OAI211_X1 U6172 ( .C1(n5003), .C2(n4977), .A(n4976), .B(n4975), .ZN(U3131)
         );
  INV_X1 U6173 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4980) );
  AOI22_X1 U6174 ( .A1(n4997), .A2(n6432), .B1(n6485), .B2(n4996), .ZN(n4979)
         );
  AOI22_X1 U6175 ( .A1(n6487), .A2(n4999), .B1(n6486), .B2(n4998), .ZN(n4978)
         );
  OAI211_X1 U6176 ( .C1(n5003), .C2(n4980), .A(n4979), .B(n4978), .ZN(U3129)
         );
  INV_X1 U6177 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4983) );
  AOI22_X1 U6178 ( .A1(n4997), .A2(n6412), .B1(n6402), .B2(n4996), .ZN(n4982)
         );
  AOI22_X1 U6179 ( .A1(n6403), .A2(n4999), .B1(n5851), .B2(n4998), .ZN(n4981)
         );
  OAI211_X1 U6180 ( .C1(n5003), .C2(n4983), .A(n4982), .B(n4981), .ZN(U3124)
         );
  INV_X1 U6181 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4986) );
  AOI22_X1 U6182 ( .A1(n4997), .A2(n6416), .B1(n6461), .B2(n4996), .ZN(n4985)
         );
  AOI22_X1 U6183 ( .A1(n6463), .A2(n4999), .B1(n6462), .B2(n4998), .ZN(n4984)
         );
  OAI211_X1 U6184 ( .C1(n5003), .C2(n4986), .A(n4985), .B(n4984), .ZN(U3125)
         );
  INV_X1 U6185 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4989) );
  AOI22_X1 U6186 ( .A1(n4997), .A2(n6420), .B1(n6467), .B2(n4996), .ZN(n4988)
         );
  AOI22_X1 U6187 ( .A1(n6469), .A2(n4999), .B1(n6468), .B2(n4998), .ZN(n4987)
         );
  OAI211_X1 U6188 ( .C1(n5003), .C2(n4989), .A(n4988), .B(n4987), .ZN(U3126)
         );
  INV_X1 U6189 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4992) );
  AOI22_X1 U6190 ( .A1(n4997), .A2(n6438), .B1(n6436), .B2(n4996), .ZN(n4991)
         );
  AOI22_X1 U6191 ( .A1(n6437), .A2(n4999), .B1(n5881), .B2(n4998), .ZN(n4990)
         );
  OAI211_X1 U6192 ( .C1(n5003), .C2(n4992), .A(n4991), .B(n4990), .ZN(U3130)
         );
  INV_X1 U6193 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4995) );
  AOI22_X1 U6194 ( .A1(n4997), .A2(n6428), .B1(n6479), .B2(n4996), .ZN(n4994)
         );
  AOI22_X1 U6195 ( .A1(n6481), .A2(n4999), .B1(n6480), .B2(n4998), .ZN(n4993)
         );
  OAI211_X1 U6196 ( .C1(n5003), .C2(n4995), .A(n4994), .B(n4993), .ZN(U3128)
         );
  INV_X1 U6197 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n5002) );
  AOI22_X1 U6198 ( .A1(n4997), .A2(n6424), .B1(n6473), .B2(n4996), .ZN(n5001)
         );
  AOI22_X1 U6199 ( .A1(n6475), .A2(n4999), .B1(n6474), .B2(n4998), .ZN(n5000)
         );
  OAI211_X1 U6200 ( .C1(n5003), .C2(n5002), .A(n5001), .B(n5000), .ZN(U3127)
         );
  AOI21_X1 U6201 ( .B1(n5004), .B2(n5007), .A(n5006), .ZN(n6301) );
  AND2_X1 U6202 ( .A1(n5009), .A2(n5008), .ZN(n5010) );
  OR2_X1 U6203 ( .A1(n5010), .A2(n3021), .ZN(n6162) );
  INV_X1 U6204 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5011) );
  OAI22_X1 U6205 ( .A1(n6162), .A2(n5557), .B1(n5011), .B2(n5567), .ZN(n5012)
         );
  AOI21_X1 U6206 ( .B1(n6301), .B2(n4283), .A(n5012), .ZN(n5013) );
  INV_X1 U6207 ( .A(n5013), .ZN(U2852) );
  INV_X1 U6208 ( .A(n6301), .ZN(n6157) );
  AOI22_X1 U6209 ( .A1(n5583), .A2(DATAI_7_), .B1(n6250), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n5014) );
  OAI21_X1 U6210 ( .B1(n6157), .B2(n5988), .A(n5014), .ZN(U2884) );
  NOR2_X1 U6211 ( .A1(n6399), .A2(n5017), .ZN(n5852) );
  NAND3_X1 U6212 ( .A1(n6517), .A2(n6512), .A3(n5018), .ZN(n5846) );
  NOR2_X1 U6213 ( .A1(n6401), .A2(n5846), .ZN(n5041) );
  AOI21_X1 U6214 ( .B1(n5852), .B2(n3358), .A(n5041), .ZN(n5023) );
  AOI21_X1 U6215 ( .B1(n5024), .B2(STATEBS16_REG_SCAN_IN), .A(n5896), .ZN(
        n5021) );
  AOI22_X1 U6216 ( .A1(n5023), .A2(n5021), .B1(n5896), .B2(n5846), .ZN(n5019)
         );
  NAND2_X1 U6217 ( .A1(n5020), .A2(n5019), .ZN(n5040) );
  INV_X1 U6218 ( .A(n5021), .ZN(n5022) );
  OAI22_X1 U6219 ( .A1(n5023), .A2(n5022), .B1(n6633), .B2(n5846), .ZN(n5039)
         );
  AOI22_X1 U6220 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5040), .B1(n6496), 
        .B2(n5039), .ZN(n5026) );
  AOI22_X1 U6221 ( .A1(n5889), .A2(n6444), .B1(n6492), .B2(n5041), .ZN(n5025)
         );
  OAI211_X1 U6222 ( .C1(n6449), .C2(n5194), .A(n5026), .B(n5025), .ZN(U3035)
         );
  AOI22_X1 U6223 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5040), .B1(n6463), 
        .B2(n5039), .ZN(n5028) );
  AOI22_X1 U6224 ( .A1(n5889), .A2(n6416), .B1(n6461), .B2(n5041), .ZN(n5027)
         );
  OAI211_X1 U6225 ( .C1(n6419), .C2(n5194), .A(n5028), .B(n5027), .ZN(U3029)
         );
  AOI22_X1 U6226 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5040), .B1(n6403), 
        .B2(n5039), .ZN(n5030) );
  AOI22_X1 U6227 ( .A1(n5889), .A2(n6412), .B1(n6402), .B2(n5041), .ZN(n5029)
         );
  OAI211_X1 U6228 ( .C1(n6415), .C2(n5194), .A(n5030), .B(n5029), .ZN(U3028)
         );
  AOI22_X1 U6229 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5040), .B1(n6469), 
        .B2(n5039), .ZN(n5032) );
  AOI22_X1 U6230 ( .A1(n5889), .A2(n6420), .B1(n6467), .B2(n5041), .ZN(n5031)
         );
  OAI211_X1 U6231 ( .C1(n6423), .C2(n5194), .A(n5032), .B(n5031), .ZN(U3030)
         );
  AOI22_X1 U6232 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5040), .B1(n6475), 
        .B2(n5039), .ZN(n5034) );
  AOI22_X1 U6233 ( .A1(n5889), .A2(n6424), .B1(n6473), .B2(n5041), .ZN(n5033)
         );
  OAI211_X1 U6234 ( .C1(n6427), .C2(n5194), .A(n5034), .B(n5033), .ZN(U3031)
         );
  AOI22_X1 U6235 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5040), .B1(n6437), 
        .B2(n5039), .ZN(n5036) );
  AOI22_X1 U6236 ( .A1(n5889), .A2(n6438), .B1(n6436), .B2(n5041), .ZN(n5035)
         );
  OAI211_X1 U6237 ( .C1(n6441), .C2(n5194), .A(n5036), .B(n5035), .ZN(U3034)
         );
  AOI22_X1 U6238 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5040), .B1(n6481), 
        .B2(n5039), .ZN(n5038) );
  AOI22_X1 U6239 ( .A1(n5889), .A2(n6428), .B1(n6479), .B2(n5041), .ZN(n5037)
         );
  OAI211_X1 U6240 ( .C1(n6431), .C2(n5194), .A(n5038), .B(n5037), .ZN(U3032)
         );
  AOI22_X1 U6241 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5040), .B1(n6487), 
        .B2(n5039), .ZN(n5043) );
  AOI22_X1 U6242 ( .A1(n5889), .A2(n6432), .B1(n6485), .B2(n5041), .ZN(n5042)
         );
  OAI211_X1 U6243 ( .C1(n6435), .C2(n5194), .A(n5043), .B(n5042), .ZN(U3033)
         );
  OR2_X1 U6244 ( .A1(n6401), .A2(n5048), .ZN(n5083) );
  OAI21_X1 U6245 ( .B1(n5045), .B2(n5044), .A(n5083), .ZN(n5050) );
  INV_X1 U6246 ( .A(n5048), .ZN(n5046) );
  AOI22_X1 U6247 ( .A1(n5047), .A2(n5050), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5046), .ZN(n5090) );
  INV_X1 U6248 ( .A(n5047), .ZN(n5051) );
  AOI21_X1 U6249 ( .B1(n5896), .B2(n5048), .A(n5112), .ZN(n5049) );
  NAND2_X1 U6250 ( .A1(n5082), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n5057) );
  INV_X1 U6251 ( .A(n6445), .ZN(n5085) );
  OAI22_X1 U6252 ( .A1(n5085), .A2(n6415), .B1(n5054), .B2(n5083), .ZN(n5055)
         );
  AOI21_X1 U6253 ( .B1(n6412), .B2(n5087), .A(n5055), .ZN(n5056) );
  OAI211_X1 U6254 ( .C1(n5090), .C2(n5910), .A(n5057), .B(n5056), .ZN(U3060)
         );
  NAND2_X1 U6255 ( .A1(n5082), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5061) );
  OAI22_X1 U6256 ( .A1(n5085), .A2(n6449), .B1(n5058), .B2(n5083), .ZN(n5059)
         );
  AOI21_X1 U6257 ( .B1(n6444), .B2(n5087), .A(n5059), .ZN(n5060) );
  OAI211_X1 U6258 ( .C1(n5090), .C2(n5941), .A(n5061), .B(n5060), .ZN(U3067)
         );
  NAND2_X1 U6259 ( .A1(n5082), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n5065) );
  OAI22_X1 U6260 ( .A1(n5085), .A2(n6419), .B1(n5062), .B2(n5083), .ZN(n5063)
         );
  AOI21_X1 U6261 ( .B1(n6416), .B2(n5087), .A(n5063), .ZN(n5064) );
  OAI211_X1 U6262 ( .C1(n5090), .C2(n5914), .A(n5065), .B(n5064), .ZN(U3061)
         );
  NAND2_X1 U6263 ( .A1(n5082), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5069) );
  OAI22_X1 U6264 ( .A1(n5085), .A2(n6427), .B1(n5066), .B2(n5083), .ZN(n5067)
         );
  AOI21_X1 U6265 ( .B1(n6424), .B2(n5087), .A(n5067), .ZN(n5068) );
  OAI211_X1 U6266 ( .C1(n5090), .C2(n5922), .A(n5069), .B(n5068), .ZN(U3063)
         );
  NAND2_X1 U6267 ( .A1(n5082), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5073) );
  OAI22_X1 U6268 ( .A1(n5085), .A2(n6441), .B1(n5070), .B2(n5083), .ZN(n5071)
         );
  AOI21_X1 U6269 ( .B1(n6438), .B2(n5087), .A(n5071), .ZN(n5072) );
  OAI211_X1 U6270 ( .C1(n5090), .C2(n5934), .A(n5073), .B(n5072), .ZN(U3066)
         );
  NAND2_X1 U6271 ( .A1(n5082), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5077) );
  OAI22_X1 U6272 ( .A1(n5085), .A2(n6431), .B1(n5074), .B2(n5083), .ZN(n5075)
         );
  AOI21_X1 U6273 ( .B1(n6428), .B2(n5087), .A(n5075), .ZN(n5076) );
  OAI211_X1 U6274 ( .C1(n5090), .C2(n5926), .A(n5077), .B(n5076), .ZN(U3064)
         );
  NAND2_X1 U6275 ( .A1(n5082), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n5081) );
  OAI22_X1 U6276 ( .A1(n5085), .A2(n6435), .B1(n5078), .B2(n5083), .ZN(n5079)
         );
  AOI21_X1 U6277 ( .B1(n6432), .B2(n5087), .A(n5079), .ZN(n5080) );
  OAI211_X1 U6278 ( .C1(n5090), .C2(n5930), .A(n5081), .B(n5080), .ZN(U3065)
         );
  NAND2_X1 U6279 ( .A1(n5082), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5089) );
  OAI22_X1 U6280 ( .A1(n5085), .A2(n6423), .B1(n5084), .B2(n5083), .ZN(n5086)
         );
  AOI21_X1 U6281 ( .B1(n6420), .B2(n5087), .A(n5086), .ZN(n5088) );
  OAI211_X1 U6282 ( .C1(n5090), .C2(n5918), .A(n5089), .B(n5088), .ZN(U3062)
         );
  INV_X1 U6283 ( .A(n5091), .ZN(n5092) );
  OAI21_X1 U6284 ( .B1(n6314), .B2(n6164), .A(n5092), .ZN(n5094) );
  NOR2_X1 U6285 ( .A1(n6168), .A2(n6335), .ZN(n5093) );
  AOI211_X1 U6286 ( .C1(n6310), .C2(n6165), .A(n5094), .B(n5093), .ZN(n5095)
         );
  OAI21_X1 U6287 ( .B1(n6297), .B2(n5096), .A(n5095), .ZN(U2980) );
  NAND2_X1 U6288 ( .A1(n4112), .A2(n5097), .ZN(n5098) );
  NAND2_X1 U6289 ( .A1(n6167), .A2(n5098), .ZN(n6209) );
  OR2_X1 U6290 ( .A1(n5100), .A2(n5099), .ZN(n6202) );
  INV_X1 U6291 ( .A(n6202), .ZN(n6219) );
  OAI22_X1 U6292 ( .A1(n6216), .A2(n4412), .B1(n6380), .B2(n6200), .ZN(n5102)
         );
  INV_X1 U6293 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6392) );
  NOR2_X1 U6294 ( .A1(n5288), .A2(n6392), .ZN(n5101) );
  AOI211_X1 U6295 ( .C1(n6219), .C2(n3358), .A(n5102), .B(n5101), .ZN(n5104)
         );
  OAI21_X1 U6296 ( .B1(n6218), .B2(n6225), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5103) );
  OAI211_X1 U6297 ( .C1(n6227), .C2(n6336), .A(n5104), .B(n5103), .ZN(U2827)
         );
  NAND2_X1 U6298 ( .A1(n5106), .A2(n5105), .ZN(n5830) );
  NOR3_X1 U6299 ( .A1(n5830), .A2(n5107), .A3(n5825), .ZN(n5108) );
  NOR2_X1 U6300 ( .A1(n5108), .A2(n5896), .ZN(n5114) );
  NOR2_X1 U6301 ( .A1(n6399), .A2(n5109), .ZN(n5195) );
  NOR2_X1 U6302 ( .A1(n5110), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5148)
         );
  AOI21_X1 U6303 ( .B1(n5195), .B2(n3358), .A(n5148), .ZN(n5115) );
  NAND3_X1 U6304 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6517), .A3(n6512), .ZN(n5187) );
  INV_X1 U6305 ( .A(n5187), .ZN(n5111) );
  NOR2_X1 U6306 ( .A1(n6408), .A2(n5111), .ZN(n5113) );
  INV_X1 U6307 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5121) );
  INV_X1 U6308 ( .A(n5114), .ZN(n5116) );
  OAI22_X1 U6309 ( .A1(n5116), .A2(n5115), .B1(n5187), .B2(n6633), .ZN(n5152)
         );
  NAND3_X1 U6310 ( .A1(n5835), .A2(n5117), .A3(n5826), .ZN(n5193) );
  AOI22_X1 U6311 ( .A1(n5149), .A2(n6493), .B1(n6492), .B2(n5148), .ZN(n5118)
         );
  OAI21_X1 U6312 ( .B1(n6501), .B2(n5193), .A(n5118), .ZN(n5119) );
  AOI21_X1 U6313 ( .B1(n5152), .B2(n6496), .A(n5119), .ZN(n5120) );
  OAI21_X1 U6314 ( .B1(n5155), .B2(n5121), .A(n5120), .ZN(U3051) );
  INV_X1 U6315 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n5126) );
  AOI22_X1 U6316 ( .A1(n5149), .A2(n5851), .B1(n6402), .B2(n5148), .ZN(n5122)
         );
  OAI21_X1 U6317 ( .B1(n5123), .B2(n5193), .A(n5122), .ZN(n5124) );
  AOI21_X1 U6318 ( .B1(n5152), .B2(n6403), .A(n5124), .ZN(n5125) );
  OAI21_X1 U6319 ( .B1(n5155), .B2(n5126), .A(n5125), .ZN(U3044) );
  INV_X1 U6320 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n5130) );
  AOI22_X1 U6321 ( .A1(n5149), .A2(n6462), .B1(n6461), .B2(n5148), .ZN(n5127)
         );
  OAI21_X1 U6322 ( .B1(n6466), .B2(n5193), .A(n5127), .ZN(n5128) );
  AOI21_X1 U6323 ( .B1(n5152), .B2(n6463), .A(n5128), .ZN(n5129) );
  OAI21_X1 U6324 ( .B1(n5155), .B2(n5130), .A(n5129), .ZN(U3045) );
  INV_X1 U6325 ( .A(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5135) );
  AOI22_X1 U6326 ( .A1(n5149), .A2(n5881), .B1(n6436), .B2(n5148), .ZN(n5131)
         );
  OAI21_X1 U6327 ( .B1(n5132), .B2(n5193), .A(n5131), .ZN(n5133) );
  AOI21_X1 U6328 ( .B1(n5152), .B2(n6437), .A(n5133), .ZN(n5134) );
  OAI21_X1 U6329 ( .B1(n5155), .B2(n5135), .A(n5134), .ZN(U3050) );
  INV_X1 U6330 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5139) );
  AOI22_X1 U6331 ( .A1(n5149), .A2(n6474), .B1(n6473), .B2(n5148), .ZN(n5136)
         );
  OAI21_X1 U6332 ( .B1(n6478), .B2(n5193), .A(n5136), .ZN(n5137) );
  AOI21_X1 U6333 ( .B1(n5152), .B2(n6475), .A(n5137), .ZN(n5138) );
  OAI21_X1 U6334 ( .B1(n5155), .B2(n5139), .A(n5138), .ZN(U3047) );
  INV_X1 U6335 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5143) );
  AOI22_X1 U6336 ( .A1(n5149), .A2(n6480), .B1(n6479), .B2(n5148), .ZN(n5140)
         );
  OAI21_X1 U6337 ( .B1(n6484), .B2(n5193), .A(n5140), .ZN(n5141) );
  AOI21_X1 U6338 ( .B1(n5152), .B2(n6481), .A(n5141), .ZN(n5142) );
  OAI21_X1 U6339 ( .B1(n5155), .B2(n5143), .A(n5142), .ZN(U3048) );
  INV_X1 U6340 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5147) );
  AOI22_X1 U6341 ( .A1(n5149), .A2(n6468), .B1(n6467), .B2(n5148), .ZN(n5144)
         );
  OAI21_X1 U6342 ( .B1(n6472), .B2(n5193), .A(n5144), .ZN(n5145) );
  AOI21_X1 U6343 ( .B1(n5152), .B2(n6469), .A(n5145), .ZN(n5146) );
  OAI21_X1 U6344 ( .B1(n5155), .B2(n5147), .A(n5146), .ZN(U3046) );
  INV_X1 U6345 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5154) );
  AOI22_X1 U6346 ( .A1(n5149), .A2(n6486), .B1(n6485), .B2(n5148), .ZN(n5150)
         );
  OAI21_X1 U6347 ( .B1(n6490), .B2(n5193), .A(n5150), .ZN(n5151) );
  AOI21_X1 U6348 ( .B1(n5152), .B2(n6487), .A(n5151), .ZN(n5153) );
  OAI21_X1 U6349 ( .B1(n5155), .B2(n5154), .A(n5153), .ZN(U3049) );
  OAI21_X1 U6350 ( .B1(n5156), .B2(n5158), .A(n5157), .ZN(n6131) );
  AOI22_X1 U6351 ( .A1(n5583), .A2(DATAI_9_), .B1(n6250), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n5159) );
  OAI21_X1 U6352 ( .B1(n6131), .B2(n5988), .A(n5159), .ZN(U2882) );
  XNOR2_X1 U6353 ( .A(n5161), .B(n5160), .ZN(n5231) );
  INV_X1 U6354 ( .A(n6369), .ZN(n5316) );
  OAI211_X1 U6355 ( .C1(n5316), .C2(n5162), .A(n6361), .B(n6366), .ZN(n6337)
         );
  NOR2_X1 U6356 ( .A1(n3021), .A2(n5163), .ZN(n5164) );
  OR2_X1 U6357 ( .A1(n5183), .A2(n5164), .ZN(n6137) );
  OR2_X1 U6358 ( .A1(n6338), .A2(n6582), .ZN(n5227) );
  OAI21_X1 U6359 ( .B1(n6137), .B2(n6339), .A(n5227), .ZN(n5169) );
  OR2_X1 U6360 ( .A1(n5166), .A2(n5165), .ZN(n6343) );
  OAI21_X1 U6361 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6344), .ZN(n5167) );
  NOR2_X1 U6362 ( .A1(n6343), .A2(n5167), .ZN(n5168) );
  AOI211_X1 U6363 ( .C1(n6337), .C2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n5169), 
        .B(n5168), .ZN(n5170) );
  OAI21_X1 U6364 ( .B1(n5231), .B2(n6035), .A(n5170), .ZN(U3010) );
  XOR2_X1 U6365 ( .A(n5172), .B(n5171), .Z(n6300) );
  INV_X1 U6366 ( .A(n6300), .ZN(n5176) );
  OR2_X1 U6367 ( .A1(n6338), .A2(n6580), .ZN(n6303) );
  OAI21_X1 U6368 ( .B1(n6339), .B2(n6162), .A(n6303), .ZN(n5174) );
  NOR2_X1 U6369 ( .A1(n6343), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5173)
         );
  AOI211_X1 U6370 ( .C1(n6337), .C2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n5174), 
        .B(n5173), .ZN(n5175) );
  OAI21_X1 U6371 ( .B1(n5176), .B2(n6035), .A(n5175), .ZN(U3011) );
  INV_X1 U6372 ( .A(n5177), .ZN(n5179) );
  INV_X1 U6373 ( .A(n5006), .ZN(n5178) );
  AOI21_X1 U6374 ( .B1(n5179), .B2(n5178), .A(n5156), .ZN(n6146) );
  INV_X1 U6375 ( .A(n6146), .ZN(n5181) );
  AOI22_X1 U6376 ( .A1(n5583), .A2(DATAI_8_), .B1(n6250), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n5180) );
  OAI21_X1 U6377 ( .B1(n5181), .B2(n5988), .A(n5180), .ZN(U2883) );
  OAI21_X1 U6378 ( .B1(n5183), .B2(n5182), .A(n5245), .ZN(n6127) );
  OAI222_X1 U6379 ( .A1(n6131), .A2(n6236), .B1(n5567), .B2(n5184), .C1(n5557), 
        .C2(n6127), .ZN(U2850) );
  INV_X1 U6380 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6138) );
  OAI22_X1 U6381 ( .A1(n6137), .A2(n5557), .B1(n6138), .B2(n5567), .ZN(n5185)
         );
  AOI21_X1 U6382 ( .B1(n6146), .B2(n4283), .A(n5185), .ZN(n5186) );
  INV_X1 U6383 ( .A(n5186), .ZN(U2851) );
  NOR2_X1 U6384 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5187), .ZN(n5219)
         );
  INV_X1 U6385 ( .A(n5219), .ZN(n5192) );
  AOI21_X1 U6386 ( .B1(n5194), .B2(n5193), .A(n5844), .ZN(n5188) );
  OAI21_X1 U6387 ( .B1(n5188), .B2(n5195), .A(n6623), .ZN(n5191) );
  NOR2_X1 U6388 ( .A1(n6397), .A2(n5189), .ZN(n5906) );
  INV_X1 U6389 ( .A(n5906), .ZN(n5190) );
  INV_X1 U6390 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5200) );
  AOI22_X1 U6391 ( .A1(n5220), .A2(n6468), .B1(n6467), .B2(n5219), .ZN(n5199)
         );
  INV_X1 U6392 ( .A(n5195), .ZN(n5197) );
  NAND3_X1 U6393 ( .A1(n5854), .A2(n6396), .A3(n6517), .ZN(n5196) );
  OAI21_X1 U6394 ( .B1(n5197), .B2(n5896), .A(n5196), .ZN(n5221) );
  AOI22_X1 U6395 ( .A1(n5222), .A2(n6420), .B1(n6469), .B2(n5221), .ZN(n5198)
         );
  OAI211_X1 U6396 ( .C1(n5226), .C2(n5200), .A(n5199), .B(n5198), .ZN(U3038)
         );
  INV_X1 U6397 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5203) );
  AOI22_X1 U6398 ( .A1(n5220), .A2(n6462), .B1(n6461), .B2(n5219), .ZN(n5202)
         );
  AOI22_X1 U6399 ( .A1(n5222), .A2(n6416), .B1(n6463), .B2(n5221), .ZN(n5201)
         );
  OAI211_X1 U6400 ( .C1(n5226), .C2(n5203), .A(n5202), .B(n5201), .ZN(U3037)
         );
  INV_X1 U6401 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5206) );
  AOI22_X1 U6402 ( .A1(n5220), .A2(n6486), .B1(n6485), .B2(n5219), .ZN(n5205)
         );
  AOI22_X1 U6403 ( .A1(n5222), .A2(n6432), .B1(n6487), .B2(n5221), .ZN(n5204)
         );
  OAI211_X1 U6404 ( .C1(n5226), .C2(n5206), .A(n5205), .B(n5204), .ZN(U3041)
         );
  INV_X1 U6405 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5209) );
  AOI22_X1 U6406 ( .A1(n5220), .A2(n5851), .B1(n6402), .B2(n5219), .ZN(n5208)
         );
  AOI22_X1 U6407 ( .A1(n5222), .A2(n6412), .B1(n6403), .B2(n5221), .ZN(n5207)
         );
  OAI211_X1 U6408 ( .C1(n5226), .C2(n5209), .A(n5208), .B(n5207), .ZN(U3036)
         );
  INV_X1 U6409 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5212) );
  AOI22_X1 U6410 ( .A1(n5220), .A2(n6480), .B1(n6479), .B2(n5219), .ZN(n5211)
         );
  AOI22_X1 U6411 ( .A1(n5222), .A2(n6428), .B1(n6481), .B2(n5221), .ZN(n5210)
         );
  OAI211_X1 U6412 ( .C1(n5226), .C2(n5212), .A(n5211), .B(n5210), .ZN(U3040)
         );
  INV_X1 U6413 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5215) );
  AOI22_X1 U6414 ( .A1(n5220), .A2(n6474), .B1(n6473), .B2(n5219), .ZN(n5214)
         );
  AOI22_X1 U6415 ( .A1(n5222), .A2(n6424), .B1(n6475), .B2(n5221), .ZN(n5213)
         );
  OAI211_X1 U6416 ( .C1(n5226), .C2(n5215), .A(n5214), .B(n5213), .ZN(U3039)
         );
  INV_X1 U6417 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5218) );
  AOI22_X1 U6418 ( .A1(n5220), .A2(n6493), .B1(n6492), .B2(n5219), .ZN(n5217)
         );
  AOI22_X1 U6419 ( .A1(n5222), .A2(n6444), .B1(n6496), .B2(n5221), .ZN(n5216)
         );
  OAI211_X1 U6420 ( .C1(n5226), .C2(n5218), .A(n5217), .B(n5216), .ZN(U3043)
         );
  INV_X1 U6421 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5225) );
  AOI22_X1 U6422 ( .A1(n5220), .A2(n5881), .B1(n6436), .B2(n5219), .ZN(n5224)
         );
  AOI22_X1 U6423 ( .A1(n5222), .A2(n6438), .B1(n6437), .B2(n5221), .ZN(n5223)
         );
  OAI211_X1 U6424 ( .C1(n5226), .C2(n5225), .A(n5224), .B(n5223), .ZN(U3042)
         );
  NAND2_X1 U6425 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5228)
         );
  OAI211_X1 U6426 ( .C1(n6324), .C2(n6143), .A(n5228), .B(n5227), .ZN(n5229)
         );
  AOI21_X1 U6427 ( .B1(n6146), .B2(n6319), .A(n5229), .ZN(n5230) );
  OAI21_X1 U6428 ( .B1(n6297), .B2(n5231), .A(n5230), .ZN(U2978) );
  OR2_X1 U6429 ( .A1(n6210), .A2(REIP_REG_1__SCAN_IN), .ZN(n6222) );
  NAND3_X1 U6430 ( .A1(n5247), .A2(REIP_REG_2__SCAN_IN), .A3(n6222), .ZN(n6211) );
  INV_X1 U6431 ( .A(n6174), .ZN(n5232) );
  NAND2_X1 U6432 ( .A1(n5247), .A2(n5232), .ZN(n6154) );
  NAND2_X1 U6433 ( .A1(n6152), .A2(n6154), .ZN(n6187) );
  AOI21_X1 U6434 ( .B1(n6573), .B2(n6211), .A(n6187), .ZN(n5233) );
  AOI21_X1 U6435 ( .B1(n6220), .B2(EBX_REG_3__SCAN_IN), .A(n5233), .ZN(n5234)
         );
  OAI21_X1 U6436 ( .B1(n5235), .B2(n6200), .A(n5234), .ZN(n5238) );
  OAI22_X1 U6437 ( .A1(n6206), .A2(n5236), .B1(n5832), .B2(n6202), .ZN(n5237)
         );
  AOI211_X1 U6438 ( .C1(PHYADDRPOINTER_REG_3__SCAN_IN), .C2(n6218), .A(n5238), 
        .B(n5237), .ZN(n5239) );
  OAI21_X1 U6439 ( .B1(n5240), .B2(n6227), .A(n5239), .ZN(U2824) );
  AOI21_X1 U6440 ( .B1(n5242), .B2(n5157), .A(n5241), .ZN(n5277) );
  INV_X1 U6441 ( .A(n5277), .ZN(n5263) );
  AOI22_X1 U6442 ( .A1(n5583), .A2(DATAI_10_), .B1(n6250), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5243) );
  OAI21_X1 U6443 ( .B1(n5263), .B2(n5988), .A(n5243), .ZN(U2881) );
  NOR2_X1 U6444 ( .A1(n5288), .A2(n5289), .ZN(n6142) );
  INV_X1 U6445 ( .A(n5249), .ZN(n6120) );
  NOR2_X1 U6446 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6120), .ZN(n6130) );
  OAI21_X1 U6447 ( .B1(n6142), .B2(n6130), .A(REIP_REG_10__SCAN_IN), .ZN(n5256) );
  INV_X1 U6448 ( .A(n5275), .ZN(n5254) );
  NAND2_X1 U6449 ( .A1(n5245), .A2(n5244), .ZN(n5246) );
  NAND2_X1 U6450 ( .A1(n5301), .A2(n5246), .ZN(n6340) );
  OAI22_X1 U6451 ( .A1(n6216), .A2(n4152), .B1(n6200), .B2(n6340), .ZN(n5253)
         );
  INV_X1 U6452 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5251) );
  NAND2_X1 U6453 ( .A1(n5248), .A2(n5247), .ZN(n6179) );
  INV_X1 U6454 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6585) );
  NAND3_X1 U6455 ( .A1(n5249), .A2(REIP_REG_9__SCAN_IN), .A3(n6585), .ZN(n5250) );
  OAI211_X1 U6456 ( .C1(n6205), .C2(n5251), .A(n6179), .B(n5250), .ZN(n5252)
         );
  AOI211_X1 U6457 ( .C1(n6225), .C2(n5254), .A(n5253), .B(n5252), .ZN(n5255)
         );
  OAI211_X1 U6458 ( .C1(n5263), .C2(n6167), .A(n5256), .B(n5255), .ZN(U2817)
         );
  XNOR2_X1 U6459 ( .A(n2999), .B(n6355), .ZN(n5258) );
  XNOR2_X1 U6460 ( .A(n5257), .B(n5258), .ZN(n6352) );
  NAND2_X1 U6461 ( .A1(n6352), .A2(n6332), .ZN(n5262) );
  INV_X1 U6462 ( .A(REIP_REG_9__SCAN_IN), .ZN(n5259) );
  NOR2_X1 U6463 ( .A1(n6338), .A2(n5259), .ZN(n6349) );
  AND2_X1 U6464 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5260)
         );
  AOI211_X1 U6465 ( .C1(n6132), .C2(n6310), .A(n6349), .B(n5260), .ZN(n5261)
         );
  OAI211_X1 U6466 ( .C1(n6335), .C2(n6131), .A(n5262), .B(n5261), .ZN(U2977)
         );
  OAI222_X1 U6467 ( .A1(n6340), .A2(n5557), .B1(n5567), .B2(n4152), .C1(n6236), 
        .C2(n5263), .ZN(U2849) );
  AND2_X1 U6468 ( .A1(n5265), .A2(n5264), .ZN(n5267) );
  OR2_X1 U6469 ( .A1(n5267), .A2(n5266), .ZN(n6237) );
  AOI22_X1 U6470 ( .A1(n5583), .A2(DATAI_11_), .B1(n6250), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5268) );
  OAI21_X1 U6471 ( .B1(n6237), .B2(n5988), .A(n5268), .ZN(U2880) );
  INV_X1 U6472 ( .A(n5270), .ZN(n5272) );
  NOR2_X1 U6473 ( .A1(n5272), .A2(n5271), .ZN(n5273) );
  XNOR2_X1 U6474 ( .A(n5269), .B(n5273), .ZN(n6342) );
  INV_X1 U6475 ( .A(n6342), .ZN(n5279) );
  AOI22_X1 U6476 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6376), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5274) );
  OAI21_X1 U6477 ( .B1(n5275), .B2(n6324), .A(n5274), .ZN(n5276) );
  AOI21_X1 U6478 ( .B1(n5277), .B2(n6319), .A(n5276), .ZN(n5278) );
  OAI21_X1 U6479 ( .B1(n5279), .B2(n6297), .A(n5278), .ZN(U2976) );
  XOR2_X1 U6480 ( .A(n5280), .B(n5266), .Z(n5328) );
  INV_X1 U6481 ( .A(n5328), .ZN(n5295) );
  OR2_X1 U6482 ( .A1(n5303), .A2(n5281), .ZN(n5282) );
  NAND2_X1 U6483 ( .A1(n5364), .A2(n5282), .ZN(n5317) );
  INV_X1 U6484 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5283) );
  OAI22_X1 U6485 ( .A1(n5317), .A2(n5557), .B1(n5283), .B2(n5567), .ZN(n5284)
         );
  INV_X1 U6486 ( .A(n5284), .ZN(n5285) );
  OAI21_X1 U6487 ( .B1(n5295), .B2(n6236), .A(n5285), .ZN(U2847) );
  AOI22_X1 U6488 ( .A1(n5583), .A2(DATAI_12_), .B1(n6250), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5286) );
  OAI21_X1 U6489 ( .B1(n5295), .B2(n5988), .A(n5286), .ZN(U2879) );
  INV_X1 U6490 ( .A(n5290), .ZN(n5287) );
  NOR3_X1 U6491 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6120), .A3(n5287), .ZN(n6115) );
  AOI21_X1 U6492 ( .B1(n5290), .B2(n5289), .A(n5288), .ZN(n6121) );
  AOI22_X1 U6493 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n6218), .B1(
        REIP_REG_12__SCAN_IN), .B2(n6121), .ZN(n5291) );
  OAI211_X1 U6494 ( .C1(n6200), .C2(n5317), .A(n5291), .B(n6179), .ZN(n5293)
         );
  OAI22_X1 U6495 ( .A1(n6206), .A2(n5326), .B1(n6216), .B2(n5283), .ZN(n5292)
         );
  NOR3_X1 U6496 ( .A1(n6115), .A2(n5293), .A3(n5292), .ZN(n5294) );
  OAI21_X1 U6497 ( .B1(n5295), .B2(n6167), .A(n5294), .ZN(U2815) );
  NAND2_X1 U6498 ( .A1(n5297), .A2(n5296), .ZN(n5299) );
  XOR2_X1 U6499 ( .A(n5299), .B(n5298), .Z(n6298) );
  AND2_X1 U6500 ( .A1(n5301), .A2(n5300), .ZN(n5302) );
  NOR2_X1 U6501 ( .A1(n5303), .A2(n5302), .ZN(n6234) );
  AOI21_X1 U6502 ( .B1(n5797), .B2(n6372), .A(n5304), .ZN(n6046) );
  OAI21_X1 U6503 ( .B1(n5797), .B2(n5796), .A(n5305), .ZN(n6034) );
  NOR2_X1 U6504 ( .A1(n5318), .A2(n6034), .ZN(n5314) );
  AOI21_X1 U6505 ( .B1(n6046), .B2(n5318), .A(n5314), .ZN(n5307) );
  NOR2_X1 U6506 ( .A1(n6338), .A2(n6587), .ZN(n5306) );
  AOI211_X1 U6507 ( .C1(n6234), .C2(n6382), .A(n5307), .B(n5306), .ZN(n5308)
         );
  OAI21_X1 U6508 ( .B1(n6298), .B2(n6035), .A(n5308), .ZN(U3007) );
  INV_X1 U6509 ( .A(n5310), .ZN(n5311) );
  NOR2_X1 U6510 ( .A1(n5312), .A2(n5311), .ZN(n5313) );
  XNOR2_X1 U6511 ( .A(n5309), .B(n5313), .ZN(n5330) );
  AOI211_X1 U6512 ( .C1(n5316), .C2(n5315), .A(n4161), .B(n5314), .ZN(n5322)
         );
  NAND2_X1 U6513 ( .A1(n6376), .A2(REIP_REG_12__SCAN_IN), .ZN(n5325) );
  INV_X1 U6514 ( .A(n5325), .ZN(n5321) );
  NOR2_X1 U6515 ( .A1(n5317), .A2(n6339), .ZN(n5320) );
  NOR3_X1 U6516 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6046), .A3(n5318), 
        .ZN(n5319) );
  NOR4_X1 U6517 ( .A1(n5322), .A2(n5321), .A3(n5320), .A4(n5319), .ZN(n5323)
         );
  OAI21_X1 U6518 ( .B1(n5330), .B2(n6035), .A(n5323), .ZN(U3006) );
  NAND2_X1 U6519 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5324)
         );
  OAI211_X1 U6520 ( .C1(n6324), .C2(n5326), .A(n5325), .B(n5324), .ZN(n5327)
         );
  AOI21_X1 U6521 ( .B1(n5328), .B2(n6319), .A(n5327), .ZN(n5329) );
  OAI21_X1 U6522 ( .B1(n5330), .B2(n6297), .A(n5329), .ZN(U2974) );
  AOI21_X1 U6523 ( .B1(n6534), .B2(n5331), .A(n5842), .ZN(n5341) );
  INV_X1 U6524 ( .A(n6052), .ZN(n5840) );
  NOR2_X1 U6525 ( .A1(n5332), .A2(n5840), .ZN(n5338) );
  INV_X1 U6526 ( .A(n5333), .ZN(n5336) );
  NAND3_X1 U6527 ( .A1(n4484), .A2(n6534), .A3(n5340), .ZN(n5334) );
  OAI21_X1 U6528 ( .B1(n5336), .B2(n5335), .A(n5334), .ZN(n5337) );
  INV_X1 U6529 ( .A(n5842), .ZN(n6058) );
  OAI21_X1 U6530 ( .B1(n5338), .B2(n5337), .A(n6058), .ZN(n5339) );
  OAI21_X1 U6531 ( .B1(n5341), .B2(n5340), .A(n5339), .ZN(U3459) );
  OAI21_X1 U6532 ( .B1(n5342), .B2(n5344), .A(n5343), .ZN(n5696) );
  AOI22_X1 U6533 ( .A1(n5583), .A2(DATAI_14_), .B1(n6250), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5345) );
  OAI21_X1 U6534 ( .B1(n5696), .B2(n5988), .A(n5345), .ZN(U2877) );
  NAND2_X1 U6535 ( .A1(n5362), .A2(n5346), .ZN(n5347) );
  NAND2_X1 U6536 ( .A1(n5478), .A2(n5347), .ZN(n5805) );
  OAI22_X1 U6537 ( .A1(n5805), .A2(n5557), .B1(n5348), .B2(n5567), .ZN(n5349)
         );
  INV_X1 U6538 ( .A(n5349), .ZN(n5350) );
  OAI21_X1 U6539 ( .B1(n5696), .B2(n6236), .A(n5350), .ZN(U2845) );
  NAND2_X1 U6540 ( .A1(n6152), .A2(n5351), .ZN(n6097) );
  AOI21_X1 U6541 ( .B1(n6592), .B2(n5352), .A(n6097), .ZN(n5355) );
  AOI22_X1 U6542 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6220), .B1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n6218), .ZN(n5353) );
  OAI211_X1 U6543 ( .C1(n5805), .C2(n6200), .A(n5353), .B(n6179), .ZN(n5354)
         );
  AOI211_X1 U6544 ( .C1(n5697), .C2(n6225), .A(n5355), .B(n5354), .ZN(n5356)
         );
  OAI21_X1 U6545 ( .B1(n5696), .B2(n6167), .A(n5356), .ZN(U2813) );
  NAND2_X1 U6546 ( .A1(n5357), .A2(n5358), .ZN(n5359) );
  AND2_X1 U6547 ( .A1(n5360), .A2(n5359), .ZN(n6114) );
  INV_X1 U6548 ( .A(n6114), .ZN(n5367) );
  AOI22_X1 U6549 ( .A1(n5583), .A2(DATAI_13_), .B1(n6250), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5361) );
  OAI21_X1 U6550 ( .B1(n5367), .B2(n5988), .A(n5361), .ZN(U2878) );
  INV_X1 U6551 ( .A(n5362), .ZN(n5363) );
  AOI21_X1 U6552 ( .B1(n5365), .B2(n5364), .A(n5363), .ZN(n6109) );
  AOI22_X1 U6553 ( .A1(n6109), .A2(n5569), .B1(EBX_REG_13__SCAN_IN), .B2(n5504), .ZN(n5366) );
  OAI21_X1 U6554 ( .B1(n5367), .B2(n6236), .A(n5366), .ZN(U2846) );
  AND2_X1 U6555 ( .A1(n5394), .A2(n4295), .ZN(n5368) );
  NAND2_X1 U6556 ( .A1(n5369), .A2(n5368), .ZN(n5371) );
  AOI22_X1 U6557 ( .A1(n6247), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6250), .ZN(n5370) );
  NAND2_X1 U6558 ( .A1(n5371), .A2(n5370), .ZN(U2860) );
  AOI21_X1 U6559 ( .B1(n5372), .B2(n6052), .A(n5842), .ZN(n5379) );
  NAND2_X1 U6560 ( .A1(n3358), .A2(n5373), .ZN(n5376) );
  NAND2_X1 U6561 ( .A1(n5374), .A2(n6503), .ZN(n5375) );
  NAND2_X1 U6562 ( .A1(n5376), .A2(n5375), .ZN(n6506) );
  OAI22_X1 U6563 ( .A1(n6542), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5838), .ZN(n5377) );
  AOI21_X1 U6564 ( .B1(n6506), .B2(n6052), .A(n5377), .ZN(n5378) );
  OAI22_X1 U6565 ( .A1(n5379), .A2(n6503), .B1(n5842), .B2(n5378), .ZN(U3461)
         );
  INV_X1 U6566 ( .A(n5381), .ZN(n5389) );
  INV_X1 U6567 ( .A(n5382), .ZN(n5383) );
  NAND2_X1 U6568 ( .A1(n5383), .A2(REIP_REG_30__SCAN_IN), .ZN(n5385) );
  AOI22_X1 U6569 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        EBX_REG_30__SCAN_IN), .B2(n6220), .ZN(n5384) );
  OAI211_X1 U6570 ( .C1(n5386), .C2(n6206), .A(n5385), .B(n5384), .ZN(n5388)
         );
  NOR3_X1 U6571 ( .A1(n5415), .A2(REIP_REG_30__SCAN_IN), .A3(n6793), .ZN(n5387) );
  AOI211_X1 U6572 ( .C1(n5389), .C2(n6177), .A(n5388), .B(n5387), .ZN(n5390)
         );
  OAI21_X1 U6573 ( .B1(n5397), .B2(n6167), .A(n5390), .ZN(U2797) );
  AOI22_X1 U6574 ( .A1(n6247), .A2(DATAI_30_), .B1(n6250), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5396) );
  AND2_X1 U6575 ( .A1(n5392), .A2(n5391), .ZN(n5393) );
  NAND2_X1 U6576 ( .A1(n6251), .A2(DATAI_14_), .ZN(n5395) );
  OAI211_X1 U6577 ( .C1(n5397), .C2(n5988), .A(n5396), .B(n5395), .ZN(U2861)
         );
  NAND2_X1 U6578 ( .A1(n5399), .A2(n5398), .ZN(n5404) );
  INV_X1 U6579 ( .A(n5400), .ZN(n5401) );
  NOR2_X1 U6580 ( .A1(n5402), .A2(n5401), .ZN(n5403) );
  AOI21_X1 U6581 ( .B1(n5406), .B2(n5404), .A(n5403), .ZN(n5408) );
  OR2_X1 U6582 ( .A1(n5406), .A2(n5405), .ZN(n5407) );
  AND2_X1 U6583 ( .A1(n5408), .A2(n5407), .ZN(n6522) );
  INV_X1 U6584 ( .A(n6522), .ZN(n5411) );
  AOI21_X1 U6585 ( .B1(n5409), .B2(n6558), .A(READY_N), .ZN(n6631) );
  OR2_X1 U6586 ( .A1(n5410), .A2(n6631), .ZN(n6524) );
  AND2_X1 U6587 ( .A1(n6524), .A2(n6539), .ZN(n6062) );
  MUX2_X1 U6588 ( .A(MORE_REG_SCAN_IN), .B(n5411), .S(n6062), .Z(U3471) );
  AOI21_X1 U6589 ( .B1(n5414), .B2(n5412), .A(n5413), .ZN(n5585) );
  INV_X1 U6590 ( .A(n5585), .ZN(n5573) );
  NOR2_X1 U6591 ( .A1(n5415), .A2(REIP_REG_29__SCAN_IN), .ZN(n5420) );
  AOI22_X1 U6592 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n6220), .ZN(n5417) );
  NAND2_X1 U6593 ( .A1(n6225), .A2(n5588), .ZN(n5416) );
  OAI211_X1 U6594 ( .C1(n5418), .C2(n6793), .A(n5417), .B(n5416), .ZN(n5419)
         );
  AOI211_X1 U6595 ( .C1(n5486), .C2(n6177), .A(n5420), .B(n5419), .ZN(n5421)
         );
  OAI21_X1 U6596 ( .B1(n5573), .B2(n6167), .A(n5421), .ZN(U2798) );
  INV_X1 U6597 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6808) );
  NOR2_X1 U6598 ( .A1(n5424), .A2(n5423), .ZN(n5425) );
  OR2_X1 U6599 ( .A1(n5426), .A2(n5425), .ZN(n5714) );
  AOI22_X1 U6600 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        EBX_REG_28__SCAN_IN), .B2(n6220), .ZN(n5427) );
  OAI21_X1 U6601 ( .B1(n6206), .B2(n5592), .A(n5427), .ZN(n5428) );
  AOI21_X1 U6602 ( .B1(n5429), .B2(REIP_REG_28__SCAN_IN), .A(n5428), .ZN(n5430) );
  OAI21_X1 U6603 ( .B1(n5714), .B2(n6200), .A(n5430), .ZN(n5431) );
  AOI21_X1 U6604 ( .B1(n5432), .B2(n6808), .A(n5431), .ZN(n5433) );
  OAI21_X1 U6605 ( .B1(n5602), .B2(n6167), .A(n5433), .ZN(U2799) );
  AND2_X1 U6606 ( .A1(n5944), .A2(REIP_REG_27__SCAN_IN), .ZN(n5439) );
  AOI22_X1 U6607 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6220), .B1(n5435), .B2(n6225), .ZN(n5436) );
  OAI21_X1 U6608 ( .B1(n5437), .B2(n6205), .A(n5436), .ZN(n5438) );
  NOR2_X1 U6609 ( .A1(n5439), .A2(n5438), .ZN(n5444) );
  INV_X1 U6610 ( .A(n5943), .ZN(n5442) );
  INV_X1 U6611 ( .A(n5440), .ZN(n5441) );
  NAND3_X1 U6612 ( .A1(n5442), .A2(n6748), .A3(n5441), .ZN(n5443) );
  OAI211_X1 U6613 ( .C1(n5489), .C2(n6200), .A(n5444), .B(n5443), .ZN(n5445)
         );
  INV_X1 U6614 ( .A(n5445), .ZN(n5446) );
  OAI21_X1 U6615 ( .B1(n5434), .B2(n6167), .A(n5446), .ZN(U2800) );
  INV_X1 U6616 ( .A(n5447), .ZN(n5449) );
  AOI21_X1 U6617 ( .B1(n5450), .B2(n5449), .A(n5448), .ZN(n5634) );
  INV_X1 U6618 ( .A(n5634), .ZN(n5582) );
  INV_X1 U6619 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6726) );
  NAND2_X1 U6620 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5965), .ZN(n5963) );
  INV_X1 U6621 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6660) );
  OAI21_X1 U6622 ( .B1(n6726), .B2(n5963), .A(n6660), .ZN(n5458) );
  INV_X1 U6623 ( .A(n5451), .ZN(n5953) );
  AND2_X1 U6624 ( .A1(n5519), .A2(n5452), .ZN(n5454) );
  OR2_X1 U6625 ( .A1(n5454), .A2(n5453), .ZN(n5744) );
  INV_X1 U6626 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5509) );
  OAI22_X1 U6627 ( .A1(n6216), .A2(n5509), .B1(n5632), .B2(n6205), .ZN(n5455)
         );
  AOI21_X1 U6628 ( .B1(n6225), .B2(n5630), .A(n5455), .ZN(n5456) );
  OAI21_X1 U6629 ( .B1(n5744), .B2(n6200), .A(n5456), .ZN(n5457) );
  AOI21_X1 U6630 ( .B1(n5458), .B2(n5953), .A(n5457), .ZN(n5459) );
  OAI21_X1 U6631 ( .B1(n5582), .B2(n6167), .A(n5459), .ZN(U2804) );
  OAI21_X1 U6632 ( .B1(n5460), .B2(n5462), .A(n5461), .ZN(n5654) );
  NAND2_X1 U6633 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5978) );
  INV_X1 U6634 ( .A(REIP_REG_20__SCAN_IN), .ZN(n5463) );
  OAI21_X1 U6635 ( .B1(n6083), .B2(n5978), .A(n5463), .ZN(n5472) );
  INV_X1 U6636 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5464) );
  OAI22_X1 U6637 ( .A1(n5464), .A2(n6205), .B1(n5656), .B2(n6206), .ZN(n5471)
         );
  INV_X1 U6638 ( .A(n5465), .ZN(n5537) );
  MUX2_X1 U6639 ( .A(n5537), .B(n5467), .S(n5466), .Z(n5469) );
  XNOR2_X1 U6640 ( .A(n5469), .B(n5468), .ZN(n5771) );
  INV_X1 U6641 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5529) );
  OAI22_X1 U6642 ( .A1(n5771), .A2(n6200), .B1(n6216), .B2(n5529), .ZN(n5470)
         );
  AOI211_X1 U6643 ( .C1(n5472), .C2(n5971), .A(n5471), .B(n5470), .ZN(n5473)
         );
  OAI21_X1 U6644 ( .B1(n5654), .B2(n6167), .A(n5473), .ZN(U2807) );
  AOI21_X1 U6645 ( .B1(n5475), .B2(n5343), .A(n5474), .ZN(n5476) );
  INV_X1 U6646 ( .A(n5476), .ZN(n5693) );
  INV_X1 U6647 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5481) );
  NAND2_X1 U6648 ( .A1(n6104), .A2(n5481), .ZN(n6096) );
  AND2_X1 U6649 ( .A1(n5478), .A2(n5477), .ZN(n5479) );
  NOR2_X1 U6650 ( .A1(n5563), .A2(n5479), .ZN(n6044) );
  INV_X1 U6651 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5566) );
  NOR2_X1 U6652 ( .A1(n6216), .A2(n5566), .ZN(n5483) );
  AOI22_X1 U6653 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n6218), .B1(n5688), 
        .B2(n6225), .ZN(n5480) );
  OAI211_X1 U6654 ( .C1(n5481), .C2(n6097), .A(n5480), .B(n6179), .ZN(n5482)
         );
  AOI211_X1 U6655 ( .C1(n6044), .C2(n6177), .A(n5483), .B(n5482), .ZN(n5484)
         );
  OAI211_X1 U6656 ( .C1(n5693), .C2(n6167), .A(n6096), .B(n5484), .ZN(U2812)
         );
  OAI22_X1 U6657 ( .A1(n5708), .A2(n5557), .B1(n5485), .B2(n5567), .ZN(U2828)
         );
  AOI22_X1 U6658 ( .A1(n5486), .A2(n5569), .B1(n5504), .B2(EBX_REG_29__SCAN_IN), .ZN(n5487) );
  OAI21_X1 U6659 ( .B1(n5573), .B2(n6236), .A(n5487), .ZN(U2830) );
  INV_X1 U6660 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5488) );
  OAI222_X1 U6661 ( .A1(n5488), .A2(n5567), .B1(n5557), .B2(n5714), .C1(n5602), 
        .C2(n6236), .ZN(U2831) );
  INV_X1 U6662 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5490) );
  OAI222_X1 U6663 ( .A1(n6236), .A2(n5434), .B1(n5567), .B2(n5490), .C1(n5489), 
        .C2(n5557), .ZN(U2832) );
  NAND2_X1 U6664 ( .A1(n5500), .A2(n5491), .ZN(n5492) );
  NAND2_X1 U6665 ( .A1(n5493), .A2(n5492), .ZN(n5945) );
  INV_X1 U6666 ( .A(n6007), .ZN(n5496) );
  OAI222_X1 U6667 ( .A1(n5557), .A2(n5945), .B1(n5567), .B2(n5497), .C1(n6236), 
        .C2(n5496), .ZN(U2833) );
  NAND2_X1 U6668 ( .A1(n4354), .A2(n5498), .ZN(n5499) );
  INV_X1 U6669 ( .A(n5991), .ZN(n5506) );
  INV_X1 U6670 ( .A(n5500), .ZN(n5501) );
  AOI21_X1 U6671 ( .B1(n5503), .B2(n5502), .A(n5501), .ZN(n6022) );
  AOI22_X1 U6672 ( .A1(n6022), .A2(n5569), .B1(EBX_REG_25__SCAN_IN), .B2(n5504), .ZN(n5505) );
  OAI21_X1 U6673 ( .B1(n5506), .B2(n6236), .A(n5505), .ZN(U2834) );
  OAI222_X1 U6674 ( .A1(n6236), .A2(n5620), .B1(n5567), .B2(n5508), .C1(n5507), 
        .C2(n5557), .ZN(U2835) );
  OAI22_X1 U6675 ( .A1(n5744), .A2(n5557), .B1(n5509), .B2(n5567), .ZN(n5510)
         );
  INV_X1 U6676 ( .A(n5510), .ZN(n5511) );
  OAI21_X1 U6677 ( .B1(n5582), .B2(n6236), .A(n5511), .ZN(U2836) );
  AND2_X1 U6678 ( .A1(n5513), .A2(n5514), .ZN(n5515) );
  OR2_X1 U6679 ( .A1(n5515), .A2(n5447), .ZN(n5959) );
  NAND2_X1 U6680 ( .A1(n5516), .A2(n5517), .ZN(n5518) );
  NAND2_X1 U6681 ( .A1(n5519), .A2(n5518), .ZN(n5969) );
  OAI22_X1 U6682 ( .A1(n5969), .A2(n5557), .B1(n5520), .B2(n5567), .ZN(n5521)
         );
  INV_X1 U6683 ( .A(n5521), .ZN(n5522) );
  OAI21_X1 U6684 ( .B1(n5959), .B2(n6236), .A(n5522), .ZN(U2837) );
  NAND2_X1 U6685 ( .A1(n5461), .A2(n5523), .ZN(n5524) );
  INV_X1 U6686 ( .A(n5997), .ZN(n5528) );
  OR2_X1 U6687 ( .A1(n3019), .A2(n5525), .ZN(n5526) );
  NAND2_X1 U6688 ( .A1(n5516), .A2(n5526), .ZN(n5972) );
  OAI222_X1 U6689 ( .A1(n6236), .A2(n5528), .B1(n5567), .B2(n5527), .C1(n5972), 
        .C2(n5557), .ZN(U2838) );
  OAI222_X1 U6690 ( .A1(n5654), .A2(n6236), .B1(n5567), .B2(n5529), .C1(n5557), 
        .C2(n5771), .ZN(U2839) );
  AND2_X1 U6691 ( .A1(n5531), .A2(n5532), .ZN(n5533) );
  OR2_X1 U6692 ( .A1(n5533), .A2(n5460), .ZN(n5984) );
  MUX2_X1 U6693 ( .A(n5537), .B(n5536), .S(n5535), .Z(n5544) );
  NOR2_X1 U6694 ( .A1(n5534), .A2(n5544), .ZN(n5546) );
  XNOR2_X1 U6695 ( .A(n5546), .B(n5538), .ZN(n6029) );
  INV_X1 U6696 ( .A(n6029), .ZN(n5540) );
  OAI222_X1 U6697 ( .A1(n6236), .A2(n5984), .B1(n5557), .B2(n5540), .C1(n5539), 
        .C2(n5567), .ZN(U2840) );
  NAND2_X1 U6698 ( .A1(n5541), .A2(n5542), .ZN(n5543) );
  INV_X1 U6699 ( .A(n6241), .ZN(n5548) );
  INV_X1 U6700 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5547) );
  AND2_X1 U6701 ( .A1(n5534), .A2(n5544), .ZN(n5545) );
  OR2_X1 U6702 ( .A1(n5546), .A2(n5545), .ZN(n6079) );
  OAI222_X1 U6703 ( .A1(n5548), .A2(n6236), .B1(n5567), .B2(n5547), .C1(n5557), 
        .C2(n6079), .ZN(U2841) );
  NAND2_X1 U6704 ( .A1(n5550), .A2(n5551), .ZN(n5552) );
  NAND2_X1 U6705 ( .A1(n5541), .A2(n5552), .ZN(n6088) );
  NAND2_X1 U6706 ( .A1(n5563), .A2(n5562), .ZN(n5555) );
  INV_X1 U6707 ( .A(n5553), .ZN(n5554) );
  NAND2_X1 U6708 ( .A1(n5555), .A2(n5554), .ZN(n5556) );
  NAND2_X1 U6709 ( .A1(n5556), .A2(n5534), .ZN(n6095) );
  OAI22_X1 U6710 ( .A1(n6095), .A2(n5557), .B1(n6085), .B2(n5567), .ZN(n5558)
         );
  INV_X1 U6711 ( .A(n5558), .ZN(n5559) );
  OAI21_X1 U6712 ( .B1(n6088), .B2(n6236), .A(n5559), .ZN(U2842) );
  OR2_X1 U6713 ( .A1(n5474), .A2(n5560), .ZN(n5561) );
  AND2_X1 U6714 ( .A1(n5550), .A2(n5561), .ZN(n6249) );
  INV_X1 U6715 ( .A(n6249), .ZN(n5565) );
  XNOR2_X1 U6716 ( .A(n5563), .B(n5562), .ZN(n6107) );
  INV_X1 U6717 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5564) );
  OAI222_X1 U6718 ( .A1(n5565), .A2(n6236), .B1(n5557), .B2(n6107), .C1(n5564), 
        .C2(n5567), .ZN(U2843) );
  NOR2_X1 U6719 ( .A1(n5567), .A2(n5566), .ZN(n5568) );
  AOI21_X1 U6720 ( .B1(n6044), .B2(n5569), .A(n5568), .ZN(n5570) );
  OAI21_X1 U6721 ( .B1(n5693), .B2(n6236), .A(n5570), .ZN(U2844) );
  AOI22_X1 U6722 ( .A1(n6247), .A2(DATAI_29_), .B1(n6250), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U6723 ( .A1(n6251), .A2(DATAI_13_), .ZN(n5571) );
  OAI211_X1 U6724 ( .C1(n5573), .C2(n5988), .A(n5572), .B(n5571), .ZN(U2862)
         );
  AOI22_X1 U6725 ( .A1(n6247), .A2(DATAI_28_), .B1(n6250), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U6726 ( .A1(n6251), .A2(DATAI_12_), .ZN(n5574) );
  OAI211_X1 U6727 ( .C1(n5602), .C2(n5988), .A(n5575), .B(n5574), .ZN(U2863)
         );
  AOI22_X1 U6728 ( .A1(n6247), .A2(DATAI_27_), .B1(n6250), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5577) );
  NAND2_X1 U6729 ( .A1(n6251), .A2(DATAI_11_), .ZN(n5576) );
  OAI211_X1 U6730 ( .C1(n5434), .C2(n5988), .A(n5577), .B(n5576), .ZN(U2864)
         );
  AOI22_X1 U6731 ( .A1(n6251), .A2(DATAI_8_), .B1(n6250), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U6732 ( .A1(n6247), .A2(DATAI_24_), .ZN(n5578) );
  OAI211_X1 U6733 ( .C1(n5620), .C2(n5988), .A(n5579), .B(n5578), .ZN(U2867)
         );
  AOI22_X1 U6734 ( .A1(n6247), .A2(DATAI_23_), .B1(n6250), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U6735 ( .A1(n6251), .A2(DATAI_7_), .ZN(n5580) );
  OAI211_X1 U6736 ( .C1(n5582), .C2(n5988), .A(n5581), .B(n5580), .ZN(U2868)
         );
  AOI22_X1 U6737 ( .A1(n5583), .A2(DATAI_15_), .B1(n6250), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5584) );
  OAI21_X1 U6738 ( .B1(n5693), .B2(n5988), .A(n5584), .ZN(U2876) );
  NAND2_X1 U6739 ( .A1(n5585), .A2(n6319), .ZN(n5590) );
  OAI22_X1 U6740 ( .A1(n6314), .A2(n5586), .B1(n6338), .B2(n6793), .ZN(n5587)
         );
  AOI21_X1 U6741 ( .B1(n6310), .B2(n5588), .A(n5587), .ZN(n5589) );
  OAI211_X1 U6742 ( .C1(n5591), .C2(n6297), .A(n5590), .B(n5589), .ZN(U2957)
         );
  NOR2_X1 U6743 ( .A1(n6338), .A2(n6808), .ZN(n5715) );
  NOR2_X1 U6744 ( .A1(n6324), .A2(n5592), .ZN(n5593) );
  AOI211_X1 U6745 ( .C1(PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n6330), .A(n5715), 
        .B(n5593), .ZN(n5601) );
  INV_X1 U6746 ( .A(n4260), .ZN(n5594) );
  NAND3_X1 U6747 ( .A1(n5594), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n2999), .ZN(n5597) );
  XNOR2_X1 U6748 ( .A(n5599), .B(n5598), .ZN(n5713) );
  NAND2_X1 U6749 ( .A1(n5713), .A2(n6332), .ZN(n5600) );
  OAI211_X1 U6750 ( .C1(n5602), .C2(n6335), .A(n5601), .B(n5600), .ZN(U2958)
         );
  AOI21_X1 U6751 ( .B1(n5604), .B2(n4085), .A(n5603), .ZN(n6021) );
  NAND2_X1 U6752 ( .A1(n5991), .A2(n6319), .ZN(n5609) );
  INV_X1 U6753 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5605) );
  OAI22_X1 U6754 ( .A1(n6314), .A2(n5606), .B1(n6338), .B2(n5605), .ZN(n5607)
         );
  AOI21_X1 U6755 ( .B1(n6310), .B2(n5952), .A(n5607), .ZN(n5608) );
  OAI211_X1 U6756 ( .C1(n6021), .C2(n6297), .A(n5609), .B(n5608), .ZN(U2961)
         );
  OR2_X2 U6757 ( .A1(n5659), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5660)
         );
  OAI21_X1 U6758 ( .B1(n5610), .B2(n5661), .A(n2999), .ZN(n5611) );
  NAND2_X1 U6759 ( .A1(n5660), .A2(n5611), .ZN(n5651) );
  INV_X1 U6760 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5612) );
  XNOR2_X1 U6761 ( .A(n2999), .B(n5612), .ZN(n5650) );
  OR2_X2 U6762 ( .A1(n5651), .A2(n5650), .ZN(n5626) );
  OR2_X1 U6763 ( .A1(n2999), .A2(n5612), .ZN(n5613) );
  XNOR2_X1 U6764 ( .A(n2999), .B(n5759), .ZN(n5645) );
  NOR2_X1 U6765 ( .A1(n2999), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5636)
         );
  NAND2_X1 U6766 ( .A1(n5643), .A2(n5636), .ZN(n5627) );
  INV_X1 U6767 ( .A(n5627), .ZN(n5615) );
  NAND2_X1 U6768 ( .A1(n5615), .A2(n5614), .ZN(n5618) );
  NOR2_X2 U6769 ( .A1(n5643), .A2(n5616), .ZN(n5637) );
  NAND4_X1 U6770 ( .A1(n5637), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .A4(n2999), .ZN(n5617) );
  NAND2_X1 U6771 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  XNOR2_X1 U6772 ( .A(n5619), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5739)
         );
  INV_X1 U6773 ( .A(n5620), .ZN(n5624) );
  NOR2_X1 U6774 ( .A1(n6338), .A2(n6771), .ZN(n5736) );
  AOI21_X1 U6775 ( .B1(n6330), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5736), 
        .ZN(n5621) );
  OAI21_X1 U6776 ( .B1(n5622), .B2(n6324), .A(n5621), .ZN(n5623) );
  AOI21_X1 U6777 ( .B1(n5624), .B2(n6319), .A(n5623), .ZN(n5625) );
  OAI21_X1 U6778 ( .B1(n5739), .B2(n6297), .A(n5625), .ZN(U2962) );
  NAND2_X1 U6779 ( .A1(n5741), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5628) );
  OAI21_X1 U6780 ( .B1(n5653), .B2(n5628), .A(n5627), .ZN(n5629) );
  XNOR2_X1 U6781 ( .A(n5629), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5747)
         );
  NAND2_X1 U6782 ( .A1(n6310), .A2(n5630), .ZN(n5631) );
  NAND2_X1 U6783 ( .A1(n6376), .A2(REIP_REG_23__SCAN_IN), .ZN(n5743) );
  OAI211_X1 U6784 ( .C1(n6314), .C2(n5632), .A(n5631), .B(n5743), .ZN(n5633)
         );
  AOI21_X1 U6785 ( .B1(n5634), .B2(n6319), .A(n5633), .ZN(n5635) );
  OAI21_X1 U6786 ( .B1(n5747), .B2(n6297), .A(n5635), .ZN(U2963) );
  AOI21_X1 U6787 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n2999), .A(n5636), 
        .ZN(n5638) );
  XOR2_X1 U6788 ( .A(n5638), .B(n5637), .Z(n5755) );
  INV_X1 U6789 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U6790 ( .A1(n6376), .A2(REIP_REG_22__SCAN_IN), .ZN(n5750) );
  OAI21_X1 U6791 ( .B1(n6314), .B2(n5639), .A(n5750), .ZN(n5641) );
  NOR2_X1 U6792 ( .A1(n5959), .A2(n6335), .ZN(n5640) );
  AOI211_X1 U6793 ( .C1(n6310), .C2(n5960), .A(n5641), .B(n5640), .ZN(n5642)
         );
  OAI21_X1 U6794 ( .B1(n5755), .B2(n6297), .A(n5642), .ZN(U2964) );
  AOI21_X1 U6795 ( .B1(n5645), .B2(n5644), .A(n5643), .ZN(n5762) );
  INV_X1 U6796 ( .A(n5970), .ZN(n5647) );
  AOI22_X1 U6797 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .B1(n6376), 
        .B2(REIP_REG_21__SCAN_IN), .ZN(n5646) );
  OAI21_X1 U6798 ( .B1(n5647), .B2(n6324), .A(n5646), .ZN(n5648) );
  AOI21_X1 U6799 ( .B1(n5997), .B2(n6319), .A(n5648), .ZN(n5649) );
  OAI21_X1 U6800 ( .B1(n5762), .B2(n6297), .A(n5649), .ZN(U2965) );
  NAND2_X1 U6801 ( .A1(n5651), .A2(n5650), .ZN(n5652) );
  NAND2_X1 U6802 ( .A1(n5653), .A2(n5652), .ZN(n5776) );
  INV_X1 U6803 ( .A(n5654), .ZN(n6000) );
  OR2_X1 U6804 ( .A1(n6338), .A2(n5463), .ZN(n5769) );
  NAND2_X1 U6805 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5655)
         );
  OAI211_X1 U6806 ( .C1(n6324), .C2(n5656), .A(n5769), .B(n5655), .ZN(n5657)
         );
  AOI21_X1 U6807 ( .B1(n6000), .B2(n6319), .A(n5657), .ZN(n5658) );
  OAI21_X1 U6808 ( .B1(n5776), .B2(n6297), .A(n5658), .ZN(U2966) );
  INV_X1 U6809 ( .A(n5659), .ZN(n5662) );
  OAI21_X1 U6810 ( .B1(n5662), .B2(n5661), .A(n5660), .ZN(n5663) );
  XNOR2_X1 U6811 ( .A(n5663), .B(n5670), .ZN(n6030) );
  NAND2_X1 U6812 ( .A1(n6030), .A2(n6332), .ZN(n5667) );
  INV_X1 U6813 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5664) );
  OAI22_X1 U6814 ( .A1(n6314), .A2(n5982), .B1(n6338), .B2(n5664), .ZN(n5665)
         );
  AOI21_X1 U6815 ( .B1(n6310), .B2(n5980), .A(n5665), .ZN(n5666) );
  OAI211_X1 U6816 ( .C1(n6335), .C2(n5984), .A(n5667), .B(n5666), .ZN(U2967)
         );
  AND2_X1 U6817 ( .A1(n2999), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5778)
         );
  INV_X1 U6818 ( .A(n5668), .ZN(n5681) );
  NAND2_X1 U6819 ( .A1(n5670), .A2(n5792), .ZN(n5671) );
  NOR3_X1 U6820 ( .A1(n3045), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5671), 
        .ZN(n5777) );
  INV_X1 U6821 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6042) );
  OR2_X1 U6822 ( .A1(n2999), .A2(n6042), .ZN(n5678) );
  INV_X1 U6823 ( .A(n5671), .ZN(n5672) );
  AOI211_X1 U6824 ( .C1(n5681), .C2(n5678), .A(n5778), .B(n5672), .ZN(n5673)
         );
  AOI211_X1 U6825 ( .C1(n5778), .C2(n5681), .A(n5777), .B(n5673), .ZN(n5795)
         );
  NAND2_X1 U6826 ( .A1(n6376), .A2(REIP_REG_17__SCAN_IN), .ZN(n5789) );
  OAI21_X1 U6827 ( .B1(n6314), .B2(n6084), .A(n5789), .ZN(n5675) );
  NOR2_X1 U6828 ( .A1(n6088), .A2(n6335), .ZN(n5674) );
  AOI211_X1 U6829 ( .C1(n6310), .C2(n6087), .A(n5675), .B(n5674), .ZN(n5676)
         );
  OAI21_X1 U6830 ( .B1(n5795), .B2(n6297), .A(n5676), .ZN(U2969) );
  INV_X1 U6831 ( .A(n5678), .ZN(n5680) );
  AND2_X1 U6832 ( .A1(n5678), .A2(n5677), .ZN(n5679) );
  OAI22_X1 U6833 ( .A1(n5681), .A2(n5680), .B1(n3008), .B2(n5679), .ZN(n6036)
         );
  INV_X1 U6834 ( .A(n6098), .ZN(n5683) );
  AOI22_X1 U6835 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6376), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5682) );
  OAI21_X1 U6836 ( .B1(n5683), .B2(n6324), .A(n5682), .ZN(n5684) );
  AOI21_X1 U6837 ( .B1(n6249), .B2(n6319), .A(n5684), .ZN(n5685) );
  OAI21_X1 U6838 ( .B1(n6036), .B2(n6297), .A(n5685), .ZN(U2970) );
  NOR2_X1 U6839 ( .A1(n6338), .A2(n5481), .ZN(n6043) );
  NOR2_X1 U6840 ( .A1(n6314), .A2(n5686), .ZN(n5687) );
  AOI211_X1 U6841 ( .C1(n6310), .C2(n5688), .A(n6043), .B(n5687), .ZN(n5692)
         );
  OAI21_X1 U6842 ( .B1(n5690), .B2(n5689), .A(n3045), .ZN(n6048) );
  NAND2_X1 U6843 ( .A1(n6048), .A2(n6332), .ZN(n5691) );
  OAI211_X1 U6844 ( .C1(n5693), .C2(n6335), .A(n5692), .B(n5691), .ZN(U2971)
         );
  XNOR2_X1 U6845 ( .A(n2999), .B(n5803), .ZN(n5695) );
  XNOR2_X1 U6846 ( .A(n5694), .B(n5695), .ZN(n5809) );
  INV_X1 U6847 ( .A(n5696), .ZN(n5701) );
  INV_X1 U6848 ( .A(n5697), .ZN(n5699) );
  AOI22_X1 U6849 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6376), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5698) );
  OAI21_X1 U6850 ( .B1(n6324), .B2(n5699), .A(n5698), .ZN(n5700) );
  AOI21_X1 U6851 ( .B1(n5701), .B2(n6319), .A(n5700), .ZN(n5702) );
  OAI21_X1 U6852 ( .B1(n5809), .B2(n6297), .A(n5702), .ZN(U2972) );
  NOR3_X1 U6853 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n5704), .A3(n5703), 
        .ZN(n5706) );
  AOI211_X1 U6854 ( .C1(n5707), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5706), .B(n5705), .ZN(n5711) );
  INV_X1 U6855 ( .A(n5708), .ZN(n5709) );
  NAND2_X1 U6856 ( .A1(n5709), .A2(n6382), .ZN(n5710) );
  OAI211_X1 U6857 ( .C1(n5712), .C2(n6035), .A(n5711), .B(n5710), .ZN(U2987)
         );
  INV_X1 U6858 ( .A(n5713), .ZN(n5724) );
  INV_X1 U6859 ( .A(n5714), .ZN(n5716) );
  AOI21_X1 U6860 ( .B1(n5716), .B2(n6382), .A(n5715), .ZN(n5723) );
  OAI21_X1 U6861 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5717), .ZN(n5718) );
  INV_X1 U6862 ( .A(n5718), .ZN(n5720) );
  AOI22_X1 U6863 ( .A1(n5721), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .B1(n5720), .B2(n5719), .ZN(n5722) );
  OAI211_X1 U6864 ( .C1(n5724), .C2(n6035), .A(n5723), .B(n5722), .ZN(U2990)
         );
  XNOR2_X1 U6865 ( .A(n2999), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5725)
         );
  XNOR2_X1 U6866 ( .A(n4260), .B(n5725), .ZN(n6006) );
  INV_X1 U6867 ( .A(n6006), .ZN(n5732) );
  INV_X1 U6868 ( .A(n6027), .ZN(n5730) );
  AOI211_X1 U6869 ( .C1(n5595), .C2(n6026), .A(n5726), .B(n6019), .ZN(n5729)
         );
  INV_X1 U6870 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5727) );
  OAI22_X1 U6871 ( .A1(n5945), .A2(n6339), .B1(n6338), .B2(n5727), .ZN(n5728)
         );
  AOI211_X1 U6872 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5730), .A(n5729), .B(n5728), .ZN(n5731) );
  OAI21_X1 U6873 ( .B1(n5732), .B2(n6035), .A(n5731), .ZN(U2992) );
  NAND3_X1 U6874 ( .A1(n5760), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n5741), .ZN(n5733) );
  AOI21_X1 U6875 ( .B1(n5734), .B2(n5733), .A(n6027), .ZN(n5735) );
  AOI211_X1 U6876 ( .C1(n6382), .C2(n5737), .A(n5736), .B(n5735), .ZN(n5738)
         );
  OAI21_X1 U6877 ( .B1(n5739), .B2(n6035), .A(n5738), .ZN(U2994) );
  INV_X1 U6878 ( .A(n5740), .ZN(n5753) );
  NAND3_X1 U6879 ( .A1(n5760), .A2(n5741), .A3(n5614), .ZN(n5742) );
  OAI211_X1 U6880 ( .C1(n5744), .C2(n6339), .A(n5743), .B(n5742), .ZN(n5745)
         );
  AOI21_X1 U6881 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5753), .A(n5745), 
        .ZN(n5746) );
  OAI21_X1 U6882 ( .B1(n5747), .B2(n6035), .A(n5746), .ZN(U2995) );
  INV_X1 U6883 ( .A(n5748), .ZN(n5749) );
  NAND2_X1 U6884 ( .A1(n5749), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5751) );
  OAI211_X1 U6885 ( .C1(n5969), .C2(n6339), .A(n5751), .B(n5750), .ZN(n5752)
         );
  AOI21_X1 U6886 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5753), .A(n5752), 
        .ZN(n5754) );
  OAI21_X1 U6887 ( .B1(n5755), .B2(n6035), .A(n5754), .ZN(U2996) );
  NOR2_X1 U6888 ( .A1(n5756), .A2(n5759), .ZN(n5758) );
  INV_X1 U6889 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6750) );
  OAI22_X1 U6890 ( .A1(n5972), .A2(n6339), .B1(n6750), .B2(n6338), .ZN(n5757)
         );
  AOI211_X1 U6891 ( .C1(n5760), .C2(n5759), .A(n5758), .B(n5757), .ZN(n5761)
         );
  OAI21_X1 U6892 ( .B1(n5762), .B2(n6035), .A(n5761), .ZN(U2997) );
  NOR2_X1 U6893 ( .A1(n6046), .A2(n5763), .ZN(n5793) );
  NAND2_X1 U6894 ( .A1(n5767), .A2(n5793), .ZN(n6033) );
  NOR2_X1 U6895 ( .A1(n5764), .A2(n6033), .ZN(n5773) );
  AOI21_X1 U6896 ( .B1(n6372), .B2(n5765), .A(n5788), .ZN(n5766) );
  OAI21_X1 U6897 ( .B1(n5768), .B2(n5767), .A(n5766), .ZN(n6028) );
  NAND2_X1 U6898 ( .A1(n6028), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5770) );
  OAI211_X1 U6899 ( .C1(n5771), .C2(n6339), .A(n5770), .B(n5769), .ZN(n5772)
         );
  AOI21_X1 U6900 ( .B1(n5774), .B2(n5773), .A(n5772), .ZN(n5775) );
  OAI21_X1 U6901 ( .B1(n5776), .B2(n6035), .A(n5775), .ZN(U2998) );
  AOI21_X1 U6902 ( .B1(n5668), .B2(n5778), .A(n5777), .ZN(n5779) );
  XNOR2_X1 U6903 ( .A(n5779), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6011)
         );
  NOR2_X1 U6904 ( .A1(n5780), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5781)
         );
  OAI21_X1 U6905 ( .B1(n5781), .B2(n5788), .A(INSTADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n5785) );
  NOR2_X1 U6906 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6046), .ZN(n5782)
         );
  AOI22_X1 U6907 ( .A1(n5783), .A2(n5782), .B1(n6376), .B2(
        REIP_REG_18__SCAN_IN), .ZN(n5784) );
  OAI211_X1 U6908 ( .C1(n6339), .C2(n6079), .A(n5785), .B(n5784), .ZN(n5786)
         );
  AOI21_X1 U6909 ( .B1(n6011), .B2(n6383), .A(n5786), .ZN(n5787) );
  INV_X1 U6910 ( .A(n5787), .ZN(U3000) );
  NAND2_X1 U6911 ( .A1(n5788), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5790) );
  OAI211_X1 U6912 ( .C1(n6339), .C2(n6095), .A(n5790), .B(n5789), .ZN(n5791)
         );
  AOI21_X1 U6913 ( .B1(n5793), .B2(n5792), .A(n5791), .ZN(n5794) );
  OAI21_X1 U6914 ( .B1(n5795), .B2(n6035), .A(n5794), .ZN(U3001) );
  NAND2_X1 U6915 ( .A1(n5798), .A2(n5796), .ZN(n6387) );
  NAND2_X1 U6916 ( .A1(n6372), .A2(n5797), .ZN(n5800) );
  OR3_X1 U6917 ( .A1(n6371), .A2(n5798), .A3(n5816), .ZN(n5799) );
  AOI211_X1 U6918 ( .C1(n5800), .C2(n5799), .A(INSTADDRPOINTER_REG_13__SCAN_IN), .B(n5815), .ZN(n5814) );
  AOI211_X1 U6919 ( .C1(n5815), .C2(n6387), .A(n5814), .B(n6034), .ZN(n5801)
         );
  OAI21_X1 U6920 ( .B1(n5804), .B2(n6385), .A(n5801), .ZN(n5813) );
  INV_X1 U6921 ( .A(n6046), .ZN(n5802) );
  AND3_X1 U6922 ( .A1(n5804), .A2(n5803), .A3(n5802), .ZN(n5807) );
  OAI22_X1 U6923 ( .A1(n5805), .A2(n6339), .B1(n6592), .B2(n6338), .ZN(n5806)
         );
  AOI211_X1 U6924 ( .C1(n5813), .C2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n5807), .B(n5806), .ZN(n5808) );
  OAI21_X1 U6925 ( .B1(n5809), .B2(n6035), .A(n5808), .ZN(U3004) );
  OAI21_X1 U6926 ( .B1(n5812), .B2(n5811), .A(n5810), .ZN(n6015) );
  INV_X1 U6927 ( .A(n6015), .ZN(n5820) );
  OAI21_X1 U6928 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5814), .A(n5813), 
        .ZN(n5819) );
  NOR4_X1 U6929 ( .A1(n6385), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n5816), 
        .A4(n5815), .ZN(n5817) );
  NOR2_X1 U6930 ( .A1(n6338), .A2(n6590), .ZN(n6016) );
  AOI211_X1 U6931 ( .C1(n6109), .C2(n6382), .A(n5817), .B(n6016), .ZN(n5818)
         );
  OAI211_X1 U6932 ( .C1(n5820), .C2(n6035), .A(n5819), .B(n5818), .ZN(U3005)
         );
  OAI211_X1 U6933 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n5821), .A(n5825), .B(
        n6408), .ZN(n5822) );
  OAI21_X1 U6934 ( .B1(n5833), .B2(n5823), .A(n5822), .ZN(n5824) );
  MUX2_X1 U6935 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5824), .S(n6393), 
        .Z(U3464) );
  XNOR2_X1 U6936 ( .A(n5826), .B(n5825), .ZN(n5827) );
  INV_X1 U6937 ( .A(n4504), .ZN(n6203) );
  OAI22_X1 U6938 ( .A1(n5827), .A2(n5896), .B1(n6203), .B2(n5833), .ZN(n5828)
         );
  MUX2_X1 U6939 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5828), .S(n6393), 
        .Z(U3463) );
  NOR2_X1 U6940 ( .A1(n5830), .A2(n5829), .ZN(n5831) );
  OAI222_X1 U6941 ( .A1(n5835), .A2(n5834), .B1(n5833), .B2(n5832), .C1(n5896), 
        .C2(n5831), .ZN(n5836) );
  MUX2_X1 U6942 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5836), .S(n6393), 
        .Z(U3462) );
  INV_X1 U6943 ( .A(n5837), .ZN(n5841) );
  OAI22_X1 U6944 ( .A1(n5841), .A2(n5840), .B1(n5839), .B2(n5838), .ZN(n5843)
         );
  MUX2_X1 U6945 ( .A(n5843), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n5842), 
        .Z(U3456) );
  NOR3_X1 U6946 ( .A1(n5889), .A2(n5887), .A3(n5896), .ZN(n5845) );
  NOR2_X1 U6947 ( .A1(n5845), .A2(n5844), .ZN(n5850) );
  NOR2_X1 U6948 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5846), .ZN(n5888)
         );
  INV_X1 U6949 ( .A(n5888), .ZN(n5848) );
  AOI211_X1 U6950 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5848), .A(n6397), .B(
        n5847), .ZN(n5849) );
  NAND2_X1 U6951 ( .A1(n5886), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5860) );
  AOI22_X1 U6952 ( .A1(n6402), .A2(n5888), .B1(n6412), .B2(n5887), .ZN(n5859)
         );
  NAND2_X1 U6953 ( .A1(n5889), .A2(n5851), .ZN(n5858) );
  NAND2_X1 U6954 ( .A1(n5852), .A2(n6408), .ZN(n5856) );
  NAND2_X1 U6955 ( .A1(n5854), .A2(n5853), .ZN(n5855) );
  NAND2_X1 U6956 ( .A1(n5856), .A2(n5855), .ZN(n5890) );
  NAND2_X1 U6957 ( .A1(n6403), .A2(n5890), .ZN(n5857) );
  NAND4_X1 U6958 ( .A1(n5860), .A2(n5859), .A3(n5858), .A4(n5857), .ZN(U3020)
         );
  NAND2_X1 U6959 ( .A1(n5886), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5864) );
  AOI22_X1 U6960 ( .A1(n6461), .A2(n5888), .B1(n6416), .B2(n5887), .ZN(n5863)
         );
  NAND2_X1 U6961 ( .A1(n5889), .A2(n6462), .ZN(n5862) );
  NAND2_X1 U6962 ( .A1(n6463), .A2(n5890), .ZN(n5861) );
  NAND4_X1 U6963 ( .A1(n5864), .A2(n5863), .A3(n5862), .A4(n5861), .ZN(U3021)
         );
  NAND2_X1 U6964 ( .A1(n5886), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5868) );
  AOI22_X1 U6965 ( .A1(n6467), .A2(n5888), .B1(n6420), .B2(n5887), .ZN(n5867)
         );
  NAND2_X1 U6966 ( .A1(n5889), .A2(n6468), .ZN(n5866) );
  NAND2_X1 U6967 ( .A1(n6469), .A2(n5890), .ZN(n5865) );
  NAND4_X1 U6968 ( .A1(n5868), .A2(n5867), .A3(n5866), .A4(n5865), .ZN(U3022)
         );
  NAND2_X1 U6969 ( .A1(n5886), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5872) );
  AOI22_X1 U6970 ( .A1(n6473), .A2(n5888), .B1(n6424), .B2(n5887), .ZN(n5871)
         );
  NAND2_X1 U6971 ( .A1(n5889), .A2(n6474), .ZN(n5870) );
  NAND2_X1 U6972 ( .A1(n6475), .A2(n5890), .ZN(n5869) );
  NAND4_X1 U6973 ( .A1(n5872), .A2(n5871), .A3(n5870), .A4(n5869), .ZN(U3023)
         );
  NAND2_X1 U6974 ( .A1(n5886), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5876) );
  AOI22_X1 U6975 ( .A1(n6479), .A2(n5888), .B1(n6428), .B2(n5887), .ZN(n5875)
         );
  NAND2_X1 U6976 ( .A1(n5889), .A2(n6480), .ZN(n5874) );
  NAND2_X1 U6977 ( .A1(n6481), .A2(n5890), .ZN(n5873) );
  NAND4_X1 U6978 ( .A1(n5876), .A2(n5875), .A3(n5874), .A4(n5873), .ZN(U3024)
         );
  NAND2_X1 U6979 ( .A1(n5886), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5880) );
  AOI22_X1 U6980 ( .A1(n6485), .A2(n5888), .B1(n6432), .B2(n5887), .ZN(n5879)
         );
  NAND2_X1 U6981 ( .A1(n5889), .A2(n6486), .ZN(n5878) );
  NAND2_X1 U6982 ( .A1(n6487), .A2(n5890), .ZN(n5877) );
  NAND4_X1 U6983 ( .A1(n5880), .A2(n5879), .A3(n5878), .A4(n5877), .ZN(U3025)
         );
  NAND2_X1 U6984 ( .A1(n5886), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5885) );
  AOI22_X1 U6985 ( .A1(n6436), .A2(n5888), .B1(n6438), .B2(n5887), .ZN(n5884)
         );
  NAND2_X1 U6986 ( .A1(n5889), .A2(n5881), .ZN(n5883) );
  NAND2_X1 U6987 ( .A1(n6437), .A2(n5890), .ZN(n5882) );
  NAND4_X1 U6988 ( .A1(n5885), .A2(n5884), .A3(n5883), .A4(n5882), .ZN(U3026)
         );
  NAND2_X1 U6989 ( .A1(n5886), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5894) );
  AOI22_X1 U6990 ( .A1(n6492), .A2(n5888), .B1(n6444), .B2(n5887), .ZN(n5893)
         );
  NAND2_X1 U6991 ( .A1(n5889), .A2(n6493), .ZN(n5892) );
  NAND2_X1 U6992 ( .A1(n6496), .A2(n5890), .ZN(n5891) );
  NAND4_X1 U6993 ( .A1(n5894), .A2(n5893), .A3(n5892), .A4(n5891), .ZN(U3027)
         );
  INV_X1 U6994 ( .A(n6500), .ZN(n5895) );
  AOI21_X1 U6995 ( .B1(n5897), .B2(STATEBS16_REG_SCAN_IN), .A(n5896), .ZN(
        n5904) );
  NOR2_X1 U6996 ( .A1(n5898), .A2(n6517), .ZN(n5899) );
  NOR2_X1 U6997 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5900), .ZN(n5936)
         );
  INV_X1 U6998 ( .A(n5901), .ZN(n5903) );
  INV_X1 U6999 ( .A(n5936), .ZN(n5902) );
  AOI22_X1 U7000 ( .A1(n5904), .A2(n5903), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5902), .ZN(n5905) );
  OAI211_X1 U7001 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6633), .A(n5906), .B(n5905), .ZN(n5935) );
  AOI22_X1 U7002 ( .A1(n6402), .A2(n5936), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5935), .ZN(n5907) );
  OAI21_X1 U7003 ( .B1(n6500), .B2(n6415), .A(n5907), .ZN(n5908) );
  AOI21_X1 U7004 ( .B1(n6412), .B2(n5939), .A(n5908), .ZN(n5909) );
  OAI21_X1 U7005 ( .B1(n5942), .B2(n5910), .A(n5909), .ZN(U3100) );
  AOI22_X1 U7006 ( .A1(n6461), .A2(n5936), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5935), .ZN(n5911) );
  OAI21_X1 U7007 ( .B1(n6500), .B2(n6419), .A(n5911), .ZN(n5912) );
  AOI21_X1 U7008 ( .B1(n6416), .B2(n5939), .A(n5912), .ZN(n5913) );
  OAI21_X1 U7009 ( .B1(n5942), .B2(n5914), .A(n5913), .ZN(U3101) );
  AOI22_X1 U7010 ( .A1(n6467), .A2(n5936), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5935), .ZN(n5915) );
  OAI21_X1 U7011 ( .B1(n6500), .B2(n6423), .A(n5915), .ZN(n5916) );
  AOI21_X1 U7012 ( .B1(n6420), .B2(n5939), .A(n5916), .ZN(n5917) );
  OAI21_X1 U7013 ( .B1(n5942), .B2(n5918), .A(n5917), .ZN(U3102) );
  AOI22_X1 U7014 ( .A1(n6473), .A2(n5936), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5935), .ZN(n5919) );
  OAI21_X1 U7015 ( .B1(n6500), .B2(n6427), .A(n5919), .ZN(n5920) );
  AOI21_X1 U7016 ( .B1(n6424), .B2(n5939), .A(n5920), .ZN(n5921) );
  OAI21_X1 U7017 ( .B1(n5942), .B2(n5922), .A(n5921), .ZN(U3103) );
  AOI22_X1 U7018 ( .A1(n6479), .A2(n5936), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5935), .ZN(n5923) );
  OAI21_X1 U7019 ( .B1(n6500), .B2(n6431), .A(n5923), .ZN(n5924) );
  AOI21_X1 U7020 ( .B1(n6428), .B2(n5939), .A(n5924), .ZN(n5925) );
  OAI21_X1 U7021 ( .B1(n5942), .B2(n5926), .A(n5925), .ZN(U3104) );
  AOI22_X1 U7022 ( .A1(n6485), .A2(n5936), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5935), .ZN(n5927) );
  OAI21_X1 U7023 ( .B1(n6500), .B2(n6435), .A(n5927), .ZN(n5928) );
  AOI21_X1 U7024 ( .B1(n6432), .B2(n5939), .A(n5928), .ZN(n5929) );
  OAI21_X1 U7025 ( .B1(n5942), .B2(n5930), .A(n5929), .ZN(U3105) );
  AOI22_X1 U7026 ( .A1(n6436), .A2(n5936), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5935), .ZN(n5931) );
  OAI21_X1 U7027 ( .B1(n6500), .B2(n6441), .A(n5931), .ZN(n5932) );
  AOI21_X1 U7028 ( .B1(n6438), .B2(n5939), .A(n5932), .ZN(n5933) );
  OAI21_X1 U7029 ( .B1(n5942), .B2(n5934), .A(n5933), .ZN(U3106) );
  AOI22_X1 U7030 ( .A1(n6492), .A2(n5936), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5935), .ZN(n5937) );
  OAI21_X1 U7031 ( .B1(n6500), .B2(n6449), .A(n5937), .ZN(n5938) );
  AOI21_X1 U7032 ( .B1(n6444), .B2(n5939), .A(n5938), .ZN(n5940) );
  OAI21_X1 U7033 ( .B1(n5942), .B2(n5941), .A(n5940), .ZN(U3107) );
  AND2_X1 U7034 ( .A1(n6274), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U7035 ( .A1(EBX_REG_26__SCAN_IN), .A2(n6220), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6218), .ZN(n5950) );
  NOR2_X1 U7036 ( .A1(n6771), .A2(n5943), .ZN(n5951) );
  AOI21_X1 U7037 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5951), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5947) );
  INV_X1 U7038 ( .A(n5944), .ZN(n5946) );
  OAI22_X1 U7039 ( .A1(n5947), .A2(n5946), .B1(n5945), .B2(n6200), .ZN(n5948)
         );
  AOI21_X1 U7040 ( .B1(n6007), .B2(n6145), .A(n5948), .ZN(n5949) );
  OAI211_X1 U7041 ( .C1(n6010), .C2(n6206), .A(n5950), .B(n5949), .ZN(U2801)
         );
  AOI22_X1 U7042 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6220), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6218), .ZN(n5958) );
  AOI22_X1 U7043 ( .A1(n5952), .A2(n6225), .B1(n5951), .B2(n5605), .ZN(n5957)
         );
  AOI22_X1 U7044 ( .A1(n5991), .A2(n6145), .B1(n6177), .B2(n6022), .ZN(n5956)
         );
  OAI21_X1 U7045 ( .B1(n5954), .B2(n5953), .A(REIP_REG_25__SCAN_IN), .ZN(n5955) );
  NAND4_X1 U7046 ( .A1(n5958), .A2(n5957), .A3(n5956), .A4(n5955), .ZN(U2802)
         );
  INV_X1 U7047 ( .A(n5959), .ZN(n5994) );
  AOI22_X1 U7048 ( .A1(n6225), .A2(n5960), .B1(EBX_REG_22__SCAN_IN), .B2(n6220), .ZN(n5962) );
  NAND2_X1 U7049 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5961)
         );
  OAI211_X1 U7050 ( .C1(n5963), .C2(REIP_REG_22__SCAN_IN), .A(n5962), .B(n5961), .ZN(n5964) );
  AOI21_X1 U7051 ( .B1(n5994), .B2(n6145), .A(n5964), .ZN(n5968) );
  NAND2_X1 U7052 ( .A1(n6750), .A2(n5965), .ZN(n5974) );
  INV_X1 U7053 ( .A(n5974), .ZN(n5966) );
  OAI21_X1 U7054 ( .B1(n5971), .B2(n5966), .A(REIP_REG_22__SCAN_IN), .ZN(n5967) );
  OAI211_X1 U7055 ( .C1(n6200), .C2(n5969), .A(n5968), .B(n5967), .ZN(U2805)
         );
  AOI22_X1 U7056 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6220), .B1(n5970), .B2(n6225), .ZN(n5977) );
  AOI22_X1 U7057 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n6218), .B1(
        REIP_REG_21__SCAN_IN), .B2(n5971), .ZN(n5976) );
  NOR2_X1 U7058 ( .A1(n5972), .A2(n6200), .ZN(n5973) );
  AOI21_X1 U7059 ( .B1(n5997), .B2(n6145), .A(n5973), .ZN(n5975) );
  NAND4_X1 U7060 ( .A1(n5977), .A2(n5976), .A3(n5975), .A4(n5974), .ZN(U2806)
         );
  OAI21_X1 U7061 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n5978), .ZN(n5987) );
  INV_X1 U7062 ( .A(n5979), .ZN(n6092) );
  AOI22_X1 U7063 ( .A1(n5980), .A2(n6225), .B1(REIP_REG_19__SCAN_IN), .B2(
        n6092), .ZN(n5981) );
  OAI211_X1 U7064 ( .C1(n6205), .C2(n5982), .A(n5981), .B(n6179), .ZN(n5983)
         );
  AOI21_X1 U7065 ( .B1(EBX_REG_19__SCAN_IN), .B2(n6220), .A(n5983), .ZN(n5986)
         );
  INV_X1 U7066 ( .A(n5984), .ZN(n6003) );
  AOI22_X1 U7067 ( .A1(n6003), .A2(n6145), .B1(n6177), .B2(n6029), .ZN(n5985)
         );
  OAI211_X1 U7068 ( .C1(n6083), .C2(n5987), .A(n5986), .B(n5985), .ZN(U2808)
         );
  AOI22_X1 U7069 ( .A1(n6007), .A2(n6248), .B1(n6247), .B2(DATAI_26_), .ZN(
        n5990) );
  AOI22_X1 U7070 ( .A1(n6251), .A2(DATAI_10_), .B1(n6250), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5989) );
  NAND2_X1 U7071 ( .A1(n5990), .A2(n5989), .ZN(U2865) );
  AOI22_X1 U7072 ( .A1(n5991), .A2(n6248), .B1(n6247), .B2(DATAI_25_), .ZN(
        n5993) );
  AOI22_X1 U7073 ( .A1(n6251), .A2(DATAI_9_), .B1(n6250), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7074 ( .A1(n5993), .A2(n5992), .ZN(U2866) );
  AOI22_X1 U7075 ( .A1(n5994), .A2(n6248), .B1(n6247), .B2(DATAI_22_), .ZN(
        n5996) );
  AOI22_X1 U7076 ( .A1(n6251), .A2(DATAI_6_), .B1(n6250), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7077 ( .A1(n5996), .A2(n5995), .ZN(U2869) );
  AOI22_X1 U7078 ( .A1(n5997), .A2(n6248), .B1(n6247), .B2(DATAI_21_), .ZN(
        n5999) );
  AOI22_X1 U7079 ( .A1(n6251), .A2(DATAI_5_), .B1(n6250), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7080 ( .A1(n5999), .A2(n5998), .ZN(U2870) );
  AOI22_X1 U7081 ( .A1(n6000), .A2(n6248), .B1(n6247), .B2(DATAI_20_), .ZN(
        n6002) );
  AOI22_X1 U7082 ( .A1(n6251), .A2(DATAI_4_), .B1(n6250), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7083 ( .A1(n6002), .A2(n6001), .ZN(U2871) );
  AOI22_X1 U7084 ( .A1(n6003), .A2(n6248), .B1(n6247), .B2(DATAI_19_), .ZN(
        n6005) );
  AOI22_X1 U7085 ( .A1(n6251), .A2(DATAI_3_), .B1(n6250), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U7086 ( .A1(n6005), .A2(n6004), .ZN(U2872) );
  AOI22_X1 U7087 ( .A1(n6376), .A2(REIP_REG_26__SCAN_IN), .B1(n6330), .B2(
        PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6009) );
  AOI22_X1 U7088 ( .A1(n6007), .A2(n6319), .B1(n6332), .B2(n6006), .ZN(n6008)
         );
  OAI211_X1 U7089 ( .C1(n6324), .C2(n6010), .A(n6009), .B(n6008), .ZN(U2960)
         );
  AOI22_X1 U7090 ( .A1(n6376), .A2(REIP_REG_18__SCAN_IN), .B1(n6330), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6013) );
  AOI22_X1 U7091 ( .A1(n6011), .A2(n6332), .B1(n6319), .B2(n6241), .ZN(n6012)
         );
  OAI211_X1 U7092 ( .C1(n6324), .C2(n6077), .A(n6013), .B(n6012), .ZN(U2968)
         );
  INV_X1 U7093 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6111) );
  INV_X1 U7094 ( .A(n6118), .ZN(n6014) );
  AOI222_X1 U7095 ( .A1(n6015), .A2(n6332), .B1(n6014), .B2(n6310), .C1(n6319), 
        .C2(n6114), .ZN(n6018) );
  INV_X1 U7096 ( .A(n6016), .ZN(n6017) );
  OAI211_X1 U7097 ( .C1(n6111), .C2(n6314), .A(n6018), .B(n6017), .ZN(U2973)
         );
  OAI22_X1 U7098 ( .A1(n5605), .A2(n6338), .B1(n6019), .B2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6020) );
  INV_X1 U7099 ( .A(n6020), .ZN(n6025) );
  INV_X1 U7100 ( .A(n6021), .ZN(n6023) );
  AOI22_X1 U7101 ( .A1(n6023), .A2(n6383), .B1(n6382), .B2(n6022), .ZN(n6024)
         );
  OAI211_X1 U7102 ( .C1(n6027), .C2(n6026), .A(n6025), .B(n6024), .ZN(U2993)
         );
  AOI22_X1 U7103 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n6028), .B1(n6376), .B2(REIP_REG_19__SCAN_IN), .ZN(n6032) );
  AOI22_X1 U7104 ( .A1(n6030), .A2(n6383), .B1(n6382), .B2(n6029), .ZN(n6031)
         );
  OAI211_X1 U7105 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n6033), .A(n6032), .B(n6031), .ZN(U2999) );
  AOI21_X1 U7106 ( .B1(n6045), .B2(n6369), .A(n6034), .ZN(n6051) );
  AOI211_X1 U7107 ( .C1(n3989), .C2(n6042), .A(n6046), .B(n6045), .ZN(n6039)
         );
  OAI22_X1 U7108 ( .A1(n6036), .A2(n6035), .B1(n6107), .B2(n6339), .ZN(n6037)
         );
  AOI21_X1 U7109 ( .B1(n6039), .B2(n6038), .A(n6037), .ZN(n6041) );
  NAND2_X1 U7110 ( .A1(n6376), .A2(REIP_REG_16__SCAN_IN), .ZN(n6040) );
  OAI211_X1 U7111 ( .C1(n6051), .C2(n6042), .A(n6041), .B(n6040), .ZN(U3002)
         );
  AOI21_X1 U7112 ( .B1(n6044), .B2(n6382), .A(n6043), .ZN(n6050) );
  NOR2_X1 U7113 ( .A1(n6046), .A2(n6045), .ZN(n6047) );
  AOI22_X1 U7114 ( .A1(n6048), .A2(n6383), .B1(n3989), .B2(n6047), .ZN(n6049)
         );
  OAI211_X1 U7115 ( .C1(n6051), .C2(n3989), .A(n6050), .B(n6049), .ZN(U3003)
         );
  INV_X1 U7116 ( .A(n6186), .ZN(n6055) );
  INV_X1 U7117 ( .A(n4417), .ZN(n6054) );
  NAND4_X1 U7118 ( .A1(n6055), .A2(n6054), .A3(n6053), .A4(n6052), .ZN(n6056)
         );
  OAI21_X1 U7119 ( .B1(n6058), .B2(n6057), .A(n6056), .ZN(U3455) );
  AOI21_X1 U7120 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6569), .A(n6564), .ZN(n6060) );
  INV_X1 U7121 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6778) );
  AOI21_X1 U7122 ( .B1(n6060), .B2(n6778), .A(n6836), .ZN(U2789) );
  INV_X2 U7123 ( .A(n6836), .ZN(n6835) );
  NOR2_X1 U7124 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6061) );
  OAI21_X1 U7125 ( .B1(n6061), .B2(D_C_N_REG_SCAN_IN), .A(n6835), .ZN(n6059)
         );
  OAI21_X1 U7126 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6835), .A(n6059), .ZN(
        U2791) );
  NOR2_X1 U7127 ( .A1(n6836), .A2(n6060), .ZN(n6618) );
  OAI21_X1 U7128 ( .B1(BS16_N), .B2(n6061), .A(n6618), .ZN(n6616) );
  OAI21_X1 U7129 ( .B1(n6618), .B2(n6822), .A(n6616), .ZN(U2792) );
  OAI21_X1 U7130 ( .B1(n6062), .B2(n6802), .A(n6297), .ZN(U2793) );
  NOR4_X1 U7131 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n6066) );
  NOR4_X1 U7132 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n6065) );
  NOR4_X1 U7133 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6064) );
  NOR4_X1 U7134 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6063) );
  NAND4_X1 U7135 ( .A1(n6066), .A2(n6065), .A3(n6064), .A4(n6063), .ZN(n6072)
         );
  NOR4_X1 U7136 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n6070) );
  AOI211_X1 U7137 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_2__SCAN_IN), .B(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n6069) );
  NOR4_X1 U7138 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n6068) );
  NOR4_X1 U7139 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n6067) );
  NAND4_X1 U7140 ( .A1(n6070), .A2(n6069), .A3(n6068), .A4(n6067), .ZN(n6071)
         );
  NOR2_X1 U7141 ( .A1(n6072), .A2(n6071), .ZN(n6629) );
  INV_X1 U7142 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6820) );
  NOR3_X1 U7143 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6074) );
  OAI21_X1 U7144 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6074), .A(n6629), .ZN(n6073)
         );
  OAI21_X1 U7145 ( .B1(n6629), .B2(n6820), .A(n6073), .ZN(U2794) );
  INV_X1 U7146 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6625) );
  INV_X1 U7147 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6617) );
  AOI21_X1 U7148 ( .B1(n6625), .B2(n6617), .A(n6074), .ZN(n6075) );
  INV_X1 U7149 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6814) );
  INV_X1 U7150 ( .A(n6629), .ZN(n6627) );
  AOI22_X1 U7151 ( .A1(n6629), .A2(n6075), .B1(n6814), .B2(n6627), .ZN(U2795)
         );
  INV_X1 U7152 ( .A(n6179), .ZN(n6190) );
  AOI22_X1 U7153 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6220), .B1(
        REIP_REG_18__SCAN_IN), .B2(n6092), .ZN(n6076) );
  OAI21_X1 U7154 ( .B1(n6077), .B2(n6206), .A(n6076), .ZN(n6078) );
  AOI211_X1 U7155 ( .C1(n6218), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6190), 
        .B(n6078), .ZN(n6082) );
  NOR2_X1 U7156 ( .A1(n6079), .A2(n6200), .ZN(n6080) );
  AOI21_X1 U7157 ( .B1(n6241), .B2(n6145), .A(n6080), .ZN(n6081) );
  OAI211_X1 U7158 ( .C1(REIP_REG_18__SCAN_IN), .C2(n6083), .A(n6082), .B(n6081), .ZN(U2809) );
  OAI22_X1 U7159 ( .A1(n6216), .A2(n6085), .B1(n6084), .B2(n6205), .ZN(n6086)
         );
  AOI211_X1 U7160 ( .C1(n6225), .C2(n6087), .A(n6190), .B(n6086), .ZN(n6094)
         );
  INV_X1 U7161 ( .A(n6088), .ZN(n6244) );
  INV_X1 U7162 ( .A(n6104), .ZN(n6090) );
  NAND2_X1 U7163 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n6089) );
  INV_X1 U7164 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6597) );
  OAI21_X1 U7165 ( .B1(n6090), .B2(n6089), .A(n6597), .ZN(n6091) );
  AOI22_X1 U7166 ( .A1(n6244), .A2(n6145), .B1(n6092), .B2(n6091), .ZN(n6093)
         );
  OAI211_X1 U7167 ( .C1(n6200), .C2(n6095), .A(n6094), .B(n6093), .ZN(U2810)
         );
  INV_X1 U7168 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6595) );
  AOI21_X1 U7169 ( .B1(n6097), .B2(n6096), .A(n6595), .ZN(n6102) );
  NAND2_X1 U7170 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6100)
         );
  AOI22_X1 U7171 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6220), .B1(n6098), .B2(n6225), .ZN(n6099) );
  NAND3_X1 U7172 ( .A1(n6100), .A2(n6179), .A3(n6099), .ZN(n6101) );
  OR2_X1 U7173 ( .A1(n6102), .A2(n6101), .ZN(n6103) );
  AOI21_X1 U7174 ( .B1(n6249), .B2(n6145), .A(n6103), .ZN(n6106) );
  NAND3_X1 U7175 ( .A1(n6104), .A2(REIP_REG_15__SCAN_IN), .A3(n6595), .ZN(
        n6105) );
  OAI211_X1 U7176 ( .C1(n6107), .C2(n6200), .A(n6106), .B(n6105), .ZN(U2811)
         );
  NOR3_X1 U7177 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6120), .A3(n6108), .ZN(n6113) );
  AOI22_X1 U7178 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6220), .B1(n6177), .B2(n6109), .ZN(n6110) );
  OAI211_X1 U7179 ( .C1(n6205), .C2(n6111), .A(n6179), .B(n6110), .ZN(n6112)
         );
  AOI211_X1 U7180 ( .C1(n6114), .C2(n6145), .A(n6113), .B(n6112), .ZN(n6117)
         );
  OAI21_X1 U7181 ( .B1(n6115), .B2(n6121), .A(REIP_REG_13__SCAN_IN), .ZN(n6116) );
  OAI211_X1 U7182 ( .C1(n6206), .C2(n6118), .A(n6117), .B(n6116), .ZN(U2814)
         );
  AOI22_X1 U7183 ( .A1(EBX_REG_11__SCAN_IN), .A2(n6220), .B1(n6177), .B2(n6234), .ZN(n6126) );
  NOR2_X1 U7184 ( .A1(n6120), .A2(n6119), .ZN(n6122) );
  MUX2_X1 U7185 ( .A(n6122), .B(n6121), .S(REIP_REG_11__SCAN_IN), .Z(n6123) );
  AOI211_X1 U7186 ( .C1(n6218), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6190), 
        .B(n6123), .ZN(n6125) );
  INV_X1 U7187 ( .A(n6237), .ZN(n6294) );
  AOI22_X1 U7188 ( .A1(n6294), .A2(n6145), .B1(n6225), .B2(n6293), .ZN(n6124)
         );
  NAND3_X1 U7189 ( .A1(n6126), .A2(n6125), .A3(n6124), .ZN(U2816) );
  INV_X1 U7190 ( .A(n6127), .ZN(n6350) );
  AOI22_X1 U7191 ( .A1(n6177), .A2(n6350), .B1(REIP_REG_9__SCAN_IN), .B2(n6142), .ZN(n6136) );
  OAI21_X1 U7192 ( .B1(n6205), .B2(n6128), .A(n6179), .ZN(n6129) );
  AOI211_X1 U7193 ( .C1(EBX_REG_9__SCAN_IN), .C2(n6220), .A(n6130), .B(n6129), 
        .ZN(n6135) );
  INV_X1 U7194 ( .A(n6131), .ZN(n6133) );
  AOI22_X1 U7195 ( .A1(n6133), .A2(n6145), .B1(n6225), .B2(n6132), .ZN(n6134)
         );
  NAND3_X1 U7196 ( .A1(n6136), .A2(n6135), .A3(n6134), .ZN(U2818) );
  OAI22_X1 U7197 ( .A1(n6138), .A2(n6216), .B1(n6200), .B2(n6137), .ZN(n6139)
         );
  INV_X1 U7198 ( .A(n6139), .ZN(n6149) );
  NAND2_X1 U7199 ( .A1(n6582), .A2(n6140), .ZN(n6141) );
  AOI22_X1 U7200 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n6218), .B1(n6142), 
        .B2(n6141), .ZN(n6148) );
  INV_X1 U7201 ( .A(n6143), .ZN(n6144) );
  AOI22_X1 U7202 ( .A1(n6146), .A2(n6145), .B1(n6225), .B2(n6144), .ZN(n6147)
         );
  NAND4_X1 U7203 ( .A1(n6149), .A2(n6148), .A3(n6147), .A4(n6179), .ZN(U2819)
         );
  NOR3_X1 U7204 ( .A1(n6210), .A2(REIP_REG_7__SCAN_IN), .A3(n6150), .ZN(n6151)
         );
  AOI211_X1 U7205 ( .C1(n6218), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6190), 
        .B(n6151), .ZN(n6161) );
  OAI21_X1 U7206 ( .B1(n6154), .B2(n6153), .A(n6152), .ZN(n6183) );
  NAND3_X1 U7207 ( .A1(n6156), .A2(n6578), .A3(n6155), .ZN(n6163) );
  AOI21_X1 U7208 ( .B1(n6183), .B2(n6163), .A(n6580), .ZN(n6159) );
  OAI22_X1 U7209 ( .A1(n6157), .A2(n6167), .B1(n6299), .B2(n6206), .ZN(n6158)
         );
  AOI211_X1 U7210 ( .C1(EBX_REG_7__SCAN_IN), .C2(n6220), .A(n6159), .B(n6158), 
        .ZN(n6160) );
  OAI211_X1 U7211 ( .C1(n6200), .C2(n6162), .A(n6161), .B(n6160), .ZN(U2820)
         );
  OAI211_X1 U7212 ( .C1(n6205), .C2(n6164), .A(n6179), .B(n6163), .ZN(n6170)
         );
  INV_X1 U7213 ( .A(n6165), .ZN(n6166) );
  OAI22_X1 U7214 ( .A1(n6168), .A2(n6167), .B1(n6166), .B2(n6206), .ZN(n6169)
         );
  AOI211_X1 U7215 ( .C1(n6177), .C2(n6171), .A(n6170), .B(n6169), .ZN(n6173)
         );
  NAND2_X1 U7216 ( .A1(EBX_REG_6__SCAN_IN), .A2(n6220), .ZN(n6172) );
  OAI211_X1 U7217 ( .C1(n6183), .C2(n6578), .A(n6173), .B(n6172), .ZN(U2821)
         );
  OR2_X1 U7218 ( .A1(n6210), .A2(n6174), .ZN(n6192) );
  INV_X1 U7219 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6576) );
  OAI21_X1 U7220 ( .B1(n6192), .B2(n6188), .A(n6576), .ZN(n6175) );
  INV_X1 U7221 ( .A(n6175), .ZN(n6182) );
  AOI22_X1 U7222 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6220), .B1(n6177), .B2(n6176), 
        .ZN(n6178) );
  NAND2_X1 U7223 ( .A1(n6179), .A2(n6178), .ZN(n6180) );
  AOI21_X1 U7224 ( .B1(n6218), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n6180), 
        .ZN(n6181) );
  OAI21_X1 U7225 ( .B1(n6183), .B2(n6182), .A(n6181), .ZN(n6184) );
  AOI21_X1 U7226 ( .B1(n6309), .B2(n6209), .A(n6184), .ZN(n6185) );
  OAI21_X1 U7227 ( .B1(n6306), .B2(n6206), .A(n6185), .ZN(U2822) );
  OAI22_X1 U7228 ( .A1(n6188), .A2(n6187), .B1(n6186), .B2(n6202), .ZN(n6189)
         );
  AOI211_X1 U7229 ( .C1(n6218), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6190), 
        .B(n6189), .ZN(n6198) );
  OAI22_X1 U7230 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6192), .B1(n6216), .B2(n6191), .ZN(n6196) );
  OAI22_X1 U7231 ( .A1(n6194), .A2(n6227), .B1(n6193), .B2(n6206), .ZN(n6195)
         );
  NOR2_X1 U7232 ( .A1(n6196), .A2(n6195), .ZN(n6197) );
  OAI211_X1 U7233 ( .C1(n6200), .C2(n6199), .A(n6198), .B(n6197), .ZN(U2823)
         );
  OAI22_X1 U7234 ( .A1(n6203), .A2(n6202), .B1(n6201), .B2(n6200), .ZN(n6208)
         );
  OAI22_X1 U7235 ( .A1(n6323), .A2(n6206), .B1(n6205), .B2(n6204), .ZN(n6207)
         );
  AOI211_X1 U7236 ( .C1(n6320), .C2(n6209), .A(n6208), .B(n6207), .ZN(n6214)
         );
  NOR2_X1 U7237 ( .A1(n6210), .A2(n6625), .ZN(n6212) );
  OAI21_X1 U7238 ( .B1(REIP_REG_2__SCAN_IN), .B2(n6212), .A(n6211), .ZN(n6213)
         );
  OAI211_X1 U7239 ( .C1(n6216), .C2(n6215), .A(n6214), .B(n6213), .ZN(U2825)
         );
  AOI22_X1 U7240 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n6218), .B1(n6217), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n6231) );
  NAND2_X1 U7241 ( .A1(n4427), .A2(n6219), .ZN(n6223) );
  NAND2_X1 U7242 ( .A1(n6220), .A2(EBX_REG_1__SCAN_IN), .ZN(n6221) );
  NAND3_X1 U7243 ( .A1(n6223), .A2(n6222), .A3(n6221), .ZN(n6224) );
  AOI21_X1 U7244 ( .B1(n6225), .B2(n4550), .A(n6224), .ZN(n6226) );
  OAI21_X1 U7245 ( .B1(n6228), .B2(n6227), .A(n6226), .ZN(n6229) );
  INV_X1 U7246 ( .A(n6229), .ZN(n6230) );
  OAI211_X1 U7247 ( .C1(n6233), .C2(n6232), .A(n6231), .B(n6230), .ZN(U2826)
         );
  INV_X1 U7248 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6240) );
  INV_X1 U7249 ( .A(n6234), .ZN(n6235) );
  OAI22_X1 U7250 ( .A1(n6237), .A2(n6236), .B1(n5557), .B2(n6235), .ZN(n6238)
         );
  INV_X1 U7251 ( .A(n6238), .ZN(n6239) );
  OAI21_X1 U7252 ( .B1(n6240), .B2(n5567), .A(n6239), .ZN(U2848) );
  AOI22_X1 U7253 ( .A1(n6241), .A2(n6248), .B1(n6247), .B2(DATAI_18_), .ZN(
        n6243) );
  AOI22_X1 U7254 ( .A1(n6251), .A2(DATAI_2_), .B1(n6250), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U7255 ( .A1(n6243), .A2(n6242), .ZN(U2873) );
  AOI22_X1 U7256 ( .A1(n6244), .A2(n6248), .B1(n6247), .B2(DATAI_17_), .ZN(
        n6246) );
  AOI22_X1 U7257 ( .A1(n6251), .A2(DATAI_1_), .B1(n6250), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7258 ( .A1(n6246), .A2(n6245), .ZN(U2874) );
  AOI22_X1 U7259 ( .A1(n6249), .A2(n6248), .B1(n6247), .B2(DATAI_16_), .ZN(
        n6253) );
  AOI22_X1 U7260 ( .A1(n6251), .A2(DATAI_0_), .B1(n6250), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U7261 ( .A1(n6253), .A2(n6252), .ZN(U2875) );
  AOI22_X1 U7262 ( .A1(n6284), .A2(LWORD_REG_15__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6254) );
  OAI21_X1 U7263 ( .B1(n4400), .B2(n6286), .A(n6254), .ZN(U2908) );
  INV_X1 U7264 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6256) );
  AOI22_X1 U7265 ( .A1(n6284), .A2(LWORD_REG_14__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6255) );
  OAI21_X1 U7266 ( .B1(n6256), .B2(n6286), .A(n6255), .ZN(U2909) );
  INV_X1 U7267 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6258) );
  AOI22_X1 U7268 ( .A1(n6284), .A2(LWORD_REG_13__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6257) );
  OAI21_X1 U7269 ( .B1(n6258), .B2(n6286), .A(n6257), .ZN(U2910) );
  INV_X1 U7270 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6260) );
  AOI22_X1 U7271 ( .A1(n6284), .A2(LWORD_REG_12__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6259) );
  OAI21_X1 U7272 ( .B1(n6260), .B2(n6286), .A(n6259), .ZN(U2911) );
  INV_X1 U7273 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6262) );
  AOI22_X1 U7274 ( .A1(n6284), .A2(LWORD_REG_11__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6261) );
  OAI21_X1 U7275 ( .B1(n6262), .B2(n6286), .A(n6261), .ZN(U2912) );
  AOI22_X1 U7276 ( .A1(n6284), .A2(LWORD_REG_10__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6263) );
  OAI21_X1 U7277 ( .B1(n4402), .B2(n6286), .A(n6263), .ZN(U2913) );
  INV_X1 U7278 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6265) );
  AOI22_X1 U7279 ( .A1(n6284), .A2(LWORD_REG_9__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6264) );
  OAI21_X1 U7280 ( .B1(n6265), .B2(n6286), .A(n6264), .ZN(U2914) );
  INV_X1 U7281 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6267) );
  AOI22_X1 U7282 ( .A1(n6284), .A2(LWORD_REG_8__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6266) );
  OAI21_X1 U7283 ( .B1(n6267), .B2(n6286), .A(n6266), .ZN(U2915) );
  INV_X1 U7284 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6269) );
  AOI22_X1 U7285 ( .A1(n6284), .A2(LWORD_REG_7__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6268) );
  OAI21_X1 U7286 ( .B1(n6269), .B2(n6286), .A(n6268), .ZN(U2916) );
  INV_X1 U7287 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6271) );
  AOI22_X1 U7288 ( .A1(n6284), .A2(LWORD_REG_6__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6270) );
  OAI21_X1 U7289 ( .B1(n6271), .B2(n6286), .A(n6270), .ZN(U2917) );
  AOI22_X1 U7290 ( .A1(n6284), .A2(LWORD_REG_5__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6272) );
  OAI21_X1 U7291 ( .B1(n6273), .B2(n6286), .A(n6272), .ZN(U2918) );
  AOI22_X1 U7292 ( .A1(n6284), .A2(LWORD_REG_4__SCAN_IN), .B1(n6274), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6275) );
  OAI21_X1 U7293 ( .B1(n6276), .B2(n6286), .A(n6275), .ZN(U2919) );
  AOI22_X1 U7294 ( .A1(n6284), .A2(LWORD_REG_3__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6277) );
  OAI21_X1 U7295 ( .B1(n6278), .B2(n6286), .A(n6277), .ZN(U2920) );
  AOI22_X1 U7296 ( .A1(n6284), .A2(LWORD_REG_2__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6279) );
  OAI21_X1 U7297 ( .B1(n6280), .B2(n6286), .A(n6279), .ZN(U2921) );
  AOI22_X1 U7298 ( .A1(n6284), .A2(LWORD_REG_1__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6281) );
  OAI21_X1 U7299 ( .B1(n6282), .B2(n6286), .A(n6281), .ZN(U2922) );
  AOI22_X1 U7300 ( .A1(n6284), .A2(LWORD_REG_0__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6285) );
  OAI21_X1 U7301 ( .B1(n6287), .B2(n6286), .A(n6285), .ZN(U2923) );
  AOI22_X1 U7302 ( .A1(n6289), .A2(UWORD_REG_10__SCAN_IN), .B1(n6288), .B2(
        DATAI_10_), .ZN(n6290) );
  OAI21_X1 U7303 ( .B1(n6292), .B2(n6291), .A(n6290), .ZN(U2934) );
  AOI22_X1 U7304 ( .A1(n6376), .A2(REIP_REG_11__SCAN_IN), .B1(n6330), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6296) );
  AOI22_X1 U7305 ( .A1(n6294), .A2(n6319), .B1(n6310), .B2(n6293), .ZN(n6295)
         );
  OAI211_X1 U7306 ( .C1(n6298), .C2(n6297), .A(n6296), .B(n6295), .ZN(U2975)
         );
  INV_X1 U7307 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6305) );
  INV_X1 U7308 ( .A(n6299), .ZN(n6302) );
  AOI222_X1 U7309 ( .A1(n6302), .A2(n6310), .B1(n6319), .B2(n6301), .C1(n6332), 
        .C2(n6300), .ZN(n6304) );
  OAI211_X1 U7310 ( .C1(n6305), .C2(n6314), .A(n6304), .B(n6303), .ZN(U2979)
         );
  INV_X1 U7311 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6315) );
  INV_X1 U7312 ( .A(n6306), .ZN(n6311) );
  INV_X1 U7313 ( .A(n6307), .ZN(n6308) );
  AOI222_X1 U7314 ( .A1(n6311), .A2(n6310), .B1(n6319), .B2(n6309), .C1(n6332), 
        .C2(n6308), .ZN(n6313) );
  OAI211_X1 U7315 ( .C1(n6315), .C2(n6314), .A(n6313), .B(n6312), .ZN(U2981)
         );
  AOI22_X1 U7316 ( .A1(n6376), .A2(REIP_REG_2__SCAN_IN), .B1(n6330), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6322) );
  XNOR2_X1 U7317 ( .A(n6316), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6318)
         );
  XNOR2_X1 U7318 ( .A(n6318), .B(n6317), .ZN(n6364) );
  AOI22_X1 U7319 ( .A1(n6320), .A2(n6319), .B1(n6332), .B2(n6364), .ZN(n6321)
         );
  OAI211_X1 U7320 ( .C1(n6324), .C2(n6323), .A(n6322), .B(n6321), .ZN(U2984)
         );
  INV_X1 U7321 ( .A(n6325), .ZN(n6328) );
  INV_X1 U7322 ( .A(n6326), .ZN(n6327) );
  AOI21_X1 U7323 ( .B1(n6328), .B2(n6371), .A(n6327), .ZN(n6384) );
  OR2_X1 U7324 ( .A1(n6330), .A2(n6329), .ZN(n6331) );
  AOI22_X1 U7325 ( .A1(n6384), .A2(n6332), .B1(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6331), .ZN(n6334) );
  NAND2_X1 U7326 ( .A1(n6376), .A2(REIP_REG_0__SCAN_IN), .ZN(n6333) );
  OAI211_X1 U7327 ( .C1(n6336), .C2(n6335), .A(n6334), .B(n6333), .ZN(U2986)
         );
  AOI21_X1 U7328 ( .B1(n6344), .B2(n6369), .A(n6337), .ZN(n6356) );
  OAI22_X1 U7329 ( .A1(n6340), .A2(n6339), .B1(n6585), .B2(n6338), .ZN(n6341)
         );
  AOI21_X1 U7330 ( .B1(n6342), .B2(n6383), .A(n6341), .ZN(n6347) );
  NOR2_X1 U7331 ( .A1(n6344), .A2(n6343), .ZN(n6351) );
  OAI211_X1 U7332 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6351), .B(n6345), .ZN(n6346) );
  OAI211_X1 U7333 ( .C1(n6356), .C2(n6348), .A(n6347), .B(n6346), .ZN(U3008)
         );
  AOI21_X1 U7334 ( .B1(n6350), .B2(n6382), .A(n6349), .ZN(n6354) );
  AOI22_X1 U7335 ( .A1(n6352), .A2(n6383), .B1(n6351), .B2(n6355), .ZN(n6353)
         );
  OAI211_X1 U7336 ( .C1(n6356), .C2(n6355), .A(n6354), .B(n6353), .ZN(U3009)
         );
  NAND2_X1 U7337 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6357), .ZN(n6367)
         );
  AOI22_X1 U7338 ( .A1(n6382), .A2(n6358), .B1(n6376), .B2(REIP_REG_2__SCAN_IN), .ZN(n6362) );
  NAND3_X1 U7339 ( .A1(n6372), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(n6359), 
        .ZN(n6360) );
  NAND3_X1 U7340 ( .A1(n6362), .A2(n6361), .A3(n6360), .ZN(n6363) );
  AOI21_X1 U7341 ( .B1(n6364), .B2(n6383), .A(n6363), .ZN(n6365) );
  OAI221_X1 U7342 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6367), .C1(n4125), .C2(n6366), .A(n6365), .ZN(U3016) );
  NAND2_X1 U7343 ( .A1(n6369), .A2(n6368), .ZN(n6379) );
  AOI21_X1 U7344 ( .B1(n6372), .B2(n6371), .A(n6370), .ZN(n6386) );
  INV_X1 U7345 ( .A(n6373), .ZN(n6375) );
  AOI222_X1 U7346 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6376), .B1(n6383), .B2(
        n6375), .C1(n6374), .C2(n6382), .ZN(n6377) );
  OAI221_X1 U7347 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n6379), .C1(n6378), .C2(n6386), .A(n6377), .ZN(U3017) );
  INV_X1 U7348 ( .A(n6380), .ZN(n6381) );
  AOI22_X1 U7349 ( .A1(n6384), .A2(n6383), .B1(n6382), .B2(n6381), .ZN(n6391)
         );
  INV_X1 U7350 ( .A(n6385), .ZN(n6389) );
  INV_X1 U7351 ( .A(n6386), .ZN(n6388) );
  OAI22_X1 U7352 ( .A1(n6389), .A2(n6388), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6387), .ZN(n6390) );
  OAI211_X1 U7353 ( .C1(n6392), .C2(n6338), .A(n6391), .B(n6390), .ZN(U3018)
         );
  NOR2_X1 U7354 ( .A1(n6394), .A2(n6393), .ZN(U3019) );
  INV_X1 U7355 ( .A(n6395), .ZN(n6400) );
  NAND3_X1 U7356 ( .A1(n6397), .A2(n6396), .A3(n6517), .ZN(n6398) );
  OAI21_X1 U7357 ( .B1(n6400), .B2(n6399), .A(n6398), .ZN(n6443) );
  NAND2_X1 U7358 ( .A1(n6401), .A2(n3368), .ZN(n6409) );
  INV_X1 U7359 ( .A(n6409), .ZN(n6442) );
  AOI22_X1 U7360 ( .A1(n6403), .A2(n6443), .B1(n6402), .B2(n6442), .ZN(n6414)
         );
  OAI21_X1 U7361 ( .B1(n6445), .B2(n6404), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6406) );
  AND2_X1 U7362 ( .A1(n6406), .A2(n6405), .ZN(n6407) );
  AOI22_X1 U7363 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6409), .B1(n6408), .B2(
        n6407), .ZN(n6411) );
  NAND3_X1 U7364 ( .A1(n6517), .A2(n6411), .A3(n6410), .ZN(n6446) );
  AOI22_X1 U7365 ( .A1(n6446), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6412), 
        .B2(n6445), .ZN(n6413) );
  OAI211_X1 U7366 ( .C1(n6415), .C2(n6460), .A(n6414), .B(n6413), .ZN(U3068)
         );
  AOI22_X1 U7367 ( .A1(n6463), .A2(n6443), .B1(n6461), .B2(n6442), .ZN(n6418)
         );
  AOI22_X1 U7368 ( .A1(n6446), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6445), 
        .B2(n6416), .ZN(n6417) );
  OAI211_X1 U7369 ( .C1(n6419), .C2(n6460), .A(n6418), .B(n6417), .ZN(U3069)
         );
  AOI22_X1 U7370 ( .A1(n6469), .A2(n6443), .B1(n6467), .B2(n6442), .ZN(n6422)
         );
  AOI22_X1 U7371 ( .A1(n6446), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6445), 
        .B2(n6420), .ZN(n6421) );
  OAI211_X1 U7372 ( .C1(n6423), .C2(n6460), .A(n6422), .B(n6421), .ZN(U3070)
         );
  AOI22_X1 U7373 ( .A1(n6475), .A2(n6443), .B1(n6473), .B2(n6442), .ZN(n6426)
         );
  AOI22_X1 U7374 ( .A1(n6446), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6445), 
        .B2(n6424), .ZN(n6425) );
  OAI211_X1 U7375 ( .C1(n6427), .C2(n6460), .A(n6426), .B(n6425), .ZN(U3071)
         );
  AOI22_X1 U7376 ( .A1(n6481), .A2(n6443), .B1(n6479), .B2(n6442), .ZN(n6430)
         );
  AOI22_X1 U7377 ( .A1(n6446), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6445), 
        .B2(n6428), .ZN(n6429) );
  OAI211_X1 U7378 ( .C1(n6431), .C2(n6460), .A(n6430), .B(n6429), .ZN(U3072)
         );
  AOI22_X1 U7379 ( .A1(n6487), .A2(n6443), .B1(n6485), .B2(n6442), .ZN(n6434)
         );
  AOI22_X1 U7380 ( .A1(n6446), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6445), 
        .B2(n6432), .ZN(n6433) );
  OAI211_X1 U7381 ( .C1(n6435), .C2(n6460), .A(n6434), .B(n6433), .ZN(U3073)
         );
  AOI22_X1 U7382 ( .A1(n6437), .A2(n6443), .B1(n6436), .B2(n6442), .ZN(n6440)
         );
  AOI22_X1 U7383 ( .A1(n6446), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6445), 
        .B2(n6438), .ZN(n6439) );
  OAI211_X1 U7384 ( .C1(n6441), .C2(n6460), .A(n6440), .B(n6439), .ZN(U3074)
         );
  AOI22_X1 U7385 ( .A1(n6496), .A2(n6443), .B1(n6492), .B2(n6442), .ZN(n6448)
         );
  AOI22_X1 U7386 ( .A1(n6446), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6445), 
        .B2(n6444), .ZN(n6447) );
  OAI211_X1 U7387 ( .C1(n6449), .C2(n6460), .A(n6448), .B(n6447), .ZN(U3075)
         );
  INV_X1 U7388 ( .A(n6450), .ZN(n6455) );
  INV_X1 U7389 ( .A(n6451), .ZN(n6454) );
  AOI22_X1 U7390 ( .A1(n6455), .A2(n6462), .B1(n6461), .B2(n6454), .ZN(n6453)
         );
  AOI22_X1 U7391 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6457), .B1(n6463), 
        .B2(n6456), .ZN(n6452) );
  OAI211_X1 U7392 ( .C1(n6466), .C2(n6460), .A(n6453), .B(n6452), .ZN(U3077)
         );
  AOI22_X1 U7393 ( .A1(n6455), .A2(n6486), .B1(n6485), .B2(n6454), .ZN(n6459)
         );
  AOI22_X1 U7394 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6457), .B1(n6487), 
        .B2(n6456), .ZN(n6458) );
  OAI211_X1 U7395 ( .C1(n6490), .C2(n6460), .A(n6459), .B(n6458), .ZN(U3081)
         );
  AOI22_X1 U7396 ( .A1(n6494), .A2(n6462), .B1(n6461), .B2(n6491), .ZN(n6465)
         );
  AOI22_X1 U7397 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6497), .B1(n6463), 
        .B2(n6495), .ZN(n6464) );
  OAI211_X1 U7398 ( .C1(n6466), .C2(n6500), .A(n6465), .B(n6464), .ZN(U3109)
         );
  AOI22_X1 U7399 ( .A1(n6494), .A2(n6468), .B1(n6467), .B2(n6491), .ZN(n6471)
         );
  AOI22_X1 U7400 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6497), .B1(n6469), 
        .B2(n6495), .ZN(n6470) );
  OAI211_X1 U7401 ( .C1(n6472), .C2(n6500), .A(n6471), .B(n6470), .ZN(U3110)
         );
  AOI22_X1 U7402 ( .A1(n6494), .A2(n6474), .B1(n6473), .B2(n6491), .ZN(n6477)
         );
  AOI22_X1 U7403 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6497), .B1(n6475), 
        .B2(n6495), .ZN(n6476) );
  OAI211_X1 U7404 ( .C1(n6478), .C2(n6500), .A(n6477), .B(n6476), .ZN(U3111)
         );
  AOI22_X1 U7405 ( .A1(n6494), .A2(n6480), .B1(n6479), .B2(n6491), .ZN(n6483)
         );
  AOI22_X1 U7406 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6497), .B1(n6481), 
        .B2(n6495), .ZN(n6482) );
  OAI211_X1 U7407 ( .C1(n6484), .C2(n6500), .A(n6483), .B(n6482), .ZN(U3112)
         );
  AOI22_X1 U7408 ( .A1(n6494), .A2(n6486), .B1(n6485), .B2(n6491), .ZN(n6489)
         );
  AOI22_X1 U7409 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6497), .B1(n6487), 
        .B2(n6495), .ZN(n6488) );
  OAI211_X1 U7410 ( .C1(n6490), .C2(n6500), .A(n6489), .B(n6488), .ZN(U3113)
         );
  AOI22_X1 U7411 ( .A1(n6494), .A2(n6493), .B1(n6492), .B2(n6491), .ZN(n6499)
         );
  AOI22_X1 U7412 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6497), .B1(n6496), 
        .B2(n6495), .ZN(n6498) );
  OAI211_X1 U7413 ( .C1(n6501), .C2(n6500), .A(n6499), .B(n6498), .ZN(U3115)
         );
  INV_X1 U7414 ( .A(n6502), .ZN(n6508) );
  OAI21_X1 U7415 ( .B1(n6504), .B2(n6503), .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .ZN(n6505) );
  NOR2_X1 U7416 ( .A1(n6506), .A2(n6505), .ZN(n6509) );
  OAI22_X1 U7417 ( .A1(n6508), .A2(n6507), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6509), .ZN(n6511) );
  NAND2_X1 U7418 ( .A1(n6509), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6510) );
  OAI211_X1 U7419 ( .C1(n6513), .C2(n6512), .A(n6511), .B(n6510), .ZN(n6515)
         );
  NAND2_X1 U7420 ( .A1(n6513), .A2(n6512), .ZN(n6514) );
  NAND2_X1 U7421 ( .A1(n6515), .A2(n6514), .ZN(n6516) );
  OAI21_X1 U7422 ( .B1(n6518), .B2(n6517), .A(n6516), .ZN(n6520) );
  NAND2_X1 U7423 ( .A1(n6518), .A2(n6517), .ZN(n6519) );
  AOI21_X1 U7424 ( .B1(n6520), .B2(n6519), .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .ZN(n6528) );
  INV_X1 U7425 ( .A(MORE_REG_SCAN_IN), .ZN(n6747) );
  AND2_X1 U7426 ( .A1(n6802), .A2(n6747), .ZN(n6523) );
  OAI211_X1 U7427 ( .C1(n6524), .C2(n6523), .A(n6522), .B(n6521), .ZN(n6525)
         );
  OAI22_X1 U7428 ( .A1(n6538), .A2(n6545), .B1(n6768), .B2(n6529), .ZN(n6533)
         );
  OR2_X1 U7429 ( .A1(n6531), .A2(n6530), .ZN(n6532) );
  AOI21_X1 U7430 ( .B1(READY_N), .B2(n6633), .A(n6619), .ZN(n6543) );
  AOI211_X1 U7431 ( .C1(n6535), .C2(n6534), .A(STATE2_REG_0__SCAN_IN), .B(
        n6619), .ZN(n6536) );
  AOI211_X1 U7432 ( .C1(n6539), .C2(n6538), .A(n6537), .B(n6536), .ZN(n6540)
         );
  OAI221_X1 U7433 ( .B1(n6636), .B2(n6543), .C1(n6636), .C2(n6541), .A(n6540), 
        .ZN(U3148) );
  NOR2_X1 U7434 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6551) );
  NOR3_X1 U7435 ( .A1(n6551), .A2(n6543), .A3(n6542), .ZN(n6547) );
  AOI221_X1 U7436 ( .B1(READY_N), .B2(n6545), .C1(n6544), .C2(n6545), .A(n6619), .ZN(n6546) );
  OR3_X1 U7437 ( .A1(n6548), .A2(n6547), .A3(n6546), .ZN(U3149) );
  OAI211_X1 U7438 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6768), .A(n6620), .B(
        n6635), .ZN(n6550) );
  OAI21_X1 U7439 ( .B1(n6551), .B2(n6550), .A(n6549), .ZN(U3150) );
  AND2_X1 U7440 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6552), .ZN(U3151) );
  AND2_X1 U7441 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6552), .ZN(U3152) );
  AND2_X1 U7442 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6552), .ZN(U3153) );
  AND2_X1 U7443 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6552), .ZN(U3154) );
  AND2_X1 U7444 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6552), .ZN(U3155) );
  AND2_X1 U7445 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6552), .ZN(U3156) );
  AND2_X1 U7446 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6552), .ZN(U3157) );
  AND2_X1 U7447 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6552), .ZN(U3158) );
  AND2_X1 U7448 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6552), .ZN(U3159) );
  AND2_X1 U7449 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6552), .ZN(U3160) );
  AND2_X1 U7450 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6552), .ZN(U3161) );
  AND2_X1 U7451 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6552), .ZN(U3162) );
  AND2_X1 U7452 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6552), .ZN(U3163) );
  AND2_X1 U7453 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6552), .ZN(U3164) );
  AND2_X1 U7454 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6552), .ZN(U3165) );
  AND2_X1 U7455 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6552), .ZN(U3166) );
  AND2_X1 U7456 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6552), .ZN(U3167) );
  AND2_X1 U7457 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6552), .ZN(U3168) );
  AND2_X1 U7458 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6552), .ZN(U3169) );
  AND2_X1 U7459 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6552), .ZN(U3170) );
  AND2_X1 U7460 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6552), .ZN(U3171) );
  AND2_X1 U7461 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6552), .ZN(U3172) );
  AND2_X1 U7462 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6552), .ZN(U3173) );
  AND2_X1 U7463 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6552), .ZN(U3174) );
  AND2_X1 U7464 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6552), .ZN(U3175) );
  AND2_X1 U7465 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6552), .ZN(U3176) );
  AND2_X1 U7466 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6552), .ZN(U3177) );
  AND2_X1 U7467 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6552), .ZN(U3178) );
  AND2_X1 U7468 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6552), .ZN(U3179) );
  AND2_X1 U7469 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6552), .ZN(U3180) );
  INV_X1 U7470 ( .A(n6567), .ZN(n6554) );
  AOI22_X1 U7471 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6568) );
  INV_X1 U7472 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6563) );
  INV_X1 U7473 ( .A(HOLD), .ZN(n6775) );
  NOR2_X1 U7474 ( .A1(n6563), .A2(n6775), .ZN(n6555) );
  INV_X1 U7475 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6562) );
  OAI21_X1 U7476 ( .B1(n6555), .B2(n6562), .A(n6835), .ZN(n6553) );
  OAI211_X1 U7477 ( .C1(NA_N), .C2(n6569), .A(n6564), .B(n6567), .ZN(n6559) );
  OAI211_X1 U7478 ( .C1(n6554), .C2(n6568), .A(n6553), .B(n6559), .ZN(U3181)
         );
  NOR2_X1 U7479 ( .A1(n6564), .A2(n6562), .ZN(n6556) );
  OAI22_X1 U7480 ( .A1(n6556), .A2(n6555), .B1(n6569), .B2(n6775), .ZN(n6557)
         );
  OAI211_X1 U7481 ( .C1(n6563), .C2(n6768), .A(n6558), .B(n6557), .ZN(U3182)
         );
  INV_X1 U7482 ( .A(NA_N), .ZN(n6676) );
  NAND2_X1 U7483 ( .A1(READY_N), .A2(n6676), .ZN(n6561) );
  OAI221_X1 U7484 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(STATE_REG_1__SCAN_IN), 
        .C1(REQUESTPENDING_REG_SCAN_IN), .C2(n6561), .A(n6569), .ZN(n6560) );
  OAI211_X1 U7485 ( .C1(n6564), .C2(HOLD), .A(n6560), .B(n6559), .ZN(n6566) );
  OR4_X1 U7486 ( .A1(n6564), .A2(n6563), .A3(n6562), .A4(n6561), .ZN(n6565) );
  OAI211_X1 U7487 ( .C1(n6568), .C2(n6567), .A(n6566), .B(n6565), .ZN(U3183)
         );
  NOR2_X1 U7488 ( .A1(n6569), .A2(n6835), .ZN(n6609) );
  NAND2_X1 U7489 ( .A1(n6569), .A2(n6836), .ZN(n6611) );
  INV_X1 U7490 ( .A(n6611), .ZN(n6612) );
  AOI22_X1 U7491 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6835), .ZN(n6570) );
  OAI21_X1 U7492 ( .B1(n6625), .B2(n6614), .A(n6570), .ZN(U3184) );
  AOI22_X1 U7493 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6835), .ZN(n6571) );
  OAI21_X1 U7494 ( .B1(n6573), .B2(n6611), .A(n6571), .ZN(U3185) );
  AOI22_X1 U7495 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6835), .ZN(n6572) );
  OAI21_X1 U7496 ( .B1(n6573), .B2(n6614), .A(n6572), .ZN(U3186) );
  AOI22_X1 U7497 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6835), .ZN(n6574) );
  OAI21_X1 U7498 ( .B1(n6576), .B2(n6611), .A(n6574), .ZN(U3187) );
  AOI22_X1 U7499 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6835), .ZN(n6575) );
  OAI21_X1 U7500 ( .B1(n6576), .B2(n6614), .A(n6575), .ZN(U3188) );
  AOI22_X1 U7501 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6835), .ZN(n6577) );
  OAI21_X1 U7502 ( .B1(n6578), .B2(n6614), .A(n6577), .ZN(U3189) );
  AOI22_X1 U7503 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6835), .ZN(n6579) );
  OAI21_X1 U7504 ( .B1(n6580), .B2(n6614), .A(n6579), .ZN(U3190) );
  AOI22_X1 U7505 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6835), .ZN(n6581) );
  OAI21_X1 U7506 ( .B1(n6582), .B2(n6614), .A(n6581), .ZN(U3191) );
  AOI22_X1 U7507 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6835), .ZN(n6583) );
  OAI21_X1 U7508 ( .B1(n6585), .B2(n6611), .A(n6583), .ZN(U3192) );
  AOI22_X1 U7509 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6835), .ZN(n6584) );
  OAI21_X1 U7510 ( .B1(n6585), .B2(n6614), .A(n6584), .ZN(U3193) );
  AOI22_X1 U7511 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6835), .ZN(n6586) );
  OAI21_X1 U7512 ( .B1(n6587), .B2(n6614), .A(n6586), .ZN(U3194) );
  AOI22_X1 U7513 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6835), .ZN(n6588) );
  OAI21_X1 U7514 ( .B1(n6590), .B2(n6611), .A(n6588), .ZN(U3195) );
  AOI22_X1 U7515 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6835), .ZN(n6589) );
  OAI21_X1 U7516 ( .B1(n6590), .B2(n6614), .A(n6589), .ZN(U3196) );
  AOI22_X1 U7517 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6835), .ZN(n6591) );
  OAI21_X1 U7518 ( .B1(n6592), .B2(n6614), .A(n6591), .ZN(U3197) );
  AOI22_X1 U7519 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6835), .ZN(n6593) );
  OAI21_X1 U7520 ( .B1(n6595), .B2(n6611), .A(n6593), .ZN(U3198) );
  AOI22_X1 U7521 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6835), .ZN(n6594) );
  OAI21_X1 U7522 ( .B1(n6595), .B2(n6614), .A(n6594), .ZN(U3199) );
  AOI22_X1 U7523 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6835), .ZN(n6596) );
  OAI21_X1 U7524 ( .B1(n6597), .B2(n6614), .A(n6596), .ZN(U3200) );
  AOI22_X1 U7525 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6835), .ZN(n6598) );
  OAI21_X1 U7526 ( .B1(n5664), .B2(n6611), .A(n6598), .ZN(U3201) );
  AOI22_X1 U7527 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6835), .ZN(n6599) );
  OAI21_X1 U7528 ( .B1(n5664), .B2(n6614), .A(n6599), .ZN(U3202) );
  AOI22_X1 U7529 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6835), .ZN(n6600) );
  OAI21_X1 U7530 ( .B1(n6750), .B2(n6611), .A(n6600), .ZN(U3203) );
  AOI22_X1 U7531 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6835), .ZN(n6601) );
  OAI21_X1 U7532 ( .B1(n6750), .B2(n6614), .A(n6601), .ZN(U3204) );
  AOI22_X1 U7533 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6835), .ZN(n6602) );
  OAI21_X1 U7534 ( .B1(n6660), .B2(n6611), .A(n6602), .ZN(U3205) );
  AOI22_X1 U7535 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6835), .ZN(n6603) );
  OAI21_X1 U7536 ( .B1(n6660), .B2(n6614), .A(n6603), .ZN(U3206) );
  AOI22_X1 U7537 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6835), .ZN(n6604) );
  OAI21_X1 U7538 ( .B1(n6771), .B2(n6614), .A(n6604), .ZN(U3207) );
  AOI22_X1 U7539 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6835), .ZN(n6605) );
  OAI21_X1 U7540 ( .B1(n5605), .B2(n6614), .A(n6605), .ZN(U3208) );
  AOI22_X1 U7541 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6835), .ZN(n6606) );
  OAI21_X1 U7542 ( .B1(n6748), .B2(n6611), .A(n6606), .ZN(U3209) );
  AOI22_X1 U7543 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6835), .ZN(n6607) );
  OAI21_X1 U7544 ( .B1(n6808), .B2(n6611), .A(n6607), .ZN(U3210) );
  AOI22_X1 U7545 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6835), .ZN(n6608) );
  OAI21_X1 U7546 ( .B1(n6808), .B2(n6614), .A(n6608), .ZN(U3211) );
  AOI22_X1 U7547 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6609), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6835), .ZN(n6610) );
  OAI21_X1 U7548 ( .B1(n6787), .B2(n6611), .A(n6610), .ZN(U3212) );
  AOI22_X1 U7549 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6612), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6835), .ZN(n6613) );
  OAI21_X1 U7550 ( .B1(n6787), .B2(n6614), .A(n6613), .ZN(U3213) );
  MUX2_X1 U7551 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6835), .Z(U3446) );
  MUX2_X1 U7552 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6835), .Z(U3447) );
  MUX2_X1 U7553 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6835), .Z(U3448) );
  OAI21_X1 U7554 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6618), .A(n6616), .ZN(
        n6615) );
  INV_X1 U7555 ( .A(n6615), .ZN(U3451) );
  OAI21_X1 U7556 ( .B1(n6618), .B2(n6617), .A(n6616), .ZN(U3452) );
  INV_X1 U7557 ( .A(n6619), .ZN(n6622) );
  OAI211_X1 U7558 ( .C1(n6623), .C2(n6622), .A(n6621), .B(n6620), .ZN(U3453)
         );
  AOI21_X1 U7559 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6624) );
  OAI22_X1 U7560 ( .A1(REIP_REG_0__SCAN_IN), .A2(n6625), .B1(
        REIP_REG_1__SCAN_IN), .B2(n6624), .ZN(n6626) );
  INV_X1 U7561 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6815) );
  AOI22_X1 U7562 ( .A1(n6629), .A2(n6626), .B1(n6815), .B2(n6627), .ZN(U3468)
         );
  NOR2_X1 U7563 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6628) );
  INV_X1 U7564 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6790) );
  AOI22_X1 U7565 ( .A1(n6629), .A2(n6628), .B1(n6790), .B2(n6627), .ZN(U3469)
         );
  INV_X1 U7566 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6705) );
  OAI22_X1 U7567 ( .A1(n6835), .A2(n6705), .B1(W_R_N_REG_SCAN_IN), .B2(n6836), 
        .ZN(n6630) );
  INV_X1 U7568 ( .A(n6630), .ZN(U3470) );
  INV_X1 U7569 ( .A(n6631), .ZN(n6632) );
  AOI211_X1 U7570 ( .C1(n6634), .C2(n6822), .A(n6633), .B(n6632), .ZN(n6637)
         );
  OAI21_X1 U7571 ( .B1(n6637), .B2(n6636), .A(n6635), .ZN(n6641) );
  AOI211_X1 U7572 ( .C1(n6284), .C2(n6768), .A(n6639), .B(n6638), .ZN(n6640)
         );
  MUX2_X1 U7573 ( .A(n6641), .B(REQUESTPENDING_REG_SCAN_IN), .S(n6640), .Z(
        U3472) );
  INV_X1 U7574 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6688) );
  INV_X1 U7575 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6784) );
  AOI22_X1 U7576 ( .A1(n6836), .A2(n6688), .B1(n6784), .B2(n6835), .ZN(U3473)
         );
  AOI22_X1 U7577 ( .A1(keyinput_f46), .A2(W_R_N_REG_SCAN_IN), .B1(DATAI_10_), 
        .B2(keyinput_f21), .ZN(n6642) );
  OAI221_X1 U7578 ( .B1(keyinput_f46), .B2(W_R_N_REG_SCAN_IN), .C1(DATAI_10_), 
        .C2(keyinput_f21), .A(n6642), .ZN(n6703) );
  AOI22_X1 U7579 ( .A1(keyinput_f41), .A2(D_C_N_REG_SCAN_IN), .B1(DATAI_1_), 
        .B2(keyinput_f30), .ZN(n6643) );
  OAI221_X1 U7580 ( .B1(keyinput_f41), .B2(D_C_N_REG_SCAN_IN), .C1(DATAI_1_), 
        .C2(keyinput_f30), .A(n6643), .ZN(n6702) );
  AOI22_X1 U7581 ( .A1(keyinput_f40), .A2(M_IO_N_REG_SCAN_IN), .B1(n6747), 
        .B2(keyinput_f44), .ZN(n6644) );
  OAI221_X1 U7582 ( .B1(keyinput_f40), .B2(M_IO_N_REG_SCAN_IN), .C1(n6747), 
        .C2(keyinput_f44), .A(n6644), .ZN(n6654) );
  OAI22_X1 U7583 ( .A1(DATAI_29_), .A2(keyinput_f2), .B1(DATAI_25_), .B2(
        keyinput_f6), .ZN(n6645) );
  AOI221_X1 U7584 ( .B1(DATAI_29_), .B2(keyinput_f2), .C1(keyinput_f6), .C2(
        DATAI_25_), .A(n6645), .ZN(n6652) );
  OAI22_X1 U7585 ( .A1(REIP_REG_28__SCAN_IN), .A2(keyinput_f54), .B1(
        CODEFETCH_REG_SCAN_IN), .B2(keyinput_f39), .ZN(n6646) );
  AOI221_X1 U7586 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_f54), .C1(
        keyinput_f39), .C2(CODEFETCH_REG_SCAN_IN), .A(n6646), .ZN(n6651) );
  OAI22_X1 U7587 ( .A1(DATAI_31_), .A2(keyinput_f0), .B1(
        BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_f49), .ZN(n6647) );
  AOI221_X1 U7588 ( .B1(DATAI_31_), .B2(keyinput_f0), .C1(keyinput_f49), .C2(
        BYTEENABLE_REG_2__SCAN_IN), .A(n6647), .ZN(n6650) );
  OAI22_X1 U7589 ( .A1(REIP_REG_27__SCAN_IN), .A2(keyinput_f55), .B1(
        REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_f42), .ZN(n6648) );
  AOI221_X1 U7590 ( .B1(REIP_REG_27__SCAN_IN), .B2(keyinput_f55), .C1(
        keyinput_f42), .C2(REQUESTPENDING_REG_SCAN_IN), .A(n6648), .ZN(n6649)
         );
  NAND4_X1 U7591 ( .A1(n6652), .A2(n6651), .A3(n6650), .A4(n6649), .ZN(n6653)
         );
  AOI211_X1 U7592 ( .C1(keyinput_f20), .C2(DATAI_11_), .A(n6654), .B(n6653), 
        .ZN(n6655) );
  OAI21_X1 U7593 ( .B1(keyinput_f20), .B2(DATAI_11_), .A(n6655), .ZN(n6701) );
  AOI22_X1 U7594 ( .A1(DATAI_21_), .A2(keyinput_f10), .B1(REIP_REG_19__SCAN_IN), .B2(keyinput_f63), .ZN(n6656) );
  OAI221_X1 U7595 ( .B1(DATAI_21_), .B2(keyinput_f10), .C1(
        REIP_REG_19__SCAN_IN), .C2(keyinput_f63), .A(n6656), .ZN(n6666) );
  AOI22_X1 U7596 ( .A1(DATAI_27_), .A2(keyinput_f4), .B1(REIP_REG_20__SCAN_IN), 
        .B2(keyinput_f62), .ZN(n6657) );
  OAI221_X1 U7597 ( .B1(DATAI_27_), .B2(keyinput_f4), .C1(REIP_REG_20__SCAN_IN), .C2(keyinput_f62), .A(n6657), .ZN(n6665) );
  INV_X1 U7598 ( .A(DATAI_8_), .ZN(n6659) );
  AOI22_X1 U7599 ( .A1(n6660), .A2(keyinput_f59), .B1(keyinput_f23), .B2(n6659), .ZN(n6658) );
  OAI221_X1 U7600 ( .B1(n6660), .B2(keyinput_f59), .C1(n6659), .C2(
        keyinput_f23), .A(n6658), .ZN(n6664) );
  AOI22_X1 U7601 ( .A1(n6662), .A2(keyinput_f24), .B1(n6769), .B2(keyinput_f1), 
        .ZN(n6661) );
  OAI221_X1 U7602 ( .B1(n6662), .B2(keyinput_f24), .C1(n6769), .C2(keyinput_f1), .A(n6661), .ZN(n6663) );
  NOR4_X1 U7603 ( .A1(n6666), .A2(n6665), .A3(n6664), .A4(n6663), .ZN(n6699)
         );
  AOI22_X1 U7604 ( .A1(keyinput_f47), .A2(BYTEENABLE_REG_0__SCAN_IN), .B1(
        DATAI_2_), .B2(keyinput_f29), .ZN(n6667) );
  OAI221_X1 U7605 ( .B1(keyinput_f47), .B2(BYTEENABLE_REG_0__SCAN_IN), .C1(
        DATAI_2_), .C2(keyinput_f29), .A(n6667), .ZN(n6674) );
  AOI22_X1 U7606 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(DATAI_13_), .B2(
        keyinput_f18), .ZN(n6668) );
  OAI221_X1 U7607 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(DATAI_13_), .C2(
        keyinput_f18), .A(n6668), .ZN(n6673) );
  AOI22_X1 U7608 ( .A1(DATAI_16_), .A2(keyinput_f15), .B1(REIP_REG_25__SCAN_IN), .B2(keyinput_f57), .ZN(n6669) );
  OAI221_X1 U7609 ( .B1(DATAI_16_), .B2(keyinput_f15), .C1(
        REIP_REG_25__SCAN_IN), .C2(keyinput_f57), .A(n6669), .ZN(n6672) );
  AOI22_X1 U7610 ( .A1(DATAI_22_), .A2(keyinput_f9), .B1(DATAI_14_), .B2(
        keyinput_f17), .ZN(n6670) );
  OAI221_X1 U7611 ( .B1(DATAI_22_), .B2(keyinput_f9), .C1(DATAI_14_), .C2(
        keyinput_f17), .A(n6670), .ZN(n6671) );
  NOR4_X1 U7612 ( .A1(n6674), .A2(n6673), .A3(n6672), .A4(n6671), .ZN(n6698)
         );
  AOI22_X1 U7613 ( .A1(n6771), .A2(keyinput_f58), .B1(keyinput_f33), .B2(n6676), .ZN(n6675) );
  OAI221_X1 U7614 ( .B1(n6771), .B2(keyinput_f58), .C1(n6676), .C2(
        keyinput_f33), .A(n6675), .ZN(n6686) );
  AOI22_X1 U7615 ( .A1(n4677), .A2(keyinput_f13), .B1(keyinput_f48), .B2(n6820), .ZN(n6677) );
  OAI221_X1 U7616 ( .B1(n4677), .B2(keyinput_f13), .C1(n6820), .C2(
        keyinput_f48), .A(n6677), .ZN(n6685) );
  INV_X1 U7617 ( .A(DATAI_19_), .ZN(n6680) );
  INV_X1 U7618 ( .A(DATAI_12_), .ZN(n6679) );
  AOI22_X1 U7619 ( .A1(n6680), .A2(keyinput_f12), .B1(n6679), .B2(keyinput_f19), .ZN(n6678) );
  OAI221_X1 U7620 ( .B1(n6680), .B2(keyinput_f12), .C1(n6679), .C2(
        keyinput_f19), .A(n6678), .ZN(n6684) );
  AOI22_X1 U7621 ( .A1(n6792), .A2(keyinput_f51), .B1(keyinput_f3), .B2(n6682), 
        .ZN(n6681) );
  OAI221_X1 U7622 ( .B1(n6792), .B2(keyinput_f51), .C1(n6682), .C2(keyinput_f3), .A(n6681), .ZN(n6683) );
  NOR4_X1 U7623 ( .A1(n6686), .A2(n6685), .A3(n6684), .A4(n6683), .ZN(n6697)
         );
  AOI22_X1 U7624 ( .A1(n6688), .A2(keyinput_f32), .B1(n6822), .B2(keyinput_f43), .ZN(n6687) );
  OAI221_X1 U7625 ( .B1(n6688), .B2(keyinput_f32), .C1(n6822), .C2(
        keyinput_f43), .A(n6687), .ZN(n6695) );
  AOI22_X1 U7626 ( .A1(n6807), .A2(keyinput_f5), .B1(keyinput_f25), .B2(n6777), 
        .ZN(n6689) );
  OAI221_X1 U7627 ( .B1(n6807), .B2(keyinput_f5), .C1(n6777), .C2(keyinput_f25), .A(n6689), .ZN(n6694) );
  AOI22_X1 U7628 ( .A1(n6802), .A2(keyinput_f45), .B1(n6774), .B2(keyinput_f16), .ZN(n6690) );
  OAI221_X1 U7629 ( .B1(n6802), .B2(keyinput_f45), .C1(n6774), .C2(
        keyinput_f16), .A(n6690), .ZN(n6693) );
  AOI22_X1 U7630 ( .A1(n4664), .A2(keyinput_f14), .B1(keyinput_f31), .B2(n6818), .ZN(n6691) );
  OAI221_X1 U7631 ( .B1(n4664), .B2(keyinput_f14), .C1(n6818), .C2(
        keyinput_f31), .A(n6691), .ZN(n6692) );
  NOR4_X1 U7632 ( .A1(n6695), .A2(n6694), .A3(n6693), .A4(n6692), .ZN(n6696)
         );
  NAND4_X1 U7633 ( .A1(n6699), .A2(n6698), .A3(n6697), .A4(n6696), .ZN(n6700)
         );
  NOR4_X1 U7634 ( .A1(n6703), .A2(n6702), .A3(n6701), .A4(n6700), .ZN(n6728)
         );
  AOI22_X1 U7635 ( .A1(n6793), .A2(keyinput_f53), .B1(keyinput_f37), .B2(n6705), .ZN(n6704) );
  OAI221_X1 U7636 ( .B1(n6793), .B2(keyinput_f53), .C1(n6705), .C2(
        keyinput_f37), .A(n6704), .ZN(n6724) );
  AOI22_X1 U7637 ( .A1(n6785), .A2(keyinput_f26), .B1(keyinput_f38), .B2(n6778), .ZN(n6706) );
  OAI221_X1 U7638 ( .B1(n6785), .B2(keyinput_f26), .C1(n6778), .C2(
        keyinput_f38), .A(n6706), .ZN(n6723) );
  XOR2_X1 U7639 ( .A(keyinput_f34), .B(BS16_N), .Z(n6709) );
  AOI22_X1 U7640 ( .A1(n4681), .A2(keyinput_f8), .B1(n6787), .B2(keyinput_f52), 
        .ZN(n6707) );
  OAI221_X1 U7641 ( .B1(n4681), .B2(keyinput_f8), .C1(n6787), .C2(keyinput_f52), .A(n6707), .ZN(n6708) );
  AOI211_X1 U7642 ( .C1(n6814), .C2(keyinput_f50), .A(n6709), .B(n6708), .ZN(
        n6710) );
  OAI21_X1 U7643 ( .B1(n6814), .B2(keyinput_f50), .A(n6710), .ZN(n6722) );
  OAI22_X1 U7644 ( .A1(n6712), .A2(keyinput_f28), .B1(n6775), .B2(keyinput_f36), .ZN(n6711) );
  AOI221_X1 U7645 ( .B1(n6712), .B2(keyinput_f28), .C1(keyinput_f36), .C2(
        n6775), .A(n6711), .ZN(n6720) );
  OAI22_X1 U7646 ( .A1(n6750), .A2(keyinput_f61), .B1(n5727), .B2(keyinput_f56), .ZN(n6713) );
  AOI221_X1 U7647 ( .B1(n6750), .B2(keyinput_f61), .C1(keyinput_f56), .C2(
        n5727), .A(n6713), .ZN(n6719) );
  INV_X1 U7648 ( .A(DATAI_9_), .ZN(n6805) );
  OAI22_X1 U7649 ( .A1(n6805), .A2(keyinput_f22), .B1(n6715), .B2(keyinput_f27), .ZN(n6714) );
  AOI221_X1 U7650 ( .B1(n6805), .B2(keyinput_f22), .C1(keyinput_f27), .C2(
        n6715), .A(n6714), .ZN(n6718) );
  INV_X1 U7651 ( .A(DATAI_20_), .ZN(n6789) );
  OAI22_X1 U7652 ( .A1(n6768), .A2(keyinput_f35), .B1(n6789), .B2(keyinput_f11), .ZN(n6716) );
  AOI221_X1 U7653 ( .B1(n6768), .B2(keyinput_f35), .C1(keyinput_f11), .C2(
        n6789), .A(n6716), .ZN(n6717) );
  NAND4_X1 U7654 ( .A1(n6720), .A2(n6719), .A3(n6718), .A4(n6717), .ZN(n6721)
         );
  NOR4_X1 U7655 ( .A1(n6724), .A2(n6723), .A3(n6722), .A4(n6721), .ZN(n6727)
         );
  NOR2_X1 U7656 ( .A1(n6726), .A2(keyinput_f60), .ZN(n6725) );
  AOI221_X1 U7657 ( .B1(n6728), .B2(n6727), .C1(keyinput_f60), .C2(n6726), .A(
        n6725), .ZN(n6834) );
  AOI22_X1 U7658 ( .A1(D_C_N_REG_SCAN_IN), .A2(keyinput_g41), .B1(DATAI_7_), 
        .B2(keyinput_g24), .ZN(n6729) );
  OAI221_X1 U7659 ( .B1(D_C_N_REG_SCAN_IN), .B2(keyinput_g41), .C1(DATAI_7_), 
        .C2(keyinput_g24), .A(n6729), .ZN(n6736) );
  AOI22_X1 U7660 ( .A1(REIP_REG_19__SCAN_IN), .A2(keyinput_g63), .B1(
        REIP_REG_23__SCAN_IN), .B2(keyinput_g59), .ZN(n6730) );
  OAI221_X1 U7661 ( .B1(REIP_REG_19__SCAN_IN), .B2(keyinput_g63), .C1(
        REIP_REG_23__SCAN_IN), .C2(keyinput_g59), .A(n6730), .ZN(n6735) );
  AOI22_X1 U7662 ( .A1(DATAI_24_), .A2(keyinput_g7), .B1(DATAI_10_), .B2(
        keyinput_g21), .ZN(n6731) );
  OAI221_X1 U7663 ( .B1(DATAI_24_), .B2(keyinput_g7), .C1(DATAI_10_), .C2(
        keyinput_g21), .A(n6731), .ZN(n6734) );
  AOI22_X1 U7664 ( .A1(W_R_N_REG_SCAN_IN), .A2(keyinput_g46), .B1(DATAI_3_), 
        .B2(keyinput_g28), .ZN(n6732) );
  OAI221_X1 U7665 ( .B1(W_R_N_REG_SCAN_IN), .B2(keyinput_g46), .C1(DATAI_3_), 
        .C2(keyinput_g28), .A(n6732), .ZN(n6733) );
  NOR4_X1 U7666 ( .A1(n6736), .A2(n6735), .A3(n6734), .A4(n6733), .ZN(n6766)
         );
  XOR2_X1 U7667 ( .A(DATAI_25_), .B(keyinput_g6), .Z(n6743) );
  AOI22_X1 U7668 ( .A1(DATAI_21_), .A2(keyinput_g10), .B1(DATAI_13_), .B2(
        keyinput_g18), .ZN(n6737) );
  OAI221_X1 U7669 ( .B1(DATAI_21_), .B2(keyinput_g10), .C1(DATAI_13_), .C2(
        keyinput_g18), .A(n6737), .ZN(n6742) );
  AOI22_X1 U7670 ( .A1(DATAI_16_), .A2(keyinput_g15), .B1(REIP_REG_20__SCAN_IN), .B2(keyinput_g62), .ZN(n6738) );
  OAI221_X1 U7671 ( .B1(DATAI_16_), .B2(keyinput_g15), .C1(
        REIP_REG_20__SCAN_IN), .C2(keyinput_g62), .A(n6738), .ZN(n6741) );
  AOI22_X1 U7672 ( .A1(NA_N), .A2(keyinput_g33), .B1(DATAI_28_), .B2(
        keyinput_g3), .ZN(n6739) );
  OAI221_X1 U7673 ( .B1(NA_N), .B2(keyinput_g33), .C1(DATAI_28_), .C2(
        keyinput_g3), .A(n6739), .ZN(n6740) );
  NOR4_X1 U7674 ( .A1(n6743), .A2(n6742), .A3(n6741), .A4(n6740), .ZN(n6765)
         );
  AOI22_X1 U7675 ( .A1(READREQUEST_REG_SCAN_IN), .A2(keyinput_g37), .B1(
        DATAI_12_), .B2(keyinput_g19), .ZN(n6744) );
  OAI221_X1 U7676 ( .B1(READREQUEST_REG_SCAN_IN), .B2(keyinput_g37), .C1(
        DATAI_12_), .C2(keyinput_g19), .A(n6744), .ZN(n6754) );
  AOI22_X1 U7677 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_g32), .B1(
        DATAI_4_), .B2(keyinput_g27), .ZN(n6745) );
  OAI221_X1 U7678 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_g32), .C1(
        DATAI_4_), .C2(keyinput_g27), .A(n6745), .ZN(n6753) );
  AOI22_X1 U7679 ( .A1(n6748), .A2(keyinput_g55), .B1(keyinput_g44), .B2(n6747), .ZN(n6746) );
  OAI221_X1 U7680 ( .B1(n6748), .B2(keyinput_g55), .C1(n6747), .C2(
        keyinput_g44), .A(n6746), .ZN(n6752) );
  AOI22_X1 U7681 ( .A1(n6750), .A2(keyinput_g61), .B1(keyinput_g56), .B2(n5727), .ZN(n6749) );
  OAI221_X1 U7682 ( .B1(n6750), .B2(keyinput_g61), .C1(n5727), .C2(
        keyinput_g56), .A(n6749), .ZN(n6751) );
  NOR4_X1 U7683 ( .A1(n6754), .A2(n6753), .A3(n6752), .A4(n6751), .ZN(n6764)
         );
  AOI22_X1 U7684 ( .A1(DATAI_2_), .A2(keyinput_g29), .B1(DATAI_8_), .B2(
        keyinput_g23), .ZN(n6755) );
  OAI221_X1 U7685 ( .B1(DATAI_2_), .B2(keyinput_g29), .C1(DATAI_8_), .C2(
        keyinput_g23), .A(n6755), .ZN(n6762) );
  AOI22_X1 U7686 ( .A1(DATAI_19_), .A2(keyinput_g12), .B1(REIP_REG_25__SCAN_IN), .B2(keyinput_g57), .ZN(n6756) );
  OAI221_X1 U7687 ( .B1(DATAI_19_), .B2(keyinput_g12), .C1(
        REIP_REG_25__SCAN_IN), .C2(keyinput_g57), .A(n6756), .ZN(n6761) );
  AOI22_X1 U7688 ( .A1(BS16_N), .A2(keyinput_g34), .B1(DATAI_14_), .B2(
        keyinput_g17), .ZN(n6757) );
  OAI221_X1 U7689 ( .B1(BS16_N), .B2(keyinput_g34), .C1(DATAI_14_), .C2(
        keyinput_g17), .A(n6757), .ZN(n6760) );
  AOI22_X1 U7690 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_g42), .B1(
        DATAI_1_), .B2(keyinput_g30), .ZN(n6758) );
  OAI221_X1 U7691 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_g42), .C1(
        DATAI_1_), .C2(keyinput_g30), .A(n6758), .ZN(n6759) );
  NOR4_X1 U7692 ( .A1(n6762), .A2(n6761), .A3(n6760), .A4(n6759), .ZN(n6763)
         );
  NAND4_X1 U7693 ( .A1(n6766), .A2(n6765), .A3(n6764), .A4(n6763), .ZN(n6832)
         );
  AOI22_X1 U7694 ( .A1(n6769), .A2(keyinput_g1), .B1(n6768), .B2(keyinput_g35), 
        .ZN(n6767) );
  OAI221_X1 U7695 ( .B1(n6769), .B2(keyinput_g1), .C1(n6768), .C2(keyinput_g35), .A(n6767), .ZN(n6782) );
  AOI22_X1 U7696 ( .A1(n6772), .A2(keyinput_g2), .B1(n6771), .B2(keyinput_g58), 
        .ZN(n6770) );
  OAI221_X1 U7697 ( .B1(n6772), .B2(keyinput_g2), .C1(n6771), .C2(keyinput_g58), .A(n6770), .ZN(n6781) );
  AOI22_X1 U7698 ( .A1(n6775), .A2(keyinput_g36), .B1(n6774), .B2(keyinput_g16), .ZN(n6773) );
  OAI221_X1 U7699 ( .B1(n6775), .B2(keyinput_g36), .C1(n6774), .C2(
        keyinput_g16), .A(n6773), .ZN(n6780) );
  AOI22_X1 U7700 ( .A1(n6778), .A2(keyinput_g38), .B1(n6777), .B2(keyinput_g25), .ZN(n6776) );
  OAI221_X1 U7701 ( .B1(n6778), .B2(keyinput_g38), .C1(n6777), .C2(
        keyinput_g25), .A(n6776), .ZN(n6779) );
  NOR4_X1 U7702 ( .A1(n6782), .A2(n6781), .A3(n6780), .A4(n6779), .ZN(n6830)
         );
  AOI22_X1 U7703 ( .A1(n6785), .A2(keyinput_g26), .B1(keyinput_g40), .B2(n6784), .ZN(n6783) );
  OAI221_X1 U7704 ( .B1(n6785), .B2(keyinput_g26), .C1(n6784), .C2(
        keyinput_g40), .A(n6783), .ZN(n6797) );
  AOI22_X1 U7705 ( .A1(n4664), .A2(keyinput_g14), .B1(n6787), .B2(keyinput_g52), .ZN(n6786) );
  OAI221_X1 U7706 ( .B1(n4664), .B2(keyinput_g14), .C1(n6787), .C2(
        keyinput_g52), .A(n6786), .ZN(n6796) );
  AOI22_X1 U7707 ( .A1(n6790), .A2(keyinput_g47), .B1(n6789), .B2(keyinput_g11), .ZN(n6788) );
  OAI221_X1 U7708 ( .B1(n6790), .B2(keyinput_g47), .C1(n6789), .C2(
        keyinput_g11), .A(n6788), .ZN(n6795) );
  AOI22_X1 U7709 ( .A1(n6793), .A2(keyinput_g53), .B1(n6792), .B2(keyinput_g51), .ZN(n6791) );
  OAI221_X1 U7710 ( .B1(n6793), .B2(keyinput_g53), .C1(n6792), .C2(
        keyinput_g51), .A(n6791), .ZN(n6794) );
  NOR4_X1 U7711 ( .A1(n6797), .A2(n6796), .A3(n6795), .A4(n6794), .ZN(n6829)
         );
  AOI22_X1 U7712 ( .A1(n6799), .A2(keyinput_g4), .B1(keyinput_g13), .B2(n4677), 
        .ZN(n6798) );
  OAI221_X1 U7713 ( .B1(n6799), .B2(keyinput_g4), .C1(n4677), .C2(keyinput_g13), .A(n6798), .ZN(n6812) );
  AOI22_X1 U7714 ( .A1(n6802), .A2(keyinput_g45), .B1(n6801), .B2(keyinput_g0), 
        .ZN(n6800) );
  OAI221_X1 U7715 ( .B1(n6802), .B2(keyinput_g45), .C1(n6801), .C2(keyinput_g0), .A(n6800), .ZN(n6811) );
  AOI22_X1 U7716 ( .A1(n6805), .A2(keyinput_g22), .B1(keyinput_g39), .B2(n6804), .ZN(n6803) );
  OAI221_X1 U7717 ( .B1(n6805), .B2(keyinput_g22), .C1(n6804), .C2(
        keyinput_g39), .A(n6803), .ZN(n6810) );
  AOI22_X1 U7718 ( .A1(n6808), .A2(keyinput_g54), .B1(keyinput_g5), .B2(n6807), 
        .ZN(n6806) );
  OAI221_X1 U7719 ( .B1(n6808), .B2(keyinput_g54), .C1(n6807), .C2(keyinput_g5), .A(n6806), .ZN(n6809) );
  NOR4_X1 U7720 ( .A1(n6812), .A2(n6811), .A3(n6810), .A4(n6809), .ZN(n6828)
         );
  AOI22_X1 U7721 ( .A1(n6815), .A2(keyinput_g49), .B1(keyinput_g50), .B2(n6814), .ZN(n6813) );
  OAI221_X1 U7722 ( .B1(n6815), .B2(keyinput_g49), .C1(n6814), .C2(
        keyinput_g50), .A(n6813), .ZN(n6826) );
  INV_X1 U7723 ( .A(DATAI_11_), .ZN(n6817) );
  AOI22_X1 U7724 ( .A1(n6818), .A2(keyinput_g31), .B1(n6817), .B2(keyinput_g20), .ZN(n6816) );
  OAI221_X1 U7725 ( .B1(n6818), .B2(keyinput_g31), .C1(n6817), .C2(
        keyinput_g20), .A(n6816), .ZN(n6825) );
  AOI22_X1 U7726 ( .A1(n4689), .A2(keyinput_g9), .B1(keyinput_g48), .B2(n6820), 
        .ZN(n6819) );
  OAI221_X1 U7727 ( .B1(n4689), .B2(keyinput_g9), .C1(n6820), .C2(keyinput_g48), .A(n6819), .ZN(n6824) );
  AOI22_X1 U7728 ( .A1(n4681), .A2(keyinput_g8), .B1(n6822), .B2(keyinput_g43), 
        .ZN(n6821) );
  OAI221_X1 U7729 ( .B1(n4681), .B2(keyinput_g8), .C1(n6822), .C2(keyinput_g43), .A(n6821), .ZN(n6823) );
  NOR4_X1 U7730 ( .A1(n6826), .A2(n6825), .A3(n6824), .A4(n6823), .ZN(n6827)
         );
  NAND4_X1 U7731 ( .A1(n6830), .A2(n6829), .A3(n6828), .A4(n6827), .ZN(n6831)
         );
  OAI22_X1 U7732 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput_g60), .B1(n6832), 
        .B2(n6831), .ZN(n6833) );
  AOI211_X1 U7733 ( .C1(REIP_REG_22__SCAN_IN), .C2(keyinput_g60), .A(n6834), 
        .B(n6833), .ZN(n6838) );
  AOI22_X1 U7734 ( .A1(n6836), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6835), .ZN(n6837) );
  XNOR2_X1 U7735 ( .A(n6838), .B(n6837), .ZN(U3445) );
  OR2_X1 U3439 ( .A1(n4069), .A2(n4124), .ZN(n3204) );
  CLKBUF_X1 U34460 ( .A(n3230), .Z(n3232) );
  AND4_X1 U3450 ( .A1(n3152), .A2(n3151), .A3(n3150), .A4(n3149), .ZN(n3153)
         );
  CLKBUF_X1 U3454 ( .A(n3187), .Z(n3212) );
  CLKBUF_X1 U3798 ( .A(n3221), .Z(n5374) );
  CLKBUF_X3 U4177 ( .A(n3194), .Z(n3313) );
  CLKBUF_X1 U4183 ( .A(n3357), .Z(n3358) );
  CLKBUF_X1 U4198 ( .A(n6283), .Z(n6274) );
endmodule

