

module b21_C_AntiSAT_k_128_3 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073;

  AND2_X1 U4801 ( .A1(n8594), .A2(n4344), .ZN(n8499) );
  NAND2_X1 U4802 ( .A1(n4603), .A2(n4601), .ZN(n8191) );
  CLKBUF_X1 U4803 ( .A(n5041), .Z(n5480) );
  INV_X2 U4804 ( .A(n5461), .ZN(n5617) );
  NAND2_X1 U4805 ( .A1(n7866), .A2(n7407), .ZN(n8375) );
  CLKBUF_X1 U4806 ( .A(n5812), .Z(n6224) );
  AND4_X1 U4807 ( .A1(n5755), .A2(n5754), .A3(n5753), .A4(n5752), .ZN(n7581)
         );
  NAND2_X1 U4808 ( .A1(n6700), .A2(n5746), .ZN(n5792) );
  OR2_X1 U4809 ( .A1(n5734), .A2(n5976), .ZN(n5735) );
  OR2_X1 U4810 ( .A1(n5732), .A2(n7997), .ZN(n7809) );
  CLKBUF_X2 U4811 ( .A(n5835), .Z(n4298) );
  AND2_X1 U4812 ( .A1(n7475), .A2(n7341), .ZN(n7367) );
  XNOR2_X1 U4813 ( .A(n5739), .B(n5738), .ZN(n5741) );
  INV_X1 U4814 ( .A(n5581), .ZN(n6268) );
  NAND2_X1 U4815 ( .A1(n5773), .A2(n5772), .ZN(n7754) );
  AND4_X1 U4816 ( .A1(n5767), .A2(n5766), .A3(n5765), .A4(n5764), .ZN(n8373)
         );
  AOI22_X1 U4817 ( .A1(n8191), .A2(n7963), .B1(n8204), .B2(n8008), .ZN(n8176)
         );
  NAND2_X1 U4818 ( .A1(n5737), .A2(n5736), .ZN(n7580) );
  AND4_X1 U4819 ( .A1(n4956), .A2(n5192), .A3(n5149), .A4(n5152), .ZN(n4296)
         );
  XNOR2_X2 U4820 ( .A(n4977), .B(P1_IR_REG_28__SCAN_IN), .ZN(n5657) );
  INV_X1 U4821 ( .A(n6498), .ZN(n6478) );
  OAI211_X4 U4823 ( .C1(n6302), .C2(n9508), .A(n5098), .B(n5097), .ZN(n6457)
         );
  AND2_X1 U4824 ( .A1(n5741), .A2(n7580), .ZN(n5835) );
  OR2_X2 U4825 ( .A1(n6212), .A2(n5719), .ZN(n5732) );
  AOI21_X2 U4826 ( .B1(n7529), .B2(n7927), .A(n7528), .ZN(n8342) );
  NAND2_X2 U4827 ( .A1(n7499), .A2(n4725), .ZN(n7529) );
  INV_X1 U4828 ( .A(n5041), .ZN(n4299) );
  NAND4_X2 U4829 ( .A1(n5856), .A2(n5855), .A3(n5854), .A4(n5853), .ZN(n9683)
         );
  OAI22_X2 U4830 ( .A1(n7269), .A2(n7884), .B1(n7268), .B2(n9681), .ZN(n7270)
         );
  AOI21_X1 U4831 ( .B1(n4310), .B2(n7630), .A(n9431), .ZN(n7634) );
  NAND2_X1 U4832 ( .A1(n4786), .A2(n4784), .ZN(n8563) );
  NAND2_X1 U4833 ( .A1(n8546), .A2(n4787), .ZN(n4786) );
  OR2_X1 U4834 ( .A1(n8537), .A2(n4842), .ZN(n8545) );
  XNOR2_X1 U4835 ( .A(n4545), .B(n6097), .ZN(n7742) );
  AOI21_X1 U4836 ( .B1(n4785), .B2(n4789), .A(n4328), .ZN(n4784) );
  AND2_X1 U4837 ( .A1(n5346), .A2(n5347), .ZN(n7167) );
  AND2_X1 U4838 ( .A1(n7432), .A2(n7431), .ZN(n7433) );
  NAND2_X1 U4839 ( .A1(n7367), .A2(n7820), .ZN(n7366) );
  NAND2_X1 U4840 ( .A1(n7103), .A2(n5845), .ZN(n7066) );
  INV_X4 U4841 ( .A(n9653), .ZN(n9405) );
  INV_X1 U4842 ( .A(n7215), .ZN(n9755) );
  OAI21_X1 U4843 ( .B1(n5227), .B2(n5228), .A(n4878), .ZN(n5215) );
  NAND2_X1 U4844 ( .A1(n8750), .A2(n8754), .ZN(n6483) );
  NAND2_X1 U4845 ( .A1(n7844), .A2(n7865), .ZN(n7201) );
  INV_X2 U4846 ( .A(n5041), .ZN(n5605) );
  NAND2_X1 U4847 ( .A1(n6442), .A2(n5057), .ZN(n5161) );
  OR2_X1 U4848 ( .A1(n6336), .A2(n4350), .ZN(n6357) );
  OR2_X1 U4849 ( .A1(n7990), .A2(n5719), .ZN(n5725) );
  NAND2_X1 U4850 ( .A1(n6439), .A2(n5057), .ZN(n5041) );
  NAND2_X4 U4851 ( .A1(n5654), .A2(n8830), .ZN(n6336) );
  INV_X2 U4852 ( .A(n8023), .ZN(n7191) );
  INV_X1 U4853 ( .A(n8373), .ZN(n8025) );
  NAND2_X1 U4854 ( .A1(n5648), .A2(n6837), .ZN(n6439) );
  CLKBUF_X3 U4855 ( .A(n5085), .Z(n8625) );
  AND2_X1 U4856 ( .A1(n5019), .A2(n9362), .ZN(n5085) );
  CLKBUF_X2 U4857 ( .A(n5066), .Z(n6302) );
  NAND2_X1 U4858 ( .A1(n5627), .A2(n4995), .ZN(n5057) );
  OR2_X1 U4859 ( .A1(n4611), .A2(n4610), .ZN(n7751) );
  NAND2_X1 U4860 ( .A1(n5066), .A2(n5746), .ZN(n5093) );
  XNOR2_X1 U4861 ( .A(n4993), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5627) );
  AOI21_X1 U4862 ( .B1(n4872), .B2(n4620), .A(n4335), .ZN(n4619) );
  XNOR2_X1 U4863 ( .A(n4775), .B(P1_IR_REG_22__SCAN_IN), .ZN(n5046) );
  INV_X2 U4864 ( .A(n5792), .ZN(n7565) );
  INV_X2 U4865 ( .A(n5793), .ZN(n7566) );
  OAI21_X1 U4866 ( .B1(n4983), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4775) );
  AND2_X1 U4867 ( .A1(n5015), .A2(n9355), .ZN(n5018) );
  NAND2_X1 U4868 ( .A1(n9355), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5017) );
  AND2_X1 U4869 ( .A1(n4990), .A2(n4975), .ZN(n4978) );
  NAND2_X1 U4870 ( .A1(n5014), .A2(n4319), .ZN(n9355) );
  INV_X2 U4871 ( .A(n7619), .ZN(n7626) );
  NAND2_X2 U4872 ( .A1(n6229), .A2(n7998), .ZN(n6700) );
  NAND2_X1 U4873 ( .A1(n4982), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4989) );
  NAND2_X1 U4874 ( .A1(n4799), .A2(n4694), .ZN(n5011) );
  MUX2_X1 U4875 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5735), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5736) );
  NAND2_X1 U4876 ( .A1(n5737), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5739) );
  AND2_X1 U4877 ( .A1(n5876), .A2(n4349), .ZN(n5974) );
  NAND2_X2 U4878 ( .A1(n4666), .A2(n4664), .ZN(n4859) );
  AND4_X1 U4879 ( .A1(n5698), .A2(n4753), .A3(n5687), .A4(n4429), .ZN(n5706)
         );
  AND2_X1 U4880 ( .A1(n4800), .A2(n4969), .ZN(n4694) );
  NOR2_X1 U4881 ( .A1(n4971), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4800) );
  INV_X1 U4882 ( .A(n5825), .ZN(n5687) );
  AND2_X1 U4883 ( .A1(n4578), .A2(n4756), .ZN(n4755) );
  AND2_X1 U4884 ( .A1(n4958), .A2(n4957), .ZN(n5150) );
  XNOR2_X1 U4885 ( .A(n4452), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6298) );
  NOR2_X1 U4886 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4728) );
  NOR2_X1 U4887 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4727) );
  INV_X1 U4888 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4988) );
  INV_X1 U4889 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4735) );
  NOR2_X1 U4890 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4956) );
  NOR2_X1 U4891 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4578) );
  NOR2_X1 U4892 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5693) );
  NOR2_X1 U4893 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5692) );
  NOR2_X1 U4894 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5694) );
  INV_X2 U4895 ( .A(n8889), .ZN(n6456) );
  AND3_X2 U4896 ( .A1(n5072), .A2(n5071), .A3(n5070), .ZN(n6435) );
  AND2_X1 U4897 ( .A1(n4755), .A2(n4754), .ZN(n4753) );
  INV_X1 U4898 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4754) );
  OR2_X1 U4899 ( .A1(n8402), .A2(n8006), .ZN(n7835) );
  NOR2_X1 U4900 ( .A1(n4597), .A2(n7596), .ZN(n4595) );
  OR2_X1 U4901 ( .A1(n9252), .A2(n9023), .ZN(n8827) );
  NAND2_X1 U4902 ( .A1(n9308), .A2(n9198), .ZN(n4722) );
  NAND2_X1 U4903 ( .A1(n8299), .A2(n4744), .ZN(n4743) );
  NOR2_X1 U4904 ( .A1(n8275), .A2(n4745), .ZN(n4744) );
  INV_X1 U4905 ( .A(n7948), .ZN(n4745) );
  INV_X1 U4906 ( .A(n6700), .ZN(n6514) );
  MUX2_X1 U4907 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5700), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n5703) );
  NAND2_X1 U4908 ( .A1(n5722), .A2(n5721), .ZN(n5724) );
  NOR2_X1 U4909 ( .A1(n9252), .A2(n9256), .ZN(n4480) );
  AND2_X1 U4910 ( .A1(n9002), .A2(n9003), .ZN(n9027) );
  OR2_X1 U4911 ( .A1(n6994), .A2(n4706), .ZN(n4705) );
  INV_X1 U4912 ( .A(n6927), .ZN(n4706) );
  INV_X1 U4913 ( .A(n5568), .ZN(n4655) );
  AND2_X1 U4914 ( .A1(n4641), .A2(n4836), .ZN(n4640) );
  NAND2_X1 U4915 ( .A1(n5290), .A2(n4902), .ZN(n4641) );
  INV_X1 U4916 ( .A(n7580), .ZN(n5740) );
  OR2_X1 U4917 ( .A1(n8414), .A2(n8008), .ZN(n7967) );
  NOR2_X1 U4918 ( .A1(n4444), .A2(n8422), .ZN(n4443) );
  INV_X1 U4919 ( .A(n4445), .ZN(n4444) );
  OR2_X1 U4920 ( .A1(n8422), .A2(n8242), .ZN(n7958) );
  OR2_X1 U4921 ( .A1(n7338), .A2(n7467), .ZN(n7890) );
  NAND2_X1 U4922 ( .A1(n8373), .A2(n7751), .ZN(n8374) );
  NAND2_X1 U4923 ( .A1(n7381), .A2(n7841), .ZN(n7857) );
  AOI21_X1 U4924 ( .B1(n9706), .B2(n9713), .A(n9714), .ZN(n8391) );
  AND2_X1 U4925 ( .A1(n5687), .A2(n4755), .ZN(n5876) );
  AND2_X1 U4926 ( .A1(n4783), .A2(n6983), .ZN(n4780) );
  INV_X1 U4927 ( .A(n6984), .ZN(n4778) );
  INV_X1 U4928 ( .A(n5020), .ZN(n5019) );
  INV_X1 U4929 ( .A(n5086), .ZN(n5581) );
  NAND2_X1 U4930 ( .A1(n5602), .A2(n5601), .ZN(n7541) );
  INV_X1 U4931 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4991) );
  NAND2_X1 U4932 ( .A1(n5429), .A2(n5428), .ZN(n4634) );
  NAND2_X1 U4933 ( .A1(n4920), .A2(n4919), .ZN(n4923) );
  NAND2_X1 U4934 ( .A1(n4912), .A2(n4911), .ZN(n5351) );
  AOI21_X1 U4935 ( .B1(n4640), .B2(n4638), .A(n4637), .ZN(n4636) );
  INV_X1 U4936 ( .A(n4908), .ZN(n4637) );
  INV_X1 U4937 ( .A(n4902), .ZN(n4638) );
  NAND2_X1 U4938 ( .A1(n4494), .A2(n4895), .ZN(n5291) );
  AOI21_X1 U4939 ( .B1(n7742), .B2(n7741), .A(n6100), .ZN(n6116) );
  AND2_X1 U4940 ( .A1(n8492), .A2(n7580), .ZN(n5779) );
  NAND2_X1 U4941 ( .A1(n5895), .A2(n7121), .ZN(n7648) );
  NAND2_X1 U4942 ( .A1(n4555), .A2(n4552), .ZN(n5895) );
  NOR2_X1 U4943 ( .A1(n4554), .A2(n7122), .ZN(n4552) );
  AOI21_X1 U4944 ( .B1(n7980), .B2(n4390), .A(n4389), .ZN(n4387) );
  AND2_X1 U4945 ( .A1(n4393), .A2(n6858), .ZN(n4390) );
  AND2_X1 U4946 ( .A1(n4391), .A2(n6858), .ZN(n4389) );
  AOI21_X1 U4947 ( .B1(n8162), .B2(n6224), .A(n6176), .ZN(n8006) );
  INV_X1 U4948 ( .A(n5779), .ZN(n5834) );
  NAND2_X1 U4949 ( .A1(n9354), .A2(n7565), .ZN(n4623) );
  AND2_X1 U4950 ( .A1(n8153), .A2(n7613), .ZN(n8398) );
  AOI21_X1 U4951 ( .B1(n4741), .B2(n4738), .A(n4330), .ZN(n4737) );
  INV_X1 U4952 ( .A(n4741), .ZN(n4739) );
  NAND2_X1 U4953 ( .A1(n5720), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5722) );
  NAND2_X1 U4954 ( .A1(n4559), .A2(n4557), .ZN(n5720) );
  OAI21_X1 U4955 ( .B1(n7594), .B2(n4338), .A(n4589), .ZN(n4588) );
  NOR2_X1 U4956 ( .A1(n4590), .A2(n7598), .ZN(n4589) );
  OR2_X1 U4957 ( .A1(n8445), .A2(n8277), .ZN(n7948) );
  NOR2_X1 U4958 ( .A1(n7771), .A2(n7714), .ZN(n7590) );
  OR2_X1 U4959 ( .A1(n8465), .A2(n8331), .ZN(n4837) );
  NAND2_X1 U4960 ( .A1(n7855), .A2(n7841), .ZN(n7384) );
  NAND2_X1 U4961 ( .A1(n6075), .A2(n6074), .ZN(n8440) );
  OR2_X1 U4962 ( .A1(n5732), .A2(n8394), .ZN(n9801) );
  AND2_X1 U4963 ( .A1(n5699), .A2(n4430), .ZN(n4429) );
  INV_X1 U4964 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4430) );
  INV_X2 U4965 ( .A(n4859), .ZN(n5746) );
  INV_X1 U4966 ( .A(n5107), .ZN(n5105) );
  OR2_X1 U4967 ( .A1(n5551), .A2(n8598), .ZN(n5607) );
  INV_X1 U4968 ( .A(n5578), .ZN(n5658) );
  AND2_X1 U4969 ( .A1(n5020), .A2(n9362), .ZN(n5086) );
  AND2_X1 U4970 ( .A1(n8827), .A2(n8861), .ZN(n8979) );
  INV_X1 U4971 ( .A(n8977), .ZN(n4698) );
  NOR2_X1 U4972 ( .A1(n9057), .A2(n9262), .ZN(n9031) );
  OR2_X1 U4973 ( .A1(n9282), .A2(n8966), .ZN(n8997) );
  NAND2_X1 U4974 ( .A1(n9107), .A2(n4823), .ZN(n9091) );
  OR2_X1 U4975 ( .A1(n9297), .A2(n9136), .ZN(n8992) );
  AOI21_X1 U4976 ( .B1(n4718), .B2(n4715), .A(n4714), .ZN(n4713) );
  NOR2_X1 U4977 ( .A1(n9163), .A2(n8961), .ZN(n4714) );
  NOR2_X1 U4978 ( .A1(n8962), .A2(n4719), .ZN(n4715) );
  INV_X1 U4979 ( .A(n8962), .ZN(n4717) );
  OR2_X1 U4980 ( .A1(n9322), .A2(n9210), .ZN(n9204) );
  AOI21_X1 U4981 ( .B1(n9322), .B2(n8958), .A(n8957), .ZN(n9203) );
  NAND2_X1 U4982 ( .A1(n9473), .A2(n4509), .ZN(n8981) );
  NAND2_X1 U4983 ( .A1(n4691), .A2(n4312), .ZN(n4690) );
  INV_X1 U4984 ( .A(n4692), .ZN(n4691) );
  AOI21_X1 U4985 ( .B1(n8763), .B2(n7312), .A(n4336), .ZN(n4692) );
  OAI22_X1 U4986 ( .A1(n7014), .A2(n7013), .B1(n9395), .B2(n7025), .ZN(n7309)
         );
  NOR2_X1 U4987 ( .A1(n7012), .A2(n8880), .ZN(n7013) );
  INV_X1 U4988 ( .A(n8635), .ZN(n5412) );
  INV_X1 U4989 ( .A(n6302), .ZN(n5411) );
  INV_X1 U4990 ( .A(n9208), .ZN(n9401) );
  NAND2_X1 U4991 ( .A1(n8637), .A2(n8636), .ZN(n9252) );
  MUX2_X1 U4992 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5012), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5015) );
  INV_X4 U4993 ( .A(n5746), .ZN(n7548) );
  NAND2_X1 U4994 ( .A1(n6006), .A2(n6005), .ZN(n8451) );
  AOI21_X1 U4995 ( .B1(n7806), .B2(n7981), .A(n7979), .ZN(n7807) );
  OAI21_X1 U4996 ( .B1(n8654), .B2(n8738), .A(n8655), .ZN(n8664) );
  AOI21_X1 U4997 ( .B1(n7873), .B2(n4307), .A(n7872), .ZN(n4421) );
  OR2_X1 U4998 ( .A1(n7863), .A2(n7986), .ZN(n4425) );
  INV_X1 U4999 ( .A(n7918), .ZN(n4406) );
  AND2_X1 U5000 ( .A1(n8696), .A2(n8741), .ZN(n4500) );
  OAI21_X1 U5001 ( .B1(n8697), .B2(n8741), .A(n9222), .ZN(n4499) );
  INV_X1 U5002 ( .A(n4405), .ZN(n4404) );
  AOI21_X1 U5003 ( .B1(n4405), .B2(n4403), .A(n4402), .ZN(n4401) );
  INV_X1 U5004 ( .A(n7914), .ZN(n4403) );
  INV_X1 U5005 ( .A(n4419), .ZN(n4418) );
  OAI22_X1 U5006 ( .A1(n7953), .A2(n7989), .B1(n7940), .B2(n7986), .ZN(n4419)
         );
  INV_X1 U5007 ( .A(n7940), .ZN(n4420) );
  INV_X1 U5008 ( .A(n7959), .ZN(n4417) );
  OAI21_X1 U5009 ( .B1(n8730), .B2(n4485), .A(n8729), .ZN(n8733) );
  NOR2_X1 U5010 ( .A1(n4752), .A2(n7206), .ZN(n4749) );
  NAND2_X1 U5011 ( .A1(n8025), .A2(n9729), .ZN(n7854) );
  NAND2_X1 U5012 ( .A1(n5711), .A2(n4550), .ZN(n4549) );
  INV_X1 U5013 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4550) );
  AOI21_X1 U5014 ( .B1(n4649), .B2(n4646), .A(n4340), .ZN(n4645) );
  INV_X1 U5015 ( .A(n4917), .ZN(n4646) );
  INV_X1 U5016 ( .A(n4923), .ZN(n4651) );
  INV_X1 U5017 ( .A(n4649), .ZN(n4647) );
  NOR2_X1 U5018 ( .A1(n4639), .A2(n4493), .ZN(n4492) );
  INV_X1 U5019 ( .A(n4895), .ZN(n4493) );
  INV_X1 U5020 ( .A(n4640), .ZN(n4639) );
  NAND2_X1 U5021 ( .A1(n4905), .A2(n4904), .ZN(n4908) );
  NAND2_X1 U5022 ( .A1(n4892), .A2(n4495), .ZN(n4494) );
  INV_X1 U5023 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5149) );
  OR2_X1 U5024 ( .A1(n5885), .A2(n5884), .ZN(n5900) );
  NAND2_X1 U5025 ( .A1(n4623), .A2(n4622), .ZN(n7988) );
  AND2_X1 U5026 ( .A1(n7803), .A2(n7558), .ZN(n4622) );
  NAND2_X1 U5027 ( .A1(n4392), .A2(n4396), .ZN(n4391) );
  NAND2_X1 U5028 ( .A1(n4397), .A2(n7986), .ZN(n4396) );
  NAND2_X1 U5029 ( .A1(n4393), .A2(n7979), .ZN(n4392) );
  INV_X1 U5030 ( .A(n7988), .ZN(n4397) );
  NAND2_X1 U5031 ( .A1(n8072), .A2(n4369), .ZN(n8081) );
  AND2_X1 U5032 ( .A1(n8182), .A2(n7969), .ZN(n4741) );
  NOR2_X1 U5033 ( .A1(n4605), .A2(n8211), .ZN(n4604) );
  INV_X1 U5034 ( .A(n4606), .ZN(n4605) );
  AND2_X1 U5035 ( .A1(n8231), .A2(n7943), .ZN(n4760) );
  NOR2_X1 U5036 ( .A1(n8231), .A2(n4607), .ZN(n4606) );
  INV_X1 U5037 ( .A(n7600), .ZN(n4607) );
  OR2_X1 U5038 ( .A1(n8434), .A2(n8278), .ZN(n7953) );
  AOI21_X1 U5039 ( .B1(n8314), .B2(n8313), .A(n7944), .ZN(n8292) );
  INV_X1 U5040 ( .A(n4837), .ZN(n4586) );
  AND2_X1 U5041 ( .A1(n9762), .A2(n9755), .ZN(n4428) );
  NAND2_X1 U5042 ( .A1(n8023), .A2(n9741), .ZN(n7865) );
  NAND2_X1 U5043 ( .A1(n7411), .A2(n7458), .ZN(n7846) );
  NOR2_X1 U5044 ( .A1(n7401), .A2(n7211), .ZN(n7402) );
  NAND2_X1 U5045 ( .A1(n7412), .A2(n8367), .ZN(n7407) );
  NAND2_X1 U5046 ( .A1(n4559), .A2(n5715), .ZN(n6033) );
  INV_X1 U5047 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5955) );
  INV_X1 U5048 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5712) );
  INV_X1 U5049 ( .A(n4549), .ZN(n4548) );
  NOR2_X1 U5050 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n4426) );
  INV_X1 U5051 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5958) );
  INV_X1 U5052 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4731) );
  NAND2_X1 U5053 ( .A1(n4733), .A2(n4735), .ZN(n4729) );
  INV_X1 U5054 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4736) );
  INV_X1 U5055 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4662) );
  NOR2_X1 U5056 ( .A1(P1_RD_REG_SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n4846) );
  NAND2_X1 U5057 ( .A1(n4793), .A2(n4795), .ZN(n4794) );
  INV_X1 U5058 ( .A(n4838), .ZN(n4795) );
  INV_X1 U5059 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5320) );
  OAI21_X1 U5060 ( .B1(n8523), .B2(n8522), .A(n4381), .ZN(n5485) );
  OR2_X1 U5061 ( .A1(n5465), .A2(n5464), .ZN(n4381) );
  OR2_X1 U5062 ( .A1(n9256), .A2(n9049), .ZN(n9002) );
  AND2_X1 U5063 ( .A1(n8745), .A2(n9077), .ZN(n8998) );
  INV_X1 U5064 ( .A(n8991), .ZN(n4815) );
  OR2_X1 U5065 ( .A1(n9287), .A2(n9135), .ZN(n8994) );
  OR2_X1 U5066 ( .A1(n9294), .A2(n8963), .ZN(n8796) );
  NOR2_X1 U5067 ( .A1(n4689), .A2(n4688), .ZN(n4687) );
  NAND2_X1 U5068 ( .A1(n4693), .A2(n7312), .ZN(n4688) );
  NOR2_X1 U5069 ( .A1(n4690), .A2(n8956), .ZN(n4686) );
  OR2_X1 U5070 ( .A1(n5321), .A2(n5320), .ZN(n5339) );
  INV_X1 U5071 ( .A(n4704), .ZN(n4703) );
  OAI22_X1 U5072 ( .A1(n6843), .A2(n4705), .B1(n7112), .B2(n8882), .ZN(n4704)
         );
  NAND2_X1 U5073 ( .A1(n4834), .A2(n8820), .ZN(n4833) );
  INV_X1 U5074 ( .A(n6924), .ZN(n4834) );
  INV_X1 U5075 ( .A(n8758), .ZN(n6843) );
  NAND2_X1 U5076 ( .A1(n8656), .A2(n8754), .ZN(n4810) );
  OAI21_X1 U5077 ( .B1(n7541), .B2(n4630), .A(n4628), .ZN(n7551) );
  INV_X1 U5078 ( .A(n4631), .ZN(n4630) );
  AOI21_X1 U5079 ( .B1(n4631), .B2(n4629), .A(n4373), .ZN(n4628) );
  NOR2_X1 U5080 ( .A1(n4632), .A2(n7547), .ZN(n4631) );
  XNOR2_X1 U5081 ( .A(n7551), .B(n7550), .ZN(n7564) );
  XNOR2_X1 U5082 ( .A(n4979), .B(P1_IR_REG_27__SCAN_IN), .ZN(n6284) );
  AND2_X1 U5083 ( .A1(n5570), .A2(n5548), .ZN(n5568) );
  NAND2_X1 U5084 ( .A1(n4931), .A2(n4930), .ZN(n5410) );
  AND2_X1 U5085 ( .A1(n5367), .A2(n4650), .ZN(n4649) );
  NAND2_X1 U5086 ( .A1(n5350), .A2(n4917), .ZN(n4650) );
  INV_X1 U5087 ( .A(n4492), .ZN(n4491) );
  NAND2_X1 U5088 ( .A1(n4492), .A2(n4490), .ZN(n4489) );
  INV_X1 U5089 ( .A(n4495), .ZN(n4490) );
  NAND2_X1 U5090 ( .A1(n4899), .A2(n4898), .ZN(n4902) );
  NAND2_X1 U5091 ( .A1(n5252), .A2(n4839), .ZN(n4892) );
  INV_X1 U5092 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U5093 ( .A1(n7515), .A2(n4533), .ZN(n9433) );
  NOR2_X1 U5094 ( .A1(n9429), .A2(n4534), .ZN(n4533) );
  INV_X1 U5095 ( .A(n5954), .ZN(n4534) );
  OR2_X1 U5096 ( .A1(n7649), .A2(n4532), .ZN(n4531) );
  INV_X1 U5097 ( .A(n7390), .ZN(n4532) );
  AOI21_X1 U5098 ( .B1(n7390), .B2(n4530), .A(n4317), .ZN(n4529) );
  INV_X1 U5099 ( .A(n7480), .ZN(n4526) );
  NOR2_X1 U5100 ( .A1(n5907), .A2(n5906), .ZN(n4530) );
  INV_X1 U5101 ( .A(n6039), .ZN(n6007) );
  AND2_X1 U5102 ( .A1(n5824), .A2(n5805), .ZN(n4547) );
  AND2_X1 U5103 ( .A1(n6147), .A2(n6146), .ZN(n8008) );
  AND2_X1 U5104 ( .A1(n6134), .A2(n6133), .ZN(n7773) );
  NAND2_X1 U5105 ( .A1(n6704), .A2(n4511), .ZN(n9367) );
  NAND2_X1 U5106 ( .A1(n6737), .A2(n4512), .ZN(n4511) );
  NOR2_X1 U5107 ( .A1(n8033), .A2(n4524), .ZN(n8048) );
  AND2_X1 U5108 ( .A1(n6735), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4524) );
  OR2_X1 U5109 ( .A1(n8048), .A2(n8049), .ZN(n4523) );
  AND2_X1 U5110 ( .A1(n4523), .A2(n4522), .ZN(n8062) );
  NAND2_X1 U5111 ( .A1(n6734), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4522) );
  OR2_X1 U5112 ( .A1(n6762), .A2(n6761), .ZN(n4517) );
  AND2_X1 U5113 ( .A1(n4517), .A2(n4516), .ZN(n6773) );
  NAND2_X1 U5114 ( .A1(n6727), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4516) );
  OR2_X1 U5115 ( .A1(n6773), .A2(n6772), .ZN(n4515) );
  XNOR2_X1 U5116 ( .A(n8081), .B(n8082), .ZN(n8074) );
  NOR2_X1 U5117 ( .A1(n8074), .A2(n9448), .ZN(n8083) );
  XNOR2_X1 U5118 ( .A(n4513), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8144) );
  NAND2_X1 U5119 ( .A1(n8137), .A2(n4375), .ZN(n4513) );
  NAND2_X1 U5120 ( .A1(n7563), .A2(n7562), .ZN(n8397) );
  AOI21_X1 U5121 ( .B1(n4571), .B2(n4570), .A(n4326), .ZN(n4569) );
  INV_X1 U5122 ( .A(n4577), .ZN(n4570) );
  INV_X1 U5123 ( .A(n7969), .ZN(n4740) );
  NAND2_X1 U5124 ( .A1(n8192), .A2(n4741), .ZN(n8181) );
  OR2_X1 U5125 ( .A1(n8215), .A2(n8414), .ZN(n8199) );
  OR2_X1 U5126 ( .A1(n8419), .A2(n7773), .ZN(n8194) );
  AND2_X1 U5127 ( .A1(n8194), .A2(n7960), .ZN(n8211) );
  INV_X1 U5128 ( .A(n8211), .ZN(n8207) );
  NAND2_X1 U5129 ( .A1(n8229), .A2(n8242), .ZN(n4608) );
  NAND2_X1 U5130 ( .A1(n4761), .A2(n4760), .ZN(n8230) );
  AND2_X1 U5131 ( .A1(n7958), .A2(n7961), .ZN(n8231) );
  NAND2_X1 U5132 ( .A1(n8429), .A2(n4606), .ZN(n4609) );
  OR2_X1 U5133 ( .A1(n8240), .A2(n8250), .ZN(n4761) );
  NAND2_X1 U5134 ( .A1(n4743), .A2(n4742), .ZN(n8263) );
  AND2_X1 U5135 ( .A1(n8264), .A2(n4308), .ZN(n4742) );
  AOI21_X1 U5136 ( .B1(n4595), .B2(n4592), .A(n4324), .ZN(n4591) );
  INV_X1 U5137 ( .A(n4599), .ZN(n4592) );
  INV_X1 U5138 ( .A(n4595), .ZN(n4593) );
  AND3_X1 U5139 ( .A1(n6054), .A2(n6053), .A3(n6052), .ZN(n8277) );
  NOR2_X1 U5140 ( .A1(n8293), .A2(n4600), .ZN(n4599) );
  INV_X1 U5141 ( .A(n7593), .ZN(n4600) );
  OAI22_X1 U5142 ( .A1(n8293), .A2(n4598), .B1(n8277), .B2(n8291), .ZN(n4597)
         );
  INV_X1 U5143 ( .A(n7592), .ZN(n4598) );
  NAND2_X1 U5144 ( .A1(n8292), .A2(n8293), .ZN(n8299) );
  AND2_X1 U5145 ( .A1(n8451), .A2(n8011), .ZN(n7592) );
  OR2_X1 U5146 ( .A1(n8307), .A2(n8451), .ZN(n8305) );
  OR2_X1 U5147 ( .A1(n8394), .A2(n7799), .ZN(n7182) );
  AOI21_X1 U5148 ( .B1(n7525), .B2(n4402), .A(n7524), .ZN(n8345) );
  NAND2_X1 U5149 ( .A1(n8345), .A2(n4409), .ZN(n8347) );
  AND4_X1 U5150 ( .A1(n5988), .A2(n5987), .A3(n5986), .A4(n5985), .ZN(n8331)
         );
  NAND2_X1 U5151 ( .A1(n4726), .A2(n8015), .ZN(n4725) );
  AND2_X1 U5152 ( .A1(n7909), .A2(n7439), .ZN(n7811) );
  INV_X1 U5153 ( .A(n4581), .ZN(n4580) );
  OAI21_X1 U5154 ( .B1(n7275), .B2(n4582), .A(n7819), .ZN(n4581) );
  NAND2_X1 U5155 ( .A1(n4583), .A2(n7275), .ZN(n7340) );
  AND4_X1 U5156 ( .A1(n5869), .A2(n5868), .A3(n5867), .A4(n5866), .ZN(n7256)
         );
  INV_X1 U5157 ( .A(n8372), .ZN(n8266) );
  NAND2_X1 U5158 ( .A1(n8376), .A2(n8374), .ZN(n7200) );
  NAND2_X1 U5159 ( .A1(n7585), .A2(n7180), .ZN(n7209) );
  AND2_X1 U5160 ( .A1(n8471), .A2(n7179), .ZN(n7180) );
  OR2_X1 U5161 ( .A1(n6516), .A2(n6752), .ZN(n8371) );
  NAND2_X1 U5162 ( .A1(n6168), .A2(n6167), .ZN(n8402) );
  NAND2_X1 U5163 ( .A1(n6154), .A2(n6153), .ZN(n8407) );
  NAND2_X1 U5164 ( .A1(n6108), .A2(n6107), .ZN(n8422) );
  NAND2_X1 U5165 ( .A1(n6047), .A2(n6046), .ZN(n8445) );
  AND3_X1 U5166 ( .A1(n5810), .A2(n5809), .A3(n5808), .ZN(n9750) );
  INV_X1 U5167 ( .A(n7751), .ZN(n9729) );
  OR2_X1 U5168 ( .A1(n7999), .A2(n7177), .ZN(n8473) );
  NOR2_X1 U5169 ( .A1(n8392), .A2(n8391), .ZN(n8475) );
  INV_X1 U5170 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4756) );
  INV_X1 U5171 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5714) );
  AND2_X1 U5172 ( .A1(n5846), .A2(n5828), .ZN(n6729) );
  NAND2_X1 U5173 ( .A1(n5295), .A2(n5294), .ZN(n7311) );
  NAND2_X1 U5174 ( .A1(n5000), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5394) );
  INV_X1 U5175 ( .A(n5374), .ZN(n5000) );
  NAND2_X1 U5176 ( .A1(n4385), .A2(n4384), .ZN(n4764) );
  INV_X1 U5177 ( .A(n5489), .ZN(n4384) );
  NAND2_X1 U5178 ( .A1(n5490), .A2(n8574), .ZN(n4385) );
  NAND2_X1 U5179 ( .A1(n4996), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5236) );
  AND2_X1 U5180 ( .A1(n5059), .A2(n5058), .ZN(n5060) );
  NAND2_X1 U5181 ( .A1(n5208), .A2(n4297), .ZN(n5059) );
  NAND2_X1 U5182 ( .A1(n5002), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5432) );
  OR2_X1 U5183 ( .A1(n5432), .A2(n8568), .ZN(n5452) );
  OR2_X1 U5184 ( .A1(n5310), .A2(n4782), .ZN(n4781) );
  INV_X1 U5185 ( .A(n5314), .ZN(n4782) );
  AND2_X1 U5186 ( .A1(n5289), .A2(n5314), .ZN(n4783) );
  OR2_X1 U5187 ( .A1(n5452), .A2(n5451), .ZN(n5471) );
  NAND2_X1 U5188 ( .A1(n4762), .A2(n4322), .ZN(n5269) );
  NAND2_X1 U5189 ( .A1(n5103), .A2(n5104), .ZN(n5107) );
  AND3_X1 U5190 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5173) );
  OAI21_X1 U5191 ( .B1(n4506), .B2(n4505), .A(n4501), .ZN(n8777) );
  NAND2_X1 U5192 ( .A1(n8832), .A2(n8828), .ZN(n4505) );
  INV_X1 U5193 ( .A(n4502), .ZN(n4501) );
  AND3_X1 U5194 ( .A1(n5045), .A2(n5044), .A3(n5043), .ZN(n8647) );
  NOR2_X1 U5195 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4958) );
  NOR2_X1 U5196 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4957) );
  AOI21_X1 U5197 ( .B1(n6397), .B2(n4457), .A(n4460), .ZN(n4456) );
  INV_X1 U5198 ( .A(n6395), .ZN(n4457) );
  OR2_X1 U5199 ( .A1(n6394), .A2(n4458), .ZN(n4455) );
  INV_X1 U5200 ( .A(n6397), .ZN(n4458) );
  NAND2_X1 U5201 ( .A1(n9609), .A2(n7140), .ZN(n8893) );
  AND2_X1 U5202 ( .A1(n5585), .A2(n5584), .ZN(n9024) );
  OR2_X1 U5203 ( .A1(n9040), .A2(n9046), .ZN(n4699) );
  NAND2_X1 U5204 ( .A1(n9118), .A2(n4475), .ZN(n9057) );
  NOR2_X1 U5205 ( .A1(n4477), .A2(n9267), .ZN(n4475) );
  INV_X1 U5206 ( .A(n4670), .ZN(n9056) );
  OAI21_X1 U5207 ( .B1(n9098), .B2(n4672), .A(n4671), .ZN(n4670) );
  AOI21_X1 U5208 ( .B1(n4674), .B2(n9079), .A(n8973), .ZN(n4671) );
  NAND2_X1 U5209 ( .A1(n9079), .A2(n4678), .ZN(n4672) );
  NAND2_X1 U5210 ( .A1(n4825), .A2(n4824), .ZN(n9107) );
  INV_X1 U5211 ( .A(n9109), .ZN(n4825) );
  NOR2_X1 U5212 ( .A1(n9144), .A2(n9294), .ZN(n9137) );
  NOR2_X1 U5213 ( .A1(n9133), .A2(n4818), .ZN(n4817) );
  INV_X1 U5214 ( .A(n8992), .ZN(n4818) );
  NAND2_X1 U5215 ( .A1(n9164), .A2(n8991), .ZN(n4819) );
  NOR2_X1 U5216 ( .A1(n4724), .A2(n4720), .ZN(n4719) );
  INV_X1 U5217 ( .A(n4722), .ZN(n4720) );
  AND2_X1 U5218 ( .A1(n8747), .A2(n9149), .ZN(n9166) );
  NAND2_X1 U5219 ( .A1(n4342), .A2(n4722), .ZN(n4718) );
  NAND2_X1 U5220 ( .A1(n4723), .A2(n4313), .ZN(n4721) );
  NAND2_X1 U5221 ( .A1(n8986), .A2(n4806), .ZN(n4805) );
  NOR2_X1 U5222 ( .A1(n8987), .A2(n4807), .ZN(n4806) );
  INV_X1 U5223 ( .A(n8985), .ZN(n4807) );
  OR2_X1 U5224 ( .A1(n9223), .A2(n9319), .ZN(n9212) );
  OR2_X1 U5225 ( .A1(n8651), .A2(n8987), .ZN(n9189) );
  OAI21_X1 U5226 ( .B1(n7305), .B2(n4803), .A(n4801), .ZN(n9205) );
  INV_X1 U5227 ( .A(n4802), .ZN(n4801) );
  OAI21_X1 U5228 ( .B1(n4303), .B2(n4803), .A(n8983), .ZN(n4802) );
  INV_X1 U5229 ( .A(n8981), .ZN(n4803) );
  NAND2_X1 U5230 ( .A1(n7305), .A2(n4303), .ZN(n8982) );
  INV_X1 U5231 ( .A(n4312), .ZN(n4689) );
  INV_X1 U5232 ( .A(n7312), .ZN(n4685) );
  NAND2_X1 U5233 ( .A1(n4831), .A2(n8670), .ZN(n4830) );
  NAND2_X1 U5234 ( .A1(n6924), .A2(n4305), .ZN(n4827) );
  AND4_X1 U5235 ( .A1(n5263), .A2(n5262), .A3(n5261), .A4(n5260), .ZN(n6996)
         );
  OR2_X1 U5236 ( .A1(n8683), .A2(n6925), .ZN(n8759) );
  NAND2_X1 U5237 ( .A1(n4707), .A2(n6843), .ZN(n6928) );
  INV_X1 U5238 ( .A(n6844), .ZN(n4707) );
  NAND2_X1 U5239 ( .A1(n6579), .A2(n4318), .ZN(n6643) );
  AND2_X1 U5240 ( .A1(n9488), .A2(n6445), .ZN(n9232) );
  INV_X1 U5241 ( .A(n9231), .ZN(n9392) );
  AND2_X1 U5242 ( .A1(n6447), .A2(n6446), .ZN(n9208) );
  INV_X1 U5243 ( .A(n9232), .ZN(n9394) );
  AND2_X1 U5244 ( .A1(n4483), .A2(n4482), .ZN(n9251) );
  NAND2_X1 U5245 ( .A1(n5577), .A2(n5576), .ZN(n9262) );
  NAND2_X1 U5246 ( .A1(n5497), .A2(n5496), .ZN(n9278) );
  INV_X1 U5247 ( .A(n5338), .ZN(n4510) );
  NAND2_X1 U5248 ( .A1(n5275), .A2(n5274), .ZN(n7012) );
  INV_X1 U5249 ( .A(n6993), .ZN(n7112) );
  NAND2_X1 U5250 ( .A1(n5233), .A2(n5232), .ZN(n6970) );
  NAND2_X1 U5251 ( .A1(n4634), .A2(n4941), .ZN(n5448) );
  NAND2_X1 U5252 ( .A1(n4648), .A2(n4917), .ZN(n5368) );
  OR2_X1 U5253 ( .A1(n5351), .A2(n5350), .ZN(n4648) );
  NAND2_X1 U5254 ( .A1(n4868), .A2(n4867), .ZN(n5167) );
  NAND2_X1 U5255 ( .A1(n4625), .A2(n4624), .ZN(n5133) );
  AOI21_X1 U5256 ( .B1(n4626), .B2(n5119), .A(n4337), .ZN(n4624) );
  XNOR2_X1 U5257 ( .A(n4857), .B(SI_3_), .ZN(n5119) );
  AND4_X1 U5258 ( .A1(n5839), .A2(n5838), .A3(n5837), .A4(n5836), .ZN(n7453)
         );
  OAI21_X1 U5259 ( .B1(n7692), .B2(n4541), .A(n4539), .ZN(n7632) );
  XOR2_X1 U5260 ( .A(n6115), .B(n6116), .Z(n7641) );
  NAND2_X1 U5261 ( .A1(n5710), .A2(n5709), .ZN(n8427) );
  NAND2_X1 U5262 ( .A1(n4537), .A2(n4535), .ZN(n6219) );
  AOI21_X1 U5263 ( .B1(n4539), .B2(n4541), .A(n4536), .ZN(n4535) );
  INV_X1 U5264 ( .A(n6166), .ZN(n4536) );
  INV_X1 U5265 ( .A(n7066), .ZN(n4551) );
  OAI211_X1 U5266 ( .C1(n6700), .C2(n6737), .A(n5731), .B(n5730), .ZN(n7673)
         );
  NAND2_X1 U5267 ( .A1(n6073), .A2(n4546), .ZN(n6096) );
  NOR2_X1 U5268 ( .A1(n4306), .A2(n4355), .ZN(n4546) );
  NAND2_X1 U5269 ( .A1(n7155), .A2(n5805), .ZN(n6939) );
  NAND2_X1 U5270 ( .A1(n6234), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9693) );
  OR3_X1 U5271 ( .A1(n6226), .A2(n9790), .A3(n6699), .ZN(n9431) );
  INV_X1 U5272 ( .A(n7790), .ZN(n9682) );
  INV_X1 U5273 ( .A(n8022), .ZN(n7411) );
  NAND2_X1 U5274 ( .A1(n6211), .A2(n9790), .ZN(n9687) );
  AOI21_X1 U5275 ( .B1(n4613), .B2(n7799), .A(n4612), .ZN(n7993) );
  NAND2_X1 U5276 ( .A1(n6858), .A2(n8395), .ZN(n7997) );
  NAND2_X1 U5277 ( .A1(n6160), .A2(n6159), .ZN(n8007) );
  INV_X1 U5278 ( .A(n7773), .ZN(n8233) );
  INV_X1 U5279 ( .A(n6737), .ZN(n9370) );
  AND2_X1 U5280 ( .A1(n6518), .A2(n6517), .ZN(n8151) );
  INV_X1 U5281 ( .A(n4431), .ZN(n8388) );
  AND2_X1 U5282 ( .A1(n7805), .A2(n4434), .ZN(n4433) );
  NOR3_X1 U5283 ( .A1(n8159), .A2(n7805), .A3(n4434), .ZN(n4432) );
  OAI21_X1 U5284 ( .B1(n4576), .B2(n4569), .A(n4567), .ZN(n4566) );
  NAND2_X1 U5285 ( .A1(n4568), .A2(n4569), .ZN(n4567) );
  NAND2_X1 U5286 ( .A1(n7839), .A2(n4572), .ZN(n4568) );
  INV_X1 U5287 ( .A(n8402), .ZN(n8164) );
  OR2_X1 U5288 ( .A1(n5722), .A2(n5721), .ZN(n5723) );
  OR2_X1 U5289 ( .A1(n7999), .A2(n8389), .ZN(n8218) );
  INV_X1 U5290 ( .A(n8321), .ZN(n8252) );
  AND4_X1 U5291 ( .A1(n5326), .A2(n5325), .A3(n5324), .A4(n5323), .ZN(n7314)
         );
  OR2_X1 U5292 ( .A1(n5651), .A2(n4773), .ZN(n4386) );
  OR2_X1 U5293 ( .A1(n5650), .A2(n8619), .ZN(n4773) );
  AND4_X1 U5294 ( .A1(n5362), .A2(n5361), .A3(n5360), .A4(n5359), .ZN(n9210)
         );
  NAND2_X1 U5295 ( .A1(n5393), .A2(n5392), .ZN(n9312) );
  INV_X1 U5296 ( .A(n5127), .ZN(n4766) );
  NAND2_X1 U5297 ( .A1(n5431), .A2(n5430), .ZN(n9297) );
  AND4_X1 U5298 ( .A1(n5302), .A2(n5301), .A3(n5300), .A4(n5299), .ZN(n7327)
         );
  INV_X1 U5299 ( .A(n6641), .ZN(n6634) );
  AND2_X1 U5300 ( .A1(n8596), .A2(n8592), .ZN(n5567) );
  AND2_X1 U5301 ( .A1(n6323), .A2(n5649), .ZN(n8595) );
  INV_X1 U5302 ( .A(n9228), .ZN(n9322) );
  NAND2_X1 U5303 ( .A1(n5506), .A2(n5505), .ZN(n9113) );
  NAND2_X1 U5304 ( .A1(n5026), .A2(n5025), .ZN(n9126) );
  OR2_X1 U5305 ( .A1(n9102), .A2(n5658), .ZN(n5026) );
  NAND2_X1 U5306 ( .A1(n5479), .A2(n5478), .ZN(n9106) );
  OR2_X1 U5307 ( .A1(n9120), .A2(n5658), .ZN(n5479) );
  INV_X1 U5308 ( .A(n7314), .ZN(n8878) );
  XNOR2_X1 U5309 ( .A(n8893), .B(n8900), .ZN(n7142) );
  NOR2_X1 U5310 ( .A1(n7142), .A2(n7141), .ZN(n8894) );
  AOI21_X1 U5311 ( .B1(n9354), .B2(n5229), .A(n8632), .ZN(n8945) );
  AOI21_X1 U5312 ( .B1(n4697), .B2(n9046), .A(n4358), .ZN(n4696) );
  INV_X1 U5313 ( .A(n5011), .ZN(n5014) );
  MUX2_X1 U5314 ( .A(n8668), .B(n8667), .S(n8738), .Z(n8682) );
  NAND2_X1 U5315 ( .A1(n4424), .A2(n4423), .ZN(n7888) );
  NOR2_X1 U5316 ( .A1(n7878), .A2(n7877), .ZN(n4423) );
  NAND2_X1 U5317 ( .A1(n4497), .A2(n4325), .ZN(n8705) );
  AND2_X1 U5318 ( .A1(n4407), .A2(n4399), .ZN(n4398) );
  MUX2_X1 U5319 ( .A(n8714), .B(n8713), .S(n8741), .Z(n8721) );
  AND2_X1 U5320 ( .A1(n4416), .A2(n4413), .ZN(n4412) );
  AND2_X1 U5321 ( .A1(n8211), .A2(n7961), .ZN(n4416) );
  INV_X1 U5322 ( .A(n4314), .ZN(n4414) );
  OR2_X1 U5323 ( .A1(n7941), .A2(n4415), .ZN(n4410) );
  NAND2_X1 U5324 ( .A1(n4417), .A2(n4320), .ZN(n4415) );
  INV_X1 U5325 ( .A(n7811), .ZN(n7343) );
  INV_X1 U5326 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5715) );
  INV_X1 U5327 ( .A(n4705), .ZN(n4702) );
  INV_X1 U5328 ( .A(n7545), .ZN(n4632) );
  INV_X1 U5329 ( .A(n7540), .ZN(n4629) );
  NAND2_X1 U5330 ( .A1(n4973), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4990) );
  AND2_X1 U5331 ( .A1(n4694), .A2(n4972), .ZN(n4465) );
  NAND2_X1 U5332 ( .A1(n4494), .A2(n4492), .ZN(n4635) );
  NOR2_X1 U5333 ( .A1(n4896), .A2(n4496), .ZN(n4495) );
  INV_X1 U5334 ( .A(n4891), .ZN(n4496) );
  NOR2_X1 U5335 ( .A1(n5191), .A2(n4618), .ZN(n4617) );
  INV_X1 U5336 ( .A(n5168), .ZN(n4618) );
  INV_X1 U5337 ( .A(n4871), .ZN(n4620) );
  AND2_X1 U5338 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5813) );
  OR2_X1 U5339 ( .A1(n8471), .A2(n7178), .ZN(n6230) );
  INV_X1 U5340 ( .A(n7775), .ZN(n4544) );
  AOI21_X1 U5341 ( .B1(n4394), .B2(n4395), .A(n7986), .ZN(n4393) );
  INV_X1 U5342 ( .A(n4311), .ZN(n4738) );
  INV_X1 U5343 ( .A(n6031), .ZN(n4559) );
  NOR2_X1 U5344 ( .A1(n4591), .A2(n8264), .ZN(n4590) );
  NOR2_X1 U5345 ( .A1(n8434), .A2(n7597), .ZN(n7598) );
  NOR2_X1 U5346 ( .A1(n8427), .A2(n8434), .ZN(n4445) );
  AND2_X1 U5347 ( .A1(n8375), .A2(n7201), .ZN(n7192) );
  NAND2_X1 U5348 ( .A1(n7201), .A2(n7193), .ZN(n7194) );
  OR2_X1 U5349 ( .A1(n8366), .A2(n8367), .ZN(n7401) );
  INV_X1 U5350 ( .A(n8375), .ZN(n7860) );
  NAND2_X1 U5351 ( .A1(n8024), .A2(n9734), .ZN(n7866) );
  NOR2_X1 U5352 ( .A1(n7673), .A2(n7586), .ZN(n7293) );
  NOR2_X1 U5353 ( .A1(n8419), .A2(n4442), .ZN(n4441) );
  INV_X1 U5354 ( .A(n4443), .ZN(n4442) );
  AND2_X1 U5355 ( .A1(n4747), .A2(n7227), .ZN(n4746) );
  AND2_X1 U5356 ( .A1(n7880), .A2(n7879), .ZN(n7230) );
  OAI21_X1 U5357 ( .B1(n6203), .B2(n6202), .A(n9706), .ZN(n8390) );
  INV_X1 U5358 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U5359 ( .A1(n6181), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6206) );
  INV_X1 U5360 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6205) );
  AND2_X1 U5361 ( .A1(n5715), .A2(n4558), .ZN(n4557) );
  INV_X1 U5362 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4558) );
  NOR2_X1 U5363 ( .A1(n5908), .A2(n4549), .ZN(n5939) );
  NAND2_X1 U5364 ( .A1(n5876), .A2(n4426), .ZN(n5908) );
  NAND2_X1 U5365 ( .A1(n5876), .A2(n5877), .ZN(n5896) );
  NOR2_X1 U5366 ( .A1(n8740), .A2(n8739), .ZN(n4508) );
  OR2_X1 U5367 ( .A1(n8735), .A2(n8734), .ZN(n8736) );
  NOR2_X1 U5368 ( .A1(n8861), .A2(n8738), .ZN(n4507) );
  OAI211_X1 U5369 ( .C1(n8742), .C2(n8741), .A(n4503), .B(n8743), .ZN(n4502)
         );
  NAND2_X1 U5370 ( .A1(n4321), .A2(n4504), .ZN(n4503) );
  INV_X1 U5371 ( .A(n8828), .ZN(n4504) );
  NOR2_X1 U5372 ( .A1(n7138), .A2(n4461), .ZN(n7139) );
  AND2_X1 U5373 ( .A1(n7145), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4461) );
  OR2_X1 U5374 ( .A1(n9262), .A2(n9024), .ZN(n9001) );
  OR2_X1 U5375 ( .A1(n9267), .A2(n9080), .ZN(n8974) );
  NOR2_X1 U5376 ( .A1(n9278), .A2(n9282), .ZN(n4478) );
  NAND2_X1 U5377 ( .A1(n4474), .A2(n9163), .ZN(n4473) );
  NOR2_X1 U5378 ( .A1(n9308), .A2(n9312), .ZN(n4474) );
  NAND2_X1 U5379 ( .A1(n4999), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5357) );
  NAND2_X1 U5380 ( .A1(n7315), .A2(n8689), .ZN(n7316) );
  NOR2_X1 U5381 ( .A1(n7015), .A2(n7311), .ZN(n7315) );
  AND2_X1 U5382 ( .A1(n6656), .A2(n4466), .ZN(n7002) );
  AND2_X1 U5383 ( .A1(n4467), .A2(n9417), .ZN(n4466) );
  NOR2_X1 U5384 ( .A1(n4468), .A2(n7112), .ZN(n4467) );
  INV_X1 U5385 ( .A(n4469), .ZN(n4468) );
  NOR2_X1 U5386 ( .A1(n6840), .A2(n6970), .ZN(n4469) );
  NAND2_X1 U5387 ( .A1(n5197), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5234) );
  INV_X1 U5388 ( .A(n4810), .ZN(n4811) );
  XNOR2_X1 U5389 ( .A(n6457), .B(n6456), .ZN(n8752) );
  NAND3_X1 U5390 ( .A1(n4970), .A2(n4988), .A3(n4985), .ZN(n4971) );
  INV_X1 U5391 ( .A(n4657), .ZN(n4656) );
  AOI21_X1 U5392 ( .B1(n4657), .B2(n4659), .A(n4655), .ZN(n4654) );
  AND2_X1 U5393 ( .A1(n5601), .A2(n5574), .ZN(n5599) );
  INV_X1 U5394 ( .A(n5521), .ZN(n4661) );
  AOI21_X1 U5395 ( .B1(n5517), .B2(n4660), .A(n4658), .ZN(n4657) );
  INV_X1 U5396 ( .A(n5541), .ZN(n4658) );
  NAND2_X1 U5397 ( .A1(n4799), .A2(n4969), .ZN(n4982) );
  OAI21_X1 U5398 ( .B1(n5410), .B2(n5409), .A(n4936), .ZN(n5429) );
  AND2_X1 U5399 ( .A1(n4941), .A2(n4940), .ZN(n5428) );
  INV_X1 U5400 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4962) );
  INV_X1 U5401 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4963) );
  INV_X1 U5402 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4964) );
  INV_X1 U5403 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n4959) );
  NAND2_X1 U5404 ( .A1(n4643), .A2(n4642), .ZN(n5032) );
  AOI21_X1 U5405 ( .B1(n4645), .B2(n4647), .A(n4360), .ZN(n4642) );
  INV_X1 U5406 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5335) );
  NOR2_X1 U5407 ( .A1(n5253), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5272) );
  INV_X1 U5408 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5192) );
  OAI21_X1 U5409 ( .B1(n7554), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n4860), .ZN(
        n4861) );
  NAND2_X1 U5410 ( .A1(n7554), .A2(n6249), .ZN(n4860) );
  NAND2_X1 U5411 ( .A1(n4665), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4664) );
  AND2_X1 U5412 ( .A1(n6166), .A2(n6165), .ZN(n7629) );
  OR2_X1 U5413 ( .A1(n5964), .A2(n5963), .ZN(n5989) );
  AND2_X1 U5414 ( .A1(n4540), .A2(n7629), .ZN(n4539) );
  OR2_X1 U5415 ( .A1(n4543), .A2(n4541), .ZN(n4540) );
  NAND2_X1 U5416 ( .A1(n4542), .A2(n6152), .ZN(n4541) );
  INV_X1 U5417 ( .A(n6088), .ZN(n6086) );
  AND2_X1 U5418 ( .A1(n6699), .A2(n7997), .ZN(n7177) );
  INV_X1 U5419 ( .A(n8473), .ZN(n7585) );
  OR2_X1 U5420 ( .A1(n6037), .A2(n7713), .ZN(n6039) );
  AND2_X1 U5421 ( .A1(n7691), .A2(n4544), .ZN(n4543) );
  NAND2_X1 U5422 ( .A1(n4544), .A2(n6136), .ZN(n4542) );
  OAI21_X1 U5423 ( .B1(n7798), .B2(n7797), .A(n7983), .ZN(n7802) );
  XNOR2_X1 U5424 ( .A(n4614), .B(n8219), .ZN(n4613) );
  NOR2_X1 U5425 ( .A1(n7839), .A2(n7832), .ZN(n4615) );
  NOR2_X1 U5426 ( .A1(n7833), .A2(n8394), .ZN(n4612) );
  INV_X1 U5427 ( .A(n4298), .ZN(n6411) );
  AND4_X1 U5428 ( .A1(n5890), .A2(n5889), .A3(n5888), .A4(n5887), .ZN(n7277)
         );
  NOR2_X1 U5429 ( .A1(n9367), .A2(n9368), .ZN(n9366) );
  NOR2_X1 U5430 ( .A1(n8062), .A2(n8063), .ZN(n8061) );
  AND2_X1 U5431 ( .A1(n4515), .A2(n4514), .ZN(n6784) );
  NAND2_X1 U5432 ( .A1(n6724), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4514) );
  NOR2_X1 U5433 ( .A1(n6782), .A2(n4519), .ZN(n6718) );
  NOR2_X1 U5434 ( .A1(n4521), .A2(n4520), .ZN(n4519) );
  NOR2_X1 U5435 ( .A1(n6718), .A2(n6717), .ZN(n6824) );
  NOR2_X1 U5436 ( .A1(n6824), .A2(n4518), .ZN(n6826) );
  AND2_X1 U5437 ( .A1(n6825), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4518) );
  NOR2_X1 U5438 ( .A1(n6826), .A2(n6827), .ZN(n6871) );
  NOR2_X1 U5439 ( .A1(n8084), .A2(n8083), .ZN(n8086) );
  NOR2_X1 U5440 ( .A1(n8121), .A2(n4378), .ZN(n8125) );
  NAND2_X1 U5441 ( .A1(n8125), .A2(n8124), .ZN(n8137) );
  NAND2_X1 U5442 ( .A1(n4436), .A2(n4435), .ZN(n4434) );
  INV_X1 U5443 ( .A(n8397), .ZN(n4435) );
  OR2_X1 U5444 ( .A1(n8159), .A2(n8397), .ZN(n8153) );
  NAND2_X1 U5445 ( .A1(n8182), .A2(n4577), .ZN(n4573) );
  OR2_X1 U5446 ( .A1(n6171), .A2(n6170), .ZN(n7612) );
  AND2_X1 U5447 ( .A1(n7835), .A2(n7834), .ZN(n8157) );
  OR2_X1 U5448 ( .A1(n8407), .A2(n8007), .ZN(n4577) );
  NOR2_X1 U5449 ( .A1(n8199), .A2(n8407), .ZN(n8177) );
  AND2_X1 U5450 ( .A1(n7967), .A2(n7969), .ZN(n8193) );
  INV_X1 U5451 ( .A(n4602), .ZN(n4601) );
  OAI22_X1 U5452 ( .A1(n8211), .A2(n4608), .B1(n8233), .B2(n8419), .ZN(n4602)
         );
  AOI21_X1 U5453 ( .B1(n4760), .B2(n8250), .A(n4759), .ZN(n4758) );
  INV_X1 U5454 ( .A(n7958), .ZN(n4759) );
  NAND2_X1 U5455 ( .A1(n8279), .A2(n4445), .ZN(n8244) );
  AND2_X1 U5456 ( .A1(n8287), .A2(n7595), .ZN(n8279) );
  NAND2_X1 U5457 ( .A1(n8279), .A2(n8262), .ZN(n8256) );
  INV_X1 U5458 ( .A(n6050), .ZN(n6048) );
  NOR2_X1 U5459 ( .A1(n8305), .A2(n8445), .ZN(n8287) );
  AND2_X1 U5460 ( .A1(n7947), .A2(n7934), .ZN(n8313) );
  NOR2_X1 U5461 ( .A1(n8355), .A2(n8462), .ZN(n4438) );
  NOR3_X1 U5462 ( .A1(n8355), .A2(n8462), .A3(n8455), .ZN(n4439) );
  INV_X1 U5463 ( .A(n4585), .ZN(n4584) );
  OAI21_X1 U5464 ( .B1(n4409), .B2(n4304), .A(n4587), .ZN(n4585) );
  OR2_X1 U5465 ( .A1(n8462), .A2(n8012), .ZN(n4587) );
  AND2_X1 U5466 ( .A1(n7945), .A2(n7935), .ZN(n7533) );
  AND4_X1 U5467 ( .A1(n5995), .A2(n5994), .A3(n5993), .A4(n5992), .ZN(n8344)
         );
  INV_X1 U5468 ( .A(n4382), .ZN(n7499) );
  OAI21_X1 U5469 ( .B1(n7445), .B2(n7913), .A(n4383), .ZN(n4382) );
  NAND2_X1 U5470 ( .A1(n7466), .A2(n7446), .ZN(n4383) );
  NAND2_X1 U5471 ( .A1(n7366), .A2(n7342), .ZN(n7344) );
  AND4_X1 U5472 ( .A1(n5918), .A2(n5917), .A3(n5916), .A4(n5915), .ZN(n7488)
         );
  AND4_X1 U5473 ( .A1(n4428), .A2(n9769), .A3(n4427), .A4(n7456), .ZN(n7282)
         );
  AND4_X1 U5474 ( .A1(n5905), .A2(n5904), .A3(n5903), .A4(n5902), .ZN(n7467)
         );
  NAND2_X1 U5475 ( .A1(n4372), .A2(n4428), .ZN(n7261) );
  NAND2_X1 U5476 ( .A1(n7456), .A2(n9755), .ZN(n7246) );
  AND4_X1 U5477 ( .A1(n5784), .A2(n5783), .A3(n5782), .A4(n5781), .ZN(n7412)
         );
  OR2_X1 U5478 ( .A1(n5834), .A2(n5780), .ZN(n5782) );
  NAND2_X1 U5479 ( .A1(n7293), .A2(n9729), .ZN(n8366) );
  NAND2_X1 U5480 ( .A1(n6138), .A2(n6137), .ZN(n8414) );
  INV_X1 U5481 ( .A(n9801), .ZN(n9791) );
  INV_X1 U5482 ( .A(n9790), .ZN(n9799) );
  INV_X1 U5483 ( .A(n7999), .ZN(n9708) );
  NAND2_X1 U5484 ( .A1(n6206), .A2(n6205), .ZN(n6208) );
  AND3_X1 U5485 ( .A1(n5958), .A2(n5955), .A3(n5712), .ZN(n5713) );
  AND2_X1 U5486 ( .A1(n5960), .A2(n5996), .ZN(n8073) );
  NOR2_X1 U5487 ( .A1(n4730), .A2(n4729), .ZN(n5806) );
  AND2_X1 U5488 ( .A1(n4733), .A2(n4734), .ZN(n4732) );
  INV_X1 U5489 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5976) );
  OAI21_X1 U5490 ( .B1(n4846), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n4663), .ZN(
        n4848) );
  NAND2_X1 U5491 ( .A1(n4668), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4663) );
  NAND2_X1 U5492 ( .A1(n5349), .A2(n5348), .ZN(n7168) );
  NAND2_X1 U5493 ( .A1(n4793), .A2(n8584), .ZN(n4792) );
  AND2_X1 U5494 ( .A1(n5593), .A2(n5592), .ZN(n5650) );
  NAND2_X1 U5495 ( .A1(n4998), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5321) );
  INV_X1 U5496 ( .A(n5297), .ZN(n4998) );
  OR2_X1 U5497 ( .A1(n5499), .A2(n5498), .ZN(n5530) );
  NAND2_X1 U5498 ( .A1(n4771), .A2(n4770), .ZN(n4769) );
  INV_X1 U5499 ( .A(n5125), .ZN(n4770) );
  INV_X1 U5500 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5220) );
  NOR2_X1 U5501 ( .A1(n8516), .A2(n4788), .ZN(n4787) );
  INV_X1 U5502 ( .A(n4792), .ZN(n4788) );
  INV_X1 U5503 ( .A(n8516), .ZN(n4785) );
  NAND2_X1 U5504 ( .A1(n4791), .A2(n4790), .ZN(n4789) );
  NAND2_X1 U5505 ( .A1(n4334), .A2(n4838), .ZN(n4790) );
  NAND2_X1 U5506 ( .A1(n4794), .A2(n4796), .ZN(n4791) );
  INV_X1 U5507 ( .A(n5471), .ZN(n5003) );
  NAND2_X1 U5508 ( .A1(n4997), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5297) );
  INV_X1 U5509 ( .A(n5277), .ZN(n4997) );
  NAND2_X1 U5510 ( .A1(n5001), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U5511 ( .A1(n5164), .A2(n5163), .ZN(n6627) );
  AND2_X1 U5512 ( .A1(n5173), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5197) );
  AND2_X1 U5513 ( .A1(n6355), .A2(n6353), .ZN(n6323) );
  NOR2_X1 U5514 ( .A1(n9562), .A2(n4448), .ZN(n9576) );
  NOR2_X1 U5515 ( .A1(n6252), .A2(n4449), .ZN(n4448) );
  INV_X1 U5516 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n4449) );
  NAND2_X1 U5517 ( .A1(n9576), .A2(n9577), .ZN(n9575) );
  NAND2_X1 U5518 ( .A1(n6394), .A2(n6395), .ZN(n6396) );
  NOR2_X1 U5519 ( .A1(n4459), .A2(n4454), .ZN(n4453) );
  INV_X1 U5520 ( .A(n4456), .ZN(n4454) );
  INV_X1 U5521 ( .A(n6428), .ZN(n4459) );
  NOR2_X1 U5522 ( .A1(n6687), .A2(n4462), .ZN(n6691) );
  AND2_X1 U5523 ( .A1(n6688), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4462) );
  NOR2_X1 U5524 ( .A1(n6691), .A2(n6690), .ZN(n7138) );
  XNOR2_X1 U5525 ( .A(n7139), .B(n9608), .ZN(n9611) );
  NOR2_X1 U5526 ( .A1(n8925), .A2(n4377), .ZN(n9626) );
  NOR2_X1 U5527 ( .A1(n9626), .A2(n9625), .ZN(n9624) );
  OR2_X1 U5528 ( .A1(n9272), .A2(n8971), .ZN(n9062) );
  NAND2_X1 U5529 ( .A1(n4820), .A2(n4821), .ZN(n9063) );
  AOI21_X1 U5530 ( .B1(n4823), .B2(n9110), .A(n4822), .ZN(n4821) );
  INV_X1 U5531 ( .A(n8998), .ZN(n4822) );
  NAND2_X1 U5532 ( .A1(n9062), .A2(n8745), .ZN(n9079) );
  NAND2_X1 U5533 ( .A1(n4678), .A2(n4676), .ZN(n4675) );
  INV_X1 U5534 ( .A(n8968), .ZN(n4676) );
  NAND2_X1 U5535 ( .A1(n9118), .A2(n4478), .ZN(n9086) );
  NAND2_X1 U5536 ( .A1(n9118), .A2(n9105), .ZN(n9099) );
  AOI21_X1 U5537 ( .B1(n4817), .B2(n4815), .A(n4814), .ZN(n4813) );
  INV_X1 U5538 ( .A(n4817), .ZN(n4816) );
  INV_X1 U5539 ( .A(n8993), .ZN(n4814) );
  AND2_X1 U5540 ( .A1(n9137), .A2(n9123), .ZN(n9118) );
  AOI21_X1 U5541 ( .B1(n4300), .B2(n4716), .A(n4333), .ZN(n4709) );
  AND2_X1 U5542 ( .A1(n9181), .A2(n8988), .ZN(n4804) );
  NOR2_X1 U5543 ( .A1(n9212), .A2(n4472), .ZN(n9174) );
  INV_X1 U5544 ( .A(n4474), .ZN(n4472) );
  NOR2_X1 U5545 ( .A1(n9212), .A2(n9312), .ZN(n9191) );
  NOR2_X1 U5546 ( .A1(n4686), .A2(n4332), .ZN(n4681) );
  NOR2_X1 U5547 ( .A1(n8676), .A2(n4829), .ZN(n4826) );
  NAND2_X1 U5548 ( .A1(n6998), .A2(n6997), .ZN(n7014) );
  NAND2_X1 U5549 ( .A1(n4833), .A2(n4831), .ZN(n9390) );
  INV_X1 U5550 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5257) );
  OR2_X1 U5551 ( .A1(n5258), .A2(n5257), .ZN(n5277) );
  NAND2_X1 U5552 ( .A1(n4833), .A2(n8669), .ZN(n7000) );
  NAND2_X1 U5553 ( .A1(n6656), .A2(n4469), .ZN(n6932) );
  AND2_X1 U5554 ( .A1(n8669), .A2(n8820), .ZN(n8758) );
  AND4_X1 U5555 ( .A1(n5204), .A2(n5203), .A3(n5202), .A4(n5201), .ZN(n6839)
         );
  OR2_X1 U5556 ( .A1(n6653), .A2(n8755), .ZN(n6838) );
  NAND2_X1 U5557 ( .A1(n6656), .A2(n6664), .ZN(n6852) );
  NOR2_X1 U5558 ( .A1(n6587), .A2(n6634), .ZN(n6656) );
  NAND2_X1 U5559 ( .A1(n4463), .A2(n6539), .ZN(n6587) );
  OAI21_X1 U5560 ( .B1(n6485), .B2(n4810), .A(n4808), .ZN(n6647) );
  INV_X1 U5561 ( .A(n4809), .ZN(n4808) );
  AND4_X1 U5562 ( .A1(n5148), .A2(n5147), .A3(n5146), .A4(n5145), .ZN(n6538)
         );
  NAND2_X1 U5563 ( .A1(n6529), .A2(n6478), .ZN(n6490) );
  AND2_X1 U5564 ( .A1(n6596), .A2(n4464), .ZN(n6529) );
  INV_X1 U5565 ( .A(n6527), .ZN(n4464) );
  NAND2_X1 U5566 ( .A1(n6464), .A2(n6463), .ZN(n8842) );
  INV_X1 U5567 ( .A(n8752), .ZN(n6523) );
  OR2_X1 U5568 ( .A1(n5066), .A2(n9495), .ZN(n5072) );
  NAND2_X1 U5569 ( .A1(n5069), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5070) );
  OR2_X1 U5570 ( .A1(n5096), .A2(n6246), .ZN(n5071) );
  OR2_X1 U5571 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(n5010), .ZN(n5013) );
  NAND2_X1 U5572 ( .A1(n4633), .A2(n7545), .ZN(n7561) );
  NAND2_X1 U5573 ( .A1(n7541), .A2(n7540), .ZN(n4633) );
  XNOR2_X1 U5574 ( .A(n7541), .B(n7540), .ZN(n7512) );
  CLKBUF_X1 U5575 ( .A(n6284), .Z(n6285) );
  XNOR2_X1 U5576 ( .A(n5600), .B(n5599), .ZN(n7494) );
  XNOR2_X1 U5577 ( .A(n5569), .B(n5568), .ZN(n7398) );
  NAND2_X1 U5578 ( .A1(n4653), .A2(n4657), .ZN(n5569) );
  NAND2_X1 U5579 ( .A1(n5518), .A2(n4660), .ZN(n4653) );
  OAI21_X1 U5580 ( .B1(n5467), .B2(n5466), .A(n4950), .ZN(n5492) );
  AND2_X1 U5581 ( .A1(n5493), .A2(n4955), .ZN(n5491) );
  NAND2_X1 U5582 ( .A1(n4652), .A2(n4923), .ZN(n5387) );
  NAND2_X1 U5583 ( .A1(n4644), .A2(n4649), .ZN(n4652) );
  NAND2_X1 U5584 ( .A1(n5351), .A2(n4917), .ZN(n4644) );
  AND2_X1 U5585 ( .A1(n4489), .A2(n4636), .ZN(n4488) );
  OR2_X1 U5586 ( .A1(n5292), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5316) );
  OAI21_X1 U5587 ( .B1(n5291), .B2(n5290), .A(n4902), .ZN(n5315) );
  NAND2_X1 U5588 ( .A1(n4892), .A2(n4891), .ZN(n5271) );
  CLKBUF_X1 U5589 ( .A(n5033), .Z(n5034) );
  NAND2_X1 U5590 ( .A1(n4621), .A2(n4871), .ZN(n5190) );
  NAND2_X1 U5591 ( .A1(n5167), .A2(n5168), .ZN(n4621) );
  AND2_X1 U5592 ( .A1(n5155), .A2(n5154), .ZN(n6392) );
  NAND2_X1 U5593 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4452) );
  NAND2_X1 U5594 ( .A1(n7515), .A2(n5954), .ZN(n9430) );
  INV_X1 U5595 ( .A(n7338), .ZN(n9782) );
  AND2_X1 U5596 ( .A1(n6228), .A2(n6227), .ZN(n9428) );
  INV_X1 U5597 ( .A(n8367), .ZN(n9734) );
  AND4_X1 U5598 ( .A1(n6025), .A2(n6024), .A3(n6023), .A4(n6022), .ZN(n7714)
         );
  OR2_X1 U5599 ( .A1(n6117), .A2(n8009), .ZN(n6114) );
  NAND2_X1 U5600 ( .A1(n7156), .A2(n5801), .ZN(n7155) );
  NAND2_X1 U5601 ( .A1(n4555), .A2(n4553), .ZN(n7125) );
  OR2_X1 U5602 ( .A1(n5751), .A2(n4512), .ZN(n5744) );
  AND4_X1 U5603 ( .A1(n5932), .A2(n5931), .A3(n5930), .A4(n5929), .ZN(n7518)
         );
  NAND2_X1 U5604 ( .A1(n4527), .A2(n4525), .ZN(n5937) );
  NAND2_X1 U5605 ( .A1(n6096), .A2(n6098), .ZN(n4545) );
  OAI21_X1 U5606 ( .B1(n7648), .B2(n7649), .A(n4528), .ZN(n7391) );
  INV_X1 U5607 ( .A(n4530), .ZN(n4528) );
  NAND2_X1 U5608 ( .A1(n9428), .A2(n8266), .ZN(n7789) );
  INV_X1 U5609 ( .A(n9693), .ZN(n7782) );
  INV_X1 U5610 ( .A(n9431), .ZN(n9674) );
  INV_X1 U5611 ( .A(n7772), .ZN(n9678) );
  NAND2_X1 U5612 ( .A1(n5999), .A2(n5998), .ZN(n7793) );
  INV_X1 U5613 ( .A(n9687), .ZN(n9435) );
  INV_X1 U5614 ( .A(n7256), .ZN(n8020) );
  NAND4_X1 U5615 ( .A1(n5819), .A2(n5818), .A3(n5817), .A4(n5816), .ZN(n8022)
         );
  NAND2_X1 U5616 ( .A1(n7603), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5819) );
  INV_X1 U5617 ( .A(n7412), .ZN(n8024) );
  INV_X2 U5618 ( .A(P2_U3966), .ZN(n8026) );
  INV_X1 U5619 ( .A(n4523), .ZN(n8047) );
  INV_X1 U5620 ( .A(n4517), .ZN(n6760) );
  INV_X1 U5621 ( .A(n4515), .ZN(n6771) );
  INV_X1 U5622 ( .A(n8151), .ZN(n9697) );
  AND2_X1 U5623 ( .A1(n8187), .A2(n8186), .ZN(n8410) );
  NOR2_X1 U5624 ( .A1(n8196), .A2(n4740), .ZN(n8183) );
  AND2_X1 U5625 ( .A1(n4609), .A2(n4608), .ZN(n8208) );
  AND2_X1 U5626 ( .A1(n8235), .A2(n8234), .ZN(n8425) );
  AND2_X1 U5627 ( .A1(n4761), .A2(n7943), .ZN(n8232) );
  NAND2_X1 U5628 ( .A1(n8429), .A2(n7600), .ZN(n8225) );
  AND2_X1 U5629 ( .A1(n8268), .A2(n8267), .ZN(n8437) );
  OAI21_X1 U5630 ( .B1(n7594), .B2(n4593), .A(n4591), .ZN(n8255) );
  INV_X1 U5631 ( .A(n8440), .ZN(n7595) );
  NAND2_X1 U5632 ( .A1(n8299), .A2(n7948), .ZN(n8274) );
  INV_X1 U5633 ( .A(n4743), .ZN(n8273) );
  NAND2_X1 U5634 ( .A1(n4596), .A2(n4594), .ZN(n8272) );
  INV_X1 U5635 ( .A(n4597), .ZN(n4594) );
  NAND2_X1 U5636 ( .A1(n7594), .A2(n4599), .ZN(n4596) );
  AOI21_X1 U5637 ( .B1(n7594), .B2(n7593), .A(n7592), .ZN(n8286) );
  NAND2_X1 U5638 ( .A1(n8347), .A2(n4837), .ZN(n8323) );
  NAND2_X1 U5639 ( .A1(n7340), .A2(n7339), .ZN(n7476) );
  NAND2_X1 U5640 ( .A1(n7225), .A2(n7871), .ZN(n7242) );
  OR2_X1 U5641 ( .A1(n7379), .A2(n9801), .ZN(n8358) );
  INV_X1 U5642 ( .A(n8218), .ZN(n8369) );
  NOR2_X1 U5643 ( .A1(n5792), .A2(n6263), .ZN(n4610) );
  INV_X1 U5644 ( .A(n8363), .ZN(n8311) );
  INV_X1 U5645 ( .A(n8358), .ZN(n8370) );
  NAND2_X1 U5646 ( .A1(n8383), .A2(n7183), .ZN(n8321) );
  OAI21_X1 U5647 ( .B1(n8388), .B2(n9801), .A(n4331), .ZN(n8476) );
  AND2_X1 U5648 ( .A1(n4566), .A2(n9806), .ZN(n4564) );
  AND2_X2 U5649 ( .A1(n8475), .A2(n8474), .ZN(n9809) );
  NOR2_X1 U5650 ( .A1(n8473), .A2(n8472), .ZN(n8474) );
  AND2_X1 U5651 ( .A1(n6231), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9715) );
  INV_X1 U5652 ( .A(n9715), .ZN(n9710) );
  NAND2_X1 U5653 ( .A1(n5708), .A2(n5707), .ZN(n7998) );
  MUX2_X1 U5654 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5705), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5708) );
  AND2_X1 U5655 ( .A1(n6185), .A2(n5704), .ZN(n7399) );
  INV_X1 U5656 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n9922) );
  XNOR2_X1 U5657 ( .A(n6182), .B(P2_IR_REG_24__SCAN_IN), .ZN(n7133) );
  NAND2_X1 U5658 ( .A1(n6208), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6182) );
  INV_X1 U5659 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7627) );
  INV_X1 U5660 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6905) );
  NAND2_X1 U5661 ( .A1(n4301), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5718) );
  INV_X1 U5662 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6860) );
  INV_X1 U5663 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4560) );
  NAND2_X1 U5664 ( .A1(n5724), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4561) );
  INV_X1 U5665 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6804) );
  INV_X1 U5666 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6594) );
  INV_X1 U5667 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6407) );
  INV_X1 U5668 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6373) );
  INV_X1 U5669 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6343) );
  INV_X1 U5670 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6315) );
  INV_X1 U5671 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6312) );
  INV_X1 U5672 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6283) );
  INV_X1 U5673 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U5674 ( .A1(n5729), .A2(n5728), .ZN(n6737) );
  AND2_X1 U5675 ( .A1(n5616), .A2(n5615), .ZN(n9049) );
  OR2_X1 U5676 ( .A1(n5666), .A2(n5658), .ZN(n5616) );
  INV_X1 U5677 ( .A(n4764), .ZN(n8506) );
  AND4_X1 U5678 ( .A1(n5225), .A2(n5224), .A3(n5223), .A4(n5222), .ZN(n9393)
         );
  AND2_X1 U5679 ( .A1(n4769), .A2(n5127), .ZN(n6365) );
  AOI21_X1 U5680 ( .B1(n8546), .B2(n4792), .A(n4789), .ZN(n8515) );
  NAND2_X1 U5681 ( .A1(n5414), .A2(n5413), .ZN(n9302) );
  AND4_X1 U5682 ( .A1(n5131), .A2(n5130), .A3(n5129), .A4(n5128), .ZN(n6574)
         );
  AND2_X1 U5683 ( .A1(n4763), .A2(n4764), .ZN(n8557) );
  OAI211_X1 U5684 ( .C1(n6302), .C2(n6248), .A(n5136), .B(n5135), .ZN(n6560)
         );
  AND4_X1 U5685 ( .A1(n5240), .A2(n5239), .A3(n5238), .A4(n5237), .ZN(n6926)
         );
  OAI21_X1 U5686 ( .B1(n5066), .B2(n6297), .A(n5056), .ZN(n6436) );
  AND2_X1 U5687 ( .A1(n5061), .A2(n5060), .ZN(n4772) );
  NAND2_X1 U5688 ( .A1(n6948), .A2(n4783), .ZN(n4776) );
  NAND2_X1 U5689 ( .A1(n5469), .A2(n5468), .ZN(n9287) );
  INV_X1 U5690 ( .A(n8615), .ZN(n8578) );
  NAND2_X1 U5691 ( .A1(n5108), .A2(n5107), .ZN(n5109) );
  INV_X1 U5692 ( .A(n8599), .ZN(n8611) );
  OR2_X1 U5693 ( .A1(n5665), .A2(n9488), .ZN(n8599) );
  AND2_X1 U5694 ( .A1(n5607), .A2(n5552), .ZN(n9059) );
  NAND2_X1 U5695 ( .A1(n5677), .A2(n6321), .ZN(n8612) );
  OR2_X1 U5696 ( .A1(n5665), .A2(n9522), .ZN(n8615) );
  INV_X1 U5697 ( .A(n8604), .ZN(n8617) );
  INV_X1 U5698 ( .A(n8595), .ZN(n8619) );
  INV_X1 U5699 ( .A(n9488), .ZN(n9522) );
  MUX2_X1 U5700 ( .A(n8836), .B(n8835), .S(n9646), .Z(n8871) );
  AND2_X1 U5701 ( .A1(n5664), .A2(n5663), .ZN(n9023) );
  INV_X1 U5702 ( .A(n9049), .ZN(n9009) );
  NAND2_X1 U5703 ( .A1(n6267), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5074) );
  NAND2_X1 U5704 ( .A1(n9589), .A2(n9590), .ZN(n9588) );
  NAND2_X1 U5705 ( .A1(n9575), .A2(n4447), .ZN(n9589) );
  OR2_X1 U5706 ( .A1(n9571), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4447) );
  NOR2_X1 U5707 ( .A1(n8894), .A2(n8895), .ZN(n8898) );
  OR2_X1 U5708 ( .A1(n6293), .A2(n9522), .ZN(n9543) );
  XNOR2_X1 U5709 ( .A(n4450), .B(n9947), .ZN(n8936) );
  OR2_X1 U5710 ( .A1(n9624), .A2(n4451), .ZN(n4450) );
  AND2_X1 U5711 ( .A1(n9630), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4451) );
  INV_X1 U5712 ( .A(n9549), .ZN(n9635) );
  AND2_X1 U5713 ( .A1(n8624), .A2(n8623), .ZN(n9248) );
  AND2_X1 U5714 ( .A1(n9029), .A2(n8978), .ZN(n9255) );
  NAND2_X1 U5715 ( .A1(n4699), .A2(n4697), .ZN(n8978) );
  NAND2_X1 U5716 ( .A1(n4699), .A2(n8977), .ZN(n9028) );
  AND2_X1 U5717 ( .A1(n9033), .A2(n9032), .ZN(n9257) );
  AND2_X1 U5718 ( .A1(n9107), .A2(n8997), .ZN(n9093) );
  AND2_X1 U5719 ( .A1(n4679), .A2(n4680), .ZN(n9085) );
  NAND2_X1 U5720 ( .A1(n9098), .A2(n8968), .ZN(n4679) );
  INV_X1 U5721 ( .A(n9287), .ZN(n9123) );
  NAND2_X1 U5722 ( .A1(n5450), .A2(n5449), .ZN(n9294) );
  NAND2_X1 U5723 ( .A1(n4819), .A2(n8992), .ZN(n9132) );
  NAND2_X1 U5724 ( .A1(n4710), .A2(n4713), .ZN(n9143) );
  NAND2_X1 U5725 ( .A1(n9190), .A2(n4711), .ZN(n4710) );
  INV_X1 U5726 ( .A(n9302), .ZN(n9163) );
  NAND2_X1 U5727 ( .A1(n4712), .A2(n4718), .ZN(n9157) );
  NAND2_X1 U5728 ( .A1(n8960), .A2(n4719), .ZN(n4712) );
  OAI21_X1 U5729 ( .B1(n8960), .B2(n4313), .A(n4723), .ZN(n9173) );
  NAND2_X1 U5730 ( .A1(n8986), .A2(n8985), .ZN(n9197) );
  NAND2_X1 U5731 ( .A1(n5372), .A2(n5371), .ZN(n9319) );
  NAND2_X1 U5732 ( .A1(n8982), .A2(n8981), .ZN(n9230) );
  AND2_X1 U5733 ( .A1(n5356), .A2(n5355), .ZN(n9228) );
  NAND2_X1 U5734 ( .A1(n7305), .A2(n8675), .ZN(n7306) );
  NAND2_X1 U5735 ( .A1(n4683), .A2(n4690), .ZN(n8953) );
  NAND2_X1 U5736 ( .A1(n7313), .A2(n4684), .ZN(n4683) );
  NOR2_X1 U5737 ( .A1(n4689), .A2(n4685), .ZN(n4684) );
  OAI21_X1 U5738 ( .B1(n7313), .B2(n8763), .A(n7312), .ZN(n7328) );
  NAND2_X1 U5739 ( .A1(n4827), .A2(n4828), .ZN(n7009) );
  INV_X1 U5740 ( .A(n9644), .ZN(n9404) );
  NAND2_X1 U5741 ( .A1(n6928), .A2(n6927), .ZN(n6995) );
  AND2_X1 U5742 ( .A1(n5219), .A2(n5218), .ZN(n6993) );
  AND2_X1 U5743 ( .A1(n6579), .A2(n6578), .ZN(n6580) );
  AND3_X1 U5744 ( .A1(n5172), .A2(n5171), .A3(n5170), .ZN(n6641) );
  INV_X1 U5745 ( .A(n9646), .ZN(n4797) );
  NAND2_X1 U5746 ( .A1(n6659), .A2(n9644), .ZN(n9653) );
  NOR3_X1 U5747 ( .A1(n9251), .A2(n9250), .A3(n4481), .ZN(n9253) );
  AND2_X1 U5748 ( .A1(n9252), .A2(n9330), .ZN(n4481) );
  AND2_X1 U5749 ( .A1(n9657), .A2(n9656), .ZN(n9660) );
  INV_X1 U5750 ( .A(n6320), .ZN(n9657) );
  XNOR2_X1 U5751 ( .A(n7557), .B(n7556), .ZN(n9354) );
  INV_X1 U5752 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5016) );
  INV_X1 U5753 ( .A(n5018), .ZN(n9362) );
  CLKBUF_X1 U5754 ( .A(n5657), .Z(n9488) );
  INV_X1 U5755 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n9965) );
  XNOR2_X1 U5756 ( .A(n5492), .B(n5491), .ZN(n7072) );
  INV_X1 U5757 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n6981) );
  INV_X1 U5758 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6903) );
  INV_X1 U5759 ( .A(n5648), .ZN(n8830) );
  INV_X1 U5760 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6836) );
  INV_X1 U5761 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6806) );
  INV_X1 U5762 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6511) );
  INV_X1 U5763 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6405) );
  INV_X1 U5764 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U5765 ( .A1(n4627), .A2(n4856), .ZN(n5118) );
  AND2_X1 U5766 ( .A1(n6219), .A2(n6218), .ZN(n6239) );
  AND2_X1 U5767 ( .A1(n4555), .A2(n5872), .ZN(n9689) );
  INV_X1 U5768 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8150) );
  AND2_X1 U5769 ( .A1(n5651), .A2(n8595), .ZN(n5684) );
  NAND2_X1 U5770 ( .A1(n6036), .A2(n6035), .ZN(n8462) );
  AND2_X1 U5771 ( .A1(n4713), .A2(n4327), .ZN(n4300) );
  INV_X1 U5772 ( .A(n7986), .ZN(n7989) );
  OR2_X1 U5773 ( .A1(n6031), .A2(n4329), .ZN(n4301) );
  NAND2_X4 U5774 ( .A1(n5725), .A2(n7182), .ZN(n5763) );
  NAND2_X1 U5775 ( .A1(n5980), .A2(n5979), .ZN(n8355) );
  AND2_X1 U5776 ( .A1(n4708), .A2(n4709), .ZN(n4302) );
  NAND2_X1 U5777 ( .A1(n8166), .A2(n4573), .ZN(n4572) );
  AND2_X1 U5778 ( .A1(n8764), .A2(n8675), .ZN(n4303) );
  OR2_X1 U5779 ( .A1(n8325), .A2(n4586), .ZN(n4304) );
  AND2_X1 U5780 ( .A1(n8685), .A2(n4831), .ZN(n4305) );
  NOR2_X1 U5781 ( .A1(n6072), .A2(n7682), .ZN(n4306) );
  NAND2_X1 U5782 ( .A1(n5550), .A2(n5549), .ZN(n9267) );
  NAND2_X1 U5783 ( .A1(n7867), .A2(n4425), .ZN(n4307) );
  INV_X1 U5784 ( .A(n4716), .ZN(n4711) );
  NAND2_X1 U5785 ( .A1(n4718), .A2(n4717), .ZN(n4716) );
  AND2_X1 U5786 ( .A1(n7920), .A2(n7927), .ZN(n7919) );
  INV_X1 U5787 ( .A(n7919), .ZN(n4402) );
  INV_X1 U5788 ( .A(n8669), .ZN(n4832) );
  AND2_X1 U5789 ( .A1(n7988), .A2(n7984), .ZN(n7981) );
  INV_X1 U5790 ( .A(n7981), .ZN(n4394) );
  NAND2_X1 U5791 ( .A1(n8440), .A2(n8297), .ZN(n4308) );
  NAND2_X1 U5792 ( .A1(n5962), .A2(n5961), .ZN(n9449) );
  INV_X1 U5793 ( .A(n9449), .ZN(n4726) );
  NAND2_X1 U5794 ( .A1(n4551), .A2(n4339), .ZN(n4555) );
  XNOR2_X1 U5795 ( .A(n4561), .B(n4560), .ZN(n6858) );
  INV_X1 U5796 ( .A(n5751), .ZN(n5811) );
  OR2_X1 U5797 ( .A1(n7698), .A2(n6000), .ZN(n4309) );
  INV_X2 U5798 ( .A(n5208), .ZN(n5461) );
  AND2_X1 U5799 ( .A1(n4538), .A2(n4542), .ZN(n4310) );
  NAND2_X1 U5800 ( .A1(n5941), .A2(n5940), .ZN(n7430) );
  INV_X1 U5801 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4734) );
  NAND2_X1 U5802 ( .A1(n6183), .A2(n5699), .ZN(n5704) );
  AND2_X2 U5803 ( .A1(n8545), .A2(n5404), .ZN(n8546) );
  AND2_X1 U5804 ( .A1(n8193), .A2(n8194), .ZN(n4311) );
  NAND2_X1 U5805 ( .A1(n9329), .A2(n8878), .ZN(n4312) );
  NOR2_X1 U5806 ( .A1(n9312), .A2(n9182), .ZN(n4313) );
  AND2_X1 U5807 ( .A1(n7953), .A2(n7940), .ZN(n8264) );
  INV_X1 U5808 ( .A(n9473), .ZN(n8955) );
  AOI21_X1 U5809 ( .B1(n6404), .B2(n5229), .A(n4510), .ZN(n9473) );
  INV_X1 U5810 ( .A(n7839), .ZN(n4576) );
  AND2_X1 U5811 ( .A1(n4736), .A2(n4735), .ZN(n5727) );
  OAI21_X1 U5812 ( .B1(n9098), .B2(n4677), .A(n4673), .ZN(n9071) );
  NOR2_X1 U5813 ( .A1(n7943), .A2(n7989), .ZN(n4314) );
  NAND2_X1 U5814 ( .A1(n4981), .A2(n4980), .ZN(n9282) );
  INV_X1 U5815 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4733) );
  XNOR2_X1 U5816 ( .A(n8407), .B(n8007), .ZN(n8182) );
  NAND2_X1 U5817 ( .A1(n6085), .A2(n6084), .ZN(n8434) );
  AND2_X1 U5818 ( .A1(n5849), .A2(n5848), .ZN(n9762) );
  NOR2_X1 U5819 ( .A1(n8546), .A2(n4838), .ZN(n4315) );
  INV_X1 U5820 ( .A(n8584), .ZN(n4796) );
  AND4_X1 U5821 ( .A1(n5745), .A2(n5744), .A3(n5743), .A4(n5742), .ZN(n7185)
         );
  NOR2_X1 U5822 ( .A1(n8683), .A2(n4832), .ZN(n4831) );
  AND2_X1 U5823 ( .A1(n9001), .A2(n8779), .ZN(n9046) );
  INV_X1 U5824 ( .A(n9046), .ZN(n4700) );
  NAND2_X1 U5825 ( .A1(n5527), .A2(n5526), .ZN(n9272) );
  INV_X1 U5826 ( .A(n9110), .ZN(n4824) );
  AND2_X1 U5827 ( .A1(n9278), .A2(n9113), .ZN(n4316) );
  NAND2_X1 U5828 ( .A1(n6018), .A2(n6017), .ZN(n8455) );
  AND2_X1 U5829 ( .A1(n5921), .A2(n5920), .ZN(n4317) );
  NAND2_X1 U5830 ( .A1(n8209), .A2(n4311), .ZN(n8192) );
  NAND2_X1 U5831 ( .A1(n6123), .A2(n6122), .ZN(n8419) );
  AND2_X1 U5832 ( .A1(n6582), .A2(n6578), .ZN(n4318) );
  NOR2_X1 U5833 ( .A1(n5013), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n4319) );
  NOR2_X1 U5834 ( .A1(n4314), .A2(n4420), .ZN(n4320) );
  INV_X1 U5835 ( .A(n4678), .ZN(n4677) );
  NOR2_X1 U5836 ( .A1(n8967), .A2(n4316), .ZN(n4678) );
  AND2_X1 U5837 ( .A1(n8643), .A2(n8741), .ZN(n4321) );
  NAND2_X1 U5838 ( .A1(n8279), .A2(n4443), .ZN(n4446) );
  AND2_X1 U5839 ( .A1(n5250), .A2(n6946), .ZN(n4322) );
  AND2_X1 U5840 ( .A1(n4819), .A2(n4817), .ZN(n4323) );
  INV_X1 U5841 ( .A(n9256), .ZN(n8942) );
  NAND2_X1 U5842 ( .A1(n5604), .A2(n5603), .ZN(n9256) );
  AND2_X1 U5843 ( .A1(n7595), .A2(n8297), .ZN(n4324) );
  INV_X1 U5844 ( .A(n4724), .ZN(n4723) );
  NOR2_X1 U5845 ( .A1(n9195), .A2(n9211), .ZN(n4724) );
  AND2_X1 U5846 ( .A1(n8703), .A2(n8704), .ZN(n4325) );
  AND2_X1 U5847 ( .A1(n8164), .A2(n8006), .ZN(n4326) );
  INV_X1 U5848 ( .A(n7979), .ZN(n4395) );
  AND2_X1 U5849 ( .A1(n7805), .A2(n7804), .ZN(n7979) );
  NAND2_X1 U5850 ( .A1(n9297), .A2(n9167), .ZN(n4327) );
  NOR2_X1 U5851 ( .A1(n5427), .A2(n5426), .ZN(n4328) );
  INV_X1 U5852 ( .A(n4829), .ZN(n4828) );
  OAI21_X1 U5853 ( .B1(n8783), .B2(n4830), .A(n8784), .ZN(n4829) );
  INV_X1 U5854 ( .A(n4477), .ZN(n4476) );
  NAND2_X1 U5855 ( .A1(n4478), .A2(n9076), .ZN(n4477) );
  INV_X1 U5856 ( .A(n8956), .ZN(n4693) );
  NOR2_X1 U5857 ( .A1(n9473), .A2(n8954), .ZN(n8956) );
  INV_X1 U5858 ( .A(n7871), .ZN(n4752) );
  INV_X1 U5859 ( .A(n4554), .ZN(n4553) );
  OR2_X1 U5860 ( .A1(n4556), .A2(n4343), .ZN(n4554) );
  INV_X1 U5861 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U5862 ( .A1(n4557), .A2(n5716), .ZN(n4329) );
  NOR2_X1 U5863 ( .A1(n8407), .A2(n8169), .ZN(n4330) );
  AND2_X1 U5864 ( .A1(n8387), .A2(n9439), .ZN(n4331) );
  AND2_X1 U5865 ( .A1(n9473), .A2(n8954), .ZN(n4332) );
  AND2_X1 U5866 ( .A1(n9148), .A2(n9136), .ZN(n4333) );
  XOR2_X1 U5867 ( .A(n5048), .B(n5620), .Z(n4334) );
  INV_X1 U5868 ( .A(n4334), .ZN(n4793) );
  AND2_X1 U5869 ( .A1(n4873), .A2(SI_7_), .ZN(n4335) );
  AND2_X1 U5870 ( .A1(n8689), .A2(n7314), .ZN(n4336) );
  INV_X1 U5871 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5645) );
  AND2_X1 U5872 ( .A1(n4858), .A2(SI_3_), .ZN(n4337) );
  OR2_X1 U5873 ( .A1(n4593), .A2(n8264), .ZN(n4338) );
  INV_X1 U5874 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4985) );
  NOR2_X1 U5875 ( .A1(n7065), .A2(n5871), .ZN(n4339) );
  INV_X1 U5876 ( .A(n4674), .ZN(n4673) );
  NAND2_X1 U5877 ( .A1(n4675), .A2(n8970), .ZN(n4674) );
  OR2_X1 U5878 ( .A1(n4927), .A2(n4651), .ZN(n4340) );
  AND2_X1 U5879 ( .A1(n5713), .A2(n4548), .ZN(n4341) );
  INV_X1 U5880 ( .A(n4572), .ZN(n4571) );
  NAND2_X1 U5881 ( .A1(n9172), .A2(n4721), .ZN(n4342) );
  AND2_X1 U5882 ( .A1(n5875), .A2(n5874), .ZN(n4343) );
  AND2_X1 U5883 ( .A1(n8496), .A2(n8497), .ZN(n4344) );
  AND2_X1 U5884 ( .A1(n4569), .A2(n7839), .ZN(n4345) );
  OR2_X1 U5885 ( .A1(n8499), .A2(n4386), .ZN(n4346) );
  AND2_X1 U5886 ( .A1(n4636), .A2(n5330), .ZN(n4347) );
  NOR2_X1 U5887 ( .A1(n9027), .A2(n4698), .ZN(n4697) );
  AND2_X1 U5888 ( .A1(n4395), .A2(n7978), .ZN(n4348) );
  AND2_X1 U5889 ( .A1(n7922), .A2(n7921), .ZN(n8341) );
  INV_X1 U5890 ( .A(n8341), .ZN(n4409) );
  AND2_X1 U5891 ( .A1(n4341), .A2(n4426), .ZN(n4349) );
  OR2_X1 U5892 ( .A1(n4798), .A2(n4797), .ZN(n4350) );
  INV_X1 U5893 ( .A(n7339), .ZN(n4582) );
  AND2_X1 U5894 ( .A1(n4743), .A2(n4308), .ZN(n4351) );
  AND2_X1 U5895 ( .A1(n7343), .A2(n7342), .ZN(n4352) );
  AND2_X1 U5896 ( .A1(n4571), .A2(n4576), .ZN(n4353) );
  AND2_X1 U5897 ( .A1(n9092), .A2(n8997), .ZN(n4823) );
  INV_X1 U5898 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4969) );
  NAND2_X1 U5899 ( .A1(n7942), .A2(n4418), .ZN(n4354) );
  NOR2_X1 U5900 ( .A1(n7501), .A2(n7793), .ZN(n4440) );
  INV_X1 U5901 ( .A(n5763), .ZN(n6124) );
  NAND2_X1 U5902 ( .A1(n6948), .A2(n5289), .ZN(n6862) );
  NAND2_X1 U5903 ( .A1(n7568), .A2(n7567), .ZN(n8152) );
  INV_X1 U5904 ( .A(n8152), .ZN(n4436) );
  INV_X1 U5905 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n4512) );
  NAND2_X1 U5906 ( .A1(n6667), .A2(n5214), .ZN(n6887) );
  NAND2_X1 U5907 ( .A1(n4682), .A2(n4681), .ZN(n9221) );
  XOR2_X1 U5908 ( .A(n6081), .B(n6082), .Z(n4355) );
  OR2_X1 U5909 ( .A1(n8964), .A2(n8963), .ZN(n4356) );
  AND4_X1 U5910 ( .A1(n5970), .A2(n5969), .A3(n5968), .A4(n5967), .ZN(n7788)
         );
  AND4_X1 U5911 ( .A1(n5344), .A2(n5343), .A3(n5342), .A4(n5341), .ZN(n8954)
         );
  INV_X1 U5912 ( .A(n8954), .ZN(n4509) );
  NAND2_X1 U5913 ( .A1(n5040), .A2(n5039), .ZN(n9308) );
  INV_X1 U5914 ( .A(n8689), .ZN(n9329) );
  AND2_X1 U5915 ( .A1(n5319), .A2(n5318), .ZN(n8689) );
  AND2_X1 U5916 ( .A1(n5537), .A2(n5536), .ZN(n8971) );
  OR2_X1 U5917 ( .A1(n9123), .A2(n9135), .ZN(n4357) );
  NOR3_X1 U5918 ( .A1(n9212), .A2(n9297), .A3(n4473), .ZN(n4470) );
  NAND2_X1 U5919 ( .A1(n9118), .A2(n4476), .ZN(n4479) );
  INV_X1 U5920 ( .A(n4437), .ZN(n8332) );
  NAND2_X1 U5921 ( .A1(n4440), .A2(n4438), .ZN(n4437) );
  AND2_X1 U5922 ( .A1(n9256), .A2(n9009), .ZN(n4358) );
  INV_X1 U5923 ( .A(n4471), .ZN(n9158) );
  NOR2_X1 U5924 ( .A1(n9212), .A2(n4473), .ZN(n4471) );
  INV_X1 U5925 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5711) );
  AND2_X1 U5926 ( .A1(n4440), .A2(n8465), .ZN(n4359) );
  AND2_X1 U5927 ( .A1(n4926), .A2(SI_17_), .ZN(n4360) );
  AND2_X1 U5928 ( .A1(n5447), .A2(n4941), .ZN(n4361) );
  OR2_X1 U5929 ( .A1(n7721), .A2(n7724), .ZN(n4362) );
  INV_X1 U5930 ( .A(n8967), .ZN(n4680) );
  AND2_X1 U5931 ( .A1(n4805), .A2(n8988), .ZN(n4363) );
  OR2_X1 U5932 ( .A1(n5908), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n4364) );
  OR2_X1 U5933 ( .A1(n7990), .A2(n8395), .ZN(n7986) );
  INV_X1 U5934 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n4520) );
  INV_X1 U5935 ( .A(n7268), .ZN(n4427) );
  XNOR2_X1 U5936 ( .A(n6180), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U5937 ( .A1(n4428), .A2(n7456), .ZN(n4365) );
  NAND2_X1 U5938 ( .A1(n5654), .A2(n4797), .ZN(n8741) );
  AND2_X1 U5939 ( .A1(n6656), .A2(n4467), .ZN(n4366) );
  NAND2_X1 U5940 ( .A1(n4776), .A2(n4781), .ZN(n6982) );
  INV_X1 U5941 ( .A(n9608), .ZN(n7143) );
  AND2_X1 U5942 ( .A1(n5337), .A2(n5352), .ZN(n9608) );
  INV_X1 U5943 ( .A(n6983), .ZN(n4779) );
  NAND2_X1 U5944 ( .A1(n4669), .A2(n6540), .ZN(n6579) );
  INV_X1 U5945 ( .A(n4660), .ZN(n4659) );
  NOR2_X1 U5946 ( .A1(n5542), .A2(n4661), .ZN(n4660) );
  AND2_X1 U5947 ( .A1(n6862), .A2(n5310), .ZN(n4367) );
  NAND2_X1 U5948 ( .A1(n6396), .A2(n6397), .ZN(n4368) );
  OR2_X1 U5949 ( .A1(n8073), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4369) );
  AND2_X1 U5950 ( .A1(n4455), .A2(n4456), .ZN(n4370) );
  OR2_X1 U5951 ( .A1(n4982), .A2(n4971), .ZN(n4371) );
  AND2_X1 U5952 ( .A1(n9769), .A2(n7456), .ZN(n4372) );
  AND2_X1 U5953 ( .A1(n7546), .A2(SI_29_), .ZN(n4373) );
  AND2_X1 U5954 ( .A1(n4774), .A2(n6627), .ZN(n4374) );
  NAND2_X1 U5955 ( .A1(n5703), .A2(n5702), .ZN(n6229) );
  OR2_X1 U5956 ( .A1(n8138), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4375) );
  NAND2_X1 U5957 ( .A1(n5106), .A2(n5105), .ZN(n6364) );
  INV_X1 U5958 ( .A(n6364), .ZN(n4768) );
  AND2_X1 U5959 ( .A1(n8396), .A2(n9456), .ZN(n9795) );
  AND2_X1 U5960 ( .A1(n4767), .A2(n6365), .ZN(n4376) );
  AND2_X1 U5961 ( .A1(n8930), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4377) );
  OR2_X1 U5962 ( .A1(n6490), .A2(n6560), .ZN(n6547) );
  INV_X1 U5963 ( .A(n6547), .ZN(n4463) );
  INV_X1 U5964 ( .A(n6858), .ZN(n8394) );
  AND2_X1 U5965 ( .A1(n8122), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4378) );
  OR2_X1 U5966 ( .A1(n7989), .A2(n8394), .ZN(n4379) );
  INV_X1 U5967 ( .A(n6721), .ZN(n4521) );
  INV_X1 U5968 ( .A(n8219), .ZN(n8395) );
  AND2_X1 U5969 ( .A1(n5724), .A2(n5723), .ZN(n8219) );
  XNOR2_X1 U5970 ( .A(n5718), .B(n5717), .ZN(n7799) );
  INV_X1 U5971 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4667) );
  NOR2_X4 U5972 ( .A1(n6336), .A2(n4798), .ZN(n9409) );
  NAND2_X1 U5973 ( .A1(n4380), .A2(n8738), .ZN(n4484) );
  NAND2_X1 U5974 ( .A1(n8718), .A2(n8719), .ZN(n4380) );
  NAND2_X1 U5975 ( .A1(n6485), .A2(n6484), .ZN(n4812) );
  NOR2_X1 U5976 ( .A1(n4508), .A2(n4507), .ZN(n4506) );
  AOI21_X1 U5977 ( .B1(n8695), .B2(n4500), .A(n4499), .ZN(n4498) );
  NAND2_X1 U5978 ( .A1(n8702), .A2(n4498), .ZN(n4497) );
  NAND3_X1 U5979 ( .A1(n5490), .A2(n8574), .A3(n5489), .ZN(n8505) );
  NAND2_X1 U5980 ( .A1(n8575), .A2(n8577), .ZN(n5490) );
  OAI21_X1 U5981 ( .B1(n4781), .B2(n4779), .A(n4778), .ZN(n4777) );
  NAND2_X2 U5982 ( .A1(n8210), .A2(n8211), .ZN(n8209) );
  NAND2_X1 U5983 ( .A1(n4616), .A2(n4619), .ZN(n5227) );
  AOI21_X1 U5984 ( .B1(n7996), .B2(n7995), .A(n7994), .ZN(n8003) );
  OAI21_X1 U5985 ( .B1(n7167), .B2(n7170), .A(n7168), .ZN(n5366) );
  NAND2_X2 U5986 ( .A1(n5269), .A2(n5268), .ZN(n6948) );
  NAND2_X1 U5987 ( .A1(n5685), .A2(n4346), .ZN(P1_U3218) );
  OAI21_X1 U5988 ( .B1(n8605), .B2(n8608), .A(n8606), .ZN(n8538) );
  AND2_X2 U5989 ( .A1(n4987), .A2(n5027), .ZN(n5648) );
  BUF_X4 U5990 ( .A(n5102), .Z(n5622) );
  INV_X1 U5991 ( .A(n7572), .ZN(n5111) );
  NAND2_X1 U5992 ( .A1(n8593), .A2(n5567), .ZN(n8594) );
  NAND2_X1 U5993 ( .A1(n6571), .A2(n6627), .ZN(n5188) );
  NAND2_X1 U5994 ( .A1(n5084), .A2(n5083), .ZN(n7572) );
  INV_X1 U5995 ( .A(n4799), .ZN(n5029) );
  AND2_X2 U5996 ( .A1(n4968), .A2(n4967), .ZN(n4799) );
  NAND2_X1 U5997 ( .A1(n8530), .A2(n8531), .ZN(n8593) );
  NAND2_X1 U5998 ( .A1(n5188), .A2(n6628), .ZN(n6630) );
  NAND3_X1 U5999 ( .A1(n4763), .A2(n4764), .A3(n8556), .ZN(n8555) );
  AOI21_X2 U6000 ( .B1(n6948), .B2(n4780), .A(n4777), .ZN(n5346) );
  NAND3_X1 U6001 ( .A1(n5060), .A2(n6324), .A3(n5061), .ZN(n6325) );
  OR2_X1 U6002 ( .A1(n7987), .A2(n4379), .ZN(n4388) );
  NAND2_X1 U6003 ( .A1(n4388), .A2(n4387), .ZN(n4843) );
  NAND2_X1 U6004 ( .A1(n4400), .A2(n4398), .ZN(n7924) );
  NAND2_X1 U6005 ( .A1(n4401), .A2(n4404), .ZN(n4399) );
  NAND2_X1 U6006 ( .A1(n7915), .A2(n4401), .ZN(n4400) );
  AOI21_X1 U6007 ( .B1(n7914), .B2(n7343), .A(n4406), .ZN(n4405) );
  NOR2_X1 U6008 ( .A1(n4409), .A2(n4408), .ZN(n4407) );
  NOR2_X1 U6009 ( .A1(n7920), .A2(n7989), .ZN(n4408) );
  NAND2_X1 U6010 ( .A1(n7956), .A2(n4417), .ZN(n4411) );
  NAND3_X1 U6011 ( .A1(n4411), .A2(n4412), .A3(n4410), .ZN(n7965) );
  NAND3_X1 U6012 ( .A1(n4354), .A2(n4417), .A3(n4414), .ZN(n4413) );
  NAND2_X1 U6013 ( .A1(n4422), .A2(n4421), .ZN(n4424) );
  NAND3_X1 U6014 ( .A1(n7862), .A2(n7861), .A3(n7873), .ZN(n4422) );
  AND3_X1 U6015 ( .A1(n4753), .A2(n5698), .A3(n5687), .ZN(n6183) );
  AOI211_X1 U6016 ( .C1(n7805), .C2(n8159), .A(n4432), .B(n4433), .ZN(n4431)
         );
  NAND2_X1 U6017 ( .A1(n4439), .A2(n4440), .ZN(n8307) );
  INV_X1 U6018 ( .A(n4440), .ZN(n8352) );
  NAND2_X1 U6019 ( .A1(n8279), .A2(n4441), .ZN(n8215) );
  INV_X1 U6020 ( .A(n4446), .ZN(n8226) );
  NAND2_X1 U6021 ( .A1(n4455), .A2(n4453), .ZN(n6607) );
  AND2_X1 U6022 ( .A1(n6427), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4460) );
  NAND2_X1 U6023 ( .A1(n4799), .A2(n4465), .ZN(n4973) );
  INV_X1 U6024 ( .A(n4470), .ZN(n9144) );
  INV_X1 U6025 ( .A(n4479), .ZN(n9072) );
  NAND2_X1 U6026 ( .A1(n9031), .A2(n4480), .ZN(n4482) );
  NAND2_X1 U6027 ( .A1(n9031), .A2(n8942), .ZN(n9033) );
  INV_X1 U6028 ( .A(n4482), .ZN(n9012) );
  AOI21_X1 U6029 ( .B1(n9033), .B2(n9252), .A(n9242), .ZN(n4483) );
  NAND2_X1 U6030 ( .A1(n4484), .A2(n9092), .ZN(n4486) );
  AOI21_X1 U6031 ( .B1(n8727), .B2(n8741), .A(n4486), .ZN(n4485) );
  AOI21_X1 U6032 ( .B1(n8733), .B2(n8732), .A(n8731), .ZN(n8734) );
  OR2_X1 U6033 ( .A1(n4892), .A2(n4491), .ZN(n4487) );
  NAND2_X1 U6034 ( .A1(n4487), .A2(n4488), .ZN(n5331) );
  NAND2_X1 U6035 ( .A1(n7648), .A2(n4529), .ZN(n4527) );
  OAI21_X1 U6036 ( .B1(n7648), .B2(n4531), .A(n4529), .ZN(n7482) );
  AOI21_X1 U6037 ( .B1(n4531), .B2(n4529), .A(n4526), .ZN(n4525) );
  NAND2_X2 U6038 ( .A1(n7517), .A2(n7516), .ZN(n7515) );
  NAND2_X1 U6039 ( .A1(n7692), .A2(n4539), .ZN(n4537) );
  NAND2_X1 U6040 ( .A1(n7692), .A2(n4543), .ZN(n4538) );
  NAND2_X1 U6041 ( .A1(n7692), .A2(n7691), .ZN(n7776) );
  NAND2_X1 U6042 ( .A1(n7155), .A2(n4547), .ZN(n6938) );
  INV_X1 U6043 ( .A(n5872), .ZN(n4556) );
  AND2_X1 U6044 ( .A1(n8399), .A2(n8400), .ZN(n4574) );
  NAND2_X1 U6045 ( .A1(n8176), .A2(n4345), .ZN(n4563) );
  NAND3_X1 U6046 ( .A1(n4565), .A2(n4564), .A3(n4563), .ZN(n4575) );
  NAND2_X1 U6047 ( .A1(n4562), .A2(n4353), .ZN(n4565) );
  INV_X1 U6048 ( .A(n8176), .ZN(n4562) );
  OAI21_X1 U6049 ( .B1(n8176), .B2(n8182), .A(n4577), .ZN(n8158) );
  NAND3_X1 U6050 ( .A1(n4565), .A2(n4566), .A3(n4563), .ZN(n8401) );
  NAND2_X1 U6051 ( .A1(n4575), .A2(n4574), .ZN(n8477) );
  NAND2_X1 U6052 ( .A1(n5687), .A2(n4578), .ZN(n5861) );
  INV_X1 U6053 ( .A(n7270), .ZN(n4583) );
  NAND2_X1 U6054 ( .A1(n4579), .A2(n4580), .ZN(n7475) );
  NAND2_X1 U6055 ( .A1(n7270), .A2(n7339), .ZN(n4579) );
  OAI21_X1 U6056 ( .B1(n8345), .B2(n4304), .A(n4584), .ZN(n7589) );
  INV_X1 U6057 ( .A(n7589), .ZN(n7591) );
  INV_X1 U6058 ( .A(n4588), .ZN(n8251) );
  NAND2_X1 U6059 ( .A1(n8429), .A2(n4604), .ZN(n4603) );
  INV_X1 U6060 ( .A(n4609), .ZN(n8224) );
  OAI22_X1 U6061 ( .A1(n5793), .A2(n6264), .B1(n6700), .B2(n6741), .ZN(n4611)
         );
  NAND2_X1 U6063 ( .A1(n7366), .A2(n4352), .ZN(n7432) );
  INV_X1 U6064 ( .A(n7185), .ZN(n7184) );
  NAND2_X2 U6065 ( .A1(n9433), .A2(n5973), .ZN(n7698) );
  NAND2_X1 U6066 ( .A1(n5789), .A2(n7078), .ZN(n7156) );
  NAND2_X1 U6067 ( .A1(n7197), .A2(n7196), .ZN(n7463) );
  NAND2_X1 U6068 ( .A1(n7433), .A2(n7913), .ZN(n7498) );
  NOR2_X2 U6069 ( .A1(n5697), .A2(n5696), .ZN(n5698) );
  NAND2_X1 U6070 ( .A1(n7674), .A2(n5761), .ZN(n7753) );
  NAND3_X1 U6071 ( .A1(n7981), .A2(n4615), .A3(n4348), .ZN(n4614) );
  NAND2_X1 U6072 ( .A1(n5167), .A2(n4617), .ZN(n4616) );
  NAND2_X1 U6073 ( .A1(n4623), .A2(n7558), .ZN(n7805) );
  NAND3_X1 U6074 ( .A1(n5094), .A2(n5095), .A3(n5119), .ZN(n4625) );
  NAND2_X1 U6075 ( .A1(n5094), .A2(n5095), .ZN(n4627) );
  INV_X1 U6076 ( .A(n4856), .ZN(n4626) );
  NAND2_X1 U6077 ( .A1(n4634), .A2(n4361), .ZN(n4945) );
  NAND2_X1 U6078 ( .A1(n4635), .A2(n4347), .ZN(n4912) );
  NAND2_X1 U6079 ( .A1(n5351), .A2(n4645), .ZN(n4643) );
  OAI21_X1 U6080 ( .B1(n5518), .B2(n5517), .A(n5521), .ZN(n5543) );
  OAI21_X1 U6081 ( .B1(n5518), .B2(n4656), .A(n4654), .ZN(n5571) );
  NAND2_X1 U6082 ( .A1(n4662), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4668) );
  INV_X1 U6083 ( .A(n4668), .ZN(n4665) );
  NAND2_X1 U6084 ( .A1(n4846), .A2(n4667), .ZN(n4666) );
  INV_X1 U6085 ( .A(n6541), .ZN(n4669) );
  NAND2_X1 U6086 ( .A1(n7313), .A2(n4687), .ZN(n4682) );
  NAND2_X1 U6087 ( .A1(n4695), .A2(n4696), .ZN(n8980) );
  NAND2_X1 U6088 ( .A1(n9040), .A2(n4697), .ZN(n4695) );
  NAND2_X1 U6089 ( .A1(n6844), .A2(n4702), .ZN(n4701) );
  NAND2_X1 U6090 ( .A1(n4701), .A2(n4703), .ZN(n9397) );
  NAND2_X1 U6091 ( .A1(n8960), .A2(n4300), .ZN(n4708) );
  INV_X1 U6092 ( .A(n7199), .ZN(n7812) );
  NAND2_X1 U6093 ( .A1(n7199), .A2(n4845), .ZN(n8376) );
  AND2_X1 U6094 ( .A1(n7855), .A2(n7857), .ZN(n4845) );
  AND2_X1 U6095 ( .A1(n7854), .A2(n8374), .ZN(n7199) );
  NAND2_X2 U6096 ( .A1(n7361), .A2(n7890), .ZN(n7466) );
  NAND4_X1 U6097 ( .A1(n4728), .A2(n4727), .A3(n5686), .A4(n4735), .ZN(n5825)
         );
  NAND3_X1 U6098 ( .A1(n4736), .A2(n4734), .A3(n4731), .ZN(n4730) );
  NAND2_X1 U6099 ( .A1(n5727), .A2(n4732), .ZN(n5790) );
  OAI21_X2 U6100 ( .B1(n8209), .B2(n4739), .A(n4737), .ZN(n8165) );
  OAI21_X2 U6101 ( .B1(n7205), .B2(n4750), .A(n4746), .ZN(n7274) );
  NAND2_X1 U6102 ( .A1(n4749), .A2(n4748), .ZN(n4747) );
  NAND2_X1 U6103 ( .A1(n4748), .A2(n7871), .ZN(n4750) );
  INV_X1 U6104 ( .A(n7817), .ZN(n4748) );
  INV_X1 U6105 ( .A(n4750), .ZN(n4751) );
  NAND2_X1 U6106 ( .A1(n7225), .A2(n4751), .ZN(n7228) );
  NAND2_X1 U6107 ( .A1(n7205), .A2(n7206), .ZN(n7225) );
  NAND3_X1 U6108 ( .A1(n5687), .A2(n5698), .A3(n4755), .ZN(n6186) );
  NAND2_X1 U6109 ( .A1(n8240), .A2(n4760), .ZN(n4757) );
  NAND2_X1 U6110 ( .A1(n4757), .A2(n4758), .ZN(n8210) );
  INV_X1 U6111 ( .A(n4761), .ZN(n8239) );
  NAND2_X1 U6112 ( .A1(n6887), .A2(n5251), .ZN(n4762) );
  NAND2_X1 U6113 ( .A1(n6668), .A2(n6669), .ZN(n6667) );
  NAND2_X1 U6114 ( .A1(n8505), .A2(n8508), .ZN(n4763) );
  OAI211_X1 U6115 ( .C1(n6364), .C2(n4766), .A(n4765), .B(n4769), .ZN(n6416)
         );
  NAND3_X1 U6116 ( .A1(n5111), .A2(n5110), .A3(n5127), .ZN(n4765) );
  NAND2_X1 U6117 ( .A1(n5111), .A2(n5110), .ZN(n6363) );
  NAND2_X1 U6118 ( .A1(n6363), .A2(n6364), .ZN(n4767) );
  INV_X1 U6119 ( .A(n5126), .ZN(n4771) );
  OAI21_X1 U6120 ( .B1(n6324), .B2(n4772), .A(n6325), .ZN(n9519) );
  NAND3_X1 U6121 ( .A1(n4774), .A2(n6572), .A3(n6627), .ZN(n6571) );
  OR2_X2 U6122 ( .A1(n5164), .A2(n5163), .ZN(n4774) );
  NAND2_X1 U6123 ( .A1(n4983), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4986) );
  NAND2_X1 U6124 ( .A1(n4986), .A2(n4985), .ZN(n5027) );
  INV_X1 U6125 ( .A(n6336), .ZN(n5028) );
  AND2_X2 U6126 ( .A1(n4299), .A2(n6357), .ZN(n5102) );
  INV_X1 U6127 ( .A(n6837), .ZN(n4798) );
  OAI21_X1 U6128 ( .B1(n5011), .B2(n5013), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5012) );
  NAND2_X1 U6129 ( .A1(n4805), .A2(n4804), .ZN(n9180) );
  OAI21_X1 U6130 ( .B1(n6484), .B2(n4810), .A(n8751), .ZN(n4809) );
  NAND2_X1 U6131 ( .A1(n4812), .A2(n4811), .ZN(n8653) );
  NAND2_X1 U6132 ( .A1(n4812), .A2(n8754), .ZN(n8654) );
  OAI21_X1 U6133 ( .B1(n9164), .B2(n4816), .A(n4813), .ZN(n9124) );
  NAND2_X1 U6134 ( .A1(n9109), .A2(n4823), .ZN(n4820) );
  NAND2_X1 U6135 ( .A1(n4826), .A2(n4827), .ZN(n7303) );
  NAND2_X1 U6136 ( .A1(n5494), .A2(n5493), .ZN(n5518) );
  OAI21_X1 U6137 ( .B1(n8872), .B2(n8871), .A(n8870), .ZN(n8877) );
  INV_X1 U6138 ( .A(n8304), .ZN(n7594) );
  OR2_X1 U6139 ( .A1(n8744), .A2(n6837), .ZN(n8872) );
  NAND2_X1 U6140 ( .A1(n5974), .A2(n5714), .ZN(n6031) );
  OAI222_X1 U6141 ( .A1(n8377), .A2(n7610), .B1(n8006), .B2(n8372), .C1(n8004), 
        .C2(n7609), .ZN(n7611) );
  INV_X1 U6142 ( .A(n8545), .ZN(n8548) );
  XNOR2_X1 U6143 ( .A(n7561), .B(n7560), .ZN(n8634) );
  INV_X1 U6144 ( .A(n7014), .ZN(n6999) );
  NAND2_X1 U6145 ( .A1(n7203), .A2(n4844), .ZN(n7204) );
  OR2_X2 U6146 ( .A1(n7911), .A2(n7441), .ZN(n7445) );
  NOR2_X1 U6147 ( .A1(n7368), .A2(n7491), .ZN(n7369) );
  AOI21_X1 U6148 ( .B1(n8499), .B2(n5684), .A(n5683), .ZN(n5685) );
  AND2_X1 U6149 ( .A1(n7641), .A2(n7640), .ZN(n7720) );
  NAND2_X1 U6150 ( .A1(n7185), .A2(n7673), .ZN(n7841) );
  INV_X1 U6151 ( .A(n7673), .ZN(n7186) );
  XNOR2_X1 U6152 ( .A(n5763), .B(n7673), .ZN(n5758) );
  INV_X1 U6153 ( .A(n5046), .ZN(n5654) );
  AND2_X1 U6154 ( .A1(n5046), .A2(n5648), .ZN(n6445) );
  NAND2_X2 U6155 ( .A1(n5924), .A2(n5923), .ZN(n7491) );
  INV_X1 U6156 ( .A(n7328), .ZN(n7330) );
  AND2_X1 U6157 ( .A1(n5797), .A2(n5796), .ZN(n4835) );
  INV_X1 U6158 ( .A(n9031), .ZN(n9041) );
  AND2_X1 U6159 ( .A1(n4908), .A2(n4907), .ZN(n4836) );
  AND2_X1 U6160 ( .A1(n5408), .A2(n5407), .ZN(n4838) );
  AND2_X1 U6161 ( .A1(n4891), .A2(n4890), .ZN(n4839) );
  INV_X1 U6162 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5738) );
  OAI21_X1 U6163 ( .B1(n7993), .B2(n4843), .A(n7992), .ZN(n7994) );
  AND2_X1 U6164 ( .A1(n4884), .A2(n4883), .ZN(n4840) );
  NAND2_X1 U6165 ( .A1(n7188), .A2(n7187), .ZN(n7292) );
  AND3_X1 U6166 ( .A1(n6080), .A2(n6079), .A3(n6078), .ZN(n8297) );
  INV_X1 U6167 ( .A(n7745), .ZN(n7599) );
  AND2_X1 U6168 ( .A1(n6095), .A2(n6094), .ZN(n8278) );
  INV_X1 U6169 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5332) );
  NOR2_X1 U6170 ( .A1(n6238), .A2(n6237), .ZN(n4841) );
  INV_X1 U6171 ( .A(n8351), .ZN(n8377) );
  AND2_X1 U6172 ( .A1(n5385), .A2(n5384), .ZN(n4842) );
  NAND2_X1 U6173 ( .A1(n7190), .A2(n7189), .ZN(n7403) );
  NAND2_X2 U6174 ( .A1(n7209), .A2(n8218), .ZN(n8383) );
  NAND2_X1 U6175 ( .A1(n8022), .A2(n9750), .ZN(n4844) );
  INV_X2 U6176 ( .A(n9669), .ZN(n9352) );
  INV_X2 U6177 ( .A(n9671), .ZN(n9334) );
  INV_X1 U6178 ( .A(n5161), .ZN(n5363) );
  INV_X1 U6179 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4970) );
  INV_X1 U6180 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4974) );
  INV_X1 U6181 ( .A(n5989), .ZN(n5981) );
  INV_X1 U6182 ( .A(n7892), .ZN(n7272) );
  INV_X1 U6183 ( .A(n5339), .ZN(n4999) );
  INV_X1 U6184 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n4903) );
  NOR2_X1 U6185 ( .A1(n5900), .A2(n6703), .ZN(n5912) );
  AND2_X1 U6186 ( .A1(n5912), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U6187 ( .A1(n5981), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5991) );
  INV_X1 U6188 ( .A(n8278), .ZN(n7597) );
  AOI21_X1 U6189 ( .B1(n7274), .B2(n7273), .A(n7272), .ZN(n7276) );
  NAND2_X1 U6190 ( .A1(n6180), .A2(n6179), .ZN(n6181) );
  INV_X1 U6191 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5699) );
  OR2_X1 U6192 ( .A1(n6324), .A2(n5588), .ZN(n5065) );
  INV_X1 U6193 ( .A(n5234), .ZN(n4996) );
  INV_X1 U6194 ( .A(n5396), .ZN(n5001) );
  INV_X1 U6195 ( .A(n5530), .ZN(n5528) );
  INV_X1 U6196 ( .A(n5473), .ZN(n5004) );
  INV_X1 U6197 ( .A(n5416), .ZN(n5002) );
  OR2_X1 U6198 ( .A1(n5357), .A2(n7148), .ZN(n5374) );
  INV_X1 U6199 ( .A(n6543), .ZN(n6540) );
  INV_X1 U6200 ( .A(n5031), .ZN(n4928) );
  INV_X1 U6201 ( .A(SI_8_), .ZN(n10017) );
  INV_X1 U6202 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5831) );
  NAND2_X1 U6203 ( .A1(n6048), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U6204 ( .A1(n6086), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6101) );
  INV_X1 U6205 ( .A(n6940), .ZN(n5824) );
  OR2_X1 U6206 ( .A1(n6021), .A2(n10019), .ZN(n6050) );
  OR2_X1 U6207 ( .A1(n7471), .A2(n9789), .ZN(n7368) );
  OR2_X1 U6208 ( .A1(n7422), .A2(n6190), .ZN(n6191) );
  OR2_X1 U6209 ( .A1(n5093), .A2(n10032), .ZN(n5098) );
  NAND2_X1 U6210 ( .A1(n5528), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U6211 ( .A1(n5004), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U6212 ( .A1(n5003), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5473) );
  INV_X1 U6213 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8549) );
  INV_X1 U6214 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7148) );
  OAI21_X1 U6215 ( .B1(n9022), .B2(n9004), .A(n9003), .ZN(n9006) );
  INV_X1 U6216 ( .A(n8971), .ZN(n8972) );
  NAND2_X1 U6217 ( .A1(n4992), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4993) );
  INV_X1 U6218 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5388) );
  OR2_X1 U6219 ( .A1(n6139), .A2(n9948), .ZN(n6171) );
  OR2_X1 U6220 ( .A1(n6076), .A2(n7686), .ZN(n6088) );
  AND2_X1 U6221 ( .A1(n6119), .A2(n4362), .ZN(n6120) );
  OR2_X1 U6222 ( .A1(n6101), .A2(n7642), .ZN(n6125) );
  INV_X1 U6223 ( .A(n8011), .ZN(n8296) );
  OR2_X1 U6224 ( .A1(n5943), .A2(n5942), .ZN(n5964) );
  INV_X1 U6225 ( .A(n7752), .ZN(n5772) );
  NAND2_X1 U6226 ( .A1(n6007), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U6227 ( .A1(n9674), .A2(n7809), .ZN(n7772) );
  AND2_X1 U6228 ( .A1(n7612), .A2(n6172), .ZN(n8162) );
  INV_X1 U6229 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6703) );
  INV_X1 U6230 ( .A(n9694), .ZN(n9700) );
  NAND2_X1 U6231 ( .A1(n6212), .A2(n5719), .ZN(n6516) );
  INV_X1 U6232 ( .A(n7230), .ZN(n7877) );
  INV_X1 U6233 ( .A(n9750), .ZN(n7458) );
  OR2_X1 U6234 ( .A1(n9801), .A2(n8395), .ZN(n8389) );
  NAND2_X1 U6235 ( .A1(n9709), .A2(n6193), .ZN(n8471) );
  NAND2_X1 U6236 ( .A1(n7181), .A2(n8395), .ZN(n8396) );
  AND2_X1 U6237 ( .A1(n7399), .A2(n6191), .ZN(n9706) );
  INV_X1 U6238 ( .A(n6183), .ZN(n6188) );
  INV_X1 U6239 ( .A(n9126), .ZN(n8966) );
  NOR2_X1 U6240 ( .A1(n5366), .A2(n5365), .ZN(n8605) );
  OR2_X1 U6241 ( .A1(n5236), .A2(n5220), .ZN(n5258) );
  INV_X1 U6242 ( .A(n6323), .ZN(n5676) );
  OR2_X1 U6243 ( .A1(n9073), .A2(n5658), .ZN(n5537) );
  OR2_X1 U6244 ( .A1(n5394), .A2(n8549), .ZN(n5396) );
  NOR2_X1 U6245 ( .A1(n9272), .A2(n8972), .ZN(n8973) );
  INV_X1 U6246 ( .A(n9282), .ZN(n9105) );
  INV_X1 U6247 ( .A(n9106), .ZN(n9135) );
  INV_X1 U6248 ( .A(n9183), .ZN(n8961) );
  INV_X1 U6249 ( .A(n7315), .ZN(n7324) );
  NOR2_X1 U6250 ( .A1(n9663), .A2(n5648), .ZN(n6328) );
  INV_X1 U6251 ( .A(n6435), .ZN(n6453) );
  AND2_X1 U6252 ( .A1(n4923), .A2(n4922), .ZN(n5367) );
  OR2_X1 U6253 ( .A1(n5034), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5253) );
  INV_X4 U6254 ( .A(n5746), .ZN(n7554) );
  NAND2_X1 U6255 ( .A1(n6121), .A2(n6120), .ZN(n7692) );
  INV_X1 U6256 ( .A(n8371), .ZN(n8328) );
  INV_X1 U6257 ( .A(n6516), .ZN(n6699) );
  AND2_X1 U6258 ( .A1(n6169), .A2(n7997), .ZN(n9790) );
  OR2_X1 U6259 ( .A1(n6697), .A2(n9710), .ZN(n7999) );
  AND2_X1 U6260 ( .A1(n6113), .A2(n6112), .ZN(n8242) );
  AND4_X1 U6261 ( .A1(n5948), .A2(n5947), .A3(n5946), .A4(n5945), .ZN(n7487)
         );
  AND2_X1 U6262 ( .A1(n6716), .A2(n7998), .ZN(n9694) );
  AND2_X1 U6263 ( .A1(n6753), .A2(n6752), .ZN(n9695) );
  AND2_X1 U6264 ( .A1(n7948), .A2(n7949), .ZN(n8293) );
  AND2_X1 U6265 ( .A1(n7892), .A2(n7881), .ZN(n7884) );
  INV_X1 U6266 ( .A(n9762), .ZN(n7874) );
  NAND2_X1 U6267 ( .A1(n7833), .A2(n7808), .ZN(n8351) );
  AND2_X1 U6268 ( .A1(n8383), .A2(n7208), .ZN(n8363) );
  NOR2_X1 U6269 ( .A1(n8473), .A2(n8471), .ZN(n8393) );
  INV_X1 U6270 ( .A(n9795), .ZN(n9806) );
  INV_X1 U6271 ( .A(n9706), .ZN(n9707) );
  INV_X1 U6272 ( .A(n5741), .ZN(n8492) );
  INV_X1 U6273 ( .A(n6267), .ZN(n8629) );
  AND2_X1 U6274 ( .A1(n5459), .A2(n5458), .ZN(n8963) );
  AND2_X1 U6275 ( .A1(n6294), .A2(n9522), .ZN(n9616) );
  INV_X1 U6276 ( .A(n9616), .ZN(n9623) );
  INV_X1 U6277 ( .A(n9543), .ZN(n9629) );
  AND2_X1 U6278 ( .A1(n9522), .A2(n6445), .ZN(n9231) );
  NAND2_X1 U6279 ( .A1(n9657), .A2(n6328), .ZN(n9644) );
  AND2_X1 U6280 ( .A1(n9653), .A2(n6358), .ZN(n9237) );
  INV_X1 U6281 ( .A(n9482), .ZN(n9332) );
  AND3_X1 U6282 ( .A1(n6331), .A2(n6330), .A3(n6329), .ZN(n6339) );
  AND2_X1 U6283 ( .A1(n6241), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5647) );
  AND2_X1 U6284 ( .A1(n5644), .A2(n5643), .ZN(n6353) );
  AND2_X1 U6285 ( .A1(n5391), .A2(n5390), .ZN(n8930) );
  AND2_X1 U6286 ( .A1(n5217), .A2(n5253), .ZN(n9600) );
  INV_X1 U6287 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9865) );
  AND2_X1 U6288 ( .A1(n7133), .A2(n6204), .ZN(n6697) );
  NAND2_X1 U6289 ( .A1(n9428), .A2(n8328), .ZN(n7790) );
  INV_X1 U6290 ( .A(n8434), .ZN(n8262) );
  INV_X1 U6291 ( .A(n8455), .ZN(n7771) );
  OR2_X1 U6292 ( .A1(n6012), .A2(n6011), .ZN(n8011) );
  NAND2_X1 U6293 ( .A1(n6229), .A2(n6751), .ZN(n9699) );
  INV_X1 U6294 ( .A(n9695), .ZN(n9698) );
  OR2_X1 U6295 ( .A1(n8362), .A2(n7224), .ZN(n8340) );
  INV_X2 U6296 ( .A(n8383), .ZN(n8362) );
  INV_X1 U6297 ( .A(n9830), .ZN(n9828) );
  AND2_X2 U6298 ( .A1(n8475), .A2(n8393), .ZN(n9830) );
  INV_X1 U6299 ( .A(n9809), .ZN(n9807) );
  NAND2_X1 U6300 ( .A1(n9708), .A2(n9707), .ZN(n9861) );
  INV_X1 U6301 ( .A(n6212), .ZN(n7624) );
  INV_X1 U6302 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9921) );
  INV_X1 U6303 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6279) );
  INV_X1 U6304 ( .A(n9407), .ZN(n9417) );
  INV_X1 U6305 ( .A(n9272), .ZN(n9076) );
  INV_X1 U6306 ( .A(n8612), .ZN(n8588) );
  INV_X1 U6307 ( .A(n7012), .ZN(n7025) );
  AND2_X1 U6308 ( .A1(n5655), .A2(n9644), .ZN(n8604) );
  NAND2_X1 U6309 ( .A1(n5558), .A2(n5557), .ZN(n9080) );
  INV_X1 U6310 ( .A(n8647), .ZN(n9198) );
  OR2_X1 U6311 ( .A1(P1_U3083), .A2(n6286), .ZN(n9621) );
  NAND2_X1 U6312 ( .A1(n9653), .A2(n9639), .ZN(n9239) );
  NAND2_X1 U6313 ( .A1(n6339), .A2(n6353), .ZN(n9671) );
  NAND2_X1 U6314 ( .A1(n6339), .A2(n6332), .ZN(n9669) );
  INV_X1 U6315 ( .A(n9660), .ZN(n9659) );
  NAND2_X1 U6316 ( .A1(n5057), .A2(n5647), .ZN(n6320) );
  INV_X1 U6317 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7426) );
  INV_X1 U6318 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6556) );
  INV_X1 U6319 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6314) );
  INV_X1 U6320 ( .A(n9357), .ZN(n9360) );
  AND2_X1 U6321 ( .A1(n6697), .A2(n9715), .ZN(P2_U3966) );
  AND2_X1 U6322 ( .A1(n6286), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  INV_X2 U6323 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  AND2_X1 U6324 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4847) );
  NAND2_X1 U6325 ( .A1(n4848), .A2(n4847), .ZN(n5749) );
  AND2_X1 U6326 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n4849) );
  NAND2_X1 U6327 ( .A1(n4859), .A2(n4849), .ZN(n5054) );
  NAND2_X1 U6328 ( .A1(n5749), .A2(n5054), .ZN(n4851) );
  INV_X1 U6329 ( .A(SI_1_), .ZN(n4850) );
  XNOR2_X1 U6330 ( .A(n4851), .B(n4850), .ZN(n5068) );
  MUX2_X1 U6331 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4859), .Z(n5067) );
  NAND2_X1 U6332 ( .A1(n5068), .A2(n5067), .ZN(n4853) );
  NAND2_X1 U6333 ( .A1(n4851), .A2(SI_1_), .ZN(n4852) );
  NAND2_X1 U6334 ( .A1(n4853), .A2(n4852), .ZN(n5094) );
  INV_X1 U6335 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6264) );
  INV_X1 U6336 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10032) );
  MUX2_X1 U6337 ( .A(n6264), .B(n10032), .S(n4859), .Z(n4854) );
  XNOR2_X1 U6338 ( .A(n4854), .B(SI_2_), .ZN(n5095) );
  INV_X1 U6339 ( .A(n4854), .ZN(n4855) );
  NAND2_X1 U6340 ( .A1(n4855), .A2(SI_2_), .ZN(n4856) );
  INV_X1 U6341 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6262) );
  INV_X1 U6342 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6245) );
  MUX2_X1 U6343 ( .A(n6262), .B(n6245), .S(n4859), .Z(n4857) );
  INV_X1 U6344 ( .A(n4857), .ZN(n4858) );
  INV_X1 U6345 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6258) );
  INV_X1 U6346 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6249) );
  XNOR2_X1 U6347 ( .A(n4861), .B(SI_4_), .ZN(n5134) );
  NAND2_X1 U6348 ( .A1(n5133), .A2(n5134), .ZN(n4864) );
  INV_X1 U6349 ( .A(n4861), .ZN(n4862) );
  NAND2_X1 U6350 ( .A1(n4862), .A2(SI_4_), .ZN(n4863) );
  NAND2_X1 U6351 ( .A1(n4864), .A2(n4863), .ZN(n5156) );
  INV_X1 U6352 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6260) );
  INV_X1 U6353 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6250) );
  MUX2_X1 U6354 ( .A(n6260), .B(n6250), .S(n7548), .Z(n4865) );
  XNOR2_X1 U6355 ( .A(n4865), .B(SI_5_), .ZN(n5157) );
  NAND2_X1 U6356 ( .A1(n5156), .A2(n5157), .ZN(n4868) );
  INV_X1 U6357 ( .A(n4865), .ZN(n4866) );
  NAND2_X1 U6358 ( .A1(n4866), .A2(SI_5_), .ZN(n4867) );
  MUX2_X1 U6359 ( .A(n6256), .B(n6253), .S(n7548), .Z(n4869) );
  XNOR2_X1 U6360 ( .A(n4869), .B(SI_6_), .ZN(n5168) );
  INV_X1 U6361 ( .A(n4869), .ZN(n4870) );
  NAND2_X1 U6362 ( .A1(n4870), .A2(SI_6_), .ZN(n4871) );
  MUX2_X1 U6363 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7548), .Z(n4873) );
  XNOR2_X1 U6364 ( .A(n4873), .B(SI_7_), .ZN(n5191) );
  INV_X1 U6365 ( .A(n5191), .ZN(n4872) );
  INV_X1 U6366 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n4874) );
  MUX2_X1 U6367 ( .A(n6279), .B(n4874), .S(n7548), .Z(n4875) );
  NAND2_X1 U6368 ( .A1(n4875), .A2(n10017), .ZN(n4878) );
  INV_X1 U6369 ( .A(n4875), .ZN(n4876) );
  NAND2_X1 U6370 ( .A1(n4876), .A2(SI_8_), .ZN(n4877) );
  NAND2_X1 U6371 ( .A1(n4878), .A2(n4877), .ZN(n5228) );
  INV_X1 U6372 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n4879) );
  MUX2_X1 U6373 ( .A(n6283), .B(n4879), .S(n7548), .Z(n4881) );
  INV_X1 U6374 ( .A(SI_9_), .ZN(n4880) );
  NAND2_X1 U6375 ( .A1(n4881), .A2(n4880), .ZN(n4884) );
  INV_X1 U6376 ( .A(n4881), .ZN(n4882) );
  NAND2_X1 U6377 ( .A1(n4882), .A2(SI_9_), .ZN(n4883) );
  NAND2_X1 U6378 ( .A1(n5215), .A2(n4840), .ZN(n4885) );
  NAND2_X1 U6379 ( .A1(n4885), .A2(n4884), .ZN(n5252) );
  INV_X1 U6380 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n4886) );
  MUX2_X1 U6381 ( .A(n6312), .B(n4886), .S(n7548), .Z(n4888) );
  INV_X1 U6382 ( .A(SI_10_), .ZN(n4887) );
  NAND2_X1 U6383 ( .A1(n4888), .A2(n4887), .ZN(n4891) );
  INV_X1 U6384 ( .A(n4888), .ZN(n4889) );
  NAND2_X1 U6385 ( .A1(n4889), .A2(SI_10_), .ZN(n4890) );
  MUX2_X1 U6386 ( .A(n6315), .B(n6314), .S(n7548), .Z(n4893) );
  XNOR2_X1 U6387 ( .A(n4893), .B(SI_11_), .ZN(n5270) );
  INV_X1 U6388 ( .A(n5270), .ZN(n4896) );
  INV_X1 U6389 ( .A(n4893), .ZN(n4894) );
  NAND2_X1 U6390 ( .A1(n4894), .A2(SI_11_), .ZN(n4895) );
  INV_X1 U6391 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n4897) );
  MUX2_X1 U6392 ( .A(n6343), .B(n4897), .S(n7554), .Z(n4899) );
  INV_X1 U6393 ( .A(SI_12_), .ZN(n4898) );
  INV_X1 U6394 ( .A(n4899), .ZN(n4900) );
  NAND2_X1 U6395 ( .A1(n4900), .A2(SI_12_), .ZN(n4901) );
  NAND2_X1 U6396 ( .A1(n4902), .A2(n4901), .ZN(n5290) );
  MUX2_X1 U6397 ( .A(n6373), .B(n4903), .S(n7554), .Z(n4905) );
  INV_X1 U6398 ( .A(SI_13_), .ZN(n4904) );
  INV_X1 U6399 ( .A(n4905), .ZN(n4906) );
  NAND2_X1 U6400 ( .A1(n4906), .A2(SI_13_), .ZN(n4907) );
  MUX2_X1 U6401 ( .A(n6407), .B(n6405), .S(n7554), .Z(n4909) );
  XNOR2_X1 U6402 ( .A(n4909), .B(SI_14_), .ZN(n5330) );
  INV_X1 U6403 ( .A(n4909), .ZN(n4910) );
  NAND2_X1 U6404 ( .A1(n4910), .A2(SI_14_), .ZN(n4911) );
  MUX2_X1 U6405 ( .A(n9921), .B(n6511), .S(n7548), .Z(n4914) );
  INV_X1 U6406 ( .A(SI_15_), .ZN(n4913) );
  NAND2_X1 U6407 ( .A1(n4914), .A2(n4913), .ZN(n4917) );
  INV_X1 U6408 ( .A(n4914), .ZN(n4915) );
  NAND2_X1 U6409 ( .A1(n4915), .A2(SI_15_), .ZN(n4916) );
  NAND2_X1 U6410 ( .A1(n4917), .A2(n4916), .ZN(n5350) );
  INV_X1 U6411 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n4918) );
  MUX2_X1 U6412 ( .A(n4918), .B(n6556), .S(n7554), .Z(n4920) );
  INV_X1 U6413 ( .A(SI_16_), .ZN(n4919) );
  INV_X1 U6414 ( .A(n4920), .ZN(n4921) );
  NAND2_X1 U6415 ( .A1(n4921), .A2(SI_16_), .ZN(n4922) );
  INV_X1 U6416 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n4924) );
  MUX2_X1 U6417 ( .A(n6594), .B(n4924), .S(n7554), .Z(n4925) );
  XNOR2_X1 U6418 ( .A(n4925), .B(SI_17_), .ZN(n5386) );
  INV_X1 U6419 ( .A(n5386), .ZN(n4927) );
  INV_X1 U6420 ( .A(n4925), .ZN(n4926) );
  MUX2_X1 U6421 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7554), .Z(n4929) );
  XNOR2_X1 U6422 ( .A(n4929), .B(SI_18_), .ZN(n5031) );
  NAND2_X1 U6423 ( .A1(n5032), .A2(n4928), .ZN(n4931) );
  NAND2_X1 U6424 ( .A1(n4929), .A2(SI_18_), .ZN(n4930) );
  MUX2_X1 U6425 ( .A(n6804), .B(n6806), .S(n7548), .Z(n4933) );
  INV_X1 U6426 ( .A(SI_19_), .ZN(n4932) );
  NAND2_X1 U6427 ( .A1(n4933), .A2(n4932), .ZN(n4936) );
  INV_X1 U6428 ( .A(n4933), .ZN(n4934) );
  NAND2_X1 U6429 ( .A1(n4934), .A2(SI_19_), .ZN(n4935) );
  NAND2_X1 U6430 ( .A1(n4936), .A2(n4935), .ZN(n5409) );
  MUX2_X1 U6431 ( .A(n6860), .B(n6836), .S(n7554), .Z(n4938) );
  INV_X1 U6432 ( .A(SI_20_), .ZN(n4937) );
  NAND2_X1 U6433 ( .A1(n4938), .A2(n4937), .ZN(n4941) );
  INV_X1 U6434 ( .A(n4938), .ZN(n4939) );
  NAND2_X1 U6435 ( .A1(n4939), .A2(SI_20_), .ZN(n4940) );
  MUX2_X1 U6436 ( .A(n6905), .B(n6903), .S(n7548), .Z(n4942) );
  XNOR2_X1 U6437 ( .A(n4942), .B(SI_21_), .ZN(n5447) );
  INV_X1 U6438 ( .A(n4942), .ZN(n4943) );
  NAND2_X1 U6439 ( .A1(n4943), .A2(SI_21_), .ZN(n4944) );
  NAND2_X1 U6440 ( .A1(n4945), .A2(n4944), .ZN(n5467) );
  MUX2_X1 U6441 ( .A(n7627), .B(n6981), .S(n7554), .Z(n4947) );
  INV_X1 U6442 ( .A(SI_22_), .ZN(n4946) );
  NAND2_X1 U6443 ( .A1(n4947), .A2(n4946), .ZN(n4950) );
  INV_X1 U6444 ( .A(n4947), .ZN(n4948) );
  NAND2_X1 U6445 ( .A1(n4948), .A2(SI_22_), .ZN(n4949) );
  NAND2_X1 U6446 ( .A1(n4950), .A2(n4949), .ZN(n5466) );
  INV_X1 U6447 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n4951) );
  MUX2_X1 U6448 ( .A(n4951), .B(n9965), .S(n7554), .Z(n4953) );
  INV_X1 U6449 ( .A(SI_23_), .ZN(n4952) );
  NAND2_X1 U6450 ( .A1(n4953), .A2(n4952), .ZN(n5493) );
  INV_X1 U6451 ( .A(n4953), .ZN(n4954) );
  NAND2_X1 U6452 ( .A1(n4954), .A2(SI_23_), .ZN(n4955) );
  NAND2_X1 U6453 ( .A1(n4296), .A2(n5150), .ZN(n5033) );
  INV_X1 U6454 ( .A(n5033), .ZN(n4968) );
  NOR2_X1 U6455 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4961) );
  NOR2_X1 U6456 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4960) );
  NAND4_X1 U6457 ( .A1(n4961), .A2(n4960), .A3(n5388), .A4(n4959), .ZN(n4966)
         );
  NAND4_X1 U6458 ( .A1(n4964), .A2(n4963), .A3(n5335), .A4(n4962), .ZN(n4965)
         );
  NOR2_X1 U6459 ( .A1(n4966), .A2(n4965), .ZN(n4967) );
  INV_X1 U6460 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4972) );
  NAND2_X1 U6461 ( .A1(n4991), .A2(n4974), .ZN(n5007) );
  NAND2_X1 U6462 ( .A1(n5007), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4975) );
  NAND2_X1 U6463 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n4976) );
  NAND2_X1 U6464 ( .A1(n4978), .A2(n4976), .ZN(n4977) );
  INV_X1 U6465 ( .A(n4978), .ZN(n4979) );
  NAND2_X2 U6466 ( .A1(n5657), .A2(n6284), .ZN(n5066) );
  NAND2_X2 U6467 ( .A1(n5066), .A2(n7548), .ZN(n5096) );
  INV_X2 U6468 ( .A(n5096), .ZN(n5229) );
  NAND2_X1 U6469 ( .A1(n7072), .A2(n5229), .ZN(n4981) );
  BUF_X4 U6470 ( .A(n5093), .Z(n8635) );
  OR2_X1 U6471 ( .A1(n8635), .A2(n9965), .ZN(n4980) );
  NAND2_X1 U6472 ( .A1(n4989), .A2(n4988), .ZN(n4983) );
  INV_X1 U6473 ( .A(n4986), .ZN(n4984) );
  NAND2_X1 U6474 ( .A1(n4984), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n4987) );
  XNOR2_X1 U6475 ( .A(n4989), .B(n4988), .ZN(n6837) );
  INV_X1 U6476 ( .A(n6439), .ZN(n6442) );
  NAND2_X1 U6477 ( .A1(n4990), .A2(n4991), .ZN(n4992) );
  XNOR2_X1 U6478 ( .A(n4990), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U6479 ( .A1(n5011), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4994) );
  XNOR2_X1 U6480 ( .A(n4994), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5642) );
  AND2_X1 U6481 ( .A1(n5625), .A2(n5642), .ZN(n4995) );
  INV_X1 U6482 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8568) );
  INV_X1 U6483 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5451) );
  INV_X1 U6484 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5005) );
  NAND2_X1 U6485 ( .A1(n5473), .A2(n5005), .ZN(n5006) );
  NAND2_X1 U6486 ( .A1(n5499), .A2(n5006), .ZN(n9102) );
  INV_X1 U6487 ( .A(n5007), .ZN(n5009) );
  NOR2_X1 U6488 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5008) );
  NAND2_X1 U6489 ( .A1(n5009), .A2(n5008), .ZN(n5010) );
  XNOR2_X2 U6490 ( .A(n5017), .B(n5016), .ZN(n5020) );
  AND2_X4 U6491 ( .A1(n5019), .A2(n5018), .ZN(n5578) );
  INV_X1 U6492 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5023) );
  AND2_X4 U6493 ( .A1(n5020), .A2(n5018), .ZN(n6267) );
  NAND2_X1 U6494 ( .A1(n8625), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5022) );
  INV_X2 U6495 ( .A(n5581), .ZN(n8626) );
  NAND2_X1 U6496 ( .A1(n8626), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5021) );
  OAI211_X1 U6497 ( .C1(n5023), .C2(n8629), .A(n5022), .B(n5021), .ZN(n5024)
         );
  INV_X1 U6498 ( .A(n5024), .ZN(n5025) );
  NAND2_X1 U6499 ( .A1(n5029), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5030) );
  XNOR2_X2 U6500 ( .A(n5030), .B(n4969), .ZN(n9646) );
  INV_X2 U6501 ( .A(n5102), .ZN(n5590) );
  OAI22_X1 U6502 ( .A1(n9105), .A2(n5461), .B1(n8966), .B2(n5590), .ZN(n8508)
         );
  XNOR2_X1 U6503 ( .A(n5032), .B(n5031), .ZN(n6678) );
  NAND2_X1 U6504 ( .A1(n6678), .A2(n5229), .ZN(n5040) );
  INV_X1 U6505 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5035) );
  NAND2_X1 U6506 ( .A1(n5272), .A2(n5035), .ZN(n5292) );
  NOR2_X1 U6507 ( .A1(n5316), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5333) );
  NOR2_X1 U6508 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5036) );
  NAND2_X1 U6509 ( .A1(n5333), .A2(n5036), .ZN(n5369) );
  OR2_X1 U6510 ( .A1(n5369), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n5037) );
  NAND2_X1 U6511 ( .A1(n5037), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U6512 ( .A1(n5389), .A2(n5388), .ZN(n5390) );
  NAND2_X1 U6513 ( .A1(n5390), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5038) );
  XNOR2_X1 U6514 ( .A(n5038), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9630) );
  AOI22_X1 U6515 ( .A1(n5412), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9630), .B2(
        n5411), .ZN(n5039) );
  INV_X1 U6516 ( .A(n9308), .ZN(n9179) );
  INV_X1 U6517 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n10030) );
  NAND2_X1 U6518 ( .A1(n5396), .A2(n10030), .ZN(n5042) );
  NAND2_X1 U6519 ( .A1(n5416), .A2(n5042), .ZN(n9176) );
  OR2_X1 U6520 ( .A1(n9176), .A2(n5658), .ZN(n5045) );
  AOI22_X1 U6521 ( .A1(n8625), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n6268), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5044) );
  NAND2_X1 U6522 ( .A1(n6267), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5043) );
  OAI22_X1 U6523 ( .A1(n9179), .A2(n5480), .B1(n8647), .B2(n5461), .ZN(n5048)
         );
  NAND2_X1 U6524 ( .A1(n5046), .A2(n9646), .ZN(n5047) );
  AND2_X2 U6525 ( .A1(n5047), .A2(n6439), .ZN(n5588) );
  INV_X2 U6526 ( .A(n5588), .ZN(n5620) );
  NAND2_X1 U6527 ( .A1(n5578), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5052) );
  NAND2_X1 U6528 ( .A1(n5085), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5051) );
  NAND2_X1 U6529 ( .A1(n6267), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5050) );
  NAND2_X1 U6530 ( .A1(n5086), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5049) );
  NAND4_X2 U6531 ( .A1(n5052), .A2(n5051), .A3(n5050), .A4(n5049), .ZN(n8892)
         );
  NAND2_X1 U6532 ( .A1(n8892), .A2(n5102), .ZN(n5061) );
  INV_X2 U6533 ( .A(n5161), .ZN(n5208) );
  INV_X1 U6534 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U6535 ( .A1(n7548), .A2(SI_0_), .ZN(n5053) );
  INV_X1 U6536 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9932) );
  NAND2_X1 U6537 ( .A1(n5053), .A2(n9932), .ZN(n5055) );
  AND2_X1 U6538 ( .A1(n5055), .A2(n5054), .ZN(n9365) );
  NAND2_X1 U6539 ( .A1(n5066), .A2(n9365), .ZN(n5056) );
  OR2_X1 U6540 ( .A1(n5057), .A2(n6297), .ZN(n5058) );
  INV_X1 U6541 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5064) );
  NAND2_X1 U6542 ( .A1(n8892), .A2(n5363), .ZN(n5063) );
  NAND2_X1 U6543 ( .A1(n4297), .A2(n4299), .ZN(n5062) );
  OAI211_X1 U6544 ( .C1(n5064), .C2(n5057), .A(n5063), .B(n5062), .ZN(n6324)
         );
  NAND2_X2 U6545 ( .A1(n6325), .A2(n5065), .ZN(n6344) );
  INV_X1 U6546 ( .A(n6298), .ZN(n9495) );
  XNOR2_X1 U6547 ( .A(n5068), .B(n5067), .ZN(n6246) );
  INV_X1 U6548 ( .A(n5093), .ZN(n5069) );
  NAND2_X1 U6549 ( .A1(n5578), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5076) );
  NAND2_X1 U6550 ( .A1(n5086), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5075) );
  NAND2_X1 U6551 ( .A1(n5085), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5073) );
  NAND4_X2 U6552 ( .A1(n5076), .A2(n5075), .A3(n5074), .A4(n5073), .ZN(n8891)
         );
  NAND2_X1 U6553 ( .A1(n8891), .A2(n5208), .ZN(n5077) );
  OAI21_X1 U6554 ( .B1(n6435), .B2(n5041), .A(n5077), .ZN(n5078) );
  XNOR2_X1 U6555 ( .A(n5078), .B(n5588), .ZN(n5081) );
  NAND2_X1 U6556 ( .A1(n6344), .A2(n5081), .ZN(n5080) );
  NAND2_X1 U6557 ( .A1(n8891), .A2(n5622), .ZN(n5079) );
  OAI21_X1 U6558 ( .B1(n6435), .B2(n5161), .A(n5079), .ZN(n6345) );
  NAND2_X1 U6559 ( .A1(n5080), .A2(n6345), .ZN(n5084) );
  INV_X1 U6560 ( .A(n5081), .ZN(n6346) );
  INV_X1 U6561 ( .A(n6344), .ZN(n5082) );
  NAND2_X1 U6562 ( .A1(n6346), .A2(n5082), .ZN(n5083) );
  NAND2_X1 U6563 ( .A1(n5578), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5090) );
  NAND2_X1 U6564 ( .A1(n5085), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5089) );
  NAND2_X1 U6565 ( .A1(n6267), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5088) );
  NAND2_X1 U6566 ( .A1(n5086), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5087) );
  NAND4_X1 U6567 ( .A1(n5090), .A2(n5089), .A3(n5088), .A4(n5087), .ZN(n8889)
         );
  NAND2_X1 U6568 ( .A1(n8889), .A2(n5208), .ZN(n5100) );
  INV_X1 U6569 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5092) );
  OR2_X1 U6570 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5116) );
  NAND2_X1 U6571 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5116), .ZN(n5091) );
  XNOR2_X1 U6572 ( .A(n5092), .B(n5091), .ZN(n9508) );
  XNOR2_X1 U6573 ( .A(n5094), .B(n5095), .ZN(n6263) );
  OR2_X1 U6574 ( .A1(n5096), .A2(n6263), .ZN(n5097) );
  NAND2_X1 U6575 ( .A1(n6457), .A2(n5605), .ZN(n5099) );
  NAND2_X1 U6576 ( .A1(n5100), .A2(n5099), .ZN(n5101) );
  XNOR2_X1 U6577 ( .A(n5101), .B(n5588), .ZN(n5106) );
  NAND2_X1 U6578 ( .A1(n6457), .A2(n5208), .ZN(n5104) );
  NAND2_X1 U6579 ( .A1(n8889), .A2(n5102), .ZN(n5103) );
  INV_X1 U6580 ( .A(n5106), .ZN(n5108) );
  NAND2_X1 U6581 ( .A1(n6364), .A2(n5109), .ZN(n7574) );
  INV_X1 U6582 ( .A(n7574), .ZN(n5110) );
  INV_X1 U6583 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U6584 ( .A1(n5578), .A2(n6473), .ZN(n5115) );
  NAND2_X1 U6585 ( .A1(n8625), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5114) );
  NAND2_X1 U6586 ( .A1(n8626), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U6587 ( .A1(n6267), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5112) );
  AND4_X2 U6588 ( .A1(n5115), .A2(n5114), .A3(n5113), .A4(n5112), .ZN(n6482)
         );
  OAI21_X1 U6589 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(n5116), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5117) );
  XNOR2_X1 U6590 ( .A(n5117), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6390) );
  INV_X1 U6591 ( .A(n6390), .ZN(n6288) );
  XNOR2_X1 U6592 ( .A(n5118), .B(n5119), .ZN(n6261) );
  OR2_X1 U6593 ( .A1(n5096), .A2(n6261), .ZN(n5121) );
  OR2_X1 U6594 ( .A1(n8635), .A2(n6245), .ZN(n5120) );
  OAI211_X2 U6595 ( .C1(n6302), .C2(n6288), .A(n5121), .B(n5120), .ZN(n6498)
         );
  NAND2_X1 U6596 ( .A1(n6498), .A2(n5605), .ZN(n5122) );
  OAI21_X1 U6597 ( .B1(n6482), .B2(n5161), .A(n5122), .ZN(n5123) );
  XNOR2_X1 U6598 ( .A(n5123), .B(n5620), .ZN(n5126) );
  NAND2_X1 U6599 ( .A1(n6498), .A2(n5208), .ZN(n5124) );
  OAI21_X1 U6600 ( .B1(n6482), .B2(n5590), .A(n5124), .ZN(n5125) );
  NAND2_X1 U6601 ( .A1(n5126), .A2(n5125), .ZN(n5127) );
  NAND2_X1 U6602 ( .A1(n8625), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5131) );
  NAND2_X1 U6603 ( .A1(n6268), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5130) );
  XNOR2_X1 U6604 ( .A(n6473), .B(P1_REG3_REG_4__SCAN_IN), .ZN(n6414) );
  NAND2_X1 U6605 ( .A1(n5578), .A2(n6414), .ZN(n5129) );
  NAND2_X1 U6606 ( .A1(n6267), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5128) );
  OR2_X1 U6607 ( .A1(n5150), .A2(n5332), .ZN(n5132) );
  XNOR2_X1 U6608 ( .A(n5132), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9531) );
  INV_X1 U6609 ( .A(n9531), .ZN(n6248) );
  XNOR2_X1 U6610 ( .A(n5134), .B(n5133), .ZN(n6257) );
  OR2_X1 U6611 ( .A1(n5096), .A2(n6257), .ZN(n5136) );
  OR2_X1 U6612 ( .A1(n8635), .A2(n6249), .ZN(n5135) );
  NAND2_X1 U6613 ( .A1(n6560), .A2(n5605), .ZN(n5137) );
  OAI21_X1 U6614 ( .B1(n6574), .B2(n5461), .A(n5137), .ZN(n5138) );
  XNOR2_X1 U6615 ( .A(n5138), .B(n5588), .ZN(n5140) );
  NAND2_X1 U6616 ( .A1(n6560), .A2(n5208), .ZN(n5139) );
  OAI21_X1 U6617 ( .B1(n6574), .B2(n5590), .A(n5139), .ZN(n5141) );
  XNOR2_X1 U6618 ( .A(n5140), .B(n5141), .ZN(n6417) );
  NAND2_X1 U6619 ( .A1(n6416), .A2(n6417), .ZN(n6415) );
  INV_X1 U6620 ( .A(n5140), .ZN(n5142) );
  OR2_X1 U6621 ( .A1(n5142), .A2(n5141), .ZN(n5143) );
  NAND2_X1 U6622 ( .A1(n6415), .A2(n5143), .ZN(n5164) );
  NAND2_X1 U6623 ( .A1(n8625), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U6624 ( .A1(n8626), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5147) );
  AOI21_X1 U6625 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5144) );
  NOR2_X1 U6626 ( .A1(n5144), .A2(n5173), .ZN(n6570) );
  NAND2_X1 U6627 ( .A1(n5578), .A2(n6570), .ZN(n5146) );
  NAND2_X1 U6628 ( .A1(n6267), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5145) );
  NAND2_X1 U6629 ( .A1(n5150), .A2(n5149), .ZN(n5151) );
  NOR2_X1 U6630 ( .A1(n5151), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5193) );
  INV_X1 U6631 ( .A(n5193), .ZN(n5155) );
  NAND2_X1 U6632 ( .A1(n5151), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5153) );
  MUX2_X1 U6633 ( .A(n5153), .B(P1_IR_REG_31__SCAN_IN), .S(n5152), .Z(n5154)
         );
  INV_X1 U6634 ( .A(n6392), .ZN(n9542) );
  OR2_X1 U6635 ( .A1(n8635), .A2(n6250), .ZN(n5159) );
  XNOR2_X1 U6636 ( .A(n5156), .B(n5157), .ZN(n6259) );
  OR2_X1 U6637 ( .A1(n5096), .A2(n6259), .ZN(n5158) );
  OAI211_X1 U6638 ( .C1(n6302), .C2(n9542), .A(n5159), .B(n5158), .ZN(n9641)
         );
  NAND2_X1 U6639 ( .A1(n9641), .A2(n5605), .ZN(n5160) );
  OAI21_X1 U6640 ( .B1(n6538), .B2(n5161), .A(n5160), .ZN(n5162) );
  XNOR2_X1 U6641 ( .A(n5162), .B(n5588), .ZN(n5163) );
  OR2_X1 U6642 ( .A1(n6538), .A2(n5590), .ZN(n5166) );
  NAND2_X1 U6643 ( .A1(n9641), .A2(n5208), .ZN(n5165) );
  AND2_X1 U6644 ( .A1(n5166), .A2(n5165), .ZN(n6572) );
  XNOR2_X1 U6645 ( .A(n5167), .B(n5168), .ZN(n6255) );
  OR2_X1 U6646 ( .A1(n6255), .A2(n5096), .ZN(n5172) );
  OR2_X1 U6647 ( .A1(n5193), .A2(n5332), .ZN(n5169) );
  XNOR2_X1 U6648 ( .A(n5169), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9567) );
  INV_X1 U6649 ( .A(n9567), .ZN(n6252) );
  OR2_X1 U6650 ( .A1(n6302), .A2(n6252), .ZN(n5171) );
  OR2_X1 U6651 ( .A1(n8635), .A2(n6253), .ZN(n5170) );
  NAND2_X1 U6652 ( .A1(n6267), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U6653 ( .A1(n8625), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5177) );
  NOR2_X1 U6654 ( .A1(n5173), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5174) );
  NOR2_X1 U6655 ( .A1(n5197), .A2(n5174), .ZN(n6637) );
  NAND2_X1 U6656 ( .A1(n5578), .A2(n6637), .ZN(n5176) );
  NAND2_X1 U6657 ( .A1(n6268), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5175) );
  NAND4_X1 U6658 ( .A1(n5178), .A2(n5177), .A3(n5176), .A4(n5175), .ZN(n8885)
         );
  NAND2_X1 U6659 ( .A1(n8885), .A2(n5617), .ZN(n5179) );
  OAI21_X1 U6660 ( .B1(n6641), .B2(n5480), .A(n5179), .ZN(n5180) );
  XNOR2_X1 U6661 ( .A(n5180), .B(n5588), .ZN(n5183) );
  OR2_X1 U6662 ( .A1(n6641), .A2(n5461), .ZN(n5182) );
  NAND2_X1 U6663 ( .A1(n8885), .A2(n5622), .ZN(n5181) );
  AND2_X1 U6664 ( .A1(n5182), .A2(n5181), .ZN(n5184) );
  NAND2_X1 U6665 ( .A1(n5183), .A2(n5184), .ZN(n5189) );
  INV_X1 U6666 ( .A(n5183), .ZN(n5186) );
  INV_X1 U6667 ( .A(n5184), .ZN(n5185) );
  NAND2_X1 U6668 ( .A1(n5186), .A2(n5185), .ZN(n5187) );
  AND2_X1 U6669 ( .A1(n5189), .A2(n5187), .ZN(n6628) );
  NAND2_X1 U6670 ( .A1(n6630), .A2(n5189), .ZN(n6668) );
  XNOR2_X1 U6671 ( .A(n5190), .B(n5191), .ZN(n6265) );
  NAND2_X1 U6672 ( .A1(n6265), .A2(n5229), .ZN(n5196) );
  NAND2_X1 U6673 ( .A1(n5193), .A2(n5192), .ZN(n5230) );
  NAND2_X1 U6674 ( .A1(n5230), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5194) );
  XNOR2_X1 U6675 ( .A(n5194), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9571) );
  AOI22_X1 U6676 ( .A1(n5412), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5411), .B2(
        n9571), .ZN(n5195) );
  NAND2_X1 U6677 ( .A1(n5196), .A2(n5195), .ZN(n6840) );
  NAND2_X1 U6678 ( .A1(n6840), .A2(n5605), .ZN(n5206) );
  NAND2_X1 U6679 ( .A1(n8625), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5204) );
  NAND2_X1 U6680 ( .A1(n8626), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5203) );
  NAND2_X1 U6681 ( .A1(n6267), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5202) );
  INV_X1 U6682 ( .A(n5197), .ZN(n5199) );
  INV_X1 U6683 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6684 ( .A1(n5199), .A2(n5198), .ZN(n5200) );
  NAND2_X1 U6685 ( .A1(n5234), .A2(n5200), .ZN(n6660) );
  INV_X1 U6686 ( .A(n6660), .ZN(n6670) );
  NAND2_X1 U6687 ( .A1(n5578), .A2(n6670), .ZN(n5201) );
  OR2_X1 U6688 ( .A1(n6839), .A2(n5461), .ZN(n5205) );
  NAND2_X1 U6689 ( .A1(n5206), .A2(n5205), .ZN(n5207) );
  XNOR2_X1 U6690 ( .A(n5207), .B(n5588), .ZN(n5213) );
  NAND2_X1 U6691 ( .A1(n6840), .A2(n5208), .ZN(n5210) );
  OR2_X1 U6692 ( .A1(n6839), .A2(n5590), .ZN(n5209) );
  NAND2_X1 U6693 ( .A1(n5210), .A2(n5209), .ZN(n5211) );
  XNOR2_X1 U6694 ( .A(n5213), .B(n5211), .ZN(n6669) );
  INV_X1 U6695 ( .A(n5211), .ZN(n5212) );
  NAND2_X1 U6696 ( .A1(n5213), .A2(n5212), .ZN(n5214) );
  XNOR2_X1 U6697 ( .A(n5215), .B(n4840), .ZN(n6280) );
  NAND2_X1 U6698 ( .A1(n6280), .A2(n5229), .ZN(n5219) );
  NAND2_X1 U6699 ( .A1(n5034), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5216) );
  MUX2_X1 U6700 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5216), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n5217) );
  AOI22_X1 U6701 ( .A1(n5412), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5411), .B2(
        n9600), .ZN(n5218) );
  NAND2_X1 U6702 ( .A1(n5236), .A2(n5220), .ZN(n5221) );
  AND2_X1 U6703 ( .A1(n5258), .A2(n5221), .ZN(n6933) );
  NAND2_X1 U6704 ( .A1(n5578), .A2(n6933), .ZN(n5225) );
  NAND2_X1 U6705 ( .A1(n8625), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6706 ( .A1(n8626), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5223) );
  NAND2_X1 U6707 ( .A1(n6267), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5222) );
  OAI22_X1 U6708 ( .A1(n6993), .A2(n5480), .B1(n9393), .B2(n5461), .ZN(n5226)
         );
  XNOR2_X1 U6709 ( .A(n5226), .B(n5620), .ZN(n5249) );
  OAI22_X1 U6710 ( .A1(n6993), .A2(n5461), .B1(n9393), .B2(n5590), .ZN(n5248)
         );
  NAND2_X1 U6711 ( .A1(n5249), .A2(n5248), .ZN(n6914) );
  XNOR2_X1 U6712 ( .A(n5227), .B(n5228), .ZN(n6276) );
  NAND2_X1 U6713 ( .A1(n6276), .A2(n5229), .ZN(n5233) );
  OAI21_X1 U6714 ( .B1(n5230), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5231) );
  XNOR2_X1 U6715 ( .A(n5231), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9584) );
  AOI22_X1 U6716 ( .A1(n5412), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5411), .B2(
        n9584), .ZN(n5232) );
  NAND2_X1 U6717 ( .A1(n6970), .A2(n5605), .ZN(n5242) );
  NAND2_X1 U6718 ( .A1(n8625), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U6719 ( .A1(n6267), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5239) );
  INV_X1 U6720 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6893) );
  NAND2_X1 U6721 ( .A1(n5234), .A2(n6893), .ZN(n5235) );
  AND2_X1 U6722 ( .A1(n5236), .A2(n5235), .ZN(n6894) );
  NAND2_X1 U6723 ( .A1(n5578), .A2(n6894), .ZN(n5238) );
  NAND2_X1 U6724 ( .A1(n8626), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5237) );
  OR2_X1 U6725 ( .A1(n6926), .A2(n5461), .ZN(n5241) );
  NAND2_X1 U6726 ( .A1(n5242), .A2(n5241), .ZN(n5243) );
  XNOR2_X1 U6727 ( .A(n5243), .B(n5588), .ZN(n5247) );
  INV_X1 U6728 ( .A(n5247), .ZN(n6889) );
  NOR2_X1 U6729 ( .A1(n6926), .A2(n5590), .ZN(n5244) );
  AOI21_X1 U6730 ( .B1(n6970), .B2(n5617), .A(n5244), .ZN(n6888) );
  INV_X1 U6731 ( .A(n6888), .ZN(n5245) );
  NAND2_X1 U6732 ( .A1(n6889), .A2(n5245), .ZN(n5246) );
  AND2_X1 U6733 ( .A1(n6914), .A2(n5246), .ZN(n5251) );
  NAND3_X1 U6734 ( .A1(n6914), .A2(n6888), .A3(n5247), .ZN(n5250) );
  OR2_X1 U6735 ( .A1(n5249), .A2(n5248), .ZN(n6946) );
  XNOR2_X1 U6736 ( .A(n5252), .B(n4839), .ZN(n6309) );
  NAND2_X1 U6737 ( .A1(n6309), .A2(n5229), .ZN(n5256) );
  NAND2_X1 U6738 ( .A1(n5253), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5254) );
  XNOR2_X1 U6739 ( .A(n5254), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6427) );
  AOI22_X1 U6740 ( .A1(n5412), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5411), .B2(
        n6427), .ZN(n5255) );
  NAND2_X1 U6741 ( .A1(n5256), .A2(n5255), .ZN(n9407) );
  NAND2_X1 U6742 ( .A1(n9407), .A2(n5605), .ZN(n5265) );
  NAND2_X1 U6743 ( .A1(n8625), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5263) );
  NAND2_X1 U6744 ( .A1(n6268), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U6745 ( .A1(n5258), .A2(n5257), .ZN(n5259) );
  AND2_X1 U6746 ( .A1(n5277), .A2(n5259), .ZN(n9403) );
  NAND2_X1 U6747 ( .A1(n5578), .A2(n9403), .ZN(n5261) );
  NAND2_X1 U6748 ( .A1(n6267), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5260) );
  OR2_X1 U6749 ( .A1(n6996), .A2(n5461), .ZN(n5264) );
  NAND2_X1 U6750 ( .A1(n5265), .A2(n5264), .ZN(n5266) );
  XNOR2_X1 U6751 ( .A(n5266), .B(n5588), .ZN(n5288) );
  NOR2_X1 U6752 ( .A1(n6996), .A2(n5590), .ZN(n5267) );
  AOI21_X1 U6753 ( .B1(n9407), .B2(n5617), .A(n5267), .ZN(n5287) );
  XNOR2_X1 U6754 ( .A(n5288), .B(n5287), .ZN(n6945) );
  INV_X1 U6755 ( .A(n6945), .ZN(n5268) );
  XNOR2_X1 U6756 ( .A(n5271), .B(n5270), .ZN(n6313) );
  NAND2_X1 U6757 ( .A1(n6313), .A2(n5229), .ZN(n5275) );
  OR2_X1 U6758 ( .A1(n5272), .A2(n5332), .ZN(n5273) );
  XNOR2_X1 U6759 ( .A(n5273), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6608) );
  AOI22_X1 U6760 ( .A1(n5412), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5411), .B2(
        n6608), .ZN(n5274) );
  NAND2_X1 U6761 ( .A1(n7012), .A2(n5605), .ZN(n5284) );
  NAND2_X1 U6762 ( .A1(n8625), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5282) );
  INV_X1 U6763 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5276) );
  NAND2_X1 U6764 ( .A1(n5277), .A2(n5276), .ZN(n5278) );
  AND2_X1 U6765 ( .A1(n5297), .A2(n5278), .ZN(n7023) );
  NAND2_X1 U6766 ( .A1(n5578), .A2(n7023), .ZN(n5281) );
  NAND2_X1 U6767 ( .A1(n6267), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U6768 ( .A1(n8626), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5279) );
  NAND4_X1 U6769 ( .A1(n5282), .A2(n5281), .A3(n5280), .A4(n5279), .ZN(n8880)
         );
  NAND2_X1 U6770 ( .A1(n8880), .A2(n5617), .ZN(n5283) );
  NAND2_X1 U6771 ( .A1(n5284), .A2(n5283), .ZN(n5285) );
  XNOR2_X1 U6772 ( .A(n5285), .B(n5620), .ZN(n5309) );
  AND2_X1 U6773 ( .A1(n8880), .A2(n5622), .ZN(n5286) );
  AOI21_X1 U6774 ( .B1(n7012), .B2(n5617), .A(n5286), .ZN(n5307) );
  XNOR2_X1 U6775 ( .A(n5309), .B(n5307), .ZN(n6863) );
  NAND2_X1 U6776 ( .A1(n5288), .A2(n5287), .ZN(n6861) );
  AND2_X1 U6777 ( .A1(n6863), .A2(n6861), .ZN(n5289) );
  XNOR2_X1 U6778 ( .A(n5291), .B(n5290), .ZN(n6317) );
  NAND2_X1 U6779 ( .A1(n6317), .A2(n5229), .ZN(n5295) );
  NAND2_X1 U6780 ( .A1(n5292), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5293) );
  XNOR2_X1 U6781 ( .A(n5293), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6688) );
  AOI22_X1 U6782 ( .A1(n5412), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5411), .B2(
        n6688), .ZN(n5294) );
  NAND2_X1 U6783 ( .A1(n7311), .A2(n5605), .ZN(n5304) );
  NAND2_X1 U6784 ( .A1(n6267), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5302) );
  NAND2_X1 U6785 ( .A1(n8625), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5301) );
  INV_X1 U6786 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5296) );
  NAND2_X1 U6787 ( .A1(n5297), .A2(n5296), .ZN(n5298) );
  AND2_X1 U6788 ( .A1(n5321), .A2(n5298), .ZN(n7017) );
  NAND2_X1 U6789 ( .A1(n5578), .A2(n7017), .ZN(n5300) );
  NAND2_X1 U6790 ( .A1(n8626), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5299) );
  OR2_X1 U6791 ( .A1(n7327), .A2(n5461), .ZN(n5303) );
  NAND2_X1 U6792 ( .A1(n5304), .A2(n5303), .ZN(n5305) );
  XNOR2_X1 U6793 ( .A(n5305), .B(n5620), .ZN(n5311) );
  NOR2_X1 U6794 ( .A1(n7327), .A2(n5590), .ZN(n5306) );
  AOI21_X1 U6795 ( .B1(n7311), .B2(n5617), .A(n5306), .ZN(n5312) );
  XNOR2_X1 U6796 ( .A(n5311), .B(n5312), .ZN(n6906) );
  INV_X1 U6797 ( .A(n5307), .ZN(n5308) );
  NAND2_X1 U6798 ( .A1(n5309), .A2(n5308), .ZN(n6907) );
  AND2_X1 U6799 ( .A1(n6906), .A2(n6907), .ZN(n5310) );
  INV_X1 U6800 ( .A(n5311), .ZN(n5313) );
  NAND2_X1 U6801 ( .A1(n5313), .A2(n5312), .ZN(n5314) );
  XNOR2_X1 U6802 ( .A(n5315), .B(n4836), .ZN(n5938) );
  NAND2_X1 U6803 ( .A1(n5938), .A2(n5229), .ZN(n5319) );
  NAND2_X1 U6804 ( .A1(n5316), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5317) );
  XNOR2_X1 U6805 ( .A(n5317), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7145) );
  AOI22_X1 U6806 ( .A1(n5412), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5411), .B2(
        n7145), .ZN(n5318) );
  NAND2_X1 U6807 ( .A1(n6267), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6808 ( .A1(n8625), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U6809 ( .A1(n5321), .A2(n5320), .ZN(n5322) );
  AND2_X1 U6810 ( .A1(n5339), .A2(n5322), .ZN(n6986) );
  NAND2_X1 U6811 ( .A1(n5578), .A2(n6986), .ZN(n5324) );
  NAND2_X1 U6812 ( .A1(n8626), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5323) );
  OAI22_X1 U6813 ( .A1(n8689), .A2(n5480), .B1(n7314), .B2(n5461), .ZN(n5327)
         );
  XNOR2_X1 U6814 ( .A(n5327), .B(n5620), .ZN(n5329) );
  OAI22_X1 U6815 ( .A1(n8689), .A2(n5461), .B1(n7314), .B2(n5590), .ZN(n5328)
         );
  OR2_X1 U6816 ( .A1(n5329), .A2(n5328), .ZN(n6983) );
  AND2_X1 U6817 ( .A1(n5329), .A2(n5328), .ZN(n6984) );
  XNOR2_X1 U6818 ( .A(n5331), .B(n5330), .ZN(n6404) );
  OR2_X1 U6819 ( .A1(n5333), .A2(n5332), .ZN(n5336) );
  INV_X1 U6820 ( .A(n5336), .ZN(n5334) );
  NAND2_X1 U6821 ( .A1(n5334), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5337) );
  NAND2_X1 U6822 ( .A1(n5336), .A2(n5335), .ZN(n5352) );
  AOI22_X1 U6823 ( .A1(n5412), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5411), .B2(
        n9608), .ZN(n5338) );
  NAND2_X1 U6824 ( .A1(n8625), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5344) );
  NAND2_X1 U6825 ( .A1(n6267), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5343) );
  INV_X1 U6826 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n10020) );
  NAND2_X1 U6827 ( .A1(n5339), .A2(n10020), .ZN(n5340) );
  AND2_X1 U6828 ( .A1(n5357), .A2(n5340), .ZN(n7317) );
  NAND2_X1 U6829 ( .A1(n5578), .A2(n7317), .ZN(n5342) );
  NAND2_X1 U6830 ( .A1(n8626), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5341) );
  OAI22_X1 U6831 ( .A1(n9473), .A2(n5480), .B1(n8954), .B2(n5461), .ZN(n5345)
         );
  XNOR2_X1 U6832 ( .A(n5345), .B(n5588), .ZN(n5347) );
  AOI22_X1 U6833 ( .A1(n8955), .A2(n5617), .B1(n5622), .B2(n4509), .ZN(n7170)
         );
  INV_X1 U6834 ( .A(n5346), .ZN(n5349) );
  INV_X1 U6835 ( .A(n5347), .ZN(n5348) );
  XNOR2_X1 U6836 ( .A(n5351), .B(n5350), .ZN(n6510) );
  NAND2_X1 U6837 ( .A1(n6510), .A2(n5229), .ZN(n5356) );
  NAND2_X1 U6838 ( .A1(n5352), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5354) );
  INV_X1 U6839 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5353) );
  XNOR2_X1 U6840 ( .A(n5354), .B(n5353), .ZN(n8900) );
  INV_X1 U6841 ( .A(n8900), .ZN(n7149) );
  AOI22_X1 U6842 ( .A1(n5412), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5411), .B2(
        n7149), .ZN(n5355) );
  NAND2_X1 U6843 ( .A1(n6267), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6844 ( .A1(n8625), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6845 ( .A1(n5357), .A2(n7148), .ZN(n5358) );
  AND2_X1 U6846 ( .A1(n5374), .A2(n5358), .ZN(n9226) );
  NAND2_X1 U6847 ( .A1(n5578), .A2(n9226), .ZN(n5360) );
  NAND2_X1 U6848 ( .A1(n8626), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5359) );
  OAI22_X1 U6849 ( .A1(n9228), .A2(n5480), .B1(n9210), .B2(n5461), .ZN(n5364)
         );
  XNOR2_X1 U6850 ( .A(n5364), .B(n5620), .ZN(n5365) );
  INV_X1 U6851 ( .A(n9210), .ZN(n8958) );
  AOI22_X1 U6852 ( .A1(n9322), .A2(n5617), .B1(n5622), .B2(n8958), .ZN(n8608)
         );
  NAND2_X1 U6853 ( .A1(n5366), .A2(n5365), .ZN(n8606) );
  XNOR2_X1 U6854 ( .A(n5368), .B(n5367), .ZN(n6508) );
  NAND2_X1 U6855 ( .A1(n6508), .A2(n5229), .ZN(n5372) );
  NAND2_X1 U6856 ( .A1(n5369), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5370) );
  XNOR2_X1 U6857 ( .A(n5370), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8919) );
  AOI22_X1 U6858 ( .A1(n5412), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5411), .B2(
        n8919), .ZN(n5371) );
  INV_X1 U6859 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U6860 ( .A1(n5374), .A2(n5373), .ZN(n5375) );
  AND2_X1 U6861 ( .A1(n5394), .A2(n5375), .ZN(n9214) );
  NAND2_X1 U6862 ( .A1(n9214), .A2(n5578), .ZN(n5379) );
  NAND2_X1 U6863 ( .A1(n8625), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U6864 ( .A1(n6268), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U6865 ( .A1(n6267), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5376) );
  NAND4_X1 U6866 ( .A1(n5379), .A2(n5378), .A3(n5377), .A4(n5376), .ZN(n9233)
         );
  AOI22_X1 U6867 ( .A1(n9319), .A2(n5617), .B1(n5622), .B2(n9233), .ZN(n5384)
         );
  NAND2_X1 U6868 ( .A1(n9319), .A2(n5605), .ZN(n5381) );
  NAND2_X1 U6869 ( .A1(n9233), .A2(n5617), .ZN(n5380) );
  NAND2_X1 U6870 ( .A1(n5381), .A2(n5380), .ZN(n5382) );
  XNOR2_X1 U6871 ( .A(n5382), .B(n5620), .ZN(n5383) );
  XOR2_X1 U6872 ( .A(n5384), .B(n5383), .Z(n8539) );
  NOR2_X1 U6873 ( .A1(n8538), .A2(n8539), .ZN(n8537) );
  INV_X1 U6874 ( .A(n5383), .ZN(n5385) );
  XNOR2_X1 U6875 ( .A(n5387), .B(n5386), .ZN(n6557) );
  NAND2_X1 U6876 ( .A1(n6557), .A2(n5229), .ZN(n5393) );
  OR2_X1 U6877 ( .A1(n5389), .A2(n5388), .ZN(n5391) );
  AOI22_X1 U6878 ( .A1(n5412), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5411), .B2(
        n8930), .ZN(n5392) );
  NAND2_X1 U6879 ( .A1(n9312), .A2(n5605), .ZN(n5402) );
  NAND2_X1 U6880 ( .A1(n5394), .A2(n8549), .ZN(n5395) );
  NAND2_X1 U6881 ( .A1(n5396), .A2(n5395), .ZN(n9192) );
  NAND2_X1 U6882 ( .A1(n8625), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U6883 ( .A1(n6267), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5397) );
  AND2_X1 U6884 ( .A1(n5398), .A2(n5397), .ZN(n5400) );
  NAND2_X1 U6885 ( .A1(n8626), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5399) );
  OAI211_X1 U6886 ( .C1(n9192), .C2(n5658), .A(n5400), .B(n5399), .ZN(n9182)
         );
  NAND2_X1 U6887 ( .A1(n9182), .A2(n5617), .ZN(n5401) );
  NAND2_X1 U6888 ( .A1(n5402), .A2(n5401), .ZN(n5403) );
  XNOR2_X1 U6889 ( .A(n5403), .B(n5620), .ZN(n5405) );
  INV_X1 U6890 ( .A(n9312), .ZN(n9195) );
  INV_X1 U6891 ( .A(n9182), .ZN(n9211) );
  OAI22_X1 U6892 ( .A1(n9195), .A2(n5461), .B1(n9211), .B2(n5590), .ZN(n5406)
         );
  XNOR2_X1 U6893 ( .A(n5405), .B(n5406), .ZN(n8547) );
  INV_X1 U6894 ( .A(n8547), .ZN(n5404) );
  INV_X1 U6895 ( .A(n5405), .ZN(n5408) );
  INV_X1 U6896 ( .A(n5406), .ZN(n5407) );
  OAI22_X1 U6897 ( .A1(n9179), .A2(n5461), .B1(n8647), .B2(n5590), .ZN(n8584)
         );
  XNOR2_X1 U6898 ( .A(n5410), .B(n5409), .ZN(n6803) );
  NAND2_X1 U6899 ( .A1(n6803), .A2(n5229), .ZN(n5414) );
  AOI22_X1 U6900 ( .A1(n5412), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4797), .B2(
        n5411), .ZN(n5413) );
  NAND2_X1 U6901 ( .A1(n9302), .A2(n5605), .ZN(n5424) );
  INV_X1 U6902 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U6903 ( .A1(n5416), .A2(n5415), .ZN(n5417) );
  NAND2_X1 U6904 ( .A1(n5432), .A2(n5417), .ZN(n9160) );
  OR2_X1 U6905 ( .A1(n9160), .A2(n5658), .ZN(n5422) );
  INV_X1 U6906 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8931) );
  NAND2_X1 U6907 ( .A1(n8625), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U6908 ( .A1(n6268), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5418) );
  OAI211_X1 U6909 ( .C1(n8629), .C2(n8931), .A(n5419), .B(n5418), .ZN(n5420)
         );
  INV_X1 U6910 ( .A(n5420), .ZN(n5421) );
  NAND2_X1 U6911 ( .A1(n5422), .A2(n5421), .ZN(n9183) );
  NAND2_X1 U6912 ( .A1(n9183), .A2(n5617), .ZN(n5423) );
  NAND2_X1 U6913 ( .A1(n5424), .A2(n5423), .ZN(n5425) );
  XNOR2_X1 U6914 ( .A(n5425), .B(n5620), .ZN(n5427) );
  OAI22_X1 U6915 ( .A1(n9163), .A2(n5461), .B1(n8961), .B2(n5590), .ZN(n5426)
         );
  XNOR2_X1 U6916 ( .A(n5427), .B(n5426), .ZN(n8516) );
  XNOR2_X1 U6917 ( .A(n5429), .B(n5428), .ZN(n6835) );
  NAND2_X1 U6918 ( .A1(n6835), .A2(n5229), .ZN(n5431) );
  OR2_X1 U6919 ( .A1(n8635), .A2(n6836), .ZN(n5430) );
  NAND2_X1 U6920 ( .A1(n9297), .A2(n5605), .ZN(n5441) );
  NAND2_X1 U6921 ( .A1(n5432), .A2(n8568), .ZN(n5433) );
  NAND2_X1 U6922 ( .A1(n5452), .A2(n5433), .ZN(n9145) );
  OR2_X1 U6923 ( .A1(n9145), .A2(n5658), .ZN(n5439) );
  INV_X1 U6924 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U6925 ( .A1(n6268), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U6926 ( .A1(n8625), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5434) );
  OAI211_X1 U6927 ( .C1(n8629), .C2(n5436), .A(n5435), .B(n5434), .ZN(n5437)
         );
  INV_X1 U6928 ( .A(n5437), .ZN(n5438) );
  NAND2_X1 U6929 ( .A1(n5439), .A2(n5438), .ZN(n9167) );
  NAND2_X1 U6930 ( .A1(n9167), .A2(n5617), .ZN(n5440) );
  NAND2_X1 U6931 ( .A1(n5441), .A2(n5440), .ZN(n5442) );
  XNOR2_X1 U6932 ( .A(n5442), .B(n5620), .ZN(n5446) );
  NAND2_X1 U6933 ( .A1(n9297), .A2(n5617), .ZN(n5444) );
  NAND2_X1 U6934 ( .A1(n9167), .A2(n5622), .ZN(n5443) );
  NAND2_X1 U6935 ( .A1(n5444), .A2(n5443), .ZN(n5445) );
  NAND2_X1 U6936 ( .A1(n5446), .A2(n5445), .ZN(n8565) );
  NOR2_X1 U6937 ( .A1(n5446), .A2(n5445), .ZN(n8564) );
  AOI21_X2 U6938 ( .B1(n8563), .B2(n8565), .A(n8564), .ZN(n8523) );
  XNOR2_X1 U6939 ( .A(n5448), .B(n5447), .ZN(n6902) );
  NAND2_X1 U6940 ( .A1(n6902), .A2(n5229), .ZN(n5450) );
  OR2_X1 U6941 ( .A1(n8635), .A2(n6903), .ZN(n5449) );
  NAND2_X1 U6942 ( .A1(n5452), .A2(n5451), .ZN(n5453) );
  AND2_X1 U6943 ( .A1(n5471), .A2(n5453), .ZN(n8524) );
  NAND2_X1 U6944 ( .A1(n8524), .A2(n5578), .ZN(n5459) );
  INV_X1 U6945 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U6946 ( .A1(n6268), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U6947 ( .A1(n8625), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5454) );
  OAI211_X1 U6948 ( .C1(n8629), .C2(n5456), .A(n5455), .B(n5454), .ZN(n5457)
         );
  INV_X1 U6949 ( .A(n5457), .ZN(n5458) );
  NOR2_X1 U6950 ( .A1(n8963), .A2(n5590), .ZN(n5460) );
  AOI21_X1 U6951 ( .B1(n9294), .B2(n5617), .A(n5460), .ZN(n5463) );
  INV_X1 U6952 ( .A(n9294), .ZN(n8964) );
  OAI22_X1 U6953 ( .A1(n8964), .A2(n5480), .B1(n8963), .B2(n5461), .ZN(n5462)
         );
  XNOR2_X1 U6954 ( .A(n5462), .B(n5620), .ZN(n5465) );
  XOR2_X1 U6955 ( .A(n5463), .B(n5465), .Z(n8522) );
  INV_X1 U6956 ( .A(n5463), .ZN(n5464) );
  XNOR2_X1 U6957 ( .A(n5467), .B(n5466), .ZN(n6980) );
  NAND2_X1 U6958 ( .A1(n6980), .A2(n5229), .ZN(n5469) );
  OR2_X1 U6959 ( .A1(n8635), .A2(n6981), .ZN(n5468) );
  INV_X1 U6960 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U6961 ( .A1(n5471), .A2(n5470), .ZN(n5472) );
  NAND2_X1 U6962 ( .A1(n5473), .A2(n5472), .ZN(n9120) );
  INV_X1 U6963 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U6964 ( .A1(n8625), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U6965 ( .A1(n6268), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5474) );
  OAI211_X1 U6966 ( .C1(n8629), .C2(n5476), .A(n5475), .B(n5474), .ZN(n5477)
         );
  INV_X1 U6967 ( .A(n5477), .ZN(n5478) );
  AOI22_X1 U6968 ( .A1(n9287), .A2(n5617), .B1(n5622), .B2(n9106), .ZN(n5486)
         );
  NAND2_X1 U6969 ( .A1(n5485), .A2(n5486), .ZN(n8575) );
  OAI22_X1 U6970 ( .A1(n9123), .A2(n5480), .B1(n9135), .B2(n5161), .ZN(n5481)
         );
  XNOR2_X1 U6971 ( .A(n5481), .B(n5620), .ZN(n8577) );
  NAND2_X1 U6972 ( .A1(n9282), .A2(n5605), .ZN(n5483) );
  NAND2_X1 U6973 ( .A1(n9126), .A2(n5617), .ZN(n5482) );
  NAND2_X1 U6974 ( .A1(n5483), .A2(n5482), .ZN(n5484) );
  XNOR2_X1 U6975 ( .A(n5484), .B(n5588), .ZN(n5489) );
  INV_X1 U6976 ( .A(n5485), .ZN(n5488) );
  INV_X1 U6977 ( .A(n5486), .ZN(n5487) );
  NAND2_X1 U6978 ( .A1(n5488), .A2(n5487), .ZN(n8574) );
  NAND2_X1 U6979 ( .A1(n5492), .A2(n5491), .ZN(n5494) );
  INV_X1 U6980 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n5495) );
  INV_X1 U6981 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7135) );
  MUX2_X1 U6982 ( .A(n5495), .B(n7135), .S(n7548), .Z(n5519) );
  XNOR2_X1 U6983 ( .A(n5519), .B(SI_24_), .ZN(n5516) );
  XNOR2_X1 U6984 ( .A(n5518), .B(n5516), .ZN(n7132) );
  NAND2_X1 U6985 ( .A1(n7132), .A2(n5229), .ZN(n5497) );
  OR2_X1 U6986 ( .A1(n8635), .A2(n7135), .ZN(n5496) );
  NAND2_X1 U6987 ( .A1(n9278), .A2(n4299), .ZN(n5508) );
  INV_X1 U6988 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U6989 ( .A1(n5499), .A2(n5498), .ZN(n5500) );
  AND2_X1 U6990 ( .A1(n5530), .A2(n5500), .ZN(n9088) );
  NAND2_X1 U6991 ( .A1(n9088), .A2(n5578), .ZN(n5506) );
  INV_X1 U6992 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U6993 ( .A1(n8625), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U6994 ( .A1(n6268), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5501) );
  OAI211_X1 U6995 ( .C1(n8629), .C2(n5503), .A(n5502), .B(n5501), .ZN(n5504)
         );
  INV_X1 U6996 ( .A(n5504), .ZN(n5505) );
  NAND2_X1 U6997 ( .A1(n9113), .A2(n5617), .ZN(n5507) );
  NAND2_X1 U6998 ( .A1(n5508), .A2(n5507), .ZN(n5509) );
  XNOR2_X1 U6999 ( .A(n5509), .B(n5620), .ZN(n5513) );
  NAND2_X1 U7000 ( .A1(n9278), .A2(n5617), .ZN(n5511) );
  NAND2_X1 U7001 ( .A1(n9113), .A2(n5622), .ZN(n5510) );
  NAND2_X1 U7002 ( .A1(n5511), .A2(n5510), .ZN(n5512) );
  NOR2_X1 U7003 ( .A1(n5513), .A2(n5512), .ZN(n5514) );
  AOI21_X1 U7004 ( .B1(n5513), .B2(n5512), .A(n5514), .ZN(n8556) );
  INV_X1 U7005 ( .A(n5514), .ZN(n5515) );
  NAND2_X1 U7006 ( .A1(n8555), .A2(n5515), .ZN(n8530) );
  INV_X1 U7007 ( .A(n5516), .ZN(n5517) );
  INV_X1 U7008 ( .A(n5519), .ZN(n5520) );
  NAND2_X1 U7009 ( .A1(n5520), .A2(SI_24_), .ZN(n5521) );
  MUX2_X1 U7010 ( .A(n9922), .B(n7426), .S(n7554), .Z(n5523) );
  INV_X1 U7011 ( .A(SI_25_), .ZN(n5522) );
  NAND2_X1 U7012 ( .A1(n5523), .A2(n5522), .ZN(n5541) );
  INV_X1 U7013 ( .A(n5523), .ZN(n5524) );
  NAND2_X1 U7014 ( .A1(n5524), .A2(SI_25_), .ZN(n5525) );
  NAND2_X1 U7015 ( .A1(n5541), .A2(n5525), .ZN(n5542) );
  XNOR2_X1 U7016 ( .A(n5543), .B(n5542), .ZN(n7421) );
  NAND2_X1 U7017 ( .A1(n7421), .A2(n5229), .ZN(n5527) );
  OR2_X1 U7018 ( .A1(n8635), .A2(n7426), .ZN(n5526) );
  INV_X1 U7019 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U7020 ( .A1(n5530), .A2(n5529), .ZN(n5531) );
  NAND2_X1 U7021 ( .A1(n5551), .A2(n5531), .ZN(n9073) );
  INV_X1 U7022 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U7023 ( .A1(n8625), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U7024 ( .A1(n6268), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5532) );
  OAI211_X1 U7025 ( .C1(n5534), .C2(n8629), .A(n5533), .B(n5532), .ZN(n5535)
         );
  INV_X1 U7026 ( .A(n5535), .ZN(n5536) );
  OAI22_X1 U7027 ( .A1(n9076), .A2(n5461), .B1(n8971), .B2(n5590), .ZN(n5564)
         );
  NAND2_X1 U7028 ( .A1(n9272), .A2(n5605), .ZN(n5539) );
  NAND2_X1 U7029 ( .A1(n8972), .A2(n5617), .ZN(n5538) );
  NAND2_X1 U7030 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  XNOR2_X1 U7031 ( .A(n5540), .B(n5620), .ZN(n5563) );
  XOR2_X1 U7032 ( .A(n5564), .B(n5563), .Z(n8531) );
  INV_X1 U7033 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5544) );
  INV_X1 U7034 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7427) );
  MUX2_X1 U7035 ( .A(n5544), .B(n7427), .S(n7554), .Z(n5546) );
  INV_X1 U7036 ( .A(SI_26_), .ZN(n5545) );
  NAND2_X1 U7037 ( .A1(n5546), .A2(n5545), .ZN(n5570) );
  INV_X1 U7038 ( .A(n5546), .ZN(n5547) );
  NAND2_X1 U7039 ( .A1(n5547), .A2(SI_26_), .ZN(n5548) );
  NAND2_X1 U7040 ( .A1(n7398), .A2(n5229), .ZN(n5550) );
  OR2_X1 U7041 ( .A1(n8635), .A2(n7427), .ZN(n5549) );
  NAND2_X1 U7042 ( .A1(n9267), .A2(n4299), .ZN(n5560) );
  INV_X1 U7043 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U7044 ( .A1(n5551), .A2(n8598), .ZN(n5552) );
  NAND2_X1 U7045 ( .A1(n9059), .A2(n5578), .ZN(n5558) );
  INV_X1 U7046 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U7047 ( .A1(n8625), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U7048 ( .A1(n6268), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5553) );
  OAI211_X1 U7049 ( .C1(n8629), .C2(n5555), .A(n5554), .B(n5553), .ZN(n5556)
         );
  INV_X1 U7050 ( .A(n5556), .ZN(n5557) );
  NAND2_X1 U7051 ( .A1(n9080), .A2(n5617), .ZN(n5559) );
  NAND2_X1 U7052 ( .A1(n5560), .A2(n5559), .ZN(n5561) );
  XNOR2_X1 U7053 ( .A(n5561), .B(n5620), .ZN(n5598) );
  AND2_X1 U7054 ( .A1(n9080), .A2(n5622), .ZN(n5562) );
  AOI21_X1 U7055 ( .B1(n9267), .B2(n5617), .A(n5562), .ZN(n5596) );
  XNOR2_X1 U7056 ( .A(n5598), .B(n5596), .ZN(n8596) );
  INV_X1 U7057 ( .A(n5563), .ZN(n5566) );
  INV_X1 U7058 ( .A(n5564), .ZN(n5565) );
  NAND2_X1 U7059 ( .A1(n5566), .A2(n5565), .ZN(n8592) );
  NAND2_X1 U7060 ( .A1(n5571), .A2(n5570), .ZN(n5600) );
  INV_X1 U7061 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7511) );
  INV_X1 U7062 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5575) );
  MUX2_X1 U7063 ( .A(n7511), .B(n5575), .S(n7554), .Z(n5572) );
  INV_X1 U7064 ( .A(SI_27_), .ZN(n9964) );
  NAND2_X1 U7065 ( .A1(n5572), .A2(n9964), .ZN(n5601) );
  INV_X1 U7066 ( .A(n5572), .ZN(n5573) );
  NAND2_X1 U7067 ( .A1(n5573), .A2(SI_27_), .ZN(n5574) );
  NAND2_X1 U7068 ( .A1(n7494), .A2(n5229), .ZN(n5577) );
  OR2_X1 U7069 ( .A1(n8635), .A2(n5575), .ZN(n5576) );
  NAND2_X1 U7070 ( .A1(n9262), .A2(n5605), .ZN(n5587) );
  XNOR2_X1 U7071 ( .A(n5607), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9042) );
  NAND2_X1 U7072 ( .A1(n9042), .A2(n5578), .ZN(n5585) );
  INV_X1 U7073 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U7074 ( .A1(n6267), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U7075 ( .A1(n8625), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5579) );
  OAI211_X1 U7076 ( .C1(n5582), .C2(n5581), .A(n5580), .B(n5579), .ZN(n5583)
         );
  INV_X1 U7077 ( .A(n5583), .ZN(n5584) );
  INV_X1 U7078 ( .A(n9024), .ZN(n9066) );
  NAND2_X1 U7079 ( .A1(n9066), .A2(n5617), .ZN(n5586) );
  NAND2_X1 U7080 ( .A1(n5587), .A2(n5586), .ZN(n5589) );
  XNOR2_X1 U7081 ( .A(n5589), .B(n5588), .ZN(n5593) );
  INV_X1 U7082 ( .A(n5593), .ZN(n5595) );
  NOR2_X1 U7083 ( .A1(n9024), .A2(n5590), .ZN(n5591) );
  AOI21_X1 U7084 ( .B1(n9262), .B2(n5617), .A(n5591), .ZN(n5592) );
  INV_X1 U7085 ( .A(n5592), .ZN(n5594) );
  AOI21_X1 U7086 ( .B1(n5595), .B2(n5594), .A(n5650), .ZN(n8496) );
  INV_X1 U7087 ( .A(n5596), .ZN(n5597) );
  NAND2_X1 U7088 ( .A1(n5598), .A2(n5597), .ZN(n8497) );
  NAND2_X1 U7089 ( .A1(n5600), .A2(n5599), .ZN(n5602) );
  MUX2_X1 U7090 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7548), .Z(n7542) );
  INV_X1 U7091 ( .A(SI_28_), .ZN(n7543) );
  XNOR2_X1 U7092 ( .A(n7542), .B(n7543), .ZN(n7540) );
  NAND2_X1 U7093 ( .A1(n7512), .A2(n5229), .ZN(n5604) );
  INV_X1 U7094 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10040) );
  OR2_X1 U7095 ( .A1(n8635), .A2(n10040), .ZN(n5603) );
  NAND2_X1 U7096 ( .A1(n9256), .A2(n4299), .ZN(n5619) );
  INV_X1 U7097 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8500) );
  INV_X1 U7098 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5606) );
  OAI21_X1 U7099 ( .B1(n5607), .B2(n8500), .A(n5606), .ZN(n5610) );
  INV_X1 U7100 ( .A(n5607), .ZN(n5609) );
  AND2_X1 U7101 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5608) );
  NAND2_X1 U7102 ( .A1(n5609), .A2(n5608), .ZN(n9013) );
  NAND2_X1 U7103 ( .A1(n5610), .A2(n9013), .ZN(n5666) );
  INV_X1 U7104 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7105 ( .A1(n8625), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U7106 ( .A1(n6268), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5611) );
  OAI211_X1 U7107 ( .C1(n8629), .C2(n5613), .A(n5612), .B(n5611), .ZN(n5614)
         );
  INV_X1 U7108 ( .A(n5614), .ZN(n5615) );
  NAND2_X1 U7109 ( .A1(n9009), .A2(n5617), .ZN(n5618) );
  NAND2_X1 U7110 ( .A1(n5619), .A2(n5618), .ZN(n5621) );
  XNOR2_X1 U7111 ( .A(n5621), .B(n5620), .ZN(n5624) );
  AOI22_X1 U7112 ( .A1(n9256), .A2(n5617), .B1(n5622), .B2(n9009), .ZN(n5623)
         );
  XNOR2_X1 U7113 ( .A(n5624), .B(n5623), .ZN(n5651) );
  INV_X1 U7114 ( .A(n5625), .ZN(n7424) );
  NAND2_X1 U7115 ( .A1(n7424), .A2(P1_B_REG_SCAN_IN), .ZN(n5626) );
  MUX2_X1 U7116 ( .A(n5626), .B(P1_B_REG_SCAN_IN), .S(n5642), .Z(n5628) );
  NAND2_X1 U7117 ( .A1(n5628), .A2(n5627), .ZN(n9656) );
  INV_X1 U7118 ( .A(n9656), .ZN(n5641) );
  NOR4_X1 U7119 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5637) );
  NOR4_X1 U7120 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5636) );
  INV_X1 U7121 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9996) );
  INV_X1 U7122 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9658) );
  INV_X1 U7123 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9924) );
  INV_X1 U7124 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9960) );
  NAND4_X1 U7125 ( .A1(n9996), .A2(n9658), .A3(n9924), .A4(n9960), .ZN(n5634)
         );
  NOR4_X1 U7126 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5632) );
  NOR4_X1 U7127 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n5631) );
  NOR4_X1 U7128 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5630) );
  NOR4_X1 U7129 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5629) );
  NAND4_X1 U7130 ( .A1(n5632), .A2(n5631), .A3(n5630), .A4(n5629), .ZN(n5633)
         );
  NOR4_X1 U7131 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5634), .A4(n5633), .ZN(n5635) );
  NAND3_X1 U7132 ( .A1(n5637), .A2(n5636), .A3(n5635), .ZN(n5638) );
  NAND2_X1 U7133 ( .A1(n5641), .A2(n5638), .ZN(n6329) );
  INV_X1 U7134 ( .A(n6329), .ZN(n5639) );
  OAI22_X1 U7135 ( .A1(n9656), .A2(P1_D_REG_1__SCAN_IN), .B1(n5627), .B2(n5625), .ZN(n6330) );
  NOR2_X1 U7136 ( .A1(n5639), .A2(n6330), .ZN(n6355) );
  INV_X1 U7137 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5640) );
  NAND2_X1 U7138 ( .A1(n5641), .A2(n5640), .ZN(n5644) );
  INV_X1 U7139 ( .A(n5627), .ZN(n7428) );
  INV_X1 U7140 ( .A(n5642), .ZN(n7136) );
  NAND2_X1 U7141 ( .A1(n7428), .A2(n7136), .ZN(n5643) );
  NAND2_X1 U7142 ( .A1(n4371), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5646) );
  XNOR2_X1 U7143 ( .A(n5646), .B(n5645), .ZN(n6241) );
  NAND2_X1 U7144 ( .A1(n6837), .A2(n9646), .ZN(n5668) );
  NAND2_X1 U7145 ( .A1(n5028), .A2(n5668), .ZN(n9479) );
  INV_X2 U7146 ( .A(n9479), .ZN(n9330) );
  OR2_X1 U7147 ( .A1(n9330), .A2(n6445), .ZN(n5667) );
  NOR2_X1 U7148 ( .A1(n6320), .A2(n5667), .ZN(n5649) );
  NAND3_X1 U7149 ( .A1(n5651), .A2(n5650), .A3(n8595), .ZN(n5682) );
  NOR2_X1 U7150 ( .A1(n6336), .A2(n6837), .ZN(n9640) );
  INV_X1 U7151 ( .A(n9640), .ZN(n5652) );
  OR2_X1 U7152 ( .A1(n6320), .A2(n5652), .ZN(n5653) );
  OR2_X1 U7153 ( .A1(n5676), .A2(n5653), .ZN(n5655) );
  OR2_X1 U7154 ( .A1(n8741), .A2(n4798), .ZN(n9663) );
  INV_X1 U7155 ( .A(n6445), .ZN(n8776) );
  OR2_X1 U7156 ( .A1(n8776), .A2(n5668), .ZN(n6441) );
  NOR2_X1 U7157 ( .A1(n6320), .A2(n6441), .ZN(n8873) );
  INV_X1 U7158 ( .A(n8873), .ZN(n5656) );
  OR2_X1 U7159 ( .A1(n5676), .A2(n5656), .ZN(n5665) );
  NOR2_X1 U7160 ( .A1(n9024), .A2(n8599), .ZN(n5680) );
  OR2_X1 U7161 ( .A1(n9013), .A2(n5658), .ZN(n5664) );
  INV_X1 U7162 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7163 ( .A1(n8625), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U7164 ( .A1(n6268), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5659) );
  OAI211_X1 U7165 ( .C1(n8629), .C2(n5661), .A(n5660), .B(n5659), .ZN(n5662)
         );
  INV_X1 U7166 ( .A(n5662), .ZN(n5663) );
  INV_X1 U7167 ( .A(n5666), .ZN(n9034) );
  INV_X1 U7168 ( .A(n5667), .ZN(n5671) );
  AND2_X1 U7169 ( .A1(n6445), .A2(n5668), .ZN(n6319) );
  INV_X1 U7170 ( .A(n6319), .ZN(n5669) );
  NAND3_X1 U7171 ( .A1(n5669), .A2(n5057), .A3(n6241), .ZN(n5670) );
  AOI21_X1 U7172 ( .B1(n5676), .B2(n5671), .A(n5670), .ZN(n5672) );
  OR2_X1 U7173 ( .A1(n5672), .A2(P1_U3084), .ZN(n5677) );
  INV_X1 U7174 ( .A(n6441), .ZN(n5673) );
  NOR2_X1 U7175 ( .A1(n9640), .A2(n5673), .ZN(n5674) );
  NOR2_X1 U7176 ( .A1(n5674), .A2(n6320), .ZN(n5675) );
  NAND2_X1 U7177 ( .A1(n5676), .A2(n5675), .ZN(n6321) );
  AOI22_X1 U7178 ( .A1(n9034), .A2(n8612), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n5678) );
  OAI21_X1 U7179 ( .B1(n9023), .B2(n8615), .A(n5678), .ZN(n5679) );
  AOI211_X1 U7180 ( .C1(n9256), .C2(n8617), .A(n5680), .B(n5679), .ZN(n5681)
         );
  NAND2_X1 U7181 ( .A1(n5682), .A2(n5681), .ZN(n5683) );
  NOR2_X1 U7182 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5691) );
  NOR2_X1 U7183 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5690) );
  NOR2_X1 U7184 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5689) );
  NOR2_X1 U7185 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5688) );
  NAND4_X1 U7186 ( .A1(n5691), .A2(n5690), .A3(n5689), .A4(n5688), .ZN(n5697)
         );
  NOR2_X1 U7187 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5695) );
  NAND4_X1 U7188 ( .A1(n5695), .A2(n5694), .A3(n5693), .A4(n5692), .ZN(n5696)
         );
  OR2_X1 U7189 ( .A1(n5706), .A2(n5976), .ZN(n5700) );
  INV_X1 U7190 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5701) );
  AND2_X2 U7191 ( .A1(n5706), .A2(n5701), .ZN(n5734) );
  INV_X1 U7192 ( .A(n5734), .ZN(n5702) );
  NAND2_X1 U7193 ( .A1(n5704), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5705) );
  INV_X1 U7194 ( .A(n5706), .ZN(n5707) );
  NAND2_X1 U7195 ( .A1(n7072), .A2(n7565), .ZN(n5710) );
  NAND2_X1 U7196 ( .A1(n7566), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5709) );
  NOR2_X1 U7197 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5716) );
  OAI21_X2 U7198 ( .B1(n4301), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6180) );
  INV_X1 U7199 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5717) );
  INV_X1 U7200 ( .A(n7799), .ZN(n5719) );
  INV_X1 U7201 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U7202 ( .A1(n6212), .A2(n8219), .ZN(n7833) );
  NAND2_X1 U7203 ( .A1(n5732), .A2(n7833), .ZN(n7990) );
  XNOR2_X1 U7204 ( .A(n8427), .B(n5763), .ZN(n6115) );
  NAND2_X1 U7205 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5726) );
  MUX2_X1 U7206 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5726), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5729) );
  INV_X1 U7207 ( .A(n5727), .ZN(n5728) );
  INV_X1 U7208 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6244) );
  OR2_X1 U7209 ( .A1(n5793), .A2(n6244), .ZN(n5731) );
  OR2_X1 U7210 ( .A1(n5792), .A2(n6246), .ZN(n5730) );
  INV_X1 U7211 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U7212 ( .A1(n5734), .A2(n5733), .ZN(n5737) );
  AND2_X2 U7213 ( .A1(n5740), .A2(n8492), .ZN(n5812) );
  NAND2_X1 U7214 ( .A1(n5812), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5745) );
  NAND2_X1 U7215 ( .A1(n5741), .A2(n5740), .ZN(n5751) );
  NAND2_X1 U7216 ( .A1(n5779), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U7217 ( .A1(n5835), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5742) );
  NAND2_X1 U7218 ( .A1(n7809), .A2(n7184), .ZN(n5759) );
  XNOR2_X1 U7219 ( .A(n5758), .B(n5759), .ZN(n7675) );
  NAND2_X1 U7220 ( .A1(n5746), .A2(SI_0_), .ZN(n5748) );
  INV_X1 U7221 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5747) );
  NAND2_X1 U7222 ( .A1(n5748), .A2(n5747), .ZN(n5750) );
  AND2_X1 U7223 ( .A1(n5750), .A2(n5749), .ZN(n8495) );
  MUX2_X1 U7224 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8495), .S(n6700), .Z(n7586) );
  OR2_X1 U7225 ( .A1(n5763), .A2(n7586), .ZN(n5757) );
  NAND2_X1 U7226 ( .A1(n5812), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5755) );
  NAND2_X1 U7227 ( .A1(n5811), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U7228 ( .A1(n5779), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U7229 ( .A1(n5835), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5752) );
  INV_X1 U7230 ( .A(n7586), .ZN(n9717) );
  OR2_X1 U7231 ( .A1(n7581), .A2(n9717), .ZN(n7376) );
  INV_X1 U7232 ( .A(n7376), .ZN(n5756) );
  NAND2_X1 U7233 ( .A1(n7809), .A2(n5756), .ZN(n7582) );
  AND2_X1 U7234 ( .A1(n5757), .A2(n7582), .ZN(n7676) );
  NAND2_X1 U7235 ( .A1(n7675), .A2(n7676), .ZN(n7674) );
  INV_X1 U7236 ( .A(n5758), .ZN(n5760) );
  NAND2_X1 U7237 ( .A1(n5760), .A2(n5759), .ZN(n5761) );
  INV_X1 U7238 ( .A(n7753), .ZN(n5773) );
  OR2_X1 U7239 ( .A1(n5727), .A2(n5976), .ZN(n5762) );
  XNOR2_X1 U7240 ( .A(n5762), .B(n4733), .ZN(n6741) );
  XNOR2_X1 U7241 ( .A(n5763), .B(n7751), .ZN(n5768) );
  NAND2_X1 U7242 ( .A1(n5812), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5767) );
  NAND2_X1 U7243 ( .A1(n5811), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5766) );
  NAND2_X1 U7244 ( .A1(n5779), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U7245 ( .A1(n5835), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5764) );
  AND2_X1 U7246 ( .A1(n7809), .A2(n8025), .ZN(n5769) );
  NAND2_X1 U7247 ( .A1(n5768), .A2(n5769), .ZN(n5774) );
  INV_X1 U7248 ( .A(n5768), .ZN(n7077) );
  INV_X1 U7249 ( .A(n5769), .ZN(n5770) );
  NAND2_X1 U7250 ( .A1(n7077), .A2(n5770), .ZN(n5771) );
  NAND2_X1 U7251 ( .A1(n5774), .A2(n5771), .ZN(n7752) );
  NAND2_X1 U7252 ( .A1(n7754), .A2(n5774), .ZN(n5789) );
  OR3_X1 U7253 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n5775) );
  NAND2_X1 U7254 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5775), .ZN(n5776) );
  XNOR2_X1 U7255 ( .A(n5776), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6735) );
  INV_X1 U7256 ( .A(n6735), .ZN(n8032) );
  OR2_X1 U7257 ( .A1(n5792), .A2(n6261), .ZN(n5778) );
  OR2_X1 U7258 ( .A1(n5793), .A2(n6262), .ZN(n5777) );
  OAI211_X1 U7259 ( .C1(n6700), .C2(n8032), .A(n5778), .B(n5777), .ZN(n8367)
         );
  XNOR2_X1 U7260 ( .A(n5763), .B(n8367), .ZN(n7158) );
  NAND2_X1 U7261 ( .A1(n5812), .A2(n8368), .ZN(n5784) );
  NAND2_X1 U7262 ( .A1(n5811), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5783) );
  INV_X1 U7263 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U7264 ( .A1(n5835), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5781) );
  AND2_X1 U7265 ( .A1(n7809), .A2(n8024), .ZN(n5785) );
  NAND2_X1 U7266 ( .A1(n7158), .A2(n5785), .ZN(n5800) );
  INV_X1 U7267 ( .A(n7158), .ZN(n5787) );
  INV_X1 U7268 ( .A(n5785), .ZN(n5786) );
  NAND2_X1 U7269 ( .A1(n5787), .A2(n5786), .ZN(n5788) );
  AND2_X1 U7270 ( .A1(n5800), .A2(n5788), .ZN(n7078) );
  NAND2_X1 U7271 ( .A1(n5790), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5791) );
  XNOR2_X1 U7272 ( .A(n5791), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6734) );
  INV_X1 U7273 ( .A(n6734), .ZN(n8046) );
  OR2_X1 U7274 ( .A1(n5792), .A2(n6257), .ZN(n5795) );
  OR2_X1 U7275 ( .A1(n5793), .A2(n6258), .ZN(n5794) );
  OAI211_X1 U7276 ( .C1(n6700), .C2(n8046), .A(n5795), .B(n5794), .ZN(n7211)
         );
  XNOR2_X1 U7277 ( .A(n5763), .B(n7211), .ZN(n5802) );
  NAND2_X1 U7278 ( .A1(n7604), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5799) );
  INV_X1 U7279 ( .A(n5813), .ZN(n5814) );
  OAI21_X1 U7280 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5814), .ZN(n7162) );
  INV_X1 U7281 ( .A(n7162), .ZN(n7416) );
  NAND2_X1 U7282 ( .A1(n5812), .A2(n7416), .ZN(n5798) );
  NAND2_X1 U7283 ( .A1(n5811), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5797) );
  NAND2_X1 U7284 ( .A1(n5835), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5796) );
  NAND3_X1 U7285 ( .A1(n5799), .A2(n5798), .A3(n4835), .ZN(n8023) );
  NAND2_X1 U7286 ( .A1(n7809), .A2(n8023), .ZN(n5803) );
  XNOR2_X1 U7287 ( .A(n5802), .B(n5803), .ZN(n7157) );
  AND2_X1 U7288 ( .A1(n7157), .A2(n5800), .ZN(n5801) );
  INV_X1 U7289 ( .A(n5802), .ZN(n5804) );
  NAND2_X1 U7290 ( .A1(n5804), .A2(n5803), .ZN(n5805) );
  OR2_X1 U7291 ( .A1(n5792), .A2(n6259), .ZN(n5810) );
  OR2_X1 U7292 ( .A1(n5793), .A2(n6260), .ZN(n5809) );
  OR2_X1 U7293 ( .A1(n5806), .A2(n5976), .ZN(n5807) );
  XNOR2_X1 U7294 ( .A(n5807), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6732) );
  NAND2_X1 U7295 ( .A1(n6514), .A2(n6732), .ZN(n5808) );
  XNOR2_X1 U7296 ( .A(n5763), .B(n7458), .ZN(n5820) );
  INV_X2 U7297 ( .A(n5751), .ZN(n7603) );
  NAND2_X1 U7298 ( .A1(n5813), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5832) );
  INV_X1 U7299 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8058) );
  NAND2_X1 U7300 ( .A1(n5814), .A2(n8058), .ZN(n5815) );
  AND2_X1 U7301 ( .A1(n5832), .A2(n5815), .ZN(n7459) );
  NAND2_X1 U7302 ( .A1(n5812), .A2(n7459), .ZN(n5818) );
  NAND2_X1 U7303 ( .A1(n7604), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5817) );
  NAND2_X1 U7304 ( .A1(n4298), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5816) );
  AND2_X1 U7305 ( .A1(n7809), .A2(n8022), .ZN(n5821) );
  NAND2_X1 U7306 ( .A1(n5820), .A2(n5821), .ZN(n5840) );
  INV_X1 U7307 ( .A(n5820), .ZN(n7100) );
  INV_X1 U7308 ( .A(n5821), .ZN(n5822) );
  NAND2_X1 U7309 ( .A1(n7100), .A2(n5822), .ZN(n5823) );
  NAND2_X1 U7310 ( .A1(n5840), .A2(n5823), .ZN(n6940) );
  NAND2_X1 U7311 ( .A1(n5825), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5827) );
  INV_X1 U7312 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U7313 ( .A1(n5827), .A2(n5826), .ZN(n5846) );
  OR2_X1 U7314 ( .A1(n5827), .A2(n5826), .ZN(n5828) );
  INV_X1 U7315 ( .A(n6729), .ZN(n6802) );
  OR2_X1 U7316 ( .A1(n5792), .A2(n6255), .ZN(n5830) );
  OR2_X1 U7317 ( .A1(n5793), .A2(n6256), .ZN(n5829) );
  OAI211_X1 U7318 ( .C1(n6700), .C2(n6802), .A(n5830), .B(n5829), .ZN(n7215)
         );
  XNOR2_X1 U7319 ( .A(n5763), .B(n7215), .ZN(n5842) );
  NAND2_X1 U7320 ( .A1(n7603), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5839) );
  NOR2_X1 U7321 ( .A1(n5832), .A2(n5831), .ZN(n5850) );
  INV_X1 U7322 ( .A(n5850), .ZN(n5851) );
  NAND2_X1 U7323 ( .A1(n5832), .A2(n5831), .ZN(n5833) );
  AND2_X1 U7324 ( .A1(n5851), .A2(n5833), .ZN(n7212) );
  NAND2_X1 U7325 ( .A1(n6224), .A2(n7212), .ZN(n5838) );
  INV_X4 U7326 ( .A(n5834), .ZN(n7604) );
  NAND2_X1 U7327 ( .A1(n7604), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U7328 ( .A1(n4298), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5836) );
  INV_X1 U7329 ( .A(n7453), .ZN(n8021) );
  NAND2_X1 U7330 ( .A1(n7809), .A2(n8021), .ZN(n5843) );
  XNOR2_X1 U7331 ( .A(n5842), .B(n5843), .ZN(n7110) );
  AND2_X1 U7332 ( .A1(n7110), .A2(n5840), .ZN(n5841) );
  NAND2_X1 U7333 ( .A1(n6938), .A2(n5841), .ZN(n7103) );
  INV_X1 U7334 ( .A(n5842), .ZN(n5844) );
  NAND2_X1 U7335 ( .A1(n5844), .A2(n5843), .ZN(n5845) );
  NAND2_X1 U7336 ( .A1(n5846), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5847) );
  XNOR2_X1 U7337 ( .A(n5847), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6727) );
  AOI22_X1 U7338 ( .A1(n7566), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6514), .B2(
        n6727), .ZN(n5849) );
  NAND2_X1 U7339 ( .A1(n6265), .A2(n7565), .ZN(n5848) );
  XNOR2_X1 U7340 ( .A(n5763), .B(n7874), .ZN(n9677) );
  NAND2_X1 U7341 ( .A1(n7603), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5856) );
  NAND2_X1 U7342 ( .A1(n5850), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5885) );
  INV_X1 U7343 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6759) );
  NAND2_X1 U7344 ( .A1(n5851), .A2(n6759), .ZN(n5852) );
  AND2_X1 U7345 ( .A1(n5885), .A2(n5852), .ZN(n7244) );
  NAND2_X1 U7346 ( .A1(n6224), .A2(n7244), .ZN(n5855) );
  NAND2_X1 U7347 ( .A1(n7604), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U7348 ( .A1(n4298), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5853) );
  AND2_X1 U7349 ( .A1(n7809), .A2(n9683), .ZN(n5857) );
  NAND2_X1 U7350 ( .A1(n9677), .A2(n5857), .ZN(n5870) );
  INV_X1 U7351 ( .A(n9677), .ZN(n5859) );
  INV_X1 U7352 ( .A(n5857), .ZN(n5858) );
  NAND2_X1 U7353 ( .A1(n5859), .A2(n5858), .ZN(n5860) );
  NAND2_X1 U7354 ( .A1(n5870), .A2(n5860), .ZN(n7065) );
  NAND2_X1 U7355 ( .A1(n6276), .A2(n7565), .ZN(n5864) );
  NAND2_X1 U7356 ( .A1(n5861), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5862) );
  XNOR2_X1 U7357 ( .A(n5862), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6724) );
  AOI22_X1 U7358 ( .A1(n7566), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6514), .B2(
        n6724), .ZN(n5863) );
  NAND2_X1 U7359 ( .A1(n5864), .A2(n5863), .ZN(n7238) );
  XNOR2_X1 U7360 ( .A(n5763), .B(n7238), .ZN(n5875) );
  INV_X1 U7361 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5883) );
  XNOR2_X1 U7362 ( .A(n5885), .B(n5883), .ZN(n9692) );
  INV_X1 U7363 ( .A(n9692), .ZN(n5865) );
  NAND2_X1 U7364 ( .A1(n6224), .A2(n5865), .ZN(n5869) );
  NAND2_X1 U7365 ( .A1(n7603), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7366 ( .A1(n7604), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U7367 ( .A1(n4298), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U7368 ( .A1(n7809), .A2(n8020), .ZN(n5873) );
  XNOR2_X1 U7369 ( .A(n5875), .B(n5873), .ZN(n9675) );
  INV_X1 U7370 ( .A(n9675), .ZN(n5871) );
  OR2_X1 U7371 ( .A1(n5871), .A2(n5870), .ZN(n5872) );
  INV_X1 U7372 ( .A(n5873), .ZN(n5874) );
  NAND2_X1 U7373 ( .A1(n6280), .A2(n7565), .ZN(n5881) );
  OR2_X1 U7374 ( .A1(n5876), .A2(n5976), .ZN(n5878) );
  MUX2_X1 U7375 ( .A(n5878), .B(P2_IR_REG_31__SCAN_IN), .S(n5877), .Z(n5879)
         );
  AND2_X1 U7376 ( .A1(n5879), .A2(n5896), .ZN(n6721) );
  AOI22_X1 U7377 ( .A1(n7566), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6514), .B2(
        n6721), .ZN(n5880) );
  NAND2_X1 U7378 ( .A1(n5881), .A2(n5880), .ZN(n7268) );
  XNOR2_X1 U7379 ( .A(n5763), .B(n7268), .ZN(n5891) );
  NAND2_X1 U7380 ( .A1(n7603), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5890) );
  INV_X1 U7381 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5882) );
  OAI21_X1 U7382 ( .B1(n5885), .B2(n5883), .A(n5882), .ZN(n5886) );
  NAND2_X1 U7383 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5884) );
  AND2_X1 U7384 ( .A1(n5886), .A2(n5900), .ZN(n7126) );
  NAND2_X1 U7385 ( .A1(n6224), .A2(n7126), .ZN(n5889) );
  NAND2_X1 U7386 ( .A1(n7604), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U7387 ( .A1(n4298), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5887) );
  INV_X1 U7388 ( .A(n7277), .ZN(n9681) );
  AND2_X1 U7389 ( .A1(n7809), .A2(n9681), .ZN(n5892) );
  AND2_X1 U7390 ( .A1(n5891), .A2(n5892), .ZN(n7122) );
  INV_X1 U7391 ( .A(n5891), .ZN(n5894) );
  INV_X1 U7392 ( .A(n5892), .ZN(n5893) );
  NAND2_X1 U7393 ( .A1(n5894), .A2(n5893), .ZN(n7121) );
  NAND2_X1 U7394 ( .A1(n6309), .A2(n7565), .ZN(n5899) );
  NAND2_X1 U7395 ( .A1(n5896), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5897) );
  XNOR2_X1 U7396 ( .A(n5897), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6825) );
  AOI22_X1 U7397 ( .A1(n7566), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6514), .B2(
        n6825), .ZN(n5898) );
  NAND2_X1 U7398 ( .A1(n5899), .A2(n5898), .ZN(n7338) );
  XNOR2_X1 U7399 ( .A(n5763), .B(n9782), .ZN(n5907) );
  NAND2_X1 U7400 ( .A1(n7603), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5905) );
  INV_X1 U7401 ( .A(n5912), .ZN(n5913) );
  NAND2_X1 U7402 ( .A1(n5900), .A2(n6703), .ZN(n5901) );
  AND2_X1 U7403 ( .A1(n5913), .A2(n5901), .ZN(n7281) );
  NAND2_X1 U7404 ( .A1(n5812), .A2(n7281), .ZN(n5904) );
  NAND2_X1 U7405 ( .A1(n7604), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U7406 ( .A1(n4298), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5902) );
  INV_X1 U7407 ( .A(n7467), .ZN(n8019) );
  NAND2_X1 U7408 ( .A1(n7809), .A2(n8019), .ZN(n5906) );
  XNOR2_X1 U7409 ( .A(n5907), .B(n5906), .ZN(n7649) );
  NAND2_X1 U7410 ( .A1(n6313), .A2(n7565), .ZN(n5911) );
  NAND2_X1 U7411 ( .A1(n5908), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5909) );
  XNOR2_X1 U7412 ( .A(n5909), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6878) );
  AOI22_X1 U7413 ( .A1(n7566), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6514), .B2(
        n6878), .ZN(n5910) );
  NAND2_X1 U7414 ( .A1(n5911), .A2(n5910), .ZN(n9789) );
  XNOR2_X1 U7415 ( .A(n9789), .B(n5763), .ZN(n5921) );
  NAND2_X1 U7416 ( .A1(n7603), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5918) );
  INV_X1 U7417 ( .A(n5925), .ZN(n5927) );
  INV_X1 U7418 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7392) );
  NAND2_X1 U7419 ( .A1(n5913), .A2(n7392), .ZN(n5914) );
  AND2_X1 U7420 ( .A1(n5927), .A2(n5914), .ZN(n7472) );
  NAND2_X1 U7421 ( .A1(n6224), .A2(n7472), .ZN(n5917) );
  NAND2_X1 U7422 ( .A1(n7604), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U7423 ( .A1(n4298), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5915) );
  INV_X1 U7424 ( .A(n7488), .ZN(n8018) );
  NAND2_X1 U7425 ( .A1(n7809), .A2(n8018), .ZN(n5919) );
  XNOR2_X1 U7426 ( .A(n5921), .B(n5919), .ZN(n7390) );
  INV_X1 U7427 ( .A(n5919), .ZN(n5920) );
  NAND2_X1 U7428 ( .A1(n6317), .A2(n7565), .ZN(n5924) );
  NAND2_X1 U7429 ( .A1(n4364), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5922) );
  XNOR2_X1 U7430 ( .A(n5922), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6963) );
  AOI22_X1 U7431 ( .A1(n7566), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6514), .B2(
        n6963), .ZN(n5923) );
  XNOR2_X1 U7432 ( .A(n7491), .B(n6124), .ZN(n5933) );
  NAND2_X1 U7433 ( .A1(n7603), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5932) );
  NAND2_X1 U7434 ( .A1(n5925), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5943) );
  INV_X1 U7435 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U7436 ( .A1(n5927), .A2(n5926), .ZN(n5928) );
  AND2_X1 U7437 ( .A1(n5943), .A2(n5928), .ZN(n7484) );
  NAND2_X1 U7438 ( .A1(n6224), .A2(n7484), .ZN(n5931) );
  NAND2_X1 U7439 ( .A1(n7604), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5930) );
  NAND2_X1 U7440 ( .A1(n4298), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5929) );
  INV_X1 U7441 ( .A(n7518), .ZN(n8017) );
  NAND2_X1 U7442 ( .A1(n7809), .A2(n8017), .ZN(n5934) );
  NAND2_X1 U7443 ( .A1(n5933), .A2(n5934), .ZN(n7480) );
  INV_X1 U7444 ( .A(n5933), .ZN(n5936) );
  INV_X1 U7445 ( .A(n5934), .ZN(n5935) );
  NAND2_X1 U7446 ( .A1(n5936), .A2(n5935), .ZN(n7481) );
  NAND2_X1 U7447 ( .A1(n5937), .A2(n7481), .ZN(n7517) );
  NAND2_X1 U7448 ( .A1(n5938), .A2(n7565), .ZN(n5941) );
  OR2_X1 U7449 ( .A1(n5939), .A2(n5976), .ZN(n5956) );
  XNOR2_X1 U7450 ( .A(n5956), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7091) );
  AOI22_X1 U7451 ( .A1(n7566), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6514), .B2(
        n7091), .ZN(n5940) );
  XNOR2_X1 U7452 ( .A(n7430), .B(n5763), .ZN(n5949) );
  NAND2_X1 U7453 ( .A1(n7603), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5948) );
  INV_X1 U7454 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5942) );
  NAND2_X1 U7455 ( .A1(n5943), .A2(n5942), .ZN(n5944) );
  AND2_X1 U7456 ( .A1(n5964), .A2(n5944), .ZN(n7521) );
  NAND2_X1 U7457 ( .A1(n5812), .A2(n7521), .ZN(n5947) );
  NAND2_X1 U7458 ( .A1(n7604), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7459 ( .A1(n4298), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5945) );
  INV_X1 U7460 ( .A(n7487), .ZN(n8016) );
  AND2_X1 U7461 ( .A1(n7809), .A2(n8016), .ZN(n5950) );
  NAND2_X1 U7462 ( .A1(n5949), .A2(n5950), .ZN(n5954) );
  INV_X1 U7463 ( .A(n5949), .ZN(n5952) );
  INV_X1 U7464 ( .A(n5950), .ZN(n5951) );
  NAND2_X1 U7465 ( .A1(n5952), .A2(n5951), .ZN(n5953) );
  AND2_X1 U7466 ( .A1(n5954), .A2(n5953), .ZN(n7516) );
  NAND2_X1 U7467 ( .A1(n6404), .A2(n7565), .ZN(n5962) );
  NAND2_X1 U7468 ( .A1(n5956), .A2(n5955), .ZN(n5957) );
  NAND2_X1 U7469 ( .A1(n5957), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5959) );
  OR2_X1 U7470 ( .A1(n5959), .A2(n5958), .ZN(n5960) );
  NAND2_X1 U7471 ( .A1(n5959), .A2(n5958), .ZN(n5996) );
  AOI22_X1 U7472 ( .A1(n7566), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8073), .B2(
        n6514), .ZN(n5961) );
  XNOR2_X1 U7473 ( .A(n9449), .B(n6124), .ZN(n5972) );
  INV_X1 U7474 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U7475 ( .A1(n5964), .A2(n5963), .ZN(n5965) );
  NAND2_X1 U7476 ( .A1(n5989), .A2(n5965), .ZN(n9438) );
  INV_X1 U7477 ( .A(n9438), .ZN(n5966) );
  NAND2_X1 U7478 ( .A1(n6224), .A2(n5966), .ZN(n5970) );
  NAND2_X1 U7479 ( .A1(n7603), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7480 ( .A1(n7604), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7481 ( .A1(n4298), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5967) );
  INV_X1 U7482 ( .A(n7788), .ZN(n8015) );
  NAND2_X1 U7483 ( .A1(n7809), .A2(n8015), .ZN(n5971) );
  XNOR2_X1 U7484 ( .A(n5972), .B(n5971), .ZN(n9429) );
  NAND2_X1 U7485 ( .A1(n5972), .A2(n5971), .ZN(n5973) );
  NAND2_X1 U7486 ( .A1(n6508), .A2(n7565), .ZN(n5980) );
  NOR2_X1 U7487 ( .A1(n5974), .A2(n5976), .ZN(n5975) );
  MUX2_X1 U7488 ( .A(n5976), .B(n5975), .S(P2_IR_REG_16__SCAN_IN), .Z(n5977)
         );
  INV_X1 U7489 ( .A(n5977), .ZN(n5978) );
  AND2_X1 U7490 ( .A1(n5978), .A2(n6031), .ZN(n8107) );
  AOI22_X1 U7491 ( .A1(n8107), .A2(n6514), .B1(n7566), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n5979) );
  XNOR2_X1 U7492 ( .A(n8355), .B(n5763), .ZN(n7703) );
  NAND2_X1 U7493 ( .A1(n7603), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5988) );
  INV_X1 U7494 ( .A(n5991), .ZN(n5982) );
  NAND2_X1 U7495 ( .A1(n5982), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6037) );
  INV_X1 U7496 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U7497 ( .A1(n5991), .A2(n5983), .ZN(n5984) );
  AND2_X1 U7498 ( .A1(n6037), .A2(n5984), .ZN(n8354) );
  NAND2_X1 U7499 ( .A1(n5812), .A2(n8354), .ZN(n5987) );
  NAND2_X1 U7500 ( .A1(n7604), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7501 ( .A1(n4298), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5985) );
  INV_X1 U7502 ( .A(n8331), .ZN(n8013) );
  AND2_X1 U7503 ( .A1(n7809), .A2(n8013), .ZN(n6003) );
  INV_X1 U7504 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U7505 ( .A1(n5989), .A2(n9938), .ZN(n5990) );
  AND2_X1 U7506 ( .A1(n5991), .A2(n5990), .ZN(n7503) );
  NAND2_X1 U7507 ( .A1(n5812), .A2(n7503), .ZN(n5995) );
  NAND2_X1 U7508 ( .A1(n7603), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U7509 ( .A1(n7604), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U7510 ( .A1(n4298), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5992) );
  INV_X1 U7511 ( .A(n8344), .ZN(n8014) );
  AND2_X1 U7512 ( .A1(n7809), .A2(n8014), .ZN(n7700) );
  NAND2_X1 U7513 ( .A1(n6510), .A2(n7565), .ZN(n5999) );
  NAND2_X1 U7514 ( .A1(n5996), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5997) );
  XNOR2_X1 U7515 ( .A(n5997), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8091) );
  AOI22_X1 U7516 ( .A1(n8091), .A2(n6514), .B1(n7566), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5998) );
  XNOR2_X1 U7517 ( .A(n7793), .B(n5763), .ZN(n7699) );
  OAI22_X1 U7518 ( .A1(n7703), .A2(n6003), .B1(n7700), .B2(n7699), .ZN(n6000)
         );
  NAND2_X1 U7519 ( .A1(n7699), .A2(n7700), .ZN(n6001) );
  INV_X1 U7520 ( .A(n6003), .ZN(n7702) );
  NAND2_X1 U7521 ( .A1(n6001), .A2(n7702), .ZN(n6004) );
  INV_X1 U7522 ( .A(n6001), .ZN(n6002) );
  AOI22_X1 U7523 ( .A1(n7703), .A2(n6004), .B1(n6003), .B2(n6002), .ZN(n7657)
         );
  NAND2_X1 U7524 ( .A1(n6803), .A2(n7565), .ZN(n6006) );
  AOI22_X1 U7525 ( .A1(n8219), .A2(n6514), .B1(n7566), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n6005) );
  XNOR2_X1 U7526 ( .A(n8451), .B(n5763), .ZN(n6015) );
  INV_X1 U7527 ( .A(n6015), .ZN(n6013) );
  INV_X1 U7528 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7713) );
  INV_X1 U7529 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10019) );
  NAND2_X1 U7530 ( .A1(n6021), .A2(n10019), .ZN(n6008) );
  NAND2_X1 U7531 ( .A1(n6050), .A2(n6008), .ZN(n8308) );
  INV_X1 U7532 ( .A(n6224), .ZN(n6141) );
  INV_X1 U7533 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n6009) );
  OAI22_X1 U7534 ( .A1(n8308), .A2(n6141), .B1(n6411), .B2(n6009), .ZN(n6012)
         );
  INV_X1 U7535 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8139) );
  INV_X1 U7536 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6010) );
  OAI22_X1 U7537 ( .A1(n5751), .A2(n8139), .B1(n5834), .B2(n6010), .ZN(n6011)
         );
  NAND2_X1 U7538 ( .A1(n7809), .A2(n8011), .ZN(n6014) );
  NAND2_X1 U7539 ( .A1(n6013), .A2(n6014), .ZN(n6068) );
  INV_X1 U7540 ( .A(n6068), .ZN(n6045) );
  XNOR2_X1 U7541 ( .A(n6015), .B(n6014), .ZN(n7671) );
  NAND2_X1 U7542 ( .A1(n6678), .A2(n7565), .ZN(n6018) );
  NAND2_X1 U7543 ( .A1(n6033), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6016) );
  XNOR2_X1 U7544 ( .A(n6016), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8138) );
  AOI22_X1 U7545 ( .A1(n8138), .A2(n6514), .B1(n7566), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n6017) );
  XNOR2_X1 U7546 ( .A(n8455), .B(n5763), .ZN(n6026) );
  NAND2_X1 U7547 ( .A1(n7603), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6025) );
  INV_X1 U7548 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7549 ( .A1(n6039), .A2(n6019), .ZN(n6020) );
  AND2_X1 U7550 ( .A1(n6021), .A2(n6020), .ZN(n7768) );
  NAND2_X1 U7551 ( .A1(n6224), .A2(n7768), .ZN(n6024) );
  NAND2_X1 U7552 ( .A1(n7604), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7553 ( .A1(n4298), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6022) );
  INV_X1 U7554 ( .A(n7714), .ZN(n8327) );
  AND2_X1 U7555 ( .A1(n7809), .A2(n8327), .ZN(n6027) );
  NAND2_X1 U7556 ( .A1(n6026), .A2(n6027), .ZN(n6030) );
  AND2_X1 U7557 ( .A1(n7671), .A2(n6030), .ZN(n6044) );
  INV_X1 U7558 ( .A(n6026), .ZN(n7660) );
  INV_X1 U7559 ( .A(n6027), .ZN(n6028) );
  NAND2_X1 U7560 ( .A1(n7660), .A2(n6028), .ZN(n6029) );
  AND2_X1 U7561 ( .A1(n6030), .A2(n6029), .ZN(n6067) );
  INV_X1 U7562 ( .A(n6067), .ZN(n7759) );
  NAND2_X1 U7563 ( .A1(n6557), .A2(n7565), .ZN(n6036) );
  NAND2_X1 U7564 ( .A1(n6031), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6032) );
  MUX2_X1 U7565 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6032), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n6034) );
  AND2_X1 U7566 ( .A1(n6034), .A2(n6033), .ZN(n8122) );
  AOI22_X1 U7567 ( .A1(n8122), .A2(n6514), .B1(n7566), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n6035) );
  XNOR2_X1 U7568 ( .A(n8462), .B(n5763), .ZN(n6062) );
  NAND2_X1 U7569 ( .A1(n7603), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7570 ( .A1(n6037), .A2(n7713), .ZN(n6038) );
  AND2_X1 U7571 ( .A1(n6039), .A2(n6038), .ZN(n8334) );
  NAND2_X1 U7572 ( .A1(n5812), .A2(n8334), .ZN(n6042) );
  NAND2_X1 U7573 ( .A1(n7604), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U7574 ( .A1(n4298), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6040) );
  NAND4_X1 U7575 ( .A1(n6043), .A2(n6042), .A3(n6041), .A4(n6040), .ZN(n8012)
         );
  AND2_X1 U7576 ( .A1(n7809), .A2(n8012), .ZN(n6063) );
  NAND2_X1 U7577 ( .A1(n6062), .A2(n6063), .ZN(n6066) );
  OR2_X1 U7578 ( .A1(n7759), .A2(n6066), .ZN(n7659) );
  AND2_X1 U7579 ( .A1(n6044), .A2(n7659), .ZN(n7665) );
  OR2_X1 U7580 ( .A1(n6045), .A2(n7665), .ZN(n6061) );
  AND2_X1 U7581 ( .A1(n7657), .A2(n6061), .ZN(n7681) );
  NAND2_X1 U7582 ( .A1(n6835), .A2(n7565), .ZN(n6047) );
  NAND2_X1 U7583 ( .A1(n7566), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6046) );
  XNOR2_X1 U7584 ( .A(n8445), .B(n5763), .ZN(n6056) );
  INV_X1 U7585 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7586 ( .A1(n6050), .A2(n6049), .ZN(n6051) );
  NAND2_X1 U7587 ( .A1(n6076), .A2(n6051), .ZN(n8288) );
  OR2_X1 U7588 ( .A1(n8288), .A2(n6141), .ZN(n6054) );
  AOI22_X1 U7589 ( .A1(n7603), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n7604), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7590 ( .A1(n4298), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6052) );
  INV_X1 U7591 ( .A(n8277), .ZN(n8010) );
  AND2_X1 U7592 ( .A1(n7809), .A2(n8010), .ZN(n6057) );
  NAND2_X1 U7593 ( .A1(n6056), .A2(n6057), .ZN(n6060) );
  AND2_X1 U7594 ( .A1(n7681), .A2(n6060), .ZN(n6055) );
  NAND2_X1 U7595 ( .A1(n4309), .A2(n6055), .ZN(n6073) );
  INV_X1 U7596 ( .A(n6060), .ZN(n6072) );
  INV_X1 U7597 ( .A(n6056), .ZN(n7683) );
  INV_X1 U7598 ( .A(n6057), .ZN(n6058) );
  NAND2_X1 U7599 ( .A1(n7683), .A2(n6058), .ZN(n6059) );
  NAND2_X1 U7600 ( .A1(n6060), .A2(n6059), .ZN(n7733) );
  INV_X1 U7601 ( .A(n7733), .ZN(n6071) );
  INV_X1 U7602 ( .A(n6061), .ZN(n6070) );
  INV_X1 U7603 ( .A(n6062), .ZN(n7761) );
  INV_X1 U7604 ( .A(n6063), .ZN(n6064) );
  NAND2_X1 U7605 ( .A1(n7761), .A2(n6064), .ZN(n6065) );
  AND2_X1 U7606 ( .A1(n6066), .A2(n6065), .ZN(n7712) );
  AND2_X1 U7607 ( .A1(n7712), .A2(n6067), .ZN(n7658) );
  AND2_X1 U7608 ( .A1(n7658), .A2(n6068), .ZN(n6069) );
  OR2_X1 U7609 ( .A1(n6070), .A2(n6069), .ZN(n7731) );
  AND2_X1 U7610 ( .A1(n6071), .A2(n7731), .ZN(n7682) );
  NAND2_X1 U7611 ( .A1(n6902), .A2(n7565), .ZN(n6075) );
  NAND2_X1 U7612 ( .A1(n7566), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6074) );
  XNOR2_X1 U7613 ( .A(n8440), .B(n6124), .ZN(n6081) );
  INV_X1 U7614 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7686) );
  NAND2_X1 U7615 ( .A1(n6076), .A2(n7686), .ZN(n6077) );
  AND2_X1 U7616 ( .A1(n6088), .A2(n6077), .ZN(n8281) );
  NAND2_X1 U7617 ( .A1(n8281), .A2(n6224), .ZN(n6080) );
  AOI22_X1 U7618 ( .A1(n7603), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n7604), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7619 ( .A1(n4298), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6078) );
  INV_X1 U7620 ( .A(n8297), .ZN(n8265) );
  AND2_X1 U7621 ( .A1(n8265), .A2(n7809), .ZN(n6082) );
  INV_X1 U7622 ( .A(n6081), .ZN(n6083) );
  NAND2_X1 U7623 ( .A1(n6083), .A2(n6082), .ZN(n6098) );
  NAND2_X1 U7624 ( .A1(n6980), .A2(n7565), .ZN(n6085) );
  NAND2_X1 U7625 ( .A1(n7566), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6084) );
  XNOR2_X1 U7626 ( .A(n8434), .B(n6124), .ZN(n6097) );
  INV_X1 U7627 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7628 ( .A1(n6088), .A2(n6087), .ZN(n6089) );
  NAND2_X1 U7629 ( .A1(n6101), .A2(n6089), .ZN(n8259) );
  OR2_X1 U7630 ( .A1(n8259), .A2(n6141), .ZN(n6095) );
  INV_X1 U7631 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7632 ( .A1(n7603), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7633 ( .A1(n7604), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6090) );
  OAI211_X1 U7634 ( .C1(n6092), .C2(n6411), .A(n6091), .B(n6090), .ZN(n6093)
         );
  INV_X1 U7635 ( .A(n6093), .ZN(n6094) );
  NAND2_X1 U7636 ( .A1(n7597), .A2(n7809), .ZN(n7741) );
  AND2_X1 U7637 ( .A1(n6098), .A2(n6097), .ZN(n6099) );
  AND2_X1 U7638 ( .A1(n6096), .A2(n6099), .ZN(n6100) );
  INV_X1 U7639 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7642) );
  NAND2_X1 U7640 ( .A1(n6101), .A2(n7642), .ZN(n6102) );
  AND2_X1 U7641 ( .A1(n6125), .A2(n6102), .ZN(n8246) );
  INV_X1 U7642 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7643 ( .A1(n7603), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7644 ( .A1(n7604), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6103) );
  OAI211_X1 U7645 ( .C1(n6105), .C2(n6411), .A(n6104), .B(n6103), .ZN(n6106)
         );
  AOI21_X1 U7646 ( .B1(n8246), .B2(n6224), .A(n6106), .ZN(n7745) );
  INV_X1 U7647 ( .A(n7809), .ZN(n6177) );
  NOR2_X1 U7648 ( .A1(n7745), .A2(n6177), .ZN(n7640) );
  NAND2_X1 U7649 ( .A1(n7132), .A2(n7565), .ZN(n6108) );
  NAND2_X1 U7650 ( .A1(n7566), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6107) );
  XNOR2_X1 U7651 ( .A(n8422), .B(n5763), .ZN(n6117) );
  XNOR2_X1 U7652 ( .A(n6125), .B(P2_REG3_REG_24__SCAN_IN), .ZN(n8227) );
  NAND2_X1 U7653 ( .A1(n8227), .A2(n6224), .ZN(n6113) );
  INV_X1 U7654 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9876) );
  NAND2_X1 U7655 ( .A1(n7603), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U7656 ( .A1(n7604), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6109) );
  OAI211_X1 U7657 ( .C1(n9876), .C2(n6411), .A(n6110), .B(n6109), .ZN(n6111)
         );
  INV_X1 U7658 ( .A(n6111), .ZN(n6112) );
  INV_X1 U7659 ( .A(n8242), .ZN(n8009) );
  NAND3_X1 U7660 ( .A1(n7641), .A2(n7640), .A3(n6114), .ZN(n6121) );
  NOR2_X1 U7661 ( .A1(n8242), .A2(n6177), .ZN(n6118) );
  AND2_X1 U7662 ( .A1(n6116), .A2(n6115), .ZN(n7719) );
  OAI21_X1 U7663 ( .B1(n6118), .B2(n6117), .A(n7719), .ZN(n6119) );
  INV_X1 U7664 ( .A(n6117), .ZN(n7721) );
  INV_X1 U7665 ( .A(n6118), .ZN(n7724) );
  NAND2_X1 U7666 ( .A1(n7421), .A2(n7565), .ZN(n6123) );
  OR2_X1 U7667 ( .A1(n5793), .A2(n9922), .ZN(n6122) );
  XNOR2_X1 U7668 ( .A(n8419), .B(n6124), .ZN(n7774) );
  INV_X1 U7669 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n7726) );
  OAI21_X1 U7670 ( .B1(n6125), .B2(n7726), .A(n9962), .ZN(n6128) );
  INV_X1 U7671 ( .A(n6125), .ZN(n6127) );
  AND2_X1 U7672 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_24__SCAN_IN), 
        .ZN(n6126) );
  NAND2_X1 U7673 ( .A1(n6127), .A2(n6126), .ZN(n6139) );
  NAND2_X1 U7674 ( .A1(n6128), .A2(n6139), .ZN(n8217) );
  OR2_X1 U7675 ( .A1(n8217), .A2(n6141), .ZN(n6134) );
  INV_X1 U7676 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7677 ( .A1(n4298), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U7678 ( .A1(n7604), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6129) );
  OAI211_X1 U7679 ( .C1(n5751), .C2(n6131), .A(n6130), .B(n6129), .ZN(n6132)
         );
  INV_X1 U7680 ( .A(n6132), .ZN(n6133) );
  NAND2_X1 U7681 ( .A1(n8233), .A2(n7809), .ZN(n6135) );
  NOR2_X1 U7682 ( .A1(n7774), .A2(n6135), .ZN(n6136) );
  AOI21_X1 U7683 ( .B1(n7774), .B2(n6135), .A(n6136), .ZN(n7691) );
  NAND2_X1 U7684 ( .A1(n7398), .A2(n7565), .ZN(n6138) );
  NAND2_X1 U7685 ( .A1(n7566), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6137) );
  XNOR2_X1 U7686 ( .A(n8414), .B(n5763), .ZN(n6148) );
  INV_X1 U7687 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U7688 ( .A1(n6139), .A2(n9948), .ZN(n6140) );
  NAND2_X1 U7689 ( .A1(n6171), .A2(n6140), .ZN(n7779) );
  OR2_X1 U7690 ( .A1(n7779), .A2(n6141), .ZN(n6147) );
  INV_X1 U7691 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7692 ( .A1(n7603), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6143) );
  NAND2_X1 U7693 ( .A1(n7604), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6142) );
  OAI211_X1 U7694 ( .C1(n6144), .C2(n6411), .A(n6143), .B(n6142), .ZN(n6145)
         );
  INV_X1 U7695 ( .A(n6145), .ZN(n6146) );
  NOR2_X1 U7696 ( .A1(n8008), .A2(n6177), .ZN(n6149) );
  NAND2_X1 U7697 ( .A1(n6148), .A2(n6149), .ZN(n6152) );
  INV_X1 U7698 ( .A(n6148), .ZN(n7631) );
  INV_X1 U7699 ( .A(n6149), .ZN(n6150) );
  NAND2_X1 U7700 ( .A1(n7631), .A2(n6150), .ZN(n6151) );
  NAND2_X1 U7701 ( .A1(n6152), .A2(n6151), .ZN(n7775) );
  NAND2_X1 U7702 ( .A1(n7494), .A2(n7565), .ZN(n6154) );
  NAND2_X1 U7703 ( .A1(n7566), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6153) );
  XNOR2_X1 U7704 ( .A(n8407), .B(n5763), .ZN(n6161) );
  XNOR2_X1 U7705 ( .A(n6171), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8178) );
  NAND2_X1 U7706 ( .A1(n8178), .A2(n6224), .ZN(n6160) );
  INV_X1 U7707 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6157) );
  NAND2_X1 U7708 ( .A1(n7603), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U7709 ( .A1(n4298), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6155) );
  OAI211_X1 U7710 ( .C1(n5834), .C2(n6157), .A(n6156), .B(n6155), .ZN(n6158)
         );
  INV_X1 U7711 ( .A(n6158), .ZN(n6159) );
  AND2_X1 U7712 ( .A1(n8007), .A2(n7809), .ZN(n6162) );
  NAND2_X1 U7713 ( .A1(n6161), .A2(n6162), .ZN(n6166) );
  INV_X1 U7714 ( .A(n6161), .ZN(n6164) );
  INV_X1 U7715 ( .A(n6162), .ZN(n6163) );
  NAND2_X1 U7716 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  NAND2_X1 U7717 ( .A1(n7512), .A2(n7565), .ZN(n6168) );
  NAND2_X1 U7718 ( .A1(n7566), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6167) );
  INV_X1 U7719 ( .A(n5732), .ZN(n6169) );
  NAND2_X1 U7720 ( .A1(n8402), .A2(n9799), .ZN(n6215) );
  NAND2_X1 U7721 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6170) );
  INV_X1 U7722 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7635) );
  INV_X1 U7723 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6235) );
  OAI21_X1 U7724 ( .B1(n6171), .B2(n7635), .A(n6235), .ZN(n6172) );
  INV_X1 U7725 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7726 ( .A1(n7603), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7727 ( .A1(n7604), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6173) );
  OAI211_X1 U7728 ( .C1(n6175), .C2(n6411), .A(n6174), .B(n6173), .ZN(n6176)
         );
  OR2_X1 U7729 ( .A1(n8006), .A2(n6177), .ZN(n6178) );
  XNOR2_X1 U7730 ( .A(n6178), .B(n5763), .ZN(n6216) );
  MUX2_X1 U7731 ( .A(n6215), .B(n8402), .S(n6216), .Z(n6214) );
  INV_X1 U7732 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U7733 ( .A1(n6188), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6184) );
  MUX2_X1 U7734 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6184), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6185) );
  OR2_X1 U7735 ( .A1(n7133), .A2(n7399), .ZN(n9709) );
  NAND2_X1 U7736 ( .A1(n6186), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6187) );
  MUX2_X1 U7737 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6187), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6189) );
  AND2_X1 U7738 ( .A1(n6189), .A2(n6188), .ZN(n7422) );
  XNOR2_X1 U7739 ( .A(n7133), .B(P2_B_REG_SCAN_IN), .ZN(n6190) );
  INV_X1 U7740 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U7741 ( .A1(n9706), .A2(n6192), .ZN(n6193) );
  INV_X1 U7742 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9713) );
  NOR2_X1 U7743 ( .A1(n7422), .A2(n7399), .ZN(n9714) );
  NOR4_X1 U7744 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6197) );
  NOR4_X1 U7745 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6196) );
  NOR4_X1 U7746 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n6195) );
  NOR4_X1 U7747 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6194) );
  NAND4_X1 U7748 ( .A1(n6197), .A2(n6196), .A3(n6195), .A4(n6194), .ZN(n6203)
         );
  NOR2_X1 U7749 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .ZN(
        n6201) );
  NOR4_X1 U7750 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6200) );
  NOR4_X1 U7751 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6199) );
  NOR4_X1 U7752 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n6198) );
  NAND4_X1 U7753 ( .A1(n6201), .A2(n6200), .A3(n6199), .A4(n6198), .ZN(n6202)
         );
  NAND2_X1 U7754 ( .A1(n8391), .A2(n8390), .ZN(n7178) );
  INV_X1 U7755 ( .A(n6230), .ZN(n6209) );
  AND2_X1 U7756 ( .A1(n7399), .A2(n7422), .ZN(n6204) );
  OR2_X1 U7757 ( .A1(n6206), .A2(n6205), .ZN(n6207) );
  NAND2_X1 U7758 ( .A1(n6208), .A2(n6207), .ZN(n6231) );
  NAND2_X1 U7759 ( .A1(n6209), .A2(n9708), .ZN(n6226) );
  OR2_X1 U7760 ( .A1(n7999), .A2(n8394), .ZN(n6210) );
  NAND2_X1 U7761 ( .A1(n6226), .A2(n6210), .ZN(n6211) );
  OAI21_X1 U7762 ( .B1(n8164), .B2(n9687), .A(n9431), .ZN(n6213) );
  OAI21_X1 U7763 ( .B1(n6219), .B2(n6214), .A(n6213), .ZN(n6240) );
  INV_X1 U7764 ( .A(n6215), .ZN(n6217) );
  MUX2_X1 U7765 ( .A(n8164), .B(n6217), .S(n6216), .Z(n6218) );
  INV_X1 U7766 ( .A(n7612), .ZN(n6225) );
  INV_X1 U7767 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6222) );
  NAND2_X1 U7768 ( .A1(n7603), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6221) );
  NAND2_X1 U7769 ( .A1(n7604), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6220) );
  OAI211_X1 U7770 ( .C1(n6222), .C2(n6411), .A(n6221), .B(n6220), .ZN(n6223)
         );
  AOI21_X1 U7771 ( .B1(n6225), .B2(n6224), .A(n6223), .ZN(n8168) );
  INV_X1 U7772 ( .A(n6226), .ZN(n6228) );
  INV_X1 U7773 ( .A(n7997), .ZN(n6227) );
  INV_X1 U7774 ( .A(n6229), .ZN(n6752) );
  OR2_X2 U7775 ( .A1(n6516), .A2(n6229), .ZN(n8372) );
  INV_X1 U7776 ( .A(n8007), .ZN(n8169) );
  OAI22_X1 U7777 ( .A1(n8168), .A2(n7790), .B1(n7789), .B2(n8169), .ZN(n6238)
         );
  NAND2_X1 U7778 ( .A1(n6230), .A2(n8389), .ZN(n7584) );
  INV_X1 U7779 ( .A(n6231), .ZN(n6513) );
  OR2_X1 U7780 ( .A1(n7177), .A2(n6513), .ZN(n6232) );
  NOR2_X1 U7781 ( .A1(n6697), .A2(n6232), .ZN(n6233) );
  NAND2_X1 U7782 ( .A1(n7584), .A2(n6233), .ZN(n6234) );
  INV_X1 U7783 ( .A(n8162), .ZN(n6236) );
  OAI22_X1 U7784 ( .A1(n9693), .A2(n6236), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6235), .ZN(n6237) );
  OAI21_X1 U7785 ( .B1(n6240), .B2(n6239), .A(n4841), .ZN(P2_U3222) );
  INV_X1 U7786 ( .A(n6241), .ZN(n7073) );
  NOR2_X1 U7787 ( .A1(n5057), .A2(n7073), .ZN(n6286) );
  NAND2_X1 U7788 ( .A1(n5057), .A2(n8776), .ZN(n6242) );
  NAND2_X1 U7789 ( .A1(n6242), .A2(n6241), .ZN(n6303) );
  NAND2_X1 U7790 ( .A1(n6303), .A2(n6302), .ZN(n6243) );
  NAND2_X1 U7791 ( .A1(n6243), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X2 U7792 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  AND2_X1 U7793 ( .A1(n7548), .A2(P2_U3152), .ZN(n8491) );
  INV_X1 U7794 ( .A(n8491), .ZN(n7628) );
  NOR2_X1 U7795 ( .A1(n7554), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7619) );
  OAI222_X1 U7796 ( .A1(n7628), .A2(n6244), .B1(n7626), .B2(n6246), .C1(
        P2_U3152), .C2(n6737), .ZN(P2_U3357) );
  NOR2_X1 U7797 ( .A1(n7548), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9357) );
  AND2_X1 U7798 ( .A1(n7554), .A2(P1_U3084), .ZN(n7071) );
  INV_X2 U7799 ( .A(n7071), .ZN(n9364) );
  OAI222_X1 U7800 ( .A1(n9360), .A2(n6245), .B1(n9364), .B2(n6261), .C1(
        P1_U3084), .C2(n6288), .ZN(P1_U3350) );
  OAI222_X1 U7801 ( .A1(n9360), .A2(n10032), .B1(n9364), .B2(n6263), .C1(
        P1_U3084), .C2(n9508), .ZN(P1_U3351) );
  INV_X1 U7802 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6247) );
  OAI222_X1 U7803 ( .A1(n9360), .A2(n6247), .B1(n9364), .B2(n6246), .C1(
        P1_U3084), .C2(n9495), .ZN(P1_U3352) );
  OAI222_X1 U7804 ( .A1(n9360), .A2(n6249), .B1(n9364), .B2(n6257), .C1(
        P1_U3084), .C2(n6248), .ZN(P1_U3349) );
  OAI222_X1 U7805 ( .A1(n9360), .A2(n6250), .B1(n9364), .B2(n6259), .C1(
        P1_U3084), .C2(n9542), .ZN(P1_U3348) );
  NAND2_X1 U7806 ( .A1(n6320), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6251) );
  OAI21_X1 U7807 ( .B1(n6330), .B2(n6320), .A(n6251), .ZN(P1_U3441) );
  OAI222_X1 U7808 ( .A1(n9360), .A2(n6253), .B1(n9364), .B2(n6255), .C1(
        P1_U3084), .C2(n6252), .ZN(P1_U3347) );
  NAND2_X1 U7809 ( .A1(n6353), .A2(n9657), .ZN(n6254) );
  OAI21_X1 U7810 ( .B1(n9657), .B2(n5640), .A(n6254), .ZN(P1_U3440) );
  OAI222_X1 U7811 ( .A1(n7628), .A2(n6256), .B1(n7626), .B2(n6255), .C1(
        P2_U3152), .C2(n6802), .ZN(P2_U3352) );
  OAI222_X1 U7812 ( .A1(n7628), .A2(n6258), .B1(n7626), .B2(n6257), .C1(
        P2_U3152), .C2(n8046), .ZN(P2_U3354) );
  INV_X1 U7813 ( .A(n6732), .ZN(n8060) );
  OAI222_X1 U7814 ( .A1(n7628), .A2(n6260), .B1(n7626), .B2(n6259), .C1(
        P2_U3152), .C2(n8060), .ZN(P2_U3353) );
  OAI222_X1 U7815 ( .A1(n7628), .A2(n6262), .B1(n7626), .B2(n6261), .C1(
        P2_U3152), .C2(n8032), .ZN(P2_U3355) );
  OAI222_X1 U7816 ( .A1(n7628), .A2(n6264), .B1(n7626), .B2(n6263), .C1(
        P2_U3152), .C2(n6741), .ZN(P2_U3356) );
  INV_X1 U7817 ( .A(n6265), .ZN(n6274) );
  AOI22_X1 U7818 ( .A1(n9571), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9357), .ZN(n6266) );
  OAI21_X1 U7819 ( .B1(n6274), .B2(n9364), .A(n6266), .ZN(P1_U3346) );
  INV_X1 U7820 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U7821 ( .A1(n6267), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U7822 ( .A1(n8625), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U7823 ( .A1(n6268), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6269) );
  NAND3_X1 U7824 ( .A1(n6271), .A2(n6270), .A3(n6269), .ZN(n8944) );
  NAND2_X1 U7825 ( .A1(n8944), .A2(P1_U4006), .ZN(n6272) );
  OAI21_X1 U7826 ( .B1(P1_U4006), .B2(n6273), .A(n6272), .ZN(P1_U3586) );
  INV_X1 U7827 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6275) );
  INV_X1 U7828 ( .A(n6727), .ZN(n6770) );
  OAI222_X1 U7829 ( .A1(n7628), .A2(n6275), .B1(n7626), .B2(n6274), .C1(
        P2_U3152), .C2(n6770), .ZN(P2_U3351) );
  INV_X1 U7830 ( .A(n6276), .ZN(n6278) );
  AOI22_X1 U7831 ( .A1(n9584), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9357), .ZN(n6277) );
  OAI21_X1 U7832 ( .B1(n6278), .B2(n9364), .A(n6277), .ZN(P1_U3345) );
  INV_X1 U7833 ( .A(n6724), .ZN(n6781) );
  OAI222_X1 U7834 ( .A1(n7628), .A2(n6279), .B1(n7626), .B2(n6278), .C1(
        P2_U3152), .C2(n6781), .ZN(P2_U3350) );
  INV_X1 U7835 ( .A(n6280), .ZN(n6282) );
  AOI22_X1 U7836 ( .A1(n9600), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9357), .ZN(n6281) );
  OAI21_X1 U7837 ( .B1(n6282), .B2(n9364), .A(n6281), .ZN(P1_U3344) );
  OAI222_X1 U7838 ( .A1(n7628), .A2(n6283), .B1(n7626), .B2(n6282), .C1(n4521), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U7839 ( .A(n6285), .ZN(n9490) );
  NOR2_X1 U7840 ( .A1(n6285), .A2(P1_U3084), .ZN(n7495) );
  NAND2_X1 U7841 ( .A1(n6303), .A2(n7495), .ZN(n6293) );
  INV_X1 U7842 ( .A(n9621), .ZN(n9634) );
  NAND2_X1 U7843 ( .A1(n9634), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U7844 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6367) );
  OAI211_X1 U7845 ( .C1(n9543), .C2(n6288), .A(n6287), .B(n6367), .ZN(n6308)
         );
  INV_X1 U7846 ( .A(n9508), .ZN(n6300) );
  INV_X1 U7847 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9489) );
  NOR2_X1 U7848 ( .A1(n6297), .A2(n9489), .ZN(n9521) );
  INV_X1 U7849 ( .A(n9521), .ZN(n9500) );
  NAND2_X1 U7850 ( .A1(P1_REG2_REG_1__SCAN_IN), .A2(n6298), .ZN(n6289) );
  OAI21_X1 U7851 ( .B1(n6298), .B2(P1_REG2_REG_1__SCAN_IN), .A(n6289), .ZN(
        n9499) );
  NOR2_X1 U7852 ( .A1(n9500), .A2(n9499), .ZN(n9498) );
  AOI21_X1 U7853 ( .B1(n6298), .B2(P1_REG2_REG_1__SCAN_IN), .A(n9498), .ZN(
        n9513) );
  INV_X1 U7854 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6290) );
  MUX2_X1 U7855 ( .A(n6290), .B(P1_REG2_REG_2__SCAN_IN), .S(n9508), .Z(n6291)
         );
  INV_X1 U7856 ( .A(n6291), .ZN(n9512) );
  NOR2_X1 U7857 ( .A1(n9513), .A2(n9512), .ZN(n9511) );
  AOI21_X1 U7858 ( .B1(n6300), .B2(P1_REG2_REG_2__SCAN_IN), .A(n9511), .ZN(
        n6296) );
  NAND2_X1 U7859 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(n6390), .ZN(n6292) );
  OAI21_X1 U7860 ( .B1(n6390), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6292), .ZN(
        n6295) );
  NOR2_X1 U7861 ( .A1(n6296), .A2(n6295), .ZN(n6389) );
  INV_X1 U7862 ( .A(n6293), .ZN(n6294) );
  AOI211_X1 U7863 ( .C1(n6296), .C2(n6295), .A(n6389), .B(n9623), .ZN(n6307)
         );
  XNOR2_X1 U7864 ( .A(n6298), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9502) );
  NOR3_X1 U7865 ( .A1(n6297), .A2(n5064), .A3(n9502), .ZN(n9501) );
  AOI21_X1 U7866 ( .B1(n6298), .B2(P1_REG1_REG_1__SCAN_IN), .A(n9501), .ZN(
        n9516) );
  INV_X1 U7867 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6299) );
  MUX2_X1 U7868 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6299), .S(n9508), .Z(n9515)
         );
  NOR2_X1 U7869 ( .A1(n9516), .A2(n9515), .ZN(n9514) );
  AOI21_X1 U7870 ( .B1(n6300), .B2(P1_REG1_REG_2__SCAN_IN), .A(n9514), .ZN(
        n6305) );
  NAND2_X1 U7871 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(n6390), .ZN(n6301) );
  OAI21_X1 U7872 ( .B1(n6390), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6301), .ZN(
        n6304) );
  NOR2_X1 U7873 ( .A1(n6305), .A2(n6304), .ZN(n6381) );
  AND3_X1 U7874 ( .A1(n6303), .A2(P1_STATE_REG_SCAN_IN), .A3(n6302), .ZN(n9492) );
  NAND2_X1 U7875 ( .A1(n9492), .A2(n6285), .ZN(n9549) );
  AOI211_X1 U7876 ( .C1(n6305), .C2(n6304), .A(n6381), .B(n9549), .ZN(n6306)
         );
  OR3_X1 U7877 ( .A1(n6308), .A2(n6307), .A3(n6306), .ZN(P1_U3244) );
  INV_X1 U7878 ( .A(n6309), .ZN(n6311) );
  AOI22_X1 U7879 ( .A1(n6427), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9357), .ZN(n6310) );
  OAI21_X1 U7880 ( .B1(n6311), .B2(n9364), .A(n6310), .ZN(P1_U3343) );
  INV_X1 U7881 ( .A(n6825), .ZN(n6758) );
  OAI222_X1 U7882 ( .A1(n7628), .A2(n6312), .B1(n7626), .B2(n6311), .C1(n6758), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7883 ( .A(n6313), .ZN(n6316) );
  INV_X1 U7884 ( .A(n6608), .ZN(n6429) );
  OAI222_X1 U7885 ( .A1(n9364), .A2(n6316), .B1(n6429), .B2(P1_U3084), .C1(
        n6314), .C2(n9360), .ZN(P1_U3342) );
  INV_X1 U7886 ( .A(n6878), .ZN(n6831) );
  OAI222_X1 U7887 ( .A1(P2_U3152), .A2(n6831), .B1(n7626), .B2(n6316), .C1(
        n6315), .C2(n7628), .ZN(P2_U3347) );
  INV_X1 U7888 ( .A(n6317), .ZN(n6342) );
  AOI22_X1 U7889 ( .A1(n6688), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9357), .ZN(n6318) );
  OAI21_X1 U7890 ( .B1(n6342), .B2(n9364), .A(n6318), .ZN(P1_U3341) );
  OR2_X1 U7891 ( .A1(n6320), .A2(n6319), .ZN(n6352) );
  INV_X1 U7892 ( .A(n6352), .ZN(n6322) );
  OAI211_X1 U7893 ( .C1(n6323), .C2(n9330), .A(n6322), .B(n6321), .ZN(n7575)
         );
  AOI22_X1 U7894 ( .A1(n8578), .A2(n8891), .B1(n7575), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6327) );
  AOI22_X1 U7895 ( .A1(n8617), .A2(n4297), .B1(n8595), .B2(n9519), .ZN(n6326)
         );
  NAND2_X1 U7896 ( .A1(n6327), .A2(n6326), .ZN(P1_U3230) );
  NOR2_X1 U7897 ( .A1(n6352), .A2(n6328), .ZN(n6331) );
  INV_X1 U7898 ( .A(n6353), .ZN(n6332) );
  INV_X1 U7899 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6338) );
  INV_X1 U7900 ( .A(n4297), .ZN(n6443) );
  INV_X1 U7901 ( .A(n8891), .ZN(n8838) );
  NOR2_X1 U7902 ( .A1(n8892), .A2(n6443), .ZN(n6461) );
  INV_X1 U7903 ( .A(n6461), .ZN(n6333) );
  NAND2_X1 U7904 ( .A1(n6443), .A2(n8892), .ZN(n8837) );
  NAND2_X1 U7905 ( .A1(n6333), .A2(n8837), .ZN(n8753) );
  NAND3_X1 U7906 ( .A1(n8753), .A2(n6441), .A3(n6336), .ZN(n6334) );
  OAI21_X1 U7907 ( .B1(n8838), .B2(n9394), .A(n6334), .ZN(n6361) );
  INV_X1 U7908 ( .A(n6361), .ZN(n6335) );
  OAI21_X1 U7909 ( .B1(n6443), .B2(n6336), .A(n6335), .ZN(n6340) );
  NAND2_X1 U7910 ( .A1(n6340), .A2(n9352), .ZN(n6337) );
  OAI21_X1 U7911 ( .B1(n9352), .B2(n6338), .A(n6337), .ZN(P1_U3454) );
  NAND2_X1 U7912 ( .A1(n6340), .A2(n9334), .ZN(n6341) );
  OAI21_X1 U7913 ( .B1(n9334), .B2(n5064), .A(n6341), .ZN(P1_U3523) );
  INV_X1 U7914 ( .A(n6963), .ZN(n6886) );
  OAI222_X1 U7915 ( .A1(n7628), .A2(n6343), .B1(n7626), .B2(n6342), .C1(
        P2_U3152), .C2(n6886), .ZN(P2_U3346) );
  XNOR2_X1 U7916 ( .A(n6345), .B(n6344), .ZN(n6347) );
  XNOR2_X1 U7917 ( .A(n6347), .B(n6346), .ZN(n6350) );
  AOI22_X1 U7918 ( .A1(n6453), .A2(n8617), .B1(n8611), .B2(n8892), .ZN(n6349)
         );
  AOI22_X1 U7919 ( .A1(n8578), .A2(n8889), .B1(n7575), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6348) );
  OAI211_X1 U7920 ( .C1(n6350), .C2(n8619), .A(n6349), .B(n6348), .ZN(P1_U3220) );
  INV_X1 U7921 ( .A(n5938), .ZN(n6372) );
  AOI22_X1 U7922 ( .A1(n7145), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9357), .ZN(n6351) );
  OAI21_X1 U7923 ( .B1(n6372), .B2(n9364), .A(n6351), .ZN(P1_U3340) );
  NOR2_X1 U7924 ( .A1(n6353), .A2(n6352), .ZN(n6354) );
  NAND2_X1 U7925 ( .A1(n6355), .A2(n6354), .ZN(n6659) );
  INV_X1 U7926 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6356) );
  OAI22_X1 U7927 ( .A1(n9653), .A2(n9489), .B1(n6356), .B2(n9644), .ZN(n6360)
         );
  INV_X1 U7928 ( .A(n6357), .ZN(n6358) );
  INV_X1 U7929 ( .A(n9237), .ZN(n8948) );
  NAND2_X2 U7930 ( .A1(n9653), .A2(n9640), .ZN(n9217) );
  AOI21_X1 U7931 ( .B1(n8948), .B2(n9217), .A(n6443), .ZN(n6359) );
  AOI211_X1 U7932 ( .C1(n9653), .C2(n6361), .A(n6360), .B(n6359), .ZN(n6362)
         );
  INV_X1 U7933 ( .A(n6362), .ZN(P1_U3291) );
  INV_X1 U7934 ( .A(n6363), .ZN(n7573) );
  NOR3_X1 U7935 ( .A1(n7573), .A2(n4768), .A3(n6365), .ZN(n6366) );
  OAI21_X1 U7936 ( .B1(n6366), .B2(n4376), .A(n8595), .ZN(n6371) );
  INV_X1 U7937 ( .A(n6367), .ZN(n6369) );
  OAI22_X1 U7938 ( .A1(n6574), .A2(n8615), .B1(n8599), .B2(n6456), .ZN(n6368)
         );
  AOI211_X1 U7939 ( .C1(n6498), .C2(n8617), .A(n6369), .B(n6368), .ZN(n6370)
         );
  OAI211_X1 U7940 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8588), .A(n6371), .B(
        n6370), .ZN(P1_U3216) );
  INV_X1 U7941 ( .A(n7091), .ZN(n7086) );
  OAI222_X1 U7942 ( .A1(n7628), .A2(n6373), .B1(n7626), .B2(n6372), .C1(n7086), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U7943 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6374) );
  MUX2_X1 U7944 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6374), .S(n6427), .Z(n6383)
         );
  NOR2_X1 U7945 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n9600), .ZN(n6375) );
  AOI21_X1 U7946 ( .B1(n9600), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6375), .ZN(
        n9602) );
  NOR2_X1 U7947 ( .A1(n9584), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6376) );
  AOI21_X1 U7948 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9584), .A(n6376), .ZN(
        n9587) );
  NOR2_X1 U7949 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n9571), .ZN(n6377) );
  AOI21_X1 U7950 ( .B1(n9571), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6377), .ZN(
        n9574) );
  NOR2_X1 U7951 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(n9567), .ZN(n6378) );
  AOI21_X1 U7952 ( .B1(n9567), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6378), .ZN(
        n9560) );
  NAND2_X1 U7953 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6392), .ZN(n6379) );
  OAI21_X1 U7954 ( .B1(n6392), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6379), .ZN(
        n9551) );
  NOR2_X1 U7955 ( .A1(P1_REG1_REG_4__SCAN_IN), .A2(n9531), .ZN(n6380) );
  AOI21_X1 U7956 ( .B1(n9531), .B2(P1_REG1_REG_4__SCAN_IN), .A(n6380), .ZN(
        n9530) );
  AOI21_X1 U7957 ( .B1(n6390), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6381), .ZN(
        n9529) );
  NAND2_X1 U7958 ( .A1(n9530), .A2(n9529), .ZN(n9528) );
  OAI21_X1 U7959 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9531), .A(n9528), .ZN(
        n9552) );
  NOR2_X1 U7960 ( .A1(n9551), .A2(n9552), .ZN(n9550) );
  AOI21_X1 U7961 ( .B1(n6392), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9550), .ZN(
        n9559) );
  NAND2_X1 U7962 ( .A1(n9560), .A2(n9559), .ZN(n9558) );
  OAI21_X1 U7963 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n9567), .A(n9558), .ZN(
        n9573) );
  NAND2_X1 U7964 ( .A1(n9574), .A2(n9573), .ZN(n9572) );
  OAI21_X1 U7965 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n9571), .A(n9572), .ZN(
        n9586) );
  NAND2_X1 U7966 ( .A1(n9587), .A2(n9586), .ZN(n9585) );
  OAI21_X1 U7967 ( .B1(n9584), .B2(P1_REG1_REG_8__SCAN_IN), .A(n9585), .ZN(
        n9603) );
  NAND2_X1 U7968 ( .A1(n9602), .A2(n9603), .ZN(n9601) );
  OAI21_X1 U7969 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9600), .A(n9601), .ZN(
        n6382) );
  NAND2_X1 U7970 ( .A1(n6382), .A2(n6383), .ZN(n6422) );
  OAI21_X1 U7971 ( .B1(n6383), .B2(n6382), .A(n6422), .ZN(n6402) );
  INV_X1 U7972 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6384) );
  NOR2_X1 U7973 ( .A1(n9621), .A2(n6384), .ZN(n6401) );
  INV_X1 U7974 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6385) );
  XNOR2_X1 U7975 ( .A(n6427), .B(n6385), .ZN(n6397) );
  NAND2_X1 U7976 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n9600), .ZN(n6395) );
  OAI21_X1 U7977 ( .B1(n9600), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6395), .ZN(
        n9596) );
  NOR2_X1 U7978 ( .A1(n9584), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6386) );
  AOI21_X1 U7979 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9584), .A(n6386), .ZN(
        n9590) );
  NOR2_X1 U7980 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n9571), .ZN(n6387) );
  AOI21_X1 U7981 ( .B1(n9571), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6387), .ZN(
        n9577) );
  NOR2_X1 U7982 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6392), .ZN(n6388) );
  AOI21_X1 U7983 ( .B1(n6392), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6388), .ZN(
        n9548) );
  AOI21_X1 U7984 ( .B1(n6390), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6389), .ZN(
        n9534) );
  NOR2_X1 U7985 ( .A1(P1_REG2_REG_4__SCAN_IN), .A2(n9531), .ZN(n6391) );
  AOI21_X1 U7986 ( .B1(n9531), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6391), .ZN(
        n9535) );
  NAND2_X1 U7987 ( .A1(n9534), .A2(n9535), .ZN(n9533) );
  OAI21_X1 U7988 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9531), .A(n9533), .ZN(
        n9547) );
  NAND2_X1 U7989 ( .A1(n9548), .A2(n9547), .ZN(n9546) );
  OAI21_X1 U7990 ( .B1(n6392), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9546), .ZN(
        n9564) );
  NAND2_X1 U7991 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(n9567), .ZN(n6393) );
  OAI21_X1 U7992 ( .B1(n9567), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6393), .ZN(
        n9563) );
  NOR2_X1 U7993 ( .A1(n9564), .A2(n9563), .ZN(n9562) );
  OAI21_X1 U7994 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9584), .A(n9588), .ZN(
        n9597) );
  NOR2_X1 U7995 ( .A1(n9596), .A2(n9597), .ZN(n9595) );
  INV_X1 U7996 ( .A(n9595), .ZN(n6394) );
  OAI211_X1 U7997 ( .C1(n6397), .C2(n6396), .A(n9616), .B(n4368), .ZN(n6399)
         );
  NAND2_X1 U7998 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6951) );
  NAND2_X1 U7999 ( .A1(n9629), .A2(n6427), .ZN(n6398) );
  NAND3_X1 U8000 ( .A1(n6399), .A2(n6951), .A3(n6398), .ZN(n6400) );
  AOI211_X1 U8001 ( .C1(n6402), .C2(n9635), .A(n6401), .B(n6400), .ZN(n6403)
         );
  INV_X1 U8002 ( .A(n6403), .ZN(P1_U3251) );
  INV_X1 U8003 ( .A(n6404), .ZN(n6406) );
  OAI222_X1 U8004 ( .A1(n9364), .A2(n6406), .B1(n7143), .B2(P1_U3084), .C1(
        n6405), .C2(n9360), .ZN(P1_U3339) );
  INV_X1 U8005 ( .A(n8073), .ZN(n7095) );
  OAI222_X1 U8006 ( .A1(n7628), .A2(n6407), .B1(n7626), .B2(n6406), .C1(n7095), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8007 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6413) );
  INV_X1 U8008 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6410) );
  NAND2_X1 U8009 ( .A1(n7603), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6409) );
  NAND2_X1 U8010 ( .A1(n7604), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6408) );
  OAI211_X1 U8011 ( .C1(n6411), .C2(n6410), .A(n6409), .B(n6408), .ZN(n7803)
         );
  NAND2_X1 U8012 ( .A1(n7803), .A2(P2_U3966), .ZN(n6412) );
  OAI21_X1 U8013 ( .B1(n6413), .B2(P2_U3966), .A(n6412), .ZN(P2_U3583) );
  INV_X1 U8014 ( .A(n6414), .ZN(n6491) );
  OAI21_X1 U8015 ( .B1(n6417), .B2(n6416), .A(n6415), .ZN(n6418) );
  NAND2_X1 U8016 ( .A1(n6418), .A2(n8595), .ZN(n6421) );
  INV_X1 U8017 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9954) );
  NOR2_X1 U8018 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9954), .ZN(n9538) );
  OAI22_X1 U8019 ( .A1(n6538), .A2(n8615), .B1(n8599), .B2(n6482), .ZN(n6419)
         );
  AOI211_X1 U8020 ( .C1(n6560), .C2(n8617), .A(n9538), .B(n6419), .ZN(n6420)
         );
  OAI211_X1 U8021 ( .C1(n8588), .C2(n6491), .A(n6421), .B(n6420), .ZN(P1_U3228) );
  INV_X1 U8022 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6434) );
  OAI21_X1 U8023 ( .B1(n6427), .B2(P1_REG1_REG_10__SCAN_IN), .A(n6422), .ZN(
        n6424) );
  INV_X1 U8024 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7008) );
  AOI22_X1 U8025 ( .A1(n6608), .A2(P1_REG1_REG_11__SCAN_IN), .B1(n7008), .B2(
        n6429), .ZN(n6423) );
  NAND2_X1 U8026 ( .A1(n6423), .A2(n6424), .ZN(n6604) );
  OAI21_X1 U8027 ( .B1(n6424), .B2(n6423), .A(n6604), .ZN(n6425) );
  NAND2_X1 U8028 ( .A1(n6425), .A2(n9635), .ZN(n6433) );
  NOR2_X1 U8029 ( .A1(n6608), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6426) );
  AOI21_X1 U8030 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6608), .A(n6426), .ZN(
        n6428) );
  OAI21_X1 U8031 ( .B1(n6428), .B2(n4370), .A(n6607), .ZN(n6431) );
  NOR2_X1 U8032 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5276), .ZN(n6865) );
  NOR2_X1 U8033 ( .A1(n9543), .A2(n6429), .ZN(n6430) );
  AOI211_X1 U8034 ( .C1(n9616), .C2(n6431), .A(n6865), .B(n6430), .ZN(n6432)
         );
  OAI211_X1 U8035 ( .C1(n9621), .C2(n6434), .A(n6433), .B(n6432), .ZN(P1_U3252) );
  XNOR2_X2 U8036 ( .A(n6435), .B(n8891), .ZN(n6437) );
  AND2_X1 U8037 ( .A1(n8892), .A2(n4297), .ZN(n6438) );
  NAND2_X1 U8038 ( .A1(n6437), .A2(n6438), .ZN(n6455) );
  OAI21_X1 U8039 ( .B1(n6437), .B2(n6438), .A(n6455), .ZN(n9664) );
  INV_X1 U8040 ( .A(n9664), .ZN(n9667) );
  AOI21_X1 U8041 ( .B1(n5654), .B2(n6439), .A(n4797), .ZN(n6440) );
  NAND2_X1 U8042 ( .A1(n6441), .A2(n6440), .ZN(n9398) );
  NAND2_X1 U8043 ( .A1(n6442), .A2(n4797), .ZN(n6469) );
  NAND2_X1 U8044 ( .A1(n9398), .A2(n6469), .ZN(n9639) );
  NAND2_X1 U8045 ( .A1(n6435), .A2(n6443), .ZN(n6527) );
  OAI211_X1 U8046 ( .C1(n6443), .C2(n6435), .A(n9409), .B(n6527), .ZN(n9662)
         );
  INV_X1 U8047 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6444) );
  OAI22_X1 U8048 ( .A1(n9662), .A2(n4797), .B1(n9644), .B2(n6444), .ZN(n6450)
         );
  INV_X1 U8049 ( .A(n8892), .ZN(n6449) );
  XNOR2_X1 U8050 ( .A(n6437), .B(n6461), .ZN(n6448) );
  NAND2_X1 U8051 ( .A1(n5046), .A2(n4797), .ZN(n6447) );
  OR2_X1 U8052 ( .A1(n8830), .A2(n6837), .ZN(n6446) );
  OAI222_X1 U8053 ( .A1(n9392), .A2(n6449), .B1(n9394), .B2(n6456), .C1(n6448), 
        .C2(n9208), .ZN(n9665) );
  AOI211_X1 U8054 ( .C1(n9667), .C2(n9639), .A(n6450), .B(n9665), .ZN(n6452)
         );
  INV_X1 U8055 ( .A(n9217), .ZN(n9406) );
  AOI22_X1 U8056 ( .A1(n9406), .A2(n6453), .B1(n9405), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6451) );
  OAI21_X1 U8057 ( .B1(n6452), .B2(n9405), .A(n6451), .ZN(P1_U3290) );
  INV_X1 U8058 ( .A(n9398), .ZN(n9668) );
  NAND2_X1 U8059 ( .A1(n8891), .A2(n6453), .ZN(n6454) );
  NAND2_X1 U8060 ( .A1(n6455), .A2(n6454), .ZN(n6520) );
  INV_X1 U8061 ( .A(n6520), .ZN(n6458) );
  NAND2_X1 U8062 ( .A1(n6458), .A2(n8752), .ZN(n6521) );
  INV_X1 U8063 ( .A(n6457), .ZN(n6596) );
  NAND2_X1 U8064 ( .A1(n6456), .A2(n6596), .ZN(n6459) );
  NAND2_X1 U8065 ( .A1(n6521), .A2(n6459), .ZN(n6460) );
  INV_X1 U8066 ( .A(n6482), .ZN(n8888) );
  NAND2_X1 U8067 ( .A1(n6478), .A2(n8888), .ZN(n8750) );
  NAND2_X1 U8068 ( .A1(n6482), .A2(n6498), .ZN(n8754) );
  NAND2_X1 U8069 ( .A1(n6460), .A2(n6483), .ZN(n6480) );
  OAI21_X1 U8070 ( .B1(n6460), .B2(n6483), .A(n6480), .ZN(n6497) );
  OAI22_X1 U8071 ( .A1(n6456), .A2(n9392), .B1(n6574), .B2(n9394), .ZN(n6468)
         );
  INV_X1 U8072 ( .A(n6437), .ZN(n6462) );
  NAND2_X1 U8073 ( .A1(n6462), .A2(n6461), .ZN(n6464) );
  NAND2_X1 U8074 ( .A1(n8838), .A2(n6453), .ZN(n6463) );
  NAND2_X1 U8075 ( .A1(n8842), .A2(n6523), .ZN(n6465) );
  NAND2_X1 U8076 ( .A1(n6456), .A2(n6457), .ZN(n8839) );
  NAND2_X1 U8077 ( .A1(n6465), .A2(n8839), .ZN(n6485) );
  XNOR2_X1 U8078 ( .A(n6485), .B(n6483), .ZN(n6466) );
  NOR2_X1 U8079 ( .A1(n6466), .A2(n9208), .ZN(n6467) );
  AOI211_X1 U8080 ( .C1(n9668), .C2(n6497), .A(n6468), .B(n6467), .ZN(n6501)
         );
  INV_X1 U8081 ( .A(n6469), .ZN(n6470) );
  NAND2_X1 U8082 ( .A1(n9653), .A2(n6470), .ZN(n7333) );
  INV_X1 U8083 ( .A(n7333), .ZN(n9413) );
  INV_X1 U8084 ( .A(n6529), .ZN(n6472) );
  INV_X1 U8085 ( .A(n6490), .ZN(n6471) );
  AOI21_X1 U8086 ( .B1(n6498), .B2(n6472), .A(n6471), .ZN(n6499) );
  NAND2_X1 U8087 ( .A1(n6499), .A2(n9237), .ZN(n6475) );
  AOI22_X1 U8088 ( .A1(n9405), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9404), .B2(
        n6473), .ZN(n6474) );
  OAI211_X1 U8089 ( .C1(n6478), .C2(n9217), .A(n6475), .B(n6474), .ZN(n6476)
         );
  AOI21_X1 U8090 ( .B1(n9413), .B2(n6497), .A(n6476), .ZN(n6477) );
  OAI21_X1 U8091 ( .B1(n6501), .B2(n9405), .A(n6477), .ZN(P1_U3288) );
  NAND2_X1 U8092 ( .A1(n6482), .A2(n6478), .ZN(n6479) );
  NAND2_X1 U8093 ( .A1(n6480), .A2(n6479), .ZN(n6481) );
  NAND2_X1 U8094 ( .A1(n6574), .A2(n6560), .ZN(n8656) );
  INV_X1 U8095 ( .A(n6560), .ZN(n6535) );
  INV_X1 U8096 ( .A(n6574), .ZN(n8887) );
  NAND2_X1 U8097 ( .A1(n6535), .A2(n8887), .ZN(n8751) );
  NAND2_X1 U8098 ( .A1(n8656), .A2(n8751), .ZN(n6486) );
  NAND2_X1 U8099 ( .A1(n6481), .A2(n6486), .ZN(n6537) );
  OAI21_X1 U8100 ( .B1(n6481), .B2(n6486), .A(n6537), .ZN(n6559) );
  OAI22_X1 U8101 ( .A1(n6538), .A2(n9394), .B1(n6482), .B2(n9392), .ZN(n6489)
         );
  INV_X1 U8102 ( .A(n6483), .ZN(n6484) );
  XNOR2_X1 U8103 ( .A(n6486), .B(n8654), .ZN(n6487) );
  NOR2_X1 U8104 ( .A1(n6487), .A2(n9208), .ZN(n6488) );
  AOI211_X1 U8105 ( .C1(n9668), .C2(n6559), .A(n6489), .B(n6488), .ZN(n6563)
         );
  AOI21_X1 U8106 ( .B1(n6560), .B2(n6490), .A(n4463), .ZN(n6561) );
  NOR2_X1 U8107 ( .A1(n9217), .A2(n6535), .ZN(n6494) );
  INV_X1 U8108 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6492) );
  OAI22_X1 U8109 ( .A1(n9653), .A2(n6492), .B1(n6491), .B2(n9644), .ZN(n6493)
         );
  AOI211_X1 U8110 ( .C1(n6561), .C2(n9237), .A(n6494), .B(n6493), .ZN(n6496)
         );
  NAND2_X1 U8111 ( .A1(n6559), .A2(n9413), .ZN(n6495) );
  OAI211_X1 U8112 ( .C1(n6563), .C2(n9405), .A(n6496), .B(n6495), .ZN(P1_U3287) );
  INV_X1 U8113 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6504) );
  INV_X1 U8114 ( .A(n6497), .ZN(n6502) );
  AOI22_X1 U8115 ( .A1(n6499), .A2(n9409), .B1(n9330), .B2(n6498), .ZN(n6500)
         );
  OAI211_X1 U8116 ( .C1(n6502), .C2(n9663), .A(n6501), .B(n6500), .ZN(n6505)
         );
  NAND2_X1 U8117 ( .A1(n6505), .A2(n9352), .ZN(n6503) );
  OAI21_X1 U8118 ( .B1(n9352), .B2(n6504), .A(n6503), .ZN(P1_U3463) );
  INV_X1 U8119 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6507) );
  NAND2_X1 U8120 ( .A1(n6505), .A2(n9334), .ZN(n6506) );
  OAI21_X1 U8121 ( .B1(n9334), .B2(n6507), .A(n6506), .ZN(P1_U3526) );
  INV_X1 U8122 ( .A(n6508), .ZN(n6555) );
  AOI22_X1 U8123 ( .A1(n8107), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8491), .ZN(n6509) );
  OAI21_X1 U8124 ( .B1(n6555), .B2(n7626), .A(n6509), .ZN(P2_U3342) );
  INV_X1 U8125 ( .A(n6510), .ZN(n6512) );
  OAI222_X1 U8126 ( .A1(n9360), .A2(n6511), .B1(n9364), .B2(n6512), .C1(
        P1_U3084), .C2(n8900), .ZN(P1_U3338) );
  INV_X1 U8127 ( .A(n8091), .ZN(n8082) );
  OAI222_X1 U8128 ( .A1(n7628), .A2(n9921), .B1(n7626), .B2(n6512), .C1(
        P2_U3152), .C2(n8082), .ZN(P2_U3343) );
  NAND2_X1 U8129 ( .A1(n6513), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8002) );
  NAND2_X1 U8130 ( .A1(n7999), .A2(n8002), .ZN(n6515) );
  NAND2_X1 U8131 ( .A1(n6515), .A2(n6514), .ZN(n6518) );
  OR2_X1 U8132 ( .A1(n7999), .A2(n6516), .ZN(n6517) );
  NOR2_X1 U8133 ( .A1(n9697), .A2(P2_U3966), .ZN(P2_U3151) );
  NAND2_X1 U8134 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8026), .ZN(n6519) );
  OAI21_X1 U8135 ( .B1(n8168), .B2(n8026), .A(n6519), .ZN(P2_U3581) );
  INV_X1 U8136 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6532) );
  INV_X1 U8137 ( .A(n6521), .ZN(n6522) );
  AOI21_X1 U8138 ( .B1(n6523), .B2(n6520), .A(n6522), .ZN(n6597) );
  XNOR2_X1 U8139 ( .A(n8842), .B(n6523), .ZN(n6526) );
  AOI22_X1 U8140 ( .A1(n8888), .A2(n9232), .B1(n9231), .B2(n8891), .ZN(n6524)
         );
  OAI21_X1 U8141 ( .B1(n6597), .B2(n9398), .A(n6524), .ZN(n6525) );
  AOI21_X1 U8142 ( .B1(n9401), .B2(n6526), .A(n6525), .ZN(n6602) );
  AND2_X1 U8143 ( .A1(n6527), .A2(n6457), .ZN(n6528) );
  NOR2_X1 U8144 ( .A1(n6529), .A2(n6528), .ZN(n6600) );
  AOI22_X1 U8145 ( .A1(n6600), .A2(n9409), .B1(n9330), .B2(n6457), .ZN(n6530)
         );
  OAI211_X1 U8146 ( .C1(n6597), .C2(n9663), .A(n6602), .B(n6530), .ZN(n6533)
         );
  NAND2_X1 U8147 ( .A1(n6533), .A2(n9352), .ZN(n6531) );
  OAI21_X1 U8148 ( .B1(n9352), .B2(n6532), .A(n6531), .ZN(P1_U3460) );
  NAND2_X1 U8149 ( .A1(n6533), .A2(n9334), .ZN(n6534) );
  OAI21_X1 U8150 ( .B1(n9334), .B2(n6299), .A(n6534), .ZN(P1_U3525) );
  INV_X1 U8151 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6551) );
  NAND2_X1 U8152 ( .A1(n6574), .A2(n6535), .ZN(n6536) );
  NAND2_X1 U8153 ( .A1(n6537), .A2(n6536), .ZN(n6541) );
  NAND2_X1 U8154 ( .A1(n6538), .A2(n9641), .ZN(n6646) );
  INV_X1 U8155 ( .A(n9641), .ZN(n6539) );
  INV_X1 U8156 ( .A(n6538), .ZN(n8886) );
  NAND2_X1 U8157 ( .A1(n6539), .A2(n8886), .ZN(n6648) );
  AND2_X1 U8158 ( .A1(n6646), .A2(n6648), .ZN(n6543) );
  NAND2_X1 U8159 ( .A1(n6541), .A2(n6543), .ZN(n6542) );
  NAND2_X1 U8160 ( .A1(n6579), .A2(n6542), .ZN(n9651) );
  NAND2_X1 U8161 ( .A1(n9398), .A2(n9663), .ZN(n9482) );
  XNOR2_X1 U8162 ( .A(n6647), .B(n6540), .ZN(n6546) );
  NAND2_X1 U8163 ( .A1(n8885), .A2(n9232), .ZN(n6544) );
  OAI21_X1 U8164 ( .B1(n6574), .B2(n9392), .A(n6544), .ZN(n6545) );
  AOI21_X1 U8165 ( .B1(n6546), .B2(n9401), .A(n6545), .ZN(n9649) );
  INV_X1 U8166 ( .A(n9409), .ZN(n9242) );
  AOI21_X1 U8167 ( .B1(n6547), .B2(n9641), .A(n9242), .ZN(n6548) );
  AND2_X1 U8168 ( .A1(n6548), .A2(n6587), .ZN(n9647) );
  AOI21_X1 U8169 ( .B1(n9330), .B2(n9641), .A(n9647), .ZN(n6549) );
  OAI211_X1 U8170 ( .C1(n9651), .C2(n9332), .A(n9649), .B(n6549), .ZN(n6552)
         );
  NAND2_X1 U8171 ( .A1(n6552), .A2(n9352), .ZN(n6550) );
  OAI21_X1 U8172 ( .B1(n9352), .B2(n6551), .A(n6550), .ZN(P1_U3469) );
  INV_X1 U8173 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U8174 ( .A1(n6552), .A2(n9334), .ZN(n6553) );
  OAI21_X1 U8175 ( .B1(n9334), .B2(n6554), .A(n6553), .ZN(P1_U3528) );
  INV_X1 U8176 ( .A(n8919), .ZN(n8907) );
  OAI222_X1 U8177 ( .A1(n9360), .A2(n6556), .B1(n8907), .B2(P1_U3084), .C1(
        n9364), .C2(n6555), .ZN(P1_U3337) );
  INV_X1 U8178 ( .A(n6557), .ZN(n6593) );
  AOI22_X1 U8179 ( .A1(n8930), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9357), .ZN(n6558) );
  OAI21_X1 U8180 ( .B1(n6593), .B2(n9364), .A(n6558), .ZN(P1_U3336) );
  INV_X1 U8181 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6566) );
  INV_X1 U8182 ( .A(n6559), .ZN(n6564) );
  AOI22_X1 U8183 ( .A1(n6561), .A2(n9409), .B1(n9330), .B2(n6560), .ZN(n6562)
         );
  OAI211_X1 U8184 ( .C1(n6564), .C2(n9663), .A(n6563), .B(n6562), .ZN(n6567)
         );
  NAND2_X1 U8185 ( .A1(n6567), .A2(n9334), .ZN(n6565) );
  OAI21_X1 U8186 ( .B1(n9334), .B2(n6566), .A(n6565), .ZN(P1_U3527) );
  INV_X1 U8187 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6569) );
  NAND2_X1 U8188 ( .A1(n6567), .A2(n9352), .ZN(n6568) );
  OAI21_X1 U8189 ( .B1(n9352), .B2(n6569), .A(n6568), .ZN(P1_U3466) );
  INV_X1 U8190 ( .A(n6570), .ZN(n9643) );
  CLKBUF_X1 U8191 ( .A(n6571), .Z(n6632) );
  OAI21_X1 U8192 ( .B1(n6572), .B2(n4374), .A(n6632), .ZN(n6573) );
  NAND2_X1 U8193 ( .A1(n6573), .A2(n8595), .ZN(n6577) );
  AND2_X1 U8194 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9554) );
  INV_X1 U8195 ( .A(n8885), .ZN(n6655) );
  OAI22_X1 U8196 ( .A1(n6655), .A2(n8615), .B1(n8599), .B2(n6574), .ZN(n6575)
         );
  AOI211_X1 U8197 ( .C1(n9641), .C2(n8617), .A(n9554), .B(n6575), .ZN(n6576)
         );
  OAI211_X1 U8198 ( .C1(n8588), .C2(n9643), .A(n6577), .B(n6576), .ZN(P1_U3225) );
  NAND2_X1 U8199 ( .A1(n8886), .A2(n9641), .ZN(n6578) );
  NAND2_X1 U8200 ( .A1(n6641), .A2(n8885), .ZN(n8661) );
  NAND2_X1 U8201 ( .A1(n6655), .A2(n6634), .ZN(n6649) );
  NAND2_X1 U8202 ( .A1(n8661), .A2(n6649), .ZN(n6582) );
  OAI21_X1 U8203 ( .B1(n6580), .B2(n6582), .A(n6643), .ZN(n6617) );
  INV_X1 U8204 ( .A(n8653), .ZN(n6581) );
  NAND2_X1 U8205 ( .A1(n8751), .A2(n6648), .ZN(n8659) );
  OAI21_X1 U8206 ( .B1(n6581), .B2(n8659), .A(n6646), .ZN(n6583) );
  XNOR2_X1 U8207 ( .A(n6583), .B(n6582), .ZN(n6585) );
  INV_X1 U8208 ( .A(n6839), .ZN(n8884) );
  AOI22_X1 U8209 ( .A1(n9232), .A2(n8884), .B1(n8886), .B2(n9231), .ZN(n6584)
         );
  OAI21_X1 U8210 ( .B1(n6585), .B2(n9208), .A(n6584), .ZN(n6586) );
  AOI21_X1 U8211 ( .B1(n6617), .B2(n9668), .A(n6586), .ZN(n6620) );
  AOI21_X1 U8212 ( .B1(n6634), .B2(n6587), .A(n6656), .ZN(n6618) );
  NAND2_X1 U8213 ( .A1(n6618), .A2(n9237), .ZN(n6589) );
  AOI22_X1 U8214 ( .A1(n9405), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n6637), .B2(
        n9404), .ZN(n6588) );
  OAI211_X1 U8215 ( .C1(n6641), .C2(n9217), .A(n6589), .B(n6588), .ZN(n6590)
         );
  AOI21_X1 U8216 ( .B1(n6617), .B2(n9413), .A(n6590), .ZN(n6591) );
  OAI21_X1 U8217 ( .B1(n6620), .B2(n9405), .A(n6591), .ZN(P1_U3285) );
  INV_X2 U8218 ( .A(P1_U4006), .ZN(n8890) );
  NAND2_X1 U8219 ( .A1(n8890), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6592) );
  OAI21_X1 U8220 ( .B1(n9023), .B2(n8890), .A(n6592), .ZN(P1_U3584) );
  INV_X1 U8221 ( .A(n8122), .ZN(n8118) );
  OAI222_X1 U8222 ( .A1(n7628), .A2(n6594), .B1(n7626), .B2(n6593), .C1(n8118), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  AOI22_X1 U8223 ( .A1(n9404), .A2(P1_REG3_REG_2__SCAN_IN), .B1(
        P1_REG2_REG_2__SCAN_IN), .B2(n9405), .ZN(n6595) );
  OAI21_X1 U8224 ( .B1(n9217), .B2(n6596), .A(n6595), .ZN(n6599) );
  NOR2_X1 U8225 ( .A1(n6597), .A2(n7333), .ZN(n6598) );
  AOI211_X1 U8226 ( .C1(n6600), .C2(n9237), .A(n6599), .B(n6598), .ZN(n6601)
         );
  OAI21_X1 U8227 ( .B1(n9405), .B2(n6602), .A(n6601), .ZN(P1_U3289) );
  INV_X1 U8228 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6616) );
  INV_X1 U8229 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6603) );
  MUX2_X1 U8230 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6603), .S(n6688), .Z(n6606)
         );
  OAI21_X1 U8231 ( .B1(n6608), .B2(P1_REG1_REG_11__SCAN_IN), .A(n6604), .ZN(
        n6605) );
  NAND2_X1 U8232 ( .A1(n6606), .A2(n6605), .ZN(n6683) );
  OAI21_X1 U8233 ( .B1(n6606), .B2(n6605), .A(n6683), .ZN(n6613) );
  OAI21_X1 U8234 ( .B1(n6608), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6607), .ZN(
        n6611) );
  NAND2_X1 U8235 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6688), .ZN(n6609) );
  OAI21_X1 U8236 ( .B1(n6688), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6609), .ZN(
        n6610) );
  NOR2_X1 U8237 ( .A1(n6610), .A2(n6611), .ZN(n6687) );
  AOI211_X1 U8238 ( .C1(n6611), .C2(n6610), .A(n6687), .B(n9623), .ZN(n6612)
         );
  AOI21_X1 U8239 ( .B1(n9635), .B2(n6613), .A(n6612), .ZN(n6615) );
  AND2_X1 U8240 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6909) );
  AOI21_X1 U8241 ( .B1(n9629), .B2(n6688), .A(n6909), .ZN(n6614) );
  OAI211_X1 U8242 ( .C1(n9621), .C2(n6616), .A(n6615), .B(n6614), .ZN(P1_U3253) );
  INV_X1 U8243 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6623) );
  INV_X1 U8244 ( .A(n6617), .ZN(n6621) );
  AOI22_X1 U8245 ( .A1(n6618), .A2(n9409), .B1(n9330), .B2(n6634), .ZN(n6619)
         );
  OAI211_X1 U8246 ( .C1(n6621), .C2(n9663), .A(n6620), .B(n6619), .ZN(n6624)
         );
  NAND2_X1 U8247 ( .A1(n6624), .A2(n9334), .ZN(n6622) );
  OAI21_X1 U8248 ( .B1(n9334), .B2(n6623), .A(n6622), .ZN(P1_U3529) );
  INV_X1 U8249 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6626) );
  NAND2_X1 U8250 ( .A1(n6624), .A2(n9352), .ZN(n6625) );
  OAI21_X1 U8251 ( .B1(n9352), .B2(n6626), .A(n6625), .ZN(P1_U3472) );
  INV_X1 U8252 ( .A(n6627), .ZN(n6629) );
  NOR2_X1 U8253 ( .A1(n6629), .A2(n6628), .ZN(n6633) );
  INV_X1 U8254 ( .A(n6630), .ZN(n6631) );
  AOI21_X1 U8255 ( .B1(n6633), .B2(n6632), .A(n6631), .ZN(n6640) );
  AOI22_X1 U8256 ( .A1(n6634), .A2(n8617), .B1(n8611), .B2(n8886), .ZN(n6639)
         );
  INV_X1 U8257 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6635) );
  NOR2_X1 U8258 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6635), .ZN(n9566) );
  NOR2_X1 U8259 ( .A1(n8615), .A2(n6839), .ZN(n6636) );
  AOI211_X1 U8260 ( .C1(n6637), .C2(n8612), .A(n9566), .B(n6636), .ZN(n6638)
         );
  OAI211_X1 U8261 ( .C1(n6640), .C2(n8619), .A(n6639), .B(n6638), .ZN(P1_U3237) );
  NAND2_X1 U8262 ( .A1(n6641), .A2(n6655), .ZN(n6642) );
  NAND2_X1 U8263 ( .A1(n6643), .A2(n6642), .ZN(n6644) );
  OR2_X1 U8264 ( .A1(n6840), .A2(n6839), .ZN(n8665) );
  NAND2_X1 U8265 ( .A1(n6840), .A2(n6839), .ZN(n8819) );
  NAND2_X1 U8266 ( .A1(n8665), .A2(n8819), .ZN(n8755) );
  NAND2_X1 U8267 ( .A1(n6644), .A2(n8755), .ZN(n6842) );
  OAI21_X1 U8268 ( .B1(n6644), .B2(n8755), .A(n6842), .ZN(n6645) );
  INV_X1 U8269 ( .A(n6645), .ZN(n6810) );
  AND2_X1 U8270 ( .A1(n6649), .A2(n6646), .ZN(n8660) );
  NAND2_X1 U8271 ( .A1(n6647), .A2(n8660), .ZN(n6651) );
  NAND2_X1 U8272 ( .A1(n8661), .A2(n6648), .ZN(n6650) );
  NAND2_X1 U8273 ( .A1(n6650), .A2(n6649), .ZN(n8812) );
  NAND2_X1 U8274 ( .A1(n6651), .A2(n8812), .ZN(n6653) );
  INV_X1 U8275 ( .A(n6838), .ZN(n6652) );
  AOI21_X1 U8276 ( .B1(n8755), .B2(n6653), .A(n6652), .ZN(n6654) );
  OAI222_X1 U8277 ( .A1(n9392), .A2(n6655), .B1(n9394), .B2(n6926), .C1(n9208), 
        .C2(n6654), .ZN(n6807) );
  INV_X1 U8278 ( .A(n6840), .ZN(n6664) );
  INV_X1 U8279 ( .A(n6656), .ZN(n6658) );
  INV_X1 U8280 ( .A(n6852), .ZN(n6657) );
  AOI211_X1 U8281 ( .C1(n6840), .C2(n6658), .A(n9242), .B(n6657), .ZN(n6808)
         );
  NOR2_X1 U8282 ( .A1(n6659), .A2(n4797), .ZN(n9412) );
  NAND2_X1 U8283 ( .A1(n6808), .A2(n9412), .ZN(n6663) );
  NOR2_X1 U8284 ( .A1(n9644), .A2(n6660), .ZN(n6661) );
  AOI21_X1 U8285 ( .B1(n9405), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6661), .ZN(
        n6662) );
  OAI211_X1 U8286 ( .C1(n6664), .C2(n9217), .A(n6663), .B(n6662), .ZN(n6665)
         );
  AOI21_X1 U8287 ( .B1(n6807), .B2(n9653), .A(n6665), .ZN(n6666) );
  OAI21_X1 U8288 ( .B1(n6810), .B2(n9239), .A(n6666), .ZN(P1_U3284) );
  OAI21_X1 U8289 ( .B1(n6669), .B2(n6668), .A(n6667), .ZN(n6676) );
  INV_X1 U8290 ( .A(n6926), .ZN(n8883) );
  NOR2_X1 U8291 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5198), .ZN(n9570) );
  AOI21_X1 U8292 ( .B1(n8578), .B2(n8883), .A(n9570), .ZN(n6674) );
  NAND2_X1 U8293 ( .A1(n8617), .A2(n6840), .ZN(n6673) );
  NAND2_X1 U8294 ( .A1(n8612), .A2(n6670), .ZN(n6672) );
  NAND2_X1 U8295 ( .A1(n8611), .A2(n8885), .ZN(n6671) );
  NAND4_X1 U8296 ( .A1(n6674), .A2(n6673), .A3(n6672), .A4(n6671), .ZN(n6675)
         );
  AOI21_X1 U8297 ( .B1(n6676), .B2(n8595), .A(n6675), .ZN(n6677) );
  INV_X1 U8298 ( .A(n6677), .ZN(P1_U3211) );
  INV_X1 U8299 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6679) );
  INV_X1 U8300 ( .A(n6678), .ZN(n6680) );
  INV_X1 U8301 ( .A(n9630), .ZN(n8928) );
  OAI222_X1 U8302 ( .A1(n9360), .A2(n6679), .B1(n9364), .B2(n6680), .C1(
        P1_U3084), .C2(n8928), .ZN(P1_U3335) );
  INV_X1 U8303 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6681) );
  INV_X1 U8304 ( .A(n8138), .ZN(n8128) );
  OAI222_X1 U8305 ( .A1(n7628), .A2(n6681), .B1(n7626), .B2(n6680), .C1(
        P2_U3152), .C2(n8128), .ZN(P2_U3340) );
  INV_X1 U8306 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6696) );
  INV_X1 U8307 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6682) );
  MUX2_X1 U8308 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6682), .S(n7145), .Z(n6686)
         );
  OR2_X1 U8309 ( .A1(n6688), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6684) );
  NAND2_X1 U8310 ( .A1(n6684), .A2(n6683), .ZN(n6685) );
  NAND2_X1 U8311 ( .A1(n6686), .A2(n6685), .ZN(n7144) );
  OAI21_X1 U8312 ( .B1(n6686), .B2(n6685), .A(n7144), .ZN(n6693) );
  INV_X1 U8313 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6689) );
  MUX2_X1 U8314 ( .A(n6689), .B(P1_REG2_REG_13__SCAN_IN), .S(n7145), .Z(n6690)
         );
  AOI211_X1 U8315 ( .C1(n6691), .C2(n6690), .A(n7138), .B(n9623), .ZN(n6692)
         );
  AOI21_X1 U8316 ( .B1(n9635), .B2(n6693), .A(n6692), .ZN(n6695) );
  AND2_X1 U8317 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6988) );
  AOI21_X1 U8318 ( .B1(n9629), .B2(n7145), .A(n6988), .ZN(n6694) );
  OAI211_X1 U8319 ( .C1(n9621), .C2(n6696), .A(n6695), .B(n6694), .ZN(P1_U3254) );
  NOR2_X1 U8320 ( .A1(n6229), .A2(P2_U3152), .ZN(n7513) );
  INV_X1 U8321 ( .A(n8002), .ZN(n7032) );
  AOI21_X1 U8322 ( .B1(n6697), .B2(n7513), .A(n7032), .ZN(n6698) );
  OAI21_X1 U8323 ( .B1(n7999), .B2(n6699), .A(n6698), .ZN(n6701) );
  AND2_X1 U8324 ( .A1(n6701), .A2(n6700), .ZN(n6716) );
  INV_X1 U8325 ( .A(n6716), .ZN(n6702) );
  NAND2_X1 U8326 ( .A1(n6702), .A2(n8026), .ZN(n6751) );
  NOR2_X1 U8327 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6703), .ZN(n6720) );
  INV_X1 U8328 ( .A(n6741), .ZN(n9381) );
  NAND2_X1 U8329 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9368) );
  NAND2_X1 U8330 ( .A1(n9370), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6704) );
  AOI21_X1 U8331 ( .B1(n9370), .B2(P2_REG1_REG_1__SCAN_IN), .A(n9366), .ZN(
        n9379) );
  INV_X1 U8332 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6705) );
  MUX2_X1 U8333 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6705), .S(n6741), .Z(n9378)
         );
  NOR2_X1 U8334 ( .A1(n9379), .A2(n9378), .ZN(n9377) );
  AOI21_X1 U8335 ( .B1(n9381), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9377), .ZN(
        n8035) );
  OR2_X1 U8336 ( .A1(n6735), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6707) );
  NAND2_X1 U8337 ( .A1(n6735), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6706) );
  NAND2_X1 U8338 ( .A1(n6707), .A2(n6706), .ZN(n8034) );
  NOR2_X1 U8339 ( .A1(n8035), .A2(n8034), .ZN(n8033) );
  OR2_X1 U8340 ( .A1(n6734), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6709) );
  NAND2_X1 U8341 ( .A1(n6734), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U8342 ( .A1(n6709), .A2(n6708), .ZN(n8049) );
  OR2_X1 U8343 ( .A1(n6732), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6711) );
  NAND2_X1 U8344 ( .A1(n6732), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6710) );
  NAND2_X1 U8345 ( .A1(n6711), .A2(n6710), .ZN(n8063) );
  AOI21_X1 U8346 ( .B1(n6732), .B2(P2_REG1_REG_5__SCAN_IN), .A(n8061), .ZN(
        n6794) );
  NAND2_X1 U8347 ( .A1(n6729), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6712) );
  OAI21_X1 U8348 ( .B1(n6729), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6712), .ZN(
        n6793) );
  NOR2_X1 U8349 ( .A1(n6794), .A2(n6793), .ZN(n6792) );
  AOI21_X1 U8350 ( .B1(n6729), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6792), .ZN(
        n6762) );
  NAND2_X1 U8351 ( .A1(n6727), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6713) );
  OAI21_X1 U8352 ( .B1(n6727), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6713), .ZN(
        n6761) );
  INV_X1 U8353 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6714) );
  MUX2_X1 U8354 ( .A(n6714), .B(P2_REG1_REG_8__SCAN_IN), .S(n6724), .Z(n6772)
         );
  MUX2_X1 U8355 ( .A(n4520), .B(P2_REG1_REG_9__SCAN_IN), .S(n6721), .Z(n6783)
         );
  NOR2_X1 U8356 ( .A1(n6784), .A2(n6783), .ZN(n6782) );
  INV_X1 U8357 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6715) );
  MUX2_X1 U8358 ( .A(n6715), .B(P2_REG1_REG_10__SCAN_IN), .S(n6825), .Z(n6717)
         );
  AOI211_X1 U8359 ( .C1(n6718), .C2(n6717), .A(n6824), .B(n9700), .ZN(n6719)
         );
  AOI211_X1 U8360 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n9697), .A(n6720), .B(
        n6719), .ZN(n6757) );
  NAND2_X1 U8361 ( .A1(n6721), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6748) );
  INV_X1 U8362 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6722) );
  MUX2_X1 U8363 ( .A(n6722), .B(P2_REG2_REG_9__SCAN_IN), .S(n6721), .Z(n6723)
         );
  INV_X1 U8364 ( .A(n6723), .ZN(n6788) );
  NAND2_X1 U8365 ( .A1(n6724), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6747) );
  INV_X1 U8366 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6725) );
  MUX2_X1 U8367 ( .A(n6725), .B(P2_REG2_REG_8__SCAN_IN), .S(n6724), .Z(n6726)
         );
  INV_X1 U8368 ( .A(n6726), .ZN(n6777) );
  NAND2_X1 U8369 ( .A1(n6727), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6746) );
  INV_X1 U8370 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6728) );
  MUX2_X1 U8371 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6728), .S(n6727), .Z(n6766)
         );
  NAND2_X1 U8372 ( .A1(n6729), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6745) );
  INV_X1 U8373 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6730) );
  MUX2_X1 U8374 ( .A(n6730), .B(P2_REG2_REG_6__SCAN_IN), .S(n6729), .Z(n6731)
         );
  INV_X1 U8375 ( .A(n6731), .ZN(n6798) );
  NAND2_X1 U8376 ( .A1(n6732), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6744) );
  INV_X1 U8377 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6733) );
  MUX2_X1 U8378 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n6733), .S(n6732), .Z(n8056)
         );
  NAND2_X1 U8379 ( .A1(n6734), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6743) );
  INV_X1 U8380 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9993) );
  MUX2_X1 U8381 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9993), .S(n6734), .Z(n8042)
         );
  NAND2_X1 U8382 ( .A1(n6735), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6742) );
  MUX2_X1 U8383 ( .A(n5780), .B(P2_REG2_REG_3__SCAN_IN), .S(n6735), .Z(n6736)
         );
  INV_X1 U8384 ( .A(n6736), .ZN(n8030) );
  INV_X1 U8385 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7301) );
  MUX2_X1 U8386 ( .A(n7301), .B(P2_REG2_REG_2__SCAN_IN), .S(n6741), .Z(n9384)
         );
  NAND2_X1 U8387 ( .A1(n9370), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6740) );
  INV_X1 U8388 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6738) );
  MUX2_X1 U8389 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6738), .S(n6737), .Z(n6739)
         );
  INV_X1 U8390 ( .A(n6739), .ZN(n9372) );
  NAND3_X1 U8391 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n9372), .ZN(n9371) );
  NAND2_X1 U8392 ( .A1(n6740), .A2(n9371), .ZN(n9385) );
  NAND2_X1 U8393 ( .A1(n9384), .A2(n9385), .ZN(n9383) );
  OAI21_X1 U8394 ( .B1(n6741), .B2(n7301), .A(n9383), .ZN(n8029) );
  NAND2_X1 U8395 ( .A1(n8030), .A2(n8029), .ZN(n8028) );
  NAND2_X1 U8396 ( .A1(n6742), .A2(n8028), .ZN(n8043) );
  NAND2_X1 U8397 ( .A1(n8042), .A2(n8043), .ZN(n8041) );
  NAND2_X1 U8398 ( .A1(n6743), .A2(n8041), .ZN(n8057) );
  NAND2_X1 U8399 ( .A1(n8056), .A2(n8057), .ZN(n8055) );
  NAND2_X1 U8400 ( .A1(n6744), .A2(n8055), .ZN(n6799) );
  NAND2_X1 U8401 ( .A1(n6798), .A2(n6799), .ZN(n6797) );
  NAND2_X1 U8402 ( .A1(n6745), .A2(n6797), .ZN(n6767) );
  NAND2_X1 U8403 ( .A1(n6766), .A2(n6767), .ZN(n6765) );
  NAND2_X1 U8404 ( .A1(n6746), .A2(n6765), .ZN(n6778) );
  NAND2_X1 U8405 ( .A1(n6777), .A2(n6778), .ZN(n6776) );
  NAND2_X1 U8406 ( .A1(n6747), .A2(n6776), .ZN(n6789) );
  NAND2_X1 U8407 ( .A1(n6788), .A2(n6789), .ZN(n6787) );
  NAND2_X1 U8408 ( .A1(n6748), .A2(n6787), .ZN(n6755) );
  INV_X1 U8409 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6749) );
  MUX2_X1 U8410 ( .A(n6749), .B(P2_REG2_REG_10__SCAN_IN), .S(n6825), .Z(n6750)
         );
  INV_X1 U8411 ( .A(n6750), .ZN(n6754) );
  INV_X1 U8412 ( .A(n7998), .ZN(n7569) );
  NAND2_X1 U8413 ( .A1(n6751), .A2(n7569), .ZN(n8142) );
  INV_X1 U8414 ( .A(n8142), .ZN(n6753) );
  NAND2_X1 U8415 ( .A1(n6754), .A2(n6755), .ZN(n6816) );
  OAI211_X1 U8416 ( .C1(n6755), .C2(n6754), .A(n9695), .B(n6816), .ZN(n6756)
         );
  OAI211_X1 U8417 ( .C1(n9699), .C2(n6758), .A(n6757), .B(n6756), .ZN(P2_U3255) );
  NOR2_X1 U8418 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6759), .ZN(n6764) );
  AOI211_X1 U8419 ( .C1(n6762), .C2(n6761), .A(n6760), .B(n9700), .ZN(n6763)
         );
  AOI211_X1 U8420 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n9697), .A(n6764), .B(
        n6763), .ZN(n6769) );
  OAI211_X1 U8421 ( .C1(n6767), .C2(n6766), .A(n9695), .B(n6765), .ZN(n6768)
         );
  OAI211_X1 U8422 ( .C1(n9699), .C2(n6770), .A(n6769), .B(n6768), .ZN(P2_U3252) );
  NAND2_X1 U8423 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n9685) );
  INV_X1 U8424 ( .A(n9685), .ZN(n6775) );
  AOI211_X1 U8425 ( .C1(n6773), .C2(n6772), .A(n6771), .B(n9700), .ZN(n6774)
         );
  AOI211_X1 U8426 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n9697), .A(n6775), .B(
        n6774), .ZN(n6780) );
  OAI211_X1 U8427 ( .C1(n6778), .C2(n6777), .A(n9695), .B(n6776), .ZN(n6779)
         );
  OAI211_X1 U8428 ( .C1(n9699), .C2(n6781), .A(n6780), .B(n6779), .ZN(P2_U3253) );
  NAND2_X1 U8429 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7127) );
  INV_X1 U8430 ( .A(n7127), .ZN(n6786) );
  AOI211_X1 U8431 ( .C1(n6784), .C2(n6783), .A(n6782), .B(n9700), .ZN(n6785)
         );
  AOI211_X1 U8432 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n9697), .A(n6786), .B(
        n6785), .ZN(n6791) );
  OAI211_X1 U8433 ( .C1(n6789), .C2(n6788), .A(n9695), .B(n6787), .ZN(n6790)
         );
  OAI211_X1 U8434 ( .C1(n9699), .C2(n4521), .A(n6791), .B(n6790), .ZN(P2_U3254) );
  NAND2_X1 U8435 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7105) );
  INV_X1 U8436 ( .A(n7105), .ZN(n6796) );
  AOI211_X1 U8437 ( .C1(n6794), .C2(n6793), .A(n6792), .B(n9700), .ZN(n6795)
         );
  AOI211_X1 U8438 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n9697), .A(n6796), .B(
        n6795), .ZN(n6801) );
  OAI211_X1 U8439 ( .C1(n6799), .C2(n6798), .A(n9695), .B(n6797), .ZN(n6800)
         );
  OAI211_X1 U8440 ( .C1(n9699), .C2(n6802), .A(n6801), .B(n6800), .ZN(P2_U3251) );
  INV_X1 U8441 ( .A(n6803), .ZN(n6805) );
  OAI222_X1 U8442 ( .A1(n7628), .A2(n6804), .B1(n7626), .B2(n6805), .C1(
        P2_U3152), .C2(n8395), .ZN(P2_U3339) );
  OAI222_X1 U8443 ( .A1(n9360), .A2(n6806), .B1(n9364), .B2(n6805), .C1(
        P1_U3084), .C2(n9646), .ZN(P1_U3334) );
  INV_X1 U8444 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6812) );
  AOI211_X1 U8445 ( .C1(n9330), .C2(n6840), .A(n6808), .B(n6807), .ZN(n6809)
         );
  OAI21_X1 U8446 ( .B1(n9332), .B2(n6810), .A(n6809), .ZN(n6813) );
  NAND2_X1 U8447 ( .A1(n6813), .A2(n9352), .ZN(n6811) );
  OAI21_X1 U8448 ( .B1(n9352), .B2(n6812), .A(n6811), .ZN(P1_U3475) );
  INV_X1 U8449 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6815) );
  NAND2_X1 U8450 ( .A1(n6813), .A2(n9334), .ZN(n6814) );
  OAI21_X1 U8451 ( .B1(n9334), .B2(n6815), .A(n6814), .ZN(P1_U3530) );
  NAND2_X1 U8452 ( .A1(n6825), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6817) );
  NAND2_X1 U8453 ( .A1(n6817), .A2(n6816), .ZN(n6821) );
  INV_X1 U8454 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6818) );
  MUX2_X1 U8455 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n6818), .S(n6878), .Z(n6819)
         );
  INV_X1 U8456 ( .A(n6819), .ZN(n6820) );
  NOR2_X1 U8457 ( .A1(n6821), .A2(n6820), .ZN(n6879) );
  AOI21_X1 U8458 ( .B1(n6821), .B2(n6820), .A(n6879), .ZN(n6834) );
  NOR2_X1 U8459 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7392), .ZN(n6822) );
  AOI21_X1 U8460 ( .B1(n9697), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6822), .ZN(
        n6830) );
  INV_X1 U8461 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6823) );
  MUX2_X1 U8462 ( .A(n6823), .B(P2_REG1_REG_11__SCAN_IN), .S(n6878), .Z(n6827)
         );
  AOI21_X1 U8463 ( .B1(n6827), .B2(n6826), .A(n6871), .ZN(n6828) );
  NAND2_X1 U8464 ( .A1(n9694), .A2(n6828), .ZN(n6829) );
  OAI211_X1 U8465 ( .C1(n9699), .C2(n6831), .A(n6830), .B(n6829), .ZN(n6832)
         );
  INV_X1 U8466 ( .A(n6832), .ZN(n6833) );
  OAI21_X1 U8467 ( .B1(n9698), .B2(n6834), .A(n6833), .ZN(P2_U3256) );
  INV_X1 U8468 ( .A(n6835), .ZN(n6859) );
  OAI222_X1 U8469 ( .A1(n9364), .A2(n6859), .B1(n6837), .B2(P1_U3084), .C1(
        n6836), .C2(n9360), .ZN(P1_U3333) );
  NAND2_X1 U8470 ( .A1(n6838), .A2(n8819), .ZN(n6924) );
  OR2_X1 U8471 ( .A1(n6970), .A2(n6926), .ZN(n8669) );
  NAND2_X1 U8472 ( .A1(n6970), .A2(n6926), .ZN(n8820) );
  XNOR2_X1 U8473 ( .A(n6924), .B(n8758), .ZN(n6848) );
  OAI22_X1 U8474 ( .A1(n9393), .A2(n9394), .B1(n6839), .B2(n9392), .ZN(n6847)
         );
  OR2_X1 U8475 ( .A1(n6840), .A2(n8884), .ZN(n6841) );
  NAND2_X1 U8476 ( .A1(n6842), .A2(n6841), .ZN(n6844) );
  NAND2_X1 U8477 ( .A1(n6844), .A2(n8758), .ZN(n6845) );
  NAND2_X1 U8478 ( .A1(n6928), .A2(n6845), .ZN(n6974) );
  NOR2_X1 U8479 ( .A1(n6974), .A2(n9398), .ZN(n6846) );
  AOI211_X1 U8480 ( .C1(n6848), .C2(n9401), .A(n6847), .B(n6846), .ZN(n6973)
         );
  INV_X1 U8481 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6850) );
  INV_X1 U8482 ( .A(n6894), .ZN(n6849) );
  OAI22_X1 U8483 ( .A1(n9653), .A2(n6850), .B1(n6849), .B2(n9644), .ZN(n6851)
         );
  AOI21_X1 U8484 ( .B1(n9406), .B2(n6970), .A(n6851), .ZN(n6855) );
  NAND2_X1 U8485 ( .A1(n6852), .A2(n6970), .ZN(n6853) );
  AND2_X1 U8486 ( .A1(n6932), .A2(n6853), .ZN(n6971) );
  NAND2_X1 U8487 ( .A1(n6971), .A2(n9237), .ZN(n6854) );
  OAI211_X1 U8488 ( .C1(n6974), .C2(n7333), .A(n6855), .B(n6854), .ZN(n6856)
         );
  INV_X1 U8489 ( .A(n6856), .ZN(n6857) );
  OAI21_X1 U8490 ( .B1(n6973), .B2(n9405), .A(n6857), .ZN(P1_U3283) );
  OAI222_X1 U8491 ( .A1(n7628), .A2(n6860), .B1(n7626), .B2(n6859), .C1(n6858), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  AND2_X1 U8492 ( .A1(n6948), .A2(n6861), .ZN(n6864) );
  OAI211_X1 U8493 ( .C1(n6864), .C2(n6863), .A(n8595), .B(n6862), .ZN(n6869)
         );
  INV_X1 U8494 ( .A(n6996), .ZN(n8881) );
  AOI21_X1 U8495 ( .B1(n8611), .B2(n8881), .A(n6865), .ZN(n6866) );
  OAI21_X1 U8496 ( .B1(n7327), .B2(n8615), .A(n6866), .ZN(n6867) );
  AOI21_X1 U8497 ( .B1(n7023), .B2(n8612), .A(n6867), .ZN(n6868) );
  OAI211_X1 U8498 ( .C1(n7025), .C2(n8604), .A(n6869), .B(n6868), .ZN(P1_U3234) );
  INV_X1 U8499 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6870) );
  MUX2_X1 U8500 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6870), .S(n6963), .Z(n6873)
         );
  AOI21_X1 U8501 ( .B1(n6878), .B2(P2_REG1_REG_11__SCAN_IN), .A(n6871), .ZN(
        n6872) );
  NAND2_X1 U8502 ( .A1(n6872), .A2(n6873), .ZN(n6962) );
  OAI21_X1 U8503 ( .B1(n6873), .B2(n6872), .A(n6962), .ZN(n6877) );
  NAND2_X1 U8504 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7485) );
  INV_X1 U8505 ( .A(n7485), .ZN(n6876) );
  INV_X1 U8506 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6874) );
  NOR2_X1 U8507 ( .A1(n8151), .A2(n6874), .ZN(n6875) );
  AOI211_X1 U8508 ( .C1(n9694), .C2(n6877), .A(n6876), .B(n6875), .ZN(n6885)
         );
  NOR2_X1 U8509 ( .A1(n6878), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6880) );
  NOR2_X1 U8510 ( .A1(n6880), .A2(n6879), .ZN(n6883) );
  INV_X1 U8511 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6881) );
  MUX2_X1 U8512 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n6881), .S(n6963), .Z(n6882)
         );
  NAND2_X1 U8513 ( .A1(n6882), .A2(n6883), .ZN(n6957) );
  OAI211_X1 U8514 ( .C1(n6883), .C2(n6882), .A(n9695), .B(n6957), .ZN(n6884)
         );
  OAI211_X1 U8515 ( .C1(n9699), .C2(n6886), .A(n6885), .B(n6884), .ZN(P2_U3257) );
  NOR2_X1 U8516 ( .A1(n6887), .A2(n6888), .ZN(n6890) );
  NOR2_X1 U8517 ( .A1(n6890), .A2(n6889), .ZN(n6917) );
  INV_X1 U8518 ( .A(n6917), .ZN(n6892) );
  AND2_X1 U8519 ( .A1(n6887), .A2(n6888), .ZN(n6916) );
  OAI21_X1 U8520 ( .B1(n6890), .B2(n6916), .A(n6889), .ZN(n6891) );
  OAI21_X1 U8521 ( .B1(n6892), .B2(n6916), .A(n6891), .ZN(n6900) );
  INV_X1 U8522 ( .A(n9393), .ZN(n8882) );
  NOR2_X1 U8523 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6893), .ZN(n9583) );
  AOI21_X1 U8524 ( .B1(n8578), .B2(n8882), .A(n9583), .ZN(n6898) );
  NAND2_X1 U8525 ( .A1(n8617), .A2(n6970), .ZN(n6897) );
  NAND2_X1 U8526 ( .A1(n8612), .A2(n6894), .ZN(n6896) );
  NAND2_X1 U8527 ( .A1(n8611), .A2(n8884), .ZN(n6895) );
  NAND4_X1 U8528 ( .A1(n6898), .A2(n6897), .A3(n6896), .A4(n6895), .ZN(n6899)
         );
  AOI21_X1 U8529 ( .B1(n6900), .B2(n8595), .A(n6899), .ZN(n6901) );
  INV_X1 U8530 ( .A(n6901), .ZN(P1_U3219) );
  INV_X1 U8531 ( .A(n6902), .ZN(n6904) );
  OAI222_X1 U8532 ( .A1(n9364), .A2(n6904), .B1(n8830), .B2(P1_U3084), .C1(
        n6903), .C2(n9360), .ZN(P1_U3332) );
  OAI222_X1 U8533 ( .A1(n7628), .A2(n6905), .B1(n7626), .B2(n6904), .C1(n7799), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  INV_X1 U8534 ( .A(n7311), .ZN(n9480) );
  AOI21_X1 U8535 ( .B1(n6862), .B2(n6907), .A(n6906), .ZN(n6908) );
  OAI21_X1 U8536 ( .B1(n4367), .B2(n6908), .A(n8595), .ZN(n6913) );
  INV_X1 U8537 ( .A(n8880), .ZN(n9395) );
  AOI21_X1 U8538 ( .B1(n8578), .B2(n8878), .A(n6909), .ZN(n6910) );
  OAI21_X1 U8539 ( .B1(n9395), .B2(n8599), .A(n6910), .ZN(n6911) );
  AOI21_X1 U8540 ( .B1(n7017), .B2(n8612), .A(n6911), .ZN(n6912) );
  OAI211_X1 U8541 ( .C1(n9480), .C2(n8604), .A(n6913), .B(n6912), .ZN(P1_U3222) );
  AND2_X1 U8542 ( .A1(n6946), .A2(n6914), .ZN(n6915) );
  OAI21_X1 U8543 ( .B1(n6917), .B2(n6916), .A(n6915), .ZN(n6947) );
  INV_X1 U8544 ( .A(n6947), .ZN(n6919) );
  NOR3_X1 U8545 ( .A1(n6917), .A2(n6916), .A3(n6915), .ZN(n6918) );
  OAI21_X1 U8546 ( .B1(n6919), .B2(n6918), .A(n8595), .ZN(n6923) );
  AND2_X1 U8547 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9599) );
  AOI21_X1 U8548 ( .B1(n8578), .B2(n8881), .A(n9599), .ZN(n6920) );
  OAI21_X1 U8549 ( .B1(n6926), .B2(n8599), .A(n6920), .ZN(n6921) );
  AOI21_X1 U8550 ( .B1(n6933), .B2(n8612), .A(n6921), .ZN(n6922) );
  OAI211_X1 U8551 ( .C1(n6993), .C2(n8604), .A(n6923), .B(n6922), .ZN(P1_U3229) );
  INV_X1 U8552 ( .A(n8820), .ZN(n8670) );
  AND2_X1 U8553 ( .A1(n6993), .A2(n8882), .ZN(n8683) );
  NAND2_X1 U8554 ( .A1(n7112), .A2(n9393), .ZN(n9389) );
  INV_X1 U8555 ( .A(n9389), .ZN(n6925) );
  XNOR2_X1 U8556 ( .A(n7000), .B(n8759), .ZN(n6931) );
  OAI22_X1 U8557 ( .A1(n6926), .A2(n9392), .B1(n6996), .B2(n9394), .ZN(n6930)
         );
  NAND2_X1 U8558 ( .A1(n6970), .A2(n8883), .ZN(n6927) );
  XNOR2_X1 U8559 ( .A(n6995), .B(n8759), .ZN(n7116) );
  NOR2_X1 U8560 ( .A1(n7116), .A2(n9398), .ZN(n6929) );
  AOI211_X1 U8561 ( .C1(n9401), .C2(n6931), .A(n6930), .B(n6929), .ZN(n7115)
         );
  AOI21_X1 U8562 ( .B1(n7112), .B2(n6932), .A(n4366), .ZN(n7113) );
  AOI22_X1 U8563 ( .A1(n9405), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n6933), .B2(
        n9404), .ZN(n6934) );
  OAI21_X1 U8564 ( .B1(n6993), .B2(n9217), .A(n6934), .ZN(n6936) );
  NOR2_X1 U8565 ( .A1(n7116), .A2(n7333), .ZN(n6935) );
  AOI211_X1 U8566 ( .C1(n7113), .C2(n9237), .A(n6936), .B(n6935), .ZN(n6937)
         );
  OAI21_X1 U8567 ( .B1(n7115), .B2(n9405), .A(n6937), .ZN(P1_U3282) );
  INV_X1 U8568 ( .A(n6938), .ZN(n7102) );
  AOI211_X1 U8569 ( .C1(n6940), .C2(n6939), .A(n9431), .B(n7102), .ZN(n6944)
         );
  AOI22_X1 U8570 ( .A1(n9682), .A2(n8021), .B1(n9435), .B2(n7458), .ZN(n6942)
         );
  AOI22_X1 U8571 ( .A1(n7782), .A2(n7459), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n6941) );
  OAI211_X1 U8572 ( .C1(n7191), .C2(n7789), .A(n6942), .B(n6941), .ZN(n6943)
         );
  OR2_X1 U8573 ( .A1(n6944), .A2(n6943), .ZN(P2_U3229) );
  AND3_X1 U8574 ( .A1(n6947), .A2(n6946), .A3(n6945), .ZN(n6950) );
  INV_X1 U8575 ( .A(n6948), .ZN(n6949) );
  OAI21_X1 U8576 ( .B1(n6950), .B2(n6949), .A(n8595), .ZN(n6956) );
  INV_X1 U8577 ( .A(n6951), .ZN(n6952) );
  AOI21_X1 U8578 ( .B1(n8578), .B2(n8880), .A(n6952), .ZN(n6953) );
  OAI21_X1 U8579 ( .B1(n9393), .B2(n8599), .A(n6953), .ZN(n6954) );
  AOI21_X1 U8580 ( .B1(n9403), .B2(n8612), .A(n6954), .ZN(n6955) );
  OAI211_X1 U8581 ( .C1(n9417), .C2(n8604), .A(n6956), .B(n6955), .ZN(P1_U3215) );
  NAND2_X1 U8582 ( .A1(n6963), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6958) );
  NAND2_X1 U8583 ( .A1(n6958), .A2(n6957), .ZN(n6960) );
  INV_X1 U8584 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7085) );
  AOI22_X1 U8585 ( .A1(n7091), .A2(n7085), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7086), .ZN(n6959) );
  NOR2_X1 U8586 ( .A1(n6960), .A2(n6959), .ZN(n7084) );
  AOI21_X1 U8587 ( .B1(n6960), .B2(n6959), .A(n7084), .ZN(n6969) );
  AND2_X1 U8588 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7520) );
  NOR2_X1 U8589 ( .A1(n9699), .A2(n7086), .ZN(n6961) );
  AOI211_X1 U8590 ( .C1(P2_ADDR_REG_13__SCAN_IN), .C2(n9697), .A(n7520), .B(
        n6961), .ZN(n6968) );
  INV_X1 U8591 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9462) );
  AOI22_X1 U8592 ( .A1(n7091), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n9462), .B2(
        n7086), .ZN(n6965) );
  OAI21_X1 U8593 ( .B1(n6963), .B2(P2_REG1_REG_12__SCAN_IN), .A(n6962), .ZN(
        n6964) );
  NAND2_X1 U8594 ( .A1(n6965), .A2(n6964), .ZN(n7090) );
  OAI21_X1 U8595 ( .B1(n6965), .B2(n6964), .A(n7090), .ZN(n6966) );
  NAND2_X1 U8596 ( .A1(n6966), .A2(n9694), .ZN(n6967) );
  OAI211_X1 U8597 ( .C1(n6969), .C2(n9698), .A(n6968), .B(n6967), .ZN(P2_U3258) );
  INV_X1 U8598 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6976) );
  AOI22_X1 U8599 ( .A1(n6971), .A2(n9409), .B1(n9330), .B2(n6970), .ZN(n6972)
         );
  OAI211_X1 U8600 ( .C1(n9663), .C2(n6974), .A(n6973), .B(n6972), .ZN(n6977)
         );
  NAND2_X1 U8601 ( .A1(n6977), .A2(n9334), .ZN(n6975) );
  OAI21_X1 U8602 ( .B1(n9334), .B2(n6976), .A(n6975), .ZN(P1_U3531) );
  INV_X1 U8603 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6979) );
  NAND2_X1 U8604 ( .A1(n6977), .A2(n9352), .ZN(n6978) );
  OAI21_X1 U8605 ( .B1(n9352), .B2(n6979), .A(n6978), .ZN(P1_U3478) );
  INV_X1 U8606 ( .A(n6980), .ZN(n7625) );
  OAI222_X1 U8607 ( .A1(n9360), .A2(n6981), .B1(n9364), .B2(n7625), .C1(
        P1_U3084), .C2(n5654), .ZN(P1_U3331) );
  NOR2_X1 U8608 ( .A1(n4779), .A2(n6984), .ZN(n6985) );
  XNOR2_X1 U8609 ( .A(n6982), .B(n6985), .ZN(n6992) );
  INV_X1 U8610 ( .A(n6986), .ZN(n7332) );
  NOR2_X1 U8611 ( .A1(n8599), .A2(n7327), .ZN(n6987) );
  AOI211_X1 U8612 ( .C1(n8578), .C2(n4509), .A(n6988), .B(n6987), .ZN(n6989)
         );
  OAI21_X1 U8613 ( .B1(n8588), .B2(n7332), .A(n6989), .ZN(n6990) );
  AOI21_X1 U8614 ( .B1(n9329), .B2(n8617), .A(n6990), .ZN(n6991) );
  OAI21_X1 U8615 ( .B1(n6992), .B2(n8619), .A(n6991), .ZN(P1_U3232) );
  INV_X1 U8616 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7005) );
  NOR2_X1 U8617 ( .A1(n6993), .A2(n9393), .ZN(n6994) );
  OR2_X1 U8618 ( .A1(n9407), .A2(n6996), .ZN(n8685) );
  NAND2_X1 U8619 ( .A1(n9407), .A2(n6996), .ZN(n8687) );
  NAND2_X1 U8620 ( .A1(n8685), .A2(n8687), .ZN(n9396) );
  NAND2_X1 U8621 ( .A1(n9397), .A2(n9396), .ZN(n6998) );
  NAND2_X1 U8622 ( .A1(n9417), .A2(n6996), .ZN(n6997) );
  XNOR2_X1 U8623 ( .A(n7012), .B(n8880), .ZN(n8761) );
  XOR2_X1 U8624 ( .A(n6999), .B(n8761), .Z(n7031) );
  INV_X1 U8625 ( .A(n8685), .ZN(n8783) );
  NAND2_X1 U8626 ( .A1(n8687), .A2(n9389), .ZN(n8671) );
  NAND2_X1 U8627 ( .A1(n8671), .A2(n8685), .ZN(n8784) );
  XNOR2_X1 U8628 ( .A(n7009), .B(n8761), .ZN(n7001) );
  INV_X1 U8629 ( .A(n7327), .ZN(n8879) );
  AOI222_X1 U8630 ( .A1(n9401), .A2(n7001), .B1(n8881), .B2(n9231), .C1(n8879), 
        .C2(n9232), .ZN(n7026) );
  INV_X1 U8631 ( .A(n7002), .ZN(n9410) );
  NAND2_X1 U8632 ( .A1(n7002), .A2(n7025), .ZN(n7015) );
  INV_X1 U8633 ( .A(n7015), .ZN(n7016) );
  AOI21_X1 U8634 ( .B1(n7012), .B2(n9410), .A(n7016), .ZN(n7029) );
  AOI22_X1 U8635 ( .A1(n7029), .A2(n9409), .B1(n9330), .B2(n7012), .ZN(n7003)
         );
  OAI211_X1 U8636 ( .C1(n7031), .C2(n9332), .A(n7026), .B(n7003), .ZN(n7006)
         );
  NAND2_X1 U8637 ( .A1(n7006), .A2(n9352), .ZN(n7004) );
  OAI21_X1 U8638 ( .B1(n9352), .B2(n7005), .A(n7004), .ZN(P1_U3487) );
  NAND2_X1 U8639 ( .A1(n7006), .A2(n9334), .ZN(n7007) );
  OAI21_X1 U8640 ( .B1(n9334), .B2(n7008), .A(n7007), .ZN(P1_U3534) );
  AND2_X1 U8641 ( .A1(n7012), .A2(n9395), .ZN(n8676) );
  OR2_X1 U8642 ( .A1(n7012), .A2(n9395), .ZN(n7302) );
  NAND2_X1 U8643 ( .A1(n7303), .A2(n7302), .ZN(n7010) );
  OR2_X1 U8644 ( .A1(n7311), .A2(n7327), .ZN(n8678) );
  NAND2_X1 U8645 ( .A1(n7311), .A2(n7327), .ZN(n8691) );
  NAND2_X1 U8646 ( .A1(n8678), .A2(n8691), .ZN(n7310) );
  XNOR2_X1 U8647 ( .A(n7010), .B(n7310), .ZN(n7011) );
  AOI222_X1 U8648 ( .A1(n9401), .A2(n7011), .B1(n8878), .B2(n9232), .C1(n8880), 
        .C2(n9231), .ZN(n9478) );
  INV_X1 U8649 ( .A(n7310), .ZN(n8763) );
  XNOR2_X1 U8650 ( .A(n7309), .B(n8763), .ZN(n9483) );
  INV_X1 U8651 ( .A(n9239), .ZN(n9030) );
  NAND2_X1 U8652 ( .A1(n9483), .A2(n9030), .ZN(n7022) );
  OAI211_X1 U8653 ( .C1(n7016), .C2(n9480), .A(n9409), .B(n7324), .ZN(n9477)
         );
  INV_X1 U8654 ( .A(n9477), .ZN(n7020) );
  AOI22_X1 U8655 ( .A1(n9405), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7017), .B2(
        n9404), .ZN(n7018) );
  OAI21_X1 U8656 ( .B1(n9480), .B2(n9217), .A(n7018), .ZN(n7019) );
  AOI21_X1 U8657 ( .B1(n7020), .B2(n9412), .A(n7019), .ZN(n7021) );
  OAI211_X1 U8658 ( .C1(n9405), .C2(n9478), .A(n7022), .B(n7021), .ZN(P1_U3279) );
  AOI22_X1 U8659 ( .A1(n9405), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7023), .B2(
        n9404), .ZN(n7024) );
  OAI21_X1 U8660 ( .B1(n7025), .B2(n9217), .A(n7024), .ZN(n7028) );
  NOR2_X1 U8661 ( .A1(n7026), .A2(n9405), .ZN(n7027) );
  AOI211_X1 U8662 ( .C1(n7029), .C2(n9237), .A(n7028), .B(n7027), .ZN(n7030)
         );
  OAI21_X1 U8663 ( .B1(n9239), .B2(n7031), .A(n7030), .ZN(P1_U3280) );
  INV_X1 U8664 ( .A(n7072), .ZN(n7034) );
  AOI21_X1 U8665 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8491), .A(n7032), .ZN(
        n7033) );
  OAI21_X1 U8666 ( .B1(n7034), .B2(n7626), .A(n7033), .ZN(P2_U3335) );
  INV_X1 U8667 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10062) );
  NOR2_X1 U8668 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7035) );
  AOI21_X1 U8669 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7035), .ZN(n9839) );
  NOR2_X1 U8670 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7036) );
  AOI21_X1 U8671 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7036), .ZN(n9842) );
  NOR2_X1 U8672 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7037) );
  AOI21_X1 U8673 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7037), .ZN(n9845) );
  NOR2_X1 U8674 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7038) );
  AOI21_X1 U8675 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7038), .ZN(n9848) );
  NOR2_X1 U8676 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7039) );
  AOI21_X1 U8677 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7039), .ZN(n9851) );
  NOR2_X1 U8678 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7045) );
  XOR2_X1 U8679 ( .A(n9865), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10073) );
  NAND2_X1 U8680 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7043) );
  XOR2_X1 U8681 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10071) );
  NAND2_X1 U8682 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7041) );
  XOR2_X1 U8683 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10069) );
  AOI21_X1 U8684 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9831) );
  INV_X1 U8685 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9835) );
  NAND3_X1 U8686 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9833) );
  OAI21_X1 U8687 ( .B1(n9831), .B2(n9835), .A(n9833), .ZN(n10068) );
  NAND2_X1 U8688 ( .A1(n10069), .A2(n10068), .ZN(n7040) );
  NAND2_X1 U8689 ( .A1(n7041), .A2(n7040), .ZN(n10070) );
  NAND2_X1 U8690 ( .A1(n10071), .A2(n10070), .ZN(n7042) );
  NAND2_X1 U8691 ( .A1(n7043), .A2(n7042), .ZN(n10072) );
  NOR2_X1 U8692 ( .A1(n10073), .A2(n10072), .ZN(n7044) );
  NOR2_X1 U8693 ( .A1(n7045), .A2(n7044), .ZN(n7046) );
  NOR2_X1 U8694 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7046), .ZN(n10057) );
  AND2_X1 U8695 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7046), .ZN(n10056) );
  NOR2_X1 U8696 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10056), .ZN(n7047) );
  NOR2_X1 U8697 ( .A1(n10057), .A2(n7047), .ZN(n7048) );
  NAND2_X1 U8698 ( .A1(n7048), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7050) );
  XOR2_X1 U8699 ( .A(n7048), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10055) );
  NAND2_X1 U8700 ( .A1(n10055), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7049) );
  NAND2_X1 U8701 ( .A1(n7050), .A2(n7049), .ZN(n7051) );
  NAND2_X1 U8702 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7051), .ZN(n7053) );
  INV_X1 U8703 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9582) );
  XNOR2_X1 U8704 ( .A(n9582), .B(n7051), .ZN(n10059) );
  NAND2_X1 U8705 ( .A1(n10059), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7052) );
  NAND2_X1 U8706 ( .A1(n7053), .A2(n7052), .ZN(n7054) );
  NAND2_X1 U8707 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7054), .ZN(n7056) );
  INV_X1 U8708 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10037) );
  XNOR2_X1 U8709 ( .A(n10037), .B(n7054), .ZN(n10064) );
  NAND2_X1 U8710 ( .A1(n10064), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7055) );
  NAND2_X1 U8711 ( .A1(n7056), .A2(n7055), .ZN(n7057) );
  AND2_X1 U8712 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7057), .ZN(n7058) );
  INV_X1 U8713 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10067) );
  XNOR2_X1 U8714 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7057), .ZN(n10066) );
  NOR2_X1 U8715 ( .A1(n10067), .A2(n10066), .ZN(n10065) );
  NOR2_X1 U8716 ( .A1(n7058), .A2(n10065), .ZN(n9860) );
  NAND2_X1 U8717 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7059) );
  OAI21_X1 U8718 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7059), .ZN(n9859) );
  NOR2_X1 U8719 ( .A1(n9860), .A2(n9859), .ZN(n9858) );
  AOI21_X1 U8720 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9858), .ZN(n9857) );
  NAND2_X1 U8721 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7060) );
  OAI21_X1 U8722 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7060), .ZN(n9856) );
  NOR2_X1 U8723 ( .A1(n9857), .A2(n9856), .ZN(n9855) );
  AOI21_X1 U8724 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9855), .ZN(n9854) );
  NOR2_X1 U8725 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7061) );
  AOI21_X1 U8726 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7061), .ZN(n9853) );
  NAND2_X1 U8727 ( .A1(n9854), .A2(n9853), .ZN(n9852) );
  OAI21_X1 U8728 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9852), .ZN(n9850) );
  NAND2_X1 U8729 ( .A1(n9851), .A2(n9850), .ZN(n9849) );
  OAI21_X1 U8730 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9849), .ZN(n9847) );
  NAND2_X1 U8731 ( .A1(n9848), .A2(n9847), .ZN(n9846) );
  OAI21_X1 U8732 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9846), .ZN(n9844) );
  NAND2_X1 U8733 ( .A1(n9845), .A2(n9844), .ZN(n9843) );
  OAI21_X1 U8734 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9843), .ZN(n9841) );
  NAND2_X1 U8735 ( .A1(n9842), .A2(n9841), .ZN(n9840) );
  OAI21_X1 U8736 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9840), .ZN(n9838) );
  NAND2_X1 U8737 ( .A1(n9839), .A2(n9838), .ZN(n9837) );
  OAI21_X1 U8738 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9837), .ZN(n10061) );
  NOR2_X1 U8739 ( .A1(n10062), .A2(n10061), .ZN(n7062) );
  NAND2_X1 U8740 ( .A1(n10062), .A2(n10061), .ZN(n10060) );
  OAI21_X1 U8741 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7062), .A(n10060), .ZN(
        n7064) );
  XNOR2_X1 U8742 ( .A(n4667), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7063) );
  XNOR2_X1 U8743 ( .A(n7064), .B(n7063), .ZN(ADD_1071_U4) );
  NOR2_X1 U8744 ( .A1(n7066), .A2(n7065), .ZN(n9676) );
  AOI211_X1 U8745 ( .C1(n7066), .C2(n7065), .A(n9431), .B(n9676), .ZN(n7070)
         );
  AOI22_X1 U8746 ( .A1(n9682), .A2(n8020), .B1(n9435), .B2(n7874), .ZN(n7068)
         );
  AOI22_X1 U8747 ( .A1(n7782), .A2(n7244), .B1(P2_REG3_REG_7__SCAN_IN), .B2(
        P2_U3152), .ZN(n7067) );
  OAI211_X1 U8748 ( .C1(n7453), .C2(n7789), .A(n7068), .B(n7067), .ZN(n7069)
         );
  OR2_X1 U8749 ( .A1(n7070), .A2(n7069), .ZN(P2_U3215) );
  NAND2_X1 U8750 ( .A1(n7072), .A2(n7071), .ZN(n7074) );
  NAND2_X1 U8751 ( .A1(n7073), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8876) );
  OAI211_X1 U8752 ( .C1(n9965), .C2(n9360), .A(n7074), .B(n8876), .ZN(P1_U3330) );
  INV_X1 U8753 ( .A(n7789), .ZN(n9684) );
  INV_X1 U8754 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8368) );
  MUX2_X1 U8755 ( .A(P2_U3152), .B(n7782), .S(n8368), .Z(n7076) );
  OAI22_X1 U8756 ( .A1(n7790), .A2(n7191), .B1(n9734), .B2(n9687), .ZN(n7075)
         );
  AOI211_X1 U8757 ( .C1(n9684), .C2(n8025), .A(n7076), .B(n7075), .ZN(n7083)
         );
  NOR3_X1 U8758 ( .A1(n7772), .A2(n7077), .A3(n8373), .ZN(n7081) );
  INV_X1 U8759 ( .A(n7078), .ZN(n7079) );
  AOI21_X1 U8760 ( .B1(n7754), .B2(n7079), .A(n9431), .ZN(n7080) );
  OAI21_X1 U8761 ( .B1(n7081), .B2(n7080), .A(n7156), .ZN(n7082) );
  NAND2_X1 U8762 ( .A1(n7083), .A2(n7082), .ZN(P2_U3220) );
  AOI21_X1 U8763 ( .B1(n7086), .B2(n7085), .A(n7084), .ZN(n7089) );
  INV_X1 U8764 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7087) );
  AOI22_X1 U8765 ( .A1(n8073), .A2(n7087), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7095), .ZN(n7088) );
  NOR2_X1 U8766 ( .A1(n7089), .A2(n7088), .ZN(n8069) );
  AOI21_X1 U8767 ( .B1(n7089), .B2(n7088), .A(n8069), .ZN(n7099) );
  INV_X1 U8768 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9455) );
  AOI22_X1 U8769 ( .A1(n8073), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n9455), .B2(
        n7095), .ZN(n7093) );
  OAI21_X1 U8770 ( .B1(n7091), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7090), .ZN(
        n7092) );
  NAND2_X1 U8771 ( .A1(n7093), .A2(n7092), .ZN(n8072) );
  OAI21_X1 U8772 ( .B1(n7093), .B2(n7092), .A(n8072), .ZN(n7097) );
  NAND2_X1 U8773 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n9425) );
  NAND2_X1 U8774 ( .A1(n9697), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7094) );
  OAI211_X1 U8775 ( .C1(n9699), .C2(n7095), .A(n9425), .B(n7094), .ZN(n7096)
         );
  AOI21_X1 U8776 ( .B1(n7097), .B2(n9694), .A(n7096), .ZN(n7098) );
  OAI21_X1 U8777 ( .B1(n7099), .B2(n9698), .A(n7098), .ZN(P2_U3259) );
  NOR3_X1 U8778 ( .A1(n7772), .A2(n7100), .A3(n7411), .ZN(n7101) );
  AOI21_X1 U8779 ( .B1(n7102), .B2(n9674), .A(n7101), .ZN(n7111) );
  INV_X1 U8780 ( .A(n7103), .ZN(n7108) );
  OAI22_X1 U8781 ( .A1(n7789), .A2(n7411), .B1(n9755), .B2(n9687), .ZN(n7107)
         );
  INV_X1 U8782 ( .A(n9683), .ZN(n7231) );
  NAND2_X1 U8783 ( .A1(n7782), .A2(n7212), .ZN(n7104) );
  OAI211_X1 U8784 ( .C1(n7790), .C2(n7231), .A(n7105), .B(n7104), .ZN(n7106)
         );
  AOI211_X1 U8785 ( .C1(n7108), .C2(n9674), .A(n7107), .B(n7106), .ZN(n7109)
         );
  OAI21_X1 U8786 ( .B1(n7111), .B2(n7110), .A(n7109), .ZN(P2_U3241) );
  INV_X1 U8787 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7118) );
  AOI22_X1 U8788 ( .A1(n7113), .A2(n9409), .B1(n9330), .B2(n7112), .ZN(n7114)
         );
  OAI211_X1 U8789 ( .C1(n9663), .C2(n7116), .A(n7115), .B(n7114), .ZN(n7119)
         );
  NAND2_X1 U8790 ( .A1(n7119), .A2(n9334), .ZN(n7117) );
  OAI21_X1 U8791 ( .B1(n9334), .B2(n7118), .A(n7117), .ZN(P1_U3532) );
  INV_X1 U8792 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10041) );
  NAND2_X1 U8793 ( .A1(n7119), .A2(n9352), .ZN(n7120) );
  OAI21_X1 U8794 ( .B1(n9352), .B2(n10041), .A(n7120), .ZN(P1_U3481) );
  INV_X1 U8795 ( .A(n7121), .ZN(n7123) );
  NOR2_X1 U8796 ( .A1(n7123), .A2(n7122), .ZN(n7124) );
  XNOR2_X1 U8797 ( .A(n7125), .B(n7124), .ZN(n7131) );
  AOI22_X1 U8798 ( .A1(n9682), .A2(n8019), .B1(n9435), .B2(n7268), .ZN(n7130)
         );
  INV_X1 U8799 ( .A(n7126), .ZN(n7260) );
  OAI21_X1 U8800 ( .B1(n9693), .B2(n7260), .A(n7127), .ZN(n7128) );
  AOI21_X1 U8801 ( .B1(n9684), .B2(n8020), .A(n7128), .ZN(n7129) );
  OAI211_X1 U8802 ( .C1(n7131), .C2(n9431), .A(n7130), .B(n7129), .ZN(P2_U3233) );
  INV_X1 U8803 ( .A(n7132), .ZN(n7137) );
  AOI22_X1 U8804 ( .A1(n7133), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n8491), .ZN(n7134) );
  OAI21_X1 U8805 ( .B1(n7137), .B2(n7626), .A(n7134), .ZN(P2_U3334) );
  OAI222_X1 U8806 ( .A1(n9364), .A2(n7137), .B1(P1_U3084), .B2(n7136), .C1(
        n7135), .C2(n9360), .ZN(P1_U3329) );
  NAND2_X1 U8807 ( .A1(n7139), .A2(n7143), .ZN(n7140) );
  INV_X1 U8808 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9610) );
  NAND2_X1 U8809 ( .A1(n9611), .A2(n9610), .ZN(n9609) );
  INV_X1 U8810 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7141) );
  AOI211_X1 U8811 ( .C1(n7142), .C2(n7141), .A(n8894), .B(n9623), .ZN(n7154)
         );
  INV_X1 U8812 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9476) );
  AOI22_X1 U8813 ( .A1(n9608), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n9476), .B2(
        n7143), .ZN(n9614) );
  OAI21_X1 U8814 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n7145), .A(n7144), .ZN(
        n9613) );
  NAND2_X1 U8815 ( .A1(n9614), .A2(n9613), .ZN(n9612) );
  OAI21_X1 U8816 ( .B1(n9608), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9612), .ZN(
        n8899) );
  XNOR2_X1 U8817 ( .A(n8899), .B(n8900), .ZN(n7147) );
  INV_X1 U8818 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7146) );
  NOR2_X1 U8819 ( .A1(n7146), .A2(n7147), .ZN(n8901) );
  AOI211_X1 U8820 ( .C1(n7147), .C2(n7146), .A(n8901), .B(n9549), .ZN(n7153)
         );
  INV_X1 U8821 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7151) );
  NOR2_X1 U8822 ( .A1(n7148), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8610) );
  AOI21_X1 U8823 ( .B1(n9629), .B2(n7149), .A(n8610), .ZN(n7150) );
  OAI21_X1 U8824 ( .B1(n9621), .B2(n7151), .A(n7150), .ZN(n7152) );
  OR3_X1 U8825 ( .A1(n7154), .A2(n7153), .A3(n7152), .ZN(P1_U3256) );
  OAI21_X1 U8826 ( .B1(n7157), .B2(n7156), .A(n7155), .ZN(n7165) );
  INV_X1 U8827 ( .A(n7157), .ZN(n7159) );
  NAND3_X1 U8828 ( .A1(n9678), .A2(n7159), .A3(n7158), .ZN(n7160) );
  AOI21_X1 U8829 ( .B1(n7160), .B2(n7789), .A(n7412), .ZN(n7164) );
  AOI22_X1 U8830 ( .A1(n9682), .A2(n8022), .B1(n9435), .B2(n7211), .ZN(n7161)
         );
  NAND2_X1 U8831 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n8044) );
  OAI211_X1 U8832 ( .C1(n7162), .C2(n9693), .A(n7161), .B(n8044), .ZN(n7163)
         );
  AOI211_X1 U8833 ( .C1(n9674), .C2(n7165), .A(n7164), .B(n7163), .ZN(n7166)
         );
  INV_X1 U8834 ( .A(n7166), .ZN(P2_U3232) );
  INV_X1 U8835 ( .A(n7167), .ZN(n7169) );
  NAND2_X1 U8836 ( .A1(n7169), .A2(n7168), .ZN(n7171) );
  XNOR2_X1 U8837 ( .A(n7171), .B(n7170), .ZN(n7176) );
  NOR2_X1 U8838 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10020), .ZN(n9607) );
  AOI21_X1 U8839 ( .B1(n8578), .B2(n8958), .A(n9607), .ZN(n7173) );
  NAND2_X1 U8840 ( .A1(n8612), .A2(n7317), .ZN(n7172) );
  OAI211_X1 U8841 ( .C1(n7314), .C2(n8599), .A(n7173), .B(n7172), .ZN(n7174)
         );
  AOI21_X1 U8842 ( .B1(n8955), .B2(n8617), .A(n7174), .ZN(n7175) );
  OAI21_X1 U8843 ( .B1(n7176), .B2(n8619), .A(n7175), .ZN(P1_U3213) );
  INV_X1 U8844 ( .A(n7178), .ZN(n7179) );
  XNOR2_X1 U8845 ( .A(n7182), .B(n6212), .ZN(n7181) );
  OR2_X1 U8846 ( .A1(n7182), .A2(n8395), .ZN(n7224) );
  NAND2_X1 U8847 ( .A1(n8396), .A2(n7224), .ZN(n7183) );
  NAND2_X1 U8848 ( .A1(n7184), .A2(n7186), .ZN(n7855) );
  NAND2_X1 U8849 ( .A1(n7384), .A2(n7376), .ZN(n7188) );
  NAND2_X1 U8850 ( .A1(n7185), .A2(n7186), .ZN(n7187) );
  NAND2_X1 U8851 ( .A1(n7292), .A2(n7812), .ZN(n7190) );
  NAND2_X1 U8852 ( .A1(n8373), .A2(n9729), .ZN(n7189) );
  NAND2_X1 U8853 ( .A1(n7191), .A2(n7211), .ZN(n7844) );
  INV_X1 U8854 ( .A(n7211), .ZN(n9741) );
  NAND2_X1 U8855 ( .A1(n7403), .A2(n7192), .ZN(n7197) );
  NAND2_X1 U8856 ( .A1(n7191), .A2(n9741), .ZN(n7195) );
  NAND2_X1 U8857 ( .A1(n7412), .A2(n9734), .ZN(n7404) );
  INV_X1 U8858 ( .A(n7404), .ZN(n7193) );
  AND2_X1 U8859 ( .A1(n7195), .A2(n7194), .ZN(n7196) );
  NOR2_X1 U8860 ( .A1(n8022), .A2(n7458), .ZN(n7198) );
  NAND2_X1 U8861 ( .A1(n7846), .A2(n4844), .ZN(n7814) );
  OAI22_X1 U8862 ( .A1(n7463), .A2(n7198), .B1(n9750), .B2(n7814), .ZN(n7220)
         );
  NAND2_X1 U8863 ( .A1(n7453), .A2(n7215), .ZN(n7871) );
  NAND2_X1 U8864 ( .A1(n8021), .A2(n9755), .ZN(n7867) );
  AND2_X1 U8865 ( .A1(n7871), .A2(n7867), .ZN(n7206) );
  INV_X1 U8866 ( .A(n7206), .ZN(n7815) );
  XNOR2_X1 U8867 ( .A(n7220), .B(n7815), .ZN(n9754) );
  NAND2_X1 U8868 ( .A1(n8394), .A2(n5719), .ZN(n7808) );
  NAND2_X1 U8869 ( .A1(n7581), .A2(n7586), .ZN(n7381) );
  NAND2_X1 U8870 ( .A1(n7860), .A2(n7200), .ZN(n8379) );
  INV_X1 U8871 ( .A(n7407), .ZN(n7849) );
  NOR2_X1 U8872 ( .A1(n7201), .A2(n7849), .ZN(n7202) );
  NAND2_X1 U8873 ( .A1(n8379), .A2(n7202), .ZN(n7409) );
  NAND2_X1 U8874 ( .A1(n7409), .A2(n7865), .ZN(n7452) );
  INV_X1 U8875 ( .A(n7452), .ZN(n7203) );
  NAND2_X1 U8876 ( .A1(n7204), .A2(n7846), .ZN(n7205) );
  OAI21_X1 U8877 ( .B1(n7206), .B2(n7205), .A(n7225), .ZN(n7207) );
  AOI222_X1 U8878 ( .A1(n8351), .A2(n7207), .B1(n9683), .B2(n8328), .C1(n8022), 
        .C2(n8266), .ZN(n9757) );
  MUX2_X1 U8879 ( .A(n6730), .B(n9757), .S(n8383), .Z(n7217) );
  NOR2_X1 U8880 ( .A1(n5732), .A2(n6858), .ZN(n7208) );
  INV_X1 U8881 ( .A(n7209), .ZN(n7210) );
  NAND2_X1 U8882 ( .A1(n7210), .A2(n8395), .ZN(n7379) );
  AND2_X1 U8883 ( .A1(n7402), .A2(n9750), .ZN(n7456) );
  OAI21_X1 U8884 ( .B1(n7456), .B2(n9755), .A(n7246), .ZN(n9756) );
  INV_X1 U8885 ( .A(n7212), .ZN(n7213) );
  OAI22_X1 U8886 ( .A1(n8358), .A2(n9756), .B1(n7213), .B2(n8218), .ZN(n7214)
         );
  AOI21_X1 U8887 ( .B1(n8363), .B2(n7215), .A(n7214), .ZN(n7216) );
  OAI211_X1 U8888 ( .C1(n8321), .C2(n9754), .A(n7217), .B(n7216), .ZN(P2_U3290) );
  NOR2_X1 U8889 ( .A1(n7453), .A2(n9755), .ZN(n7219) );
  NAND2_X1 U8890 ( .A1(n7453), .A2(n9755), .ZN(n7218) );
  OAI21_X1 U8891 ( .B1(n7220), .B2(n7219), .A(n7218), .ZN(n7241) );
  XNOR2_X1 U8892 ( .A(n9683), .B(n9762), .ZN(n7817) );
  NOR2_X1 U8893 ( .A1(n7874), .A2(n9683), .ZN(n7221) );
  AOI21_X1 U8894 ( .B1(n7241), .B2(n7817), .A(n7221), .ZN(n7222) );
  NAND2_X1 U8895 ( .A1(n7256), .A2(n7238), .ZN(n7880) );
  INV_X1 U8896 ( .A(n7238), .ZN(n9769) );
  NAND2_X1 U8897 ( .A1(n9769), .A2(n8020), .ZN(n7879) );
  NAND2_X1 U8898 ( .A1(n7222), .A2(n7877), .ZN(n7254) );
  OR2_X1 U8899 ( .A1(n7222), .A2(n7877), .ZN(n7223) );
  NAND2_X1 U8900 ( .A1(n7254), .A2(n7223), .ZN(n9768) );
  NAND2_X1 U8901 ( .A1(n9683), .A2(n9762), .ZN(n7226) );
  AND2_X1 U8902 ( .A1(n7228), .A2(n7226), .ZN(n7229) );
  AND2_X1 U8903 ( .A1(n7230), .A2(n7226), .ZN(n7227) );
  OAI21_X1 U8904 ( .B1(n7230), .B2(n7229), .A(n7274), .ZN(n7233) );
  OAI22_X1 U8905 ( .A1(n7231), .A2(n8372), .B1(n8371), .B2(n7277), .ZN(n7232)
         );
  AOI21_X1 U8906 ( .B1(n7233), .B2(n8351), .A(n7232), .ZN(n7234) );
  OAI21_X1 U8907 ( .B1(n9768), .B2(n8396), .A(n7234), .ZN(n9771) );
  MUX2_X1 U8908 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9771), .S(n8383), .Z(n7235)
         );
  INV_X1 U8909 ( .A(n7235), .ZN(n7240) );
  NAND2_X1 U8910 ( .A1(n4365), .A2(n7238), .ZN(n7236) );
  NAND2_X1 U8911 ( .A1(n7261), .A2(n7236), .ZN(n9770) );
  OAI22_X1 U8912 ( .A1(n8358), .A2(n9770), .B1(n9692), .B2(n8218), .ZN(n7237)
         );
  AOI21_X1 U8913 ( .B1(n8363), .B2(n7238), .A(n7237), .ZN(n7239) );
  OAI211_X1 U8914 ( .C1(n9768), .C2(n8340), .A(n7240), .B(n7239), .ZN(P2_U3288) );
  XNOR2_X1 U8915 ( .A(n7241), .B(n7817), .ZN(n9766) );
  INV_X1 U8916 ( .A(n9766), .ZN(n7252) );
  XNOR2_X1 U8917 ( .A(n7242), .B(n7817), .ZN(n7243) );
  OAI222_X1 U8918 ( .A1(n8372), .A2(n7453), .B1(n8371), .B2(n7256), .C1(n8377), 
        .C2(n7243), .ZN(n9764) );
  NAND2_X1 U8919 ( .A1(n9764), .A2(n8383), .ZN(n7251) );
  INV_X1 U8920 ( .A(n7244), .ZN(n7245) );
  OAI22_X1 U8921 ( .A1(n8383), .A2(n6728), .B1(n7245), .B2(n8218), .ZN(n7249)
         );
  INV_X1 U8922 ( .A(n7246), .ZN(n7247) );
  OAI21_X1 U8923 ( .B1(n7247), .B2(n9762), .A(n4365), .ZN(n9763) );
  NOR2_X1 U8924 ( .A1(n8358), .A2(n9763), .ZN(n7248) );
  AOI211_X1 U8925 ( .C1(n8363), .C2(n7874), .A(n7249), .B(n7248), .ZN(n7250)
         );
  OAI211_X1 U8926 ( .C1(n7252), .C2(n8321), .A(n7251), .B(n7250), .ZN(P2_U3289) );
  OR2_X1 U8927 ( .A1(n7256), .A2(n9769), .ZN(n7253) );
  NAND2_X1 U8928 ( .A1(n7254), .A2(n7253), .ZN(n7269) );
  OR2_X1 U8929 ( .A1(n7268), .A2(n7277), .ZN(n7892) );
  NAND2_X1 U8930 ( .A1(n7268), .A2(n7277), .ZN(n7881) );
  XOR2_X1 U8931 ( .A(n7269), .B(n7884), .Z(n9775) );
  NAND2_X1 U8932 ( .A1(n7274), .A2(n7880), .ZN(n7255) );
  XNOR2_X1 U8933 ( .A(n7255), .B(n7884), .ZN(n7258) );
  OAI22_X1 U8934 ( .A1(n7256), .A2(n8372), .B1(n8371), .B2(n7467), .ZN(n7257)
         );
  AOI21_X1 U8935 ( .B1(n7258), .B2(n8351), .A(n7257), .ZN(n7259) );
  OAI21_X1 U8936 ( .B1(n9775), .B2(n8396), .A(n7259), .ZN(n9777) );
  NAND2_X1 U8937 ( .A1(n9777), .A2(n8383), .ZN(n7267) );
  OAI22_X1 U8938 ( .A1(n8383), .A2(n6722), .B1(n7260), .B2(n8218), .ZN(n7265)
         );
  INV_X1 U8939 ( .A(n7261), .ZN(n7263) );
  INV_X1 U8940 ( .A(n7282), .ZN(n7262) );
  OAI21_X1 U8941 ( .B1(n4427), .B2(n7263), .A(n7262), .ZN(n9776) );
  NOR2_X1 U8942 ( .A1(n9776), .A2(n8358), .ZN(n7264) );
  AOI211_X1 U8943 ( .C1(n8363), .C2(n7268), .A(n7265), .B(n7264), .ZN(n7266)
         );
  OAI211_X1 U8944 ( .C1(n9775), .C2(n8340), .A(n7267), .B(n7266), .ZN(P2_U3287) );
  NAND2_X1 U8945 ( .A1(n7338), .A2(n7467), .ZN(n7889) );
  NAND2_X1 U8946 ( .A1(n7890), .A2(n7889), .ZN(n7275) );
  INV_X1 U8947 ( .A(n7275), .ZN(n7885) );
  NAND2_X1 U8948 ( .A1(n7270), .A2(n7885), .ZN(n7271) );
  NAND2_X1 U8949 ( .A1(n7340), .A2(n7271), .ZN(n9781) );
  AND2_X1 U8950 ( .A1(n7880), .A2(n7881), .ZN(n7273) );
  AOI21_X1 U8951 ( .B1(n7276), .B2(n7275), .A(n8377), .ZN(n7279) );
  OR2_X2 U8952 ( .A1(n7276), .A2(n7275), .ZN(n7361) );
  OR2_X1 U8953 ( .A1(n8372), .A2(n7277), .ZN(n7278) );
  OAI21_X1 U8954 ( .B1(n8371), .B2(n7488), .A(n7278), .ZN(n7651) );
  AOI21_X1 U8955 ( .B1(n7279), .B2(n7361), .A(n7651), .ZN(n7280) );
  OAI21_X1 U8956 ( .B1(n9781), .B2(n8396), .A(n7280), .ZN(n9784) );
  NAND2_X1 U8957 ( .A1(n9784), .A2(n8383), .ZN(n7286) );
  INV_X1 U8958 ( .A(n7281), .ZN(n7652) );
  OAI22_X1 U8959 ( .A1(n8383), .A2(n6749), .B1(n7652), .B2(n8218), .ZN(n7284)
         );
  NAND2_X1 U8960 ( .A1(n7282), .A2(n9782), .ZN(n7471) );
  OAI21_X1 U8961 ( .B1(n7282), .B2(n9782), .A(n7471), .ZN(n9783) );
  NOR2_X1 U8962 ( .A1(n9783), .A2(n8358), .ZN(n7283) );
  AOI211_X1 U8963 ( .C1(n8363), .C2(n7338), .A(n7284), .B(n7283), .ZN(n7285)
         );
  OAI211_X1 U8964 ( .C1(n9781), .C2(n8340), .A(n7286), .B(n7285), .ZN(P2_U3286) );
  INV_X1 U8965 ( .A(n7581), .ZN(n8027) );
  NAND2_X1 U8966 ( .A1(n8027), .A2(n9717), .ZN(n7853) );
  NAND2_X1 U8967 ( .A1(n7381), .A2(n7853), .ZN(n9719) );
  INV_X1 U8968 ( .A(n9719), .ZN(n7291) );
  AOI22_X1 U8969 ( .A1(n8328), .A2(n7184), .B1(n8351), .B2(n9719), .ZN(n9716)
         );
  INV_X1 U8970 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7287) );
  OAI22_X1 U8971 ( .A1(n8362), .A2(n9716), .B1(n7287), .B2(n8218), .ZN(n7288)
         );
  AOI21_X1 U8972 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n8362), .A(n7288), .ZN(
        n7290) );
  OAI21_X1 U8973 ( .B1(n8370), .B2(n8363), .A(n7586), .ZN(n7289) );
  OAI211_X1 U8974 ( .C1(n7291), .C2(n8321), .A(n7290), .B(n7289), .ZN(P2_U3296) );
  XNOR2_X1 U8975 ( .A(n7292), .B(n7812), .ZN(n9731) );
  AOI22_X1 U8976 ( .A1(n8252), .A2(n9731), .B1(n8363), .B2(n7751), .ZN(n7300)
         );
  INV_X1 U8977 ( .A(n7293), .ZN(n7377) );
  INV_X1 U8978 ( .A(n8366), .ZN(n7294) );
  AOI211_X1 U8979 ( .C1(n7751), .C2(n7377), .A(n7294), .B(n9801), .ZN(n9726)
         );
  INV_X1 U8980 ( .A(n7379), .ZN(n7298) );
  INV_X1 U8981 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7296) );
  OAI21_X1 U8982 ( .B1(n4845), .B2(n7199), .A(n8376), .ZN(n7295) );
  AOI222_X1 U8983 ( .A1(n8351), .A2(n7295), .B1(n7184), .B2(n8266), .C1(n8024), 
        .C2(n8328), .ZN(n9728) );
  OAI21_X1 U8984 ( .B1(n7296), .B2(n8218), .A(n9728), .ZN(n7297) );
  AOI22_X1 U8985 ( .A1(n9726), .A2(n7298), .B1(n7297), .B2(n8383), .ZN(n7299)
         );
  OAI211_X1 U8986 ( .C1(n7301), .C2(n8383), .A(n7300), .B(n7299), .ZN(P2_U3294) );
  AND2_X1 U8987 ( .A1(n8678), .A2(n7302), .ZN(n8693) );
  NAND2_X1 U8988 ( .A1(n7303), .A2(n8693), .ZN(n7304) );
  NAND2_X1 U8989 ( .A1(n7304), .A2(n8691), .ZN(n7325) );
  XNOR2_X1 U8990 ( .A(n9329), .B(n8878), .ZN(n7329) );
  NAND2_X1 U8991 ( .A1(n7325), .A2(n7329), .ZN(n7305) );
  NAND2_X1 U8992 ( .A1(n9329), .A2(n7314), .ZN(n8675) );
  NAND2_X1 U8993 ( .A1(n8955), .A2(n8954), .ZN(n8698) );
  NAND2_X1 U8994 ( .A1(n8981), .A2(n8698), .ZN(n8749) );
  AOI21_X1 U8995 ( .B1(n7306), .B2(n8749), .A(n9208), .ZN(n7308) );
  OAI22_X1 U8996 ( .A1(n7314), .A2(n9392), .B1(n9210), .B2(n9394), .ZN(n7307)
         );
  AOI21_X1 U8997 ( .B1(n7308), .B2(n8982), .A(n7307), .ZN(n9472) );
  INV_X1 U8998 ( .A(n7309), .ZN(n7313) );
  NAND2_X1 U8999 ( .A1(n7311), .A2(n8879), .ZN(n7312) );
  XNOR2_X1 U9000 ( .A(n8953), .B(n8749), .ZN(n9475) );
  NAND2_X1 U9001 ( .A1(n9475), .A2(n9030), .ZN(n7322) );
  INV_X1 U9002 ( .A(n7316), .ZN(n7323) );
  NOR2_X1 U9003 ( .A1(n7316), .A2(n8955), .ZN(n8941) );
  INV_X1 U9004 ( .A(n8941), .ZN(n9225) );
  OAI211_X1 U9005 ( .C1(n9473), .C2(n7323), .A(n9225), .B(n9409), .ZN(n9471)
         );
  INV_X1 U9006 ( .A(n9471), .ZN(n7320) );
  AOI22_X1 U9007 ( .A1(n9405), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7317), .B2(
        n9404), .ZN(n7318) );
  OAI21_X1 U9008 ( .B1(n9473), .B2(n9217), .A(n7318), .ZN(n7319) );
  AOI21_X1 U9009 ( .B1(n7320), .B2(n9412), .A(n7319), .ZN(n7321) );
  OAI211_X1 U9010 ( .C1(n9405), .C2(n9472), .A(n7322), .B(n7321), .ZN(P1_U3277) );
  AOI211_X1 U9011 ( .C1(n9329), .C2(n7324), .A(n9242), .B(n7323), .ZN(n9328)
         );
  INV_X1 U9012 ( .A(n7329), .ZN(n8766) );
  XNOR2_X1 U9013 ( .A(n7325), .B(n8766), .ZN(n7326) );
  OAI222_X1 U9014 ( .A1(n9394), .A2(n8954), .B1(n9392), .B2(n7327), .C1(n9208), 
        .C2(n7326), .ZN(n9327) );
  XNOR2_X1 U9015 ( .A(n7330), .B(n7329), .ZN(n9333) );
  NOR2_X1 U9016 ( .A1(n9333), .A2(n9398), .ZN(n7331) );
  AOI211_X1 U9017 ( .C1(n9328), .C2(n9646), .A(n9327), .B(n7331), .ZN(n7337)
         );
  OAI22_X1 U9018 ( .A1(n9653), .A2(n6689), .B1(n7332), .B2(n9644), .ZN(n7335)
         );
  NOR2_X1 U9019 ( .A1(n9333), .A2(n7333), .ZN(n7334) );
  AOI211_X1 U9020 ( .C1(n9406), .C2(n9329), .A(n7335), .B(n7334), .ZN(n7336)
         );
  OAI21_X1 U9021 ( .B1(n7337), .B2(n9405), .A(n7336), .ZN(P1_U3278) );
  NAND2_X1 U9022 ( .A1(n7338), .A2(n8019), .ZN(n7339) );
  OR2_X1 U9023 ( .A1(n9789), .A2(n7488), .ZN(n7891) );
  NAND2_X1 U9024 ( .A1(n9789), .A2(n7488), .ZN(n7898) );
  NAND2_X1 U9025 ( .A1(n7891), .A2(n7898), .ZN(n7819) );
  NAND2_X1 U9026 ( .A1(n9789), .A2(n8018), .ZN(n7341) );
  OR2_X1 U9027 ( .A1(n7491), .A2(n7518), .ZN(n7900) );
  NAND2_X1 U9028 ( .A1(n7491), .A2(n7518), .ZN(n7904) );
  NAND2_X1 U9029 ( .A1(n7900), .A2(n7904), .ZN(n7820) );
  INV_X1 U9030 ( .A(n7820), .ZN(n7363) );
  OR2_X1 U9031 ( .A1(n7491), .A2(n8017), .ZN(n7342) );
  OR2_X1 U9032 ( .A1(n7430), .A2(n7487), .ZN(n7909) );
  NAND2_X1 U9033 ( .A1(n7430), .A2(n7487), .ZN(n7439) );
  NAND2_X1 U9034 ( .A1(n7344), .A2(n7811), .ZN(n7345) );
  NAND2_X1 U9035 ( .A1(n7432), .A2(n7345), .ZN(n7354) );
  INV_X1 U9036 ( .A(n7904), .ZN(n7899) );
  AND2_X1 U9037 ( .A1(n7900), .A2(n7891), .ZN(n7903) );
  OR2_X1 U9038 ( .A1(n7899), .A2(n7903), .ZN(n7440) );
  AND2_X1 U9039 ( .A1(n7890), .A2(n7440), .ZN(n7346) );
  NAND2_X1 U9040 ( .A1(n7361), .A2(n7346), .ZN(n7349) );
  INV_X1 U9041 ( .A(n7440), .ZN(n7347) );
  AND2_X1 U9042 ( .A1(n7898), .A2(n7904), .ZN(n7438) );
  OR2_X1 U9043 ( .A1(n7347), .A2(n7438), .ZN(n7348) );
  NAND2_X1 U9044 ( .A1(n7349), .A2(n7348), .ZN(n7350) );
  XNOR2_X1 U9045 ( .A(n7350), .B(n7811), .ZN(n7352) );
  OAI22_X1 U9046 ( .A1(n7518), .A2(n8372), .B1(n8371), .B2(n7788), .ZN(n7351)
         );
  AOI21_X1 U9047 ( .B1(n7352), .B2(n8351), .A(n7351), .ZN(n7353) );
  OAI21_X1 U9048 ( .B1(n7354), .B2(n8396), .A(n7353), .ZN(n9459) );
  INV_X1 U9049 ( .A(n9459), .ZN(n7360) );
  INV_X1 U9050 ( .A(n7354), .ZN(n9461) );
  INV_X1 U9051 ( .A(n8340), .ZN(n8364) );
  INV_X1 U9052 ( .A(n7430), .ZN(n9457) );
  AND2_X1 U9053 ( .A1(n7369), .A2(n9457), .ZN(n7434) );
  NOR2_X1 U9054 ( .A1(n7369), .A2(n9457), .ZN(n7355) );
  OR2_X1 U9055 ( .A1(n7434), .A2(n7355), .ZN(n9458) );
  AOI22_X1 U9056 ( .A1(n8362), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7521), .B2(
        n8369), .ZN(n7357) );
  NAND2_X1 U9057 ( .A1(n8363), .A2(n7430), .ZN(n7356) );
  OAI211_X1 U9058 ( .C1(n9458), .C2(n8358), .A(n7357), .B(n7356), .ZN(n7358)
         );
  AOI21_X1 U9059 ( .B1(n9461), .B2(n8364), .A(n7358), .ZN(n7359) );
  OAI21_X1 U9060 ( .B1(n7360), .B2(n8362), .A(n7359), .ZN(P2_U3283) );
  NAND2_X1 U9061 ( .A1(n7466), .A2(n7898), .ZN(n7362) );
  NAND2_X1 U9062 ( .A1(n7362), .A2(n7891), .ZN(n7364) );
  XNOR2_X1 U9063 ( .A(n7364), .B(n7363), .ZN(n7365) );
  OAI222_X1 U9064 ( .A1(n8371), .A2(n7487), .B1(n8372), .B2(n7488), .C1(n8377), 
        .C2(n7365), .ZN(n9803) );
  INV_X1 U9065 ( .A(n9803), .ZN(n7375) );
  OAI21_X1 U9066 ( .B1(n7367), .B2(n7820), .A(n7366), .ZN(n9805) );
  INV_X1 U9067 ( .A(n7491), .ZN(n9800) );
  INV_X1 U9068 ( .A(n7368), .ZN(n7470) );
  INV_X1 U9069 ( .A(n7369), .ZN(n7370) );
  OAI21_X1 U9070 ( .B1(n9800), .B2(n7470), .A(n7370), .ZN(n9802) );
  AOI22_X1 U9071 ( .A1(n8362), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7484), .B2(
        n8369), .ZN(n7372) );
  NAND2_X1 U9072 ( .A1(n8363), .A2(n7491), .ZN(n7371) );
  OAI211_X1 U9073 ( .C1(n9802), .C2(n8358), .A(n7372), .B(n7371), .ZN(n7373)
         );
  AOI21_X1 U9074 ( .B1(n9805), .B2(n8252), .A(n7373), .ZN(n7374) );
  OAI21_X1 U9075 ( .B1(n7375), .B2(n8362), .A(n7374), .ZN(P2_U3284) );
  XNOR2_X1 U9076 ( .A(n7384), .B(n7376), .ZN(n9724) );
  OAI211_X1 U9077 ( .C1(n7186), .C2(n9717), .A(n9791), .B(n7377), .ZN(n9721)
         );
  INV_X1 U9078 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7378) );
  OAI22_X1 U9079 ( .A1(n7379), .A2(n9721), .B1(n7378), .B2(n8218), .ZN(n7380)
         );
  AOI21_X1 U9080 ( .B1(n8252), .B2(n9724), .A(n7380), .ZN(n7389) );
  INV_X1 U9081 ( .A(n7381), .ZN(n7385) );
  INV_X1 U9082 ( .A(n7855), .ZN(n7382) );
  OAI21_X1 U9083 ( .B1(n7857), .B2(n7382), .A(n8351), .ZN(n7383) );
  AOI21_X1 U9084 ( .B1(n7385), .B2(n7384), .A(n7383), .ZN(n7387) );
  OAI22_X1 U9085 ( .A1(n7581), .A2(n8372), .B1(n8371), .B2(n8373), .ZN(n7386)
         );
  NOR2_X1 U9086 ( .A1(n7387), .A2(n7386), .ZN(n9722) );
  MUX2_X1 U9087 ( .A(n6738), .B(n9722), .S(n8383), .Z(n7388) );
  OAI211_X1 U9088 ( .C1(n7186), .C2(n8311), .A(n7389), .B(n7388), .ZN(P2_U3295) );
  XNOR2_X1 U9089 ( .A(n7391), .B(n7390), .ZN(n7397) );
  INV_X1 U9090 ( .A(n7472), .ZN(n7393) );
  OAI22_X1 U9091 ( .A1(n9693), .A2(n7393), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7392), .ZN(n7395) );
  OAI22_X1 U9092 ( .A1(n7467), .A2(n7789), .B1(n7790), .B2(n7518), .ZN(n7394)
         );
  AOI211_X1 U9093 ( .C1(n9435), .C2(n9789), .A(n7395), .B(n7394), .ZN(n7396)
         );
  OAI21_X1 U9094 ( .B1(n7397), .B2(n9431), .A(n7396), .ZN(P2_U3238) );
  INV_X1 U9095 ( .A(n7398), .ZN(n7429) );
  AOI22_X1 U9096 ( .A1(n7399), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n8491), .ZN(n7400) );
  OAI21_X1 U9097 ( .B1(n7429), .B2(n7626), .A(n7400), .ZN(P2_U3332) );
  INV_X1 U9098 ( .A(n7401), .ZN(n8365) );
  INV_X1 U9099 ( .A(n7402), .ZN(n7457) );
  OAI21_X1 U9100 ( .B1(n9741), .B2(n8365), .A(n7457), .ZN(n9742) );
  OAI22_X1 U9101 ( .A1(n8311), .A2(n9741), .B1(n9742), .B2(n8358), .ZN(n7420)
         );
  NAND2_X1 U9102 ( .A1(n7403), .A2(n8375), .ZN(n7405) );
  NAND2_X1 U9103 ( .A1(n7405), .A2(n7404), .ZN(n7406) );
  XNOR2_X1 U9104 ( .A(n7406), .B(n7201), .ZN(n9745) );
  NAND2_X1 U9105 ( .A1(n8252), .A2(n9745), .ZN(n7418) );
  NAND2_X1 U9106 ( .A1(n8379), .A2(n7407), .ZN(n7408) );
  NAND2_X1 U9107 ( .A1(n7408), .A2(n7201), .ZN(n7410) );
  NAND3_X1 U9108 ( .A1(n7410), .A2(n7409), .A3(n8351), .ZN(n7415) );
  OAI22_X1 U9109 ( .A1(n7412), .A2(n8372), .B1(n8371), .B2(n7411), .ZN(n7413)
         );
  INV_X1 U9110 ( .A(n7413), .ZN(n7414) );
  NAND2_X1 U9111 ( .A1(n7415), .A2(n7414), .ZN(n9743) );
  AOI22_X1 U9112 ( .A1(n8383), .A2(n9743), .B1(n7416), .B2(n8369), .ZN(n7417)
         );
  OAI211_X1 U9113 ( .C1(n9993), .C2(n8383), .A(n7418), .B(n7417), .ZN(n7419)
         );
  OR2_X1 U9114 ( .A1(n7420), .A2(n7419), .ZN(P2_U3292) );
  INV_X1 U9115 ( .A(n7421), .ZN(n7425) );
  INV_X1 U9116 ( .A(n7422), .ZN(n7423) );
  OAI222_X1 U9117 ( .A1(n7628), .A2(n9922), .B1(n7626), .B2(n7425), .C1(n7423), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI222_X1 U9118 ( .A1(n9360), .A2(n7426), .B1(n9364), .B2(n7425), .C1(n7424), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  OAI222_X1 U9119 ( .A1(n9364), .A2(n7429), .B1(P1_U3084), .B2(n7428), .C1(
        n7427), .C2(n9360), .ZN(P1_U3327) );
  NAND2_X1 U9120 ( .A1(n7430), .A2(n8016), .ZN(n7431) );
  XNOR2_X1 U9121 ( .A(n9449), .B(n7788), .ZN(n7913) );
  INV_X1 U9122 ( .A(n7913), .ZN(n7822) );
  OAI21_X1 U9123 ( .B1(n7433), .B2(n7913), .A(n7498), .ZN(n9454) );
  NAND2_X1 U9124 ( .A1(n7434), .A2(n4726), .ZN(n7501) );
  OR2_X1 U9125 ( .A1(n7434), .A2(n4726), .ZN(n7435) );
  NAND2_X1 U9126 ( .A1(n7501), .A2(n7435), .ZN(n9452) );
  OAI22_X1 U9127 ( .A1(n8383), .A2(n7087), .B1(n9438), .B2(n8218), .ZN(n7436)
         );
  AOI21_X1 U9128 ( .B1(n8363), .B2(n9449), .A(n7436), .ZN(n7437) );
  OAI21_X1 U9129 ( .B1(n9452), .B2(n8358), .A(n7437), .ZN(n7450) );
  AND2_X1 U9130 ( .A1(n7438), .A2(n7439), .ZN(n7444) );
  NAND2_X1 U9131 ( .A1(n7466), .A2(n7444), .ZN(n7442) );
  INV_X1 U9132 ( .A(n7439), .ZN(n7911) );
  AND2_X1 U9133 ( .A1(n7811), .A2(n7440), .ZN(n7441) );
  AND2_X1 U9134 ( .A1(n7442), .A2(n7445), .ZN(n7443) );
  AOI21_X1 U9135 ( .B1(n7443), .B2(n7913), .A(n8377), .ZN(n7448) );
  AND2_X1 U9136 ( .A1(n7444), .A2(n7822), .ZN(n7446) );
  OR2_X1 U9137 ( .A1(n8371), .A2(n8344), .ZN(n7447) );
  OAI21_X1 U9138 ( .B1(n8372), .B2(n7487), .A(n7447), .ZN(n9427) );
  AOI21_X1 U9139 ( .B1(n7448), .B2(n7499), .A(n9427), .ZN(n9451) );
  NOR2_X1 U9140 ( .A1(n9451), .A2(n8362), .ZN(n7449) );
  AOI211_X1 U9141 ( .C1(n8252), .C2(n9454), .A(n7450), .B(n7449), .ZN(n7451)
         );
  INV_X1 U9142 ( .A(n7451), .ZN(P2_U3282) );
  XNOR2_X1 U9143 ( .A(n7452), .B(n7814), .ZN(n7455) );
  OAI22_X1 U9144 ( .A1(n7191), .A2(n8372), .B1(n8371), .B2(n7453), .ZN(n7454)
         );
  AOI21_X1 U9145 ( .B1(n7455), .B2(n8351), .A(n7454), .ZN(n9749) );
  AND2_X1 U9146 ( .A1(n8383), .A2(n8395), .ZN(n8319) );
  AOI211_X1 U9147 ( .C1(n7458), .C2(n7457), .A(n9801), .B(n7456), .ZN(n9747)
         );
  INV_X1 U9148 ( .A(n7459), .ZN(n7460) );
  OAI22_X1 U9149 ( .A1(n8383), .A2(n6733), .B1(n7460), .B2(n8218), .ZN(n7462)
         );
  NOR2_X1 U9150 ( .A1(n8311), .A2(n9750), .ZN(n7461) );
  AOI211_X1 U9151 ( .C1(n8319), .C2(n9747), .A(n7462), .B(n7461), .ZN(n7465)
         );
  XNOR2_X1 U9152 ( .A(n7463), .B(n7814), .ZN(n9752) );
  NAND2_X1 U9153 ( .A1(n8252), .A2(n9752), .ZN(n7464) );
  OAI211_X1 U9154 ( .C1(n8362), .C2(n9749), .A(n7465), .B(n7464), .ZN(P2_U3291) );
  XNOR2_X1 U9155 ( .A(n7466), .B(n7819), .ZN(n7469) );
  OAI22_X1 U9156 ( .A1(n7467), .A2(n8372), .B1(n8371), .B2(n7518), .ZN(n7468)
         );
  AOI21_X1 U9157 ( .B1(n7469), .B2(n8351), .A(n7468), .ZN(n9794) );
  AOI21_X1 U9158 ( .B1(n9789), .B2(n7471), .A(n7470), .ZN(n9792) );
  INV_X1 U9159 ( .A(n9789), .ZN(n7474) );
  AOI22_X1 U9160 ( .A1(n8362), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7472), .B2(
        n8369), .ZN(n7473) );
  OAI21_X1 U9161 ( .B1(n8311), .B2(n7474), .A(n7473), .ZN(n7478) );
  OAI21_X1 U9162 ( .B1(n7476), .B2(n7819), .A(n7475), .ZN(n9796) );
  NOR2_X1 U9163 ( .A1(n9796), .A2(n8321), .ZN(n7477) );
  AOI211_X1 U9164 ( .C1(n8370), .C2(n9792), .A(n7478), .B(n7477), .ZN(n7479)
         );
  OAI21_X1 U9165 ( .B1(n8362), .B2(n9794), .A(n7479), .ZN(P2_U3285) );
  NAND2_X1 U9166 ( .A1(n7481), .A2(n7480), .ZN(n7483) );
  XOR2_X1 U9167 ( .A(n7483), .B(n7482), .Z(n7493) );
  INV_X1 U9168 ( .A(n7484), .ZN(n7486) );
  OAI21_X1 U9169 ( .B1(n9693), .B2(n7486), .A(n7485), .ZN(n7490) );
  OAI22_X1 U9170 ( .A1(n7488), .A2(n7789), .B1(n7790), .B2(n7487), .ZN(n7489)
         );
  AOI211_X1 U9171 ( .C1(n9435), .C2(n7491), .A(n7490), .B(n7489), .ZN(n7492)
         );
  OAI21_X1 U9172 ( .B1(n7493), .B2(n9431), .A(n7492), .ZN(P2_U3226) );
  INV_X1 U9173 ( .A(n7494), .ZN(n7510) );
  AOI21_X1 U9174 ( .B1(n9357), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7495), .ZN(
        n7496) );
  OAI21_X1 U9175 ( .B1(n7510), .B2(n9364), .A(n7496), .ZN(P1_U3326) );
  OR2_X1 U9176 ( .A1(n9449), .A2(n8015), .ZN(n7497) );
  NAND2_X1 U9177 ( .A1(n7498), .A2(n7497), .ZN(n7525) );
  NOR2_X1 U9178 ( .A1(n7793), .A2(n8344), .ZN(n7528) );
  INV_X1 U9179 ( .A(n7528), .ZN(n7920) );
  NAND2_X1 U9180 ( .A1(n7793), .A2(n8344), .ZN(n7927) );
  XNOR2_X1 U9181 ( .A(n7525), .B(n4402), .ZN(n9447) );
  INV_X1 U9182 ( .A(n9447), .ZN(n7509) );
  XNOR2_X1 U9183 ( .A(n7529), .B(n7919), .ZN(n7500) );
  OAI222_X1 U9184 ( .A1(n8372), .A2(n7788), .B1(n8371), .B2(n8331), .C1(n8377), 
        .C2(n7500), .ZN(n9445) );
  INV_X1 U9185 ( .A(n7501), .ZN(n7502) );
  INV_X1 U9186 ( .A(n7793), .ZN(n9443) );
  OAI21_X1 U9187 ( .B1(n7502), .B2(n9443), .A(n8352), .ZN(n9444) );
  INV_X1 U9188 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7504) );
  INV_X1 U9189 ( .A(n7503), .ZN(n7787) );
  OAI22_X1 U9190 ( .A1(n8383), .A2(n7504), .B1(n7787), .B2(n8218), .ZN(n7505)
         );
  AOI21_X1 U9191 ( .B1(n8363), .B2(n7793), .A(n7505), .ZN(n7506) );
  OAI21_X1 U9192 ( .B1(n9444), .B2(n8358), .A(n7506), .ZN(n7507) );
  AOI21_X1 U9193 ( .B1(n9445), .B2(n8383), .A(n7507), .ZN(n7508) );
  OAI21_X1 U9194 ( .B1(n7509), .B2(n8321), .A(n7508), .ZN(P2_U3281) );
  OAI222_X1 U9195 ( .A1(n7628), .A2(n7511), .B1(n7626), .B2(n7510), .C1(n7998), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U9196 ( .A(n7512), .ZN(n7623) );
  AOI21_X1 U9197 ( .B1(n8491), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n7513), .ZN(
        n7514) );
  OAI21_X1 U9198 ( .B1(n7623), .B2(n7626), .A(n7514), .ZN(P2_U3330) );
  OAI211_X1 U9199 ( .C1(n7517), .C2(n7516), .A(n7515), .B(n9674), .ZN(n7523)
         );
  OAI22_X1 U9200 ( .A1(n7518), .A2(n7789), .B1(n7790), .B2(n7788), .ZN(n7519)
         );
  AOI211_X1 U9201 ( .C1(n7782), .C2(n7521), .A(n7520), .B(n7519), .ZN(n7522)
         );
  OAI211_X1 U9202 ( .C1(n9457), .C2(n9687), .A(n7523), .B(n7522), .ZN(P2_U3236) );
  NOR2_X1 U9203 ( .A1(n7793), .A2(n8014), .ZN(n7524) );
  OR2_X1 U9204 ( .A1(n8355), .A2(n8331), .ZN(n7922) );
  AND2_X1 U9205 ( .A1(n8355), .A2(n8331), .ZN(n7530) );
  INV_X1 U9206 ( .A(n7530), .ZN(n7921) );
  INV_X1 U9207 ( .A(n8355), .ZN(n8465) );
  XNOR2_X1 U9208 ( .A(n8462), .B(n8012), .ZN(n8325) );
  OR2_X1 U9209 ( .A1(n8455), .A2(n7714), .ZN(n7945) );
  NAND2_X1 U9210 ( .A1(n8455), .A2(n7714), .ZN(n7935) );
  XNOR2_X1 U9211 ( .A(n7589), .B(n7533), .ZN(n8459) );
  INV_X1 U9212 ( .A(n8462), .ZN(n7718) );
  INV_X1 U9213 ( .A(n8307), .ZN(n7526) );
  AOI21_X1 U9214 ( .B1(n8455), .B2(n4437), .A(n7526), .ZN(n8456) );
  AOI22_X1 U9215 ( .A1(n8362), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n7768), .B2(
        n8369), .ZN(n7527) );
  OAI21_X1 U9216 ( .B1(n7771), .B2(n8311), .A(n7527), .ZN(n7538) );
  AOI21_X1 U9217 ( .B1(n8342), .B2(n7922), .A(n7530), .ZN(n8326) );
  NAND2_X1 U9218 ( .A1(n8326), .A2(n8325), .ZN(n8324) );
  INV_X1 U9219 ( .A(n8324), .ZN(n7531) );
  INV_X1 U9220 ( .A(n8012), .ZN(n8343) );
  OR2_X1 U9221 ( .A1(n8462), .A2(n8343), .ZN(n7532) );
  INV_X1 U9222 ( .A(n7532), .ZN(n7930) );
  INV_X1 U9223 ( .A(n7533), .ZN(n7825) );
  OAI21_X1 U9224 ( .B1(n7531), .B2(n7930), .A(n7825), .ZN(n7534) );
  NAND3_X1 U9225 ( .A1(n8324), .A2(n7533), .A3(n7532), .ZN(n7601) );
  AOI21_X1 U9226 ( .B1(n7534), .B2(n7601), .A(n8377), .ZN(n7536) );
  OR2_X1 U9227 ( .A1(n8372), .A2(n8343), .ZN(n7535) );
  OAI21_X1 U9228 ( .B1(n8371), .B2(n8296), .A(n7535), .ZN(n7765) );
  NOR2_X1 U9229 ( .A1(n7536), .A2(n7765), .ZN(n8458) );
  NOR2_X1 U9230 ( .A1(n8458), .A2(n8362), .ZN(n7537) );
  AOI211_X1 U9231 ( .C1(n8456), .C2(n8370), .A(n7538), .B(n7537), .ZN(n7539)
         );
  OAI21_X1 U9232 ( .B1(n8459), .B2(n8321), .A(n7539), .ZN(P2_U3278) );
  INV_X1 U9233 ( .A(n7542), .ZN(n7544) );
  NAND2_X1 U9234 ( .A1(n7544), .A2(n7543), .ZN(n7545) );
  INV_X1 U9235 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7579) );
  INV_X1 U9236 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9361) );
  MUX2_X1 U9237 ( .A(n7579), .B(n9361), .S(n7554), .Z(n7559) );
  INV_X1 U9238 ( .A(n7559), .ZN(n7546) );
  NOR2_X1 U9239 ( .A1(n7546), .A2(SI_29_), .ZN(n7547) );
  MUX2_X1 U9240 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7548), .Z(n7550) );
  INV_X1 U9241 ( .A(n7564), .ZN(n7549) );
  NAND2_X1 U9242 ( .A1(n7549), .A2(SI_30_), .ZN(n7553) );
  NAND2_X1 U9243 ( .A1(n7551), .A2(n7550), .ZN(n7552) );
  NAND2_X1 U9244 ( .A1(n7553), .A2(n7552), .ZN(n7557) );
  MUX2_X1 U9245 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7554), .Z(n7555) );
  XNOR2_X1 U9246 ( .A(n7555), .B(SI_31_), .ZN(n7556) );
  NAND2_X1 U9247 ( .A1(n7566), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7558) );
  INV_X1 U9248 ( .A(n8419), .ZN(n7697) );
  NAND2_X1 U9249 ( .A1(n8164), .A2(n8177), .ZN(n8159) );
  XNOR2_X1 U9250 ( .A(n7559), .B(SI_29_), .ZN(n7560) );
  NAND2_X1 U9251 ( .A1(n8634), .A2(n7565), .ZN(n7563) );
  NAND2_X1 U9252 ( .A1(n7566), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7562) );
  XNOR2_X1 U9253 ( .A(n7564), .B(SI_30_), .ZN(n8621) );
  NAND2_X1 U9254 ( .A1(n8621), .A2(n7565), .ZN(n7568) );
  NAND2_X1 U9255 ( .A1(n7566), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7567) );
  AOI21_X1 U9256 ( .B1(n7569), .B2(P2_B_REG_SCAN_IN), .A(n8371), .ZN(n7608) );
  NAND2_X1 U9257 ( .A1(n7608), .A2(n7803), .ZN(n9439) );
  NOR2_X1 U9258 ( .A1(n8362), .A2(n9439), .ZN(n8154) );
  AOI21_X1 U9259 ( .B1(n8362), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8154), .ZN(
        n7571) );
  NAND2_X1 U9260 ( .A1(n7805), .A2(n8363), .ZN(n7570) );
  OAI211_X1 U9261 ( .C1(n8388), .C2(n8358), .A(n7571), .B(n7570), .ZN(P2_U3265) );
  AOI21_X1 U9262 ( .B1(n7574), .B2(n7572), .A(n7573), .ZN(n7578) );
  AOI22_X1 U9263 ( .A1(n6457), .A2(n8617), .B1(n8611), .B2(n8891), .ZN(n7577)
         );
  AOI22_X1 U9264 ( .A1(n8578), .A2(n8888), .B1(n7575), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7576) );
  OAI211_X1 U9265 ( .C1(n7578), .C2(n8619), .A(n7577), .B(n7576), .ZN(P1_U3235) );
  INV_X1 U9266 ( .A(n8634), .ZN(n9363) );
  OAI222_X1 U9267 ( .A1(n7580), .A2(P2_U3152), .B1(n7626), .B2(n9363), .C1(
        n7579), .C2(n7628), .ZN(P2_U3329) );
  OAI22_X1 U9268 ( .A1(n7772), .A2(n7581), .B1(n9717), .B2(n9431), .ZN(n7583)
         );
  NAND2_X1 U9269 ( .A1(n7583), .A2(n7582), .ZN(n7588) );
  NAND2_X1 U9270 ( .A1(n7585), .A2(n7584), .ZN(n7750) );
  AOI22_X1 U9271 ( .A1(n9435), .A2(n7586), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n7750), .ZN(n7587) );
  OAI211_X1 U9272 ( .C1(n7185), .C2(n7790), .A(n7588), .B(n7587), .ZN(P2_U3234) );
  INV_X1 U9273 ( .A(n8422), .ZN(n8229) );
  OAI22_X1 U9274 ( .A1(n7591), .A2(n7590), .B1(n8327), .B2(n8455), .ZN(n8304)
         );
  INV_X1 U9275 ( .A(n8451), .ZN(n8312) );
  NAND2_X1 U9276 ( .A1(n8312), .A2(n8296), .ZN(n7593) );
  NAND2_X1 U9277 ( .A1(n8445), .A2(n8277), .ZN(n7949) );
  INV_X1 U9278 ( .A(n8445), .ZN(n8291) );
  NOR2_X1 U9279 ( .A1(n7595), .A2(n8297), .ZN(n7596) );
  NAND2_X1 U9280 ( .A1(n8434), .A2(n8278), .ZN(n7940) );
  OR2_X1 U9281 ( .A1(n8427), .A2(n7745), .ZN(n7957) );
  NAND2_X1 U9282 ( .A1(n8427), .A2(n7745), .ZN(n7943) );
  NAND2_X1 U9283 ( .A1(n7957), .A2(n7943), .ZN(n8250) );
  NAND2_X1 U9284 ( .A1(n8251), .A2(n8250), .ZN(n8429) );
  INV_X1 U9285 ( .A(n8427), .ZN(n8248) );
  NAND2_X1 U9286 ( .A1(n8427), .A2(n7599), .ZN(n7600) );
  NAND2_X1 U9287 ( .A1(n8422), .A2(n8242), .ZN(n7961) );
  NAND2_X1 U9288 ( .A1(n8419), .A2(n7773), .ZN(n7960) );
  NAND2_X1 U9289 ( .A1(n8414), .A2(n8008), .ZN(n7969) );
  INV_X1 U9290 ( .A(n8193), .ZN(n7963) );
  INV_X1 U9291 ( .A(n8414), .ZN(n8204) );
  NAND2_X1 U9292 ( .A1(n8402), .A2(n8006), .ZN(n7834) );
  INV_X1 U9293 ( .A(n8157), .ZN(n8166) );
  NOR2_X1 U9294 ( .A1(n8397), .A2(n8168), .ZN(n7797) );
  INV_X1 U9295 ( .A(n7797), .ZN(n7977) );
  NAND2_X1 U9296 ( .A1(n8397), .A2(n8168), .ZN(n7983) );
  NAND2_X1 U9297 ( .A1(n7977), .A2(n7983), .ZN(n7839) );
  NAND2_X1 U9298 ( .A1(n7601), .A2(n7935), .ZN(n8314) );
  OR2_X1 U9299 ( .A1(n8451), .A2(n8296), .ZN(n7947) );
  NAND2_X1 U9300 ( .A1(n8451), .A2(n8296), .ZN(n7934) );
  INV_X1 U9301 ( .A(n7934), .ZN(n7944) );
  XNOR2_X1 U9302 ( .A(n8440), .B(n8297), .ZN(n8275) );
  NAND2_X1 U9303 ( .A1(n8263), .A2(n7953), .ZN(n8240) );
  NAND2_X1 U9304 ( .A1(n8165), .A2(n8157), .ZN(n8171) );
  NAND2_X1 U9305 ( .A1(n8171), .A2(n7835), .ZN(n7798) );
  XNOR2_X1 U9306 ( .A(n7798), .B(n7839), .ZN(n7602) );
  INV_X1 U9307 ( .A(n7602), .ZN(n7610) );
  NAND2_X1 U9308 ( .A1(n7603), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7607) );
  NAND2_X1 U9309 ( .A1(n7604), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7606) );
  NAND2_X1 U9310 ( .A1(n4298), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7605) );
  AND3_X1 U9311 ( .A1(n7607), .A2(n7606), .A3(n7605), .ZN(n8004) );
  INV_X1 U9312 ( .A(n7608), .ZN(n7609) );
  INV_X1 U9313 ( .A(n7611), .ZN(n8400) );
  OAI21_X1 U9314 ( .B1(n7612), .B2(n8218), .A(n8400), .ZN(n7617) );
  NAND2_X1 U9315 ( .A1(n8159), .A2(n8397), .ZN(n7613) );
  INV_X1 U9316 ( .A(n8398), .ZN(n7615) );
  AOI22_X1 U9317 ( .A1(n8397), .A2(n8363), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n8362), .ZN(n7614) );
  OAI21_X1 U9318 ( .B1(n7615), .B2(n8358), .A(n7614), .ZN(n7616) );
  AOI21_X1 U9319 ( .B1(n7617), .B2(n8383), .A(n7616), .ZN(n7618) );
  OAI21_X1 U9320 ( .B1(n8401), .B2(n8321), .A(n7618), .ZN(P2_U3267) );
  INV_X1 U9321 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8622) );
  INV_X1 U9322 ( .A(n8621), .ZN(n8494) );
  OAI222_X1 U9323 ( .A1(n9360), .A2(n8622), .B1(n9364), .B2(n8494), .C1(
        P1_U3084), .C2(n5020), .ZN(P1_U3323) );
  NAND3_X1 U9324 ( .A1(n5738), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n7622) );
  NAND2_X1 U9325 ( .A1(n9354), .A2(n7619), .ZN(n7621) );
  NAND2_X1 U9326 ( .A1(n8491), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7620) );
  OAI211_X1 U9327 ( .C1(n5737), .C2(n7622), .A(n7621), .B(n7620), .ZN(P2_U3327) );
  OAI222_X1 U9328 ( .A1(n9364), .A2(n7623), .B1(P1_U3084), .B2(n9488), .C1(
        n10040), .C2(n9360), .ZN(P1_U3325) );
  OAI222_X1 U9329 ( .A1(n7628), .A2(n7627), .B1(n7626), .B2(n7625), .C1(
        P2_U3152), .C2(n7624), .ZN(P2_U3336) );
  INV_X1 U9330 ( .A(n8407), .ZN(n8180) );
  INV_X1 U9331 ( .A(n7629), .ZN(n7630) );
  NOR3_X1 U9332 ( .A1(n7631), .A2(n8008), .A3(n7772), .ZN(n7633) );
  OAI21_X1 U9333 ( .B1(n7634), .B2(n7633), .A(n7632), .ZN(n7639) );
  NOR2_X1 U9334 ( .A1(n7635), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7637) );
  OAI22_X1 U9335 ( .A1(n8006), .A2(n7790), .B1(n7789), .B2(n8008), .ZN(n7636)
         );
  AOI211_X1 U9336 ( .C1(n7782), .C2(n8178), .A(n7637), .B(n7636), .ZN(n7638)
         );
  OAI211_X1 U9337 ( .C1(n8180), .C2(n9687), .A(n7639), .B(n7638), .ZN(P2_U3216) );
  AOI22_X1 U9338 ( .A1(n7641), .A2(n9674), .B1(n9678), .B2(n7599), .ZN(n7647)
         );
  INV_X1 U9339 ( .A(n8246), .ZN(n7643) );
  OAI22_X1 U9340 ( .A1(n9693), .A2(n7643), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7642), .ZN(n7645) );
  OAI22_X1 U9341 ( .A1(n8242), .A2(n7790), .B1(n7789), .B2(n8278), .ZN(n7644)
         );
  AOI211_X1 U9342 ( .C1(n8427), .C2(n9435), .A(n7645), .B(n7644), .ZN(n7646)
         );
  OAI21_X1 U9343 ( .B1(n7647), .B2(n7720), .A(n7646), .ZN(P2_U3218) );
  XOR2_X1 U9344 ( .A(n7649), .B(n7648), .Z(n7650) );
  NAND2_X1 U9345 ( .A1(n7650), .A2(n9674), .ZN(n7656) );
  AOI22_X1 U9346 ( .A1(n9428), .A2(n7651), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n7655) );
  OR2_X1 U9347 ( .A1(n9687), .A2(n9782), .ZN(n7654) );
  OR2_X1 U9348 ( .A1(n9693), .A2(n7652), .ZN(n7653) );
  NAND4_X1 U9349 ( .A1(n7656), .A2(n7655), .A3(n7654), .A4(n7653), .ZN(
        P2_U3219) );
  NAND2_X1 U9350 ( .A1(n4309), .A2(n7657), .ZN(n7711) );
  NAND2_X1 U9351 ( .A1(n7711), .A2(n7658), .ZN(n7666) );
  AND2_X1 U9352 ( .A1(n7666), .A2(n7659), .ZN(n7762) );
  INV_X1 U9353 ( .A(n7762), .ZN(n7662) );
  NOR3_X1 U9354 ( .A1(n7660), .A2(n7714), .A3(n7772), .ZN(n7661) );
  AOI21_X1 U9355 ( .B1(n7662), .B2(n9674), .A(n7661), .ZN(n7672) );
  OR2_X1 U9356 ( .A1(n8372), .A2(n7714), .ZN(n7663) );
  OAI21_X1 U9357 ( .B1(n8371), .B2(n8277), .A(n7663), .ZN(n8315) );
  AOI22_X1 U9358 ( .A1(n9428), .A2(n8315), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n7664) );
  OAI21_X1 U9359 ( .B1(n8308), .B2(n9693), .A(n7664), .ZN(n7669) );
  NAND2_X1 U9360 ( .A1(n7666), .A2(n7665), .ZN(n7667) );
  NOR2_X1 U9361 ( .A1(n7667), .A2(n9431), .ZN(n7668) );
  AOI211_X1 U9362 ( .C1(n9435), .C2(n8451), .A(n7669), .B(n7668), .ZN(n7670)
         );
  OAI21_X1 U9363 ( .B1(n7672), .B2(n7671), .A(n7670), .ZN(P2_U3221) );
  AOI22_X1 U9364 ( .A1(n9684), .A2(n8027), .B1(n9682), .B2(n8025), .ZN(n7680)
         );
  AOI22_X1 U9365 ( .A1(n9435), .A2(n7673), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n7750), .ZN(n7679) );
  OAI21_X1 U9366 ( .B1(n7676), .B2(n7675), .A(n7674), .ZN(n7677) );
  NAND2_X1 U9367 ( .A1(n7677), .A2(n9674), .ZN(n7678) );
  NAND3_X1 U9368 ( .A1(n7680), .A2(n7679), .A3(n7678), .ZN(P2_U3224) );
  NAND2_X1 U9369 ( .A1(n4309), .A2(n7681), .ZN(n7732) );
  NAND2_X1 U9370 ( .A1(n7732), .A2(n7682), .ZN(n7735) );
  AOI21_X1 U9371 ( .B1(n7735), .B2(n4355), .A(n9431), .ZN(n7685) );
  NOR3_X1 U9372 ( .A1(n7683), .A2(n8277), .A3(n7772), .ZN(n7684) );
  OAI21_X1 U9373 ( .B1(n7685), .B2(n7684), .A(n6096), .ZN(n7690) );
  NOR2_X1 U9374 ( .A1(n7686), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7688) );
  OAI22_X1 U9375 ( .A1(n8277), .A2(n7789), .B1(n7790), .B2(n8278), .ZN(n7687)
         );
  AOI211_X1 U9376 ( .C1(n7782), .C2(n8281), .A(n7688), .B(n7687), .ZN(n7689)
         );
  OAI211_X1 U9377 ( .C1(n7595), .C2(n9687), .A(n7690), .B(n7689), .ZN(P2_U3225) );
  OAI211_X1 U9378 ( .C1(n7692), .C2(n7691), .A(n7776), .B(n9674), .ZN(n7696)
         );
  OAI22_X1 U9379 ( .A1(n8008), .A2(n8371), .B1(n8242), .B2(n8372), .ZN(n8212)
         );
  AOI22_X1 U9380 ( .A1(n9428), .A2(n8212), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n7693) );
  OAI21_X1 U9381 ( .B1(n8217), .B2(n9693), .A(n7693), .ZN(n7694) );
  INV_X1 U9382 ( .A(n7694), .ZN(n7695) );
  OAI211_X1 U9383 ( .C1(n7697), .C2(n9687), .A(n7696), .B(n7695), .ZN(P2_U3227) );
  INV_X1 U9384 ( .A(n7699), .ZN(n7701) );
  XNOR2_X1 U9385 ( .A(n7698), .B(n7699), .ZN(n7785) );
  NAND2_X1 U9386 ( .A1(n7785), .A2(n7700), .ZN(n7786) );
  OAI21_X1 U9387 ( .B1(n7701), .B2(n7698), .A(n7786), .ZN(n7705) );
  XNOR2_X1 U9388 ( .A(n7703), .B(n7702), .ZN(n7704) );
  XNOR2_X1 U9389 ( .A(n7705), .B(n7704), .ZN(n7710) );
  INV_X1 U9390 ( .A(n8354), .ZN(n7706) );
  NAND2_X1 U9391 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8088) );
  OAI21_X1 U9392 ( .B1(n9693), .B2(n7706), .A(n8088), .ZN(n7708) );
  OAI22_X1 U9393 ( .A1(n8344), .A2(n7789), .B1(n7790), .B2(n8343), .ZN(n7707)
         );
  AOI211_X1 U9394 ( .C1(n9435), .C2(n8355), .A(n7708), .B(n7707), .ZN(n7709)
         );
  OAI21_X1 U9395 ( .B1(n7710), .B2(n9431), .A(n7709), .ZN(P2_U3228) );
  NAND2_X1 U9396 ( .A1(n7711), .A2(n7712), .ZN(n7760) );
  OAI211_X1 U9397 ( .C1(n7712), .C2(n7711), .A(n7760), .B(n9674), .ZN(n7717)
         );
  NOR2_X1 U9398 ( .A1(n7713), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8106) );
  OAI22_X1 U9399 ( .A1(n7714), .A2(n7790), .B1(n7789), .B2(n8331), .ZN(n7715)
         );
  AOI211_X1 U9400 ( .C1(n7782), .C2(n8334), .A(n8106), .B(n7715), .ZN(n7716)
         );
  OAI211_X1 U9401 ( .C1(n7718), .C2(n9687), .A(n7717), .B(n7716), .ZN(P2_U3230) );
  NOR2_X1 U9402 ( .A1(n7720), .A2(n7719), .ZN(n7722) );
  XNOR2_X1 U9403 ( .A(n7722), .B(n7721), .ZN(n7725) );
  OAI22_X1 U9404 ( .A1(n7725), .A2(n9431), .B1(n8242), .B2(n7772), .ZN(n7723)
         );
  OAI21_X1 U9405 ( .B1(n7725), .B2(n7724), .A(n7723), .ZN(n7730) );
  NOR2_X1 U9406 ( .A1(n7726), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7728) );
  OAI22_X1 U9407 ( .A1(n7745), .A2(n7789), .B1(n7790), .B2(n7773), .ZN(n7727)
         );
  AOI211_X1 U9408 ( .C1(n7782), .C2(n8227), .A(n7728), .B(n7727), .ZN(n7729)
         );
  OAI211_X1 U9409 ( .C1(n8229), .C2(n9687), .A(n7730), .B(n7729), .ZN(P2_U3231) );
  NAND2_X1 U9410 ( .A1(n7732), .A2(n7731), .ZN(n7734) );
  AOI21_X1 U9411 ( .B1(n7734), .B2(n7733), .A(n9431), .ZN(n7736) );
  NAND2_X1 U9412 ( .A1(n7736), .A2(n7735), .ZN(n7740) );
  NOR2_X1 U9413 ( .A1(n9693), .A2(n8288), .ZN(n7738) );
  OAI22_X1 U9414 ( .A1(n8297), .A2(n7790), .B1(n7789), .B2(n8296), .ZN(n7737)
         );
  AOI211_X1 U9415 ( .C1(P2_REG3_REG_20__SCAN_IN), .C2(P2_U3152), .A(n7738), 
        .B(n7737), .ZN(n7739) );
  OAI211_X1 U9416 ( .C1(n8291), .C2(n9687), .A(n7740), .B(n7739), .ZN(P2_U3235) );
  NAND2_X1 U9417 ( .A1(n9678), .A2(n7597), .ZN(n7744) );
  NAND2_X1 U9418 ( .A1(n9674), .A2(n7741), .ZN(n7743) );
  MUX2_X1 U9419 ( .A(n7744), .B(n7743), .S(n7742), .Z(n7749) );
  NOR2_X1 U9420 ( .A1(n9693), .A2(n8259), .ZN(n7747) );
  OAI22_X1 U9421 ( .A1(n7745), .A2(n7790), .B1(n7789), .B2(n8297), .ZN(n7746)
         );
  AOI211_X1 U9422 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3152), .A(n7747), 
        .B(n7746), .ZN(n7748) );
  OAI211_X1 U9423 ( .C1(n8262), .C2(n9687), .A(n7749), .B(n7748), .ZN(P2_U3237) );
  AOI22_X1 U9424 ( .A1(n9682), .A2(n8024), .B1(n9684), .B2(n7184), .ZN(n7758)
         );
  AOI22_X1 U9425 ( .A1(n9435), .A2(n7751), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n7750), .ZN(n7757) );
  AOI21_X1 U9426 ( .B1(n7753), .B2(n7752), .A(n9431), .ZN(n7755) );
  NAND2_X1 U9427 ( .A1(n7755), .A2(n7754), .ZN(n7756) );
  NAND3_X1 U9428 ( .A1(n7758), .A2(n7757), .A3(n7756), .ZN(P2_U3239) );
  AOI21_X1 U9429 ( .B1(n7760), .B2(n7759), .A(n9431), .ZN(n7764) );
  NOR3_X1 U9430 ( .A1(n7761), .A2(n8343), .A3(n7772), .ZN(n7763) );
  OAI21_X1 U9431 ( .B1(n7764), .B2(n7763), .A(n7762), .ZN(n7770) );
  INV_X1 U9432 ( .A(n9428), .ZN(n7780) );
  INV_X1 U9433 ( .A(n7765), .ZN(n7766) );
  NAND2_X1 U9434 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8127) );
  OAI21_X1 U9435 ( .B1(n7780), .B2(n7766), .A(n8127), .ZN(n7767) );
  AOI21_X1 U9436 ( .B1(n7768), .B2(n7782), .A(n7767), .ZN(n7769) );
  OAI211_X1 U9437 ( .C1(n7771), .C2(n9687), .A(n7770), .B(n7769), .ZN(P2_U3240) );
  NOR3_X1 U9438 ( .A1(n7774), .A2(n7773), .A3(n7772), .ZN(n7778) );
  AOI21_X1 U9439 ( .B1(n7776), .B2(n7775), .A(n9431), .ZN(n7777) );
  OAI21_X1 U9440 ( .B1(n7778), .B2(n7777), .A(n4310), .ZN(n7784) );
  INV_X1 U9441 ( .A(n7779), .ZN(n8201) );
  AOI22_X1 U9442 ( .A1(n8007), .A2(n8328), .B1(n8233), .B2(n8266), .ZN(n8197)
         );
  OAI22_X1 U9443 ( .A1(n7780), .A2(n8197), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9948), .ZN(n7781) );
  AOI21_X1 U9444 ( .B1(n8201), .B2(n7782), .A(n7781), .ZN(n7783) );
  OAI211_X1 U9445 ( .C1(n8204), .C2(n9687), .A(n7784), .B(n7783), .ZN(P2_U3242) );
  AOI22_X1 U9446 ( .A1(n7785), .A2(n9674), .B1(n9678), .B2(n8014), .ZN(n7796)
         );
  INV_X1 U9447 ( .A(n7786), .ZN(n7795) );
  OAI22_X1 U9448 ( .A1(n9693), .A2(n7787), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9938), .ZN(n7792) );
  OAI22_X1 U9449 ( .A1(n8331), .A2(n7790), .B1(n7789), .B2(n7788), .ZN(n7791)
         );
  AOI211_X1 U9450 ( .C1(n9435), .C2(n7793), .A(n7792), .B(n7791), .ZN(n7794)
         );
  OAI21_X1 U9451 ( .B1(n7796), .B2(n7795), .A(n7794), .ZN(P2_U3243) );
  INV_X1 U9452 ( .A(n7802), .ZN(n7800) );
  NOR2_X1 U9453 ( .A1(n8152), .A2(n8004), .ZN(n7810) );
  OAI22_X1 U9454 ( .A1(n7800), .A2(n7810), .B1(n7799), .B2(n7803), .ZN(n7801)
         );
  OAI21_X1 U9455 ( .B1(n7802), .B2(n8152), .A(n7801), .ZN(n7806) );
  INV_X1 U9456 ( .A(n7803), .ZN(n7804) );
  NAND2_X1 U9457 ( .A1(n8152), .A2(n8004), .ZN(n7984) );
  XNOR2_X1 U9458 ( .A(n7807), .B(n8395), .ZN(n7996) );
  NAND2_X1 U9459 ( .A1(n7809), .A2(n7808), .ZN(n7995) );
  INV_X1 U9460 ( .A(n7810), .ZN(n7978) );
  INV_X1 U9461 ( .A(n8231), .ZN(n7830) );
  INV_X1 U9462 ( .A(n8313), .ZN(n7826) );
  INV_X1 U9463 ( .A(n8325), .ZN(n8322) );
  NOR3_X1 U9464 ( .A1(n7857), .A2(n7812), .A3(n7201), .ZN(n7813) );
  AND2_X1 U9465 ( .A1(n7855), .A2(n7853), .ZN(n7840) );
  NAND4_X1 U9466 ( .A1(n7860), .A2(n8394), .A3(n7813), .A4(n7840), .ZN(n7816)
         );
  NOR4_X1 U9467 ( .A1(n7816), .A2(n7877), .A3(n7815), .A4(n7814), .ZN(n7818)
         );
  NAND4_X1 U9468 ( .A1(n7818), .A2(n7885), .A3(n7884), .A4(n4748), .ZN(n7821)
         );
  NOR4_X1 U9469 ( .A1(n7343), .A2(n7821), .A3(n7820), .A4(n7819), .ZN(n7823)
         );
  NAND4_X1 U9470 ( .A1(n8341), .A2(n7919), .A3(n7823), .A4(n7822), .ZN(n7824)
         );
  NOR4_X1 U9471 ( .A1(n7826), .A2(n7825), .A3(n8322), .A4(n7824), .ZN(n7828)
         );
  INV_X1 U9472 ( .A(n8275), .ZN(n7827) );
  NAND4_X1 U9473 ( .A1(n8264), .A2(n8293), .A3(n7828), .A4(n7827), .ZN(n7829)
         );
  NOR4_X1 U9474 ( .A1(n8207), .A2(n7830), .A3(n8250), .A4(n7829), .ZN(n7831)
         );
  NAND4_X1 U9475 ( .A1(n8157), .A2(n8193), .A3(n7831), .A4(n8182), .ZN(n7832)
         );
  INV_X1 U9476 ( .A(n7834), .ZN(n7837) );
  INV_X1 U9477 ( .A(n7835), .ZN(n7836) );
  MUX2_X1 U9478 ( .A(n7837), .B(n7836), .S(n7986), .Z(n7838) );
  NOR2_X1 U9479 ( .A1(n7839), .A2(n7838), .ZN(n7976) );
  INV_X1 U9480 ( .A(n7840), .ZN(n7842) );
  NAND3_X1 U9481 ( .A1(n7842), .A2(n8374), .A3(n7841), .ZN(n7843) );
  NAND2_X1 U9482 ( .A1(n7843), .A2(n7854), .ZN(n7863) );
  AND2_X1 U9483 ( .A1(n7846), .A2(n7844), .ZN(n7847) );
  AND2_X1 U9484 ( .A1(n4844), .A2(n7865), .ZN(n7845) );
  MUX2_X1 U9485 ( .A(n7847), .B(n7845), .S(n7986), .Z(n7864) );
  INV_X1 U9486 ( .A(n7846), .ZN(n7850) );
  INV_X1 U9487 ( .A(n7847), .ZN(n7848) );
  OAI22_X1 U9488 ( .A1(n7864), .A2(n7850), .B1(n7849), .B2(n7848), .ZN(n7851)
         );
  NAND2_X1 U9489 ( .A1(n7851), .A2(n7871), .ZN(n7852) );
  NAND2_X1 U9490 ( .A1(n7852), .A2(n7986), .ZN(n7862) );
  AND2_X1 U9491 ( .A1(n7853), .A2(n5719), .ZN(n7856) );
  OAI211_X1 U9492 ( .C1(n7857), .C2(n7856), .A(n7855), .B(n7854), .ZN(n7858)
         );
  NAND3_X1 U9493 ( .A1(n7858), .A2(n7986), .A3(n8374), .ZN(n7859) );
  NAND3_X1 U9494 ( .A1(n7864), .A2(n7860), .A3(n7859), .ZN(n7861) );
  INV_X1 U9495 ( .A(n7864), .ZN(n7869) );
  AND2_X1 U9496 ( .A1(n7866), .A2(n7865), .ZN(n7868) );
  OAI211_X1 U9497 ( .C1(n7869), .C2(n7868), .A(n4844), .B(n7867), .ZN(n7870)
         );
  NAND2_X1 U9498 ( .A1(n7870), .A2(n7989), .ZN(n7873) );
  OAI21_X1 U9499 ( .B1(n7986), .B2(n7871), .A(n4748), .ZN(n7872) );
  AND2_X1 U9500 ( .A1(n7986), .A2(n7874), .ZN(n7876) );
  NOR2_X1 U9501 ( .A1(n7986), .A2(n7874), .ZN(n7875) );
  MUX2_X1 U9502 ( .A(n7876), .B(n7875), .S(n9683), .Z(n7878) );
  MUX2_X1 U9503 ( .A(n7880), .B(n7879), .S(n7986), .Z(n7882) );
  AND2_X1 U9504 ( .A1(n7882), .A2(n7881), .ZN(n7887) );
  NOR2_X1 U9505 ( .A1(n7986), .A2(n7272), .ZN(n7883) );
  AOI22_X1 U9506 ( .A1(n7885), .A2(n7884), .B1(n7883), .B2(n7890), .ZN(n7886)
         );
  AOI21_X1 U9507 ( .B1(n7888), .B2(n7887), .A(n7886), .ZN(n7897) );
  NAND2_X1 U9508 ( .A1(n7898), .A2(n7889), .ZN(n7895) );
  INV_X1 U9509 ( .A(n7889), .ZN(n7893) );
  OAI211_X1 U9510 ( .C1(n7893), .C2(n7892), .A(n7891), .B(n7890), .ZN(n7894)
         );
  MUX2_X1 U9511 ( .A(n7895), .B(n7894), .S(n7986), .Z(n7896) );
  OR2_X1 U9512 ( .A1(n7897), .A2(n7896), .ZN(n7902) );
  NAND2_X1 U9513 ( .A1(n7902), .A2(n7898), .ZN(n7901) );
  AOI21_X1 U9514 ( .B1(n7901), .B2(n7900), .A(n7899), .ZN(n7908) );
  INV_X1 U9515 ( .A(n7902), .ZN(n7906) );
  INV_X1 U9516 ( .A(n7903), .ZN(n7905) );
  OAI21_X1 U9517 ( .B1(n7906), .B2(n7905), .A(n7904), .ZN(n7907) );
  MUX2_X1 U9518 ( .A(n7908), .B(n7907), .S(n7989), .Z(n7915) );
  INV_X1 U9519 ( .A(n7909), .ZN(n7910) );
  MUX2_X1 U9520 ( .A(n7911), .B(n7910), .S(n7989), .Z(n7912) );
  NOR2_X1 U9521 ( .A1(n7913), .A2(n7912), .ZN(n7914) );
  NAND2_X1 U9522 ( .A1(n7986), .A2(n8015), .ZN(n7917) );
  OR2_X1 U9523 ( .A1(n7986), .A2(n8015), .ZN(n7916) );
  MUX2_X1 U9524 ( .A(n7917), .B(n7916), .S(n9449), .Z(n7918) );
  MUX2_X1 U9525 ( .A(n7922), .B(n7921), .S(n7986), .Z(n7923) );
  AND2_X1 U9526 ( .A1(n8325), .A2(n7923), .ZN(n7925) );
  NAND2_X1 U9527 ( .A1(n7924), .A2(n7925), .ZN(n7933) );
  INV_X1 U9528 ( .A(n7925), .ZN(n7928) );
  NAND2_X1 U9529 ( .A1(n8462), .A2(n8343), .ZN(n7926) );
  OAI211_X1 U9530 ( .C1(n7928), .C2(n7927), .A(n7935), .B(n7926), .ZN(n7929)
         );
  MUX2_X1 U9531 ( .A(n7930), .B(n7929), .S(n7989), .Z(n7931) );
  INV_X1 U9532 ( .A(n7931), .ZN(n7932) );
  NAND3_X1 U9533 ( .A1(n7933), .A2(n7932), .A3(n7945), .ZN(n7946) );
  NAND3_X1 U9534 ( .A1(n7946), .A2(n7935), .A3(n7934), .ZN(n7937) );
  INV_X1 U9535 ( .A(n7949), .ZN(n7936) );
  AOI21_X1 U9536 ( .B1(n7937), .B2(n7947), .A(n7936), .ZN(n7939) );
  OR2_X1 U9537 ( .A1(n8440), .A2(n8297), .ZN(n7952) );
  NAND2_X1 U9538 ( .A1(n7952), .A2(n7948), .ZN(n7938) );
  OAI211_X1 U9539 ( .C1(n7939), .C2(n7938), .A(n7986), .B(n4308), .ZN(n7941)
         );
  INV_X1 U9540 ( .A(n8250), .ZN(n7942) );
  AOI21_X1 U9541 ( .B1(n7946), .B2(n7945), .A(n7944), .ZN(n7951) );
  NAND2_X1 U9542 ( .A1(n7948), .A2(n7947), .ZN(n7950) );
  OAI211_X1 U9543 ( .C1(n7951), .C2(n7950), .A(n7949), .B(n4308), .ZN(n7954)
         );
  NAND4_X1 U9544 ( .A1(n7954), .A2(n7989), .A3(n7953), .A4(n7952), .ZN(n7955)
         );
  NAND2_X1 U9545 ( .A1(n7955), .A2(n7958), .ZN(n7956) );
  AOI21_X1 U9546 ( .B1(n7958), .B2(n7957), .A(n7986), .ZN(n7959) );
  OAI21_X1 U9547 ( .B1(n8207), .B2(n7961), .A(n7960), .ZN(n7962) );
  OAI21_X1 U9548 ( .B1(n7963), .B2(n7962), .A(n7986), .ZN(n7964) );
  NAND2_X1 U9549 ( .A1(n7965), .A2(n7964), .ZN(n7968) );
  AOI21_X1 U9550 ( .B1(n7967), .B2(n8194), .A(n7986), .ZN(n7966) );
  AOI21_X1 U9551 ( .B1(n7968), .B2(n7967), .A(n7966), .ZN(n7974) );
  OAI21_X1 U9552 ( .B1(n7969), .B2(n7986), .A(n8182), .ZN(n7973) );
  NAND2_X1 U9553 ( .A1(n8007), .A2(n7989), .ZN(n7971) );
  OR2_X1 U9554 ( .A1(n8007), .A2(n7989), .ZN(n7970) );
  MUX2_X1 U9555 ( .A(n7971), .B(n7970), .S(n8407), .Z(n7972) );
  OAI211_X1 U9556 ( .C1(n7974), .C2(n7973), .A(n8157), .B(n7972), .ZN(n7975)
         );
  NAND2_X1 U9557 ( .A1(n7976), .A2(n7975), .ZN(n7982) );
  NAND3_X1 U9558 ( .A1(n7978), .A2(n7977), .A3(n7982), .ZN(n7980) );
  NAND3_X1 U9559 ( .A1(n7984), .A2(n7983), .A3(n7982), .ZN(n7985) );
  NAND2_X1 U9560 ( .A1(n4348), .A2(n7985), .ZN(n7987) );
  INV_X1 U9561 ( .A(n7990), .ZN(n7991) );
  NAND2_X1 U9562 ( .A1(n4843), .A2(n7991), .ZN(n7992) );
  NOR4_X1 U9563 ( .A1(n7999), .A2(n7998), .A3(n7997), .A4(n8372), .ZN(n8001)
         );
  OAI21_X1 U9564 ( .B1(n8002), .B2(n6212), .A(P2_B_REG_SCAN_IN), .ZN(n8000) );
  OAI22_X1 U9565 ( .A1(n8003), .A2(n8002), .B1(n8001), .B2(n8000), .ZN(
        P2_U3244) );
  INV_X1 U9566 ( .A(n8004), .ZN(n8005) );
  MUX2_X1 U9567 ( .A(n8005), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8026), .Z(
        P2_U3582) );
  INV_X1 U9568 ( .A(n8006), .ZN(n8185) );
  MUX2_X1 U9569 ( .A(n8185), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8026), .Z(
        P2_U3580) );
  MUX2_X1 U9570 ( .A(n8007), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8026), .Z(
        P2_U3579) );
  INV_X1 U9571 ( .A(n8008), .ZN(n8184) );
  MUX2_X1 U9572 ( .A(n8184), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8026), .Z(
        P2_U3578) );
  MUX2_X1 U9573 ( .A(n8233), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8026), .Z(
        P2_U3577) );
  MUX2_X1 U9574 ( .A(n8009), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8026), .Z(
        P2_U3576) );
  MUX2_X1 U9575 ( .A(n7599), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8026), .Z(
        P2_U3575) );
  MUX2_X1 U9576 ( .A(n7597), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8026), .Z(
        P2_U3574) );
  MUX2_X1 U9577 ( .A(n8265), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8026), .Z(
        P2_U3573) );
  MUX2_X1 U9578 ( .A(n8010), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8026), .Z(
        P2_U3572) );
  MUX2_X1 U9579 ( .A(n8011), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8026), .Z(
        P2_U3571) );
  MUX2_X1 U9580 ( .A(n8327), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8026), .Z(
        P2_U3570) );
  MUX2_X1 U9581 ( .A(n8012), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8026), .Z(
        P2_U3569) );
  MUX2_X1 U9582 ( .A(n8013), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8026), .Z(
        P2_U3568) );
  MUX2_X1 U9583 ( .A(n8014), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8026), .Z(
        P2_U3567) );
  MUX2_X1 U9584 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8015), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9585 ( .A(n8016), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8026), .Z(
        P2_U3565) );
  MUX2_X1 U9586 ( .A(n8017), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8026), .Z(
        P2_U3564) );
  MUX2_X1 U9587 ( .A(n8018), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8026), .Z(
        P2_U3563) );
  MUX2_X1 U9588 ( .A(n8019), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8026), .Z(
        P2_U3562) );
  MUX2_X1 U9589 ( .A(n9681), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8026), .Z(
        P2_U3561) );
  MUX2_X1 U9590 ( .A(n8020), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8026), .Z(
        P2_U3560) );
  MUX2_X1 U9591 ( .A(n9683), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8026), .Z(
        P2_U3559) );
  MUX2_X1 U9592 ( .A(n8021), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8026), .Z(
        P2_U3558) );
  MUX2_X1 U9593 ( .A(n8022), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8026), .Z(
        P2_U3557) );
  MUX2_X1 U9594 ( .A(n8023), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8026), .Z(
        P2_U3556) );
  MUX2_X1 U9595 ( .A(n8024), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8026), .Z(
        P2_U3555) );
  MUX2_X1 U9596 ( .A(n8025), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8026), .Z(
        P2_U3554) );
  MUX2_X1 U9597 ( .A(n7184), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8026), .Z(
        P2_U3553) );
  MUX2_X1 U9598 ( .A(n8027), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8026), .Z(
        P2_U3552) );
  OAI211_X1 U9599 ( .C1(n8030), .C2(n8029), .A(n9695), .B(n8028), .ZN(n8040)
         );
  NOR2_X1 U9600 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8368), .ZN(n8031) );
  AOI21_X1 U9601 ( .B1(n9697), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n8031), .ZN(
        n8039) );
  OR2_X1 U9602 ( .A1(n9699), .A2(n8032), .ZN(n8038) );
  AOI21_X1 U9603 ( .B1(n8035), .B2(n8034), .A(n8033), .ZN(n8036) );
  NAND2_X1 U9604 ( .A1(n9694), .A2(n8036), .ZN(n8037) );
  NAND4_X1 U9605 ( .A1(n8040), .A2(n8039), .A3(n8038), .A4(n8037), .ZN(
        P2_U3248) );
  OAI211_X1 U9606 ( .C1(n8043), .C2(n8042), .A(n9695), .B(n8041), .ZN(n8054)
         );
  INV_X1 U9607 ( .A(n8044), .ZN(n8045) );
  AOI21_X1 U9608 ( .B1(n9697), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n8045), .ZN(
        n8053) );
  OR2_X1 U9609 ( .A1(n9699), .A2(n8046), .ZN(n8052) );
  AOI21_X1 U9610 ( .B1(n8049), .B2(n8048), .A(n8047), .ZN(n8050) );
  NAND2_X1 U9611 ( .A1(n9694), .A2(n8050), .ZN(n8051) );
  NAND4_X1 U9612 ( .A1(n8054), .A2(n8053), .A3(n8052), .A4(n8051), .ZN(
        P2_U3249) );
  OAI211_X1 U9613 ( .C1(n8057), .C2(n8056), .A(n9695), .B(n8055), .ZN(n8068)
         );
  NOR2_X1 U9614 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8058), .ZN(n8059) );
  AOI21_X1 U9615 ( .B1(n9697), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8059), .ZN(
        n8067) );
  OR2_X1 U9616 ( .A1(n9699), .A2(n8060), .ZN(n8066) );
  AOI21_X1 U9617 ( .B1(n8063), .B2(n8062), .A(n8061), .ZN(n8064) );
  NAND2_X1 U9618 ( .A1(n9694), .A2(n8064), .ZN(n8065) );
  NAND4_X1 U9619 ( .A1(n8068), .A2(n8067), .A3(n8066), .A4(n8065), .ZN(
        P2_U3250) );
  NOR2_X1 U9620 ( .A1(n8073), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8070) );
  NOR2_X1 U9621 ( .A1(n8070), .A2(n8069), .ZN(n8090) );
  XNOR2_X1 U9622 ( .A(n8090), .B(n8091), .ZN(n8071) );
  NOR2_X1 U9623 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n8071), .ZN(n8092) );
  AOI21_X1 U9624 ( .B1(n8071), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8092), .ZN(
        n8080) );
  INV_X1 U9625 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9448) );
  AOI211_X1 U9626 ( .C1(n8074), .C2(n9448), .A(n8083), .B(n9700), .ZN(n8078)
         );
  NOR2_X1 U9627 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9938), .ZN(n8075) );
  AOI21_X1 U9628 ( .B1(n9697), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8075), .ZN(
        n8076) );
  OAI21_X1 U9629 ( .B1(n9699), .B2(n8082), .A(n8076), .ZN(n8077) );
  NOR2_X1 U9630 ( .A1(n8078), .A2(n8077), .ZN(n8079) );
  OAI21_X1 U9631 ( .B1(n8080), .B2(n9698), .A(n8079), .ZN(P2_U3260) );
  NOR2_X1 U9632 ( .A1(n8082), .A2(n8081), .ZN(n8084) );
  XOR2_X1 U9633 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8107), .Z(n8085) );
  NAND2_X1 U9634 ( .A1(n8085), .A2(n8086), .ZN(n8108) );
  OAI21_X1 U9635 ( .B1(n8086), .B2(n8085), .A(n8108), .ZN(n8087) );
  NAND2_X1 U9636 ( .A1(n8087), .A2(n9694), .ZN(n8101) );
  INV_X1 U9637 ( .A(n8088), .ZN(n8089) );
  AOI21_X1 U9638 ( .B1(n9697), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8089), .ZN(
        n8100) );
  NOR2_X1 U9639 ( .A1(n8091), .A2(n8090), .ZN(n8093) );
  NOR2_X1 U9640 ( .A1(n8093), .A2(n8092), .ZN(n8097) );
  INV_X1 U9641 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8094) );
  MUX2_X1 U9642 ( .A(n8094), .B(P2_REG2_REG_16__SCAN_IN), .S(n8107), .Z(n8095)
         );
  INV_X1 U9643 ( .A(n8095), .ZN(n8096) );
  NAND2_X1 U9644 ( .A1(n8096), .A2(n8097), .ZN(n8102) );
  OAI211_X1 U9645 ( .C1(n8097), .C2(n8096), .A(n9695), .B(n8102), .ZN(n8099)
         );
  INV_X1 U9646 ( .A(n9699), .ZN(n9382) );
  NAND2_X1 U9647 ( .A1(n9382), .A2(n8107), .ZN(n8098) );
  NAND4_X1 U9648 ( .A1(n8101), .A2(n8100), .A3(n8099), .A4(n8098), .ZN(
        P2_U3261) );
  NAND2_X1 U9649 ( .A1(n8107), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8103) );
  NAND2_X1 U9650 ( .A1(n8103), .A2(n8102), .ZN(n8105) );
  XNOR2_X1 U9651 ( .A(n8118), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n8104) );
  NAND2_X1 U9652 ( .A1(n8104), .A2(n8105), .ZN(n8117) );
  OAI211_X1 U9653 ( .C1(n8105), .C2(n8104), .A(n9695), .B(n8117), .ZN(n8116)
         );
  AOI21_X1 U9654 ( .B1(n9697), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8106), .ZN(
        n8115) );
  OR2_X1 U9655 ( .A1(n9699), .A2(n8118), .ZN(n8114) );
  XNOR2_X1 U9656 ( .A(n8122), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8111) );
  OR2_X1 U9657 ( .A1(n8107), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U9658 ( .A1(n8109), .A2(n8108), .ZN(n8110) );
  NOR2_X1 U9659 ( .A1(n8111), .A2(n8110), .ZN(n8121) );
  AOI21_X1 U9660 ( .B1(n8111), .B2(n8110), .A(n8121), .ZN(n8112) );
  NAND2_X1 U9661 ( .A1(n9694), .A2(n8112), .ZN(n8113) );
  NAND4_X1 U9662 ( .A1(n8116), .A2(n8115), .A3(n8114), .A4(n8113), .ZN(
        P2_U3262) );
  INV_X1 U9663 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8119) );
  OAI21_X1 U9664 ( .B1(n8119), .B2(n8118), .A(n8117), .ZN(n8133) );
  XNOR2_X1 U9665 ( .A(n8138), .B(n8133), .ZN(n8120) );
  NOR2_X1 U9666 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8120), .ZN(n8134) );
  AOI21_X1 U9667 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8120), .A(n8134), .ZN(
        n8132) );
  INV_X1 U9668 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8123) );
  AOI22_X1 U9669 ( .A1(n8138), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n8123), .B2(
        n8128), .ZN(n8124) );
  OAI21_X1 U9670 ( .B1(n8125), .B2(n8124), .A(n8137), .ZN(n8130) );
  NAND2_X1 U9671 ( .A1(n9697), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n8126) );
  OAI211_X1 U9672 ( .C1(n9699), .C2(n8128), .A(n8127), .B(n8126), .ZN(n8129)
         );
  AOI21_X1 U9673 ( .B1(n8130), .B2(n9694), .A(n8129), .ZN(n8131) );
  OAI21_X1 U9674 ( .B1(n8132), .B2(n9698), .A(n8131), .ZN(P2_U3263) );
  NOR2_X1 U9675 ( .A1(n8138), .A2(n8133), .ZN(n8135) );
  NOR2_X1 U9676 ( .A1(n8135), .A2(n8134), .ZN(n8136) );
  XOR2_X1 U9677 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8136), .Z(n8145) );
  INV_X1 U9678 ( .A(n8144), .ZN(n8140) );
  NAND2_X1 U9679 ( .A1(n8140), .A2(n9694), .ZN(n8141) );
  OAI211_X1 U9680 ( .C1(n8145), .C2(n8142), .A(n9699), .B(n8141), .ZN(n8143)
         );
  INV_X1 U9681 ( .A(n8143), .ZN(n8147) );
  AOI22_X1 U9682 ( .A1(n8145), .A2(n9695), .B1(n9694), .B2(n8144), .ZN(n8146)
         );
  MUX2_X1 U9683 ( .A(n8147), .B(n8146), .S(n8395), .Z(n8149) );
  NAND2_X1 U9684 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8148) );
  OAI211_X1 U9685 ( .C1(n8151), .C2(n8150), .A(n8149), .B(n8148), .ZN(P2_U3264) );
  XOR2_X1 U9686 ( .A(n8153), .B(n8152), .Z(n9441) );
  NAND2_X1 U9687 ( .A1(n9441), .A2(n8370), .ZN(n8156) );
  AOI21_X1 U9688 ( .B1(n8362), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8154), .ZN(
        n8155) );
  OAI211_X1 U9689 ( .C1(n4436), .C2(n8311), .A(n8156), .B(n8155), .ZN(P2_U3266) );
  XNOR2_X1 U9690 ( .A(n8158), .B(n8157), .ZN(n8406) );
  INV_X1 U9691 ( .A(n8177), .ZN(n8161) );
  INV_X1 U9692 ( .A(n8159), .ZN(n8160) );
  AOI21_X1 U9693 ( .B1(n8402), .B2(n8161), .A(n8160), .ZN(n8403) );
  AOI22_X1 U9694 ( .A1(n8362), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8162), .B2(
        n8369), .ZN(n8163) );
  OAI21_X1 U9695 ( .B1(n8164), .B2(n8311), .A(n8163), .ZN(n8174) );
  INV_X1 U9696 ( .A(n8165), .ZN(n8167) );
  AOI21_X1 U9697 ( .B1(n8167), .B2(n8166), .A(n8377), .ZN(n8172) );
  OAI22_X1 U9698 ( .A1(n8169), .A2(n8372), .B1(n8168), .B2(n8371), .ZN(n8170)
         );
  AOI21_X1 U9699 ( .B1(n8172), .B2(n8171), .A(n8170), .ZN(n8405) );
  NOR2_X1 U9700 ( .A1(n8405), .A2(n8362), .ZN(n8173) );
  AOI211_X1 U9701 ( .C1(n8370), .C2(n8403), .A(n8174), .B(n8173), .ZN(n8175)
         );
  OAI21_X1 U9702 ( .B1(n8406), .B2(n8321), .A(n8175), .ZN(P2_U3268) );
  XOR2_X1 U9703 ( .A(n8182), .B(n8176), .Z(n8411) );
  AOI21_X1 U9704 ( .B1(n8407), .B2(n8199), .A(n8177), .ZN(n8408) );
  AOI22_X1 U9705 ( .A1(n8362), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8178), .B2(
        n8369), .ZN(n8179) );
  OAI21_X1 U9706 ( .B1(n8180), .B2(n8311), .A(n8179), .ZN(n8189) );
  OAI211_X1 U9707 ( .C1(n8183), .C2(n8182), .A(n8181), .B(n8351), .ZN(n8187)
         );
  AOI22_X1 U9708 ( .A1(n8185), .A2(n8328), .B1(n8266), .B2(n8184), .ZN(n8186)
         );
  NOR2_X1 U9709 ( .A1(n8410), .A2(n8362), .ZN(n8188) );
  AOI211_X1 U9710 ( .C1(n8370), .C2(n8408), .A(n8189), .B(n8188), .ZN(n8190)
         );
  OAI21_X1 U9711 ( .B1(n8411), .B2(n8321), .A(n8190), .ZN(P2_U3269) );
  XNOR2_X1 U9712 ( .A(n8191), .B(n8193), .ZN(n8416) );
  INV_X1 U9713 ( .A(n8192), .ZN(n8196) );
  AOI21_X1 U9714 ( .B1(n8209), .B2(n8194), .A(n8193), .ZN(n8195) );
  OAI21_X1 U9715 ( .B1(n8196), .B2(n8195), .A(n8351), .ZN(n8198) );
  NAND2_X1 U9716 ( .A1(n8198), .A2(n8197), .ZN(n8412) );
  INV_X1 U9717 ( .A(n8199), .ZN(n8200) );
  AOI211_X1 U9718 ( .C1(n8414), .C2(n8215), .A(n9801), .B(n8200), .ZN(n8413)
         );
  NAND2_X1 U9719 ( .A1(n8413), .A2(n8319), .ZN(n8203) );
  AOI22_X1 U9720 ( .A1(n8362), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8201), .B2(
        n8369), .ZN(n8202) );
  OAI211_X1 U9721 ( .C1(n8204), .C2(n8311), .A(n8203), .B(n8202), .ZN(n8205)
         );
  AOI21_X1 U9722 ( .B1(n8412), .B2(n8383), .A(n8205), .ZN(n8206) );
  OAI21_X1 U9723 ( .B1(n8416), .B2(n8321), .A(n8206), .ZN(P2_U3270) );
  XNOR2_X1 U9724 ( .A(n8208), .B(n8207), .ZN(n8421) );
  AOI22_X1 U9725 ( .A1(n8419), .A2(n8363), .B1(n8362), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8223) );
  OAI211_X1 U9726 ( .C1(n8211), .C2(n8210), .A(n8209), .B(n8351), .ZN(n8214)
         );
  INV_X1 U9727 ( .A(n8212), .ZN(n8213) );
  NAND2_X1 U9728 ( .A1(n8214), .A2(n8213), .ZN(n8417) );
  INV_X1 U9729 ( .A(n8215), .ZN(n8216) );
  AOI211_X1 U9730 ( .C1(n8419), .C2(n4446), .A(n9801), .B(n8216), .ZN(n8418)
         );
  INV_X1 U9731 ( .A(n8418), .ZN(n8220) );
  OAI22_X1 U9732 ( .A1(n8220), .A2(n8219), .B1(n8218), .B2(n8217), .ZN(n8221)
         );
  OAI21_X1 U9733 ( .B1(n8417), .B2(n8221), .A(n8383), .ZN(n8222) );
  OAI211_X1 U9734 ( .C1(n8421), .C2(n8321), .A(n8223), .B(n8222), .ZN(P2_U3271) );
  AOI21_X1 U9735 ( .B1(n8231), .B2(n8225), .A(n8224), .ZN(n8426) );
  AOI21_X1 U9736 ( .B1(n8422), .B2(n8244), .A(n8226), .ZN(n8423) );
  AOI22_X1 U9737 ( .A1(n8362), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8227), .B2(
        n8369), .ZN(n8228) );
  OAI21_X1 U9738 ( .B1(n8229), .B2(n8311), .A(n8228), .ZN(n8237) );
  OAI211_X1 U9739 ( .C1(n8232), .C2(n8231), .A(n8230), .B(n8351), .ZN(n8235)
         );
  AOI22_X1 U9740 ( .A1(n8233), .A2(n8328), .B1(n8266), .B2(n7599), .ZN(n8234)
         );
  NOR2_X1 U9741 ( .A1(n8425), .A2(n8362), .ZN(n8236) );
  AOI211_X1 U9742 ( .C1(n8423), .C2(n8370), .A(n8237), .B(n8236), .ZN(n8238)
         );
  OAI21_X1 U9743 ( .B1(n8426), .B2(n8321), .A(n8238), .ZN(P2_U3272) );
  AOI21_X1 U9744 ( .B1(n8250), .B2(n8240), .A(n8239), .ZN(n8241) );
  OAI222_X1 U9745 ( .A1(n8372), .A2(n8278), .B1(n8371), .B2(n8242), .C1(n8377), 
        .C2(n8241), .ZN(n8243) );
  INV_X1 U9746 ( .A(n8243), .ZN(n8433) );
  INV_X1 U9747 ( .A(n8244), .ZN(n8245) );
  AOI21_X1 U9748 ( .B1(n8427), .B2(n8256), .A(n8245), .ZN(n8428) );
  AOI22_X1 U9749 ( .A1(n8362), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8246), .B2(
        n8369), .ZN(n8247) );
  OAI21_X1 U9750 ( .B1(n8248), .B2(n8311), .A(n8247), .ZN(n8249) );
  AOI21_X1 U9751 ( .B1(n8428), .B2(n8370), .A(n8249), .ZN(n8254) );
  OR2_X1 U9752 ( .A1(n8251), .A2(n8250), .ZN(n8430) );
  NAND3_X1 U9753 ( .A1(n8430), .A2(n8429), .A3(n8252), .ZN(n8253) );
  OAI211_X1 U9754 ( .C1(n8433), .C2(n8362), .A(n8254), .B(n8253), .ZN(P2_U3273) );
  XNOR2_X1 U9755 ( .A(n8255), .B(n8264), .ZN(n8438) );
  INV_X1 U9756 ( .A(n8279), .ZN(n8258) );
  INV_X1 U9757 ( .A(n8256), .ZN(n8257) );
  AOI21_X1 U9758 ( .B1(n8434), .B2(n8258), .A(n8257), .ZN(n8435) );
  INV_X1 U9759 ( .A(n8259), .ZN(n8260) );
  AOI22_X1 U9760 ( .A1(n8362), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8260), .B2(
        n8369), .ZN(n8261) );
  OAI21_X1 U9761 ( .B1(n8262), .B2(n8311), .A(n8261), .ZN(n8270) );
  OAI211_X1 U9762 ( .C1(n4351), .C2(n8264), .A(n8263), .B(n8351), .ZN(n8268)
         );
  AOI22_X1 U9763 ( .A1(n7599), .A2(n8328), .B1(n8266), .B2(n8265), .ZN(n8267)
         );
  NOR2_X1 U9764 ( .A1(n8437), .A2(n8362), .ZN(n8269) );
  AOI211_X1 U9765 ( .C1(n8435), .C2(n8370), .A(n8270), .B(n8269), .ZN(n8271)
         );
  OAI21_X1 U9766 ( .B1(n8438), .B2(n8321), .A(n8271), .ZN(P2_U3274) );
  XNOR2_X1 U9767 ( .A(n8272), .B(n8275), .ZN(n8444) );
  AOI21_X1 U9768 ( .B1(n8275), .B2(n8274), .A(n8273), .ZN(n8276) );
  OAI222_X1 U9769 ( .A1(n8371), .A2(n8278), .B1(n8372), .B2(n8277), .C1(n8377), 
        .C2(n8276), .ZN(n8439) );
  INV_X1 U9770 ( .A(n8287), .ZN(n8280) );
  AOI21_X1 U9771 ( .B1(n8440), .B2(n8280), .A(n8279), .ZN(n8441) );
  NAND2_X1 U9772 ( .A1(n8441), .A2(n8370), .ZN(n8283) );
  AOI22_X1 U9773 ( .A1(n8362), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8281), .B2(
        n8369), .ZN(n8282) );
  OAI211_X1 U9774 ( .C1(n7595), .C2(n8311), .A(n8283), .B(n8282), .ZN(n8284)
         );
  AOI21_X1 U9775 ( .B1(n8439), .B2(n8383), .A(n8284), .ZN(n8285) );
  OAI21_X1 U9776 ( .B1(n8444), .B2(n8321), .A(n8285), .ZN(P2_U3275) );
  XNOR2_X1 U9777 ( .A(n8286), .B(n8293), .ZN(n8449) );
  AOI21_X1 U9778 ( .B1(n8445), .B2(n8305), .A(n8287), .ZN(n8446) );
  INV_X1 U9779 ( .A(n8288), .ZN(n8289) );
  AOI22_X1 U9780 ( .A1(n8362), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8289), .B2(
        n8369), .ZN(n8290) );
  OAI21_X1 U9781 ( .B1(n8291), .B2(n8311), .A(n8290), .ZN(n8302) );
  INV_X1 U9782 ( .A(n8292), .ZN(n8295) );
  INV_X1 U9783 ( .A(n8293), .ZN(n8294) );
  AOI21_X1 U9784 ( .B1(n8295), .B2(n8294), .A(n8377), .ZN(n8300) );
  OAI22_X1 U9785 ( .A1(n8297), .A2(n8371), .B1(n8372), .B2(n8296), .ZN(n8298)
         );
  AOI21_X1 U9786 ( .B1(n8300), .B2(n8299), .A(n8298), .ZN(n8448) );
  NOR2_X1 U9787 ( .A1(n8448), .A2(n8362), .ZN(n8301) );
  AOI211_X1 U9788 ( .C1(n8446), .C2(n8370), .A(n8302), .B(n8301), .ZN(n8303)
         );
  OAI21_X1 U9789 ( .B1(n8321), .B2(n8449), .A(n8303), .ZN(P2_U3276) );
  XNOR2_X1 U9790 ( .A(n8304), .B(n8313), .ZN(n8454) );
  INV_X1 U9791 ( .A(n8305), .ZN(n8306) );
  AOI211_X1 U9792 ( .C1(n8451), .C2(n8307), .A(n9801), .B(n8306), .ZN(n8450)
         );
  INV_X1 U9793 ( .A(n8308), .ZN(n8309) );
  AOI22_X1 U9794 ( .A1(n8362), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8309), .B2(
        n8369), .ZN(n8310) );
  OAI21_X1 U9795 ( .B1(n8312), .B2(n8311), .A(n8310), .ZN(n8318) );
  XNOR2_X1 U9796 ( .A(n8314), .B(n8313), .ZN(n8316) );
  AOI21_X1 U9797 ( .B1(n8316), .B2(n8351), .A(n8315), .ZN(n8453) );
  NOR2_X1 U9798 ( .A1(n8453), .A2(n8362), .ZN(n8317) );
  AOI211_X1 U9799 ( .C1(n8450), .C2(n8319), .A(n8318), .B(n8317), .ZN(n8320)
         );
  OAI21_X1 U9800 ( .B1(n8454), .B2(n8321), .A(n8320), .ZN(P2_U3277) );
  XNOR2_X1 U9801 ( .A(n8323), .B(n8322), .ZN(n8464) );
  OAI211_X1 U9802 ( .C1(n8326), .C2(n8325), .A(n8324), .B(n8351), .ZN(n8330)
         );
  NAND2_X1 U9803 ( .A1(n8328), .A2(n8327), .ZN(n8329) );
  OAI211_X1 U9804 ( .C1(n8331), .C2(n8372), .A(n8330), .B(n8329), .ZN(n8460)
         );
  INV_X1 U9805 ( .A(n8460), .ZN(n8336) );
  INV_X1 U9806 ( .A(n4359), .ZN(n8333) );
  AOI211_X1 U9807 ( .C1(n8462), .C2(n8333), .A(n9801), .B(n8332), .ZN(n8461)
         );
  AOI22_X1 U9808 ( .A1(n8461), .A2(n8395), .B1(n8369), .B2(n8334), .ZN(n8335)
         );
  OAI211_X1 U9809 ( .C1(n8464), .C2(n8396), .A(n8336), .B(n8335), .ZN(n8337)
         );
  NAND2_X1 U9810 ( .A1(n8337), .A2(n8383), .ZN(n8339) );
  AOI22_X1 U9811 ( .A1(n8462), .A2(n8363), .B1(n8362), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n8338) );
  OAI211_X1 U9812 ( .C1(n8464), .C2(n8340), .A(n8339), .B(n8338), .ZN(P2_U3279) );
  XNOR2_X1 U9813 ( .A(n8342), .B(n8341), .ZN(n8350) );
  OAI22_X1 U9814 ( .A1(n8344), .A2(n8372), .B1(n8371), .B2(n8343), .ZN(n8349)
         );
  OR2_X1 U9815 ( .A1(n8345), .A2(n4409), .ZN(n8346) );
  NAND2_X1 U9816 ( .A1(n8347), .A2(n8346), .ZN(n8470) );
  NOR2_X1 U9817 ( .A1(n8470), .A2(n8396), .ZN(n8348) );
  AOI211_X1 U9818 ( .C1(n8351), .C2(n8350), .A(n8349), .B(n8348), .ZN(n8469)
         );
  INV_X1 U9819 ( .A(n8470), .ZN(n8360) );
  AND2_X1 U9820 ( .A1(n8352), .A2(n8355), .ZN(n8353) );
  OR2_X1 U9821 ( .A1(n8353), .A2(n4359), .ZN(n8466) );
  AOI22_X1 U9822 ( .A1(n8362), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8354), .B2(
        n8369), .ZN(n8357) );
  NAND2_X1 U9823 ( .A1(n8355), .A2(n8363), .ZN(n8356) );
  OAI211_X1 U9824 ( .C1(n8466), .C2(n8358), .A(n8357), .B(n8356), .ZN(n8359)
         );
  AOI21_X1 U9825 ( .B1(n8360), .B2(n8364), .A(n8359), .ZN(n8361) );
  OAI21_X1 U9826 ( .B1(n8469), .B2(n8362), .A(n8361), .ZN(P2_U3280) );
  XNOR2_X1 U9827 ( .A(n8375), .B(n7403), .ZN(n9739) );
  AOI22_X1 U9828 ( .A1(n8364), .A2(n9739), .B1(n8363), .B2(n8367), .ZN(n8386)
         );
  AOI21_X1 U9829 ( .B1(n8367), .B2(n8366), .A(n8365), .ZN(n9733) );
  AOI22_X1 U9830 ( .A1(n8370), .A2(n9733), .B1(n8369), .B2(n8368), .ZN(n8385)
         );
  INV_X1 U9831 ( .A(n8396), .ZN(n8382) );
  OAI22_X1 U9832 ( .A1(n8373), .A2(n8372), .B1(n8371), .B2(n7191), .ZN(n8381)
         );
  NAND3_X1 U9833 ( .A1(n8376), .A2(n8375), .A3(n8374), .ZN(n8378) );
  AOI21_X1 U9834 ( .B1(n8379), .B2(n8378), .A(n8377), .ZN(n8380) );
  AOI211_X1 U9835 ( .C1(n8382), .C2(n9739), .A(n8381), .B(n8380), .ZN(n9736)
         );
  MUX2_X1 U9836 ( .A(n5780), .B(n9736), .S(n8383), .Z(n8384) );
  NAND3_X1 U9837 ( .A1(n8386), .A2(n8385), .A3(n8384), .ZN(P2_U3293) );
  NAND2_X1 U9838 ( .A1(n7805), .A2(n9790), .ZN(n8387) );
  NAND2_X1 U9839 ( .A1(n8390), .A2(n8389), .ZN(n8392) );
  MUX2_X1 U9840 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8476), .S(n9830), .Z(
        P2_U3551) );
  OR3_X1 U9841 ( .A1(n6212), .A2(n8395), .A3(n8394), .ZN(n9456) );
  AOI22_X1 U9842 ( .A1(n8398), .A2(n9791), .B1(n9790), .B2(n8397), .ZN(n8399)
         );
  MUX2_X1 U9843 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8477), .S(n9830), .Z(
        P2_U3549) );
  AOI22_X1 U9844 ( .A1(n8403), .A2(n9791), .B1(n9790), .B2(n8402), .ZN(n8404)
         );
  OAI211_X1 U9845 ( .C1(n8406), .C2(n9795), .A(n8405), .B(n8404), .ZN(n8478)
         );
  MUX2_X1 U9846 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8478), .S(n9830), .Z(
        P2_U3548) );
  AOI22_X1 U9847 ( .A1(n8408), .A2(n9791), .B1(n9790), .B2(n8407), .ZN(n8409)
         );
  OAI211_X1 U9848 ( .C1(n8411), .C2(n9795), .A(n8410), .B(n8409), .ZN(n8479)
         );
  MUX2_X1 U9849 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8479), .S(n9830), .Z(
        P2_U3547) );
  AOI211_X1 U9850 ( .C1(n9790), .C2(n8414), .A(n8413), .B(n8412), .ZN(n8415)
         );
  OAI21_X1 U9851 ( .B1(n8416), .B2(n9795), .A(n8415), .ZN(n8480) );
  MUX2_X1 U9852 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8480), .S(n9830), .Z(
        P2_U3546) );
  AOI211_X1 U9853 ( .C1(n9790), .C2(n8419), .A(n8418), .B(n8417), .ZN(n8420)
         );
  OAI21_X1 U9854 ( .B1(n8421), .B2(n9795), .A(n8420), .ZN(n8481) );
  MUX2_X1 U9855 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8481), .S(n9830), .Z(
        P2_U3545) );
  AOI22_X1 U9856 ( .A1(n8423), .A2(n9791), .B1(n9790), .B2(n8422), .ZN(n8424)
         );
  OAI211_X1 U9857 ( .C1(n8426), .C2(n9795), .A(n8425), .B(n8424), .ZN(n8482)
         );
  MUX2_X1 U9858 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8482), .S(n9830), .Z(
        P2_U3544) );
  AOI22_X1 U9859 ( .A1(n8428), .A2(n9791), .B1(n9790), .B2(n8427), .ZN(n8432)
         );
  NAND3_X1 U9860 ( .A1(n8430), .A2(n8429), .A3(n9806), .ZN(n8431) );
  NAND3_X1 U9861 ( .A1(n8433), .A2(n8432), .A3(n8431), .ZN(n8483) );
  MUX2_X1 U9862 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8483), .S(n9830), .Z(
        P2_U3543) );
  AOI22_X1 U9863 ( .A1(n8435), .A2(n9791), .B1(n9790), .B2(n8434), .ZN(n8436)
         );
  OAI211_X1 U9864 ( .C1(n8438), .C2(n9795), .A(n8437), .B(n8436), .ZN(n8484)
         );
  MUX2_X1 U9865 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8484), .S(n9830), .Z(
        P2_U3542) );
  INV_X1 U9866 ( .A(n8439), .ZN(n8443) );
  AOI22_X1 U9867 ( .A1(n8441), .A2(n9791), .B1(n9790), .B2(n8440), .ZN(n8442)
         );
  OAI211_X1 U9868 ( .C1(n8444), .C2(n9795), .A(n8443), .B(n8442), .ZN(n8485)
         );
  MUX2_X1 U9869 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8485), .S(n9830), .Z(
        P2_U3541) );
  AOI22_X1 U9870 ( .A1(n8446), .A2(n9791), .B1(n9790), .B2(n8445), .ZN(n8447)
         );
  OAI211_X1 U9871 ( .C1(n8449), .C2(n9795), .A(n8448), .B(n8447), .ZN(n8486)
         );
  MUX2_X1 U9872 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8486), .S(n9830), .Z(
        P2_U3540) );
  AOI21_X1 U9873 ( .B1(n9790), .B2(n8451), .A(n8450), .ZN(n8452) );
  OAI211_X1 U9874 ( .C1(n8454), .C2(n9795), .A(n8453), .B(n8452), .ZN(n8487)
         );
  MUX2_X1 U9875 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8487), .S(n9830), .Z(
        P2_U3539) );
  AOI22_X1 U9876 ( .A1(n8456), .A2(n9791), .B1(n9790), .B2(n8455), .ZN(n8457)
         );
  OAI211_X1 U9877 ( .C1(n8459), .C2(n9795), .A(n8458), .B(n8457), .ZN(n8488)
         );
  MUX2_X1 U9878 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8488), .S(n9830), .Z(
        P2_U3538) );
  AOI211_X1 U9879 ( .C1(n9790), .C2(n8462), .A(n8461), .B(n8460), .ZN(n8463)
         );
  OAI21_X1 U9880 ( .B1(n9795), .B2(n8464), .A(n8463), .ZN(n8489) );
  MUX2_X1 U9881 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8489), .S(n9830), .Z(
        P2_U3537) );
  OAI22_X1 U9882 ( .A1(n8466), .A2(n9801), .B1(n8465), .B2(n9799), .ZN(n8467)
         );
  INV_X1 U9883 ( .A(n8467), .ZN(n8468) );
  OAI211_X1 U9884 ( .C1(n9456), .C2(n8470), .A(n8469), .B(n8468), .ZN(n8490)
         );
  MUX2_X1 U9885 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8490), .S(n9830), .Z(
        P2_U3536) );
  INV_X1 U9886 ( .A(n8471), .ZN(n8472) );
  MUX2_X1 U9887 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8476), .S(n9809), .Z(
        P2_U3519) );
  MUX2_X1 U9888 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8477), .S(n9809), .Z(
        P2_U3517) );
  MUX2_X1 U9889 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8478), .S(n9809), .Z(
        P2_U3516) );
  MUX2_X1 U9890 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8479), .S(n9809), .Z(
        P2_U3515) );
  MUX2_X1 U9891 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8480), .S(n9809), .Z(
        P2_U3514) );
  MUX2_X1 U9892 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8481), .S(n9809), .Z(
        P2_U3513) );
  MUX2_X1 U9893 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8482), .S(n9809), .Z(
        P2_U3512) );
  MUX2_X1 U9894 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8483), .S(n9809), .Z(
        P2_U3511) );
  MUX2_X1 U9895 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8484), .S(n9809), .Z(
        P2_U3510) );
  MUX2_X1 U9896 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8485), .S(n9809), .Z(
        P2_U3509) );
  MUX2_X1 U9897 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8486), .S(n9809), .Z(
        P2_U3508) );
  MUX2_X1 U9898 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8487), .S(n9809), .Z(
        P2_U3507) );
  MUX2_X1 U9899 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8488), .S(n9809), .Z(
        P2_U3505) );
  MUX2_X1 U9900 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8489), .S(n9809), .Z(
        P2_U3502) );
  MUX2_X1 U9901 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8490), .S(n9809), .Z(
        P2_U3499) );
  AOI22_X1 U9902 ( .A1(n8492), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8491), .ZN(n8493) );
  OAI21_X1 U9903 ( .B1(n8494), .B2(n7626), .A(n8493), .ZN(P2_U3328) );
  MUX2_X1 U9904 ( .A(n8495), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U9905 ( .A(n9262), .ZN(n9044) );
  AOI21_X1 U9906 ( .B1(n8594), .B2(n8497), .A(n8496), .ZN(n8498) );
  OAI21_X1 U9907 ( .B1(n8499), .B2(n8498), .A(n8595), .ZN(n8504) );
  INV_X1 U9908 ( .A(n9080), .ZN(n9048) );
  OAI22_X1 U9909 ( .A1(n9048), .A2(n8599), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8500), .ZN(n8502) );
  NOR2_X1 U9910 ( .A1(n9049), .A2(n8615), .ZN(n8501) );
  AOI211_X1 U9911 ( .C1(n9042), .C2(n8612), .A(n8502), .B(n8501), .ZN(n8503)
         );
  OAI211_X1 U9912 ( .C1(n9044), .C2(n8604), .A(n8504), .B(n8503), .ZN(P1_U3212) );
  INV_X1 U9913 ( .A(n8505), .ZN(n8507) );
  NOR2_X1 U9914 ( .A1(n8507), .A2(n8506), .ZN(n8509) );
  XNOR2_X1 U9915 ( .A(n8509), .B(n8508), .ZN(n8514) );
  NAND2_X1 U9916 ( .A1(n9113), .A2(n8578), .ZN(n8511) );
  AOI22_X1 U9917 ( .A1(n9106), .A2(n8611), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8510) );
  OAI211_X1 U9918 ( .C1(n8588), .C2(n9102), .A(n8511), .B(n8510), .ZN(n8512)
         );
  AOI21_X1 U9919 ( .B1(n9282), .B2(n8617), .A(n8512), .ZN(n8513) );
  OAI21_X1 U9920 ( .B1(n8514), .B2(n8619), .A(n8513), .ZN(P1_U3214) );
  XOR2_X1 U9921 ( .A(n8516), .B(n8515), .Z(n8521) );
  AOI22_X1 U9922 ( .A1(n8578), .A2(n9167), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3084), .ZN(n8518) );
  NAND2_X1 U9923 ( .A1(n8611), .A2(n9198), .ZN(n8517) );
  OAI211_X1 U9924 ( .C1(n8588), .C2(n9160), .A(n8518), .B(n8517), .ZN(n8519)
         );
  AOI21_X1 U9925 ( .B1(n9302), .B2(n8617), .A(n8519), .ZN(n8520) );
  OAI21_X1 U9926 ( .B1(n8521), .B2(n8619), .A(n8520), .ZN(P1_U3217) );
  XOR2_X1 U9927 ( .A(n8523), .B(n8522), .Z(n8529) );
  INV_X1 U9928 ( .A(n8524), .ZN(n9138) );
  NAND2_X1 U9929 ( .A1(n9106), .A2(n8578), .ZN(n8526) );
  AOI22_X1 U9930 ( .A1(n8611), .A2(n9167), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8525) );
  OAI211_X1 U9931 ( .C1(n8588), .C2(n9138), .A(n8526), .B(n8525), .ZN(n8527)
         );
  AOI21_X1 U9932 ( .B1(n9294), .B2(n8617), .A(n8527), .ZN(n8528) );
  OAI21_X1 U9933 ( .B1(n8529), .B2(n8619), .A(n8528), .ZN(P1_U3221) );
  OAI21_X1 U9934 ( .B1(n8531), .B2(n8530), .A(n8593), .ZN(n8532) );
  NAND2_X1 U9935 ( .A1(n8532), .A2(n8595), .ZN(n8536) );
  AOI22_X1 U9936 ( .A1(n9113), .A2(n8611), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8533) );
  OAI21_X1 U9937 ( .B1(n8588), .B2(n9073), .A(n8533), .ZN(n8534) );
  AOI21_X1 U9938 ( .B1(n8578), .B2(n9080), .A(n8534), .ZN(n8535) );
  OAI211_X1 U9939 ( .C1(n9076), .C2(n8604), .A(n8536), .B(n8535), .ZN(P1_U3223) );
  AOI21_X1 U9940 ( .B1(n8539), .B2(n8538), .A(n8537), .ZN(n8544) );
  AOI22_X1 U9941 ( .A1(n8578), .A2(n9182), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n8541) );
  NAND2_X1 U9942 ( .A1(n8612), .A2(n9214), .ZN(n8540) );
  OAI211_X1 U9943 ( .C1(n9210), .C2(n8599), .A(n8541), .B(n8540), .ZN(n8542)
         );
  AOI21_X1 U9944 ( .B1(n9319), .B2(n8617), .A(n8542), .ZN(n8543) );
  OAI21_X1 U9945 ( .B1(n8544), .B2(n8619), .A(n8543), .ZN(P1_U3224) );
  AOI21_X1 U9946 ( .B1(n8548), .B2(n8547), .A(n8546), .ZN(n8554) );
  OAI22_X1 U9947 ( .A1(n8615), .A2(n8647), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8549), .ZN(n8550) );
  AOI21_X1 U9948 ( .B1(n8611), .B2(n9233), .A(n8550), .ZN(n8551) );
  OAI21_X1 U9949 ( .B1(n8588), .B2(n9192), .A(n8551), .ZN(n8552) );
  AOI21_X1 U9950 ( .B1(n9312), .B2(n8617), .A(n8552), .ZN(n8553) );
  OAI21_X1 U9951 ( .B1(n8554), .B2(n8619), .A(n8553), .ZN(P1_U3226) );
  INV_X1 U9952 ( .A(n9278), .ZN(n9090) );
  OAI21_X1 U9953 ( .B1(n8557), .B2(n8556), .A(n8555), .ZN(n8558) );
  NAND2_X1 U9954 ( .A1(n8558), .A2(n8595), .ZN(n8562) );
  AOI22_X1 U9955 ( .A1(n9126), .A2(n8611), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8559) );
  OAI21_X1 U9956 ( .B1(n8971), .B2(n8615), .A(n8559), .ZN(n8560) );
  AOI21_X1 U9957 ( .B1(n9088), .B2(n8612), .A(n8560), .ZN(n8561) );
  OAI211_X1 U9958 ( .C1(n9090), .C2(n8604), .A(n8562), .B(n8561), .ZN(P1_U3227) );
  INV_X1 U9959 ( .A(n8564), .ZN(n8566) );
  NAND2_X1 U9960 ( .A1(n8566), .A2(n8565), .ZN(n8567) );
  XNOR2_X1 U9961 ( .A(n8563), .B(n8567), .ZN(n8573) );
  OAI22_X1 U9962 ( .A1(n8963), .A2(n8615), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8568), .ZN(n8569) );
  AOI21_X1 U9963 ( .B1(n8611), .B2(n9183), .A(n8569), .ZN(n8570) );
  OAI21_X1 U9964 ( .B1(n8588), .B2(n9145), .A(n8570), .ZN(n8571) );
  AOI21_X1 U9965 ( .B1(n9297), .B2(n8617), .A(n8571), .ZN(n8572) );
  OAI21_X1 U9966 ( .B1(n8573), .B2(n8619), .A(n8572), .ZN(P1_U3231) );
  NAND2_X1 U9967 ( .A1(n8575), .A2(n8574), .ZN(n8576) );
  XOR2_X1 U9968 ( .A(n8577), .B(n8576), .Z(n8583) );
  NAND2_X1 U9969 ( .A1(n9126), .A2(n8578), .ZN(n8580) );
  INV_X1 U9970 ( .A(n8963), .ZN(n9152) );
  AOI22_X1 U9971 ( .A1(n9152), .A2(n8611), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8579) );
  OAI211_X1 U9972 ( .C1(n8588), .C2(n9120), .A(n8580), .B(n8579), .ZN(n8581)
         );
  AOI21_X1 U9973 ( .B1(n9287), .B2(n8617), .A(n8581), .ZN(n8582) );
  OAI21_X1 U9974 ( .B1(n8583), .B2(n8619), .A(n8582), .ZN(P1_U3233) );
  XNOR2_X1 U9975 ( .A(n4334), .B(n8584), .ZN(n8585) );
  XNOR2_X1 U9976 ( .A(n4315), .B(n8585), .ZN(n8591) );
  NAND2_X1 U9977 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9622) );
  OAI21_X1 U9978 ( .B1(n8615), .B2(n8961), .A(n9622), .ZN(n8586) );
  AOI21_X1 U9979 ( .B1(n8611), .B2(n9182), .A(n8586), .ZN(n8587) );
  OAI21_X1 U9980 ( .B1(n8588), .B2(n9176), .A(n8587), .ZN(n8589) );
  AOI21_X1 U9981 ( .B1(n9308), .B2(n8617), .A(n8589), .ZN(n8590) );
  OAI21_X1 U9982 ( .B1(n8591), .B2(n8619), .A(n8590), .ZN(P1_U3236) );
  INV_X1 U9983 ( .A(n9267), .ZN(n9061) );
  AND2_X1 U9984 ( .A1(n8593), .A2(n8592), .ZN(n8597) );
  OAI211_X1 U9985 ( .C1(n8597), .C2(n8596), .A(n8595), .B(n8594), .ZN(n8603)
         );
  OAI22_X1 U9986 ( .A1(n8971), .A2(n8599), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8598), .ZN(n8601) );
  NOR2_X1 U9987 ( .A1(n9024), .A2(n8615), .ZN(n8600) );
  AOI211_X1 U9988 ( .C1(n9059), .C2(n8612), .A(n8601), .B(n8600), .ZN(n8602)
         );
  OAI211_X1 U9989 ( .C1(n9061), .C2(n8604), .A(n8603), .B(n8602), .ZN(P1_U3238) );
  INV_X1 U9990 ( .A(n8605), .ZN(n8607) );
  NAND2_X1 U9991 ( .A1(n8607), .A2(n8606), .ZN(n8609) );
  XNOR2_X1 U9992 ( .A(n8609), .B(n8608), .ZN(n8620) );
  INV_X1 U9993 ( .A(n9233), .ZN(n8787) );
  AOI21_X1 U9994 ( .B1(n8611), .B2(n4509), .A(n8610), .ZN(n8614) );
  NAND2_X1 U9995 ( .A1(n8612), .A2(n9226), .ZN(n8613) );
  OAI211_X1 U9996 ( .C1(n8787), .C2(n8615), .A(n8614), .B(n8613), .ZN(n8616)
         );
  AOI21_X1 U9997 ( .B1(n9322), .B2(n8617), .A(n8616), .ZN(n8618) );
  OAI21_X1 U9998 ( .B1(n8620), .B2(n8619), .A(n8618), .ZN(P1_U3239) );
  NAND2_X1 U9999 ( .A1(n8621), .A2(n5229), .ZN(n8624) );
  OR2_X1 U10000 ( .A1(n8635), .A2(n8622), .ZN(n8623) );
  INV_X1 U10001 ( .A(n9248), .ZN(n8949) );
  INV_X1 U10002 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9937) );
  NAND2_X1 U10003 ( .A1(n8625), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U10004 ( .A1(n8626), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8627) );
  OAI211_X1 U10005 ( .C1(n8629), .C2(n9937), .A(n8628), .B(n8627), .ZN(n9007)
         );
  INV_X1 U10006 ( .A(n9007), .ZN(n8630) );
  NOR2_X1 U10007 ( .A1(n8949), .A2(n8630), .ZN(n8772) );
  INV_X1 U10008 ( .A(n8772), .ZN(n8631) );
  NAND2_X1 U10009 ( .A1(n8631), .A2(n8944), .ZN(n8633) );
  NOR2_X1 U10010 ( .A1(n8635), .A2(n6413), .ZN(n8632) );
  INV_X1 U10011 ( .A(n8945), .ZN(n9240) );
  NAND2_X1 U10012 ( .A1(n8633), .A2(n9240), .ZN(n8832) );
  NAND2_X1 U10013 ( .A1(n8634), .A2(n5229), .ZN(n8637) );
  OR2_X1 U10014 ( .A1(n8635), .A2(n9361), .ZN(n8636) );
  NAND2_X1 U10015 ( .A1(n9252), .A2(n9023), .ZN(n8861) );
  NAND2_X1 U10016 ( .A1(n9256), .A2(n9049), .ZN(n9003) );
  MUX2_X1 U10017 ( .A(n9003), .B(n9002), .S(n8741), .Z(n8638) );
  NAND2_X1 U10018 ( .A1(n8979), .A2(n8638), .ZN(n8739) );
  OAI21_X1 U10019 ( .B1(n8739), .B2(n9001), .A(n8827), .ZN(n8640) );
  NAND2_X1 U10020 ( .A1(n8944), .A2(n9007), .ZN(n8639) );
  NAND2_X1 U10021 ( .A1(n8949), .A2(n8639), .ZN(n8828) );
  NAND2_X1 U10022 ( .A1(n8640), .A2(n8828), .ZN(n8641) );
  AND2_X1 U10023 ( .A1(n8832), .A2(n8641), .ZN(n8742) );
  INV_X1 U10024 ( .A(n8944), .ZN(n8642) );
  AND2_X1 U10025 ( .A1(n9240), .A2(n8642), .ZN(n8773) );
  INV_X1 U10026 ( .A(n8773), .ZN(n8643) );
  INV_X1 U10027 ( .A(n8741), .ZN(n8738) );
  NAND2_X1 U10028 ( .A1(n9262), .A2(n9024), .ZN(n8779) );
  XNOR2_X1 U10029 ( .A(n9278), .B(n9113), .ZN(n9092) );
  INV_X1 U10030 ( .A(n9092), .ZN(n8728) );
  AND2_X1 U10031 ( .A1(n9282), .A2(n9126), .ZN(n8967) );
  OR2_X1 U10032 ( .A1(n8728), .A2(n8967), .ZN(n8644) );
  NAND2_X1 U10033 ( .A1(n9272), .A2(n8971), .ZN(n8745) );
  INV_X1 U10034 ( .A(n9113), .ZN(n8969) );
  NAND2_X1 U10035 ( .A1(n9278), .A2(n8969), .ZN(n9077) );
  OAI21_X1 U10036 ( .B1(n9105), .B2(n8644), .A(n8998), .ZN(n8646) );
  OR2_X1 U10037 ( .A1(n9278), .A2(n8969), .ZN(n8806) );
  OAI211_X1 U10038 ( .C1(n8644), .C2(n8966), .A(n8806), .B(n9062), .ZN(n8645)
         );
  MUX2_X1 U10039 ( .A(n8646), .B(n8645), .S(n8741), .Z(n8730) );
  NAND2_X1 U10040 ( .A1(n8997), .A2(n8994), .ZN(n8803) );
  INV_X1 U10041 ( .A(n8803), .ZN(n8719) );
  OR2_X1 U10042 ( .A1(n9308), .A2(n8647), .ZN(n8748) );
  OR2_X1 U10043 ( .A1(n9312), .A2(n9211), .ZN(n8988) );
  AND2_X1 U10044 ( .A1(n8748), .A2(n8988), .ZN(n8798) );
  INV_X1 U10045 ( .A(n8798), .ZN(n8649) );
  NAND2_X1 U10046 ( .A1(n9308), .A2(n8647), .ZN(n8989) );
  AND2_X1 U10047 ( .A1(n9312), .A2(n9211), .ZN(n8987) );
  INV_X1 U10048 ( .A(n8987), .ZN(n8648) );
  AND2_X1 U10049 ( .A1(n8989), .A2(n8648), .ZN(n8794) );
  INV_X1 U10050 ( .A(n8794), .ZN(n8823) );
  MUX2_X1 U10051 ( .A(n8649), .B(n8823), .S(n8738), .Z(n8650) );
  INV_X1 U10052 ( .A(n8650), .ZN(n8708) );
  MUX2_X1 U10053 ( .A(n9233), .B(n9319), .S(n8738), .Z(n8706) );
  XNOR2_X1 U10054 ( .A(n9319), .B(n9233), .ZN(n9206) );
  INV_X1 U10055 ( .A(n8988), .ZN(n8651) );
  INV_X1 U10056 ( .A(n9189), .ZN(n9196) );
  NAND2_X1 U10057 ( .A1(n8751), .A2(n8741), .ZN(n8652) );
  NAND2_X1 U10058 ( .A1(n8653), .A2(n8652), .ZN(n8655) );
  AND2_X1 U10059 ( .A1(n8660), .A2(n8656), .ZN(n8844) );
  NAND2_X1 U10060 ( .A1(n8664), .A2(n8844), .ZN(n8658) );
  AND2_X1 U10061 ( .A1(n8812), .A2(n8665), .ZN(n8843) );
  INV_X1 U10062 ( .A(n8819), .ZN(n8657) );
  AOI21_X1 U10063 ( .B1(n8658), .B2(n8843), .A(n8657), .ZN(n8668) );
  INV_X1 U10064 ( .A(n8660), .ZN(n8663) );
  NAND2_X1 U10065 ( .A1(n8660), .A2(n8659), .ZN(n8662) );
  AND2_X1 U10066 ( .A1(n8662), .A2(n8661), .ZN(n8814) );
  OAI21_X1 U10067 ( .B1(n8664), .B2(n8663), .A(n8814), .ZN(n8666) );
  INV_X1 U10068 ( .A(n8665), .ZN(n8815) );
  AOI21_X1 U10069 ( .B1(n8666), .B2(n8819), .A(n8815), .ZN(n8667) );
  OR2_X1 U10070 ( .A1(n8683), .A2(n4832), .ZN(n8782) );
  OAI21_X1 U10071 ( .B1(n8682), .B2(n8670), .A(n4831), .ZN(n8673) );
  INV_X1 U10072 ( .A(n8671), .ZN(n8672) );
  NAND2_X1 U10073 ( .A1(n8673), .A2(n8672), .ZN(n8674) );
  NAND4_X1 U10074 ( .A1(n8674), .A2(n8685), .A3(n8678), .A4(n8761), .ZN(n8681)
         );
  AND2_X1 U10075 ( .A1(n8698), .A2(n8675), .ZN(n8786) );
  INV_X1 U10076 ( .A(n8676), .ZN(n8677) );
  AND2_X1 U10077 ( .A1(n8691), .A2(n8677), .ZN(n8785) );
  INV_X1 U10078 ( .A(n8785), .ZN(n8679) );
  NAND2_X1 U10079 ( .A1(n8679), .A2(n8678), .ZN(n8680) );
  NAND3_X1 U10080 ( .A1(n8681), .A2(n8786), .A3(n8680), .ZN(n8697) );
  OAI211_X1 U10081 ( .C1(n8682), .C2(n4832), .A(n9389), .B(n8820), .ZN(n8686)
         );
  INV_X1 U10082 ( .A(n8683), .ZN(n8684) );
  NAND3_X1 U10083 ( .A1(n8686), .A2(n8685), .A3(n8684), .ZN(n8688) );
  NAND4_X1 U10084 ( .A1(n8688), .A2(n8687), .A3(n8691), .A4(n8761), .ZN(n8696)
         );
  NAND2_X1 U10085 ( .A1(n8689), .A2(n8878), .ZN(n8690) );
  NAND2_X1 U10086 ( .A1(n8981), .A2(n8690), .ZN(n8699) );
  INV_X1 U10087 ( .A(n8691), .ZN(n8692) );
  NOR2_X1 U10088 ( .A1(n8693), .A2(n8692), .ZN(n8694) );
  OR2_X1 U10089 ( .A1(n8699), .A2(n8694), .ZN(n8790) );
  INV_X1 U10090 ( .A(n8790), .ZN(n8695) );
  NAND2_X1 U10091 ( .A1(n9322), .A2(n9210), .ZN(n8983) );
  NAND2_X1 U10092 ( .A1(n9204), .A2(n8983), .ZN(n9229) );
  INV_X1 U10093 ( .A(n9229), .ZN(n9222) );
  NAND2_X1 U10094 ( .A1(n8699), .A2(n8698), .ZN(n8701) );
  INV_X1 U10095 ( .A(n8786), .ZN(n8700) );
  NAND2_X1 U10096 ( .A1(n8700), .A2(n8981), .ZN(n8789) );
  MUX2_X1 U10097 ( .A(n8701), .B(n8789), .S(n8741), .Z(n8702) );
  NAND2_X1 U10098 ( .A1(n9319), .A2(n9233), .ZN(n8959) );
  NAND2_X1 U10099 ( .A1(n8706), .A2(n8959), .ZN(n8704) );
  MUX2_X1 U10100 ( .A(n8983), .B(n9204), .S(n8741), .Z(n8703) );
  OAI211_X1 U10101 ( .C1(n8706), .C2(n9206), .A(n9196), .B(n8705), .ZN(n8707)
         );
  NAND2_X1 U10102 ( .A1(n8708), .A2(n8707), .ZN(n8711) );
  OR2_X1 U10103 ( .A1(n9302), .A2(n8961), .ZN(n8747) );
  NAND3_X1 U10104 ( .A1(n8711), .A2(n8748), .A3(n8747), .ZN(n8709) );
  INV_X1 U10105 ( .A(n9167), .ZN(n9136) );
  NAND2_X1 U10106 ( .A1(n9297), .A2(n9136), .ZN(n8746) );
  NAND2_X1 U10107 ( .A1(n9302), .A2(n8961), .ZN(n9149) );
  NAND3_X1 U10108 ( .A1(n8709), .A2(n8746), .A3(n9149), .ZN(n8714) );
  AND2_X1 U10109 ( .A1(n8992), .A2(n8747), .ZN(n8795) );
  NAND2_X1 U10110 ( .A1(n9149), .A2(n8989), .ZN(n8797) );
  INV_X1 U10111 ( .A(n8797), .ZN(n8710) );
  NAND2_X1 U10112 ( .A1(n8711), .A2(n8710), .ZN(n8712) );
  NAND2_X1 U10113 ( .A1(n8795), .A2(n8712), .ZN(n8713) );
  INV_X1 U10114 ( .A(n8721), .ZN(n8717) );
  NAND2_X1 U10115 ( .A1(n8796), .A2(n8992), .ZN(n8716) );
  NAND2_X1 U10116 ( .A1(n9287), .A2(n9135), .ZN(n8995) );
  NAND2_X1 U10117 ( .A1(n9294), .A2(n8963), .ZN(n8993) );
  NAND2_X1 U10118 ( .A1(n8995), .A2(n8993), .ZN(n8724) );
  INV_X1 U10119 ( .A(n8724), .ZN(n8715) );
  OAI21_X1 U10120 ( .B1(n8717), .B2(n8716), .A(n8715), .ZN(n8718) );
  INV_X1 U10121 ( .A(n8796), .ZN(n8720) );
  NOR2_X1 U10122 ( .A1(n8721), .A2(n8720), .ZN(n8725) );
  INV_X1 U10123 ( .A(n8746), .ZN(n8722) );
  AND2_X1 U10124 ( .A1(n8796), .A2(n8722), .ZN(n8723) );
  OR2_X1 U10125 ( .A1(n8724), .A2(n8723), .ZN(n8801) );
  OAI21_X1 U10126 ( .B1(n8725), .B2(n8801), .A(n8994), .ZN(n8726) );
  NAND2_X1 U10127 ( .A1(n9282), .A2(n8966), .ZN(n8802) );
  NAND2_X1 U10128 ( .A1(n8726), .A2(n8802), .ZN(n8727) );
  MUX2_X1 U10129 ( .A(n9062), .B(n8745), .S(n8741), .Z(n8729) );
  NAND2_X1 U10130 ( .A1(n9267), .A2(n9080), .ZN(n8975) );
  OAI21_X1 U10131 ( .B1(n8733), .B2(n8975), .A(n9046), .ZN(n8735) );
  INV_X1 U10132 ( .A(n8974), .ZN(n8732) );
  MUX2_X1 U10133 ( .A(n9080), .B(n9267), .S(n8741), .Z(n8731) );
  OAI211_X1 U10134 ( .C1(n8738), .C2(n8779), .A(n8736), .B(n9027), .ZN(n8737)
         );
  INV_X1 U10135 ( .A(n8737), .ZN(n8740) );
  AND2_X1 U10136 ( .A1(n8945), .A2(n8944), .ZN(n8865) );
  INV_X1 U10137 ( .A(n8865), .ZN(n8743) );
  AND4_X1 U10138 ( .A1(n8777), .A2(n5648), .A3(n8743), .A4(n5654), .ZN(n8744)
         );
  NOR2_X1 U10139 ( .A1(n9248), .A2(n9007), .ZN(n8860) );
  INV_X1 U10140 ( .A(n8979), .ZN(n9005) );
  NAND2_X1 U10141 ( .A1(n8997), .A2(n8802), .ZN(n9110) );
  NAND2_X1 U10142 ( .A1(n8994), .A2(n8995), .ZN(n9125) );
  NAND2_X1 U10143 ( .A1(n8796), .A2(n8993), .ZN(n9133) );
  NAND2_X1 U10144 ( .A1(n8992), .A2(n8746), .ZN(n9151) );
  NAND2_X1 U10145 ( .A1(n8748), .A2(n8989), .ZN(n9172) );
  INV_X1 U10146 ( .A(n9172), .ZN(n9181) );
  INV_X1 U10147 ( .A(n8749), .ZN(n8764) );
  NAND2_X1 U10148 ( .A1(n8751), .A2(n8750), .ZN(n8811) );
  NOR4_X1 U10149 ( .A1(n8753), .A2(n8752), .A3(n6437), .A4(n8811), .ZN(n8757)
         );
  AND2_X1 U10150 ( .A1(n8844), .A2(n8754), .ZN(n8850) );
  INV_X1 U10151 ( .A(n8755), .ZN(n8756) );
  NAND4_X1 U10152 ( .A1(n8757), .A2(n8850), .A3(n8756), .A4(n8812), .ZN(n8760)
         );
  NOR4_X1 U10153 ( .A1(n9396), .A2(n8760), .A3(n8759), .A4(n6843), .ZN(n8762)
         );
  NAND4_X1 U10154 ( .A1(n8764), .A2(n8763), .A3(n8762), .A4(n8761), .ZN(n8765)
         );
  NOR4_X1 U10155 ( .A1(n9189), .A2(n8766), .A3(n9229), .A4(n8765), .ZN(n8767)
         );
  NAND4_X1 U10156 ( .A1(n9166), .A2(n9181), .A3(n8767), .A4(n9206), .ZN(n8768)
         );
  OR4_X1 U10157 ( .A1(n9125), .A2(n9133), .A3(n9151), .A4(n8768), .ZN(n8769)
         );
  NOR4_X1 U10158 ( .A1(n9079), .A2(n8728), .A3(n9110), .A4(n8769), .ZN(n8770)
         );
  NAND2_X1 U10159 ( .A1(n8974), .A2(n8975), .ZN(n9065) );
  NAND4_X1 U10160 ( .A1(n9027), .A2(n9046), .A3(n8770), .A4(n9065), .ZN(n8771)
         );
  NOR4_X1 U10161 ( .A1(n8865), .A2(n8860), .A3(n9005), .A4(n8771), .ZN(n8774)
         );
  NOR2_X1 U10162 ( .A1(n8773), .A2(n8772), .ZN(n8867) );
  AOI21_X1 U10163 ( .B1(n8774), .B2(n8867), .A(n5648), .ZN(n8834) );
  INV_X1 U10164 ( .A(n8834), .ZN(n8775) );
  OAI21_X1 U10165 ( .B1(n8777), .B2(n8776), .A(n8775), .ZN(n8836) );
  AND2_X1 U10166 ( .A1(n9267), .A2(n9048), .ZN(n8999) );
  NAND2_X1 U10167 ( .A1(n9001), .A2(n8999), .ZN(n8778) );
  AND3_X1 U10168 ( .A1(n9003), .A2(n8779), .A3(n8778), .ZN(n8857) );
  OR2_X1 U10169 ( .A1(n9267), .A2(n9048), .ZN(n8780) );
  AND2_X1 U10170 ( .A1(n8780), .A2(n9062), .ZN(n9000) );
  NAND2_X1 U10171 ( .A1(n8802), .A2(n9149), .ZN(n8781) );
  NOR2_X1 U10172 ( .A1(n8781), .A2(n8801), .ZN(n8810) );
  NAND2_X1 U10173 ( .A1(n9319), .A2(n8787), .ZN(n8985) );
  NOR2_X1 U10174 ( .A1(n8783), .A2(n8782), .ZN(n8792) );
  NAND4_X1 U10175 ( .A1(n8983), .A2(n8786), .A3(n8785), .A4(n8784), .ZN(n8818)
         );
  OR2_X1 U10176 ( .A1(n9319), .A2(n8787), .ZN(n8788) );
  AND2_X1 U10177 ( .A1(n8788), .A2(n9204), .ZN(n8984) );
  NAND3_X1 U10178 ( .A1(n8790), .A2(n8983), .A3(n8789), .ZN(n8791) );
  OAI211_X1 U10179 ( .C1(n8792), .C2(n8818), .A(n8984), .B(n8791), .ZN(n8793)
         );
  NAND4_X1 U10180 ( .A1(n8810), .A2(n8794), .A3(n8985), .A4(n8793), .ZN(n8807)
         );
  OAI211_X1 U10181 ( .C1(n8798), .C2(n8797), .A(n8796), .B(n8795), .ZN(n8799)
         );
  INV_X1 U10182 ( .A(n8799), .ZN(n8800) );
  NOR2_X1 U10183 ( .A1(n8801), .A2(n8800), .ZN(n8804) );
  OAI21_X1 U10184 ( .B1(n8804), .B2(n8803), .A(n8802), .ZN(n8805) );
  NAND3_X1 U10185 ( .A1(n8807), .A2(n8806), .A3(n8805), .ZN(n8808) );
  NAND2_X1 U10186 ( .A1(n8998), .A2(n8808), .ZN(n8809) );
  AND2_X1 U10187 ( .A1(n9000), .A2(n8809), .ZN(n8854) );
  NAND2_X1 U10188 ( .A1(n8998), .A2(n8810), .ZN(n8853) );
  INV_X1 U10189 ( .A(n8811), .ZN(n8845) );
  NAND3_X1 U10190 ( .A1(n6485), .A2(n8845), .A3(n8812), .ZN(n8817) );
  INV_X1 U10191 ( .A(n8850), .ZN(n8813) );
  NAND2_X1 U10192 ( .A1(n8814), .A2(n8813), .ZN(n8816) );
  AOI21_X1 U10193 ( .B1(n8817), .B2(n8816), .A(n8815), .ZN(n8824) );
  INV_X1 U10194 ( .A(n8818), .ZN(n8821) );
  NAND4_X1 U10195 ( .A1(n8985), .A2(n8821), .A3(n8820), .A4(n8819), .ZN(n8822)
         );
  OR2_X1 U10196 ( .A1(n8823), .A2(n8822), .ZN(n8851) );
  OR3_X1 U10197 ( .A1(n8853), .A2(n8824), .A3(n8851), .ZN(n8825) );
  NAND3_X1 U10198 ( .A1(n8854), .A2(n9001), .A3(n8825), .ZN(n8826) );
  AND2_X1 U10199 ( .A1(n8857), .A2(n8826), .ZN(n8829) );
  NAND2_X1 U10200 ( .A1(n8827), .A2(n9002), .ZN(n8863) );
  OAI211_X1 U10201 ( .C1(n8829), .C2(n8863), .A(n8828), .B(n8861), .ZN(n8831)
         );
  AOI211_X1 U10202 ( .C1(n8832), .C2(n8831), .A(n8830), .B(n8865), .ZN(n8833)
         );
  NOR2_X1 U10203 ( .A1(n8834), .A2(n8833), .ZN(n8835) );
  OAI211_X1 U10204 ( .C1(n6453), .C2(n8838), .A(n5648), .B(n8837), .ZN(n8840)
         );
  NAND2_X1 U10205 ( .A1(n8840), .A2(n8839), .ZN(n8841) );
  OAI22_X1 U10206 ( .A1(n8842), .A2(n8841), .B1(n6456), .B2(n6457), .ZN(n8849)
         );
  INV_X1 U10207 ( .A(n8843), .ZN(n8848) );
  INV_X1 U10208 ( .A(n8844), .ZN(n8846) );
  NOR2_X1 U10209 ( .A1(n8846), .A2(n8845), .ZN(n8847) );
  AOI211_X1 U10210 ( .C1(n8850), .C2(n8849), .A(n8848), .B(n8847), .ZN(n8852)
         );
  NOR3_X1 U10211 ( .A1(n8853), .A2(n8852), .A3(n8851), .ZN(n8856) );
  INV_X1 U10212 ( .A(n8854), .ZN(n8855) );
  NOR2_X1 U10213 ( .A1(n8856), .A2(n8855), .ZN(n8859) );
  INV_X1 U10214 ( .A(n8857), .ZN(n8858) );
  AOI21_X1 U10215 ( .B1(n9046), .B2(n8859), .A(n8858), .ZN(n8864) );
  INV_X1 U10216 ( .A(n8860), .ZN(n8862) );
  OAI211_X1 U10217 ( .C1(n8864), .C2(n8863), .A(n8862), .B(n8861), .ZN(n8866)
         );
  AOI21_X1 U10218 ( .B1(n8867), .B2(n8866), .A(n8865), .ZN(n8868) );
  XNOR2_X1 U10219 ( .A(n8868), .B(n9646), .ZN(n8869) );
  NAND2_X1 U10220 ( .A1(n8869), .A2(n6837), .ZN(n8870) );
  NAND3_X1 U10221 ( .A1(n8873), .A2(n9522), .A3(n9490), .ZN(n8874) );
  OAI211_X1 U10222 ( .C1(n5046), .C2(n8876), .A(n8874), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8875) );
  OAI21_X1 U10223 ( .B1(n8877), .B2(n8876), .A(n8875), .ZN(P1_U3240) );
  MUX2_X1 U10224 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9007), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10225 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9009), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10226 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9066), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10227 ( .A(n9080), .B(P1_DATAO_REG_26__SCAN_IN), .S(n8890), .Z(
        P1_U3581) );
  MUX2_X1 U10228 ( .A(n8972), .B(P1_DATAO_REG_25__SCAN_IN), .S(n8890), .Z(
        P1_U3580) );
  MUX2_X1 U10229 ( .A(n9113), .B(P1_DATAO_REG_24__SCAN_IN), .S(n8890), .Z(
        P1_U3579) );
  MUX2_X1 U10230 ( .A(n9126), .B(P1_DATAO_REG_23__SCAN_IN), .S(n8890), .Z(
        P1_U3578) );
  MUX2_X1 U10231 ( .A(n9106), .B(P1_DATAO_REG_22__SCAN_IN), .S(n8890), .Z(
        P1_U3577) );
  MUX2_X1 U10232 ( .A(n9152), .B(P1_DATAO_REG_21__SCAN_IN), .S(n8890), .Z(
        P1_U3576) );
  MUX2_X1 U10233 ( .A(n9167), .B(P1_DATAO_REG_20__SCAN_IN), .S(n8890), .Z(
        P1_U3575) );
  MUX2_X1 U10234 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9183), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10235 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9198), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10236 ( .A(n9182), .B(P1_DATAO_REG_17__SCAN_IN), .S(n8890), .Z(
        P1_U3572) );
  MUX2_X1 U10237 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9233), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10238 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n8958), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10239 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n4509), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10240 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8878), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10241 ( .A(n8879), .B(P1_DATAO_REG_12__SCAN_IN), .S(n8890), .Z(
        P1_U3567) );
  MUX2_X1 U10242 ( .A(n8880), .B(P1_DATAO_REG_11__SCAN_IN), .S(n8890), .Z(
        P1_U3566) );
  MUX2_X1 U10243 ( .A(n8881), .B(P1_DATAO_REG_10__SCAN_IN), .S(n8890), .Z(
        P1_U3565) );
  MUX2_X1 U10244 ( .A(n8882), .B(P1_DATAO_REG_9__SCAN_IN), .S(n8890), .Z(
        P1_U3564) );
  MUX2_X1 U10245 ( .A(n8883), .B(P1_DATAO_REG_8__SCAN_IN), .S(n8890), .Z(
        P1_U3563) );
  MUX2_X1 U10246 ( .A(n8884), .B(P1_DATAO_REG_7__SCAN_IN), .S(n8890), .Z(
        P1_U3562) );
  MUX2_X1 U10247 ( .A(n8885), .B(P1_DATAO_REG_6__SCAN_IN), .S(n8890), .Z(
        P1_U3561) );
  MUX2_X1 U10248 ( .A(n8886), .B(P1_DATAO_REG_5__SCAN_IN), .S(n8890), .Z(
        P1_U3560) );
  MUX2_X1 U10249 ( .A(n8887), .B(P1_DATAO_REG_4__SCAN_IN), .S(n8890), .Z(
        P1_U3559) );
  MUX2_X1 U10250 ( .A(n8888), .B(P1_DATAO_REG_3__SCAN_IN), .S(n8890), .Z(
        P1_U3558) );
  MUX2_X1 U10251 ( .A(n8889), .B(P1_DATAO_REG_2__SCAN_IN), .S(n8890), .Z(
        P1_U3557) );
  MUX2_X1 U10252 ( .A(n8891), .B(P1_DATAO_REG_1__SCAN_IN), .S(n8890), .Z(
        P1_U3556) );
  MUX2_X1 U10253 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n8892), .S(P1_U4006), .Z(
        P1_U3555) );
  NOR2_X1 U10254 ( .A1(n8900), .A2(n8893), .ZN(n8895) );
  NAND2_X1 U10255 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n8919), .ZN(n8896) );
  OAI21_X1 U10256 ( .B1(n8919), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8896), .ZN(
        n8897) );
  NOR2_X1 U10257 ( .A1(n8898), .A2(n8897), .ZN(n8914) );
  AOI211_X1 U10258 ( .C1(n8898), .C2(n8897), .A(n8914), .B(n9623), .ZN(n8910)
         );
  NOR2_X1 U10259 ( .A1(n8900), .A2(n8899), .ZN(n8902) );
  NOR2_X1 U10260 ( .A1(n8902), .A2(n8901), .ZN(n8904) );
  XNOR2_X1 U10261 ( .A(n8919), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n8903) );
  NOR2_X1 U10262 ( .A1(n8904), .A2(n8903), .ZN(n8918) );
  AOI211_X1 U10263 ( .C1(n8904), .C2(n8903), .A(n8918), .B(n9549), .ZN(n8909)
         );
  NAND2_X1 U10264 ( .A1(n9634), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n8906) );
  NAND2_X1 U10265 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n8905) );
  OAI211_X1 U10266 ( .C1(n9543), .C2(n8907), .A(n8906), .B(n8905), .ZN(n8908)
         );
  OR3_X1 U10267 ( .A1(n8910), .A2(n8909), .A3(n8908), .ZN(P1_U3257) );
  INV_X1 U10268 ( .A(n8930), .ZN(n8913) );
  NAND2_X1 U10269 ( .A1(n9634), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n8912) );
  NAND2_X1 U10270 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n8911) );
  OAI211_X1 U10271 ( .C1(n9543), .C2(n8913), .A(n8912), .B(n8911), .ZN(n8924)
         );
  AOI21_X1 U10272 ( .B1(n8919), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8914), .ZN(
        n8917) );
  NAND2_X1 U10273 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n8930), .ZN(n8915) );
  OAI21_X1 U10274 ( .B1(n8930), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8915), .ZN(
        n8916) );
  NOR2_X1 U10275 ( .A1(n8917), .A2(n8916), .ZN(n8925) );
  AOI211_X1 U10276 ( .C1(n8917), .C2(n8916), .A(n8925), .B(n9623), .ZN(n8923)
         );
  AOI21_X1 U10277 ( .B1(n8919), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8918), .ZN(
        n8921) );
  XNOR2_X1 U10278 ( .A(n8930), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n8920) );
  NOR2_X1 U10279 ( .A1(n8921), .A2(n8920), .ZN(n8929) );
  AOI211_X1 U10280 ( .C1(n8921), .C2(n8920), .A(n8929), .B(n9549), .ZN(n8922)
         );
  OR3_X1 U10281 ( .A1(n8924), .A2(n8923), .A3(n8922), .ZN(P1_U3258) );
  INV_X1 U10282 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9947) );
  NAND2_X1 U10283 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n9630), .ZN(n8926) );
  OAI21_X1 U10284 ( .B1(n9630), .B2(P1_REG2_REG_18__SCAN_IN), .A(n8926), .ZN(
        n9625) );
  INV_X1 U10285 ( .A(n8936), .ZN(n8934) );
  INV_X1 U10286 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8927) );
  AOI22_X1 U10287 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n9630), .B1(n8928), .B2(
        n8927), .ZN(n9633) );
  AOI21_X1 U10288 ( .B1(n8930), .B2(P1_REG1_REG_17__SCAN_IN), .A(n8929), .ZN(
        n9632) );
  NAND2_X1 U10289 ( .A1(n9633), .A2(n9632), .ZN(n9631) );
  OAI21_X1 U10290 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9630), .A(n9631), .ZN(
        n8932) );
  XOR2_X1 U10291 ( .A(n8932), .B(n8931), .Z(n8935) );
  OAI21_X1 U10292 ( .B1(n8935), .B2(n9549), .A(n9543), .ZN(n8933) );
  AOI21_X1 U10293 ( .B1(n8934), .B2(n9616), .A(n8933), .ZN(n8938) );
  AOI22_X1 U10294 ( .A1(n8936), .A2(n9616), .B1(n9635), .B2(n8935), .ZN(n8937)
         );
  MUX2_X1 U10295 ( .A(n8938), .B(n8937), .S(n9646), .Z(n8940) );
  NAND2_X1 U10296 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3084), .ZN(n8939) );
  OAI211_X1 U10297 ( .C1(n4667), .C2(n9621), .A(n8940), .B(n8939), .ZN(
        P1_U3260) );
  NAND2_X1 U10298 ( .A1(n8941), .A2(n9228), .ZN(n9223) );
  NAND2_X1 U10299 ( .A1(n9248), .A2(n9012), .ZN(n9244) );
  XNOR2_X1 U10300 ( .A(n9240), .B(n9244), .ZN(n9243) );
  NAND2_X1 U10301 ( .A1(n9490), .A2(P1_B_REG_SCAN_IN), .ZN(n8943) );
  AND2_X1 U10302 ( .A1(n9232), .A2(n8943), .ZN(n9008) );
  NAND2_X1 U10303 ( .A1(n8944), .A2(n9008), .ZN(n9246) );
  NOR2_X1 U10304 ( .A1(n9405), .A2(n9246), .ZN(n8950) );
  NOR2_X1 U10305 ( .A1(n8945), .A2(n9217), .ZN(n8946) );
  AOI211_X1 U10306 ( .C1(n9405), .C2(P1_REG2_REG_31__SCAN_IN), .A(n8950), .B(
        n8946), .ZN(n8947) );
  OAI21_X1 U10307 ( .B1(n9243), .B2(n8948), .A(n8947), .ZN(P1_U3261) );
  NAND2_X1 U10308 ( .A1(n8949), .A2(n4482), .ZN(n9245) );
  NAND3_X1 U10309 ( .A1(n9245), .A2(n9237), .A3(n9244), .ZN(n8952) );
  AOI21_X1 U10310 ( .B1(n9405), .B2(P1_REG2_REG_30__SCAN_IN), .A(n8950), .ZN(
        n8951) );
  OAI211_X1 U10311 ( .C1(n9248), .C2(n9217), .A(n8952), .B(n8951), .ZN(
        P1_U3262) );
  AOI21_X1 U10312 ( .B1(n9228), .B2(n9210), .A(n9221), .ZN(n8957) );
  OAI21_X1 U10313 ( .B1(n9203), .B2(n9206), .A(n8959), .ZN(n9190) );
  INV_X1 U10314 ( .A(n9190), .ZN(n8960) );
  NOR2_X1 U10315 ( .A1(n9302), .A2(n9183), .ZN(n8962) );
  INV_X1 U10316 ( .A(n9297), .ZN(n9148) );
  NAND2_X1 U10317 ( .A1(n4302), .A2(n9133), .ZN(n9131) );
  NAND2_X1 U10318 ( .A1(n9131), .A2(n4356), .ZN(n9117) );
  OAI21_X1 U10319 ( .B1(n9287), .B2(n9106), .A(n9117), .ZN(n8965) );
  NAND2_X1 U10320 ( .A1(n8965), .A2(n4357), .ZN(n9098) );
  NAND2_X1 U10321 ( .A1(n9105), .A2(n8966), .ZN(n8968) );
  NAND2_X1 U10322 ( .A1(n9090), .A2(n8969), .ZN(n8970) );
  NAND2_X1 U10323 ( .A1(n9056), .A2(n8974), .ZN(n8976) );
  NAND2_X1 U10324 ( .A1(n8976), .A2(n8975), .ZN(n9040) );
  NAND2_X1 U10325 ( .A1(n9044), .A2(n9024), .ZN(n8977) );
  XNOR2_X1 U10326 ( .A(n8980), .B(n8979), .ZN(n9249) );
  INV_X1 U10327 ( .A(n9249), .ZN(n9020) );
  NAND2_X1 U10328 ( .A1(n9205), .A2(n8984), .ZN(n8986) );
  NAND2_X1 U10329 ( .A1(n9180), .A2(n8989), .ZN(n9165) );
  NAND2_X1 U10330 ( .A1(n9165), .A2(n9166), .ZN(n9164) );
  INV_X1 U10331 ( .A(n9149), .ZN(n8990) );
  NOR2_X1 U10332 ( .A1(n9151), .A2(n8990), .ZN(n8991) );
  NAND2_X1 U10333 ( .A1(n9124), .A2(n8994), .ZN(n8996) );
  NAND2_X1 U10334 ( .A1(n8996), .A2(n8995), .ZN(n9109) );
  AOI21_X1 U10335 ( .B1(n9063), .B2(n9000), .A(n8999), .ZN(n9045) );
  NAND2_X1 U10336 ( .A1(n9045), .A2(n9046), .ZN(n9051) );
  NAND2_X1 U10337 ( .A1(n9051), .A2(n9001), .ZN(n9022) );
  INV_X1 U10338 ( .A(n9002), .ZN(n9004) );
  XNOR2_X1 U10339 ( .A(n9006), .B(n9005), .ZN(n9011) );
  AOI22_X1 U10340 ( .A1(n9009), .A2(n9231), .B1(n9008), .B2(n9007), .ZN(n9010)
         );
  OAI21_X1 U10341 ( .B1(n9011), .B2(n9208), .A(n9010), .ZN(n9250) );
  INV_X1 U10342 ( .A(n9252), .ZN(n9017) );
  NOR2_X1 U10343 ( .A1(n9405), .A2(n4797), .ZN(n9187) );
  NAND2_X1 U10344 ( .A1(n9251), .A2(n9187), .ZN(n9016) );
  INV_X1 U10345 ( .A(n9013), .ZN(n9014) );
  AOI22_X1 U10346 ( .A1(n9014), .A2(n9404), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9405), .ZN(n9015) );
  OAI211_X1 U10347 ( .C1(n9017), .C2(n9217), .A(n9016), .B(n9015), .ZN(n9018)
         );
  AOI21_X1 U10348 ( .B1(n9250), .B2(n9653), .A(n9018), .ZN(n9019) );
  OAI21_X1 U10349 ( .B1(n9020), .B2(n9239), .A(n9019), .ZN(P1_U3355) );
  INV_X1 U10350 ( .A(n9027), .ZN(n9021) );
  XNOR2_X1 U10351 ( .A(n9022), .B(n9021), .ZN(n9026) );
  OAI22_X1 U10352 ( .A1(n9024), .A2(n9392), .B1(n9023), .B2(n9394), .ZN(n9025)
         );
  AOI21_X1 U10353 ( .B1(n9026), .B2(n9401), .A(n9025), .ZN(n9259) );
  NAND2_X1 U10354 ( .A1(n9028), .A2(n9027), .ZN(n9029) );
  NAND2_X1 U10355 ( .A1(n9255), .A2(n9030), .ZN(n9039) );
  NAND2_X1 U10356 ( .A1(n9256), .A2(n9041), .ZN(n9032) );
  NAND2_X1 U10357 ( .A1(n9256), .A2(n9406), .ZN(n9036) );
  AOI22_X1 U10358 ( .A1(n9034), .A2(n9404), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9405), .ZN(n9035) );
  NAND2_X1 U10359 ( .A1(n9036), .A2(n9035), .ZN(n9037) );
  AOI21_X1 U10360 ( .B1(n9257), .B2(n9237), .A(n9037), .ZN(n9038) );
  OAI211_X1 U10361 ( .C1(n9405), .C2(n9259), .A(n9039), .B(n9038), .ZN(
        P1_U3263) );
  XOR2_X1 U10362 ( .A(n9040), .B(n9046), .Z(n9266) );
  AOI21_X1 U10363 ( .B1(n9262), .B2(n9057), .A(n9031), .ZN(n9263) );
  AOI22_X1 U10364 ( .A1(n9042), .A2(n9404), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9405), .ZN(n9043) );
  OAI21_X1 U10365 ( .B1(n9044), .B2(n9217), .A(n9043), .ZN(n9054) );
  INV_X1 U10366 ( .A(n9045), .ZN(n9047) );
  AOI21_X1 U10367 ( .B1(n9047), .B2(n4700), .A(n9208), .ZN(n9052) );
  OAI22_X1 U10368 ( .A1(n9049), .A2(n9394), .B1(n9048), .B2(n9392), .ZN(n9050)
         );
  AOI21_X1 U10369 ( .B1(n9052), .B2(n9051), .A(n9050), .ZN(n9265) );
  NOR2_X1 U10370 ( .A1(n9265), .A2(n9405), .ZN(n9053) );
  AOI211_X1 U10371 ( .C1(n9237), .C2(n9263), .A(n9054), .B(n9053), .ZN(n9055)
         );
  OAI21_X1 U10372 ( .B1(n9266), .B2(n9239), .A(n9055), .ZN(P1_U3264) );
  XOR2_X1 U10373 ( .A(n9065), .B(n9056), .Z(n9271) );
  INV_X1 U10374 ( .A(n9057), .ZN(n9058) );
  AOI21_X1 U10375 ( .B1(n9267), .B2(n4479), .A(n9058), .ZN(n9268) );
  AOI22_X1 U10376 ( .A1(n9059), .A2(n9404), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9405), .ZN(n9060) );
  OAI21_X1 U10377 ( .B1(n9061), .B2(n9217), .A(n9060), .ZN(n9069) );
  NAND2_X1 U10378 ( .A1(n9063), .A2(n9062), .ZN(n9064) );
  XOR2_X1 U10379 ( .A(n9065), .B(n9064), .Z(n9067) );
  AOI222_X1 U10380 ( .A1(n9401), .A2(n9067), .B1(n9066), .B2(n9232), .C1(n8972), .C2(n9231), .ZN(n9270) );
  NOR2_X1 U10381 ( .A1(n9270), .A2(n9405), .ZN(n9068) );
  AOI211_X1 U10382 ( .C1(n9237), .C2(n9268), .A(n9069), .B(n9068), .ZN(n9070)
         );
  OAI21_X1 U10383 ( .B1(n9271), .B2(n9239), .A(n9070), .ZN(P1_U3265) );
  XOR2_X1 U10384 ( .A(n9079), .B(n9071), .Z(n9276) );
  AOI21_X1 U10385 ( .B1(n9272), .B2(n9086), .A(n9072), .ZN(n9273) );
  INV_X1 U10386 ( .A(n9073), .ZN(n9074) );
  AOI22_X1 U10387 ( .A1(n9074), .A2(n9404), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9405), .ZN(n9075) );
  OAI21_X1 U10388 ( .B1(n9076), .B2(n9217), .A(n9075), .ZN(n9083) );
  NAND2_X1 U10389 ( .A1(n9091), .A2(n9077), .ZN(n9078) );
  XOR2_X1 U10390 ( .A(n9079), .B(n9078), .Z(n9081) );
  AOI222_X1 U10391 ( .A1(n9401), .A2(n9081), .B1(n9113), .B2(n9231), .C1(n9080), .C2(n9232), .ZN(n9275) );
  NOR2_X1 U10392 ( .A1(n9275), .A2(n9405), .ZN(n9082) );
  AOI211_X1 U10393 ( .C1(n9273), .C2(n9237), .A(n9083), .B(n9082), .ZN(n9084)
         );
  OAI21_X1 U10394 ( .B1(n9276), .B2(n9239), .A(n9084), .ZN(P1_U3266) );
  XNOR2_X1 U10395 ( .A(n9085), .B(n9092), .ZN(n9281) );
  INV_X1 U10396 ( .A(n9086), .ZN(n9087) );
  AOI211_X1 U10397 ( .C1(n9278), .C2(n9099), .A(n9242), .B(n9087), .ZN(n9277)
         );
  AOI22_X1 U10398 ( .A1(n9088), .A2(n9404), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9405), .ZN(n9089) );
  OAI21_X1 U10399 ( .B1(n9090), .B2(n9217), .A(n9089), .ZN(n9096) );
  OAI21_X1 U10400 ( .B1(n9093), .B2(n9092), .A(n9091), .ZN(n9094) );
  AOI222_X1 U10401 ( .A1(n9401), .A2(n9094), .B1(n8972), .B2(n9232), .C1(n9126), .C2(n9231), .ZN(n9280) );
  NOR2_X1 U10402 ( .A1(n9280), .A2(n9405), .ZN(n9095) );
  AOI211_X1 U10403 ( .C1(n9277), .C2(n9187), .A(n9096), .B(n9095), .ZN(n9097)
         );
  OAI21_X1 U10404 ( .B1(n9281), .B2(n9239), .A(n9097), .ZN(P1_U3267) );
  XNOR2_X1 U10405 ( .A(n9098), .B(n9110), .ZN(n9286) );
  INV_X1 U10406 ( .A(n9118), .ZN(n9101) );
  INV_X1 U10407 ( .A(n9099), .ZN(n9100) );
  AOI21_X1 U10408 ( .B1(n9282), .B2(n9101), .A(n9100), .ZN(n9283) );
  INV_X1 U10409 ( .A(n9102), .ZN(n9103) );
  AOI22_X1 U10410 ( .A1(n9103), .A2(n9404), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9405), .ZN(n9104) );
  OAI21_X1 U10411 ( .B1(n9105), .B2(n9217), .A(n9104), .ZN(n9115) );
  AND2_X1 U10412 ( .A1(n9106), .A2(n9231), .ZN(n9112) );
  INV_X1 U10413 ( .A(n9107), .ZN(n9108) );
  AOI211_X1 U10414 ( .C1(n9110), .C2(n9109), .A(n9208), .B(n9108), .ZN(n9111)
         );
  AOI211_X1 U10415 ( .C1(n9232), .C2(n9113), .A(n9112), .B(n9111), .ZN(n9285)
         );
  NOR2_X1 U10416 ( .A1(n9285), .A2(n9405), .ZN(n9114) );
  AOI211_X1 U10417 ( .C1(n9283), .C2(n9237), .A(n9115), .B(n9114), .ZN(n9116)
         );
  OAI21_X1 U10418 ( .B1(n9286), .B2(n9239), .A(n9116), .ZN(P1_U3268) );
  XNOR2_X1 U10419 ( .A(n9117), .B(n9125), .ZN(n9291) );
  INV_X1 U10420 ( .A(n9137), .ZN(n9119) );
  AOI21_X1 U10421 ( .B1(n9287), .B2(n9119), .A(n9118), .ZN(n9288) );
  INV_X1 U10422 ( .A(n9120), .ZN(n9121) );
  AOI22_X1 U10423 ( .A1(n9121), .A2(n9404), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9405), .ZN(n9122) );
  OAI21_X1 U10424 ( .B1(n9123), .B2(n9217), .A(n9122), .ZN(n9129) );
  XOR2_X1 U10425 ( .A(n9125), .B(n9124), .Z(n9127) );
  AOI222_X1 U10426 ( .A1(n9401), .A2(n9127), .B1(n9152), .B2(n9231), .C1(n9126), .C2(n9232), .ZN(n9290) );
  NOR2_X1 U10427 ( .A1(n9290), .A2(n9405), .ZN(n9128) );
  AOI211_X1 U10428 ( .C1(n9288), .C2(n9237), .A(n9129), .B(n9128), .ZN(n9130)
         );
  OAI21_X1 U10429 ( .B1(n9291), .B2(n9239), .A(n9130), .ZN(P1_U3269) );
  OAI21_X1 U10430 ( .B1(n4302), .B2(n9133), .A(n9131), .ZN(n9296) );
  AOI22_X1 U10431 ( .A1(n9294), .A2(n9406), .B1(n9405), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9142) );
  AOI21_X1 U10432 ( .B1(n9133), .B2(n9132), .A(n4323), .ZN(n9134) );
  OAI222_X1 U10433 ( .A1(n9392), .A2(n9136), .B1(n9394), .B2(n9135), .C1(n9208), .C2(n9134), .ZN(n9292) );
  AOI211_X1 U10434 ( .C1(n9294), .C2(n9144), .A(n9242), .B(n9137), .ZN(n9293)
         );
  INV_X1 U10435 ( .A(n9293), .ZN(n9139) );
  OAI22_X1 U10436 ( .A1(n9139), .A2(n4797), .B1(n9644), .B2(n9138), .ZN(n9140)
         );
  OAI21_X1 U10437 ( .B1(n9292), .B2(n9140), .A(n9653), .ZN(n9141) );
  OAI211_X1 U10438 ( .C1(n9296), .C2(n9239), .A(n9142), .B(n9141), .ZN(
        P1_U3270) );
  XNOR2_X1 U10439 ( .A(n9143), .B(n9151), .ZN(n9301) );
  AOI21_X1 U10440 ( .B1(n9297), .B2(n9158), .A(n4470), .ZN(n9298) );
  INV_X1 U10441 ( .A(n9145), .ZN(n9146) );
  AOI22_X1 U10442 ( .A1(n9405), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9146), .B2(
        n9404), .ZN(n9147) );
  OAI21_X1 U10443 ( .B1(n9148), .B2(n9217), .A(n9147), .ZN(n9155) );
  NAND2_X1 U10444 ( .A1(n9164), .A2(n9149), .ZN(n9150) );
  XOR2_X1 U10445 ( .A(n9151), .B(n9150), .Z(n9153) );
  AOI222_X1 U10446 ( .A1(n9401), .A2(n9153), .B1(n9152), .B2(n9232), .C1(n9183), .C2(n9231), .ZN(n9300) );
  NOR2_X1 U10447 ( .A1(n9300), .A2(n9405), .ZN(n9154) );
  AOI211_X1 U10448 ( .C1(n9298), .C2(n9237), .A(n9155), .B(n9154), .ZN(n9156)
         );
  OAI21_X1 U10449 ( .B1(n9301), .B2(n9239), .A(n9156), .ZN(P1_U3271) );
  XNOR2_X1 U10450 ( .A(n9157), .B(n9166), .ZN(n9306) );
  INV_X1 U10451 ( .A(n9174), .ZN(n9159) );
  AOI21_X1 U10452 ( .B1(n9302), .B2(n9159), .A(n4471), .ZN(n9303) );
  INV_X1 U10453 ( .A(n9160), .ZN(n9161) );
  AOI22_X1 U10454 ( .A1(n9405), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9161), .B2(
        n9404), .ZN(n9162) );
  OAI21_X1 U10455 ( .B1(n9163), .B2(n9217), .A(n9162), .ZN(n9170) );
  OAI21_X1 U10456 ( .B1(n9166), .B2(n9165), .A(n9164), .ZN(n9168) );
  AOI222_X1 U10457 ( .A1(n9401), .A2(n9168), .B1(n9167), .B2(n9232), .C1(n9198), .C2(n9231), .ZN(n9305) );
  NOR2_X1 U10458 ( .A1(n9305), .A2(n9405), .ZN(n9169) );
  AOI211_X1 U10459 ( .C1(n9303), .C2(n9237), .A(n9170), .B(n9169), .ZN(n9171)
         );
  OAI21_X1 U10460 ( .B1(n9306), .B2(n9239), .A(n9171), .ZN(P1_U3272) );
  XNOR2_X1 U10461 ( .A(n9173), .B(n9172), .ZN(n9311) );
  INV_X1 U10462 ( .A(n9191), .ZN(n9175) );
  AOI211_X1 U10463 ( .C1(n9308), .C2(n9175), .A(n9242), .B(n9174), .ZN(n9307)
         );
  INV_X1 U10464 ( .A(n9176), .ZN(n9177) );
  AOI22_X1 U10465 ( .A1(n9405), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9177), .B2(
        n9404), .ZN(n9178) );
  OAI21_X1 U10466 ( .B1(n9179), .B2(n9217), .A(n9178), .ZN(n9186) );
  OAI21_X1 U10467 ( .B1(n9181), .B2(n4363), .A(n9180), .ZN(n9184) );
  AOI222_X1 U10468 ( .A1(n9401), .A2(n9184), .B1(n9183), .B2(n9232), .C1(n9182), .C2(n9231), .ZN(n9310) );
  NOR2_X1 U10469 ( .A1(n9310), .A2(n9405), .ZN(n9185) );
  AOI211_X1 U10470 ( .C1(n9307), .C2(n9187), .A(n9186), .B(n9185), .ZN(n9188)
         );
  OAI21_X1 U10471 ( .B1(n9311), .B2(n9239), .A(n9188), .ZN(P1_U3273) );
  XNOR2_X1 U10472 ( .A(n9190), .B(n9189), .ZN(n9316) );
  AOI21_X1 U10473 ( .B1(n9312), .B2(n9212), .A(n9191), .ZN(n9313) );
  INV_X1 U10474 ( .A(n9192), .ZN(n9193) );
  AOI22_X1 U10475 ( .A1(n9405), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9193), .B2(
        n9404), .ZN(n9194) );
  OAI21_X1 U10476 ( .B1(n9195), .B2(n9217), .A(n9194), .ZN(n9201) );
  XNOR2_X1 U10477 ( .A(n9197), .B(n9196), .ZN(n9199) );
  AOI222_X1 U10478 ( .A1(n9401), .A2(n9199), .B1(n9198), .B2(n9232), .C1(n9233), .C2(n9231), .ZN(n9315) );
  NOR2_X1 U10479 ( .A1(n9315), .A2(n9405), .ZN(n9200) );
  AOI211_X1 U10480 ( .C1(n9313), .C2(n9237), .A(n9201), .B(n9200), .ZN(n9202)
         );
  OAI21_X1 U10481 ( .B1(n9316), .B2(n9239), .A(n9202), .ZN(P1_U3274) );
  XNOR2_X1 U10482 ( .A(n9203), .B(n9206), .ZN(n9321) );
  NAND2_X1 U10483 ( .A1(n9205), .A2(n9204), .ZN(n9207) );
  XNOR2_X1 U10484 ( .A(n9207), .B(n9206), .ZN(n9209) );
  OAI222_X1 U10485 ( .A1(n9394), .A2(n9211), .B1(n9392), .B2(n9210), .C1(n9209), .C2(n9208), .ZN(n9317) );
  INV_X1 U10486 ( .A(n9319), .ZN(n9218) );
  INV_X1 U10487 ( .A(n9212), .ZN(n9213) );
  AOI211_X1 U10488 ( .C1(n9319), .C2(n9223), .A(n9242), .B(n9213), .ZN(n9318)
         );
  NAND2_X1 U10489 ( .A1(n9318), .A2(n9412), .ZN(n9216) );
  AOI22_X1 U10490 ( .A1(n9405), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9214), .B2(
        n9404), .ZN(n9215) );
  OAI211_X1 U10491 ( .C1(n9218), .C2(n9217), .A(n9216), .B(n9215), .ZN(n9219)
         );
  AOI21_X1 U10492 ( .B1(n9317), .B2(n9653), .A(n9219), .ZN(n9220) );
  OAI21_X1 U10493 ( .B1(n9321), .B2(n9239), .A(n9220), .ZN(P1_U3275) );
  XNOR2_X1 U10494 ( .A(n9221), .B(n9222), .ZN(n9326) );
  INV_X1 U10495 ( .A(n9223), .ZN(n9224) );
  AOI21_X1 U10496 ( .B1(n9322), .B2(n9225), .A(n9224), .ZN(n9323) );
  AOI22_X1 U10497 ( .A1(n9405), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9226), .B2(
        n9404), .ZN(n9227) );
  OAI21_X1 U10498 ( .B1(n9228), .B2(n9217), .A(n9227), .ZN(n9236) );
  XNOR2_X1 U10499 ( .A(n9230), .B(n9229), .ZN(n9234) );
  AOI222_X1 U10500 ( .A1(n9401), .A2(n9234), .B1(n9233), .B2(n9232), .C1(n4509), .C2(n9231), .ZN(n9325) );
  NOR2_X1 U10501 ( .A1(n9325), .A2(n9405), .ZN(n9235) );
  AOI211_X1 U10502 ( .C1(n9323), .C2(n9237), .A(n9236), .B(n9235), .ZN(n9238)
         );
  OAI21_X1 U10503 ( .B1(n9326), .B2(n9239), .A(n9238), .ZN(P1_U3276) );
  NAND2_X1 U10504 ( .A1(n9240), .A2(n9330), .ZN(n9241) );
  OAI211_X1 U10505 ( .C1(n9243), .C2(n9242), .A(n9241), .B(n9246), .ZN(n9335)
         );
  MUX2_X1 U10506 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9335), .S(n9334), .Z(
        P1_U3554) );
  NAND3_X1 U10507 ( .A1(n9245), .A2(n9409), .A3(n9244), .ZN(n9247) );
  OAI211_X1 U10508 ( .C1(n9248), .C2(n9479), .A(n9247), .B(n9246), .ZN(n9336)
         );
  MUX2_X1 U10509 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9336), .S(n9334), .Z(
        P1_U3553) );
  NAND2_X1 U10510 ( .A1(n9249), .A2(n9482), .ZN(n9254) );
  NAND2_X1 U10511 ( .A1(n9254), .A2(n9253), .ZN(n9337) );
  MUX2_X1 U10512 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9337), .S(n9334), .Z(
        P1_U3552) );
  NAND2_X1 U10513 ( .A1(n9255), .A2(n9482), .ZN(n9261) );
  AOI22_X1 U10514 ( .A1(n9257), .A2(n9409), .B1(n9330), .B2(n9256), .ZN(n9258)
         );
  AND2_X1 U10515 ( .A1(n9259), .A2(n9258), .ZN(n9260) );
  NAND2_X1 U10516 ( .A1(n9261), .A2(n9260), .ZN(n9338) );
  MUX2_X1 U10517 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9338), .S(n9334), .Z(
        P1_U3551) );
  AOI22_X1 U10518 ( .A1(n9263), .A2(n9409), .B1(n9330), .B2(n9262), .ZN(n9264)
         );
  OAI211_X1 U10519 ( .C1(n9266), .C2(n9332), .A(n9265), .B(n9264), .ZN(n9339)
         );
  MUX2_X1 U10520 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9339), .S(n9334), .Z(
        P1_U3550) );
  AOI22_X1 U10521 ( .A1(n9268), .A2(n9409), .B1(n9330), .B2(n9267), .ZN(n9269)
         );
  OAI211_X1 U10522 ( .C1(n9271), .C2(n9332), .A(n9270), .B(n9269), .ZN(n9340)
         );
  MUX2_X1 U10523 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9340), .S(n9334), .Z(
        P1_U3549) );
  AOI22_X1 U10524 ( .A1(n9273), .A2(n9409), .B1(n9330), .B2(n9272), .ZN(n9274)
         );
  OAI211_X1 U10525 ( .C1(n9276), .C2(n9332), .A(n9275), .B(n9274), .ZN(n9341)
         );
  MUX2_X1 U10526 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9341), .S(n9334), .Z(
        P1_U3548) );
  AOI21_X1 U10527 ( .B1(n9330), .B2(n9278), .A(n9277), .ZN(n9279) );
  OAI211_X1 U10528 ( .C1(n9281), .C2(n9332), .A(n9280), .B(n9279), .ZN(n9342)
         );
  MUX2_X1 U10529 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9342), .S(n9334), .Z(
        P1_U3547) );
  AOI22_X1 U10530 ( .A1(n9283), .A2(n9409), .B1(n9330), .B2(n9282), .ZN(n9284)
         );
  OAI211_X1 U10531 ( .C1(n9286), .C2(n9332), .A(n9285), .B(n9284), .ZN(n9343)
         );
  MUX2_X1 U10532 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9343), .S(n9334), .Z(
        P1_U3546) );
  AOI22_X1 U10533 ( .A1(n9288), .A2(n9409), .B1(n9330), .B2(n9287), .ZN(n9289)
         );
  OAI211_X1 U10534 ( .C1(n9291), .C2(n9332), .A(n9290), .B(n9289), .ZN(n9344)
         );
  MUX2_X1 U10535 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9344), .S(n9334), .Z(
        P1_U3545) );
  AOI211_X1 U10536 ( .C1(n9330), .C2(n9294), .A(n9293), .B(n9292), .ZN(n9295)
         );
  OAI21_X1 U10537 ( .B1(n9296), .B2(n9332), .A(n9295), .ZN(n9345) );
  MUX2_X1 U10538 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9345), .S(n9334), .Z(
        P1_U3544) );
  AOI22_X1 U10539 ( .A1(n9298), .A2(n9409), .B1(n9330), .B2(n9297), .ZN(n9299)
         );
  OAI211_X1 U10540 ( .C1(n9301), .C2(n9332), .A(n9300), .B(n9299), .ZN(n9346)
         );
  MUX2_X1 U10541 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9346), .S(n9334), .Z(
        P1_U3543) );
  AOI22_X1 U10542 ( .A1(n9303), .A2(n9409), .B1(n9330), .B2(n9302), .ZN(n9304)
         );
  OAI211_X1 U10543 ( .C1(n9306), .C2(n9332), .A(n9305), .B(n9304), .ZN(n9347)
         );
  MUX2_X1 U10544 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9347), .S(n9334), .Z(
        P1_U3542) );
  AOI21_X1 U10545 ( .B1(n9330), .B2(n9308), .A(n9307), .ZN(n9309) );
  OAI211_X1 U10546 ( .C1(n9311), .C2(n9332), .A(n9310), .B(n9309), .ZN(n9348)
         );
  MUX2_X1 U10547 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9348), .S(n9334), .Z(
        P1_U3541) );
  AOI22_X1 U10548 ( .A1(n9313), .A2(n9409), .B1(n9330), .B2(n9312), .ZN(n9314)
         );
  OAI211_X1 U10549 ( .C1(n9316), .C2(n9332), .A(n9315), .B(n9314), .ZN(n9349)
         );
  MUX2_X1 U10550 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9349), .S(n9334), .Z(
        P1_U3540) );
  AOI211_X1 U10551 ( .C1(n9330), .C2(n9319), .A(n9318), .B(n9317), .ZN(n9320)
         );
  OAI21_X1 U10552 ( .B1(n9321), .B2(n9332), .A(n9320), .ZN(n9350) );
  MUX2_X1 U10553 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9350), .S(n9334), .Z(
        P1_U3539) );
  AOI22_X1 U10554 ( .A1(n9323), .A2(n9409), .B1(n9330), .B2(n9322), .ZN(n9324)
         );
  OAI211_X1 U10555 ( .C1(n9326), .C2(n9332), .A(n9325), .B(n9324), .ZN(n9351)
         );
  MUX2_X1 U10556 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9351), .S(n9334), .Z(
        P1_U3538) );
  AOI211_X1 U10557 ( .C1(n9330), .C2(n9329), .A(n9328), .B(n9327), .ZN(n9331)
         );
  OAI21_X1 U10558 ( .B1(n9333), .B2(n9332), .A(n9331), .ZN(n9353) );
  MUX2_X1 U10559 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9353), .S(n9334), .Z(
        P1_U3536) );
  MUX2_X1 U10560 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9335), .S(n9352), .Z(
        P1_U3522) );
  MUX2_X1 U10561 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9336), .S(n9352), .Z(
        P1_U3521) );
  MUX2_X1 U10562 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9337), .S(n9352), .Z(
        P1_U3520) );
  MUX2_X1 U10563 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9338), .S(n9352), .Z(
        P1_U3519) );
  MUX2_X1 U10564 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9339), .S(n9352), .Z(
        P1_U3518) );
  MUX2_X1 U10565 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9340), .S(n9352), .Z(
        P1_U3517) );
  MUX2_X1 U10566 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9341), .S(n9352), .Z(
        P1_U3516) );
  MUX2_X1 U10567 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9342), .S(n9352), .Z(
        P1_U3515) );
  MUX2_X1 U10568 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9343), .S(n9352), .Z(
        P1_U3514) );
  MUX2_X1 U10569 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9344), .S(n9352), .Z(
        P1_U3513) );
  MUX2_X1 U10570 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9345), .S(n9352), .Z(
        P1_U3512) );
  MUX2_X1 U10571 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9346), .S(n9352), .Z(
        P1_U3511) );
  MUX2_X1 U10572 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9347), .S(n9352), .Z(
        P1_U3510) );
  MUX2_X1 U10573 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9348), .S(n9352), .Z(
        P1_U3508) );
  MUX2_X1 U10574 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9349), .S(n9352), .Z(
        P1_U3505) );
  MUX2_X1 U10575 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9350), .S(n9352), .Z(
        P1_U3502) );
  MUX2_X1 U10576 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9351), .S(n9352), .Z(
        P1_U3499) );
  MUX2_X1 U10577 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9353), .S(n9352), .Z(
        P1_U3493) );
  INV_X1 U10578 ( .A(n9354), .ZN(n9359) );
  NOR4_X1 U10579 ( .A1(n9355), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n5332), .ZN(n9356) );
  AOI21_X1 U10580 ( .B1(n9357), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9356), .ZN(
        n9358) );
  OAI21_X1 U10581 ( .B1(n9359), .B2(n9364), .A(n9358), .ZN(P1_U3322) );
  OAI222_X1 U10582 ( .A1(n9364), .A2(n9363), .B1(n9362), .B2(P1_U3084), .C1(
        n9361), .C2(n9360), .ZN(P1_U3324) );
  MUX2_X1 U10583 ( .A(n9365), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10584 ( .A1(n9697), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9376) );
  AOI211_X1 U10585 ( .C1(n9368), .C2(n9367), .A(n9366), .B(n9700), .ZN(n9369)
         );
  AOI21_X1 U10586 ( .B1(n9382), .B2(n9370), .A(n9369), .ZN(n9375) );
  AND2_X1 U10587 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9373) );
  OAI211_X1 U10588 ( .C1(n9373), .C2(n9372), .A(n9695), .B(n9371), .ZN(n9374)
         );
  NAND3_X1 U10589 ( .A1(n9376), .A2(n9375), .A3(n9374), .ZN(P2_U3246) );
  AOI22_X1 U10590 ( .A1(n9697), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9388) );
  AOI211_X1 U10591 ( .C1(n9379), .C2(n9378), .A(n9377), .B(n9700), .ZN(n9380)
         );
  AOI21_X1 U10592 ( .B1(n9382), .B2(n9381), .A(n9380), .ZN(n9387) );
  OAI211_X1 U10593 ( .C1(n9385), .C2(n9384), .A(n9695), .B(n9383), .ZN(n9386)
         );
  NAND3_X1 U10594 ( .A1(n9388), .A2(n9387), .A3(n9386), .ZN(P2_U3247) );
  NAND2_X1 U10595 ( .A1(n9390), .A2(n9389), .ZN(n9391) );
  XOR2_X1 U10596 ( .A(n9396), .B(n9391), .Z(n9402) );
  OAI22_X1 U10597 ( .A1(n9395), .A2(n9394), .B1(n9393), .B2(n9392), .ZN(n9400)
         );
  XOR2_X1 U10598 ( .A(n9397), .B(n9396), .Z(n9408) );
  NOR2_X1 U10599 ( .A1(n9408), .A2(n9398), .ZN(n9399) );
  AOI211_X1 U10600 ( .C1(n9402), .C2(n9401), .A(n9400), .B(n9399), .ZN(n9418)
         );
  AOI222_X1 U10601 ( .A1(n9407), .A2(n9406), .B1(P1_REG2_REG_10__SCAN_IN), 
        .B2(n9405), .C1(n9404), .C2(n9403), .ZN(n9415) );
  INV_X1 U10602 ( .A(n9408), .ZN(n9421) );
  OAI211_X1 U10603 ( .C1(n9417), .C2(n4366), .A(n9410), .B(n9409), .ZN(n9416)
         );
  INV_X1 U10604 ( .A(n9416), .ZN(n9411) );
  AOI22_X1 U10605 ( .A1(n9421), .A2(n9413), .B1(n9412), .B2(n9411), .ZN(n9414)
         );
  OAI211_X1 U10606 ( .C1(n9405), .C2(n9418), .A(n9415), .B(n9414), .ZN(
        P1_U3281) );
  INV_X1 U10607 ( .A(n9663), .ZN(n9422) );
  OAI21_X1 U10608 ( .B1(n9417), .B2(n9479), .A(n9416), .ZN(n9420) );
  INV_X1 U10609 ( .A(n9418), .ZN(n9419) );
  AOI211_X1 U10610 ( .C1(n9422), .C2(n9421), .A(n9420), .B(n9419), .ZN(n9424)
         );
  INV_X1 U10611 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9423) );
  AOI22_X1 U10612 ( .A1(n9352), .A2(n9424), .B1(n9423), .B2(n9669), .ZN(
        P1_U3484) );
  AOI22_X1 U10613 ( .A1(n9334), .A2(n9424), .B1(n6374), .B2(n9671), .ZN(
        P1_U3533) );
  INV_X1 U10614 ( .A(n9425), .ZN(n9426) );
  AOI21_X1 U10615 ( .B1(n9428), .B2(n9427), .A(n9426), .ZN(n9437) );
  NAND2_X1 U10616 ( .A1(n9430), .A2(n9429), .ZN(n9432) );
  AOI21_X1 U10617 ( .B1(n9433), .B2(n9432), .A(n9431), .ZN(n9434) );
  AOI21_X1 U10618 ( .B1(n9435), .B2(n9449), .A(n9434), .ZN(n9436) );
  OAI211_X1 U10619 ( .C1(n9693), .C2(n9438), .A(n9437), .B(n9436), .ZN(
        P2_U3217) );
  OAI21_X1 U10620 ( .B1(n4436), .B2(n9799), .A(n9439), .ZN(n9440) );
  AOI21_X1 U10621 ( .B1(n9441), .B2(n9791), .A(n9440), .ZN(n9464) );
  INV_X1 U10622 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9442) );
  AOI22_X1 U10623 ( .A1(n9830), .A2(n9464), .B1(n9442), .B2(n9828), .ZN(
        P2_U3550) );
  OAI22_X1 U10624 ( .A1(n9444), .A2(n9801), .B1(n9443), .B2(n9799), .ZN(n9446)
         );
  AOI211_X1 U10625 ( .C1(n9806), .C2(n9447), .A(n9446), .B(n9445), .ZN(n9466)
         );
  AOI22_X1 U10626 ( .A1(n9830), .A2(n9466), .B1(n9448), .B2(n9828), .ZN(
        P2_U3535) );
  NAND2_X1 U10627 ( .A1(n9449), .A2(n9790), .ZN(n9450) );
  OAI211_X1 U10628 ( .C1(n9801), .C2(n9452), .A(n9451), .B(n9450), .ZN(n9453)
         );
  AOI21_X1 U10629 ( .B1(n9454), .B2(n9806), .A(n9453), .ZN(n9468) );
  AOI22_X1 U10630 ( .A1(n9830), .A2(n9468), .B1(n9455), .B2(n9828), .ZN(
        P2_U3534) );
  INV_X1 U10631 ( .A(n9456), .ZN(n9787) );
  OAI22_X1 U10632 ( .A1(n9458), .A2(n9801), .B1(n9457), .B2(n9799), .ZN(n9460)
         );
  AOI211_X1 U10633 ( .C1(n9787), .C2(n9461), .A(n9460), .B(n9459), .ZN(n9470)
         );
  AOI22_X1 U10634 ( .A1(n9830), .A2(n9470), .B1(n9462), .B2(n9828), .ZN(
        P2_U3533) );
  INV_X1 U10635 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9463) );
  AOI22_X1 U10636 ( .A1(n9809), .A2(n9464), .B1(n9463), .B2(n9807), .ZN(
        P2_U3518) );
  INV_X1 U10637 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9465) );
  AOI22_X1 U10638 ( .A1(n9809), .A2(n9466), .B1(n9465), .B2(n9807), .ZN(
        P2_U3496) );
  INV_X1 U10639 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9467) );
  AOI22_X1 U10640 ( .A1(n9809), .A2(n9468), .B1(n9467), .B2(n9807), .ZN(
        P2_U3493) );
  INV_X1 U10641 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9469) );
  AOI22_X1 U10642 ( .A1(n9809), .A2(n9470), .B1(n9469), .B2(n9807), .ZN(
        P2_U3490) );
  OAI211_X1 U10643 ( .C1(n9473), .C2(n9479), .A(n9472), .B(n9471), .ZN(n9474)
         );
  AOI21_X1 U10644 ( .B1(n9475), .B2(n9482), .A(n9474), .ZN(n9485) );
  AOI22_X1 U10645 ( .A1(n9334), .A2(n9485), .B1(n9476), .B2(n9671), .ZN(
        P1_U3537) );
  OAI211_X1 U10646 ( .C1(n9480), .C2(n9479), .A(n9478), .B(n9477), .ZN(n9481)
         );
  AOI21_X1 U10647 ( .B1(n9483), .B2(n9482), .A(n9481), .ZN(n9487) );
  AOI22_X1 U10648 ( .A1(n9334), .A2(n9487), .B1(n6603), .B2(n9671), .ZN(
        P1_U3535) );
  INV_X1 U10649 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9484) );
  AOI22_X1 U10650 ( .A1(n9352), .A2(n9485), .B1(n9484), .B2(n9669), .ZN(
        P1_U3496) );
  INV_X1 U10651 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9486) );
  AOI22_X1 U10652 ( .A1(n9352), .A2(n9487), .B1(n9486), .B2(n9669), .ZN(
        P1_U3490) );
  INV_X1 U10653 ( .A(P1_WR_REG_SCAN_IN), .ZN(n10021) );
  XOR2_X1 U10654 ( .A(n10021), .B(P2_WR_REG_SCAN_IN), .Z(U123) );
  XNOR2_X1 U10655 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10656 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9919) );
  AOI21_X1 U10657 ( .B1(n9489), .B2(n9490), .A(n9488), .ZN(n9525) );
  OAI21_X1 U10658 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n9490), .A(n9525), .ZN(
        n9491) );
  XNOR2_X1 U10659 ( .A(n9491), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9493) );
  AOI22_X1 U10660 ( .A1(n9493), .A2(n9492), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3084), .ZN(n9494) );
  OAI21_X1 U10661 ( .B1(n9621), .B2(n9919), .A(n9494), .ZN(P1_U3241) );
  INV_X1 U10662 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9496) );
  OAI22_X1 U10663 ( .A1(n9621), .A2(n9496), .B1(n9543), .B2(n9495), .ZN(n9497)
         );
  INV_X1 U10664 ( .A(n9497), .ZN(n9507) );
  AOI211_X1 U10665 ( .C1(n9500), .C2(n9499), .A(n9498), .B(n9623), .ZN(n9505)
         );
  NAND2_X1 U10666 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9503) );
  AOI211_X1 U10667 ( .C1(n9503), .C2(n9502), .A(n9501), .B(n9549), .ZN(n9504)
         );
  AOI211_X1 U10668 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(P1_U3084), .A(n9505), 
        .B(n9504), .ZN(n9506) );
  NAND2_X1 U10669 ( .A1(n9507), .A2(n9506), .ZN(P1_U3242) );
  INV_X1 U10670 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9509) );
  OAI22_X1 U10671 ( .A1(n9621), .A2(n9509), .B1(n9543), .B2(n9508), .ZN(n9510)
         );
  INV_X1 U10672 ( .A(n9510), .ZN(n9527) );
  AOI211_X1 U10673 ( .C1(n9513), .C2(n9512), .A(n9511), .B(n9623), .ZN(n9518)
         );
  AOI211_X1 U10674 ( .C1(n9516), .C2(n9515), .A(n9514), .B(n9549), .ZN(n9517)
         );
  AOI211_X1 U10675 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(P1_U3084), .A(n9518), 
        .B(n9517), .ZN(n9526) );
  INV_X1 U10676 ( .A(n9519), .ZN(n9520) );
  MUX2_X1 U10677 ( .A(n9521), .B(n9520), .S(n6285), .Z(n9523) );
  NAND2_X1 U10678 ( .A1(n9523), .A2(n9522), .ZN(n9524) );
  OAI211_X1 U10679 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9525), .A(n9524), .B(
        P1_U4006), .ZN(n9539) );
  NAND3_X1 U10680 ( .A1(n9527), .A2(n9526), .A3(n9539), .ZN(P1_U3243) );
  OAI21_X1 U10681 ( .B1(n9530), .B2(n9529), .A(n9528), .ZN(n9532) );
  AOI22_X1 U10682 ( .A1(n9635), .A2(n9532), .B1(n9531), .B2(n9629), .ZN(n9541)
         );
  OAI21_X1 U10683 ( .B1(n9535), .B2(n9534), .A(n9533), .ZN(n9536) );
  AND2_X1 U10684 ( .A1(n9616), .A2(n9536), .ZN(n9537) );
  AOI211_X1 U10685 ( .C1(P1_ADDR_REG_4__SCAN_IN), .C2(n9634), .A(n9538), .B(
        n9537), .ZN(n9540) );
  NAND3_X1 U10686 ( .A1(n9541), .A2(n9540), .A3(n9539), .ZN(P1_U3245) );
  INV_X1 U10687 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9544) );
  OAI22_X1 U10688 ( .A1(n9621), .A2(n9544), .B1(n9543), .B2(n9542), .ZN(n9545)
         );
  INV_X1 U10689 ( .A(n9545), .ZN(n9557) );
  OAI21_X1 U10690 ( .B1(n9548), .B2(n9547), .A(n9546), .ZN(n9555) );
  AOI211_X1 U10691 ( .C1(n9552), .C2(n9551), .A(n9550), .B(n9549), .ZN(n9553)
         );
  AOI211_X1 U10692 ( .C1(n9616), .C2(n9555), .A(n9554), .B(n9553), .ZN(n9556)
         );
  NAND2_X1 U10693 ( .A1(n9557), .A2(n9556), .ZN(P1_U3246) );
  OAI21_X1 U10694 ( .B1(n9560), .B2(n9559), .A(n9558), .ZN(n9561) );
  AOI22_X1 U10695 ( .A1(n9561), .A2(n9635), .B1(n9634), .B2(
        P1_ADDR_REG_6__SCAN_IN), .ZN(n9569) );
  AOI211_X1 U10696 ( .C1(n9564), .C2(n9563), .A(n9562), .B(n9623), .ZN(n9565)
         );
  AOI211_X1 U10697 ( .C1(n9629), .C2(n9567), .A(n9566), .B(n9565), .ZN(n9568)
         );
  NAND2_X1 U10698 ( .A1(n9569), .A2(n9568), .ZN(P1_U3247) );
  AOI21_X1 U10699 ( .B1(n9629), .B2(n9571), .A(n9570), .ZN(n9581) );
  OAI21_X1 U10700 ( .B1(n9574), .B2(n9573), .A(n9572), .ZN(n9579) );
  OAI21_X1 U10701 ( .B1(n9577), .B2(n9576), .A(n9575), .ZN(n9578) );
  AOI22_X1 U10702 ( .A1(n9579), .A2(n9635), .B1(n9616), .B2(n9578), .ZN(n9580)
         );
  OAI211_X1 U10703 ( .C1(n9621), .C2(n9582), .A(n9581), .B(n9580), .ZN(
        P1_U3248) );
  AOI21_X1 U10704 ( .B1(n9629), .B2(n9584), .A(n9583), .ZN(n9594) );
  OAI21_X1 U10705 ( .B1(n9587), .B2(n9586), .A(n9585), .ZN(n9592) );
  OAI21_X1 U10706 ( .B1(n9590), .B2(n9589), .A(n9588), .ZN(n9591) );
  AOI22_X1 U10707 ( .A1(n9592), .A2(n9635), .B1(n9616), .B2(n9591), .ZN(n9593)
         );
  OAI211_X1 U10708 ( .C1(n9621), .C2(n10037), .A(n9594), .B(n9593), .ZN(
        P1_U3249) );
  AOI211_X1 U10709 ( .C1(n9597), .C2(n9596), .A(n9595), .B(n9623), .ZN(n9598)
         );
  AOI211_X1 U10710 ( .C1(n9629), .C2(n9600), .A(n9599), .B(n9598), .ZN(n9606)
         );
  OAI21_X1 U10711 ( .B1(n9603), .B2(n9602), .A(n9601), .ZN(n9604) );
  NAND2_X1 U10712 ( .A1(n9604), .A2(n9635), .ZN(n9605) );
  OAI211_X1 U10713 ( .C1(n10067), .C2(n9621), .A(n9606), .B(n9605), .ZN(
        P1_U3250) );
  INV_X1 U10714 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9620) );
  AOI21_X1 U10715 ( .B1(n9629), .B2(n9608), .A(n9607), .ZN(n9619) );
  OAI21_X1 U10716 ( .B1(n9611), .B2(n9610), .A(n9609), .ZN(n9617) );
  OAI21_X1 U10717 ( .B1(n9614), .B2(n9613), .A(n9612), .ZN(n9615) );
  AOI22_X1 U10718 ( .A1(n9617), .A2(n9616), .B1(n9635), .B2(n9615), .ZN(n9618)
         );
  OAI211_X1 U10719 ( .C1(n9621), .C2(n9620), .A(n9619), .B(n9618), .ZN(
        P1_U3255) );
  INV_X1 U10720 ( .A(n9622), .ZN(n9628) );
  AOI211_X1 U10721 ( .C1(n9626), .C2(n9625), .A(n9624), .B(n9623), .ZN(n9627)
         );
  AOI211_X1 U10722 ( .C1(n9630), .C2(n9629), .A(n9628), .B(n9627), .ZN(n9638)
         );
  OAI21_X1 U10723 ( .B1(n9633), .B2(n9632), .A(n9631), .ZN(n9636) );
  AOI22_X1 U10724 ( .A1(n9636), .A2(n9635), .B1(n9634), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n9637) );
  NAND2_X1 U10725 ( .A1(n9638), .A2(n9637), .ZN(P1_U3259) );
  INV_X1 U10726 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9655) );
  INV_X1 U10727 ( .A(n9639), .ZN(n9650) );
  NAND2_X1 U10728 ( .A1(n9641), .A2(n9640), .ZN(n9642) );
  OAI21_X1 U10729 ( .B1(n9644), .B2(n9643), .A(n9642), .ZN(n9645) );
  AOI21_X1 U10730 ( .B1(n9647), .B2(n9646), .A(n9645), .ZN(n9648) );
  OAI211_X1 U10731 ( .C1(n9651), .C2(n9650), .A(n9649), .B(n9648), .ZN(n9652)
         );
  INV_X1 U10732 ( .A(n9652), .ZN(n9654) );
  AOI22_X1 U10733 ( .A1(n9405), .A2(n9655), .B1(n9654), .B2(n9653), .ZN(
        P1_U3286) );
  AND2_X1 U10734 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9659), .ZN(P1_U3292) );
  AND2_X1 U10735 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9659), .ZN(P1_U3293) );
  AND2_X1 U10736 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9659), .ZN(P1_U3294) );
  AND2_X1 U10737 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9659), .ZN(P1_U3295) );
  AND2_X1 U10738 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9659), .ZN(P1_U3296) );
  AND2_X1 U10739 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9659), .ZN(P1_U3297) );
  AND2_X1 U10740 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9659), .ZN(P1_U3298) );
  AND2_X1 U10741 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9659), .ZN(P1_U3299) );
  NOR2_X1 U10742 ( .A1(n9660), .A2(n9960), .ZN(P1_U3300) );
  AND2_X1 U10743 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9659), .ZN(P1_U3301) );
  AND2_X1 U10744 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9659), .ZN(P1_U3302) );
  AND2_X1 U10745 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9659), .ZN(P1_U3303) );
  NOR2_X1 U10746 ( .A1(n9660), .A2(n9924), .ZN(P1_U3304) );
  AND2_X1 U10747 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9659), .ZN(P1_U3305) );
  AND2_X1 U10748 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9659), .ZN(P1_U3306) );
  AND2_X1 U10749 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9659), .ZN(P1_U3307) );
  AND2_X1 U10750 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9659), .ZN(P1_U3308) );
  AND2_X1 U10751 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9659), .ZN(P1_U3309) );
  AND2_X1 U10752 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9659), .ZN(P1_U3310) );
  AND2_X1 U10753 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9659), .ZN(P1_U3311) );
  AND2_X1 U10754 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9659), .ZN(P1_U3312) );
  AND2_X1 U10755 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9659), .ZN(P1_U3313) );
  AND2_X1 U10756 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9659), .ZN(P1_U3314) );
  AND2_X1 U10757 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9659), .ZN(P1_U3315) );
  AND2_X1 U10758 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9659), .ZN(P1_U3316) );
  INV_X1 U10759 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9863) );
  NOR2_X1 U10760 ( .A1(n9660), .A2(n9863), .ZN(P1_U3317) );
  NOR2_X1 U10761 ( .A1(n9660), .A2(n9996), .ZN(P1_U3318) );
  NOR2_X1 U10762 ( .A1(n9660), .A2(n9658), .ZN(P1_U3319) );
  AND2_X1 U10763 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9659), .ZN(P1_U3320) );
  INV_X1 U10764 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10031) );
  NOR2_X1 U10765 ( .A1(n9660), .A2(n10031), .ZN(P1_U3321) );
  NAND2_X1 U10766 ( .A1(n6453), .A2(n9330), .ZN(n9661) );
  OAI211_X1 U10767 ( .C1(n9664), .C2(n9663), .A(n9662), .B(n9661), .ZN(n9666)
         );
  AOI211_X1 U10768 ( .C1(n9668), .C2(n9667), .A(n9666), .B(n9665), .ZN(n9673)
         );
  INV_X1 U10769 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9670) );
  AOI22_X1 U10770 ( .A1(n9352), .A2(n9673), .B1(n9670), .B2(n9669), .ZN(
        P1_U3457) );
  INV_X1 U10771 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9672) );
  AOI22_X1 U10772 ( .A1(n9334), .A2(n9673), .B1(n9672), .B2(n9671), .ZN(
        P1_U3524) );
  OAI21_X1 U10773 ( .B1(n9676), .B2(n9675), .A(n9674), .ZN(n9680) );
  NAND3_X1 U10774 ( .A1(n9678), .A2(n9677), .A3(n9683), .ZN(n9679) );
  NAND2_X1 U10775 ( .A1(n9680), .A2(n9679), .ZN(n9690) );
  AOI22_X1 U10776 ( .A1(n9684), .A2(n9683), .B1(n9682), .B2(n9681), .ZN(n9686)
         );
  OAI211_X1 U10777 ( .C1(n9769), .C2(n9687), .A(n9686), .B(n9685), .ZN(n9688)
         );
  AOI21_X1 U10778 ( .B1(n9690), .B2(n9689), .A(n9688), .ZN(n9691) );
  OAI21_X1 U10779 ( .B1(n9693), .B2(n9692), .A(n9691), .ZN(P2_U3223) );
  AOI22_X1 U10780 ( .A1(n9695), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9694), .ZN(n9705) );
  AOI22_X1 U10781 ( .A1(n9697), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9704) );
  NOR2_X1 U10782 ( .A1(n9698), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9702) );
  OAI21_X1 U10783 ( .B1(n9700), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9699), .ZN(
        n9701) );
  OAI21_X1 U10784 ( .B1(n9702), .B2(n9701), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9703) );
  OAI211_X1 U10785 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9705), .A(n9704), .B(
        n9703), .ZN(P2_U3245) );
  AND2_X1 U10786 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9861), .ZN(P2_U3298) );
  AND2_X1 U10787 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9861), .ZN(P2_U3299) );
  AND2_X1 U10788 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9861), .ZN(P2_U3300) );
  AND2_X1 U10789 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9861), .ZN(P2_U3301) );
  AND2_X1 U10790 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9861), .ZN(P2_U3302) );
  AND2_X1 U10791 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9861), .ZN(P2_U3303) );
  AND2_X1 U10792 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9861), .ZN(P2_U3304) );
  AND2_X1 U10793 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9861), .ZN(P2_U3305) );
  AND2_X1 U10794 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9861), .ZN(P2_U3306) );
  AND2_X1 U10795 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9861), .ZN(P2_U3307) );
  AND2_X1 U10796 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9861), .ZN(P2_U3308) );
  AND2_X1 U10797 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9861), .ZN(P2_U3309) );
  AND2_X1 U10798 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9861), .ZN(P2_U3310) );
  AND2_X1 U10799 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9861), .ZN(P2_U3311) );
  AND2_X1 U10800 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9861), .ZN(P2_U3312) );
  AND2_X1 U10801 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9861), .ZN(P2_U3313) );
  AND2_X1 U10802 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9861), .ZN(P2_U3314) );
  INV_X1 U10803 ( .A(n9861), .ZN(n9711) );
  INV_X1 U10804 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10038) );
  NOR2_X1 U10805 ( .A1(n9711), .A2(n10038), .ZN(P2_U3315) );
  AND2_X1 U10806 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9861), .ZN(P2_U3316) );
  INV_X1 U10807 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n9934) );
  NOR2_X1 U10808 ( .A1(n9711), .A2(n9934), .ZN(P2_U3317) );
  AND2_X1 U10809 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9861), .ZN(P2_U3318) );
  AND2_X1 U10810 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9861), .ZN(P2_U3319) );
  AND2_X1 U10811 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9861), .ZN(P2_U3320) );
  AND2_X1 U10812 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9861), .ZN(P2_U3321) );
  AND2_X1 U10813 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9861), .ZN(P2_U3322) );
  AND2_X1 U10814 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9861), .ZN(P2_U3323) );
  AND2_X1 U10815 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9861), .ZN(P2_U3324) );
  AND2_X1 U10816 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9861), .ZN(P2_U3325) );
  AND2_X1 U10817 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9861), .ZN(P2_U3326) );
  OAI22_X1 U10818 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n9711), .B1(n9710), .B2(
        n9709), .ZN(n9712) );
  INV_X1 U10819 ( .A(n9712), .ZN(P2_U3437) );
  AOI22_X1 U10820 ( .A1(n9715), .A2(n9714), .B1(n9713), .B2(n9861), .ZN(
        P2_U3438) );
  OAI21_X1 U10821 ( .B1(n5732), .B2(n9717), .A(n9716), .ZN(n9718) );
  AOI21_X1 U10822 ( .B1(n9806), .B2(n9719), .A(n9718), .ZN(n9811) );
  INV_X1 U10823 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9720) );
  AOI22_X1 U10824 ( .A1(n9809), .A2(n9811), .B1(n9720), .B2(n9807), .ZN(
        P2_U3451) );
  OAI211_X1 U10825 ( .C1(n7186), .C2(n9799), .A(n9722), .B(n9721), .ZN(n9723)
         );
  AOI21_X1 U10826 ( .B1(n9806), .B2(n9724), .A(n9723), .ZN(n9812) );
  INV_X1 U10827 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9725) );
  AOI22_X1 U10828 ( .A1(n9809), .A2(n9812), .B1(n9725), .B2(n9807), .ZN(
        P2_U3454) );
  INV_X1 U10829 ( .A(n9726), .ZN(n9727) );
  OAI211_X1 U10830 ( .C1(n9729), .C2(n9799), .A(n9728), .B(n9727), .ZN(n9730)
         );
  AOI21_X1 U10831 ( .B1(n9806), .B2(n9731), .A(n9730), .ZN(n9813) );
  INV_X1 U10832 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9732) );
  AOI22_X1 U10833 ( .A1(n9809), .A2(n9813), .B1(n9732), .B2(n9807), .ZN(
        P2_U3457) );
  INV_X1 U10834 ( .A(n9733), .ZN(n9735) );
  OAI22_X1 U10835 ( .A1(n9735), .A2(n9801), .B1(n9734), .B2(n9799), .ZN(n9738)
         );
  INV_X1 U10836 ( .A(n9736), .ZN(n9737) );
  AOI211_X1 U10837 ( .C1(n9787), .C2(n9739), .A(n9738), .B(n9737), .ZN(n9815)
         );
  INV_X1 U10838 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9740) );
  AOI22_X1 U10839 ( .A1(n9809), .A2(n9815), .B1(n9740), .B2(n9807), .ZN(
        P2_U3460) );
  OAI22_X1 U10840 ( .A1(n9742), .A2(n9801), .B1(n9741), .B2(n9799), .ZN(n9744)
         );
  AOI211_X1 U10841 ( .C1(n9806), .C2(n9745), .A(n9744), .B(n9743), .ZN(n9817)
         );
  INV_X1 U10842 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9746) );
  AOI22_X1 U10843 ( .A1(n9809), .A2(n9817), .B1(n9746), .B2(n9807), .ZN(
        P2_U3463) );
  INV_X1 U10844 ( .A(n9747), .ZN(n9748) );
  OAI211_X1 U10845 ( .C1(n9750), .C2(n9799), .A(n9749), .B(n9748), .ZN(n9751)
         );
  AOI21_X1 U10846 ( .B1(n9806), .B2(n9752), .A(n9751), .ZN(n9819) );
  INV_X1 U10847 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9753) );
  AOI22_X1 U10848 ( .A1(n9809), .A2(n9819), .B1(n9753), .B2(n9807), .ZN(
        P2_U3466) );
  INV_X1 U10849 ( .A(n9754), .ZN(n9760) );
  OAI22_X1 U10850 ( .A1(n9756), .A2(n9801), .B1(n9755), .B2(n9799), .ZN(n9759)
         );
  INV_X1 U10851 ( .A(n9757), .ZN(n9758) );
  AOI211_X1 U10852 ( .C1(n9760), .C2(n9806), .A(n9759), .B(n9758), .ZN(n9821)
         );
  INV_X1 U10853 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9761) );
  AOI22_X1 U10854 ( .A1(n9809), .A2(n9821), .B1(n9761), .B2(n9807), .ZN(
        P2_U3469) );
  OAI22_X1 U10855 ( .A1(n9763), .A2(n9801), .B1(n9762), .B2(n9799), .ZN(n9765)
         );
  AOI211_X1 U10856 ( .C1(n9766), .C2(n9806), .A(n9765), .B(n9764), .ZN(n9823)
         );
  INV_X1 U10857 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9767) );
  AOI22_X1 U10858 ( .A1(n9809), .A2(n9823), .B1(n9767), .B2(n9807), .ZN(
        P2_U3472) );
  INV_X1 U10859 ( .A(n9768), .ZN(n9773) );
  OAI22_X1 U10860 ( .A1(n9770), .A2(n9801), .B1(n9769), .B2(n9799), .ZN(n9772)
         );
  AOI211_X1 U10861 ( .C1(n9787), .C2(n9773), .A(n9772), .B(n9771), .ZN(n9824)
         );
  INV_X1 U10862 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9774) );
  AOI22_X1 U10863 ( .A1(n9809), .A2(n9824), .B1(n9774), .B2(n9807), .ZN(
        P2_U3475) );
  INV_X1 U10864 ( .A(n9775), .ZN(n9779) );
  OAI22_X1 U10865 ( .A1(n9776), .A2(n9801), .B1(n4427), .B2(n9799), .ZN(n9778)
         );
  AOI211_X1 U10866 ( .C1(n9787), .C2(n9779), .A(n9778), .B(n9777), .ZN(n9825)
         );
  INV_X1 U10867 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9780) );
  AOI22_X1 U10868 ( .A1(n9809), .A2(n9825), .B1(n9780), .B2(n9807), .ZN(
        P2_U3478) );
  INV_X1 U10869 ( .A(n9781), .ZN(n9786) );
  OAI22_X1 U10870 ( .A1(n9783), .A2(n9801), .B1(n9782), .B2(n9799), .ZN(n9785)
         );
  AOI211_X1 U10871 ( .C1(n9787), .C2(n9786), .A(n9785), .B(n9784), .ZN(n9826)
         );
  INV_X1 U10872 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9788) );
  AOI22_X1 U10873 ( .A1(n9809), .A2(n9826), .B1(n9788), .B2(n9807), .ZN(
        P2_U3481) );
  AOI22_X1 U10874 ( .A1(n9792), .A2(n9791), .B1(n9790), .B2(n9789), .ZN(n9793)
         );
  OAI211_X1 U10875 ( .C1(n9796), .C2(n9795), .A(n9794), .B(n9793), .ZN(n9797)
         );
  INV_X1 U10876 ( .A(n9797), .ZN(n9827) );
  INV_X1 U10877 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9798) );
  AOI22_X1 U10878 ( .A1(n9809), .A2(n9827), .B1(n9798), .B2(n9807), .ZN(
        P2_U3484) );
  OAI22_X1 U10879 ( .A1(n9802), .A2(n9801), .B1(n9800), .B2(n9799), .ZN(n9804)
         );
  AOI211_X1 U10880 ( .C1(n9806), .C2(n9805), .A(n9804), .B(n9803), .ZN(n9829)
         );
  INV_X1 U10881 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9808) );
  AOI22_X1 U10882 ( .A1(n9809), .A2(n9829), .B1(n9808), .B2(n9807), .ZN(
        P2_U3487) );
  INV_X1 U10883 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9810) );
  AOI22_X1 U10884 ( .A1(n9830), .A2(n9811), .B1(n9810), .B2(n9828), .ZN(
        P2_U3520) );
  AOI22_X1 U10885 ( .A1(n9830), .A2(n9812), .B1(n4512), .B2(n9828), .ZN(
        P2_U3521) );
  AOI22_X1 U10886 ( .A1(n9830), .A2(n9813), .B1(n6705), .B2(n9828), .ZN(
        P2_U3522) );
  INV_X1 U10887 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9814) );
  AOI22_X1 U10888 ( .A1(n9830), .A2(n9815), .B1(n9814), .B2(n9828), .ZN(
        P2_U3523) );
  INV_X1 U10889 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9816) );
  AOI22_X1 U10890 ( .A1(n9830), .A2(n9817), .B1(n9816), .B2(n9828), .ZN(
        P2_U3524) );
  INV_X1 U10891 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9818) );
  AOI22_X1 U10892 ( .A1(n9830), .A2(n9819), .B1(n9818), .B2(n9828), .ZN(
        P2_U3525) );
  INV_X1 U10893 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9820) );
  AOI22_X1 U10894 ( .A1(n9830), .A2(n9821), .B1(n9820), .B2(n9828), .ZN(
        P2_U3526) );
  INV_X1 U10895 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9822) );
  AOI22_X1 U10896 ( .A1(n9830), .A2(n9823), .B1(n9822), .B2(n9828), .ZN(
        P2_U3527) );
  AOI22_X1 U10897 ( .A1(n9830), .A2(n9824), .B1(n6714), .B2(n9828), .ZN(
        P2_U3528) );
  AOI22_X1 U10898 ( .A1(n9830), .A2(n9825), .B1(n4520), .B2(n9828), .ZN(
        P2_U3529) );
  AOI22_X1 U10899 ( .A1(n9830), .A2(n9826), .B1(n6715), .B2(n9828), .ZN(
        P2_U3530) );
  AOI22_X1 U10900 ( .A1(n9830), .A2(n9827), .B1(n6823), .B2(n9828), .ZN(
        P2_U3531) );
  AOI22_X1 U10901 ( .A1(n9830), .A2(n9829), .B1(n6870), .B2(n9828), .ZN(
        P2_U3532) );
  INV_X1 U10902 ( .A(n9831), .ZN(n9832) );
  NAND2_X1 U10903 ( .A1(n9833), .A2(n9832), .ZN(n9834) );
  XOR2_X1 U10904 ( .A(n9835), .B(n9834), .Z(ADD_1071_U5) );
  INV_X1 U10905 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n9836) );
  AOI22_X1 U10906 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n9836), .B2(n9919), .ZN(ADD_1071_U46) );
  OAI21_X1 U10907 ( .B1(n9839), .B2(n9838), .A(n9837), .ZN(ADD_1071_U56) );
  OAI21_X1 U10908 ( .B1(n9842), .B2(n9841), .A(n9840), .ZN(ADD_1071_U57) );
  OAI21_X1 U10909 ( .B1(n9845), .B2(n9844), .A(n9843), .ZN(ADD_1071_U58) );
  OAI21_X1 U10910 ( .B1(n9848), .B2(n9847), .A(n9846), .ZN(ADD_1071_U59) );
  OAI21_X1 U10911 ( .B1(n9851), .B2(n9850), .A(n9849), .ZN(ADD_1071_U60) );
  OAI21_X1 U10912 ( .B1(n9854), .B2(n9853), .A(n9852), .ZN(ADD_1071_U61) );
  AOI21_X1 U10913 ( .B1(n9857), .B2(n9856), .A(n9855), .ZN(ADD_1071_U62) );
  AOI21_X1 U10914 ( .B1(n9860), .B2(n9859), .A(n9858), .ZN(ADD_1071_U63) );
  NAND2_X1 U10915 ( .A1(n9861), .A2(P2_D_REG_31__SCAN_IN), .ZN(n10054) );
  AOI22_X1 U10916 ( .A1(n4520), .A2(keyinput18), .B1(n9863), .B2(keyinput26), 
        .ZN(n9862) );
  OAI221_X1 U10917 ( .B1(n4520), .B2(keyinput18), .C1(n9863), .C2(keyinput26), 
        .A(n9862), .ZN(n9872) );
  INV_X1 U10918 ( .A(SI_14_), .ZN(n9997) );
  AOI22_X1 U10919 ( .A1(n9865), .A2(keyinput20), .B1(n9997), .B2(keyinput50), 
        .ZN(n9864) );
  OAI221_X1 U10920 ( .B1(n9865), .B2(keyinput20), .C1(n9997), .C2(keyinput50), 
        .A(n9864), .ZN(n9871) );
  AOI22_X1 U10921 ( .A1(n9932), .A2(keyinput25), .B1(n9922), .B2(keyinput28), 
        .ZN(n9866) );
  OAI221_X1 U10922 ( .B1(n9932), .B2(keyinput25), .C1(n9922), .C2(keyinput28), 
        .A(n9866), .ZN(n9870) );
  INV_X1 U10923 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9935) );
  XOR2_X1 U10924 ( .A(n9935), .B(keyinput48), .Z(n9868) );
  XNOR2_X1 U10925 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(keyinput34), .ZN(n9867) );
  NAND2_X1 U10926 ( .A1(n9868), .A2(n9867), .ZN(n9869) );
  OR4_X1 U10927 ( .A1(n9872), .A2(n9871), .A3(n9870), .A4(n9869), .ZN(n10052)
         );
  OAI22_X1 U10928 ( .A1(n6235), .A2(keyinput12), .B1(keyinput44), .B2(
        P1_DATAO_REG_20__SCAN_IN), .ZN(n9873) );
  AOI221_X1 U10929 ( .B1(n6235), .B2(keyinput12), .C1(P1_DATAO_REG_20__SCAN_IN), .C2(keyinput44), .A(n9873), .ZN(n9881) );
  OAI22_X1 U10930 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(keyinput62), .B1(
        keyinput59), .B2(P2_REG2_REG_27__SCAN_IN), .ZN(n9874) );
  AOI221_X1 U10931 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(keyinput62), .C1(
        P2_REG2_REG_27__SCAN_IN), .C2(keyinput59), .A(n9874), .ZN(n9880) );
  INV_X1 U10932 ( .A(SI_31_), .ZN(n9926) );
  OAI22_X1 U10933 ( .A1(n9876), .A2(keyinput43), .B1(n9926), .B2(keyinput38), 
        .ZN(n9875) );
  AOI221_X1 U10934 ( .B1(n9876), .B2(keyinput43), .C1(keyinput38), .C2(n9926), 
        .A(n9875), .ZN(n9879) );
  INV_X1 U10935 ( .A(SI_24_), .ZN(n9951) );
  OAI22_X1 U10936 ( .A1(n9960), .A2(keyinput47), .B1(n9951), .B2(keyinput17), 
        .ZN(n9877) );
  AOI221_X1 U10937 ( .B1(n9960), .B2(keyinput47), .C1(keyinput17), .C2(n9951), 
        .A(n9877), .ZN(n9878) );
  NAND4_X1 U10938 ( .A1(n9881), .A2(n9880), .A3(n9879), .A4(n9878), .ZN(n10051) );
  AOI22_X1 U10939 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput46), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(keyinput30), .ZN(n9882) );
  OAI221_X1 U10940 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput46), .C1(
        P1_DATAO_REG_15__SCAN_IN), .C2(keyinput30), .A(n9882), .ZN(n9889) );
  AOI22_X1 U10941 ( .A1(P2_REG2_REG_4__SCAN_IN), .A2(keyinput6), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput4), .ZN(n9883) );
  OAI221_X1 U10942 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(keyinput6), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput4), .A(n9883), .ZN(n9888) );
  AOI22_X1 U10943 ( .A1(P1_REG0_REG_27__SCAN_IN), .A2(keyinput7), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(keyinput29), .ZN(n9884) );
  OAI221_X1 U10944 ( .B1(P1_REG0_REG_27__SCAN_IN), .B2(keyinput7), .C1(
        P2_DATAO_REG_8__SCAN_IN), .C2(keyinput29), .A(n9884), .ZN(n9887) );
  AOI22_X1 U10945 ( .A1(P2_REG1_REG_20__SCAN_IN), .A2(keyinput14), .B1(
        P1_D_REG_0__SCAN_IN), .B2(keyinput49), .ZN(n9885) );
  OAI221_X1 U10946 ( .B1(P2_REG1_REG_20__SCAN_IN), .B2(keyinput14), .C1(
        P1_D_REG_0__SCAN_IN), .C2(keyinput49), .A(n9885), .ZN(n9886) );
  NOR4_X1 U10947 ( .A1(n9889), .A2(n9888), .A3(n9887), .A4(n9886), .ZN(n9917)
         );
  AOI22_X1 U10948 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(keyinput16), .B1(
        P1_D_REG_5__SCAN_IN), .B2(keyinput58), .ZN(n9890) );
  OAI221_X1 U10949 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(keyinput16), .C1(
        P1_D_REG_5__SCAN_IN), .C2(keyinput58), .A(n9890), .ZN(n9897) );
  AOI22_X1 U10950 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(keyinput8), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput39), .ZN(n9891) );
  OAI221_X1 U10951 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(keyinput8), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput39), .A(n9891), .ZN(n9896) );
  AOI22_X1 U10952 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(keyinput35), .B1(
        P1_D_REG_4__SCAN_IN), .B2(keyinput33), .ZN(n9892) );
  OAI221_X1 U10953 ( .B1(P1_REG3_REG_7__SCAN_IN), .B2(keyinput35), .C1(
        P1_D_REG_4__SCAN_IN), .C2(keyinput33), .A(n9892), .ZN(n9895) );
  AOI22_X1 U10954 ( .A1(P1_REG1_REG_1__SCAN_IN), .A2(keyinput45), .B1(
        P1_IR_REG_29__SCAN_IN), .B2(keyinput13), .ZN(n9893) );
  OAI221_X1 U10955 ( .B1(P1_REG1_REG_1__SCAN_IN), .B2(keyinput45), .C1(
        P1_IR_REG_29__SCAN_IN), .C2(keyinput13), .A(n9893), .ZN(n9894) );
  NOR4_X1 U10956 ( .A1(n9897), .A2(n9896), .A3(n9895), .A4(n9894), .ZN(n9916)
         );
  AOI22_X1 U10957 ( .A1(P2_REG0_REG_9__SCAN_IN), .A2(keyinput11), .B1(
        P1_D_REG_19__SCAN_IN), .B2(keyinput31), .ZN(n9898) );
  OAI221_X1 U10958 ( .B1(P2_REG0_REG_9__SCAN_IN), .B2(keyinput11), .C1(
        P1_D_REG_19__SCAN_IN), .C2(keyinput31), .A(n9898), .ZN(n9905) );
  AOI22_X1 U10959 ( .A1(P1_REG0_REG_17__SCAN_IN), .A2(keyinput57), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(keyinput37), .ZN(n9899) );
  OAI221_X1 U10960 ( .B1(P1_REG0_REG_17__SCAN_IN), .B2(keyinput57), .C1(
        P2_DATAO_REG_23__SCAN_IN), .C2(keyinput37), .A(n9899), .ZN(n9904) );
  AOI22_X1 U10961 ( .A1(P2_REG1_REG_25__SCAN_IN), .A2(keyinput54), .B1(SI_28_), 
        .B2(keyinput15), .ZN(n9900) );
  OAI221_X1 U10962 ( .B1(P2_REG1_REG_25__SCAN_IN), .B2(keyinput54), .C1(SI_28_), .C2(keyinput15), .A(n9900), .ZN(n9903) );
  AOI22_X1 U10963 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput40), .B1(
        P1_IR_REG_24__SCAN_IN), .B2(keyinput23), .ZN(n9901) );
  OAI221_X1 U10964 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput40), .C1(
        P1_IR_REG_24__SCAN_IN), .C2(keyinput23), .A(n9901), .ZN(n9902) );
  NOR4_X1 U10965 ( .A1(n9905), .A2(n9904), .A3(n9903), .A4(n9902), .ZN(n9915)
         );
  AOI22_X1 U10966 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(keyinput53), .B1(
        P2_REG2_REG_12__SCAN_IN), .B2(keyinput1), .ZN(n9906) );
  OAI221_X1 U10967 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(keyinput53), .C1(
        P2_REG2_REG_12__SCAN_IN), .C2(keyinput1), .A(n9906), .ZN(n9913) );
  AOI22_X1 U10968 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(keyinput21), .B1(
        P1_REG3_REG_11__SCAN_IN), .B2(keyinput2), .ZN(n9907) );
  OAI221_X1 U10969 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(keyinput21), .C1(
        P1_REG3_REG_11__SCAN_IN), .C2(keyinput2), .A(n9907), .ZN(n9912) );
  AOI22_X1 U10970 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(keyinput55), .B1(
        P2_D_REG_11__SCAN_IN), .B2(keyinput10), .ZN(n9908) );
  OAI221_X1 U10971 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(keyinput55), .C1(
        P2_D_REG_11__SCAN_IN), .C2(keyinput10), .A(n9908), .ZN(n9911) );
  AOI22_X1 U10972 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(keyinput36), .B1(SI_27_), .B2(keyinput22), .ZN(n9909) );
  OAI221_X1 U10973 ( .B1(P1_DATAO_REG_22__SCAN_IN), .B2(keyinput36), .C1(
        SI_27_), .C2(keyinput22), .A(n9909), .ZN(n9910) );
  NOR4_X1 U10974 ( .A1(n9913), .A2(n9912), .A3(n9911), .A4(n9910), .ZN(n9914)
         );
  NAND4_X1 U10975 ( .A1(n9917), .A2(n9916), .A3(n9915), .A4(n9914), .ZN(n10050) );
  AOI22_X1 U10976 ( .A1(n10020), .A2(keyinput67), .B1(keyinput85), .B2(n9919), 
        .ZN(n9918) );
  OAI221_X1 U10977 ( .B1(n10020), .B2(keyinput67), .C1(n9919), .C2(keyinput85), 
        .A(n9918), .ZN(n9930) );
  AOI22_X1 U10978 ( .A1(n9922), .A2(keyinput92), .B1(keyinput94), .B2(n9921), 
        .ZN(n9920) );
  OAI221_X1 U10979 ( .B1(n9922), .B2(keyinput92), .C1(n9921), .C2(keyinput94), 
        .A(n9920), .ZN(n9929) );
  AOI22_X1 U10980 ( .A1(n10017), .A2(keyinput88), .B1(n9924), .B2(keyinput95), 
        .ZN(n9923) );
  OAI221_X1 U10981 ( .B1(n10017), .B2(keyinput88), .C1(n9924), .C2(keyinput95), 
        .A(n9923), .ZN(n9928) );
  AOI22_X1 U10982 ( .A1(n9926), .A2(keyinput102), .B1(n7543), .B2(keyinput79), 
        .ZN(n9925) );
  OAI221_X1 U10983 ( .B1(n9926), .B2(keyinput102), .C1(n7543), .C2(keyinput79), 
        .A(n9925), .ZN(n9927) );
  NOR4_X1 U10984 ( .A1(n9930), .A2(n9929), .A3(n9928), .A4(n9927), .ZN(n9975)
         );
  AOI22_X1 U10985 ( .A1(n9932), .A2(keyinput89), .B1(keyinput66), .B2(n5276), 
        .ZN(n9931) );
  OAI221_X1 U10986 ( .B1(n9932), .B2(keyinput89), .C1(n5276), .C2(keyinput66), 
        .A(n9931), .ZN(n9945) );
  AOI22_X1 U10987 ( .A1(n9935), .A2(keyinput112), .B1(n9934), .B2(keyinput74), 
        .ZN(n9933) );
  OAI221_X1 U10988 ( .B1(n9935), .B2(keyinput112), .C1(n9934), .C2(keyinput74), 
        .A(n9933), .ZN(n9944) );
  AOI22_X1 U10989 ( .A1(n9938), .A2(keyinput103), .B1(keyinput125), .B2(n9937), 
        .ZN(n9936) );
  OAI221_X1 U10990 ( .B1(n9938), .B2(keyinput103), .C1(n9937), .C2(keyinput125), .A(n9936), .ZN(n9943) );
  INV_X1 U10991 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9939) );
  XOR2_X1 U10992 ( .A(n9939), .B(keyinput72), .Z(n9941) );
  XNOR2_X1 U10993 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput105), .ZN(n9940)
         );
  NAND2_X1 U10994 ( .A1(n9941), .A2(n9940), .ZN(n9942) );
  NOR4_X1 U10995 ( .A1(n9945), .A2(n9944), .A3(n9943), .A4(n9942), .ZN(n9974)
         );
  AOI22_X1 U10996 ( .A1(n9948), .A2(keyinput68), .B1(n9947), .B2(keyinput80), 
        .ZN(n9946) );
  OAI221_X1 U10997 ( .B1(n9948), .B2(keyinput68), .C1(n9947), .C2(keyinput80), 
        .A(n9946), .ZN(n9958) );
  INV_X1 U10998 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9950) );
  AOI22_X1 U10999 ( .A1(n9951), .A2(keyinput81), .B1(keyinput78), .B2(n9950), 
        .ZN(n9949) );
  OAI221_X1 U11000 ( .B1(n9951), .B2(keyinput81), .C1(n9950), .C2(keyinput78), 
        .A(n9949), .ZN(n9957) );
  INV_X1 U11001 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10016) );
  AOI22_X1 U11002 ( .A1(n10041), .A2(keyinput120), .B1(keyinput116), .B2(
        n10016), .ZN(n9952) );
  OAI221_X1 U11003 ( .B1(n10041), .B2(keyinput120), .C1(n10016), .C2(
        keyinput116), .A(n9952), .ZN(n9956) );
  AOI22_X1 U11004 ( .A1(n5198), .A2(keyinput99), .B1(keyinput126), .B2(n9954), 
        .ZN(n9953) );
  OAI221_X1 U11005 ( .B1(n5198), .B2(keyinput99), .C1(n9954), .C2(keyinput126), 
        .A(n9953), .ZN(n9955) );
  NOR4_X1 U11006 ( .A1(n9958), .A2(n9957), .A3(n9956), .A4(n9955), .ZN(n9973)
         );
  AOI22_X1 U11007 ( .A1(n10019), .A2(keyinput115), .B1(n9960), .B2(keyinput111), .ZN(n9959) );
  OAI221_X1 U11008 ( .B1(n10019), .B2(keyinput115), .C1(n9960), .C2(
        keyinput111), .A(n9959), .ZN(n9971) );
  INV_X1 U11009 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9962) );
  AOI22_X1 U11010 ( .A1(n9962), .A2(keyinput104), .B1(n6235), .B2(keyinput76), 
        .ZN(n9961) );
  OAI221_X1 U11011 ( .B1(n9962), .B2(keyinput104), .C1(n6235), .C2(keyinput76), 
        .A(n9961), .ZN(n9970) );
  AOI22_X1 U11012 ( .A1(n9965), .A2(keyinput101), .B1(n9964), .B2(keyinput86), 
        .ZN(n9963) );
  OAI221_X1 U11013 ( .B1(n9965), .B2(keyinput101), .C1(n9964), .C2(keyinput86), 
        .A(n9963), .ZN(n9969) );
  XNOR2_X1 U11014 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(keyinput108), .ZN(n9967)
         );
  XNOR2_X1 U11015 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput87), .ZN(n9966) );
  NAND2_X1 U11016 ( .A1(n9967), .A2(n9966), .ZN(n9968) );
  NOR4_X1 U11017 ( .A1(n9971), .A2(n9970), .A3(n9969), .A4(n9968), .ZN(n9972)
         );
  NAND4_X1 U11018 ( .A1(n9975), .A2(n9974), .A3(n9973), .A4(n9972), .ZN(n10048) );
  AOI22_X1 U11019 ( .A1(P2_D_REG_13__SCAN_IN), .A2(keyinput64), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(keyinput124), .ZN(n9976) );
  OAI221_X1 U11020 ( .B1(P2_D_REG_13__SCAN_IN), .B2(keyinput64), .C1(
        P2_DATAO_REG_28__SCAN_IN), .C2(keyinput124), .A(n9976), .ZN(n9983) );
  AOI22_X1 U11021 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(keyinput117), .B1(
        P1_ADDR_REG_4__SCAN_IN), .B2(keyinput84), .ZN(n9977) );
  OAI221_X1 U11022 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(keyinput117), .C1(
        P1_ADDR_REG_4__SCAN_IN), .C2(keyinput84), .A(n9977), .ZN(n9982) );
  AOI22_X1 U11023 ( .A1(P1_REG0_REG_17__SCAN_IN), .A2(keyinput121), .B1(
        P1_IR_REG_29__SCAN_IN), .B2(keyinput77), .ZN(n9978) );
  OAI221_X1 U11024 ( .B1(P1_REG0_REG_17__SCAN_IN), .B2(keyinput121), .C1(
        P1_IR_REG_29__SCAN_IN), .C2(keyinput77), .A(n9978), .ZN(n9981) );
  AOI22_X1 U11025 ( .A1(P2_REG0_REG_9__SCAN_IN), .A2(keyinput75), .B1(
        P1_D_REG_2__SCAN_IN), .B2(keyinput83), .ZN(n9979) );
  OAI221_X1 U11026 ( .B1(P2_REG0_REG_9__SCAN_IN), .B2(keyinput75), .C1(
        P1_D_REG_2__SCAN_IN), .C2(keyinput83), .A(n9979), .ZN(n9980) );
  NOR4_X1 U11027 ( .A1(n9983), .A2(n9982), .A3(n9981), .A4(n9980), .ZN(n10014)
         );
  AOI22_X1 U11028 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(keyinput82), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(keyinput110), .ZN(n9984) );
  OAI221_X1 U11029 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(keyinput82), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput110), .A(n9984), .ZN(n9991) );
  AOI22_X1 U11030 ( .A1(P1_WR_REG_SCAN_IN), .A2(keyinput96), .B1(
        P2_REG1_REG_13__SCAN_IN), .B2(keyinput119), .ZN(n9985) );
  OAI221_X1 U11031 ( .B1(P1_WR_REG_SCAN_IN), .B2(keyinput96), .C1(
        P2_REG1_REG_13__SCAN_IN), .C2(keyinput119), .A(n9985), .ZN(n9990) );
  AOI22_X1 U11032 ( .A1(P1_REG0_REG_27__SCAN_IN), .A2(keyinput71), .B1(
        P1_IR_REG_22__SCAN_IN), .B2(keyinput73), .ZN(n9986) );
  OAI221_X1 U11033 ( .B1(P1_REG0_REG_27__SCAN_IN), .B2(keyinput71), .C1(
        P1_IR_REG_22__SCAN_IN), .C2(keyinput73), .A(n9986), .ZN(n9989) );
  AOI22_X1 U11034 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(keyinput98), .B1(
        P1_D_REG_0__SCAN_IN), .B2(keyinput113), .ZN(n9987) );
  OAI221_X1 U11035 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(keyinput98), .C1(
        P1_D_REG_0__SCAN_IN), .C2(keyinput113), .A(n9987), .ZN(n9988) );
  NOR4_X1 U11036 ( .A1(n9991), .A2(n9990), .A3(n9989), .A4(n9988), .ZN(n10013)
         );
  AOI22_X1 U11037 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput93), .B1(n9993), 
        .B2(keyinput70), .ZN(n9992) );
  OAI221_X1 U11038 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput93), .C1(n9993), 
        .C2(keyinput70), .A(n9992), .ZN(n10002) );
  AOI22_X1 U11039 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(keyinput69), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput106), .ZN(n9994) );
  OAI221_X1 U11040 ( .B1(P1_REG3_REG_18__SCAN_IN), .B2(keyinput69), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput106), .A(n9994), .ZN(n10001) );
  AOI22_X1 U11041 ( .A1(n9997), .A2(keyinput114), .B1(n9996), .B2(keyinput122), 
        .ZN(n9995) );
  OAI221_X1 U11042 ( .B1(n9997), .B2(keyinput114), .C1(n9996), .C2(keyinput122), .A(n9995), .ZN(n10000) );
  AOI22_X1 U11043 ( .A1(n6881), .A2(keyinput65), .B1(n6157), .B2(keyinput123), 
        .ZN(n9998) );
  OAI221_X1 U11044 ( .B1(n6881), .B2(keyinput65), .C1(n6157), .C2(keyinput123), 
        .A(n9998), .ZN(n9999) );
  NOR4_X1 U11045 ( .A1(n10002), .A2(n10001), .A3(n10000), .A4(n9999), .ZN(
        n10012) );
  AOI22_X1 U11046 ( .A1(P2_REG2_REG_5__SCAN_IN), .A2(keyinput91), .B1(
        P1_D_REG_4__SCAN_IN), .B2(keyinput97), .ZN(n10003) );
  OAI221_X1 U11047 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(keyinput91), .C1(
        P1_D_REG_4__SCAN_IN), .C2(keyinput97), .A(n10003), .ZN(n10010) );
  AOI22_X1 U11048 ( .A1(P2_REG1_REG_25__SCAN_IN), .A2(keyinput118), .B1(
        P1_D_REG_6__SCAN_IN), .B2(keyinput90), .ZN(n10004) );
  OAI221_X1 U11049 ( .B1(P2_REG1_REG_25__SCAN_IN), .B2(keyinput118), .C1(
        P1_D_REG_6__SCAN_IN), .C2(keyinput90), .A(n10004), .ZN(n10009) );
  AOI22_X1 U11050 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(keyinput127), .B1(
        P1_REG1_REG_1__SCAN_IN), .B2(keyinput109), .ZN(n10005) );
  OAI221_X1 U11051 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(keyinput127), .C1(
        P1_REG1_REG_1__SCAN_IN), .C2(keyinput109), .A(n10005), .ZN(n10008) );
  AOI22_X1 U11052 ( .A1(P2_REG0_REG_24__SCAN_IN), .A2(keyinput107), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(keyinput100), .ZN(n10006) );
  OAI221_X1 U11053 ( .B1(P2_REG0_REG_24__SCAN_IN), .B2(keyinput107), .C1(
        P1_DATAO_REG_22__SCAN_IN), .C2(keyinput100), .A(n10006), .ZN(n10007)
         );
  NOR4_X1 U11054 ( .A1(n10010), .A2(n10009), .A3(n10008), .A4(n10007), .ZN(
        n10011) );
  NAND4_X1 U11055 ( .A1(n10014), .A2(n10013), .A3(n10012), .A4(n10011), .ZN(
        n10047) );
  AOI22_X1 U11056 ( .A1(n10017), .A2(keyinput24), .B1(keyinput52), .B2(n10016), 
        .ZN(n10015) );
  OAI221_X1 U11057 ( .B1(n10017), .B2(keyinput24), .C1(n10016), .C2(keyinput52), .A(n10015), .ZN(n10028) );
  AOI22_X1 U11058 ( .A1(n10020), .A2(keyinput3), .B1(keyinput51), .B2(n10019), 
        .ZN(n10018) );
  OAI221_X1 U11059 ( .B1(n10020), .B2(keyinput3), .C1(n10019), .C2(keyinput51), 
        .A(n10018), .ZN(n10027) );
  XNOR2_X1 U11060 ( .A(n10021), .B(keyinput32), .ZN(n10026) );
  XNOR2_X1 U11061 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput42), .ZN(n10024) );
  XNOR2_X1 U11062 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput9), .ZN(n10023) );
  XNOR2_X1 U11063 ( .A(P1_REG1_REG_30__SCAN_IN), .B(keyinput61), .ZN(n10022)
         );
  NAND3_X1 U11064 ( .A1(n10024), .A2(n10023), .A3(n10022), .ZN(n10025) );
  NOR4_X1 U11065 ( .A1(n10028), .A2(n10027), .A3(n10026), .A4(n10025), .ZN(
        n10046) );
  AOI22_X1 U11066 ( .A1(n6733), .A2(keyinput27), .B1(n10030), .B2(keyinput5), 
        .ZN(n10029) );
  OAI221_X1 U11067 ( .B1(n6733), .B2(keyinput27), .C1(n10030), .C2(keyinput5), 
        .A(n10029), .ZN(n10035) );
  XNOR2_X1 U11068 ( .A(n10031), .B(keyinput19), .ZN(n10034) );
  XNOR2_X1 U11069 ( .A(n10032), .B(keyinput41), .ZN(n10033) );
  OR3_X1 U11070 ( .A1(n10035), .A2(n10034), .A3(n10033), .ZN(n10044) );
  AOI22_X1 U11071 ( .A1(n10038), .A2(keyinput0), .B1(keyinput63), .B2(n10037), 
        .ZN(n10036) );
  OAI221_X1 U11072 ( .B1(n10038), .B2(keyinput0), .C1(n10037), .C2(keyinput63), 
        .A(n10036), .ZN(n10043) );
  AOI22_X1 U11073 ( .A1(n10041), .A2(keyinput56), .B1(n10040), .B2(keyinput60), 
        .ZN(n10039) );
  OAI221_X1 U11074 ( .B1(n10041), .B2(keyinput56), .C1(n10040), .C2(keyinput60), .A(n10039), .ZN(n10042) );
  NOR3_X1 U11075 ( .A1(n10044), .A2(n10043), .A3(n10042), .ZN(n10045) );
  OAI211_X1 U11076 ( .C1(n10048), .C2(n10047), .A(n10046), .B(n10045), .ZN(
        n10049) );
  NOR4_X1 U11077 ( .A1(n10052), .A2(n10051), .A3(n10050), .A4(n10049), .ZN(
        n10053) );
  XNOR2_X1 U11078 ( .A(n10054), .B(n10053), .ZN(P2_U3297) );
  XOR2_X1 U11079 ( .A(n10055), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11080 ( .A1(n10057), .A2(n10056), .ZN(n10058) );
  XOR2_X1 U11081 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10058), .Z(ADD_1071_U51) );
  XOR2_X1 U11082 ( .A(n10059), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  OAI21_X1 U11083 ( .B1(n10062), .B2(n10061), .A(n10060), .ZN(n10063) );
  XNOR2_X1 U11084 ( .A(n10063), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11085 ( .A(n10064), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  AOI21_X1 U11086 ( .B1(n10067), .B2(n10066), .A(n10065), .ZN(ADD_1071_U47) );
  XOR2_X1 U11087 ( .A(n10069), .B(n10068), .Z(ADD_1071_U54) );
  XOR2_X1 U11088 ( .A(n10071), .B(n10070), .Z(ADD_1071_U53) );
  XNOR2_X1 U11089 ( .A(n10073), .B(n10072), .ZN(ADD_1071_U52) );
  NAND2_X1 U4822 ( .A1(n6700), .A2(n7548), .ZN(n5793) );
  CLKBUF_X1 U6062 ( .A(n6436), .Z(n4297) );
endmodule

