

module b22_C_AntiSAT_k_128_5 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6472, n6473, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15413;

  INV_X4 U7220 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X4 U7221 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  AND2_X1 U7222 ( .A1(n13379), .A2(n13446), .ZN(n13445) );
  NAND3_X1 U7223 ( .A1(n7621), .A2(n7434), .A3(n7622), .ZN(n7623) );
  INV_X2 U7224 ( .A(n11080), .ZN(n11674) );
  AND2_X1 U7225 ( .A1(n12555), .A2(n12551), .ZN(n15072) );
  AND2_X2 U7226 ( .A1(n12524), .A2(n12695), .ZN(n12657) );
  NAND4_X2 U7227 ( .A1(n7780), .A2(n7779), .A3(n7778), .A4(n7777), .ZN(n13309)
         );
  INV_X1 U7228 ( .A(n7736), .ZN(n9210) );
  INV_X2 U7229 ( .A(n9207), .ZN(n8016) );
  NAND2_X1 U7230 ( .A1(n8309), .A2(n9945), .ZN(n8552) );
  CLKBUF_X1 U7231 ( .A(n9387), .Z(n9814) );
  MUX2_X1 U7232 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8803), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8807) );
  INV_X1 U7233 ( .A(n8248), .ZN(n7701) );
  AND3_X2 U7234 ( .A1(n9344), .A2(n9343), .A3(n9342), .ZN(n11339) );
  AOI21_X1 U7235 ( .B1(n7708), .B2(n7707), .A(n7572), .ZN(n7742) );
  NAND2_X2 U7237 ( .A1(n14456), .A2(n14459), .ZN(n9339) );
  NOR2_X1 U7238 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n6713) );
  NOR2_X1 U7239 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6712) );
  INV_X1 U7241 ( .A(n9821), .ZN(n9802) );
  NAND2_X1 U7242 ( .A1(n11651), .A2(n8915), .ZN(n8917) );
  NAND2_X1 U7243 ( .A1(n7051), .A2(n8610), .ZN(n8622) );
  OR2_X1 U7244 ( .A1(n7265), .A2(n6530), .ZN(n7262) );
  AND2_X1 U7245 ( .A1(n8221), .A2(n6863), .ZN(n8993) );
  OR2_X1 U7246 ( .A1(n12455), .A2(n6928), .ZN(n6924) );
  INV_X1 U7247 ( .A(n8956), .ZN(n10646) );
  NAND2_X1 U7248 ( .A1(n12662), .A2(n12663), .ZN(n12902) );
  INV_X1 U7249 ( .A(n10901), .ZN(n8324) );
  INV_X1 U7250 ( .A(n12265), .ZN(n9299) );
  INV_X1 U7251 ( .A(n11339), .ZN(n10982) );
  NAND2_X1 U7252 ( .A1(n8785), .A2(n12599), .ZN(n12130) );
  INV_X1 U7253 ( .A(n7702), .ZN(n8246) );
  INV_X1 U7254 ( .A(n14040), .ZN(n10810) );
  INV_X1 U7255 ( .A(n9387), .ZN(n9791) );
  NAND2_X1 U7256 ( .A1(n12550), .A2(n12553), .ZN(n12547) );
  NAND2_X1 U7257 ( .A1(n8711), .A2(n8710), .ZN(n12464) );
  NAND2_X1 U7258 ( .A1(n7966), .A2(n7965), .ZN(n13744) );
  NAND2_X1 U7259 ( .A1(n9717), .A2(n9716), .ZN(n14351) );
  NAND2_X1 U7260 ( .A1(n9629), .A2(n9628), .ZN(n14385) );
  AND4_X1 U7261 ( .A1(n9392), .A2(n9391), .A3(n9390), .A4(n9389), .ZN(n11194)
         );
  NAND2_X1 U7262 ( .A1(n14448), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9294) );
  NAND4_X1 U7263 ( .A1(n8330), .A2(n8329), .A3(n8328), .A4(n8327), .ZN(n15074)
         );
  OAI21_X1 U7264 ( .B1(n11503), .B2(n7365), .A(n7362), .ZN(n11812) );
  NAND4_X1 U7265 ( .A1(n9429), .A2(n9428), .A3(n9427), .A4(n9426), .ZN(n14034)
         );
  OAI211_X1 U7266 ( .C1(n9207), .C2(n9956), .A(n7746), .B(n7745), .ZN(n10915)
         );
  OAI21_X2 U7267 ( .B1(n13100), .B2(n7402), .A(n7399), .ZN(n12977) );
  CLKBUF_X1 U7268 ( .A(n9177), .Z(n6472) );
  INV_X1 U7269 ( .A(n8996), .ZN(n9177) );
  NAND2_X1 U7270 ( .A1(n9299), .A2(n14453), .ZN(n9812) );
  CLKBUF_X3 U7271 ( .A(n9812), .Z(n6475) );
  NAND2_X2 U7272 ( .A1(n8807), .A2(n8808), .ZN(n11607) );
  INV_X1 U7273 ( .A(n13684), .ZN(n13512) );
  INV_X1 U7274 ( .A(n11981), .ZN(n10537) );
  AOI21_X2 U7275 ( .B1(n7087), .B2(n7084), .A(n6586), .ZN(n7083) );
  OAI21_X2 U7276 ( .B1(n14290), .B2(n6819), .A(n6645), .ZN(n14254) );
  OAI21_X2 U7277 ( .B1(n9887), .B2(n9886), .A(n9885), .ZN(n9898) );
  INV_X4 U7278 ( .A(n8671), .ZN(n12489) );
  XNOR2_X2 U7279 ( .A(n7573), .B(SI_2_), .ZN(n7741) );
  NOR4_X2 U7280 ( .A1(n9253), .A2(n9252), .A3(n7267), .A4(n9251), .ZN(n9255)
         );
  XNOR2_X2 U7281 ( .A(n8308), .B(P3_IR_REG_2__SCAN_IN), .ZN(n10259) );
  OAI21_X2 U7282 ( .B1(n7256), .B2(n6525), .A(n6708), .ZN(n13593) );
  NAND2_X2 U7283 ( .A1(n12214), .A2(n7257), .ZN(n7256) );
  BUF_X4 U7284 ( .A(n8534), .Z(n8765) );
  OAI211_X2 U7285 ( .C1(n10586), .C2(n6532), .A(n6766), .B(n10657), .ZN(n10669) );
  OR2_X1 U7286 ( .A1(n7782), .A2(n6532), .ZN(n6766) );
  NAND2_X2 U7287 ( .A1(n10446), .A2(n7360), .ZN(n10586) );
  BUF_X4 U7288 ( .A(n7753), .Z(n9209) );
  INV_X2 U7289 ( .A(n12657), .ZN(n12675) );
  XNOR2_X1 U7290 ( .A(n13688), .B(n13412), .ZN(n13517) );
  OAI222_X1 U7292 ( .A1(n13178), .A2(n13177), .B1(P3_U3151), .B2(n13176), .C1(
        n13175), .C2(n13174), .ZN(P3_U3266) );
  NAND2_X1 U7293 ( .A1(n8275), .A2(n13176), .ZN(n8298) );
  NAND2_X2 U7294 ( .A1(n12532), .A2(n8883), .ZN(n15111) );
  XNOR2_X2 U7295 ( .A(n8506), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8505) );
  OAI222_X1 U7296 ( .A1(n14464), .A2(n12280), .B1(P1_U3086), .B2(n12265), .C1(
        n12482), .C2(n14474), .ZN(P1_U3325) );
  XNOR2_X2 U7298 ( .A(n7234), .B(n10626), .ZN(n10434) );
  NAND2_X1 U7299 ( .A1(n7050), .A2(n12488), .ZN(n13117) );
  NAND2_X1 U7300 ( .A1(n6716), .A2(n6715), .ZN(n12950) );
  XNOR2_X1 U7301 ( .A(n9206), .B(n9205), .ZN(n12264) );
  NAND2_X1 U7302 ( .A1(n8180), .A2(n8179), .ZN(n13668) );
  NOR2_X2 U7303 ( .A1(n14182), .A2(n14351), .ZN(n7012) );
  INV_X1 U7304 ( .A(n14231), .ZN(n14437) );
  XNOR2_X1 U7305 ( .A(n8093), .B(n8092), .ZN(n8091) );
  NAND2_X1 U7306 ( .A1(n6860), .A2(SI_18_), .ZN(n7433) );
  OR2_X1 U7307 ( .A1(n11395), .A2(n11554), .ZN(n11522) );
  NAND2_X2 U7308 ( .A1(n8324), .A2(n15096), .ZN(n12542) );
  INV_X1 U7309 ( .A(n11119), .ZN(n14306) );
  INV_X1 U7310 ( .A(n14984), .ZN(n6696) );
  INV_X1 U7311 ( .A(n12711), .ZN(n11092) );
  NAND3_X1 U7313 ( .A1(n8315), .A2(n6876), .A3(n8314), .ZN(n12712) );
  NAND2_X1 U7314 ( .A1(n10521), .A2(n8887), .ZN(n8883) );
  INV_X1 U7315 ( .A(n15074), .ZN(n10909) );
  NOR2_X2 U7316 ( .A1(n15108), .A2(n10698), .ZN(n15105) );
  NAND2_X2 U7317 ( .A1(n11141), .A2(n13902), .ZN(n10801) );
  INV_X1 U7318 ( .A(n11053), .ZN(n14802) );
  INV_X2 U7319 ( .A(n7233), .ZN(n10626) );
  CLKBUF_X3 U7320 ( .A(n9338), .Z(n9825) );
  NAND4_X2 U7321 ( .A1(n7706), .A2(n7705), .A3(n7704), .A4(n7703), .ZN(n9002)
         );
  INV_X4 U7322 ( .A(n13938), .ZN(n11103) );
  OR2_X1 U7323 ( .A1(n8298), .A2(n10227), .ZN(n8290) );
  NAND2_X2 U7324 ( .A1(n7728), .A2(n7672), .ZN(n8247) );
  NAND2_X2 U7325 ( .A1(n9339), .A2(n9945), .ZN(n9633) );
  NAND2_X1 U7326 ( .A1(n9339), .A2(n9975), .ZN(n9572) );
  INV_X2 U7327 ( .A(n9339), .ZN(n9627) );
  INV_X2 U7328 ( .A(n7720), .ZN(n7728) );
  INV_X1 U7329 ( .A(n14453), .ZN(n9298) );
  INV_X1 U7330 ( .A(n11983), .ZN(n8221) );
  NAND2_X1 U7331 ( .A1(n8309), .A2(n9975), .ZN(n8412) );
  CLKBUF_X3 U7332 ( .A(n8309), .Z(n10243) );
  INV_X2 U7333 ( .A(n12846), .ZN(n12824) );
  XNOR2_X1 U7334 ( .A(n7586), .B(SI_5_), .ZN(n7786) );
  NAND2_X2 U7335 ( .A1(n8244), .A2(n13796), .ZN(n10069) );
  INV_X1 U7336 ( .A(n9924), .ZN(n6863) );
  OAI21_X1 U7337 ( .B1(n9945), .B2(n9952), .A(n6859), .ZN(n7586) );
  AND2_X1 U7339 ( .A1(n6889), .A2(n6888), .ZN(n12698) );
  AOI21_X1 U7340 ( .B1(n12689), .B2(n8879), .A(n6890), .ZN(n6889) );
  OAI21_X1 U7341 ( .B1(n12497), .B2(n7378), .A(n7377), .ZN(n7376) );
  NAND2_X1 U7342 ( .A1(n9273), .A2(n9274), .ZN(n9272) );
  XNOR2_X1 U7343 ( .A(n6717), .B(n6801), .ZN(n6800) );
  NAND2_X1 U7344 ( .A1(n13901), .A2(n13900), .ZN(n14005) );
  OR2_X1 U7345 ( .A1(n12893), .A2(n8793), .ZN(n8794) );
  OR2_X1 U7346 ( .A1(n12893), .A2(n12892), .ZN(n13058) );
  NAND2_X1 U7347 ( .A1(n12481), .A2(n12480), .ZN(n13122) );
  MUX2_X1 U7348 ( .A(n14422), .B(n14421), .S(n14845), .Z(n14423) );
  OR3_X1 U7349 ( .A1(n13681), .A2(n13680), .A3(n13679), .ZN(n13758) );
  XNOR2_X1 U7350 ( .A(n6875), .B(n6874), .ZN(n13662) );
  NAND2_X1 U7351 ( .A1(n13463), .A2(n13417), .ZN(n6875) );
  AOI21_X1 U7352 ( .B1(n7197), .B2(n7199), .A(n6632), .ZN(n7195) );
  AOI21_X1 U7353 ( .B1(n12328), .B2(n14255), .A(n12327), .ZN(n14335) );
  NAND2_X1 U7354 ( .A1(n6849), .A2(n14125), .ZN(n14341) );
  XNOR2_X1 U7355 ( .A(n12667), .B(n12905), .ZN(n12890) );
  AND2_X1 U7356 ( .A1(n14339), .A2(n14113), .ZN(n7201) );
  OR2_X1 U7357 ( .A1(n14126), .A2(n14831), .ZN(n6849) );
  NAND2_X1 U7358 ( .A1(n12950), .A2(n7218), .ZN(n12932) );
  AND2_X1 U7359 ( .A1(n6774), .A2(n6775), .ZN(n14105) );
  NAND2_X1 U7360 ( .A1(n6774), .A2(n6773), .ZN(n14104) );
  XNOR2_X1 U7361 ( .A(n8090), .B(n8082), .ZN(n13190) );
  NAND2_X1 U7362 ( .A1(n8741), .A2(n8740), .ZN(n8843) );
  NAND2_X1 U7363 ( .A1(n14141), .A2(n14140), .ZN(n14139) );
  INV_X1 U7364 ( .A(n9851), .ZN(n14417) );
  NAND2_X1 U7365 ( .A1(n8693), .A2(n8692), .ZN(n13066) );
  INV_X1 U7366 ( .A(n13439), .ZN(n6874) );
  NAND2_X1 U7367 ( .A1(n14160), .A2(n12318), .ZN(n14138) );
  AOI21_X2 U7368 ( .B1(n12264), .B2(n9209), .A(n9208), .ZN(n13754) );
  NAND2_X1 U7369 ( .A1(n7550), .A2(n12337), .ZN(n6657) );
  AOI21_X1 U7370 ( .B1(n14175), .B2(n14176), .A(n12317), .ZN(n14161) );
  OAI21_X1 U7371 ( .B1(n14208), .B2(n6772), .A(n6770), .ZN(n14175) );
  OAI21_X1 U7372 ( .B1(n12972), .B2(n12515), .A(n12514), .ZN(n12960) );
  NAND2_X1 U7373 ( .A1(n8665), .A2(n8664), .ZN(n12952) );
  NAND2_X1 U7374 ( .A1(n13433), .A2(n13432), .ZN(n13539) );
  NAND2_X1 U7375 ( .A1(n9781), .A2(n9780), .ZN(n14330) );
  NAND2_X1 U7376 ( .A1(n6794), .A2(n8113), .ZN(n13684) );
  AND2_X1 U7377 ( .A1(n13517), .A2(n6527), .ZN(n7265) );
  AND2_X1 U7378 ( .A1(n8158), .A2(n8157), .ZN(n13416) );
  NAND2_X1 U7379 ( .A1(n14768), .A2(n14770), .ZN(n14774) );
  NAND2_X1 U7380 ( .A1(n9737), .A2(n9736), .ZN(n14346) );
  NAND2_X1 U7381 ( .A1(n14221), .A2(n12314), .ZN(n14208) );
  XNOR2_X1 U7382 ( .A(n8688), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n8687) );
  AND2_X1 U7383 ( .A1(n14241), .A2(n12313), .ZN(n7561) );
  OAI21_X1 U7384 ( .B1(n14254), .B2(n7185), .A(n7183), .ZN(n14205) );
  NAND2_X1 U7385 ( .A1(n14241), .A2(n6486), .ZN(n14221) );
  NAND2_X1 U7386 ( .A1(n13034), .A2(n13033), .ZN(n13032) );
  AOI21_X1 U7387 ( .B1(n7237), .B2(n7239), .A(n13431), .ZN(n7235) );
  CLKBUF_X1 U7388 ( .A(n14254), .Z(n6893) );
  NAND2_X1 U7389 ( .A1(n8135), .A2(n8134), .ZN(n13495) );
  NAND2_X1 U7390 ( .A1(n14256), .A2(n7335), .ZN(n14241) );
  NAND2_X1 U7391 ( .A1(n14257), .A2(n14258), .ZN(n14256) );
  NAND2_X1 U7392 ( .A1(n12254), .A2(n12253), .ZN(n12252) );
  NAND2_X1 U7393 ( .A1(n8025), .A2(n13241), .ZN(n13248) );
  AND2_X1 U7394 ( .A1(n14294), .A2(n6509), .ZN(n14240) );
  NOR2_X1 U7395 ( .A1(n13610), .A2(n7127), .ZN(n7126) );
  AND2_X1 U7396 ( .A1(n8081), .A2(n8080), .ZN(n13536) );
  AND2_X1 U7397 ( .A1(n14225), .A2(n12313), .ZN(n6486) );
  NAND2_X1 U7398 ( .A1(n14392), .A2(n12309), .ZN(n14257) );
  NAND2_X1 U7399 ( .A1(n12211), .A2(n12210), .ZN(n12214) );
  AND2_X1 U7400 ( .A1(n14476), .A2(n6853), .ZN(n14193) );
  NAND2_X1 U7401 ( .A1(n14287), .A2(n12308), .ZN(n14282) );
  NAND2_X1 U7402 ( .A1(n9669), .A2(n9668), .ZN(n14431) );
  NAND2_X1 U7403 ( .A1(n14287), .A2(n6487), .ZN(n14392) );
  NAND2_X1 U7404 ( .A1(n7358), .A2(n11968), .ZN(n13245) );
  NAND2_X1 U7405 ( .A1(n12183), .A2(n12182), .ZN(n12181) );
  AND2_X1 U7406 ( .A1(n7995), .A2(n7359), .ZN(n7358) );
  OAI21_X2 U7407 ( .B1(n8091), .B2(n7405), .A(n8094), .ZN(n8132) );
  NAND2_X1 U7408 ( .A1(n11967), .A2(n7991), .ZN(n11968) );
  NAND2_X1 U7409 ( .A1(n12126), .A2(n8521), .ZN(n12183) );
  NAND2_X2 U7410 ( .A1(n7057), .A2(n8046), .ZN(n13710) );
  XNOR2_X1 U7411 ( .A(n14237), .B(n14259), .ZN(n14247) );
  CLKBUF_X1 U7412 ( .A(n8079), .Z(n9682) );
  NAND2_X1 U7413 ( .A1(n8624), .A2(n8623), .ZN(n8639) );
  NAND2_X1 U7414 ( .A1(n6744), .A2(n6528), .ZN(n6955) );
  NAND2_X1 U7415 ( .A1(n12010), .A2(n12009), .ZN(n12013) );
  NAND2_X1 U7416 ( .A1(n11908), .A2(n11907), .ZN(n12010) );
  XNOR2_X1 U7417 ( .A(n8045), .B(n8055), .ZN(n11900) );
  NAND2_X1 U7418 ( .A1(n12084), .A2(n12095), .ZN(n12137) );
  NAND2_X1 U7419 ( .A1(n14615), .A2(n12083), .ZN(n12084) );
  NAND2_X1 U7420 ( .A1(n14617), .A2(n14616), .ZN(n14615) );
  NAND2_X1 U7421 ( .A1(n7433), .A2(n7432), .ZN(n7070) );
  AND2_X1 U7422 ( .A1(n14270), .A2(n12308), .ZN(n6487) );
  OR2_X1 U7423 ( .A1(n11669), .A2(n11668), .ZN(n11818) );
  NAND2_X1 U7424 ( .A1(n12108), .A2(n12082), .ZN(n14617) );
  NAND2_X1 U7425 ( .A1(n8597), .A2(n8596), .ZN(n8609) );
  NAND2_X1 U7426 ( .A1(n8782), .A2(n12584), .ZN(n14667) );
  NAND2_X1 U7427 ( .A1(n11519), .A2(n11660), .ZN(n11667) );
  NAND2_X1 U7428 ( .A1(n9590), .A2(n9589), .ZN(n13828) );
  NAND2_X1 U7429 ( .A1(n11518), .A2(n11517), .ZN(n11519) );
  NAND2_X1 U7430 ( .A1(n11631), .A2(n11630), .ZN(n11632) );
  NAND2_X1 U7431 ( .A1(n7019), .A2(n8564), .ZN(n8579) );
  NAND2_X1 U7432 ( .A1(n7924), .A2(n7923), .ZN(n13221) );
  NAND2_X1 U7433 ( .A1(n11594), .A2(n7325), .ZN(n11631) );
  NAND2_X1 U7434 ( .A1(n9546), .A2(n9545), .ZN(n14602) );
  NAND2_X1 U7435 ( .A1(n11373), .A2(n11372), .ZN(n11594) );
  NAND2_X1 U7436 ( .A1(n7942), .A2(n7941), .ZN(n14868) );
  NAND2_X1 U7437 ( .A1(n11538), .A2(n11371), .ZN(n11373) );
  XNOR2_X1 U7438 ( .A(n7903), .B(n7902), .ZN(n10375) );
  AOI21_X1 U7439 ( .B1(n6477), .B2(n11369), .A(n11368), .ZN(n11540) );
  NAND2_X1 U7440 ( .A1(n9470), .A2(n9469), .ZN(n15198) );
  NAND2_X1 U7441 ( .A1(n7330), .A2(n7331), .ZN(n6477) );
  OR2_X1 U7442 ( .A1(n8507), .A2(n7023), .ZN(n6887) );
  AND2_X1 U7443 ( .A1(n11162), .A2(n11166), .ZN(n11254) );
  INV_X2 U7444 ( .A(n14964), .ZN(n14952) );
  AND2_X2 U7445 ( .A1(n9934), .A2(n14950), .ZN(n14964) );
  INV_X2 U7446 ( .A(n15122), .ZN(n15124) );
  NAND2_X1 U7447 ( .A1(n7106), .A2(n7105), .ZN(n11079) );
  NOR2_X1 U7448 ( .A1(n14015), .A2(n14274), .ZN(n14703) );
  CLKBUF_X3 U7449 ( .A(n8893), .Z(n8957) );
  INV_X2 U7450 ( .A(n8893), .ZN(n8956) );
  AND2_X1 U7451 ( .A1(n6478), .A2(n9858), .ZN(n10851) );
  AOI21_X1 U7452 ( .B1(n10849), .B2(n10850), .A(n9365), .ZN(n10852) );
  NOR2_X1 U7453 ( .A1(n10072), .A2(P2_U3088), .ZN(P2_U3947) );
  INV_X1 U7454 ( .A(n8878), .ZN(n13166) );
  OR2_X1 U7455 ( .A1(n10392), .A2(n10391), .ZN(n6730) );
  INV_X1 U7456 ( .A(n14038), .ZN(n10724) );
  OR2_X1 U7457 ( .A1(n10868), .A2(n10915), .ZN(n10926) );
  INV_X2 U7458 ( .A(n10521), .ZN(n10730) );
  NAND3_X2 U7459 ( .A1(n9337), .A2(n9336), .A3(n9335), .ZN(n14038) );
  AND4_X1 U7460 ( .A1(n8279), .A2(n8277), .A3(n8280), .A4(n8278), .ZN(n10521)
         );
  NAND2_X1 U7461 ( .A1(n10626), .A2(n8994), .ZN(n10868) );
  OAI211_X1 U7462 ( .C1(n8412), .C2(n10012), .A(n8288), .B(n8287), .ZN(n8887)
         );
  AND4_X2 U7463 ( .A1(n9348), .A2(n9346), .A3(n9347), .A4(n6776), .ZN(n11054)
         );
  NAND2_X1 U7464 ( .A1(n9331), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9336) );
  AND2_X1 U7465 ( .A1(n9334), .A2(n9333), .ZN(n9335) );
  INV_X1 U7466 ( .A(n9572), .ZN(n9338) );
  CLKBUF_X1 U7467 ( .A(n8298), .Z(n12493) );
  INV_X2 U7468 ( .A(n8298), .ZN(n8747) );
  INV_X2 U7469 ( .A(n9409), .ZN(n6476) );
  OR2_X1 U7470 ( .A1(n9812), .A2(n9349), .ZN(n6776) );
  MUX2_X1 U7472 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8809), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8810) );
  NAND2_X1 U7473 ( .A1(n10069), .A2(n9945), .ZN(n7962) );
  AND2_X1 U7474 ( .A1(n9923), .A2(n11983), .ZN(n8236) );
  NAND2_X2 U7475 ( .A1(n7672), .A2(n7720), .ZN(n8248) );
  NOR2_X1 U7476 ( .A1(n10261), .A2(n10260), .ZN(n10262) );
  AND2_X2 U7477 ( .A1(n12279), .A2(n7720), .ZN(n7702) );
  INV_X1 U7478 ( .A(n7672), .ZN(n12279) );
  NAND2_X1 U7479 ( .A1(n11977), .A2(n8771), .ZN(n8309) );
  NAND2_X2 U7480 ( .A1(n7336), .A2(n7339), .ZN(n14459) );
  NAND2_X1 U7481 ( .A1(n7646), .A2(n8198), .ZN(n11983) );
  CLKBUF_X1 U7482 ( .A(n11977), .Z(n6870) );
  OAI211_X2 U7483 ( .C1(n9329), .C2(n9328), .A(n9327), .B(n9326), .ZN(n14626)
         );
  XNOR2_X1 U7484 ( .A(n8754), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12695) );
  NAND2_X1 U7485 ( .A1(n8762), .A2(n6514), .ZN(n12529) );
  NAND2_X1 U7486 ( .A1(n6825), .A2(n8318), .ZN(n8333) );
  XNOR2_X1 U7487 ( .A(n9315), .B(n9314), .ZN(n11981) );
  MUX2_X1 U7488 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7645), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n7646) );
  NAND2_X1 U7489 ( .A1(n8198), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6765) );
  NAND2_X1 U7490 ( .A1(n6668), .A2(n6667), .ZN(n13796) );
  AOI21_X1 U7491 ( .B1(n8284), .B2(P3_IR_REG_31__SCAN_IN), .A(n8274), .ZN(
        n7208) );
  OR2_X1 U7492 ( .A1(n9296), .A2(n7502), .ZN(n6813) );
  NAND2_X1 U7493 ( .A1(n8270), .A2(n7386), .ZN(n13168) );
  NAND2_X2 U7494 ( .A1(n9945), .A2(P1_U3086), .ZN(n14474) );
  MUX2_X1 U7495 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8283), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n6877) );
  NAND2_X1 U7496 ( .A1(n7017), .A2(n7016), .ZN(n7339) );
  NAND2_X1 U7497 ( .A1(n9945), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6859) );
  NAND2_X2 U7498 ( .A1(n9975), .A2(P3_U3151), .ZN(n13175) );
  AOI21_X1 U7499 ( .B1(n8011), .B2(n7665), .A(n6568), .ZN(n7666) );
  NAND2_X1 U7500 ( .A1(n6584), .A2(n9311), .ZN(n14448) );
  NOR2_X1 U7501 ( .A1(n8508), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8527) );
  AND2_X1 U7502 ( .A1(n6704), .A2(n7639), .ZN(n7558) );
  NOR2_X1 U7503 ( .A1(n8268), .A2(P3_IR_REG_26__SCAN_IN), .ZN(n7384) );
  AND2_X1 U7504 ( .A1(n8755), .A2(n8266), .ZN(n7557) );
  NOR2_X2 U7505 ( .A1(n9393), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9431) );
  AND2_X1 U7506 ( .A1(n7649), .A2(n7647), .ZN(n7656) );
  AND4_X1 U7507 ( .A1(n7637), .A2(n7633), .A3(n7767), .A4(n7804), .ZN(n6706)
         );
  AND3_X1 U7508 ( .A1(n8265), .A2(n8264), .A3(n8263), .ZN(n8755) );
  NAND2_X1 U7509 ( .A1(n8285), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8303) );
  AND2_X1 U7510 ( .A1(n6653), .A2(n6652), .ZN(n9893) );
  AND2_X1 U7511 ( .A1(n7636), .A2(n7634), .ZN(n6705) );
  INV_X1 U7512 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9451) );
  INV_X1 U7513 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7767) );
  INV_X1 U7514 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n7655) );
  NOR2_X1 U7515 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n7371) );
  NOR2_X1 U7516 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7743) );
  INV_X1 U7517 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8833) );
  INV_X1 U7518 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8285) );
  INV_X1 U7519 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7369) );
  INV_X1 U7520 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8199) );
  NOR2_X1 U7521 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n10246) );
  NOR2_X1 U7522 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), .ZN(
        n8267) );
  INV_X1 U7523 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7327) );
  INV_X1 U7524 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9430) );
  INV_X1 U7525 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8805) );
  NOR2_X1 U7526 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n7634) );
  NOR2_X1 U7527 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n7637) );
  INV_X4 U7528 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7529 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6479) );
  INV_X1 U7530 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9432) );
  INV_X1 U7531 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n6480) );
  INV_X1 U7532 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6481) );
  NOR2_X1 U7533 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n7370) );
  NOR2_X1 U7534 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n8263) );
  NOR2_X1 U7535 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n8264) );
  NOR2_X1 U7536 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n8265) );
  INV_X1 U7537 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9562) );
  NOR2_X1 U7538 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n6484) );
  NOR2_X1 U7539 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6483) );
  INV_X1 U7540 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7063) );
  INV_X1 U7541 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n12003) );
  INV_X1 U7542 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7062) );
  INV_X1 U7543 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7568) );
  XNOR2_X1 U7544 ( .A(n6477), .B(n11374), .ZN(n11428) );
  NAND2_X1 U7545 ( .A1(n10988), .A2(n6478), .ZN(n10990) );
  NAND2_X1 U7546 ( .A1(n10724), .A2(n10982), .ZN(n6478) );
  AND3_X4 U7547 ( .A1(n9305), .A2(n7556), .A3(n9431), .ZN(n9311) );
  NAND4_X2 U7548 ( .A1(n7327), .A2(n6481), .A3(n6480), .A4(n6479), .ZN(n9393)
         );
  NOR2_X2 U7549 ( .A1(n9586), .A2(n6482), .ZN(n9305) );
  NAND4_X1 U7550 ( .A1(n9286), .A2(n9432), .A3(n9430), .A4(n9451), .ZN(n6482)
         );
  NAND4_X1 U7551 ( .A1(n6485), .A2(n6484), .A3(n6483), .A4(n9562), .ZN(n9586)
         );
  NOR2_X1 U7552 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n6485) );
  NAND2_X1 U7553 ( .A1(n12306), .A2(n7334), .ZN(n14287) );
  NAND2_X1 U7554 ( .A1(n9304), .A2(n6561), .ZN(n6654) );
  OAI21_X2 U7555 ( .B1(n7465), .B2(n7460), .A(n7458), .ZN(n12466) );
  OAI21_X2 U7556 ( .B1(n8359), .B2(n7213), .A(n7212), .ZN(n11232) );
  INV_X4 U7558 ( .A(n6476), .ZN(n9386) );
  OAI21_X2 U7559 ( .B1(n14667), .B2(n7390), .A(n7387), .ZN(n14650) );
  NAND2_X1 U7560 ( .A1(n10810), .A2(n11053), .ZN(n10850) );
  NAND4_X2 U7561 ( .A1(n7740), .A2(n7739), .A3(n7738), .A4(n7737), .ZN(n13311)
         );
  NAND2_X4 U7562 ( .A1(n8236), .A2(n6863), .ZN(n11080) );
  OAI211_X1 U7563 ( .C1(n9602), .C2(n12095), .A(n6490), .B(n9604), .ZN(n7512)
         );
  NAND2_X1 U7564 ( .A1(n6583), .A2(n12320), .ZN(n7352) );
  AND2_X1 U7565 ( .A1(n8261), .A2(n8260), .ZN(n8262) );
  NOR2_X1 U7566 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8261) );
  NOR2_X1 U7567 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n8260) );
  NAND2_X1 U7568 ( .A1(n10730), .A2(n15104), .ZN(n12532) );
  AND2_X1 U7569 ( .A1(n6797), .A2(n6537), .ZN(n7087) );
  NAND2_X1 U7570 ( .A1(n12267), .A2(n8123), .ZN(n6797) );
  INV_X1 U7571 ( .A(n7258), .ZN(n7257) );
  OAI21_X1 U7572 ( .B1(n12213), .B2(n7259), .A(n13422), .ZN(n7258) );
  AND2_X1 U7573 ( .A1(n12363), .A2(n9852), .ZN(n12341) );
  NAND2_X1 U7574 ( .A1(n7071), .A2(n7075), .ZN(n7886) );
  NAND2_X1 U7575 ( .A1(n7864), .A2(n7599), .ZN(n7071) );
  XNOR2_X1 U7576 ( .A(n7374), .B(n12859), .ZN(n12691) );
  NAND2_X1 U7577 ( .A1(n7376), .A2(n7375), .ZN(n7374) );
  NOR2_X1 U7578 ( .A1(n12684), .A2(n6535), .ZN(n7375) );
  NAND2_X1 U7579 ( .A1(n12917), .A2(n8704), .ZN(n12903) );
  AOI21_X1 U7580 ( .B1(n7429), .B2(n14127), .A(n7431), .ZN(n7428) );
  NOR2_X1 U7581 ( .A1(n14024), .A2(n14337), .ZN(n7431) );
  NOR2_X1 U7582 ( .A1(n14554), .A2(n14594), .ZN(n14557) );
  AOI21_X1 U7583 ( .B1(n7492), .B2(n7491), .A(n7489), .ZN(n7488) );
  NAND2_X1 U7584 ( .A1(n6689), .A2(n9023), .ZN(n9024) );
  AND2_X1 U7585 ( .A1(n7511), .A2(n12334), .ZN(n7506) );
  OAI21_X1 U7586 ( .B1(n7510), .B2(n7509), .A(n7508), .ZN(n7504) );
  INV_X1 U7587 ( .A(n9618), .ZN(n7508) );
  OAI21_X1 U7588 ( .B1(n6676), .B2(n6675), .A(n6540), .ZN(n7531) );
  AOI21_X1 U7589 ( .B1(n9148), .B2(n9149), .A(n9147), .ZN(n6676) );
  NOR2_X1 U7590 ( .A1(n9148), .A2(n9149), .ZN(n6675) );
  OAI21_X1 U7591 ( .B1(n7419), .B2(n7418), .A(n7920), .ZN(n7417) );
  INV_X1 U7592 ( .A(n6792), .ZN(n14482) );
  NOR2_X1 U7593 ( .A1(n8554), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8569) );
  INV_X1 U7594 ( .A(n13176), .ZN(n8276) );
  NAND2_X1 U7595 ( .A1(n6907), .A2(n15030), .ZN(n6906) );
  NOR2_X1 U7596 ( .A1(n11841), .A2(n7232), .ZN(n11957) );
  AND2_X1 U7597 ( .A1(n11842), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7232) );
  AND3_X1 U7598 ( .A1(n6956), .A2(n6634), .A3(n6958), .ZN(n12744) );
  AND2_X1 U7599 ( .A1(n6953), .A2(n6952), .ZN(n12830) );
  NAND2_X1 U7600 ( .A1(n12802), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n6952) );
  OR2_X1 U7601 ( .A1(n13090), .A2(n12974), .ZN(n12634) );
  OR2_X1 U7602 ( .A1(n8552), .A2(n10011), .ZN(n8288) );
  NAND2_X1 U7603 ( .A1(n8601), .A2(n10416), .ZN(n8287) );
  INV_X1 U7604 ( .A(n12529), .ZN(n12524) );
  XNOR2_X1 U7605 ( .A(n6746), .B(n8281), .ZN(n8771) );
  NAND2_X1 U7606 ( .A1(n6747), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6746) );
  AND2_X1 U7607 ( .A1(n7049), .A2(n8388), .ZN(n7048) );
  INV_X1 U7608 ( .A(n8391), .ZN(n7049) );
  AND2_X1 U7609 ( .A1(n7098), .A2(n7097), .ZN(n7096) );
  NAND2_X1 U7610 ( .A1(n13678), .A2(n13436), .ZN(n7157) );
  NOR2_X1 U7611 ( .A1(n7162), .A2(n7167), .ZN(n7159) );
  NOR2_X1 U7612 ( .A1(n13430), .A2(n7241), .ZN(n7240) );
  INV_X1 U7613 ( .A(n13429), .ZN(n7241) );
  INV_X1 U7614 ( .A(n13420), .ZN(n7259) );
  NAND2_X1 U7615 ( .A1(n9002), .A2(n10626), .ZN(n9237) );
  NAND2_X1 U7616 ( .A1(n9236), .A2(n7233), .ZN(n10860) );
  AND2_X2 U7617 ( .A1(n7743), .A2(n7635), .ZN(n7768) );
  INV_X1 U7618 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7635) );
  NAND2_X1 U7619 ( .A1(n14104), .A2(n12322), .ZN(n12323) );
  OR2_X1 U7620 ( .A1(n14231), .A2(n13956), .ZN(n12314) );
  AND2_X1 U7621 ( .A1(n6646), .A2(n7509), .ZN(n6645) );
  NAND2_X1 U7622 ( .A1(n6647), .A2(n12333), .ZN(n6646) );
  INV_X1 U7623 ( .A(n12332), .ZN(n6647) );
  NAND2_X1 U7624 ( .A1(n9181), .A2(n9180), .ZN(n9202) );
  XNOR2_X1 U7625 ( .A(n8061), .B(SI_20_), .ZN(n8045) );
  NAND2_X1 U7626 ( .A1(n7424), .A2(n7426), .ZN(n7421) );
  NAND2_X1 U7627 ( .A1(n7596), .A2(n7422), .ZN(n6793) );
  OAI21_X1 U7628 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14497), .A(n14496), .ZN(
        n14561) );
  AOI21_X1 U7629 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n14504), .A(n14503), .ZN(
        n14570) );
  NAND2_X1 U7630 ( .A1(n7455), .A2(n6636), .ZN(n7454) );
  OR2_X1 U7631 ( .A1(n8930), .A2(n8931), .ZN(n6940) );
  NAND2_X1 U7632 ( .A1(n10688), .A2(n7474), .ZN(n10814) );
  INV_X1 U7633 ( .A(n7472), .ZN(n7474) );
  INV_X1 U7634 ( .A(n8902), .ZN(n7473) );
  INV_X1 U7635 ( .A(n8313), .ZN(n8750) );
  NOR2_X1 U7636 ( .A1(n10406), .A2(n10225), .ZN(n10405) );
  OR2_X1 U7637 ( .A1(n10470), .A2(n10471), .ZN(n6743) );
  NOR2_X1 U7638 ( .A1(n7294), .A2(n11949), .ZN(n6915) );
  NOR2_X1 U7639 ( .A1(n12727), .A2(n12715), .ZN(n12746) );
  NAND2_X1 U7640 ( .A1(n6951), .A2(n6950), .ZN(n6835) );
  INV_X1 U7641 ( .A(n12748), .ZN(n6950) );
  OR2_X1 U7642 ( .A1(n12767), .A2(n13114), .ZN(n6744) );
  AND2_X1 U7643 ( .A1(n12933), .A2(n8675), .ZN(n7218) );
  AOI21_X1 U7644 ( .B1(n7396), .B2(n7395), .A(n7394), .ZN(n7393) );
  INV_X1 U7645 ( .A(n12613), .ZN(n7394) );
  INV_X1 U7646 ( .A(n12603), .ZN(n7395) );
  AND2_X1 U7647 ( .A1(n12578), .A2(n8432), .ZN(n12571) );
  BUF_X1 U7648 ( .A(n8371), .Z(n12479) );
  INV_X4 U7649 ( .A(n8412), .ZN(n12487) );
  INV_X1 U7650 ( .A(n8552), .ZN(n8371) );
  INV_X1 U7651 ( .A(n8282), .ZN(n8270) );
  AND2_X1 U7652 ( .A1(n6638), .A2(n8725), .ZN(n7052) );
  NAND2_X1 U7653 ( .A1(n8659), .A2(n8658), .ZN(n8662) );
  INV_X1 U7654 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8599) );
  NAND2_X1 U7655 ( .A1(n6949), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8600) );
  INV_X1 U7656 ( .A(n7032), .ZN(n7031) );
  OAI21_X1 U7657 ( .B1(n8440), .B2(n7033), .A(n8444), .ZN(n7032) );
  NAND2_X1 U7658 ( .A1(n6885), .A2(n8440), .ZN(n7030) );
  AND2_X1 U7659 ( .A1(n8415), .A2(n8403), .ZN(n8404) );
  AOI21_X1 U7660 ( .B1(n8367), .B2(n7039), .A(n7038), .ZN(n7037) );
  INV_X1 U7661 ( .A(n8353), .ZN(n7039) );
  OR2_X1 U7662 ( .A1(n8339), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8372) );
  INV_X1 U7663 ( .A(n7087), .ZN(n7085) );
  INV_X1 U7664 ( .A(n8150), .ZN(n7357) );
  NOR2_X1 U7665 ( .A1(n12304), .A2(n8074), .ZN(n8090) );
  NAND2_X1 U7666 ( .A1(n11219), .A2(n6757), .ZN(n11261) );
  NOR2_X1 U7667 ( .A1(n11263), .A2(n6758), .ZN(n6757) );
  INV_X1 U7668 ( .A(n11222), .ZN(n6758) );
  XNOR2_X1 U7669 ( .A(n13710), .B(n6809), .ZN(n8048) );
  NAND2_X1 U7670 ( .A1(n11503), .A2(n7933), .ZN(n13216) );
  NAND2_X1 U7671 ( .A1(n13524), .A2(n13512), .ZN(n13508) );
  INV_X1 U7672 ( .A(n7267), .ZN(n7260) );
  XNOR2_X1 U7673 ( .A(n13684), .B(n13485), .ZN(n7267) );
  OAI21_X1 U7674 ( .B1(n12161), .B2(n7133), .A(n7131), .ZN(n13393) );
  INV_X1 U7675 ( .A(n7134), .ZN(n7133) );
  AOI21_X1 U7676 ( .B1(n7134), .B2(n7132), .A(n12213), .ZN(n7131) );
  INV_X1 U7677 ( .A(n7135), .ZN(n7132) );
  NAND2_X1 U7678 ( .A1(n11818), .A2(n7276), .ZN(n11906) );
  AND2_X1 U7679 ( .A1(n11819), .A2(n11817), .ZN(n7276) );
  AOI21_X1 U7680 ( .B1(n6496), .B2(n7122), .A(n6543), .ZN(n7120) );
  NAND2_X1 U7681 ( .A1(n11403), .A2(n11513), .ZN(n11518) );
  NAND2_X1 U7682 ( .A1(n11246), .A2(n11245), .ZN(n7273) );
  AND2_X1 U7683 ( .A1(n9926), .A2(n9925), .ZN(n13562) );
  AND2_X1 U7684 ( .A1(n9267), .A2(n8236), .ZN(n14990) );
  INV_X1 U7685 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7671) );
  NAND2_X1 U7686 ( .A1(n6712), .A2(n6711), .ZN(n6700) );
  INV_X1 U7687 ( .A(n7340), .ZN(n6998) );
  AOI21_X1 U7688 ( .B1(n6491), .B2(n12228), .A(n7345), .ZN(n7340) );
  AND2_X1 U7689 ( .A1(n13815), .A2(n13816), .ZN(n7345) );
  OAI21_X1 U7690 ( .B1(n11613), .B2(n6968), .A(n6966), .ZN(n15194) );
  AOI21_X1 U7691 ( .B1(n6969), .B2(n6972), .A(n6967), .ZN(n6966) );
  INV_X1 U7692 ( .A(n6969), .ZN(n6968) );
  INV_X1 U7693 ( .A(n15195), .ZN(n6967) );
  NOR2_X1 U7694 ( .A1(n13837), .A2(n13836), .ZN(n13838) );
  NAND2_X1 U7695 ( .A1(n7427), .A2(n6544), .ZN(n12352) );
  NAND2_X1 U7696 ( .A1(n14146), .A2(n12340), .ZN(n14128) );
  NOR2_X1 U7697 ( .A1(n14225), .A2(n7189), .ZN(n7186) );
  OAI21_X1 U7698 ( .B1(n12329), .B2(n12330), .A(n12331), .ZN(n14292) );
  OR2_X1 U7699 ( .A1(n13828), .A2(n14713), .ZN(n12305) );
  AOI21_X1 U7700 ( .B1(n11638), .B2(n11755), .A(n7323), .ZN(n7322) );
  NAND2_X1 U7702 ( .A1(n9820), .A2(n9819), .ZN(n14327) );
  INV_X1 U7703 ( .A(n14837), .ZN(n14828) );
  AND2_X1 U7704 ( .A1(n9893), .A2(n6538), .ZN(n7564) );
  INV_X1 U7705 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9289) );
  INV_X1 U7706 ( .A(n14448), .ZN(n6812) );
  AOI21_X1 U7707 ( .B1(n14597), .B2(n6503), .A(n6575), .ZN(n14562) );
  NAND2_X1 U7708 ( .A1(n14755), .A2(n14559), .ZN(n6785) );
  NOR2_X1 U7709 ( .A1(n12409), .A2(n12410), .ZN(n12408) );
  AOI21_X1 U7710 ( .B1(n12889), .B2(n15109), .A(n8855), .ZN(n8856) );
  NAND2_X1 U7711 ( .A1(n6800), .A2(n15112), .ZN(n8857) );
  NAND2_X1 U7712 ( .A1(n8018), .A2(n8017), .ZN(n13727) );
  NAND2_X1 U7713 ( .A1(n6767), .A2(n10436), .ZN(n10446) );
  NAND2_X1 U7714 ( .A1(n10435), .A2(n7735), .ZN(n6767) );
  NAND2_X1 U7715 ( .A1(n7693), .A2(n7692), .ZN(n13625) );
  NAND2_X1 U7716 ( .A1(n9750), .A2(n9749), .ZN(n14130) );
  MUX2_X1 U7717 ( .A(n10724), .B(n11339), .S(n9399), .Z(n9370) );
  INV_X1 U7718 ( .A(n9456), .ZN(n7493) );
  NAND2_X1 U7719 ( .A1(n6691), .A2(n6690), .ZN(n9021) );
  INV_X1 U7720 ( .A(n9015), .ZN(n6822) );
  OR2_X1 U7721 ( .A1(n7493), .A2(n9458), .ZN(n7491) );
  NAND2_X1 U7722 ( .A1(n9444), .A2(n9443), .ZN(n9457) );
  AND2_X1 U7723 ( .A1(n7493), .A2(n9458), .ZN(n7492) );
  OR2_X1 U7724 ( .A1(n9021), .A2(n9020), .ZN(n7548) );
  INV_X1 U7725 ( .A(n9028), .ZN(n7535) );
  OAI22_X1 U7726 ( .A1(n9046), .A2(n6686), .B1(n9045), .B2(n9044), .ZN(n9052)
         );
  NOR2_X1 U7727 ( .A1(n6882), .A2(n6824), .ZN(n6686) );
  OAI22_X1 U7728 ( .A1(n9039), .A2(n7540), .B1(n7539), .B2(n9040), .ZN(n9046)
         );
  INV_X1 U7729 ( .A(n9045), .ZN(n6824) );
  INV_X1 U7730 ( .A(n9068), .ZN(n6684) );
  AND2_X1 U7731 ( .A1(n7505), .A2(n6612), .ZN(n7510) );
  NAND2_X1 U7732 ( .A1(n7511), .A2(n9602), .ZN(n7505) );
  INV_X1 U7733 ( .A(n9606), .ZN(n7514) );
  NAND2_X1 U7734 ( .A1(n7521), .A2(n7520), .ZN(n7519) );
  INV_X1 U7735 ( .A(n9101), .ZN(n7521) );
  INV_X1 U7736 ( .A(n9102), .ZN(n7520) );
  OAI21_X1 U7737 ( .B1(n6688), .B2(n6687), .A(n7516), .ZN(n9123) );
  OR3_X1 U7738 ( .A1(n9108), .A2(n9107), .A3(n9106), .ZN(n9121) );
  NOR2_X1 U7739 ( .A1(n9660), .A2(n9661), .ZN(n7499) );
  AOI21_X1 U7740 ( .B1(n9660), .B2(n9661), .A(n7500), .ZN(n7494) );
  INV_X1 U7741 ( .A(n9648), .ZN(n7500) );
  NAND2_X1 U7742 ( .A1(n9142), .A2(n9144), .ZN(n7542) );
  INV_X1 U7743 ( .A(n7532), .ZN(n7530) );
  INV_X1 U7744 ( .A(n9153), .ZN(n6880) );
  OR2_X1 U7745 ( .A1(n9157), .A2(n9158), .ZN(n6673) );
  AND2_X1 U7746 ( .A1(n7392), .A2(n14661), .ZN(n7391) );
  NAND2_X1 U7747 ( .A1(n14671), .A2(n12590), .ZN(n7392) );
  INV_X1 U7748 ( .A(n12593), .ZN(n7388) );
  INV_X1 U7749 ( .A(n8522), .ZN(n7023) );
  INV_X1 U7750 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8496) );
  NAND2_X1 U7751 ( .A1(n9169), .A2(n9170), .ZN(n7528) );
  OAI22_X1 U7752 ( .A1(n9179), .A2(n9178), .B1(n9169), .B2(n9170), .ZN(n7526)
         );
  OAI21_X1 U7753 ( .B1(n9164), .B2(n9163), .A(n9162), .ZN(n9165) );
  XNOR2_X1 U7754 ( .A(n9829), .B(n14626), .ZN(n9803) );
  INV_X1 U7755 ( .A(n7350), .ZN(n6775) );
  OAI21_X1 U7756 ( .B1(n14140), .B2(n7352), .A(n12321), .ZN(n7350) );
  NAND2_X1 U7757 ( .A1(n14138), .A2(n7351), .ZN(n6774) );
  INV_X1 U7758 ( .A(n7352), .ZN(n7351) );
  NAND3_X1 U7759 ( .A1(n7065), .A2(n7067), .A3(n7627), .ZN(n8061) );
  NAND2_X1 U7760 ( .A1(n7433), .A2(n7068), .ZN(n7067) );
  NOR2_X1 U7761 ( .A1(n7412), .A2(n7688), .ZN(n7068) );
  NOR2_X1 U7762 ( .A1(n7979), .A2(n7093), .ZN(n7089) );
  INV_X1 U7763 ( .A(n7996), .ZN(n7093) );
  INV_X1 U7764 ( .A(n7618), .ZN(n7091) );
  AOI21_X1 U7765 ( .B1(n7075), .B2(n7073), .A(n7417), .ZN(n7072) );
  INV_X1 U7766 ( .A(n7599), .ZN(n7073) );
  INV_X1 U7767 ( .A(n7075), .ZN(n7074) );
  INV_X1 U7768 ( .A(n7417), .ZN(n7416) );
  INV_X1 U7769 ( .A(n7605), .ZN(n7418) );
  AND2_X1 U7770 ( .A1(n7076), .A2(n7883), .ZN(n7075) );
  NAND2_X1 U7771 ( .A1(n7862), .A2(n7599), .ZN(n7076) );
  INV_X1 U7772 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7064) );
  NAND2_X1 U7773 ( .A1(n7060), .A2(n12003), .ZN(n7407) );
  NAND2_X1 U7774 ( .A1(n6852), .A2(n6570), .ZN(n6851) );
  NAND2_X1 U7775 ( .A1(n14483), .A2(n10779), .ZN(n6852) );
  INV_X1 U7776 ( .A(n6929), .ZN(n6928) );
  NOR2_X1 U7777 ( .A1(n6930), .A2(n12390), .ZN(n6929) );
  INV_X1 U7778 ( .A(n6933), .ZN(n6930) );
  INV_X1 U7779 ( .A(n6935), .ZN(n6927) );
  NAND2_X1 U7780 ( .A1(n8934), .A2(n12963), .ZN(n8935) );
  AND2_X1 U7781 ( .A1(n8569), .A2(n8568), .ZN(n8586) );
  NOR2_X1 U7782 ( .A1(n12522), .A2(n12500), .ZN(n7377) );
  INV_X1 U7783 ( .A(n12676), .ZN(n6843) );
  NAND2_X1 U7784 ( .A1(n12666), .A2(n12890), .ZN(n12674) );
  NAND2_X1 U7785 ( .A1(n10483), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7289) );
  OR2_X1 U7786 ( .A1(n10466), .A2(n10467), .ZN(n6666) );
  INV_X1 U7787 ( .A(n7289), .ZN(n7288) );
  NAND2_X1 U7788 ( .A1(n11021), .A2(n11022), .ZN(n11293) );
  INV_X1 U7789 ( .A(n7282), .ZN(n6908) );
  INV_X1 U7790 ( .A(n12835), .ZN(n7230) );
  AND2_X1 U7791 ( .A1(n6661), .A2(n6660), .ZN(n12813) );
  NAND2_X1 U7792 ( .A1(n12802), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n6660) );
  OR2_X1 U7793 ( .A1(n8840), .A2(n8848), .ZN(n12671) );
  AND2_X1 U7794 ( .A1(n8695), .A2(n8694), .ZN(n8713) );
  NOR2_X1 U7795 ( .A1(n8680), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8695) );
  OR2_X1 U7796 ( .A1(n12966), .A2(n12975), .ZN(n12643) );
  INV_X1 U7797 ( .A(n6807), .ZN(n6805) );
  INV_X1 U7798 ( .A(n8788), .ZN(n7401) );
  NOR2_X1 U7799 ( .A1(n8613), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8628) );
  NOR2_X1 U7800 ( .A1(n7217), .A2(n6808), .ZN(n6807) );
  INV_X1 U7801 ( .A(n8576), .ZN(n6808) );
  NAND2_X1 U7802 ( .A1(n6497), .A2(n13028), .ZN(n7217) );
  OR2_X1 U7803 ( .A1(n13098), .A2(n8931), .ZN(n12622) );
  OR2_X1 U7804 ( .A1(n13158), .A2(n13035), .ZN(n12614) );
  NAND2_X1 U7805 ( .A1(n11208), .A2(n11317), .ZN(n12564) );
  NAND2_X1 U7806 ( .A1(n12542), .A2(n12545), .ZN(n7216) );
  NOR3_X1 U7807 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_20__SCAN_IN), .A3(
        P3_IR_REG_13__SCAN_IN), .ZN(n8266) );
  INV_X1 U7808 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8802) );
  NAND2_X1 U7809 ( .A1(n8500), .A2(n7557), .ZN(n8759) );
  NOR2_X1 U7810 ( .A1(n7023), .A2(n10615), .ZN(n7021) );
  NAND2_X2 U7811 ( .A1(n9920), .A2(n9259), .ZN(n8181) );
  NOR2_X1 U7812 ( .A1(n8198), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n8227) );
  NAND2_X1 U7813 ( .A1(n7100), .A2(n13484), .ZN(n7250) );
  NAND2_X1 U7814 ( .A1(n12165), .A2(n7274), .ZN(n12211) );
  NOR2_X1 U7815 ( .A1(n12200), .A2(n7275), .ZN(n7274) );
  INV_X1 U7816 ( .A(n12164), .ZN(n7275) );
  INV_X1 U7817 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7662) );
  INV_X1 U7818 ( .A(n13910), .ZN(n7318) );
  NAND2_X1 U7819 ( .A1(n11773), .A2(n11774), .ZN(n6975) );
  NAND2_X1 U7820 ( .A1(n14041), .A2(n13902), .ZN(n7348) );
  INV_X1 U7821 ( .A(n7191), .ZN(n7184) );
  NOR2_X1 U7822 ( .A1(n14247), .A2(n7192), .ZN(n7191) );
  INV_X1 U7823 ( .A(n12335), .ZN(n7192) );
  OAI21_X1 U7824 ( .B1(n14247), .B2(n7190), .A(n7193), .ZN(n7189) );
  NAND2_X1 U7825 ( .A1(n6522), .A2(n12335), .ZN(n7190) );
  AND2_X1 U7826 ( .A1(n14247), .A2(n12311), .ZN(n7335) );
  AND2_X1 U7827 ( .A1(n11374), .A2(n7175), .ZN(n7174) );
  NAND2_X1 U7828 ( .A1(n7012), .A2(n7011), .ZN(n14150) );
  INV_X1 U7829 ( .A(n14346), .ZN(n7011) );
  AND2_X1 U7830 ( .A1(n10537), .A2(n11901), .ZN(n10599) );
  OAI21_X1 U7831 ( .B1(n9173), .B2(n9172), .A(n9174), .ZN(n9181) );
  AND2_X1 U7832 ( .A1(n7564), .A2(n9290), .ZN(n7503) );
  XNOR2_X1 U7833 ( .A(n8132), .B(n11605), .ZN(n8106) );
  INV_X1 U7834 ( .A(n7070), .ZN(n7069) );
  INV_X1 U7835 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8524) );
  NOR2_X1 U7836 ( .A1(n7902), .A2(n7420), .ZN(n7419) );
  NAND2_X1 U7837 ( .A1(n7823), .A2(n7593), .ZN(n7596) );
  XNOR2_X1 U7838 ( .A(n6857), .B(P3_ADDR_REG_1__SCAN_IN), .ZN(n14526) );
  INV_X1 U7839 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6857) );
  XNOR2_X1 U7840 ( .A(n6851), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n14521) );
  INV_X1 U7841 ( .A(n6851), .ZN(n14484) );
  OAI22_X1 U7842 ( .A1(n14538), .A2(n14487), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n10837), .ZN(n14488) );
  AOI21_X1 U7843 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n15045), .A(n14491), .ZN(
        n14551) );
  NOR2_X1 U7844 ( .A1(n14546), .A2(n14545), .ZN(n14491) );
  OAI21_X1 U7845 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14499), .A(n14498), .ZN(
        n14514) );
  INV_X1 U7846 ( .A(n12029), .ZN(n7455) );
  NAND2_X1 U7847 ( .A1(n6585), .A2(n6939), .ZN(n6936) );
  NAND2_X1 U7848 ( .A1(n12454), .A2(n6940), .ZN(n6938) );
  OR2_X1 U7849 ( .A1(n8920), .A2(n14675), .ZN(n7456) );
  OR2_X1 U7850 ( .A1(n8937), .A2(n8936), .ZN(n7446) );
  NAND2_X1 U7851 ( .A1(n7441), .A2(n8888), .ZN(n7440) );
  NOR2_X1 U7852 ( .A1(n8311), .A2(n8310), .ZN(n8892) );
  OAI22_X1 U7853 ( .A1(n8412), .A2(n9978), .B1(n10259), .B2(n10243), .ZN(n8311) );
  AOI21_X1 U7854 ( .B1(n12399), .B2(n12400), .A(n7463), .ZN(n7462) );
  INV_X1 U7855 ( .A(n8952), .ZN(n7463) );
  INV_X1 U7856 ( .A(n7459), .ZN(n7458) );
  OAI21_X1 U7857 ( .B1(n6531), .B2(n7460), .A(n12467), .ZN(n7459) );
  INV_X1 U7858 ( .A(n7462), .ZN(n7460) );
  NAND2_X1 U7859 ( .A1(n12373), .A2(n12429), .ZN(n7465) );
  NOR2_X1 U7860 ( .A1(n6500), .A2(n6560), .ZN(n7451) );
  NAND2_X1 U7861 ( .A1(n8513), .A2(n15376), .ZN(n8532) );
  AND4_X1 U7862 ( .A1(n8458), .A2(n8457), .A3(n8456), .A4(n8455), .ZN(n8918)
         );
  OR2_X1 U7863 ( .A1(n8298), .A2(n10226), .ZN(n8279) );
  INV_X1 U7864 ( .A(n8476), .ZN(n8299) );
  NOR2_X1 U7865 ( .A1(n10405), .A2(n10257), .ZN(n10470) );
  XNOR2_X1 U7866 ( .A(n10259), .B(n10248), .ZN(n10467) );
  NOR2_X1 U7867 ( .A1(n10409), .A2(n6903), .ZN(n10466) );
  AND2_X1 U7868 ( .A1(n6891), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n6903) );
  NOR2_X1 U7869 ( .A1(n6963), .A2(n15181), .ZN(n7224) );
  OR2_X1 U7870 ( .A1(n6517), .A2(n11284), .ZN(n7285) );
  NAND2_X1 U7871 ( .A1(n6741), .A2(n6740), .ZN(n15038) );
  NAND2_X1 U7872 ( .A1(n11276), .A2(n7222), .ZN(n6740) );
  OR2_X1 U7873 ( .A1(n11017), .A2(n7219), .ZN(n6741) );
  NAND2_X1 U7874 ( .A1(n7222), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7219) );
  NAND2_X1 U7875 ( .A1(n7285), .A2(n7284), .ZN(n7283) );
  NAND2_X1 U7876 ( .A1(n11835), .A2(n11836), .ZN(n11950) );
  OAI21_X1 U7877 ( .B1(n11291), .B2(n6914), .A(n6913), .ZN(n6912) );
  NAND2_X1 U7878 ( .A1(n6917), .A2(n11949), .ZN(n6914) );
  AOI21_X1 U7879 ( .B1(n6915), .B2(n11290), .A(n6916), .ZN(n6913) );
  NAND2_X1 U7880 ( .A1(n6959), .A2(n6510), .ZN(n6958) );
  INV_X1 U7881 ( .A(n11959), .ZN(n6957) );
  INV_X1 U7882 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8499) );
  XNOR2_X1 U7883 ( .A(n12744), .B(n12745), .ZN(n12727) );
  NOR2_X1 U7884 ( .A1(n12713), .A2(n6902), .ZN(n12733) );
  NOR2_X1 U7885 ( .A1(n11964), .A2(n11943), .ZN(n6902) );
  NAND2_X1 U7886 ( .A1(n12783), .A2(n12784), .ZN(n12807) );
  AOI21_X1 U7887 ( .B1(n12807), .B2(n6745), .A(n12809), .ZN(n12821) );
  INV_X1 U7888 ( .A(n12808), .ZN(n6745) );
  XNOR2_X1 U7889 ( .A(n6726), .B(n6725), .ZN(n6724) );
  INV_X1 U7890 ( .A(n12848), .ZN(n6725) );
  NAND2_X1 U7891 ( .A1(n6728), .A2(n6727), .ZN(n6726) );
  NAND2_X1 U7892 ( .A1(n12850), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n6727) );
  NOR2_X1 U7893 ( .A1(n12852), .A2(n12851), .ZN(n12853) );
  INV_X1 U7894 ( .A(n12676), .ZN(n12670) );
  OR2_X1 U7895 ( .A1(n8764), .A2(n12670), .ZN(n6802) );
  NAND2_X1 U7896 ( .A1(n12932), .A2(n6541), .ZN(n12917) );
  NOR2_X1 U7897 ( .A1(n12933), .A2(n7373), .ZN(n7372) );
  INV_X1 U7898 ( .A(n12649), .ZN(n7373) );
  NAND2_X1 U7899 ( .A1(n8679), .A2(n8678), .ZN(n12941) );
  INV_X1 U7900 ( .A(n12953), .ZN(n6715) );
  INV_X1 U7901 ( .A(n12947), .ZN(n6716) );
  NOR2_X1 U7902 ( .A1(n12991), .A2(n7404), .ZN(n7403) );
  INV_X1 U7903 ( .A(n12630), .ZN(n7404) );
  NAND2_X1 U7904 ( .A1(n13032), .A2(n6807), .ZN(n6803) );
  NAND2_X1 U7905 ( .A1(n13100), .A2(n8788), .ZN(n13011) );
  NAND2_X1 U7906 ( .A1(n12252), .A2(n8560), .ZN(n13034) );
  NAND2_X1 U7907 ( .A1(n12181), .A2(n8539), .ZN(n12254) );
  NAND2_X1 U7908 ( .A1(n6720), .A2(n8483), .ZN(n14645) );
  INV_X1 U7909 ( .A(n8783), .ZN(n14661) );
  OR2_X1 U7910 ( .A1(n14677), .A2(n14657), .ZN(n12590) );
  AND4_X1 U7911 ( .A1(n8439), .A2(n8438), .A3(n8437), .A4(n8436), .ZN(n14674)
         );
  OR2_X1 U7912 ( .A1(n14667), .A2(n14671), .ZN(n14668) );
  INV_X1 U7913 ( .A(n7381), .ZN(n7380) );
  AOI21_X1 U7914 ( .B1(n11566), .B2(n7381), .A(n6498), .ZN(n7379) );
  NOR2_X1 U7915 ( .A1(n8781), .A2(n7382), .ZN(n7381) );
  AND2_X1 U7916 ( .A1(n11570), .A2(n8414), .ZN(n11621) );
  NAND2_X1 U7917 ( .A1(n8413), .A2(n11566), .ZN(n11570) );
  INV_X1 U7918 ( .A(n11568), .ZN(n8413) );
  AOI21_X1 U7919 ( .B1(n15072), .B2(n7214), .A(n6572), .ZN(n7212) );
  INV_X1 U7920 ( .A(n7214), .ZN(n7213) );
  OR2_X1 U7921 ( .A1(n8361), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8377) );
  AND2_X1 U7922 ( .A1(n8968), .A2(n12657), .ZN(n15106) );
  INV_X1 U7923 ( .A(n15078), .ZN(n15112) );
  NAND2_X1 U7924 ( .A1(n15108), .A2(n10583), .ZN(n15110) );
  NAND2_X1 U7925 ( .A1(n12954), .A2(n12953), .ZN(n13077) );
  AND2_X1 U7926 ( .A1(n9916), .A2(n13165), .ZN(n8967) );
  NAND2_X1 U7927 ( .A1(n7445), .A2(n8814), .ZN(n8878) );
  AND2_X1 U7928 ( .A1(n8813), .A2(n7443), .ZN(n7442) );
  NAND2_X1 U7929 ( .A1(n7024), .A2(n12289), .ZN(n12484) );
  NAND2_X1 U7930 ( .A1(n12288), .A2(n12287), .ZN(n7024) );
  NOR2_X1 U7931 ( .A1(n8723), .A2(n7055), .ZN(n7054) );
  INV_X1 U7932 ( .A(n8707), .ZN(n7055) );
  AND2_X1 U7933 ( .A1(n8676), .A2(n8660), .ZN(n8661) );
  NAND2_X1 U7934 ( .A1(n8662), .A2(n8661), .ZN(n8677) );
  NAND2_X1 U7935 ( .A1(n7043), .A2(n7042), .ZN(n8659) );
  INV_X1 U7936 ( .A(n8642), .ZN(n7042) );
  XNOR2_X1 U7937 ( .A(n8622), .B(n11940), .ZN(n8621) );
  NAND2_X1 U7938 ( .A1(n7018), .A2(n8580), .ZN(n8594) );
  NAND2_X1 U7939 ( .A1(n8544), .A2(n8543), .ZN(n8563) );
  AND2_X1 U7940 ( .A1(n8459), .A2(n8443), .ZN(n8444) );
  INV_X1 U7941 ( .A(n8442), .ZN(n7033) );
  OR2_X1 U7942 ( .A1(n8447), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n8462) );
  AND2_X1 U7943 ( .A1(n8442), .A2(n8417), .ZN(n8440) );
  CLKBUF_X1 U7944 ( .A(n8441), .Z(n6885) );
  INV_X1 U7945 ( .A(n7046), .ZN(n7045) );
  OAI21_X1 U7946 ( .B1(n7048), .B2(n7047), .A(n8404), .ZN(n7046) );
  INV_X1 U7947 ( .A(n8401), .ZN(n7047) );
  NAND2_X1 U7948 ( .A1(n8389), .A2(n7048), .ZN(n8402) );
  AND2_X1 U7949 ( .A1(n8369), .A2(n8354), .ZN(n8367) );
  AND2_X1 U7950 ( .A1(n8353), .A2(n8336), .ZN(n8351) );
  INV_X1 U7951 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8337) );
  AND2_X2 U7952 ( .A1(n10246), .A2(n8259), .ZN(n8320) );
  CLKBUF_X1 U7953 ( .A(n10246), .Z(n6891) );
  OR2_X1 U7954 ( .A1(n8149), .A2(n8148), .ZN(n8150) );
  INV_X1 U7955 ( .A(n8171), .ZN(n7080) );
  INV_X1 U7956 ( .A(n7095), .ZN(n7355) );
  OAI21_X1 U7957 ( .B1(n8047), .B2(n13265), .A(n6580), .ZN(n7095) );
  OR2_X1 U7958 ( .A1(n13264), .A2(n13265), .ZN(n7354) );
  AND2_X1 U7959 ( .A1(n8146), .A2(n8122), .ZN(n12267) );
  INV_X1 U7960 ( .A(n13251), .ZN(n6763) );
  NAND2_X1 U7961 ( .A1(n13190), .A2(n6762), .ZN(n6761) );
  AND2_X1 U7962 ( .A1(n13251), .A2(n6858), .ZN(n6762) );
  NAND2_X1 U7963 ( .A1(n7082), .A2(n7087), .ZN(n13282) );
  NAND2_X1 U7964 ( .A1(n12266), .A2(n12267), .ZN(n7082) );
  NOR2_X1 U7965 ( .A1(n6869), .A2(n8221), .ZN(n6682) );
  OR2_X1 U7966 ( .A1(n7869), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n7904) );
  NAND2_X1 U7967 ( .A1(n7659), .A2(n7658), .ZN(n8011) );
  NOR2_X1 U7968 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n7657) );
  NOR2_X1 U7969 ( .A1(n9215), .A2(n13659), .ZN(n7101) );
  OR2_X1 U7970 ( .A1(n13668), .A2(n13296), .ZN(n9231) );
  OR2_X1 U7971 ( .A1(n7247), .A2(n7244), .ZN(n7243) );
  INV_X1 U7972 ( .A(n7250), .ZN(n7244) );
  AND2_X1 U7973 ( .A1(n13468), .A2(n7248), .ZN(n7247) );
  NAND2_X1 U7974 ( .A1(n7554), .A2(n7249), .ZN(n7248) );
  NAND2_X1 U7975 ( .A1(n7554), .A2(n7250), .ZN(n7245) );
  NAND2_X1 U7976 ( .A1(n6698), .A2(n6697), .ZN(n13453) );
  AOI21_X1 U7977 ( .B1(n7243), .B2(n7245), .A(n6699), .ZN(n6698) );
  NAND2_X1 U7978 ( .A1(n13482), .A2(n7243), .ZN(n6697) );
  NAND2_X1 U7979 ( .A1(n13524), .A2(n7098), .ZN(n13474) );
  AND2_X1 U7980 ( .A1(n13415), .A2(n7157), .ZN(n7153) );
  OR2_X1 U7981 ( .A1(n7155), .A2(n7152), .ZN(n6515) );
  INV_X1 U7982 ( .A(n7157), .ZN(n7152) );
  OR2_X1 U7983 ( .A1(n13495), .A2(n13436), .ZN(n13437) );
  NAND2_X1 U7984 ( .A1(n13539), .A2(n7263), .ZN(n7261) );
  NOR2_X1 U7985 ( .A1(n6530), .A2(n7264), .ZN(n7263) );
  INV_X1 U7986 ( .A(n13517), .ZN(n13410) );
  OR2_X1 U7987 ( .A1(n7164), .A2(n13407), .ZN(n7162) );
  NOR2_X1 U7988 ( .A1(n6542), .A2(n7165), .ZN(n7164) );
  NOR2_X1 U7989 ( .A1(n13407), .A2(n7161), .ZN(n7160) );
  INV_X1 U7990 ( .A(n13405), .ZN(n7161) );
  AOI21_X1 U7991 ( .B1(n7126), .B2(n7124), .A(n6565), .ZN(n7123) );
  INV_X1 U7992 ( .A(n7126), .ZN(n7125) );
  INV_X1 U7993 ( .A(n13642), .ZN(n7124) );
  AND2_X1 U7994 ( .A1(n6709), .A2(n13424), .ZN(n6708) );
  OR2_X1 U7995 ( .A1(n6525), .A2(n7255), .ZN(n6709) );
  INV_X1 U7996 ( .A(n7110), .ZN(n13621) );
  NAND2_X1 U7997 ( .A1(n12214), .A2(n12213), .ZN(n13421) );
  AND2_X1 U7998 ( .A1(n7138), .A2(n12162), .ZN(n7135) );
  OR2_X1 U7999 ( .A1(n7136), .A2(n12199), .ZN(n7134) );
  AOI21_X1 U8000 ( .B1(n12160), .B2(n12162), .A(n7137), .ZN(n7136) );
  NAND2_X1 U8001 ( .A1(n7143), .A2(n6494), .ZN(n7142) );
  NAND2_X1 U8002 ( .A1(n6523), .A2(n11814), .ZN(n7144) );
  NAND2_X1 U8003 ( .A1(n7907), .A2(n7906), .ZN(n11816) );
  NAND2_X1 U8004 ( .A1(n7889), .A2(n7888), .ZN(n11663) );
  AND2_X1 U8005 ( .A1(n11244), .A2(n11243), .ZN(n7566) );
  NAND2_X1 U8006 ( .A1(n7566), .A2(n11249), .ZN(n11393) );
  NOR2_X1 U8007 ( .A1(n11249), .A2(n7272), .ZN(n7271) );
  INV_X1 U8008 ( .A(n11248), .ZN(n7272) );
  NAND2_X1 U8009 ( .A1(n11158), .A2(n11157), .ZN(n11246) );
  AND2_X1 U8010 ( .A1(n10067), .A2(n8244), .ZN(n13578) );
  NAND2_X1 U8011 ( .A1(n9197), .A2(n9196), .ZN(n13380) );
  NAND2_X1 U8012 ( .A1(n13801), .A2(n9209), .ZN(n6794) );
  NAND2_X1 U8013 ( .A1(n7643), .A2(n7642), .ZN(n13568) );
  INV_X1 U8014 ( .A(n14994), .ZN(n15009) );
  AND2_X1 U8016 ( .A1(n7545), .A2(n7641), .ZN(n7129) );
  AND3_X1 U8017 ( .A1(n8202), .A2(n7654), .A3(n7653), .ZN(n9924) );
  OR2_X1 U8018 ( .A1(n8011), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n8013) );
  NAND2_X1 U8019 ( .A1(n9909), .A2(n9993), .ZN(n10539) );
  NOR2_X1 U8020 ( .A1(n7302), .A2(n6993), .ZN(n6992) );
  INV_X1 U8021 ( .A(n13842), .ZN(n6993) );
  NAND2_X1 U8022 ( .A1(n7307), .A2(n13849), .ZN(n7302) );
  AND2_X1 U8023 ( .A1(n13997), .A2(n7305), .ZN(n7304) );
  OR2_X1 U8024 ( .A1(n7306), .A2(n14729), .ZN(n7305) );
  AND2_X1 U8025 ( .A1(n13935), .A2(n7317), .ZN(n7316) );
  OR2_X1 U8026 ( .A1(n14006), .A2(n7318), .ZN(n7317) );
  OR2_X1 U8027 ( .A1(n6973), .A2(n6970), .ZN(n6969) );
  INV_X1 U8028 ( .A(n6975), .ZN(n6970) );
  AND2_X1 U8029 ( .A1(n6628), .A2(n11775), .ZN(n6973) );
  AND2_X1 U8030 ( .A1(n12042), .A2(n12041), .ZN(n6493) );
  AND2_X1 U8031 ( .A1(n13831), .A2(n13830), .ZN(n13837) );
  NAND2_X1 U8032 ( .A1(n6981), .A2(n6977), .ZN(n11460) );
  AND2_X1 U8033 ( .A1(n6979), .A2(n6978), .ZN(n6977) );
  NAND2_X1 U8034 ( .A1(n11192), .A2(n6982), .ZN(n6981) );
  NAND2_X1 U8035 ( .A1(n6984), .A2(n6980), .ZN(n6979) );
  INV_X1 U8036 ( .A(n6521), .ZN(n6983) );
  NAND2_X1 U8037 ( .A1(n6521), .A2(n6985), .ZN(n6984) );
  NAND2_X1 U8038 ( .A1(n15194), .A2(n11785), .ZN(n11786) );
  OAI21_X1 U8039 ( .B1(n11460), .B2(n11459), .A(n11458), .ZN(n11613) );
  OR2_X1 U8040 ( .A1(n14114), .A2(n14330), .ZN(n12353) );
  INV_X1 U8041 ( .A(n12341), .ZN(n12342) );
  NOR2_X1 U8042 ( .A1(n14150), .A2(n14130), .ZN(n14129) );
  NAND2_X1 U8043 ( .A1(n14129), .A2(n14118), .ZN(n14114) );
  AND2_X1 U8044 ( .A1(n9810), .A2(n9762), .ZN(n14116) );
  OR2_X1 U8045 ( .A1(n14431), .A2(n14197), .ZN(n6820) );
  NOR2_X1 U8046 ( .A1(n14191), .A2(n7329), .ZN(n7328) );
  INV_X1 U8047 ( .A(n12316), .ZN(n7329) );
  NAND2_X1 U8048 ( .A1(n14208), .A2(n14207), .ZN(n14206) );
  NAND2_X1 U8049 ( .A1(n6893), .A2(n7191), .ZN(n7187) );
  INV_X1 U8050 ( .A(n7189), .ZN(n7188) );
  AND2_X1 U8051 ( .A1(n12314), .A2(n9854), .ZN(n14225) );
  AND2_X1 U8052 ( .A1(n12307), .A2(n12305), .ZN(n7334) );
  NAND2_X1 U8053 ( .A1(n12137), .A2(n12136), .ZN(n12138) );
  NAND2_X1 U8054 ( .A1(n12138), .A2(n12330), .ZN(n12306) );
  NAND2_X1 U8055 ( .A1(n12149), .A2(n12148), .ZN(n12329) );
  NAND2_X1 U8056 ( .A1(n11755), .A2(n9856), .ZN(n11638) );
  NOR2_X1 U8057 ( .A1(n11595), .A2(n7326), .ZN(n7325) );
  INV_X1 U8058 ( .A(n11593), .ZN(n7326) );
  NAND2_X1 U8059 ( .A1(n6582), .A2(n7180), .ZN(n7178) );
  INV_X1 U8060 ( .A(n11369), .ZN(n11374) );
  OR2_X1 U8061 ( .A1(n11194), .A2(n11193), .ZN(n7180) );
  NAND2_X1 U8062 ( .A1(n14814), .A2(n14626), .ZN(n11141) );
  NAND2_X1 U8063 ( .A1(n6769), .A2(n11120), .ZN(n11122) );
  OR2_X1 U8064 ( .A1(n11122), .A2(n11121), .ZN(n11134) );
  INV_X1 U8065 ( .A(n6650), .ZN(n10987) );
  NAND2_X1 U8066 ( .A1(n10987), .A2(n10986), .ZN(n11118) );
  INV_X1 U8067 ( .A(n14626), .ZN(n11043) );
  OR2_X1 U8068 ( .A1(n9354), .A2(n11349), .ZN(n9348) );
  NAND2_X1 U8069 ( .A1(n9828), .A2(n9827), .ZN(n14089) );
  NAND2_X1 U8070 ( .A1(n9789), .A2(n9788), .ZN(n9851) );
  NAND2_X1 U8071 ( .A1(n12367), .A2(n14255), .ZN(n14328) );
  XNOR2_X1 U8072 ( .A(n6854), .B(n12365), .ZN(n6649) );
  NAND2_X1 U8073 ( .A1(n12352), .A2(n6549), .ZN(n6854) );
  INV_X1 U8074 ( .A(n14325), .ZN(n7013) );
  INV_X1 U8075 ( .A(n14614), .ZN(n14831) );
  NAND3_X1 U8076 ( .A1(n9311), .A2(n7503), .A3(n9291), .ZN(n9295) );
  NAND2_X1 U8077 ( .A1(n7503), .A2(n9311), .ZN(n9304) );
  INV_X1 U8078 ( .A(n9304), .ZN(n7338) );
  NOR2_X1 U8079 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7337) );
  NAND2_X1 U8080 ( .A1(n7564), .A2(n9311), .ZN(n7017) );
  INV_X1 U8081 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9323) );
  NAND2_X1 U8082 ( .A1(n6879), .A2(n9306), .ZN(n9608) );
  INV_X1 U8083 ( .A(n9325), .ZN(n6879) );
  XNOR2_X1 U8084 ( .A(n7823), .B(n7824), .ZN(n9969) );
  XNOR2_X1 U8085 ( .A(n14526), .B(n6871), .ZN(n14528) );
  INV_X1 U8086 ( .A(n14527), .ZN(n6871) );
  XNOR2_X1 U8087 ( .A(n14481), .B(n14480), .ZN(n14523) );
  NAND2_X1 U8088 ( .A1(n15393), .A2(n14533), .ZN(n14535) );
  XNOR2_X1 U8089 ( .A(n14521), .B(n10349), .ZN(n14534) );
  NOR2_X1 U8090 ( .A1(n14588), .A2(n14542), .ZN(n14544) );
  AOI21_X1 U8091 ( .B1(n14495), .B2(n14494), .A(n14493), .ZN(n14515) );
  NAND2_X1 U8092 ( .A1(n14758), .A2(n14564), .ZN(n14567) );
  OAI21_X1 U8093 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n14506), .A(n14505), .ZN(
        n14573) );
  AND2_X1 U8094 ( .A1(n11206), .A2(n7467), .ZN(n7466) );
  NAND2_X1 U8095 ( .A1(n11089), .A2(n8906), .ZN(n7467) );
  NAND2_X1 U8096 ( .A1(n8897), .A2(n6943), .ZN(n10688) );
  INV_X1 U8097 ( .A(n10687), .ZN(n6943) );
  OR2_X1 U8098 ( .A1(n8925), .A2(n12412), .ZN(n6944) );
  NAND2_X1 U8099 ( .A1(n8612), .A2(n8611), .ZN(n13090) );
  NOR2_X1 U8100 ( .A1(n12691), .A2(n12690), .ZN(n6890) );
  NOR2_X1 U8101 ( .A1(n12684), .A2(n6826), .ZN(n12520) );
  INV_X1 U8102 ( .A(n12688), .ZN(n6888) );
  NAND2_X1 U8103 ( .A1(n8736), .A2(n8735), .ZN(n12905) );
  NAND2_X1 U8104 ( .A1(n8721), .A2(n8720), .ZN(n12921) );
  INV_X1 U8105 ( .A(n8918), .ZN(n14657) );
  INV_X1 U8106 ( .A(n14674), .ZN(n12707) );
  NAND2_X1 U8107 ( .A1(n6729), .A2(n6960), .ZN(n11016) );
  NAND2_X1 U8108 ( .A1(n6499), .A2(n6961), .ZN(n6960) );
  NAND2_X1 U8109 ( .A1(n6730), .A2(n6558), .ZN(n6729) );
  OR2_X1 U8110 ( .A1(n11017), .A2(n15185), .ZN(n7221) );
  XNOR2_X1 U8111 ( .A(n12733), .B(n12745), .ZN(n12714) );
  OR2_X1 U8112 ( .A1(n12714), .A2(n12716), .ZN(n7280) );
  INV_X1 U8113 ( .A(n12735), .ZN(n7279) );
  INV_X1 U8114 ( .A(n6951), .ZN(n12749) );
  INV_X1 U8115 ( .A(n6835), .ZN(n12765) );
  NAND2_X1 U8116 ( .A1(n6901), .A2(n7277), .ZN(n6659) );
  NAND2_X1 U8117 ( .A1(n12735), .A2(n7281), .ZN(n7277) );
  OR2_X1 U8118 ( .A1(n12714), .A2(n7278), .ZN(n6901) );
  NAND2_X1 U8119 ( .A1(n7281), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7278) );
  OR2_X1 U8120 ( .A1(n12779), .A2(n12778), .ZN(n6661) );
  INV_X1 U8121 ( .A(n6955), .ZN(n12792) );
  INV_X1 U8122 ( .A(n6953), .ZN(n12799) );
  INV_X1 U8123 ( .A(n7298), .ZN(n12814) );
  AND2_X1 U8124 ( .A1(n12803), .A2(n12804), .ZN(n6923) );
  INV_X1 U8125 ( .A(n12855), .ZN(n15052) );
  OR2_X1 U8126 ( .A1(n12812), .A2(n15060), .ZN(n6920) );
  INV_X1 U8127 ( .A(n7229), .ZN(n12832) );
  OR2_X1 U8128 ( .A1(n12803), .A2(n12804), .ZN(n7298) );
  NAND2_X1 U8129 ( .A1(n8546), .A2(n6946), .ZN(n8598) );
  INV_X1 U8130 ( .A(n12860), .ZN(n15054) );
  NAND2_X1 U8131 ( .A1(n7383), .A2(n12573), .ZN(n11619) );
  NAND2_X1 U8132 ( .A1(n11567), .A2(n12569), .ZN(n7383) );
  NOR2_X1 U8133 ( .A1(n12871), .A2(n7559), .ZN(n8877) );
  NAND2_X1 U8134 ( .A1(n8512), .A2(n8511), .ZN(n12243) );
  NOR2_X1 U8135 ( .A1(P3_IR_REG_29__SCAN_IN), .A2(P3_IR_REG_28__SCAN_IN), .ZN(
        n7386) );
  XNOR2_X1 U8136 ( .A(n8373), .B(n8383), .ZN(n11028) );
  INV_X1 U8137 ( .A(n7366), .ZN(n7365) );
  AND2_X1 U8138 ( .A1(n7974), .A2(n7363), .ZN(n7362) );
  NAND2_X1 U8139 ( .A1(n7364), .A2(n7366), .ZN(n7363) );
  INV_X1 U8140 ( .A(n13536), .ZN(n13695) );
  AND2_X1 U8141 ( .A1(n7900), .A2(n7882), .ZN(n7367) );
  NAND2_X1 U8142 ( .A1(n8001), .A2(n8000), .ZN(n13419) );
  NOR2_X1 U8143 ( .A1(n10588), .A2(n7361), .ZN(n7360) );
  INV_X1 U8144 ( .A(n7750), .ZN(n7361) );
  INV_X1 U8145 ( .A(n8994), .ZN(n10421) );
  AOI21_X1 U8146 ( .B1(n13264), .B2(n8047), .A(n13265), .ZN(n13258) );
  NAND2_X1 U8147 ( .A1(n11900), .A2(n9209), .ZN(n7057) );
  AND2_X1 U8148 ( .A1(n13216), .A2(n7937), .ZN(n14862) );
  XNOR2_X1 U8149 ( .A(n7994), .B(n7992), .ZN(n11967) );
  INV_X1 U8150 ( .A(n9176), .ZN(n13295) );
  OR2_X1 U8151 ( .A1(n8247), .A2(n10429), .ZN(n7705) );
  NAND2_X1 U8152 ( .A1(n7702), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7704) );
  NAND2_X1 U8153 ( .A1(n7731), .A2(n7730), .ZN(n10323) );
  NAND2_X1 U8154 ( .A1(n13645), .A2(n7126), .ZN(n13613) );
  NAND2_X1 U8155 ( .A1(n13645), .A2(n13395), .ZN(n13611) );
  NAND2_X1 U8156 ( .A1(n7256), .A2(n7255), .ZN(n13615) );
  NAND2_X1 U8157 ( .A1(n10069), .A2(n6502), .ZN(n7104) );
  NOR2_X1 U8158 ( .A1(n13667), .A2(n6545), .ZN(n6814) );
  NAND2_X1 U8159 ( .A1(n6988), .A2(n13910), .ZN(n6987) );
  NAND2_X1 U8160 ( .A1(n14005), .A2(n14006), .ZN(n6988) );
  INV_X1 U8161 ( .A(n13935), .ZN(n6986) );
  NAND2_X1 U8162 ( .A1(n9770), .A2(n9769), .ZN(n14337) );
  NAND2_X1 U8163 ( .A1(n6995), .A2(n6994), .ZN(n14700) );
  OR2_X1 U8164 ( .A1(n6998), .A2(n6491), .ZN(n6994) );
  NOR2_X1 U8165 ( .A1(n6998), .A2(n6997), .ZN(n6996) );
  NAND2_X1 U8166 ( .A1(n9701), .A2(n9700), .ZN(n14356) );
  INV_X1 U8167 ( .A(n11853), .ZN(n14838) );
  NAND2_X1 U8168 ( .A1(n7300), .A2(n13893), .ZN(n13963) );
  NAND2_X1 U8169 ( .A1(n13971), .A2(n13972), .ZN(n7300) );
  NAND2_X1 U8170 ( .A1(n9612), .A2(n9611), .ZN(n14735) );
  NAND2_X1 U8171 ( .A1(n10567), .A2(n10562), .ZN(n14731) );
  NAND2_X1 U8172 ( .A1(n10570), .A2(n14611), .ZN(n15197) );
  OR2_X1 U8173 ( .A1(n9812), .A2(n10153), .ZN(n9359) );
  AND3_X1 U8174 ( .A1(n9358), .A2(n9357), .A3(n9356), .ZN(n9360) );
  AOI211_X1 U8175 ( .C1(n12353), .C2(n14327), .A(n14096), .B(n14822), .ZN(
        n14325) );
  NAND2_X1 U8176 ( .A1(n14328), .A2(n14323), .ZN(n6845) );
  NAND2_X1 U8177 ( .A1(n6649), .A2(n14631), .ZN(n6648) );
  NAND2_X1 U8178 ( .A1(n14279), .A2(n11042), .ZN(n14307) );
  NAND2_X1 U8179 ( .A1(n9339), .A2(n7170), .ZN(n9362) );
  NAND2_X1 U8180 ( .A1(n9627), .A2(n10189), .ZN(n6658) );
  NOR2_X1 U8181 ( .A1(n9975), .A2(n7406), .ZN(n7170) );
  INV_X1 U8182 ( .A(n7202), .ZN(n7198) );
  AND2_X1 U8183 ( .A1(n7430), .A2(n7429), .ZN(n14103) );
  AND2_X1 U8184 ( .A1(n7430), .A2(n6539), .ZN(n14101) );
  INV_X1 U8185 ( .A(n7201), .ZN(n7199) );
  AND2_X1 U8186 ( .A1(n6603), .A2(n9290), .ZN(n7501) );
  XNOR2_X1 U8187 ( .A(n14528), .B(n10147), .ZN(n15407) );
  NOR2_X1 U8188 ( .A1(n15408), .A2(n15407), .ZN(n15406) );
  OR2_X1 U8189 ( .A1(n15403), .A2(n15404), .ZN(n6833) );
  XNOR2_X1 U8190 ( .A(n6778), .B(n14547), .ZN(n14593) );
  INV_X1 U8191 ( .A(n14555), .ZN(n14556) );
  XOR2_X1 U8192 ( .A(n14516), .B(n14515), .Z(n14755) );
  XNOR2_X1 U8193 ( .A(n14567), .B(n14566), .ZN(n14763) );
  INV_X1 U8194 ( .A(n14565), .ZN(n14566) );
  NAND2_X1 U8195 ( .A1(n6798), .A2(n6831), .ZN(n14770) );
  INV_X1 U8196 ( .A(n14572), .ZN(n6831) );
  XNOR2_X1 U8197 ( .A(n14574), .B(n14573), .ZN(n14775) );
  OAI21_X1 U8198 ( .B1(n14636), .B2(n14635), .A(n14579), .ZN(n14580) );
  XNOR2_X1 U8199 ( .A(n14642), .B(n14641), .ZN(n14639) );
  OAI21_X1 U8200 ( .B1(n14638), .B2(n14639), .A(n11707), .ZN(n7115) );
  NAND2_X1 U8201 ( .A1(n7233), .A2(n9168), .ZN(n9004) );
  INV_X1 U8202 ( .A(n9014), .ZN(n6865) );
  NAND2_X1 U8203 ( .A1(n9475), .A2(n9474), .ZN(n9495) );
  OAI21_X1 U8204 ( .B1(n9457), .B2(n7492), .A(n6896), .ZN(n9474) );
  AND2_X1 U8205 ( .A1(n7491), .A2(n7489), .ZN(n6896) );
  OAI21_X1 U8206 ( .B1(n9029), .B2(n7534), .A(n7533), .ZN(n9034) );
  OR2_X1 U8207 ( .A1(n9027), .A2(n9028), .ZN(n7533) );
  NOR2_X1 U8208 ( .A1(n7536), .A2(n7535), .ZN(n7534) );
  NOR2_X1 U8209 ( .A1(n9038), .A2(n9041), .ZN(n7540) );
  INV_X1 U8210 ( .A(n9038), .ZN(n7539) );
  OAI21_X1 U8211 ( .B1(n11401), .B2(n9152), .A(n9049), .ZN(n9050) );
  NAND2_X1 U8212 ( .A1(n9052), .A2(n9053), .ZN(n9051) );
  NAND2_X1 U8213 ( .A1(n9533), .A2(n9535), .ZN(n6894) );
  INV_X1 U8214 ( .A(n15092), .ZN(n12534) );
  INV_X1 U8215 ( .A(n9605), .ZN(n7515) );
  NAND2_X1 U8216 ( .A1(n6684), .A2(n6683), .ZN(n6861) );
  INV_X1 U8217 ( .A(n9067), .ZN(n6683) );
  NAND2_X1 U8218 ( .A1(n7507), .A2(n6818), .ZN(n7567) );
  AND2_X1 U8219 ( .A1(n7510), .A2(n6819), .ZN(n6818) );
  AOI21_X1 U8220 ( .B1(n9084), .B2(n9083), .A(n9082), .ZN(n6687) );
  OAI21_X1 U8221 ( .B1(n9084), .B2(n9083), .A(n6576), .ZN(n6688) );
  NAND2_X1 U8222 ( .A1(n9088), .A2(n9087), .ZN(n7518) );
  AND2_X1 U8223 ( .A1(n9104), .A2(n7517), .ZN(n7516) );
  NAND2_X1 U8224 ( .A1(n7519), .A2(n6547), .ZN(n7517) );
  AND2_X1 U8225 ( .A1(n9105), .A2(n9103), .ZN(n9104) );
  INV_X1 U8226 ( .A(n7499), .ZN(n7495) );
  NOR2_X1 U8227 ( .A1(n7499), .A2(n7497), .ZN(n7496) );
  NAND2_X1 U8228 ( .A1(n9143), .A2(n7544), .ZN(n7543) );
  INV_X1 U8229 ( .A(n9144), .ZN(n7544) );
  NAND2_X1 U8230 ( .A1(n9151), .A2(n9150), .ZN(n7532) );
  NAND2_X1 U8231 ( .A1(n9702), .A2(n9704), .ZN(n7485) );
  NAND2_X1 U8232 ( .A1(n6672), .A2(n6555), .ZN(n9164) );
  NAND2_X1 U8233 ( .A1(n6674), .A2(n6673), .ZN(n6672) );
  NAND2_X1 U8234 ( .A1(n9738), .A2(n9740), .ZN(n7482) );
  OAI21_X1 U8235 ( .B1(n9803), .B2(n11901), .A(n6856), .ZN(n9330) );
  NAND2_X1 U8236 ( .A1(n9803), .A2(n11981), .ZN(n6856) );
  NAND2_X1 U8237 ( .A1(n7412), .A2(n7627), .ZN(n7411) );
  INV_X1 U8238 ( .A(n8060), .ZN(n7413) );
  AND2_X1 U8239 ( .A1(n6743), .A2(n6742), .ZN(n10261) );
  NAND2_X1 U8240 ( .A1(n10483), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n6742) );
  INV_X1 U8241 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8281) );
  INV_X1 U8242 ( .A(n11003), .ZN(n10964) );
  NAND2_X1 U8243 ( .A1(n7178), .A2(n11322), .ZN(n7175) );
  NAND2_X1 U8244 ( .A1(n11118), .A2(n6651), .ZN(n7176) );
  AND2_X1 U8245 ( .A1(n7179), .A2(n11322), .ZN(n6651) );
  NAND2_X1 U8246 ( .A1(n14802), .A2(n14040), .ZN(n10848) );
  NAND2_X1 U8247 ( .A1(n6791), .A2(n7409), .ZN(n8076) );
  INV_X1 U8248 ( .A(n7410), .ZN(n7409) );
  NAND2_X1 U8249 ( .A1(n7070), .A2(n6504), .ZN(n6791) );
  OAI21_X1 U8250 ( .B1(n7411), .B2(n8060), .A(n8059), .ZN(n7410) );
  NAND2_X1 U8251 ( .A1(n9311), .A2(n7346), .ZN(n9318) );
  NOR2_X1 U8252 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n7346) );
  NAND2_X1 U8253 ( .A1(n7425), .A2(n7423), .ZN(n7422) );
  NAND2_X1 U8254 ( .A1(n7595), .A2(n7426), .ZN(n7423) );
  OAI21_X1 U8255 ( .B1(n14523), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6559), .ZN(
        n6792) );
  INV_X1 U8256 ( .A(n7454), .ZN(n7453) );
  INV_X1 U8257 ( .A(n12682), .ZN(n7378) );
  OAI21_X1 U8258 ( .B1(n12824), .B2(P3_REG2_REG_1__SCAN_IN), .A(n6735), .ZN(
        n6734) );
  NAND2_X1 U8259 ( .A1(n12824), .A2(n10225), .ZN(n6735) );
  NOR2_X1 U8260 ( .A1(n10397), .A2(n6571), .ZN(n10399) );
  OR2_X1 U8261 ( .A1(n10399), .A2(n10400), .ZN(n7290) );
  NAND2_X1 U8262 ( .A1(n11019), .A2(n11020), .ZN(n11021) );
  NOR2_X1 U8263 ( .A1(n11027), .A2(n6899), .ZN(n11283) );
  AND2_X1 U8264 ( .A1(n11028), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n6899) );
  INV_X1 U8265 ( .A(n15039), .ZN(n7222) );
  NAND2_X1 U8266 ( .A1(n12759), .A2(n12758), .ZN(n12781) );
  NAND2_X1 U8267 ( .A1(n8520), .A2(n12603), .ZN(n7398) );
  AND2_X1 U8268 ( .A1(n12603), .A2(n12604), .ZN(n12601) );
  INV_X1 U8269 ( .A(n12573), .ZN(n7382) );
  NAND2_X1 U8270 ( .A1(n11230), .A2(n8396), .ZN(n11568) );
  AND2_X1 U8271 ( .A1(n11309), .A2(n8360), .ZN(n7214) );
  NAND2_X1 U8272 ( .A1(n8359), .A2(n8358), .ZN(n15069) );
  INV_X1 U8273 ( .A(n15072), .ZN(n8358) );
  NAND2_X1 U8274 ( .A1(n10909), .A2(n8900), .ZN(n12550) );
  NAND2_X1 U8275 ( .A1(n15088), .A2(n15107), .ZN(n12536) );
  AOI21_X1 U8276 ( .B1(n7391), .B2(n7389), .A(n7388), .ZN(n7387) );
  INV_X1 U8277 ( .A(n7391), .ZN(n7390) );
  INV_X1 U8278 ( .A(n12590), .ZN(n7389) );
  INV_X1 U8279 ( .A(n11696), .ZN(n8831) );
  INV_X1 U8280 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n7443) );
  NAND2_X1 U8281 ( .A1(n8677), .A2(n8676), .ZN(n8688) );
  INV_X1 U8282 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n6945) );
  INV_X1 U8283 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n8595) );
  AND2_X1 U8284 ( .A1(n8545), .A2(n8549), .ZN(n6948) );
  INV_X1 U8285 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8549) );
  INV_X1 U8286 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8545) );
  NOR2_X1 U8287 ( .A1(n7036), .A2(n7040), .ZN(n7035) );
  INV_X1 U8288 ( .A(n8351), .ZN(n7036) );
  INV_X1 U8289 ( .A(n8367), .ZN(n7040) );
  INV_X1 U8290 ( .A(n8369), .ZN(n7038) );
  NAND2_X1 U8291 ( .A1(n7560), .A2(n7526), .ZN(n7525) );
  OR2_X1 U8292 ( .A1(n9221), .A2(n9253), .ZN(n7552) );
  NAND2_X1 U8293 ( .A1(n7560), .A2(n7528), .ZN(n7527) );
  AND2_X1 U8294 ( .A1(n12284), .A2(n6863), .ZN(n9211) );
  INV_X1 U8295 ( .A(n13437), .ZN(n7249) );
  AND2_X1 U8296 ( .A1(n7099), .A2(n13416), .ZN(n7098) );
  AND2_X1 U8297 ( .A1(n13512), .A2(n13678), .ZN(n7099) );
  AND2_X1 U8298 ( .A1(n7695), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8037) );
  NOR2_X1 U8300 ( .A1(n7142), .A2(n7141), .ZN(n7140) );
  INV_X1 U8301 ( .A(n12004), .ZN(n7141) );
  NOR2_X1 U8302 ( .A1(n7967), .A2(n11807), .ZN(n7987) );
  OR2_X1 U8303 ( .A1(n11249), .A2(n7122), .ZN(n7121) );
  INV_X1 U8304 ( .A(n11392), .ZN(n7122) );
  NAND2_X1 U8305 ( .A1(n11002), .A2(n10966), .ZN(n10968) );
  AND2_X1 U8306 ( .A1(n9237), .A2(n9922), .ZN(n7251) );
  XNOR2_X1 U8307 ( .A(n13310), .B(n10953), .ZN(n10922) );
  NAND2_X1 U8308 ( .A1(n10923), .A2(n10922), .ZN(n10963) );
  NAND2_X1 U8309 ( .A1(n7659), .A2(n7647), .ZN(n7963) );
  OR2_X1 U8310 ( .A1(n7846), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n7865) );
  OR2_X1 U8311 ( .A1(n7787), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n7803) );
  INV_X1 U8312 ( .A(n11446), .ZN(n6980) );
  NAND2_X1 U8313 ( .A1(n6985), .A2(n11446), .ZN(n6982) );
  NAND2_X1 U8314 ( .A1(n6983), .A2(n11191), .ZN(n6978) );
  NAND2_X1 U8315 ( .A1(n9801), .A2(n9800), .ZN(n9840) );
  OR2_X1 U8316 ( .A1(n9802), .A2(n9799), .ZN(n9800) );
  NAND2_X1 U8317 ( .A1(n14417), .A2(n9802), .ZN(n9801) );
  NAND2_X1 U8318 ( .A1(n9771), .A2(n9773), .ZN(n7479) );
  INV_X1 U8319 ( .A(n10599), .ZN(n10600) );
  NOR2_X1 U8320 ( .A1(n14212), .A2(n14193), .ZN(n14181) );
  NOR2_X1 U8321 ( .A1(n14385), .A2(n7005), .ZN(n7004) );
  INV_X1 U8322 ( .A(n7006), .ZN(n7005) );
  NOR2_X1 U8323 ( .A1(n14721), .A2(n14735), .ZN(n7006) );
  OR2_X1 U8324 ( .A1(n13820), .A2(n12139), .ZN(n12136) );
  NOR2_X1 U8325 ( .A1(n12087), .A2(n14602), .ZN(n7009) );
  NOR2_X1 U8326 ( .A1(n11320), .A2(n7333), .ZN(n7332) );
  INV_X1 U8327 ( .A(n11133), .ZN(n7333) );
  NOR2_X1 U8328 ( .A1(n14813), .A2(n11447), .ZN(n11320) );
  INV_X1 U8329 ( .A(n14107), .ZN(n13937) );
  AND2_X1 U8330 ( .A1(n6775), .A2(n14106), .ZN(n6773) );
  INV_X1 U8331 ( .A(n7328), .ZN(n6772) );
  AOI21_X1 U8332 ( .B1(n7328), .B2(n6771), .A(n6506), .ZN(n6770) );
  NOR2_X1 U8333 ( .A1(n11053), .A2(n11045), .ZN(n11044) );
  AND2_X1 U8334 ( .A1(n11044), .A2(n11339), .ZN(n10994) );
  OAI21_X1 U8335 ( .B1(n8173), .B2(n8172), .A(n8175), .ZN(n9173) );
  NOR2_X1 U8336 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n6652) );
  NAND2_X1 U8337 ( .A1(n9320), .A2(n9319), .ZN(n9891) );
  INV_X1 U8338 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9319) );
  INV_X1 U8339 ( .A(n9318), .ZN(n9320) );
  AOI21_X1 U8340 ( .B1(n7092), .B2(n7996), .A(n7091), .ZN(n7090) );
  INV_X1 U8341 ( .A(n7614), .ZN(n7092) );
  INV_X1 U8342 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9286) );
  XNOR2_X1 U8343 ( .A(n7615), .B(SI_16_), .ZN(n7996) );
  AOI21_X1 U8344 ( .B1(n7416), .B2(n7418), .A(n6577), .ZN(n7414) );
  XNOR2_X1 U8345 ( .A(n7607), .B(SI_13_), .ZN(n7938) );
  INV_X1 U8346 ( .A(n7742), .ZN(n6790) );
  OAI211_X1 U8347 ( .C1(n7408), .C2(P1_DATAO_REG_1__SCAN_IN), .A(n6817), .B(
        n6816), .ZN(n7571) );
  NAND2_X1 U8348 ( .A1(n6855), .A2(n9946), .ZN(n6817) );
  NAND2_X1 U8349 ( .A1(n7061), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7408) );
  AOI21_X1 U8350 ( .B1(n7117), .B2(n6878), .A(n14479), .ZN(n14481) );
  AND2_X1 U8351 ( .A1(n14478), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n14479) );
  INV_X1 U8352 ( .A(n14524), .ZN(n6878) );
  INV_X1 U8353 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14478) );
  INV_X1 U8354 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n14480) );
  XNOR2_X1 U8355 ( .A(n6792), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n14522) );
  NOR2_X1 U8356 ( .A1(n14490), .A2(n14489), .ZN(n14546) );
  AND2_X1 U8357 ( .A1(n14520), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14489) );
  OAI21_X1 U8358 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n15067), .A(n14492), .ZN(
        n14519) );
  INV_X1 U8359 ( .A(n7440), .ZN(n7439) );
  AOI21_X1 U8360 ( .B1(n6927), .B2(n6929), .A(n6926), .ZN(n6925) );
  INV_X1 U8361 ( .A(n12389), .ZN(n6926) );
  NAND2_X1 U8362 ( .A1(n8628), .A2(n8627), .ZN(n8647) );
  INV_X1 U8363 ( .A(n12704), .ZN(n12412) );
  NOR2_X1 U8364 ( .A1(n11559), .A2(n7476), .ZN(n7475) );
  INV_X1 U8365 ( .A(n8911), .ZN(n7476) );
  AND2_X1 U8366 ( .A1(n8426), .A2(n8423), .ZN(n8434) );
  NAND2_X1 U8367 ( .A1(n12435), .A2(n6934), .ZN(n6933) );
  INV_X1 U8368 ( .A(n6936), .ZN(n6934) );
  AND2_X1 U8369 ( .A1(n12435), .A2(n6526), .ZN(n6935) );
  NOR2_X1 U8370 ( .A1(n8917), .A2(n8916), .ZN(n11878) );
  NAND2_X1 U8371 ( .A1(n8586), .A2(n8585), .ZN(n8604) );
  OR2_X1 U8372 ( .A1(n8532), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8554) );
  NAND2_X1 U8373 ( .A1(n6829), .A2(n6557), .ZN(n6826) );
  NOR2_X1 U8374 ( .A1(n12680), .A2(n6828), .ZN(n6827) );
  NAND2_X1 U8375 ( .A1(n6843), .A2(n12657), .ZN(n6842) );
  OR2_X1 U8376 ( .A1(n8860), .A2(n8847), .ZN(n12682) );
  CLKBUF_X1 U8377 ( .A(n8476), .Z(n8671) );
  NAND2_X1 U8378 ( .A1(n8747), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7206) );
  AOI22_X1 U8379 ( .A1(n10256), .A2(n10506), .B1(P3_IR_REG_1__SCAN_IN), .B2(
        n10255), .ZN(n10406) );
  NAND2_X1 U8380 ( .A1(n10228), .A2(n6733), .ZN(n10411) );
  OR2_X1 U8381 ( .A1(n6734), .A2(n10416), .ZN(n6733) );
  INV_X1 U8382 ( .A(n6666), .ZN(n10465) );
  NAND2_X1 U8383 ( .A1(n10501), .A2(n7288), .ZN(n6904) );
  AOI21_X1 U8384 ( .B1(n7286), .B2(n10484), .A(n10249), .ZN(n10397) );
  NAND2_X1 U8385 ( .A1(n10486), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10487) );
  AND2_X1 U8386 ( .A1(n6732), .A2(n6731), .ZN(n10392) );
  INV_X1 U8387 ( .A(n10265), .ZN(n6731) );
  NAND2_X1 U8388 ( .A1(n10487), .A2(n10264), .ZN(n6732) );
  NAND2_X1 U8389 ( .A1(n10399), .A2(n10400), .ZN(n7293) );
  NAND2_X1 U8390 ( .A1(n7293), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7292) );
  INV_X1 U8391 ( .A(n7290), .ZN(n10838) );
  INV_X1 U8392 ( .A(n6730), .ZN(n10393) );
  OAI21_X1 U8393 ( .B1(n10829), .B2(n10830), .A(n10828), .ZN(n10831) );
  NAND2_X1 U8394 ( .A1(n10831), .A2(n10832), .ZN(n11019) );
  AND2_X1 U8395 ( .A1(n7290), .A2(n7292), .ZN(n10841) );
  NOR2_X1 U8396 ( .A1(n10841), .A2(n10840), .ZN(n11027) );
  NOR2_X1 U8397 ( .A1(n10826), .A2(n10400), .ZN(n6962) );
  AOI22_X1 U8398 ( .A1(n15033), .A2(n15032), .B1(n15035), .B2(n11297), .ZN(
        n15050) );
  OAI211_X1 U8399 ( .C1(n7285), .C2(n6663), .A(n6507), .B(n6662), .ZN(n15047)
         );
  INV_X1 U8400 ( .A(n6907), .ZN(n6663) );
  NAND2_X1 U8401 ( .A1(n7285), .A2(n6620), .ZN(n6662) );
  NAND2_X1 U8402 ( .A1(n11286), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7282) );
  NOR2_X1 U8403 ( .A1(n15047), .A2(n15048), .ZN(n15046) );
  AND2_X1 U8404 ( .A1(n11286), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n6739) );
  AND2_X1 U8405 ( .A1(n11950), .A2(n11951), .ZN(n11953) );
  AND2_X1 U8406 ( .A1(n11953), .A2(n11954), .ZN(n12718) );
  NOR2_X1 U8407 ( .A1(n12718), .A2(n12719), .ZN(n12720) );
  OR2_X1 U8408 ( .A1(n12746), .A2(n12747), .ZN(n6951) );
  NOR2_X1 U8409 ( .A1(n6738), .A2(n6736), .ZN(n12741) );
  NOR2_X1 U8410 ( .A1(n6737), .A2(n12717), .ZN(n6736) );
  INV_X1 U8411 ( .A(n12736), .ZN(n6738) );
  INV_X1 U8412 ( .A(n12737), .ZN(n6737) );
  NAND2_X1 U8413 ( .A1(n12741), .A2(n12740), .ZN(n12759) );
  INV_X1 U8414 ( .A(n12738), .ZN(n7281) );
  NAND2_X1 U8415 ( .A1(n6955), .A2(n6954), .ZN(n6953) );
  INV_X1 U8416 ( .A(n12791), .ZN(n6954) );
  NOR2_X1 U8417 ( .A1(n6659), .A2(n6635), .ZN(n12774) );
  NAND2_X1 U8418 ( .A1(n7230), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n7227) );
  NAND2_X1 U8419 ( .A1(n12833), .A2(n7230), .ZN(n7226) );
  NAND2_X1 U8420 ( .A1(n6964), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n7229) );
  INV_X1 U8421 ( .A(n12800), .ZN(n6964) );
  AND2_X1 U8422 ( .A1(n6948), .A2(n6947), .ZN(n6946) );
  INV_X1 U8423 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n6947) );
  AND2_X1 U8424 ( .A1(n8527), .A2(n8526), .ZN(n8546) );
  NAND2_X1 U8425 ( .A1(n6802), .A2(n6554), .ZN(n6717) );
  OR2_X1 U8426 ( .A1(n8746), .A2(n12872), .ZN(n12880) );
  NAND2_X1 U8427 ( .A1(n7207), .A2(n8722), .ZN(n12888) );
  NAND2_X1 U8428 ( .A1(n8713), .A2(n8712), .ZN(n8729) );
  AND2_X1 U8429 ( .A1(n8703), .A2(n8702), .ZN(n12936) );
  AND2_X1 U8430 ( .A1(n12950), .A2(n8675), .ZN(n12934) );
  AND2_X1 U8431 ( .A1(n12643), .A2(n12642), .ZN(n12964) );
  AOI21_X1 U8432 ( .B1(n8619), .B2(n6805), .A(n6534), .ZN(n6804) );
  INV_X1 U8433 ( .A(n8619), .ZN(n6806) );
  AOI21_X1 U8434 ( .B1(n7403), .B2(n7401), .A(n7400), .ZN(n7399) );
  INV_X1 U8435 ( .A(n7403), .ZN(n7402) );
  INV_X1 U8436 ( .A(n12634), .ZN(n7400) );
  OR2_X1 U8437 ( .A1(n12516), .A2(n12515), .ZN(n12976) );
  OR2_X1 U8438 ( .A1(n8604), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8613) );
  NAND2_X1 U8439 ( .A1(n13032), .A2(n8576), .ZN(n13018) );
  INV_X1 U8440 ( .A(n13033), .ZN(n13039) );
  OR2_X1 U8441 ( .A1(n12243), .A2(n12705), .ZN(n12603) );
  NAND2_X1 U8442 ( .A1(n6719), .A2(n6621), .ZN(n12127) );
  NAND2_X1 U8443 ( .A1(n14651), .A2(n8921), .ZN(n7211) );
  NAND2_X1 U8444 ( .A1(n8485), .A2(n8484), .ZN(n8514) );
  INV_X1 U8445 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8484) );
  NAND2_X1 U8446 ( .A1(n6799), .A2(n8468), .ZN(n14656) );
  OAI21_X1 U8447 ( .B1(n14672), .B2(n14657), .A(n8467), .ZN(n6799) );
  NAND2_X1 U8448 ( .A1(n8434), .A2(n8433), .ZN(n8477) );
  NAND2_X1 U8449 ( .A1(n6721), .A2(n7209), .ZN(n11685) );
  AOI21_X1 U8450 ( .B1(n12569), .B2(n6488), .A(n7210), .ZN(n7209) );
  NAND2_X1 U8451 ( .A1(n11568), .A2(n6488), .ZN(n6721) );
  INV_X1 U8452 ( .A(n12578), .ZN(n7210) );
  NAND2_X1 U8453 ( .A1(n8780), .A2(n12567), .ZN(n11567) );
  AND2_X1 U8454 ( .A1(n15069), .A2(n8360), .ZN(n11310) );
  NAND2_X1 U8455 ( .A1(n15069), .A2(n7214), .ZN(n11308) );
  INV_X1 U8456 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8345) );
  NAND2_X1 U8457 ( .A1(n12542), .A2(n8775), .ZN(n10935) );
  INV_X1 U8458 ( .A(n15107), .ZN(n10894) );
  NAND2_X1 U8459 ( .A1(n7215), .A2(n8312), .ZN(n10897) );
  NAND2_X1 U8460 ( .A1(n8800), .A2(n8871), .ZN(n15075) );
  INV_X1 U8461 ( .A(n7216), .ZN(n12505) );
  NAND2_X1 U8462 ( .A1(n15111), .A2(n15110), .ZN(n6714) );
  NAND2_X1 U8463 ( .A1(n10580), .A2(n10579), .ZN(n10582) );
  NAND2_X1 U8464 ( .A1(n8728), .A2(n8727), .ZN(n12667) );
  NAND2_X1 U8465 ( .A1(n8626), .A2(n8625), .ZN(n12387) );
  NAND2_X1 U8466 ( .A1(n8531), .A2(n8530), .ZN(n12152) );
  AND3_X1 U8467 ( .A1(n8376), .A2(n8375), .A3(n8374), .ZN(n15147) );
  NAND2_X1 U8468 ( .A1(n7025), .A2(n8844), .ZN(n12288) );
  NAND2_X1 U8469 ( .A1(n7026), .A2(n6639), .ZN(n7025) );
  NAND2_X1 U8470 ( .A1(n8284), .A2(n6877), .ZN(n11977) );
  XNOR2_X1 U8471 ( .A(n8812), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8813) );
  OR2_X1 U8472 ( .A1(n8706), .A2(n8705), .ZN(n8708) );
  NAND2_X1 U8473 ( .A1(n8690), .A2(n8689), .ZN(n8706) );
  OR2_X1 U8474 ( .A1(n8688), .A2(n13806), .ZN(n8689) );
  NAND2_X1 U8475 ( .A1(n8687), .A2(n14473), .ZN(n8690) );
  AND2_X1 U8476 ( .A1(n6529), .A2(n8833), .ZN(n7469) );
  XNOR2_X1 U8477 ( .A(n8834), .B(n8833), .ZN(n10241) );
  NAND2_X1 U8478 ( .A1(n7470), .A2(n6529), .ZN(n8832) );
  NAND2_X1 U8479 ( .A1(n7044), .A2(n8640), .ZN(n8643) );
  CLKBUF_X1 U8480 ( .A(n8759), .Z(n8760) );
  XNOR2_X1 U8481 ( .A(n8758), .B(P3_IR_REG_20__SCAN_IN), .ZN(n8868) );
  OAI21_X1 U8482 ( .B1(n8757), .B2(n8756), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8758) );
  AND2_X1 U8483 ( .A1(n8546), .A2(n8545), .ZN(n8550) );
  NAND2_X1 U8484 ( .A1(n6886), .A2(n7020), .ZN(n8542) );
  AND2_X1 U8485 ( .A1(n6887), .A2(n8525), .ZN(n6886) );
  INV_X1 U8486 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8526) );
  AOI21_X1 U8487 ( .B1(n7031), .B2(n7033), .A(n7028), .ZN(n7027) );
  INV_X1 U8488 ( .A(n8459), .ZN(n7028) );
  AND2_X1 U8489 ( .A1(n8408), .A2(n8407), .ZN(n8418) );
  AND2_X1 U8490 ( .A1(n8384), .A2(n8383), .ZN(n8408) );
  NOR2_X1 U8491 ( .A1(n8372), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8384) );
  INV_X1 U8492 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8383) );
  INV_X1 U8493 ( .A(n7933), .ZN(n7364) );
  AND2_X1 U8494 ( .A1(n14863), .A2(n7937), .ZN(n7366) );
  NOR2_X1 U8495 ( .A1(n13555), .A2(n11674), .ZN(n6858) );
  NOR2_X1 U8496 ( .A1(n7874), .A2(n11266), .ZN(n7890) );
  OR2_X1 U8497 ( .A1(n8002), .A2(n13232), .ZN(n8020) );
  OR2_X1 U8498 ( .A1(n7926), .A2(n7925), .ZN(n7944) );
  OR2_X1 U8499 ( .A1(n7944), .A2(n7943), .ZN(n7967) );
  NAND2_X1 U8500 ( .A1(n13216), .A2(n7366), .ZN(n14861) );
  NOR2_X1 U8501 ( .A1(n8064), .A2(n12297), .ZN(n8084) );
  NAND2_X1 U8502 ( .A1(n8039), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8064) );
  AND2_X1 U8503 ( .A1(n7890), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7909) );
  NAND2_X1 U8504 ( .A1(n7909), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7926) );
  INV_X1 U8505 ( .A(n8181), .ZN(n7234) );
  NOR2_X1 U8506 ( .A1(n8020), .A2(n8019), .ZN(n8021) );
  AND2_X1 U8507 ( .A1(n8021), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7695) );
  OR2_X1 U8508 ( .A1(n7963), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n7981) );
  AOI21_X1 U8509 ( .B1(n12281), .B2(n9209), .A(n9175), .ZN(n13446) );
  INV_X1 U8510 ( .A(n13379), .ZN(n13458) );
  INV_X1 U8511 ( .A(n6515), .ZN(n7151) );
  INV_X1 U8512 ( .A(n7153), .ZN(n7150) );
  AND2_X1 U8513 ( .A1(n13684), .A2(n6840), .ZN(n13414) );
  NAND2_X1 U8514 ( .A1(n13415), .A2(n13500), .ZN(n7156) );
  AND4_X1 U8515 ( .A1(n8168), .A2(n8167), .A3(n8166), .A4(n8165), .ZN(n13484)
         );
  NAND2_X1 U8516 ( .A1(n13539), .A2(n13538), .ZN(n7266) );
  AOI21_X1 U8517 ( .B1(n7240), .B2(n7238), .A(n6578), .ZN(n7237) );
  INV_X1 U8518 ( .A(n13428), .ZN(n7238) );
  INV_X1 U8519 ( .A(n7240), .ZN(n7239) );
  NAND2_X1 U8520 ( .A1(n7108), .A2(n7107), .ZN(n13566) );
  NAND2_X1 U8521 ( .A1(n7110), .A2(n7109), .ZN(n13601) );
  INV_X1 U8522 ( .A(n13395), .ZN(n7127) );
  AOI21_X1 U8523 ( .B1(n7257), .B2(n7259), .A(n6566), .ZN(n7255) );
  NAND2_X1 U8524 ( .A1(n13643), .A2(n13642), .ZN(n13645) );
  NAND2_X1 U8525 ( .A1(n11906), .A2(n11905), .ZN(n11908) );
  NAND2_X1 U8526 ( .A1(n11667), .A2(n11666), .ZN(n11669) );
  OAI21_X1 U8527 ( .B1(n7270), .B2(n11246), .A(n7268), .ZN(n11403) );
  INV_X1 U8528 ( .A(n7271), .ZN(n7270) );
  AOI21_X1 U8529 ( .B1(n7271), .B2(n7269), .A(n6564), .ZN(n7268) );
  INV_X1 U8530 ( .A(n11245), .ZN(n7269) );
  OR2_X1 U8531 ( .A1(n7852), .A2(n7851), .ZN(n7874) );
  NAND2_X1 U8532 ( .A1(n11254), .A2(n11434), .ZN(n11395) );
  INV_X1 U8533 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7810) );
  INV_X1 U8534 ( .A(n11010), .ZN(n7106) );
  AND2_X1 U8535 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7792) );
  NAND2_X1 U8536 ( .A1(n6710), .A2(n11003), .ZN(n11002) );
  NAND2_X1 U8537 ( .A1(n6707), .A2(n10860), .ZN(n10862) );
  INV_X1 U8538 ( .A(n7251), .ZN(n6707) );
  NAND2_X1 U8539 ( .A1(n10863), .A2(n10862), .ZN(n10921) );
  NAND2_X1 U8540 ( .A1(n7251), .A2(n10860), .ZN(n10861) );
  NAND2_X1 U8541 ( .A1(n12165), .A2(n12164), .ZN(n12166) );
  AND2_X1 U8542 ( .A1(n9920), .A2(n13692), .ZN(n14994) );
  INV_X1 U8543 ( .A(n8236), .ZN(n10635) );
  NAND2_X1 U8544 ( .A1(n6671), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6670) );
  INV_X1 U8545 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8207) );
  OR2_X1 U8546 ( .A1(n8202), .A2(n8201), .ZN(n8206) );
  NAND2_X1 U8547 ( .A1(n7659), .A2(n7644), .ZN(n8202) );
  NAND2_X1 U8548 ( .A1(n6574), .A2(n7659), .ZN(n8198) );
  OAI21_X1 U8549 ( .B1(n8013), .B2(n7667), .A(n7666), .ZN(n8235) );
  INV_X1 U8550 ( .A(n6999), .ZN(n6997) );
  NAND2_X1 U8551 ( .A1(n9637), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9650) );
  INV_X1 U8552 ( .A(n7316), .ZN(n7313) );
  AOI21_X1 U8553 ( .B1(n7316), .B2(n7318), .A(n6581), .ZN(n7315) );
  NOR2_X1 U8554 ( .A1(n9650), .A2(n13983), .ZN(n9662) );
  NOR2_X1 U8555 ( .A1(n13955), .A2(n7321), .ZN(n7320) );
  INV_X1 U8556 ( .A(n13868), .ZN(n7321) );
  OR2_X1 U8557 ( .A1(n9592), .A2(n9284), .ZN(n9614) );
  NOR2_X1 U8558 ( .A1(n10540), .A2(n7349), .ZN(n10543) );
  INV_X1 U8559 ( .A(n11141), .ZN(n7347) );
  INV_X1 U8560 ( .A(n12231), .ZN(n7341) );
  AOI21_X1 U8561 ( .B1(n7344), .B2(n6493), .A(n6629), .ZN(n7343) );
  NAND2_X1 U8562 ( .A1(n6615), .A2(n7344), .ZN(n7342) );
  OR2_X1 U8563 ( .A1(n9508), .A2(n9507), .ZN(n9523) );
  NOR2_X1 U8564 ( .A1(n11924), .A2(n7000), .ZN(n6999) );
  INV_X1 U8565 ( .A(n7001), .ZN(n7000) );
  NAND2_X1 U8566 ( .A1(n11921), .A2(n11920), .ZN(n7001) );
  NAND2_X1 U8567 ( .A1(n14717), .A2(n13842), .ZN(n14730) );
  AND4_X1 U8568 ( .A1(n9561), .A2(n9560), .A3(n9559), .A4(n9558), .ZN(n12224)
         );
  OR2_X1 U8569 ( .A1(n9354), .A2(n9353), .ZN(n9357) );
  NAND2_X1 U8570 ( .A1(n14346), .A2(n12319), .ZN(n12320) );
  AND2_X1 U8571 ( .A1(n14156), .A2(n12339), .ZN(n14148) );
  NAND2_X1 U8572 ( .A1(n6657), .A2(n7181), .ZN(n14156) );
  NOR2_X1 U8573 ( .A1(n14162), .A2(n7182), .ZN(n7181) );
  INV_X1 U8574 ( .A(n12338), .ZN(n7182) );
  NAND2_X1 U8575 ( .A1(n14181), .A2(n12345), .ZN(n14182) );
  AND2_X1 U8576 ( .A1(n14190), .A2(n12336), .ZN(n7550) );
  AOI21_X1 U8577 ( .B1(n7186), .B2(n7184), .A(n6567), .ZN(n7183) );
  NOR2_X1 U8578 ( .A1(n9614), .A2(n9613), .ZN(n9621) );
  NAND2_X1 U8579 ( .A1(n14294), .A2(n7004), .ZN(n14262) );
  NOR2_X1 U8580 ( .A1(n13828), .A2(n12143), .ZN(n14294) );
  NAND2_X1 U8581 ( .A1(n14294), .A2(n14398), .ZN(n14293) );
  NAND2_X1 U8582 ( .A1(n11750), .A2(n7007), .ZN(n12143) );
  AND2_X1 U8583 ( .A1(n6495), .A2(n7008), .ZN(n7007) );
  NAND2_X1 U8584 ( .A1(n11750), .A2(n6495), .ZN(n14610) );
  NAND2_X1 U8585 ( .A1(n6655), .A2(n7513), .ZN(n12149) );
  AND2_X1 U8586 ( .A1(n9556), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9579) );
  NAND2_X1 U8587 ( .A1(n11750), .A2(n11919), .ZN(n12107) );
  AND2_X1 U8588 ( .A1(n11640), .A2(n14838), .ZN(n11750) );
  AND2_X1 U8589 ( .A1(n7551), .A2(n11379), .ZN(n7172) );
  NAND2_X1 U8590 ( .A1(n11594), .A2(n11593), .ZN(n11596) );
  AND2_X1 U8591 ( .A1(n11589), .A2(n11796), .ZN(n11640) );
  NOR2_X1 U8592 ( .A1(n11533), .A2(n15198), .ZN(n11589) );
  AND3_X1 U8593 ( .A1(n7010), .A2(n11044), .A3(n14306), .ZN(n11138) );
  NOR2_X1 U8594 ( .A1(n10982), .A2(n14809), .ZN(n7010) );
  NAND2_X1 U8595 ( .A1(n10994), .A2(n14306), .ZN(n11127) );
  XNOR2_X1 U8596 ( .A(n14040), .B(n11053), .ZN(n11048) );
  NAND2_X1 U8597 ( .A1(n11054), .A2(n11045), .ZN(n10849) );
  NAND2_X1 U8598 ( .A1(n14814), .A2(n11043), .ZN(n10594) );
  INV_X1 U8599 ( .A(n11045), .ZN(n11351) );
  AND2_X1 U8600 ( .A1(n12346), .A2(n12353), .ZN(n14329) );
  NAND2_X1 U8601 ( .A1(n9659), .A2(n9658), .ZN(n14231) );
  INV_X1 U8602 ( .A(n9633), .ZN(n9826) );
  INV_X1 U8603 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9291) );
  OAI211_X1 U8604 ( .C1(n9202), .C2(n9194), .A(n9193), .B(n9192), .ZN(n13785)
         );
  NAND2_X1 U8605 ( .A1(n9202), .A2(n9201), .ZN(n9206) );
  XNOR2_X1 U8606 ( .A(n9181), .B(n9180), .ZN(n12281) );
  XNOR2_X1 U8607 ( .A(n9173), .B(n9172), .ZN(n13790) );
  XNOR2_X1 U8608 ( .A(n9908), .B(P1_IR_REG_26__SCAN_IN), .ZN(n9993) );
  NAND2_X1 U8609 ( .A1(n9907), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9908) );
  INV_X1 U8610 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9900) );
  NAND2_X1 U8611 ( .A1(n9901), .A2(n9900), .ZN(n9907) );
  INV_X1 U8612 ( .A(n9905), .ZN(n9901) );
  XNOR2_X1 U8613 ( .A(n8112), .B(n8111), .ZN(n13801) );
  NAND2_X1 U8614 ( .A1(n9311), .A2(n7002), .ZN(n9905) );
  AND2_X1 U8615 ( .A1(n9893), .A2(n9288), .ZN(n7002) );
  XNOR2_X1 U8616 ( .A(n8106), .B(n8124), .ZN(n9715) );
  INV_X1 U8617 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n15226) );
  XNOR2_X1 U8618 ( .A(n7632), .B(n7631), .ZN(n11980) );
  NAND2_X1 U8619 ( .A1(n7070), .A2(n7623), .ZN(n7679) );
  NAND2_X1 U8620 ( .A1(n7069), .A2(n7623), .ZN(n7690) );
  NAND2_X1 U8621 ( .A1(n7433), .A2(n7623), .ZN(n7687) );
  INV_X1 U8622 ( .A(n7435), .ZN(n7437) );
  NAND2_X1 U8623 ( .A1(n7415), .A2(n7605), .ZN(n7921) );
  NAND2_X1 U8624 ( .A1(n7886), .A2(n7419), .ZN(n7415) );
  NAND2_X1 U8625 ( .A1(n7886), .A2(n7602), .ZN(n7903) );
  OR2_X1 U8626 ( .A1(n9502), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n9544) );
  AND2_X1 U8627 ( .A1(n7886), .A2(n7885), .ZN(n10221) );
  OR2_X1 U8628 ( .A1(n9466), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9587) );
  NAND2_X1 U8629 ( .A1(n7596), .A2(n7595), .ZN(n7845) );
  OR2_X1 U8630 ( .A1(n9450), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n9466) );
  NOR2_X1 U8631 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9340) );
  XNOR2_X1 U8632 ( .A(n7571), .B(SI_1_), .ZN(n7708) );
  XOR2_X1 U8633 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), .Z(
        n14524) );
  OAI22_X1 U8634 ( .A1(n14526), .A2(n14527), .B1(P1_ADDR_REG_1__SCAN_IN), .B2(
        n7118), .ZN(n7117) );
  INV_X1 U8635 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n7118) );
  XNOR2_X1 U8636 ( .A(n14522), .B(n10779), .ZN(n14531) );
  NAND2_X1 U8637 ( .A1(n6777), .A2(n14536), .ZN(n14541) );
  NOR2_X1 U8638 ( .A1(n14486), .A2(n14485), .ZN(n14538) );
  INV_X1 U8639 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14537) );
  NAND2_X1 U8640 ( .A1(n6779), .A2(n6551), .ZN(n6778) );
  OAI21_X1 U8641 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n14501), .A(n14500), .ZN(
        n14512) );
  NAND2_X1 U8642 ( .A1(n11090), .A2(n8906), .ZN(n11207) );
  NAND2_X1 U8643 ( .A1(n7452), .A2(n7454), .ZN(n12119) );
  AND2_X1 U8644 ( .A1(n7477), .A2(n6508), .ZN(n11653) );
  NAND2_X1 U8645 ( .A1(n6937), .A2(n6940), .ZN(n12381) );
  OR2_X1 U8646 ( .A1(n12455), .A2(n12454), .ZN(n6937) );
  NAND2_X1 U8647 ( .A1(n11359), .A2(n11358), .ZN(n11357) );
  AND2_X1 U8648 ( .A1(n8891), .A2(n8888), .ZN(n10650) );
  NAND2_X1 U8649 ( .A1(n7439), .A2(n8891), .ZN(n10649) );
  NAND2_X1 U8650 ( .A1(n12428), .A2(n8948), .ZN(n7461) );
  NAND2_X1 U8651 ( .A1(n10814), .A2(n8902), .ZN(n10907) );
  NAND2_X1 U8652 ( .A1(n8567), .A2(n8566), .ZN(n13041) );
  AND2_X1 U8653 ( .A1(n7465), .A2(n7464), .ZN(n12398) );
  AND2_X1 U8654 ( .A1(n10688), .A2(n8899), .ZN(n10815) );
  NAND2_X1 U8655 ( .A1(n11357), .A2(n8911), .ZN(n11558) );
  NAND2_X1 U8656 ( .A1(n6931), .A2(n6933), .ZN(n12437) );
  NAND2_X1 U8657 ( .A1(n12455), .A2(n6935), .ZN(n6931) );
  NAND2_X1 U8658 ( .A1(n6932), .A2(n6936), .ZN(n12436) );
  NAND2_X1 U8659 ( .A1(n12455), .A2(n6526), .ZN(n6932) );
  NAND2_X1 U8660 ( .A1(n8919), .A2(n7456), .ZN(n12031) );
  NAND2_X1 U8661 ( .A1(n8646), .A2(n8645), .ZN(n12966) );
  OR2_X1 U8662 ( .A1(n11088), .A2(n11089), .ZN(n11090) );
  NAND2_X1 U8663 ( .A1(n7457), .A2(n7462), .ZN(n12465) );
  NOR2_X1 U8664 ( .A1(n7449), .A2(n7448), .ZN(n7447) );
  INV_X1 U8665 ( .A(n12154), .ZN(n7448) );
  INV_X1 U8666 ( .A(n7451), .ZN(n7449) );
  AND2_X1 U8667 ( .A1(n7450), .A2(n7451), .ZN(n12155) );
  AND2_X1 U8668 ( .A1(n8960), .A2(n8967), .ZN(n12468) );
  INV_X1 U8669 ( .A(n12936), .ZN(n12904) );
  OR2_X1 U8670 ( .A1(n9916), .A2(n10027), .ZN(n12703) );
  INV_X1 U8671 ( .A(n12418), .ZN(n13021) );
  NAND4_X1 U8672 ( .A1(n8366), .A2(n8365), .A3(n8364), .A4(n8363), .ZN(n15073)
         );
  NAND4_X1 U8673 ( .A1(n8350), .A2(n8349), .A3(n8348), .A4(n8347), .ZN(n12711)
         );
  INV_X1 U8674 ( .A(n6743), .ZN(n10469) );
  NAND2_X1 U8675 ( .A1(n7223), .A2(n7225), .ZN(n10394) );
  AND2_X1 U8676 ( .A1(n7223), .A2(n7224), .ZN(n10824) );
  INV_X1 U8677 ( .A(n7285), .ZN(n15031) );
  INV_X1 U8678 ( .A(n7283), .ZN(n15029) );
  INV_X1 U8679 ( .A(n11276), .ZN(n7220) );
  INV_X1 U8680 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15067) );
  INV_X1 U8681 ( .A(n6919), .ZN(n11830) );
  INV_X1 U8682 ( .A(n6959), .ZN(n11843) );
  NAND2_X1 U8683 ( .A1(n6911), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n6910) );
  NAND2_X1 U8684 ( .A1(n6958), .A2(n6956), .ZN(n12725) );
  NOR2_X1 U8685 ( .A1(n6511), .A2(n11958), .ZN(n11960) );
  NAND2_X1 U8686 ( .A1(n8473), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8474) );
  INV_X1 U8687 ( .A(n6744), .ZN(n12789) );
  INV_X1 U8688 ( .A(n12806), .ZN(n6921) );
  INV_X1 U8689 ( .A(n12815), .ZN(n7297) );
  NAND2_X1 U8690 ( .A1(n7299), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7296) );
  INV_X1 U8691 ( .A(n12816), .ZN(n7299) );
  OAI21_X1 U8692 ( .B1(n12856), .B2(n12855), .A(n6723), .ZN(n6892) );
  AOI21_X1 U8693 ( .B1(n6724), .B2(n12862), .A(n12861), .ZN(n6723) );
  INV_X1 U8694 ( .A(n6802), .ZN(n8841) );
  AND2_X1 U8695 ( .A1(n12932), .A2(n8686), .ZN(n12919) );
  AND2_X1 U8696 ( .A1(n12931), .A2(n12930), .ZN(n13069) );
  NAND2_X1 U8697 ( .A1(n13077), .A2(n12649), .ZN(n12929) );
  NAND2_X1 U8698 ( .A1(n13011), .A2(n7403), .ZN(n12994) );
  NAND2_X1 U8699 ( .A1(n13011), .A2(n12630), .ZN(n12992) );
  NAND2_X1 U8700 ( .A1(n6803), .A2(n8619), .ZN(n12986) );
  NAND2_X1 U8701 ( .A1(n8584), .A2(n8583), .ZN(n13098) );
  NAND2_X1 U8702 ( .A1(n15083), .A2(n15080), .ZN(n13044) );
  AND2_X1 U8703 ( .A1(n15122), .A2(n14676), .ZN(n14664) );
  NAND2_X1 U8704 ( .A1(n14668), .A2(n12590), .ZN(n14662) );
  NAND2_X1 U8705 ( .A1(n11570), .A2(n6488), .ZN(n11620) );
  NOR2_X1 U8706 ( .A1(n10582), .A2(n15090), .ZN(n15083) );
  INV_X1 U8707 ( .A(n15117), .ZN(n15090) );
  NAND2_X1 U8708 ( .A1(n10581), .A2(n15090), .ZN(n15089) );
  AND2_X1 U8709 ( .A1(n15122), .A2(n15102), .ZN(n15120) );
  NAND2_X1 U8710 ( .A1(n10582), .A2(n15089), .ZN(n15122) );
  INV_X1 U8711 ( .A(n13122), .ZN(n13052) );
  NAND2_X1 U8712 ( .A1(n13167), .A2(n12487), .ZN(n7050) );
  INV_X1 U8713 ( .A(n12667), .ZN(n13129) );
  INV_X1 U8714 ( .A(n12464), .ZN(n13133) );
  NAND2_X1 U8715 ( .A1(n8603), .A2(n8602), .ZN(n13151) );
  AOI21_X1 U8716 ( .B1(n10381), .B2(n12487), .A(n8553), .ZN(n13158) );
  OR2_X1 U8717 ( .A1(n8412), .A2(n8294), .ZN(n8296) );
  AND2_X1 U8718 ( .A1(n10241), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13165) );
  INV_X1 U8719 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8273) );
  INV_X1 U8720 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n8271) );
  OR2_X1 U8721 ( .A1(n8662), .A2(n8661), .ZN(n8663) );
  INV_X1 U8722 ( .A(SI_21_), .ZN(n15362) );
  INV_X1 U8723 ( .A(n8868), .ZN(n10890) );
  INV_X1 U8724 ( .A(n8621), .ZN(n8620) );
  CLKBUF_X1 U8725 ( .A(n8880), .Z(n12859) );
  INV_X1 U8726 ( .A(SI_17_), .ZN(n10518) );
  INV_X1 U8727 ( .A(SI_15_), .ZN(n15360) );
  NAND2_X1 U8728 ( .A1(n8507), .A2(n7022), .ZN(n8523) );
  NAND2_X1 U8729 ( .A1(n8505), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7022) );
  INV_X1 U8730 ( .A(SI_13_), .ZN(n10115) );
  INV_X1 U8731 ( .A(SI_12_), .ZN(n9982) );
  OAI21_X1 U8732 ( .B1(n6885), .B2(n7033), .A(n7031), .ZN(n8460) );
  NAND2_X1 U8733 ( .A1(n7030), .A2(n8442), .ZN(n8445) );
  XNOR2_X1 U8734 ( .A(n8449), .B(n8448), .ZN(n11842) );
  NAND2_X1 U8735 ( .A1(n8402), .A2(n8401), .ZN(n8405) );
  XNOR2_X1 U8736 ( .A(n8409), .B(n7369), .ZN(n11286) );
  OR2_X1 U8737 ( .A1(n8418), .A2(n8273), .ZN(n8409) );
  NAND2_X1 U8738 ( .A1(n8389), .A2(n8388), .ZN(n8392) );
  NAND2_X1 U8739 ( .A1(n7041), .A2(n8353), .ZN(n8368) );
  NAND2_X1 U8740 ( .A1(n8352), .A2(n8351), .ZN(n7041) );
  AND2_X1 U8741 ( .A1(n8340), .A2(n8372), .ZN(n10390) );
  NAND2_X1 U8742 ( .A1(n6900), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8308) );
  OR2_X1 U8743 ( .A1(n9915), .A2(n9914), .ZN(n10072) );
  NAND2_X1 U8744 ( .A1(n13282), .A2(n8150), .ZN(n13180) );
  NAND2_X1 U8745 ( .A1(n7078), .A2(n7083), .ZN(n13182) );
  OR2_X1 U8746 ( .A1(n12266), .A2(n7085), .ZN(n7078) );
  NAND2_X1 U8747 ( .A1(n11261), .A2(n7882), .ZN(n11410) );
  NOR2_X1 U8748 ( .A1(n13444), .A2(n8233), .ZN(n8234) );
  AOI21_X1 U8749 ( .B1(n7081), .B2(n7079), .A(n6513), .ZN(n6750) );
  NAND2_X1 U8750 ( .A1(n7354), .A2(n6489), .ZN(n13210) );
  NAND2_X1 U8751 ( .A1(n7086), .A2(n12267), .ZN(n12269) );
  NAND2_X1 U8752 ( .A1(n11968), .A2(n7995), .ZN(n13229) );
  INV_X1 U8753 ( .A(n13230), .ZN(n7359) );
  NAND2_X1 U8754 ( .A1(n13191), .A2(n7547), .ZN(n13250) );
  NAND2_X1 U8755 ( .A1(n10586), .A2(n7782), .ZN(n10659) );
  AND2_X1 U8756 ( .A1(n13200), .A2(n8034), .ZN(n6867) );
  INV_X1 U8757 ( .A(n8049), .ZN(n7056) );
  NOR2_X1 U8758 ( .A1(n12295), .A2(n8071), .ZN(n12304) );
  NAND2_X1 U8759 ( .A1(n11500), .A2(n7901), .ZN(n7919) );
  NAND2_X1 U8760 ( .A1(n13248), .A2(n6759), .ZN(n13272) );
  NOR2_X1 U8761 ( .A1(n13270), .A2(n6760), .ZN(n6759) );
  INV_X1 U8762 ( .A(n8029), .ZN(n6760) );
  NAND2_X1 U8763 ( .A1(n13248), .A2(n8029), .ZN(n13271) );
  AND2_X1 U8764 ( .A1(n7821), .A2(n7800), .ZN(n7368) );
  NAND2_X1 U8765 ( .A1(n10669), .A2(n7800), .ZN(n10793) );
  AND2_X1 U8766 ( .A1(n8232), .A2(n10631), .ZN(n14860) );
  NAND2_X1 U8767 ( .A1(n8238), .A2(n14950), .ZN(n14867) );
  INV_X1 U8768 ( .A(n9923), .ZN(n10616) );
  NAND2_X1 U8769 ( .A1(n6682), .A2(n10637), .ZN(n6678) );
  OAI21_X1 U8770 ( .B1(n6682), .B2(n9265), .A(n9266), .ZN(n6677) );
  NAND2_X1 U8771 ( .A1(n9261), .A2(n9260), .ZN(n6679) );
  AND2_X1 U8772 ( .A1(n8014), .A2(n8013), .ZN(n14937) );
  XNOR2_X1 U8773 ( .A(n13387), .B(n13750), .ZN(n7102) );
  OR2_X1 U8774 ( .A1(n8183), .A2(n8254), .ZN(n13447) );
  NAND2_X1 U8775 ( .A1(n13453), .A2(n6830), .ZN(n13440) );
  NAND2_X1 U8776 ( .A1(n7097), .A2(n13296), .ZN(n6830) );
  OAI21_X1 U8777 ( .B1(n13482), .B2(n7245), .A(n7243), .ZN(n13455) );
  NAND2_X1 U8778 ( .A1(n6515), .A2(n7147), .ZN(n13479) );
  NAND2_X1 U8779 ( .A1(n7153), .A2(n13500), .ZN(n7147) );
  OAI21_X1 U8780 ( .B1(n13500), .B2(n7151), .A(n7148), .ZN(n13670) );
  NAND2_X1 U8781 ( .A1(n7246), .A2(n7554), .ZN(n13469) );
  NAND2_X1 U8782 ( .A1(n13482), .A2(n13437), .ZN(n7246) );
  NAND2_X1 U8783 ( .A1(n7261), .A2(n7262), .ZN(n13503) );
  NAND2_X1 U8784 ( .A1(n7158), .A2(n7162), .ZN(n13531) );
  NAND2_X1 U8785 ( .A1(n13565), .A2(n7160), .ZN(n7158) );
  NAND2_X1 U8786 ( .A1(n7163), .A2(n13405), .ZN(n13546) );
  OR2_X1 U8787 ( .A1(n13565), .A2(n13404), .ZN(n7163) );
  NAND2_X1 U8788 ( .A1(n7242), .A2(n13429), .ZN(n13560) );
  NAND2_X1 U8789 ( .A1(n13575), .A2(n13428), .ZN(n7242) );
  NAND2_X1 U8790 ( .A1(n13421), .A2(n13420), .ZN(n13629) );
  NAND2_X1 U8791 ( .A1(n7130), .A2(n7134), .ZN(n12202) );
  NAND2_X1 U8792 ( .A1(n12161), .A2(n7135), .ZN(n7130) );
  OAI21_X1 U8793 ( .B1(n12161), .B2(n12160), .A(n12162), .ZN(n12201) );
  NAND2_X1 U8794 ( .A1(n7139), .A2(n7142), .ZN(n12005) );
  NAND2_X1 U8795 ( .A1(n11813), .A2(n6630), .ZN(n7139) );
  OAI21_X1 U8796 ( .B1(n11813), .B2(n6523), .A(n11814), .ZN(n11904) );
  NAND2_X1 U8797 ( .A1(n11393), .A2(n11392), .ZN(n11515) );
  NAND2_X1 U8798 ( .A1(n7273), .A2(n7271), .ZN(n11402) );
  NAND2_X1 U8799 ( .A1(n7273), .A2(n11248), .ZN(n11250) );
  NOR2_X1 U8800 ( .A1(n9919), .A2(n7254), .ZN(n10617) );
  INV_X1 U8801 ( .A(n13380), .ZN(n13750) );
  OR2_X1 U8802 ( .A1(n13725), .A2(n13724), .ZN(n13773) );
  NAND2_X1 U8803 ( .A1(n7986), .A2(n7985), .ZN(n13782) );
  NAND2_X1 U8804 ( .A1(n7872), .A2(n7871), .ZN(n11554) );
  INV_X2 U8805 ( .A(n15017), .ZN(n15018) );
  AND2_X1 U8806 ( .A1(n8239), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14973) );
  AND2_X1 U8807 ( .A1(n7129), .A2(n7671), .ZN(n7128) );
  NAND2_X1 U8808 ( .A1(n6702), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7670) );
  AND2_X1 U8809 ( .A1(n7558), .A2(n7129), .ZN(n6703) );
  AND2_X1 U8810 ( .A1(n6671), .A2(n6669), .ZN(n6668) );
  NAND2_X1 U8811 ( .A1(n7546), .A2(n6562), .ZN(n6667) );
  NAND2_X1 U8812 ( .A1(n7545), .A2(n13786), .ZN(n6669) );
  INV_X1 U8813 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12285) );
  CLKBUF_X1 U8814 ( .A(n8235), .Z(n12284) );
  INV_X1 U8815 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11348) );
  INV_X1 U8816 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10791) );
  INV_X1 U8817 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10504) );
  OR2_X1 U8818 ( .A1(n7659), .A2(n13786), .ZN(n7922) );
  INV_X1 U8819 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10380) );
  INV_X1 U8820 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10222) );
  INV_X1 U8821 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10059) );
  INV_X1 U8822 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9970) );
  INV_X1 U8823 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9968) );
  INV_X1 U8824 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9958) );
  INV_X1 U8825 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9963) );
  INV_X1 U8826 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9960) );
  INV_X1 U8827 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9956) );
  AND2_X1 U8828 ( .A1(n6974), .A2(n6628), .ZN(n11776) );
  NAND2_X1 U8829 ( .A1(n11613), .A2(n11611), .ZN(n6974) );
  NAND2_X1 U8830 ( .A1(n9455), .A2(n9454), .ZN(n11536) );
  NAND2_X1 U8831 ( .A1(n11859), .A2(n11858), .ZN(n11922) );
  NAND2_X1 U8832 ( .A1(n11111), .A2(n11110), .ZN(n11112) );
  OAI21_X1 U8833 ( .B1(n13838), .B2(n6991), .A(n6989), .ZN(n13926) );
  INV_X1 U8834 ( .A(n6992), .ZN(n6991) );
  AND2_X1 U8835 ( .A1(n6992), .A2(n14013), .ZN(n6990) );
  NAND2_X1 U8836 ( .A1(n13926), .A2(n13925), .ZN(n13924) );
  NAND2_X1 U8837 ( .A1(n7311), .A2(n7310), .ZN(n7309) );
  NAND2_X1 U8838 ( .A1(n7319), .A2(n7315), .ZN(n7310) );
  NAND2_X1 U8839 ( .A1(n13944), .A2(n7312), .ZN(n7311) );
  NAND2_X1 U8840 ( .A1(n7315), .A2(n7313), .ZN(n7312) );
  NAND2_X1 U8841 ( .A1(n13944), .A2(n7315), .ZN(n7314) );
  NAND2_X1 U8842 ( .A1(n6965), .A2(n6969), .ZN(n15196) );
  NAND2_X1 U8843 ( .A1(n11613), .A2(n6971), .ZN(n6965) );
  NOR2_X1 U8844 ( .A1(n10718), .A2(n10803), .ZN(n10722) );
  NAND2_X1 U8845 ( .A1(n13978), .A2(n13868), .ZN(n13954) );
  NOR2_X1 U8846 ( .A1(n6615), .A2(n6493), .ZN(n12229) );
  NAND2_X1 U8847 ( .A1(n13838), .A2(n14012), .ZN(n14717) );
  AOI21_X1 U8848 ( .B1(n14012), .B2(n7301), .A(n14715), .ZN(n14716) );
  INV_X1 U8849 ( .A(n13837), .ZN(n7301) );
  NAND2_X1 U8850 ( .A1(n13886), .A2(n13885), .ZN(n13971) );
  OAI21_X1 U8851 ( .B1(n11192), .B2(n6983), .A(n11191), .ZN(n11445) );
  INV_X1 U8852 ( .A(n11193), .ZN(n14809) );
  NAND2_X1 U8853 ( .A1(n13980), .A2(n13979), .ZN(n13978) );
  AND2_X1 U8854 ( .A1(n7342), .A2(n6491), .ZN(n13814) );
  NAND2_X1 U8855 ( .A1(n7342), .A2(n7343), .ZN(n12230) );
  NAND2_X1 U8856 ( .A1(n11922), .A2(n7001), .ZN(n11923) );
  NAND2_X1 U8857 ( .A1(n7303), .A2(n13849), .ZN(n13998) );
  NAND2_X1 U8858 ( .A1(n14730), .A2(n14729), .ZN(n7303) );
  NAND2_X1 U8859 ( .A1(n14014), .A2(n14013), .ZN(n14012) );
  INV_X1 U8860 ( .A(n14731), .ZN(n15206) );
  OR2_X1 U8861 ( .A1(n9835), .A2(n9848), .ZN(n9886) );
  OR2_X1 U8862 ( .A1(n9812), .A2(n10173), .ZN(n9337) );
  INV_X1 U8863 ( .A(n11054), .ZN(n14041) );
  AND2_X1 U8864 ( .A1(n7427), .A2(n7428), .ZN(n12343) );
  NAND2_X1 U8865 ( .A1(n12326), .A2(n12325), .ZN(n12327) );
  NAND2_X1 U8866 ( .A1(n7200), .A2(n14113), .ZN(n14340) );
  NAND2_X1 U8867 ( .A1(n14206), .A2(n12316), .ZN(n14189) );
  NAND2_X1 U8868 ( .A1(n7187), .A2(n7186), .ZN(n7562) );
  NAND2_X1 U8869 ( .A1(n7187), .A2(n7188), .ZN(n14226) );
  NAND2_X1 U8870 ( .A1(n14256), .A2(n12311), .ZN(n14243) );
  OAI21_X1 U8871 ( .B1(n6893), .B2(n6522), .A(n12335), .ZN(n14248) );
  NAND2_X1 U8872 ( .A1(n14290), .A2(n12332), .ZN(n14271) );
  NAND2_X1 U8873 ( .A1(n12306), .A2(n12305), .ZN(n14289) );
  NAND2_X1 U8874 ( .A1(n11756), .A2(n11755), .ZN(n11758) );
  OAI211_X1 U8875 ( .C1(n11118), .C2(n7178), .A(n11322), .B(n7173), .ZN(n11375) );
  OR2_X1 U8876 ( .A1(n7179), .A2(n7178), .ZN(n7173) );
  NAND2_X1 U8877 ( .A1(n7177), .A2(n7180), .ZN(n11323) );
  NAND2_X1 U8878 ( .A1(n11118), .A2(n7179), .ZN(n7177) );
  NAND2_X1 U8879 ( .A1(n11134), .A2(n11133), .ZN(n11321) );
  INV_X1 U8880 ( .A(n14307), .ZN(n14601) );
  OR2_X1 U8881 ( .A1(n14112), .A2(n14827), .ZN(n7202) );
  NAND2_X1 U8882 ( .A1(n9491), .A2(n9490), .ZN(n11767) );
  INV_X1 U8883 ( .A(n14089), .ZN(n14413) );
  NAND2_X1 U8884 ( .A1(n6649), .A2(n14842), .ZN(n7015) );
  AOI21_X1 U8885 ( .B1(n14327), .B2(n14828), .A(n14326), .ZN(n7014) );
  NAND2_X1 U8886 ( .A1(n6848), .A2(n6847), .ZN(n6846) );
  INV_X1 U8887 ( .A(n14342), .ZN(n6847) );
  NAND2_X1 U8888 ( .A1(n14343), .A2(n14842), .ZN(n6848) );
  INV_X1 U8889 ( .A(n13828), .ZN(n14447) );
  INV_X1 U8890 ( .A(n11767), .ZN(n11796) );
  NAND2_X2 U8891 ( .A1(n6813), .A2(n6810), .ZN(n14453) );
  NOR2_X1 U8892 ( .A1(n6812), .A2(n6811), .ZN(n6810) );
  NOR2_X1 U8893 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6811) );
  NOR2_X1 U8894 ( .A1(n9292), .A2(n9290), .ZN(n7016) );
  INV_X1 U8895 ( .A(n9993), .ZN(n14465) );
  INV_X1 U8896 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11902) );
  NAND2_X1 U8897 ( .A1(n9608), .A2(n6563), .ZN(n9326) );
  INV_X1 U8898 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11346) );
  INV_X1 U8899 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11171) );
  INV_X1 U8900 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10950) );
  XNOR2_X1 U8901 ( .A(n9576), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11476) );
  INV_X1 U8902 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10377) );
  INV_X1 U8903 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10224) );
  INV_X1 U8904 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10057) );
  INV_X1 U8905 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10003) );
  INV_X1 U8906 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9972) );
  INV_X1 U8907 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9965) );
  INV_X1 U8908 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9954) );
  NOR2_X1 U8909 ( .A1(n15406), .A2(n14529), .ZN(n14585) );
  INV_X1 U8910 ( .A(n6832), .ZN(n15395) );
  INV_X1 U8911 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6834) );
  XNOR2_X1 U8912 ( .A(n14531), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15394) );
  XNOR2_X1 U8913 ( .A(n6839), .B(n14534), .ZN(n15397) );
  NAND2_X1 U8914 ( .A1(n15397), .A2(n15396), .ZN(n6777) );
  XNOR2_X1 U8915 ( .A(n14541), .B(n14540), .ZN(n14590) );
  NOR2_X1 U8916 ( .A1(n14590), .A2(n14589), .ZN(n14588) );
  OR2_X1 U8917 ( .A1(n15400), .A2(n15401), .ZN(n6779) );
  OAI211_X1 U8918 ( .C1(n14591), .C2(n6783), .A(n6781), .B(n6780), .ZN(n14595)
         );
  NOR2_X1 U8919 ( .A1(n14595), .A2(n14596), .ZN(n14594) );
  INV_X1 U8920 ( .A(n14563), .ZN(n7112) );
  NAND2_X1 U8921 ( .A1(n14761), .A2(n14568), .ZN(n14765) );
  NAND2_X1 U8922 ( .A1(n14773), .A2(n14576), .ZN(n14636) );
  OAI21_X1 U8923 ( .B1(n14774), .B2(n14775), .A(n14575), .ZN(n14576) );
  AOI21_X1 U8924 ( .B1(n7225), .B2(P3_REG1_REG_5__SCAN_IN), .A(n10823), .ZN(
        n10827) );
  INV_X1 U8925 ( .A(n7221), .ZN(n11275) );
  INV_X1 U8926 ( .A(n7280), .ZN(n12734) );
  AOI21_X1 U8927 ( .B1(n6616), .B2(n12738), .A(n6659), .ZN(n12755) );
  INV_X1 U8928 ( .A(n6661), .ZN(n12801) );
  OAI21_X1 U8929 ( .B1(n12814), .B2(n6923), .A(n11289), .ZN(n6922) );
  INV_X1 U8930 ( .A(n8875), .ZN(n8876) );
  OAI21_X1 U8931 ( .B1(n12874), .B2(n13116), .A(n8874), .ZN(n8875) );
  NOR2_X1 U8932 ( .A1(n6520), .A2(n8862), .ZN(n8863) );
  NAND2_X1 U8933 ( .A1(n10446), .A2(n7750), .ZN(n10589) );
  NAND2_X1 U8934 ( .A1(n7169), .A2(n6637), .ZN(P2_U3495) );
  NAND2_X1 U8935 ( .A1(n13756), .A2(n15018), .ZN(n7169) );
  INV_X1 U8936 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n7168) );
  XNOR2_X1 U8937 ( .A(n6987), .B(n6986), .ZN(n13915) );
  NAND2_X1 U8938 ( .A1(n6844), .A2(n6546), .ZN(P1_U3356) );
  NAND2_X1 U8939 ( .A1(n6845), .A2(n14279), .ZN(n6844) );
  AOI21_X1 U8940 ( .B1(n7201), .B2(n7198), .A(n14843), .ZN(n7197) );
  NAND2_X1 U8941 ( .A1(n14756), .A2(n14755), .ZN(n14754) );
  NAND2_X1 U8942 ( .A1(n14597), .A2(n14558), .ZN(n14756) );
  INV_X1 U8943 ( .A(n14770), .ZN(n14769) );
  XNOR2_X1 U8944 ( .A(n14644), .B(n6643), .ZN(n7113) );
  AND2_X1 U8945 ( .A1(n12571), .A2(n8414), .ZN(n6488) );
  AND2_X1 U8946 ( .A1(n7355), .A2(n13211), .ZN(n6489) );
  NAND2_X1 U8947 ( .A1(n7515), .A2(n9606), .ZN(n6490) );
  AND2_X1 U8948 ( .A1(n7343), .A2(n7341), .ZN(n6491) );
  INV_X1 U8949 ( .A(n10501), .ZN(n10260) );
  INV_X1 U8950 ( .A(n11191), .ZN(n6985) );
  NAND2_X1 U8951 ( .A1(n10860), .A2(n9237), .ZN(n9918) );
  AND2_X2 U8952 ( .A1(n7059), .A2(n7058), .ZN(n7580) );
  INV_X1 U8953 ( .A(n13431), .ZN(n7165) );
  AND2_X1 U8954 ( .A1(n6835), .A2(n6633), .ZN(n6492) );
  XNOR2_X1 U8955 ( .A(n8048), .B(n7056), .ZN(n13265) );
  INV_X1 U8956 ( .A(n13446), .ZN(n13659) );
  OR2_X1 U8957 ( .A1(n13221), .A2(n13301), .ZN(n6494) );
  AND2_X1 U8958 ( .A1(n7009), .A2(n14745), .ZN(n6495) );
  INV_X2 U8959 ( .A(n9017), .ZN(n9214) );
  AND2_X1 U8960 ( .A1(n11514), .A2(n7121), .ZN(n6496) );
  OR2_X1 U8961 ( .A1(n13151), .A2(n12457), .ZN(n6497) );
  AND2_X1 U8962 ( .A1(n12708), .A2(n11624), .ZN(n6498) );
  NOR2_X1 U8963 ( .A1(n10826), .A2(n15181), .ZN(n6499) );
  AND2_X1 U8964 ( .A1(n12120), .A2(n7453), .ZN(n6500) );
  AND2_X1 U8965 ( .A1(n8534), .A2(n10902), .ZN(n6501) );
  OAI21_X1 U8966 ( .B1(n12866), .B2(n13117), .A(n12499), .ZN(n12522) );
  AND2_X1 U8967 ( .A1(n9975), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6502) );
  AND2_X1 U8968 ( .A1(n14558), .A2(n6785), .ZN(n6503) );
  AND2_X1 U8969 ( .A1(n7623), .A2(n6619), .ZN(n6504) );
  NAND2_X1 U8970 ( .A1(n13524), .A2(n7099), .ZN(n6505) );
  INV_X1 U8971 ( .A(n12267), .ZN(n7084) );
  INV_X1 U8972 ( .A(n13668), .ZN(n7097) );
  OAI21_X1 U8973 ( .B1(n7465), .B2(n12400), .A(n6553), .ZN(n12397) );
  INV_X1 U8974 ( .A(n14337), .ZN(n14118) );
  AND2_X1 U8975 ( .A1(n14193), .A2(n13919), .ZN(n6506) );
  INV_X1 U8976 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8269) );
  AND2_X1 U8977 ( .A1(n6906), .A2(n6618), .ZN(n6507) );
  NAND2_X1 U8978 ( .A1(n8913), .A2(n11655), .ZN(n6508) );
  INV_X1 U8979 ( .A(n9533), .ZN(n7478) );
  AND2_X1 U8980 ( .A1(n7004), .A2(n7003), .ZN(n6509) );
  XNOR2_X1 U8981 ( .A(n11957), .B(n11949), .ZN(n6959) );
  INV_X1 U8982 ( .A(n13555), .ZN(n13520) );
  AND4_X1 U8983 ( .A1(n8088), .A2(n8087), .A3(n8086), .A4(n8085), .ZN(n13555)
         );
  NOR2_X1 U8984 ( .A1(n11959), .A2(n14693), .ZN(n6510) );
  INV_X1 U8985 ( .A(n7688), .ZN(n7432) );
  AND2_X1 U8986 ( .A1(n6959), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n6511) );
  INV_X1 U8987 ( .A(n12200), .ZN(n7137) );
  NOR2_X1 U8988 ( .A1(n7291), .A2(n10838), .ZN(n6512) );
  NAND2_X2 U8989 ( .A1(n12279), .A2(n7728), .ZN(n7736) );
  NAND2_X1 U8990 ( .A1(n13787), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7714) );
  INV_X2 U8991 ( .A(n9354), .ZN(n9331) );
  XOR2_X1 U8992 ( .A(n13668), .B(n6809), .Z(n6513) );
  OR2_X1 U8993 ( .A1(n8760), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n6514) );
  INV_X4 U8994 ( .A(n9017), .ZN(n9168) );
  NAND2_X1 U8995 ( .A1(n12036), .A2(n8921), .ZN(n6516) );
  INV_X1 U8996 ( .A(n9833), .ZN(n11901) );
  INV_X1 U8997 ( .A(n7512), .ZN(n7511) );
  NOR2_X1 U8998 ( .A1(n11029), .A2(n11239), .ZN(n6517) );
  NAND3_X1 U8999 ( .A1(n8500), .A2(n7557), .A3(n7385), .ZN(n6518) );
  INV_X1 U9000 ( .A(n6718), .ZN(n10863) );
  NAND2_X1 U9001 ( .A1(n9238), .A2(n10920), .ZN(n6718) );
  INV_X1 U9002 ( .A(n12334), .ZN(n7509) );
  AND3_X1 U9003 ( .A1(n7371), .A2(n7370), .A3(n7369), .ZN(n6519) );
  NOR2_X1 U9004 ( .A1(n12874), .A2(n13162), .ZN(n6520) );
  OR2_X1 U9005 ( .A1(n11190), .A2(n11189), .ZN(n6521) );
  NOR2_X1 U9006 ( .A1(n14385), .A2(n14027), .ZN(n6522) );
  AND2_X1 U9007 ( .A1(n11816), .A2(n13302), .ZN(n6523) );
  INV_X1 U9008 ( .A(n13944), .ZN(n7319) );
  NAND2_X1 U9009 ( .A1(n8335), .A2(n8334), .ZN(n8352) );
  AND2_X1 U9010 ( .A1(n6904), .A2(n6665), .ZN(n6524) );
  AND2_X1 U9011 ( .A1(n13625), .A2(n13595), .ZN(n6525) );
  NAND2_X1 U9012 ( .A1(n7771), .A2(n7770), .ZN(n14984) );
  AND2_X1 U9013 ( .A1(n6939), .A2(n6940), .ZN(n6526) );
  NAND2_X1 U9014 ( .A1(n13536), .A2(n13520), .ZN(n6527) );
  OR2_X1 U9015 ( .A1(n12788), .A2(n6492), .ZN(n6528) );
  AND2_X1 U9016 ( .A1(n8802), .A2(n7471), .ZN(n6529) );
  AND2_X1 U9017 ( .A1(n13688), .A2(n13434), .ZN(n6530) );
  AND2_X1 U9018 ( .A1(n12399), .A2(n7464), .ZN(n6531) );
  AND2_X1 U9019 ( .A1(n10656), .A2(n7784), .ZN(n6532) );
  INV_X1 U9020 ( .A(n12502), .ZN(n6801) );
  AND2_X1 U9021 ( .A1(n14813), .A2(n11447), .ZN(n6533) );
  XNOR2_X1 U9022 ( .A(n12087), .B(n14029), .ZN(n11757) );
  INV_X1 U9023 ( .A(n11757), .ZN(n7323) );
  NAND2_X1 U9024 ( .A1(n7592), .A2(n7591), .ZN(n7823) );
  AND2_X1 U9025 ( .A1(n13090), .A2(n13004), .ZN(n6534) );
  INV_X1 U9026 ( .A(n14127), .ZN(n14123) );
  AND2_X1 U9027 ( .A1(n12680), .A2(n13117), .ZN(n6535) );
  NAND2_X1 U9028 ( .A1(n7446), .A2(n8938), .ZN(n12446) );
  AND2_X1 U9029 ( .A1(n15404), .A2(n15403), .ZN(n6536) );
  AND2_X1 U9030 ( .A1(n8146), .A2(n13287), .ZN(n6537) );
  NAND2_X1 U9031 ( .A1(n9340), .A2(n7327), .ZN(n9377) );
  INV_X1 U9032 ( .A(n12228), .ZN(n7344) );
  AND3_X1 U9033 ( .A1(n9900), .A2(n9289), .A3(n9288), .ZN(n6538) );
  INV_X1 U9034 ( .A(n15030), .ZN(n7284) );
  INV_X1 U9035 ( .A(n9672), .ZN(n7497) );
  NAND2_X1 U9036 ( .A1(n14130), .A2(n14143), .ZN(n6539) );
  OR2_X1 U9037 ( .A1(n9150), .A2(n9151), .ZN(n6540) );
  NAND2_X1 U9038 ( .A1(n9310), .A2(n9309), .ZN(n14721) );
  AND2_X1 U9039 ( .A1(n12918), .A2(n8686), .ZN(n6541) );
  AND2_X1 U9040 ( .A1(n13404), .A2(n13405), .ZN(n6542) );
  INV_X1 U9041 ( .A(n12087), .ZN(n11919) );
  NAND2_X1 U9042 ( .A1(n9532), .A2(n9531), .ZN(n12087) );
  AND2_X1 U9043 ( .A1(n11554), .A2(n13304), .ZN(n6543) );
  AND2_X1 U9044 ( .A1(n7428), .A2(n12342), .ZN(n6544) );
  AND2_X1 U9045 ( .A1(n13668), .A2(n14990), .ZN(n6545) );
  INV_X1 U9046 ( .A(n9473), .ZN(n7489) );
  AND2_X1 U9047 ( .A1(n6648), .A2(n12368), .ZN(n6546) );
  AND2_X1 U9048 ( .A1(n7523), .A2(n7522), .ZN(n6547) );
  OR2_X1 U9049 ( .A1(n9034), .A2(n9033), .ZN(n6548) );
  INV_X1 U9050 ( .A(n7979), .ZN(n7436) );
  XNOR2_X1 U9051 ( .A(n7612), .B(SI_15_), .ZN(n7979) );
  OR2_X1 U9052 ( .A1(n13939), .A2(n13937), .ZN(n6549) );
  AND2_X1 U9053 ( .A1(n8299), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n6550) );
  OR2_X1 U9054 ( .A1(n14544), .A2(n14543), .ZN(n6551) );
  AND2_X1 U9055 ( .A1(n14206), .A2(n7328), .ZN(n6552) );
  AND2_X1 U9056 ( .A1(n9566), .A2(n9565), .ZN(n14745) );
  AND2_X1 U9057 ( .A1(n12399), .A2(n7461), .ZN(n6553) );
  INV_X1 U9058 ( .A(n6972), .ZN(n6971) );
  NAND2_X1 U9059 ( .A1(n6975), .A2(n11611), .ZN(n6972) );
  NAND2_X1 U9060 ( .A1(n8840), .A2(n12889), .ZN(n6554) );
  AND2_X1 U9061 ( .A1(n12622), .A2(n12625), .ZN(n12983) );
  INV_X1 U9062 ( .A(n7012), .ZN(n14166) );
  INV_X1 U9063 ( .A(n13849), .ZN(n7306) );
  OR2_X1 U9064 ( .A1(n9160), .A2(n9159), .ZN(n6555) );
  AND2_X1 U9065 ( .A1(n7298), .A2(n7297), .ZN(n6556) );
  AND2_X1 U9066 ( .A1(n6801), .A2(n6827), .ZN(n6557) );
  OR2_X1 U9067 ( .A1(n6499), .A2(n6962), .ZN(n6558) );
  NAND2_X1 U9068 ( .A1(n13417), .A2(n9231), .ZN(n13454) );
  INV_X1 U9069 ( .A(n13454), .ZN(n6699) );
  OR2_X1 U9070 ( .A1(n14481), .A2(n14480), .ZN(n6559) );
  AND2_X1 U9071 ( .A1(n8924), .A2(n14647), .ZN(n6560) );
  AND2_X1 U9072 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n6561) );
  AND2_X1 U9073 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n6562) );
  AND2_X1 U9074 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6563) );
  NOR2_X1 U9075 ( .A1(n11437), .A2(n11401), .ZN(n6564) );
  NOR2_X1 U9076 ( .A1(n13625), .A2(n13396), .ZN(n6565) );
  NOR2_X1 U9077 ( .A1(n13727), .A2(n13423), .ZN(n6566) );
  NOR2_X1 U9078 ( .A1(n14437), .A2(n13956), .ZN(n6567) );
  XNOR2_X1 U9079 ( .A(n12952), .B(n12701), .ZN(n12953) );
  AND2_X1 U9080 ( .A1(n7663), .A2(n7664), .ZN(n6568) );
  AND2_X1 U9081 ( .A1(n6748), .A2(n6752), .ZN(n6569) );
  OR2_X1 U9082 ( .A1(n14482), .A2(n7116), .ZN(n6570) );
  AND2_X1 U9083 ( .A1(n10398), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6571) );
  AND2_X1 U9084 ( .A1(n12573), .A2(n12572), .ZN(n12569) );
  AND2_X1 U9085 ( .A1(n15073), .A2(n11317), .ZN(n6572) );
  AND2_X1 U9086 ( .A1(n12120), .A2(n7455), .ZN(n6573) );
  AND2_X1 U9087 ( .A1(n7644), .A2(n6764), .ZN(n6574) );
  INV_X1 U9088 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9313) );
  INV_X1 U9089 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9290) );
  NOR2_X1 U9090 ( .A1(n14755), .A2(n14559), .ZN(n6575) );
  INV_X1 U9091 ( .A(n7167), .ZN(n7166) );
  NOR2_X1 U9092 ( .A1(n13536), .A2(n13555), .ZN(n7167) );
  INV_X1 U9093 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7471) );
  AND2_X1 U9094 ( .A1(n12305), .A2(n9855), .ZN(n12330) );
  NAND2_X1 U9095 ( .A1(n13190), .A2(n6858), .ZN(n13191) );
  AND2_X1 U9096 ( .A1(n7519), .A2(n7518), .ZN(n6576) );
  AND2_X1 U9097 ( .A1(n7606), .A2(n9982), .ZN(n6577) );
  NOR2_X1 U9098 ( .A1(n13568), .A2(n13556), .ZN(n6578) );
  INV_X1 U9099 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9952) );
  AND2_X1 U9100 ( .A1(n8274), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6579) );
  NAND2_X1 U9101 ( .A1(n8050), .A2(n8049), .ZN(n6580) );
  AND2_X1 U9102 ( .A1(n13934), .A2(n13933), .ZN(n6581) );
  NAND2_X1 U9103 ( .A1(n14813), .A2(n14035), .ZN(n6582) );
  INV_X1 U9104 ( .A(n14549), .ZN(n6784) );
  INV_X1 U9105 ( .A(n7425), .ZN(n7424) );
  OAI21_X1 U9106 ( .B1(n7595), .B2(n7426), .A(n7597), .ZN(n7425) );
  NAND2_X1 U9107 ( .A1(n13967), .A2(n14130), .ZN(n6583) );
  INV_X1 U9108 ( .A(n12428), .ZN(n7464) );
  AND2_X1 U9109 ( .A1(n7564), .A2(n7501), .ZN(n6584) );
  AND2_X1 U9110 ( .A1(n12136), .A2(n9599), .ZN(n12095) );
  INV_X1 U9111 ( .A(n12095), .ZN(n7513) );
  NAND2_X1 U9112 ( .A1(n6938), .A2(n12380), .ZN(n6585) );
  OR2_X1 U9113 ( .A1(n13179), .A2(n7357), .ZN(n6586) );
  AND2_X1 U9114 ( .A1(n7079), .A2(n6513), .ZN(n6587) );
  INV_X1 U9115 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7545) );
  NAND2_X1 U9116 ( .A1(n7144), .A2(n11903), .ZN(n7143) );
  AND2_X1 U9117 ( .A1(n13495), .A2(n13438), .ZN(n6588) );
  AND3_X1 U9118 ( .A1(n6494), .A2(n12004), .A3(n11814), .ZN(n6589) );
  AND2_X1 U9119 ( .A1(n7266), .A2(n6527), .ZN(n6590) );
  AND2_X1 U9120 ( .A1(n7156), .A2(n7154), .ZN(n6591) );
  INV_X1 U9121 ( .A(n9027), .ZN(n7536) );
  AND2_X1 U9122 ( .A1(n6508), .A2(n11652), .ZN(n6592) );
  INV_X1 U9123 ( .A(n13856), .ZN(n7307) );
  NOR2_X1 U9124 ( .A1(n7304), .A2(n13856), .ZN(n6593) );
  INV_X1 U9125 ( .A(n12199), .ZN(n7138) );
  AND2_X1 U9126 ( .A1(n7166), .A2(n7160), .ZN(n6594) );
  AND2_X1 U9127 ( .A1(n13669), .A2(n6814), .ZN(n6595) );
  AND2_X1 U9128 ( .A1(n6919), .A2(n6918), .ZN(n6596) );
  AND2_X1 U9129 ( .A1(n7319), .A2(n7316), .ZN(n6597) );
  AND2_X1 U9130 ( .A1(n8737), .A2(n8722), .ZN(n6598) );
  AND2_X1 U9131 ( .A1(n7013), .A2(n7014), .ZN(n6599) );
  OR2_X1 U9132 ( .A1(n9134), .A2(n9135), .ZN(n6600) );
  AND2_X1 U9133 ( .A1(n7283), .A2(n7282), .ZN(n6601) );
  OR2_X1 U9134 ( .A1(n9060), .A2(n9062), .ZN(n6602) );
  AND2_X1 U9135 ( .A1(n9291), .A2(n7502), .ZN(n6603) );
  AND2_X1 U9136 ( .A1(n6946), .A2(n6945), .ZN(n6604) );
  OR2_X1 U9137 ( .A1(n9061), .A2(n7537), .ZN(n6605) );
  NAND2_X1 U9138 ( .A1(n9134), .A2(n9135), .ZN(n6606) );
  NAND2_X1 U9139 ( .A1(n9772), .A2(n7481), .ZN(n6607) );
  NAND2_X1 U9140 ( .A1(n9703), .A2(n7487), .ZN(n6608) );
  NAND2_X1 U9141 ( .A1(n9534), .A2(n7478), .ZN(n6609) );
  NOR2_X1 U9142 ( .A1(n13416), .A2(n13484), .ZN(n6610) );
  AND2_X1 U9143 ( .A1(n8051), .A2(n7356), .ZN(n6611) );
  NAND2_X1 U9144 ( .A1(n7514), .A2(n9605), .ZN(n6612) );
  AND2_X1 U9145 ( .A1(n6539), .A2(n14100), .ZN(n7429) );
  INV_X1 U9146 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7502) );
  OR2_X1 U9147 ( .A1(n12464), .A2(n12921), .ZN(n6613) );
  NAND2_X1 U9148 ( .A1(n9739), .A2(n7484), .ZN(n6614) );
  INV_X1 U9149 ( .A(n7397), .ZN(n7396) );
  NAND2_X1 U9150 ( .A1(n12606), .A2(n7398), .ZN(n7397) );
  INV_X1 U9151 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6764) );
  INV_X1 U9152 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8274) );
  INV_X1 U9153 ( .A(n11949), .ZN(n7231) );
  INV_X1 U9154 ( .A(n13568), .ZN(n7107) );
  INV_X1 U9155 ( .A(n14207), .ZN(n6771) );
  XNOR2_X1 U9156 ( .A(n8355), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10400) );
  INV_X1 U9157 ( .A(n10400), .ZN(n6961) );
  XNOR2_X1 U9158 ( .A(n8419), .B(P3_IR_REG_9__SCAN_IN), .ZN(n15053) );
  INV_X1 U9159 ( .A(n15053), .ZN(n6905) );
  INV_X1 U9160 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7406) );
  INV_X1 U9161 ( .A(n13485), .ZN(n6840) );
  NAND2_X1 U9162 ( .A1(n13272), .A2(n6867), .ZN(n13264) );
  AND2_X1 U9163 ( .A1(n11922), .A2(n6999), .ZN(n6615) );
  INV_X1 U9164 ( .A(n12333), .ZN(n6819) );
  AND2_X1 U9165 ( .A1(n7280), .A2(n7279), .ZN(n6616) );
  NAND2_X1 U9166 ( .A1(n14294), .A2(n7006), .ZN(n6617) );
  AND4_X1 U9167 ( .A1(n8492), .A2(n8491), .A3(n8490), .A4(n8489), .ZN(n8921)
         );
  NAND2_X1 U9168 ( .A1(n8546), .A2(n6948), .ZN(n8581) );
  OR2_X1 U9169 ( .A1(n7282), .A2(n15053), .ZN(n6618) );
  AND2_X1 U9170 ( .A1(n7413), .A2(n7627), .ZN(n6619) );
  INV_X1 U9171 ( .A(n7108), .ZN(n13581) );
  NOR2_X1 U9172 ( .A1(n13601), .A2(n13710), .ZN(n7108) );
  AND4_X1 U9173 ( .A1(n8189), .A2(n8188), .A3(n8187), .A4(n8186), .ZN(n13444)
         );
  AND2_X1 U9174 ( .A1(n7284), .A2(n6905), .ZN(n6620) );
  OR2_X1 U9175 ( .A1(n14651), .A2(n8921), .ZN(n6621) );
  INV_X1 U9176 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7116) );
  INV_X1 U9177 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n6898) );
  INV_X1 U9178 ( .A(SI_8_), .ZN(n7426) );
  INV_X1 U9179 ( .A(n11290), .ZN(n6917) );
  INV_X1 U9180 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9946) );
  INV_X1 U9181 ( .A(n7294), .ZN(n6918) );
  AND2_X1 U9182 ( .A1(n11842), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7294) );
  INV_X1 U9183 ( .A(SI_14_), .ZN(n10129) );
  INV_X1 U9184 ( .A(n8840), .ZN(n13056) );
  NAND2_X1 U9185 ( .A1(n8744), .A2(n8743), .ZN(n8840) );
  INV_X1 U9186 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10615) );
  NOR2_X1 U9187 ( .A1(n8008), .A2(n10518), .ZN(n6622) );
  INV_X1 U9188 ( .A(n7678), .ZN(n7412) );
  NOR2_X1 U9189 ( .A1(n6918), .A2(n7231), .ZN(n6916) );
  NOR2_X1 U9190 ( .A1(n6908), .A2(n6905), .ZN(n6907) );
  OR2_X1 U9191 ( .A1(n14424), .A2(n14409), .ZN(n6623) );
  OR2_X1 U9192 ( .A1(n14976), .A2(n6863), .ZN(n6624) );
  AND2_X1 U9193 ( .A1(n7627), .A2(n7626), .ZN(n7678) );
  AND2_X1 U9194 ( .A1(n11818), .A2(n11817), .ZN(n6625) );
  AND2_X1 U9195 ( .A1(n7354), .A2(n7355), .ZN(n6626) );
  AND3_X1 U9196 ( .A1(n6976), .A2(n11111), .A3(n11110), .ZN(n11192) );
  NAND2_X1 U9197 ( .A1(n9578), .A2(n9577), .ZN(n13820) );
  INV_X1 U9198 ( .A(n13820), .ZN(n7008) );
  AND2_X1 U9199 ( .A1(n11117), .A2(n11121), .ZN(n7179) );
  INV_X1 U9200 ( .A(n11668), .ZN(n6837) );
  NAND2_X1 U9201 ( .A1(n7681), .A2(n7680), .ZN(n13603) );
  INV_X1 U9202 ( .A(n13603), .ZN(n7109) );
  NAND2_X1 U9203 ( .A1(n9636), .A2(n9635), .ZN(n14237) );
  INV_X1 U9204 ( .A(n14237), .ZN(n7003) );
  NAND2_X1 U9205 ( .A1(n7444), .A2(n8813), .ZN(n8815) );
  INV_X1 U9206 ( .A(n11121), .ZN(n11131) );
  AND2_X1 U9207 ( .A1(n11750), .A2(n7009), .ZN(n6627) );
  INV_X1 U9208 ( .A(n11964), .ZN(n12726) );
  OR2_X1 U9209 ( .A1(n11467), .A2(n11466), .ZN(n6628) );
  AND2_X1 U9210 ( .A1(n12048), .A2(n12047), .ZN(n6629) );
  NAND2_X1 U9211 ( .A1(n6664), .A2(n6917), .ZN(n6919) );
  OR2_X1 U9212 ( .A1(n11632), .A2(n11638), .ZN(n11756) );
  AND2_X1 U9213 ( .A1(n6494), .A2(n11814), .ZN(n6630) );
  NOR2_X1 U9214 ( .A1(n11822), .A2(n13221), .ZN(n7103) );
  OR2_X1 U9215 ( .A1(n11192), .A2(n6984), .ZN(n6631) );
  AND2_X1 U9216 ( .A1(n14843), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6632) );
  INV_X1 U9217 ( .A(n6756), .ZN(n11227) );
  NAND2_X1 U9218 ( .A1(n11219), .A2(n11222), .ZN(n6756) );
  NAND2_X1 U9219 ( .A1(n12766), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n6633) );
  OR2_X1 U9220 ( .A1(n11964), .A2(n14688), .ZN(n6634) );
  INV_X1 U9221 ( .A(n11071), .ZN(n7105) );
  NAND2_X1 U9222 ( .A1(n10393), .A2(n10400), .ZN(n7225) );
  AND2_X1 U9223 ( .A1(n12766), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n6635) );
  INV_X1 U9224 ( .A(n12712), .ZN(n15096) );
  NAND2_X1 U9225 ( .A1(n11118), .A2(n11117), .ZN(n11132) );
  NOR2_X1 U9226 ( .A1(n10393), .A2(n10400), .ZN(n10823) );
  INV_X1 U9227 ( .A(n10823), .ZN(n7223) );
  AND2_X1 U9228 ( .A1(n8922), .A2(n8921), .ZN(n6636) );
  OR2_X1 U9229 ( .A1(n15018), .A2(n7168), .ZN(n6637) );
  OR2_X1 U9230 ( .A1(n13797), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U9231 ( .A1(n8842), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6639) );
  OR2_X1 U9232 ( .A1(n10838), .A2(n7292), .ZN(n6640) );
  AND2_X1 U9233 ( .A1(n7221), .A2(n7220), .ZN(n6641) );
  AND2_X1 U9234 ( .A1(n12805), .A2(n6921), .ZN(n6642) );
  INV_X1 U9235 ( .A(n13311), .ZN(n6836) );
  XOR2_X1 U9236 ( .A(n7565), .B(P3_ADDR_REG_19__SCAN_IN), .Z(n6643) );
  INV_X1 U9237 ( .A(SI_23_), .ZN(n7405) );
  NAND2_X1 U9238 ( .A1(n10547), .A2(n10568), .ZN(n6644) );
  AND2_X1 U9239 ( .A1(n9994), .A2(n10539), .ZN(n10568) );
  XNOR2_X1 U9240 ( .A(n11283), .B(n11292), .ZN(n11029) );
  XNOR2_X1 U9241 ( .A(n12813), .B(n12831), .ZN(n12803) );
  NOR2_X1 U9242 ( .A1(n12831), .A2(n12830), .ZN(n12833) );
  XNOR2_X1 U9243 ( .A(n12830), .B(n12831), .ZN(n12800) );
  OAI21_X1 U9244 ( .B1(n10985), .B2(n10984), .A(n10983), .ZN(n6650) );
  NOR2_X1 U9245 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n6653) );
  OAI211_X2 U9246 ( .C1(P1_IR_REG_31__SCAN_IN), .C2(P1_IR_REG_28__SCAN_IN), 
        .A(n9295), .B(n6654), .ZN(n14456) );
  INV_X1 U9247 ( .A(n12094), .ZN(n6655) );
  NAND2_X1 U9248 ( .A1(n6656), .A2(n7172), .ZN(n11584) );
  NAND2_X1 U9249 ( .A1(n6656), .A2(n11379), .ZN(n11582) );
  NAND2_X1 U9250 ( .A1(n11531), .A2(n11378), .ZN(n6656) );
  NAND2_X1 U9251 ( .A1(n6657), .A2(n12338), .ZN(n14158) );
  OAI21_X1 U9252 ( .B1(n7550), .B2(n12337), .A(n6657), .ZN(n14360) );
  NAND3_X1 U9253 ( .A1(n14146), .A2(n12340), .A3(n7429), .ZN(n7427) );
  OAI211_X2 U9254 ( .C1(n9572), .C2(n9947), .A(n9362), .B(n6658), .ZN(n11053)
         );
  NOR2_X1 U9255 ( .A1(n12775), .A2(n12776), .ZN(n12779) );
  INV_X1 U9256 ( .A(n11291), .ZN(n6664) );
  NAND3_X1 U9257 ( .A1(n6666), .A2(n10260), .A3(n7289), .ZN(n6665) );
  NAND4_X1 U9258 ( .A1(n7659), .A2(n7644), .A3(n7545), .A4(n7558), .ZN(n6671)
         );
  NAND2_X1 U9259 ( .A1(n6821), .A2(n9156), .ZN(n6674) );
  NAND3_X1 U9260 ( .A1(n6679), .A2(n6678), .A3(n6677), .ZN(n6681) );
  NAND2_X1 U9261 ( .A1(n6680), .A2(n9271), .ZN(P2_U3328) );
  NAND2_X1 U9262 ( .A1(n6681), .A2(n9268), .ZN(n6680) );
  NAND2_X1 U9263 ( .A1(n6685), .A2(n6602), .ZN(n9068) );
  NAND3_X1 U9264 ( .A1(n9057), .A2(n6605), .A3(n9056), .ZN(n6685) );
  NAND2_X1 U9265 ( .A1(n9021), .A2(n9020), .ZN(n6689) );
  NAND2_X1 U9266 ( .A1(n6823), .A2(n6822), .ZN(n6690) );
  NAND2_X1 U9267 ( .A1(n6866), .A2(n6865), .ZN(n6691) );
  OAI211_X1 U9268 ( .C1(n9139), .C2(n6695), .A(n6692), .B(n7542), .ZN(n7541)
         );
  NAND2_X1 U9269 ( .A1(n6694), .A2(n6693), .ZN(n6692) );
  INV_X1 U9270 ( .A(n9138), .ZN(n6693) );
  NAND2_X1 U9271 ( .A1(n6695), .A2(n9139), .ZN(n6694) );
  NAND2_X1 U9272 ( .A1(n7538), .A2(n6600), .ZN(n6695) );
  OAI211_X2 U9273 ( .C1(n7962), .C2(n9947), .A(n7710), .B(n7104), .ZN(n7233)
         );
  XNOR2_X1 U9274 ( .A(n10965), .B(n6696), .ZN(n11003) );
  NAND2_X1 U9275 ( .A1(n10963), .A2(n10962), .ZN(n6710) );
  NAND2_X2 U9276 ( .A1(n13501), .A2(n13435), .ZN(n13482) );
  INV_X1 U9277 ( .A(n8201), .ZN(n6704) );
  NOR2_X4 U9278 ( .A1(n6701), .A2(n6700), .ZN(n7644) );
  NAND3_X1 U9279 ( .A1(n7656), .A2(n7640), .A3(n6713), .ZN(n6701) );
  NAND3_X1 U9280 ( .A1(n6712), .A2(n6711), .A3(n6713), .ZN(n7652) );
  NAND3_X1 U9281 ( .A1(n7644), .A2(n7659), .A3(n6703), .ZN(n6702) );
  AND3_X4 U9282 ( .A1(n7768), .A2(n6706), .A3(n6705), .ZN(n7659) );
  AOI21_X2 U9283 ( .B1(n13593), .B2(n13427), .A(n13426), .ZN(n13575) );
  OR2_X2 U9284 ( .A1(n12013), .A2(n12012), .ZN(n12165) );
  OAI21_X1 U9285 ( .B1(n11003), .B2(n6710), .A(n11002), .ZN(n11004) );
  NOR2_X2 U9286 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n6711) );
  NAND2_X1 U9287 ( .A1(n8884), .A2(n6714), .ZN(n15093) );
  NAND2_X1 U9288 ( .A1(n11074), .A2(n11149), .ZN(n11158) );
  NAND2_X1 U9289 ( .A1(n12886), .A2(n8738), .ZN(n8764) );
  INV_X1 U9290 ( .A(n10915), .ZN(n14978) );
  NAND2_X1 U9291 ( .A1(n6836), .A2(n10915), .ZN(n10920) );
  NAND2_X1 U9292 ( .A1(n14645), .A2(n7211), .ZN(n6719) );
  NAND2_X1 U9293 ( .A1(n14656), .A2(n8783), .ZN(n6720) );
  NAND3_X1 U9294 ( .A1(n7261), .A2(n7262), .A3(n7260), .ZN(n13501) );
  INV_X1 U9295 ( .A(n7962), .ZN(n7753) );
  NAND2_X1 U9296 ( .A1(n11232), .A2(n11231), .ZN(n11230) );
  AND3_X2 U9297 ( .A1(n6519), .A2(n8320), .A3(n8262), .ZN(n8500) );
  NAND3_X1 U9298 ( .A1(n7557), .A2(n6722), .A3(n7384), .ZN(n8282) );
  AND4_X2 U9299 ( .A1(n6519), .A2(n8320), .A3(n8281), .A4(n8262), .ZN(n6722)
         );
  OAI21_X2 U9300 ( .B1(n13032), .B2(n6806), .A(n6804), .ZN(n12972) );
  INV_X1 U9301 ( .A(n12845), .ZN(n6728) );
  NAND2_X1 U9302 ( .A1(n6734), .A2(n10416), .ZN(n10228) );
  XNOR2_X1 U9303 ( .A(n11278), .B(n15053), .ZN(n15059) );
  NOR2_X2 U9304 ( .A1(n15038), .A2(n6739), .ZN(n11278) );
  XNOR2_X1 U9305 ( .A(n11274), .B(n11292), .ZN(n11017) );
  XNOR2_X1 U9306 ( .A(n10259), .B(n10258), .ZN(n10471) );
  NAND3_X1 U9307 ( .A1(n8500), .A2(n7384), .A3(n7557), .ZN(n6747) );
  NAND2_X1 U9308 ( .A1(n6749), .A2(n6748), .ZN(n6755) );
  NAND2_X1 U9309 ( .A1(n6569), .A2(n6749), .ZN(n6751) );
  NAND2_X1 U9310 ( .A1(n6587), .A2(n7081), .ZN(n6748) );
  INV_X1 U9311 ( .A(n6750), .ZN(n6749) );
  NAND2_X1 U9312 ( .A1(n6753), .A2(n6751), .ZN(P2_U3192) );
  INV_X1 U9313 ( .A(n8258), .ZN(n6752) );
  AOI21_X1 U9314 ( .B1(n6755), .B2(n8234), .A(n6754), .ZN(n6753) );
  INV_X1 U9315 ( .A(n8257), .ZN(n6754) );
  NAND2_X1 U9316 ( .A1(n11261), .A2(n7367), .ZN(n11500) );
  OAI21_X2 U9317 ( .B1(n7547), .B2(n6763), .A(n6761), .ZN(n12266) );
  XNOR2_X2 U9318 ( .A(n6765), .B(n7655), .ZN(n9923) );
  NAND2_X1 U9319 ( .A1(n7368), .A2(n10669), .ZN(n10876) );
  NAND2_X1 U9320 ( .A1(n10427), .A2(n10426), .ZN(n10435) );
  AND2_X1 U9321 ( .A1(n10419), .A2(n7732), .ZN(n10427) );
  NAND2_X1 U9322 ( .A1(n6769), .A2(n6768), .ZN(n10991) );
  OR2_X1 U9323 ( .A1(n10990), .A2(n10989), .ZN(n6768) );
  NAND2_X1 U9324 ( .A1(n10990), .A2(n10989), .ZN(n6769) );
  OAI21_X1 U9325 ( .B1(n15396), .B2(n15397), .A(n6777), .ZN(SUB_1596_U58) );
  INV_X1 U9326 ( .A(n6779), .ZN(n15399) );
  INV_X1 U9327 ( .A(n6778), .ZN(n14548) );
  XNOR2_X1 U9328 ( .A(n14544), .B(n14543), .ZN(n15400) );
  NAND2_X1 U9329 ( .A1(n6784), .A2(n14553), .ZN(n6780) );
  NAND2_X1 U9330 ( .A1(n14591), .A2(n6782), .ZN(n6781) );
  NOR2_X1 U9331 ( .A1(n6784), .A2(n14553), .ZN(n6782) );
  INV_X1 U9332 ( .A(n14553), .ZN(n6783) );
  NAND2_X1 U9333 ( .A1(n14591), .A2(n14549), .ZN(n14552) );
  NAND2_X1 U9334 ( .A1(n14598), .A2(n15332), .ZN(n14597) );
  NAND2_X1 U9335 ( .A1(n6786), .A2(n7575), .ZN(n7752) );
  NAND2_X1 U9336 ( .A1(n6790), .A2(n7741), .ZN(n6786) );
  OAI211_X1 U9337 ( .C1(n6790), .C2(n6789), .A(n7576), .B(n6787), .ZN(n7579)
         );
  NAND2_X1 U9338 ( .A1(n6788), .A2(n7575), .ZN(n6787) );
  INV_X1 U9339 ( .A(n7741), .ZN(n6788) );
  INV_X1 U9340 ( .A(n7575), .ZN(n6789) );
  NAND2_X2 U9341 ( .A1(n6793), .A2(n7421), .ZN(n7864) );
  NAND3_X1 U9342 ( .A1(n7435), .A2(n7089), .A3(n6795), .ZN(n7088) );
  NAND2_X2 U9343 ( .A1(n6796), .A2(SI_14_), .ZN(n6795) );
  NAND3_X1 U9344 ( .A1(n7435), .A2(n7436), .A3(n6795), .ZN(n7094) );
  NAND2_X1 U9345 ( .A1(n7611), .A2(n6795), .ZN(n7959) );
  NAND2_X1 U9346 ( .A1(n7435), .A2(n6795), .ZN(n7980) );
  NAND2_X1 U9347 ( .A1(n7437), .A2(n6795), .ZN(n7961) );
  INV_X1 U9348 ( .A(n7610), .ZN(n6796) );
  NAND2_X1 U9349 ( .A1(n7111), .A2(n14764), .ZN(n6798) );
  NAND3_X1 U9350 ( .A1(n7111), .A2(n14572), .A3(n14764), .ZN(n14771) );
  NAND2_X1 U9351 ( .A1(n14771), .A2(n14772), .ZN(n14768) );
  NAND2_X1 U9352 ( .A1(n15093), .A2(n15092), .ZN(n7215) );
  NAND2_X1 U9353 ( .A1(n12536), .A2(n12541), .ZN(n15092) );
  NAND2_X1 U9354 ( .A1(n10895), .A2(n8325), .ZN(n10937) );
  NAND3_X1 U9355 ( .A1(n7215), .A2(n8312), .A3(n7216), .ZN(n10895) );
  NAND2_X1 U9356 ( .A1(n10937), .A2(n12547), .ZN(n10936) );
  AOI21_X2 U9357 ( .B1(n7620), .B2(n7619), .A(n6622), .ZN(n7621) );
  NAND2_X1 U9358 ( .A1(n7094), .A2(n7614), .ZN(n7997) );
  NAND2_X1 U9359 ( .A1(n7609), .A2(n7608), .ZN(n7610) );
  XNOR2_X1 U9360 ( .A(n9256), .B(n12284), .ZN(n6869) );
  NAND2_X1 U9361 ( .A1(n10936), .A2(n8343), .ZN(n15071) );
  NAND2_X1 U9362 ( .A1(n12903), .A2(n6613), .ZN(n7207) );
  NAND2_X1 U9363 ( .A1(n6815), .A2(n7353), .ZN(n8072) );
  NOR2_X1 U9364 ( .A1(n8302), .A2(n7549), .ZN(n7205) );
  NAND2_X1 U9365 ( .A1(n7206), .A2(n7203), .ZN(n12541) );
  INV_X1 U9366 ( .A(n8302), .ZN(n6838) );
  INV_X1 U9367 ( .A(n12294), .ZN(n8275) );
  NOR2_X2 U9368 ( .A1(n12294), .A2(n13176), .ZN(n8534) );
  NAND2_X1 U9369 ( .A1(n8300), .A2(n8301), .ZN(n8302) );
  NAND2_X1 U9370 ( .A1(n7207), .A2(n6598), .ZN(n12886) );
  NAND2_X1 U9372 ( .A1(n12110), .A2(n12109), .ZN(n12108) );
  NAND2_X2 U9373 ( .A1(n9298), .A2(n9299), .ZN(n9354) );
  NOR2_X1 U9374 ( .A1(n14341), .A2(n6846), .ZN(n14421) );
  OAI21_X1 U9375 ( .B1(n7864), .B2(n7862), .A(n7599), .ZN(n7884) );
  INV_X1 U9376 ( .A(n13538), .ZN(n7264) );
  NOR2_X1 U9377 ( .A1(n7204), .A2(n7549), .ZN(n7203) );
  NAND2_X1 U9378 ( .A1(n12127), .A2(n8520), .ZN(n12126) );
  INV_X1 U9379 ( .A(n15071), .ZN(n8359) );
  NAND2_X1 U9380 ( .A1(n8942), .A2(n8941), .ZN(n12429) );
  NAND2_X1 U9381 ( .A1(n6924), .A2(n6925), .ZN(n12388) );
  INV_X1 U9383 ( .A(n8759), .ZN(n7470) );
  NOR2_X1 U9384 ( .A1(n13660), .A2(n7553), .ZN(n13661) );
  NAND2_X1 U9385 ( .A1(n12466), .A2(n8955), .ZN(n9273) );
  OAI211_X1 U9386 ( .C1(n10688), .C2(n7473), .A(n10906), .B(n6942), .ZN(n6941)
         );
  OAI21_X2 U9387 ( .B1(n11878), .B2(n8918), .A(n11879), .ZN(n11892) );
  AOI21_X2 U9388 ( .B1(n12424), .B2(n8927), .A(n12408), .ZN(n12421) );
  NAND2_X1 U9389 ( .A1(n10878), .A2(n7842), .ZN(n11220) );
  NAND2_X1 U9390 ( .A1(n13264), .A2(n6489), .ZN(n6815) );
  NAND3_X1 U9391 ( .A1(n7408), .A2(n7407), .A3(n7406), .ZN(n6816) );
  OAI21_X1 U9392 ( .B1(n14205), .B2(n14207), .A(n6820), .ZN(n14192) );
  AND2_X1 U9393 ( .A1(n8999), .A2(n8998), .ZN(n6873) );
  NAND2_X1 U9394 ( .A1(n9155), .A2(n9154), .ZN(n6821) );
  INV_X1 U9395 ( .A(n9016), .ZN(n6823) );
  NAND2_X1 U9396 ( .A1(n9074), .A2(n9075), .ZN(n9073) );
  NAND2_X1 U9397 ( .A1(n6861), .A2(n6862), .ZN(n9074) );
  MUX2_X1 U9398 ( .A(n10145), .B(n13808), .S(n10069), .Z(n8994) );
  NAND2_X1 U9399 ( .A1(n8317), .A2(n8316), .ZN(n6825) );
  NAND3_X1 U9400 ( .A1(n12670), .A2(n12890), .A3(n12519), .ZN(n6828) );
  INV_X1 U9401 ( .A(n12522), .ZN(n6829) );
  NAND2_X2 U9402 ( .A1(n7034), .A2(n7037), .ZN(n8387) );
  NAND2_X2 U9403 ( .A1(n8387), .A2(n8386), .ZN(n8389) );
  XNOR2_X1 U9404 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8305) );
  NAND2_X1 U9405 ( .A1(n8276), .A2(n12294), .ZN(n8476) );
  INV_X1 U9406 ( .A(n8843), .ZN(n7026) );
  NAND2_X1 U9407 ( .A1(n8416), .A2(n8415), .ZN(n8441) );
  NAND2_X1 U9408 ( .A1(n7053), .A2(n7052), .ZN(n8741) );
  INV_X1 U9409 ( .A(n6833), .ZN(n15402) );
  OAI21_X1 U9410 ( .B1(n6536), .B2(n6834), .A(n6833), .ZN(n6832) );
  XNOR2_X1 U9411 ( .A(n14557), .B(n14556), .ZN(n14598) );
  NOR2_X1 U9412 ( .A1(n15059), .A2(n15188), .ZN(n15058) );
  INV_X1 U9413 ( .A(n6891), .ZN(n6900) );
  INV_X1 U9414 ( .A(n6892), .ZN(n12863) );
  OAI21_X1 U9415 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n14530), .A(n14584), .ZN(
        n15403) );
  INV_X1 U9416 ( .A(n14535), .ZN(n6839) );
  NAND2_X1 U9417 ( .A1(n11073), .A2(n11072), .ZN(n11074) );
  NAND2_X1 U9418 ( .A1(n12020), .A2(n12019), .ZN(n12172) );
  NAND2_X1 U9419 ( .A1(n6838), .A2(n8892), .ZN(n7204) );
  INV_X1 U9420 ( .A(n7103), .ZN(n11910) );
  NAND2_X1 U9422 ( .A1(n10852), .A2(n10851), .ZN(n10988) );
  AND2_X4 U9423 ( .A1(n12265), .A2(n9298), .ZN(n9409) );
  NAND2_X1 U9424 ( .A1(n6841), .A2(n8306), .ZN(n8317) );
  NAND2_X1 U9425 ( .A1(n8304), .A2(n8305), .ZN(n6841) );
  NAND2_X1 U9426 ( .A1(n8542), .A2(n8541), .ZN(n8544) );
  OR2_X1 U9427 ( .A1(n12674), .A2(n6842), .ZN(n12677) );
  OAI21_X1 U9428 ( .B1(n13662), .B2(n14994), .A(n13661), .ZN(n13663) );
  INV_X1 U9429 ( .A(n13478), .ZN(n7149) );
  OAI21_X1 U9430 ( .B1(n8152), .B2(n11798), .A(n8151), .ZN(n8154) );
  NAND2_X1 U9431 ( .A1(n7324), .A2(n7322), .ZN(n12081) );
  NAND2_X1 U9432 ( .A1(n14161), .A2(n14162), .ZN(n14160) );
  NAND2_X1 U9433 ( .A1(n8806), .A2(n8805), .ZN(n8808) );
  NAND2_X1 U9434 ( .A1(n7470), .A2(n7469), .ZN(n8804) );
  NAND2_X1 U9435 ( .A1(n7440), .A2(n8891), .ZN(n10728) );
  NAND2_X1 U9436 ( .A1(n8944), .A2(n12962), .ZN(n12373) );
  NAND2_X1 U9437 ( .A1(n7450), .A2(n7447), .ZN(n12153) );
  NAND2_X1 U9438 ( .A1(n7444), .A2(n7442), .ZN(n7445) );
  NAND2_X1 U9439 ( .A1(n7468), .A2(n7466), .ZN(n11205) );
  NAND2_X1 U9440 ( .A1(n7477), .A2(n6592), .ZN(n11651) );
  NAND2_X1 U9441 ( .A1(n6941), .A2(n8904), .ZN(n11088) );
  NAND2_X1 U9442 ( .A1(n11205), .A2(n8908), .ZN(n11359) );
  NAND2_X1 U9443 ( .A1(n11357), .A2(n7475), .ZN(n7477) );
  NAND2_X1 U9444 ( .A1(n10816), .A2(n8899), .ZN(n7472) );
  NAND2_X1 U9445 ( .A1(n7472), .A2(n8902), .ZN(n6942) );
  NAND2_X1 U9446 ( .A1(n12153), .A2(n6944), .ZN(n12409) );
  NAND2_X1 U9447 ( .A1(n8811), .A2(n11696), .ZN(n7444) );
  NAND2_X1 U9448 ( .A1(n7196), .A2(n7201), .ZN(n14420) );
  AOI22_X2 U9449 ( .A1(n12421), .A2(n8929), .B1(n12419), .B2(n13021), .ZN(
        n12455) );
  INV_X1 U9450 ( .A(n9633), .ZN(n6850) );
  NAND2_X1 U9451 ( .A1(n6850), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9343) );
  INV_X1 U9452 ( .A(n8268), .ZN(n7385) );
  NAND2_X1 U9453 ( .A1(n8270), .A2(n8269), .ZN(n8284) );
  NAND2_X1 U9454 ( .A1(n11377), .A2(n11376), .ZN(n11531) );
  OAI22_X1 U9455 ( .A1(n11041), .A2(n11048), .B1(n14040), .B2(n11053), .ZN(
        n10985) );
  INV_X1 U9456 ( .A(n7407), .ZN(n6855) );
  NAND2_X1 U9457 ( .A1(n7584), .A2(n7583), .ZN(n7785) );
  OAI21_X1 U9458 ( .B1(n7864), .B2(n7074), .A(n7072), .ZN(n7077) );
  NAND2_X1 U9459 ( .A1(n12081), .A2(n12080), .ZN(n12110) );
  NAND2_X1 U9460 ( .A1(n7498), .A2(n7495), .ZN(n6897) );
  XNOR2_X1 U9461 ( .A(n14562), .B(n7112), .ZN(n14760) );
  NAND2_X1 U9462 ( .A1(n14580), .A2(n14634), .ZN(n14638) );
  NAND2_X1 U9463 ( .A1(n14760), .A2(n14759), .ZN(n14758) );
  NAND2_X1 U9464 ( .A1(n14638), .A2(n14639), .ZN(n14640) );
  NAND2_X1 U9465 ( .A1(n14765), .A2(n14766), .ZN(n14764) );
  AOI21_X1 U9466 ( .B1(n6489), .B2(n13265), .A(n6611), .ZN(n7353) );
  AOI21_X1 U9467 ( .B1(n7083), .B2(n7085), .A(n7080), .ZN(n7079) );
  NAND2_X1 U9468 ( .A1(n8857), .A2(n8856), .ZN(n12871) );
  NAND2_X1 U9469 ( .A1(n14139), .A2(n12320), .ZN(n14124) );
  NAND2_X1 U9470 ( .A1(n7621), .A2(n7622), .ZN(n6860) );
  OAI21_X1 U9471 ( .B1(n13666), .B2(n14994), .A(n6595), .ZN(n13756) );
  INV_X1 U9472 ( .A(n9066), .ZN(n6862) );
  INV_X1 U9473 ( .A(n8235), .ZN(n6864) );
  NAND2_X2 U9474 ( .A1(n6864), .A2(n6863), .ZN(n10637) );
  AOI21_X1 U9475 ( .B1(n9068), .B2(n9067), .A(n9065), .ZN(n9066) );
  NAND2_X1 U9476 ( .A1(n9123), .A2(n9122), .ZN(n9129) );
  NAND2_X1 U9477 ( .A1(n9016), .A2(n9015), .ZN(n6866) );
  XNOR2_X1 U9478 ( .A(n10434), .B(n7734), .ZN(n10426) );
  INV_X1 U9479 ( .A(n9266), .ZN(n9261) );
  INV_X1 U9480 ( .A(n9044), .ZN(n6882) );
  NAND2_X1 U9481 ( .A1(n6868), .A2(n9005), .ZN(n9011) );
  NAND2_X1 U9482 ( .A1(n9006), .A2(n9007), .ZN(n6868) );
  NAND2_X1 U9483 ( .A1(n9230), .A2(n9229), .ZN(n9266) );
  NAND2_X1 U9484 ( .A1(n6881), .A2(n6880), .ZN(n9156) );
  NAND2_X1 U9485 ( .A1(n9213), .A2(n7233), .ZN(n8990) );
  INV_X1 U9486 ( .A(n8500), .ZN(n8473) );
  XNOR2_X2 U9487 ( .A(n8272), .B(n8271), .ZN(n12294) );
  NAND2_X1 U9488 ( .A1(n7115), .A2(n14640), .ZN(n7114) );
  XNOR2_X1 U9489 ( .A(n7114), .B(n7113), .ZN(SUB_1596_U4) );
  NAND3_X1 U9490 ( .A1(n14328), .A2(n7015), .A3(n6599), .ZN(n14418) );
  NAND2_X1 U9491 ( .A1(n14774), .A2(n14775), .ZN(n14773) );
  NAND2_X1 U9492 ( .A1(n7531), .A2(n7529), .ZN(n6881) );
  NAND2_X1 U9493 ( .A1(n7531), .A2(n7532), .ZN(n9155) );
  AND2_X1 U9494 ( .A1(n6873), .A2(n6872), .ZN(n9007) );
  NAND2_X1 U9495 ( .A1(n9000), .A2(n9001), .ZN(n6872) );
  OAI21_X1 U9496 ( .B1(n9129), .B2(n9128), .A(n9127), .ZN(n9131) );
  AOI21_X1 U9497 ( .B1(n9034), .B2(n9033), .A(n9032), .ZN(n6884) );
  NAND2_X2 U9498 ( .A1(n7611), .A2(n7438), .ZN(n7435) );
  XNOR2_X1 U9499 ( .A(n8076), .B(SI_22_), .ZN(n8079) );
  NAND2_X1 U9500 ( .A1(n8108), .A2(n8107), .ZN(n8112) );
  NAND2_X1 U9501 ( .A1(n7077), .A2(n7414), .ZN(n7939) );
  AOI21_X1 U9502 ( .B1(n7148), .B2(n7151), .A(n6610), .ZN(n7145) );
  NAND2_X1 U9503 ( .A1(n7146), .A2(n7145), .ZN(n13464) );
  NOR2_X1 U9504 ( .A1(n13414), .A2(n6588), .ZN(n7155) );
  NOR2_X1 U9505 ( .A1(n6550), .A2(n6501), .ZN(n6876) );
  NAND2_X1 U9506 ( .A1(n7997), .A2(n7996), .ZN(n7620) );
  INV_X1 U9507 ( .A(n7602), .ZN(n7420) );
  NAND2_X1 U9508 ( .A1(n7066), .A2(n7678), .ZN(n7065) );
  NAND2_X1 U9509 ( .A1(n14593), .A2(n14592), .ZN(n14591) );
  AOI22_X2 U9510 ( .A1(n9787), .A2(n9786), .B1(n9785), .B2(n9784), .ZN(n9890)
         );
  NAND2_X1 U9511 ( .A1(n7490), .A2(n7488), .ZN(n9472) );
  NAND2_X1 U9512 ( .A1(n6897), .A2(n7497), .ZN(n9673) );
  NAND2_X1 U9513 ( .A1(n6895), .A2(n6894), .ZN(n9549) );
  BUF_X4 U9514 ( .A(n9492), .Z(n9821) );
  NOR2_X1 U9515 ( .A1(n10637), .A2(n11983), .ZN(n9935) );
  INV_X2 U9516 ( .A(n8996), .ZN(n9213) );
  NAND2_X1 U9517 ( .A1(n6883), .A2(n6548), .ZN(n9039) );
  INV_X1 U9518 ( .A(n6884), .ZN(n6883) );
  NAND2_X1 U9519 ( .A1(n14345), .A2(n6623), .ZN(P1_U3554) );
  NAND3_X1 U9520 ( .A1(n7568), .A2(n7064), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7061) );
  INV_X1 U9521 ( .A(n7186), .ZN(n7185) );
  NAND2_X1 U9522 ( .A1(n8609), .A2(n8608), .ZN(n7051) );
  NAND2_X1 U9523 ( .A1(n8639), .A2(n8638), .ZN(n7044) );
  NAND2_X1 U9524 ( .A1(n8594), .A2(n8593), .ZN(n8597) );
  INV_X1 U9525 ( .A(n8643), .ZN(n7043) );
  NAND2_X1 U9526 ( .A1(n8498), .A2(n8497), .ZN(n8506) );
  NAND2_X1 U9527 ( .A1(n7029), .A2(n7027), .ZN(n8470) );
  NAND2_X1 U9528 ( .A1(n7176), .A2(n7174), .ZN(n11377) );
  NAND3_X1 U9529 ( .A1(n9522), .A2(n9521), .A3(n6609), .ZN(n6895) );
  NAND2_X1 U9530 ( .A1(n9603), .A2(n7511), .ZN(n7507) );
  NAND2_X1 U9531 ( .A1(n7480), .A2(n7479), .ZN(n9782) );
  NAND2_X1 U9532 ( .A1(n7486), .A2(n7485), .ZN(n9720) );
  NAND2_X1 U9533 ( .A1(n7483), .A2(n7482), .ZN(n9753) );
  NAND2_X1 U9534 ( .A1(n7567), .A2(n9620), .ZN(n9632) );
  MUX2_X1 U9535 ( .A(n10982), .B(n14038), .S(n9399), .Z(n9369) );
  INV_X1 U9536 ( .A(n7117), .ZN(n14525) );
  OAI21_X1 U9537 ( .B1(n14765), .B2(n14766), .A(n14569), .ZN(n7111) );
  NAND2_X1 U9538 ( .A1(n6909), .A2(n6911), .ZN(n11831) );
  INV_X1 U9539 ( .A(n6912), .ZN(n6909) );
  NOR2_X1 U9540 ( .A1(n6912), .A2(n6910), .ZN(n11941) );
  NAND2_X1 U9541 ( .A1(n11291), .A2(n6915), .ZN(n6911) );
  NAND4_X1 U9542 ( .A1(n6922), .A2(n12811), .A3(n6642), .A4(n6920), .ZN(
        P3_U3199) );
  NAND2_X1 U9543 ( .A1(n8932), .A2(n13022), .ZN(n6939) );
  NAND3_X1 U9544 ( .A1(n7456), .A2(n8919), .A3(n6573), .ZN(n7450) );
  NAND2_X1 U9545 ( .A1(n8546), .A2(n6604), .ZN(n6949) );
  NAND2_X1 U9546 ( .A1(n11958), .A2(n6957), .ZN(n6956) );
  INV_X1 U9547 ( .A(n7225), .ZN(n6963) );
  NAND3_X1 U9548 ( .A1(n7229), .A2(n7228), .A3(n12835), .ZN(n12836) );
  INV_X1 U9549 ( .A(n11113), .ZN(n6976) );
  AOI21_X1 U9550 ( .B1(n14014), .B2(n6990), .A(n6593), .ZN(n6989) );
  NAND2_X1 U9551 ( .A1(n11922), .A2(n6996), .ZN(n6995) );
  NAND2_X1 U9552 ( .A1(n9311), .A2(n9893), .ZN(n9903) );
  NAND2_X1 U9553 ( .A1(n11138), .A2(n11448), .ZN(n11324) );
  NOR2_X2 U9554 ( .A1(n12353), .A2(n14327), .ZN(n14096) );
  NAND2_X1 U9555 ( .A1(n8579), .A2(n8578), .ZN(n7018) );
  NAND2_X1 U9556 ( .A1(n8563), .A2(n8562), .ZN(n7019) );
  NAND2_X1 U9557 ( .A1(n8505), .A2(n7021), .ZN(n7020) );
  NAND2_X1 U9558 ( .A1(n8441), .A2(n7031), .ZN(n7029) );
  NAND2_X1 U9559 ( .A1(n8352), .A2(n7035), .ZN(n7034) );
  OAI21_X2 U9560 ( .B1(n8389), .B2(n7047), .A(n7045), .ZN(n8416) );
  NAND2_X1 U9561 ( .A1(n8708), .A2(n7054), .ZN(n7053) );
  NAND2_X1 U9562 ( .A1(n7053), .A2(n8725), .ZN(n8739) );
  NAND2_X1 U9563 ( .A1(n8708), .A2(n8707), .ZN(n8724) );
  NAND4_X1 U9564 ( .A1(n7568), .A2(n7064), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7058) );
  NAND4_X1 U9565 ( .A1(n7063), .A2(n12003), .A3(n7062), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7059) );
  NAND3_X1 U9566 ( .A1(n7062), .A2(n7063), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7060) );
  INV_X1 U9567 ( .A(n7623), .ZN(n7066) );
  NAND2_X1 U9568 ( .A1(n12266), .A2(n7083), .ZN(n7081) );
  OR2_X1 U9569 ( .A1(n12266), .A2(n8123), .ZN(n7086) );
  NAND2_X1 U9570 ( .A1(n7088), .A2(n7090), .ZN(n8010) );
  INV_X2 U9571 ( .A(n13416), .ZN(n7100) );
  NAND2_X1 U9572 ( .A1(n13379), .A2(n7101), .ZN(n13387) );
  NAND2_X1 U9573 ( .A1(n7102), .A2(n11674), .ZN(n13651) );
  NOR2_X2 U9574 ( .A1(n12172), .A2(n13782), .ZN(n12204) );
  NOR2_X2 U9575 ( .A1(n11910), .A2(n14868), .ZN(n12020) );
  NAND2_X2 U9576 ( .A1(n10069), .A2(n9975), .ZN(n9207) );
  NOR2_X2 U9577 ( .A1(n11079), .A2(n14991), .ZN(n11162) );
  NAND2_X1 U9578 ( .A1(n7566), .A2(n6496), .ZN(n7119) );
  NAND2_X1 U9579 ( .A1(n7119), .A2(n7120), .ZN(n11662) );
  OAI21_X1 U9580 ( .B1(n13643), .B2(n7125), .A(n7123), .ZN(n13591) );
  NAND4_X1 U9581 ( .A1(n7659), .A2(n7558), .A3(n7128), .A4(n7644), .ZN(n13787)
         );
  AOI21_X1 U9582 ( .B1(n11813), .B2(n6589), .A(n7140), .ZN(n12007) );
  NAND2_X1 U9583 ( .A1(n13500), .A2(n7148), .ZN(n7146) );
  AOI21_X2 U9584 ( .B1(n7150), .B2(n6515), .A(n7149), .ZN(n7148) );
  INV_X1 U9585 ( .A(n13414), .ZN(n7154) );
  AOI21_X1 U9586 ( .B1(n13565), .B2(n6594), .A(n7159), .ZN(n13409) );
  OR2_X1 U9587 ( .A1(n14237), .A2(n14259), .ZN(n7193) );
  NAND2_X1 U9588 ( .A1(n14336), .A2(n7197), .ZN(n7194) );
  NAND2_X1 U9589 ( .A1(n7194), .A2(n7195), .ZN(P1_U3523) );
  NAND2_X1 U9590 ( .A1(n14336), .A2(n7202), .ZN(n7196) );
  NAND2_X1 U9591 ( .A1(n14336), .A2(n14112), .ZN(n7200) );
  NAND2_X1 U9592 ( .A1(n7205), .A2(n7206), .ZN(n15107) );
  OAI21_X2 U9593 ( .B1(n7208), .B2(n6579), .A(n13168), .ZN(n13176) );
  OAI21_X1 U9594 ( .B1(n12800), .B2(n7227), .A(n7226), .ZN(n12845) );
  INV_X1 U9595 ( .A(n12833), .ZN(n7228) );
  NOR2_X1 U9596 ( .A1(n11279), .A2(n15058), .ZN(n11282) );
  XNOR2_X1 U9597 ( .A(n6492), .B(n12788), .ZN(n12767) );
  NOR2_X1 U9598 ( .A1(n11282), .A2(n11281), .ZN(n11841) );
  NAND2_X1 U9599 ( .A1(n11585), .A2(n11595), .ZN(n11637) );
  NOR2_X1 U9600 ( .A1(n7338), .A2(n7337), .ZN(n7336) );
  NAND2_X1 U9601 ( .A1(n11665), .A2(n11664), .ZN(n11813) );
  NAND2_X1 U9602 ( .A1(n13403), .A2(n13402), .ZN(n13565) );
  NAND2_X1 U9603 ( .A1(n13411), .A2(n13410), .ZN(n13519) );
  OAI21_X1 U9604 ( .B1(n13575), .B2(n7239), .A(n7237), .ZN(n13553) );
  NAND2_X1 U9605 ( .A1(n7236), .A2(n7235), .ZN(n13433) );
  NAND2_X1 U9606 ( .A1(n13575), .A2(n7237), .ZN(n7236) );
  NAND2_X1 U9607 ( .A1(n10861), .A2(n7252), .ZN(n9927) );
  NAND2_X1 U9608 ( .A1(n9918), .A2(n9921), .ZN(n7252) );
  NAND3_X1 U9609 ( .A1(n10922), .A2(n10863), .A3(n7253), .ZN(n9240) );
  NOR2_X1 U9610 ( .A1(n9918), .A2(n6624), .ZN(n7253) );
  NOR2_X1 U9611 ( .A1(n9918), .A2(n9917), .ZN(n7254) );
  NAND2_X1 U9612 ( .A1(n10465), .A2(n10501), .ZN(n7287) );
  OAI21_X1 U9613 ( .B1(n10465), .B2(n7288), .A(n10501), .ZN(n7286) );
  NAND3_X1 U9614 ( .A1(n6524), .A2(P3_REG2_REG_3__SCAN_IN), .A3(n7287), .ZN(
        n10484) );
  AND2_X1 U9615 ( .A1(n6524), .A2(n7287), .ZN(n10485) );
  INV_X1 U9616 ( .A(n7293), .ZN(n7291) );
  NAND2_X1 U9617 ( .A1(n12815), .A2(n7299), .ZN(n7295) );
  OAI21_X1 U9618 ( .B1(n12803), .B2(n7296), .A(n7295), .ZN(n12843) );
  NAND2_X1 U9619 ( .A1(n13963), .A2(n13964), .ZN(n13901) );
  NAND2_X1 U9620 ( .A1(n14005), .A2(n6597), .ZN(n7308) );
  OAI211_X1 U9621 ( .C1(n14005), .C2(n7314), .A(n7309), .B(n7308), .ZN(n13951)
         );
  NAND2_X1 U9622 ( .A1(n13978), .A2(n7320), .ZN(n13952) );
  NAND2_X1 U9623 ( .A1(n11632), .A2(n11755), .ZN(n7324) );
  NAND2_X1 U9624 ( .A1(n11122), .A2(n7332), .ZN(n7330) );
  AOI21_X1 U9625 ( .B1(n11121), .B2(n7332), .A(n6533), .ZN(n7331) );
  NAND2_X1 U9626 ( .A1(n9311), .A2(n9313), .ZN(n9316) );
  NAND2_X1 U9627 ( .A1(n9318), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9317) );
  NOR2_X1 U9628 ( .A1(n7348), .A2(n7347), .ZN(n7349) );
  INV_X4 U9629 ( .A(n13936), .ZN(n13902) );
  INV_X2 U9630 ( .A(n10801), .ZN(n13906) );
  INV_X1 U9631 ( .A(n8052), .ZN(n7356) );
  NAND2_X1 U9632 ( .A1(n13077), .A2(n7372), .ZN(n12931) );
  OAI21_X1 U9633 ( .B1(n11567), .B2(n7380), .A(n7379), .ZN(n11683) );
  OAI21_X1 U9634 ( .B1(n12130), .B2(n7397), .A(n7393), .ZN(n12257) );
  OAI21_X1 U9635 ( .B1(n12130), .B2(n8520), .A(n12603), .ZN(n12186) );
  NAND3_X1 U9636 ( .A1(n15087), .A2(n12536), .A3(n12541), .ZN(n8774) );
  NAND2_X1 U9637 ( .A1(n14128), .A2(n14123), .ZN(n7430) );
  INV_X1 U9638 ( .A(n9715), .ZN(n14471) );
  NAND2_X1 U9639 ( .A1(n9715), .A2(n9825), .ZN(n9717) );
  INV_X1 U9640 ( .A(SI_18_), .ZN(n7434) );
  INV_X1 U9641 ( .A(n7958), .ZN(n7438) );
  NAND2_X1 U9642 ( .A1(n8890), .A2(n8889), .ZN(n7441) );
  NAND2_X1 U9643 ( .A1(n10728), .A2(n10729), .ZN(n8896) );
  NAND3_X1 U9644 ( .A1(n7446), .A2(n8938), .A3(n12975), .ZN(n12447) );
  NAND2_X1 U9645 ( .A1(n8937), .A2(n8936), .ZN(n8938) );
  NAND3_X1 U9646 ( .A1(n8919), .A2(n7456), .A3(n7455), .ZN(n7452) );
  NAND2_X1 U9647 ( .A1(n7465), .A2(n6531), .ZN(n7457) );
  NAND2_X1 U9648 ( .A1(n11088), .A2(n8906), .ZN(n7468) );
  INV_X1 U9649 ( .A(n7477), .ZN(n11557) );
  NAND2_X1 U9650 ( .A1(n9549), .A2(n9550), .ZN(n9548) );
  NAND3_X1 U9651 ( .A1(n9758), .A2(n9757), .A3(n6607), .ZN(n7480) );
  INV_X1 U9652 ( .A(n9771), .ZN(n7481) );
  NAND3_X1 U9653 ( .A1(n9725), .A2(n9724), .A3(n6614), .ZN(n7483) );
  INV_X1 U9654 ( .A(n9738), .ZN(n7484) );
  NAND3_X1 U9655 ( .A1(n9691), .A2(n9690), .A3(n6608), .ZN(n7486) );
  INV_X1 U9656 ( .A(n9702), .ZN(n7487) );
  NAND2_X1 U9657 ( .A1(n9457), .A2(n7491), .ZN(n7490) );
  NAND2_X1 U9658 ( .A1(n9649), .A2(n7494), .ZN(n7498) );
  NAND2_X1 U9659 ( .A1(n7498), .A2(n7496), .ZN(n9671) );
  AOI21_X2 U9660 ( .B1(n9603), .B2(n7506), .A(n7504), .ZN(n9619) );
  INV_X1 U9661 ( .A(n9088), .ZN(n7522) );
  INV_X1 U9662 ( .A(n9087), .ZN(n7523) );
  NAND2_X1 U9663 ( .A1(n7524), .A2(n9224), .ZN(n9230) );
  OAI211_X1 U9664 ( .C1(n9171), .C2(n7527), .A(n7525), .B(n7552), .ZN(n7524)
         );
  NOR2_X1 U9665 ( .A1(n7530), .A2(n9154), .ZN(n7529) );
  INV_X1 U9666 ( .A(n9062), .ZN(n7537) );
  NAND3_X1 U9667 ( .A1(n9131), .A2(n9130), .A3(n6606), .ZN(n7538) );
  NAND2_X1 U9668 ( .A1(n7541), .A2(n7543), .ZN(n9148) );
  NAND3_X1 U9669 ( .A1(n7659), .A2(n7558), .A3(n7644), .ZN(n7546) );
  NAND2_X1 U9670 ( .A1(n8213), .A2(n7546), .ZN(n13800) );
  AND2_X1 U9671 ( .A1(n10717), .A2(n10716), .ZN(n10718) );
  NAND2_X1 U9672 ( .A1(n14335), .A2(n14334), .ZN(n14419) );
  INV_X1 U9673 ( .A(n14333), .ZN(n14334) );
  OAI21_X1 U9674 ( .B1(n13464), .B2(n6699), .A(n13463), .ZN(n13666) );
  OAI21_X1 U9675 ( .B1(n14332), .B2(n14819), .A(n14331), .ZN(n14333) );
  NAND2_X1 U9676 ( .A1(n8784), .A2(n6516), .ZN(n8785) );
  INV_X1 U9677 ( .A(n13658), .ZN(n13665) );
  INV_X2 U9678 ( .A(n8181), .ZN(n8159) );
  INV_X1 U9679 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9482) );
  NAND2_X1 U9680 ( .A1(n9295), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9296) );
  NAND2_X1 U9681 ( .A1(n9272), .A2(n8963), .ZN(n8988) );
  NAND2_X1 U9682 ( .A1(n8534), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8280) );
  OR2_X1 U9683 ( .A1(n12323), .A2(n12341), .ZN(n12324) );
  NAND2_X1 U9684 ( .A1(n12323), .A2(n12341), .ZN(n12364) );
  OR2_X2 U9685 ( .A1(n9571), .A2(n9570), .ZN(n9603) );
  NOR2_X1 U9686 ( .A1(n11054), .A2(n11351), .ZN(n11041) );
  NAND2_X1 U9687 ( .A1(n7668), .A2(n12284), .ZN(n9920) );
  NAND2_X4 U9688 ( .A1(n9360), .A2(n9359), .ZN(n14040) );
  NAND2_X1 U9689 ( .A1(n12265), .A2(n14453), .ZN(n9387) );
  NAND2_X1 U9690 ( .A1(n7701), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7706) );
  NOR3_X1 U9691 ( .A1(n9890), .A2(n9889), .A3(n9888), .ZN(n9897) );
  AND2_X2 U9692 ( .A1(n9935), .A2(n9923), .ZN(n8996) );
  INV_X1 U9693 ( .A(n14356), .ZN(n12345) );
  INV_X1 U9694 ( .A(n14176), .ZN(n12337) );
  OR2_X1 U9695 ( .A1(n8090), .A2(n8089), .ZN(n7547) );
  AND2_X1 U9696 ( .A1(n8299), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7549) );
  OR2_X1 U9697 ( .A1(n15198), .A2(n14032), .ZN(n7551) );
  AND2_X1 U9698 ( .A1(n13659), .A2(n14990), .ZN(n7553) );
  OR2_X1 U9699 ( .A1(n13678), .A2(n13438), .ZN(n7554) );
  AND2_X1 U9700 ( .A1(n10848), .A2(n9492), .ZN(n7555) );
  AND3_X1 U9701 ( .A1(n9287), .A2(n9306), .A3(n9323), .ZN(n7556) );
  INV_X1 U9702 ( .A(n14286), .ZN(n14631) );
  INV_X1 U9703 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n7722) );
  AND2_X1 U9704 ( .A1(n12876), .A2(n14692), .ZN(n7559) );
  INV_X1 U9705 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9314) );
  AND2_X1 U9706 ( .A1(n14860), .A2(n11080), .ZN(n13189) );
  INV_X1 U9707 ( .A(n13189), .ZN(n8233) );
  INV_X1 U9708 ( .A(n13444), .ZN(n13296) );
  AND2_X1 U9709 ( .A1(n9200), .A2(n9220), .ZN(n7560) );
  AND2_X2 U9710 ( .A1(n12358), .A2(n14611), .ZN(n14630) );
  INV_X1 U9711 ( .A(n10601), .ZN(n13812) );
  INV_X1 U9712 ( .A(n12702), .ZN(n12975) );
  OR2_X1 U9713 ( .A1(n10719), .A2(n13812), .ZN(n7563) );
  NAND2_X1 U9714 ( .A1(n8969), .A2(n12657), .ZN(n15094) );
  XNOR2_X1 U9715 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7565) );
  INV_X1 U9716 ( .A(n12307), .ZN(n14291) );
  AND2_X2 U9717 ( .A1(n10579), .A2(n8873), .ZN(n15193) );
  NAND2_X1 U9718 ( .A1(n15176), .A2(n15080), .ZN(n13162) );
  INV_X1 U9719 ( .A(n13162), .ZN(n8837) );
  AND2_X2 U9720 ( .A1(n8835), .A2(n8967), .ZN(n15176) );
  INV_X1 U9721 ( .A(n10848), .ZN(n9365) );
  NAND2_X1 U9722 ( .A1(n8996), .A2(n10323), .ZN(n9000) );
  NAND2_X1 U9723 ( .A1(n9370), .A2(n9369), .ZN(n9371) );
  NAND2_X1 U9724 ( .A1(n9011), .A2(n9010), .ZN(n9016) );
  INV_X1 U9725 ( .A(n9022), .ZN(n9023) );
  NAND2_X1 U9726 ( .A1(n7548), .A2(n9024), .ZN(n9029) );
  INV_X1 U9727 ( .A(n9053), .ZN(n9054) );
  NAND2_X1 U9728 ( .A1(n9079), .A2(n9078), .ZN(n9084) );
  INV_X1 U9729 ( .A(n9142), .ZN(n9143) );
  INV_X1 U9730 ( .A(n9158), .ZN(n9159) );
  INV_X1 U9731 ( .A(n9161), .ZN(n9162) );
  NOR2_X1 U9732 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n9287) );
  INV_X1 U9733 ( .A(n9798), .ZN(n9799) );
  INV_X1 U9734 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9288) );
  OR2_X1 U9735 ( .A1(n9223), .A2(n9222), .ZN(n9224) );
  INV_X1 U9736 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7633) );
  INV_X1 U9737 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7640) );
  INV_X1 U9738 ( .A(n9840), .ZN(n9808) );
  AND2_X1 U9739 ( .A1(n10398), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10391) );
  INV_X1 U9740 ( .A(n12601), .ZN(n8520) );
  INV_X1 U9741 ( .A(n12889), .ZN(n8848) );
  INV_X1 U9742 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8259) );
  INV_X1 U9743 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7851) );
  INV_X1 U9744 ( .A(n9002), .ZN(n9236) );
  INV_X1 U9745 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7641) );
  INV_X1 U9746 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n7638) );
  INV_X1 U9747 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7804) );
  INV_X1 U9748 ( .A(n14715), .ZN(n13836) );
  OR2_X1 U9749 ( .A1(n13841), .A2(n13840), .ZN(n13842) );
  NAND2_X1 U9750 ( .A1(n9808), .A2(n9843), .ZN(n9824) );
  INV_X1 U9751 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9507) );
  INV_X1 U9752 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9293) );
  INV_X1 U9753 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n15376) );
  XNOR2_X1 U9754 ( .A(n12952), .B(n10646), .ZN(n8941) );
  OR2_X1 U9755 ( .A1(n8729), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8745) );
  OR2_X1 U9756 ( .A1(n8647), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8666) );
  AND2_X1 U9757 ( .A1(n11028), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n11015) );
  OR2_X1 U9758 ( .A1(n8666), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8680) );
  INV_X1 U9759 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n8433) );
  INV_X1 U9760 ( .A(n8993), .ZN(n9259) );
  AND2_X1 U9761 ( .A1(n10527), .A2(n7781), .ZN(n7782) );
  INV_X1 U9762 ( .A(n8098), .ZN(n8099) );
  INV_X1 U9763 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8019) );
  NAND2_X1 U9764 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n8099), .ZN(n8138) );
  INV_X1 U9765 ( .A(n13744), .ZN(n12019) );
  OR2_X1 U9766 ( .A1(n8220), .A2(n14972), .ZN(n8242) );
  NAND2_X1 U9767 ( .A1(n13409), .A2(n13408), .ZN(n13516) );
  INV_X1 U9768 ( .A(n12020), .ZN(n12018) );
  INV_X1 U9769 ( .A(n11108), .ZN(n10802) );
  INV_X1 U9770 ( .A(n9675), .ZN(n9676) );
  AND3_X1 U9771 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n9424) );
  OR2_X1 U9772 ( .A1(n10680), .A2(n10679), .ZN(n10758) );
  INV_X1 U9773 ( .A(n14385), .ZN(n12344) );
  OR2_X1 U9774 ( .A1(n9523), .A2(n10296), .ZN(n9536) );
  NAND2_X1 U9775 ( .A1(n7624), .A2(n12262), .ZN(n7627) );
  NOR2_X1 U9776 ( .A1(n14512), .A2(n14511), .ZN(n14503) );
  AND2_X1 U9777 ( .A1(n8952), .A2(n8951), .ZN(n12399) );
  INV_X1 U9778 ( .A(n12439), .ZN(n12472) );
  NOR2_X1 U9779 ( .A1(n8745), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12872) );
  NOR2_X1 U9780 ( .A1(n11016), .A2(n11015), .ZN(n11274) );
  INV_X1 U9781 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14497) );
  INV_X1 U9782 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14501) );
  AND2_X1 U9783 ( .A1(n10254), .A2(n10244), .ZN(n10266) );
  INV_X1 U9784 ( .A(n12983), .ZN(n13028) );
  INV_X1 U9785 ( .A(n12182), .ZN(n12606) );
  OR3_X1 U9786 ( .A1(n8477), .A2(P3_REG3_REG_11__SCAN_IN), .A3(
        P3_REG3_REG_12__SCAN_IN), .ZN(n8486) );
  NOR2_X1 U9787 ( .A1(n8377), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8426) );
  INV_X1 U9788 ( .A(n12859), .ZN(n12501) );
  AND2_X1 U9789 ( .A1(n8871), .A2(n12675), .ZN(n10578) );
  AND2_X1 U9790 ( .A1(n6516), .A2(n12599), .ZN(n14649) );
  AND2_X1 U9791 ( .A1(n8827), .A2(n12690), .ZN(n15078) );
  INV_X1 U9792 ( .A(n15075), .ZN(n15116) );
  NAND2_X1 U9793 ( .A1(n8472), .A2(n8471), .ZN(n8495) );
  NAND2_X1 U9794 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8286) );
  INV_X1 U9795 ( .A(n11409), .ZN(n7900) );
  INV_X1 U9796 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n11266) );
  INV_X1 U9797 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7943) );
  AND2_X1 U9798 ( .A1(n8037), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8039) );
  AND2_X1 U9799 ( .A1(n9267), .A2(n10067), .ZN(n10629) );
  OR3_X1 U9800 ( .A1(n12195), .A2(n12194), .A3(n12193), .ZN(n13742) );
  NAND2_X1 U9801 ( .A1(n14700), .A2(n14701), .ZN(n14699) );
  AND2_X1 U9802 ( .A1(n11860), .A2(n11857), .ZN(n11858) );
  INV_X1 U9803 ( .A(n14024), .ZN(n13948) );
  OR2_X1 U9804 ( .A1(n13892), .A2(n13891), .ZN(n13893) );
  NAND2_X1 U9805 ( .A1(n11786), .A2(n11787), .ZN(n11859) );
  INV_X1 U9806 ( .A(n14703), .ZN(n14728) );
  XNOR2_X1 U9807 ( .A(n11107), .B(n10802), .ZN(n10807) );
  NOR2_X1 U9808 ( .A1(n9829), .A2(n11981), .ZN(n10564) );
  AND2_X1 U9809 ( .A1(n9621), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9637) );
  INV_X1 U9810 ( .A(n6475), .ZN(n9790) );
  INV_X1 U9811 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14517) );
  INV_X1 U9812 ( .A(n14181), .ZN(n14195) );
  NOR2_X1 U9813 ( .A1(n9536), .A2(n12050), .ZN(n9556) );
  INV_X1 U9814 ( .A(n14140), .ZN(n14147) );
  INV_X1 U9815 ( .A(n14814), .ZN(n14822) );
  NOR2_X1 U9816 ( .A1(n10572), .A2(P1_U3086), .ZN(n10595) );
  NOR2_X1 U9817 ( .A1(n9989), .A2(n14465), .ZN(n10556) );
  NOR2_X1 U9818 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n14521), .ZN(n14485) );
  OAI21_X1 U9819 ( .B1(n13129), .B2(n12477), .A(n9279), .ZN(n9280) );
  INV_X1 U9820 ( .A(n12034), .ZN(n12474) );
  AND2_X1 U9821 ( .A1(n12496), .A2(n12495), .ZN(n12866) );
  INV_X1 U9822 ( .A(n13165), .ZN(n10027) );
  AND4_X1 U9823 ( .A1(n8575), .A2(n8574), .A3(n8573), .A4(n8572), .ZN(n12418)
         );
  INV_X1 U9824 ( .A(n15094), .ZN(n15109) );
  NAND2_X1 U9825 ( .A1(n12501), .A2(n10890), .ZN(n15117) );
  AND2_X1 U9826 ( .A1(n8867), .A2(n8866), .ZN(n10579) );
  NOR2_X1 U9827 ( .A1(n15176), .A2(n8861), .ZN(n8862) );
  NAND2_X1 U9828 ( .A1(n8798), .A2(n12529), .ZN(n15169) );
  OR2_X1 U9829 ( .A1(n15075), .A2(n15166), .ZN(n14692) );
  INV_X1 U9830 ( .A(n15148), .ZN(n15166) );
  INV_X1 U9831 ( .A(n15169), .ZN(n15080) );
  AND2_X1 U9832 ( .A1(n11803), .A2(n7973), .ZN(n7974) );
  INV_X1 U9833 ( .A(n13254), .ZN(n13284) );
  AND4_X1 U9834 ( .A1(n8118), .A2(n8117), .A3(n8116), .A4(n8115), .ZN(n13485)
         );
  AND2_X1 U9835 ( .A1(n13373), .A2(n10704), .ZN(n13374) );
  INV_X1 U9836 ( .A(n14873), .ZN(n14943) );
  AND2_X1 U9837 ( .A1(n13459), .A2(n13458), .ZN(n13667) );
  INV_X1 U9838 ( .A(n13594), .ZN(n13576) );
  AND2_X1 U9839 ( .A1(n13393), .A2(n12203), .ZN(n13733) );
  INV_X1 U9840 ( .A(n14958), .ZN(n13649) );
  NAND2_X2 U9841 ( .A1(n14973), .A2(n8237), .ZN(n14950) );
  AND2_X1 U9842 ( .A1(n8215), .A2(n8214), .ZN(n14965) );
  AND2_X1 U9843 ( .A1(n9915), .A2(n10068), .ZN(n8239) );
  AND2_X1 U9844 ( .A1(n8203), .A2(n8206), .ZN(n8226) );
  AND2_X1 U9845 ( .A1(n7870), .A2(n7904), .ZN(n10108) );
  AND2_X1 U9846 ( .A1(n9579), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9591) );
  INV_X1 U9847 ( .A(n14745), .ZN(n12234) );
  INV_X1 U9848 ( .A(n14015), .ZN(n15200) );
  NOR2_X1 U9849 ( .A1(n10571), .A2(n10559), .ZN(n10567) );
  INV_X1 U9850 ( .A(n12245), .ZN(n9896) );
  AND2_X1 U9851 ( .A1(n9657), .A2(n9656), .ZN(n13956) );
  AND4_X1 U9852 ( .A1(n9585), .A2(n9584), .A3(n9583), .A4(n9582), .ZN(n12139)
         );
  OR2_X1 U9853 ( .A1(n10158), .A2(n10157), .ZN(n14781) );
  AND2_X1 U9854 ( .A1(n10161), .A2(n14459), .ZN(n14083) );
  INV_X1 U9855 ( .A(n14781), .ZN(n14074) );
  INV_X1 U9856 ( .A(n12310), .ZN(n14258) );
  NAND2_X1 U9857 ( .A1(n10569), .A2(n10568), .ZN(n14611) );
  INV_X1 U9858 ( .A(n14831), .ZN(n14255) );
  OAI21_X1 U9859 ( .B1(n10547), .B2(P1_D_REG_0__SCAN_IN), .A(n10545), .ZN(
        n11035) );
  AND2_X1 U9860 ( .A1(n14797), .A2(n14796), .ZN(n14819) );
  INV_X1 U9861 ( .A(n14819), .ZN(n14842) );
  INV_X1 U9862 ( .A(n11035), .ZN(n10598) );
  OR2_X1 U9863 ( .A1(n9993), .A2(n9992), .ZN(n10545) );
  INV_X1 U9864 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9306) );
  INV_X1 U9865 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14543) );
  AND2_X1 U9866 ( .A1(n10254), .A2(n10253), .ZN(n15028) );
  NOR2_X1 U9867 ( .A1(n8986), .A2(n8985), .ZN(n8987) );
  INV_X1 U9868 ( .A(n12468), .ZN(n12462) );
  AND2_X1 U9869 ( .A1(n8982), .A2(n8981), .ZN(n12034) );
  NAND2_X1 U9870 ( .A1(n8753), .A2(n8752), .ZN(n12889) );
  NAND2_X1 U9871 ( .A1(n8636), .A2(n8635), .ZN(n12988) );
  INV_X1 U9872 ( .A(n8921), .ZN(n14658) );
  INV_X1 U9873 ( .A(n12862), .ZN(n15060) );
  INV_X1 U9874 ( .A(n11289), .ZN(n15056) );
  INV_X1 U9875 ( .A(n15120), .ZN(n12944) );
  INV_X1 U9876 ( .A(n15193), .ZN(n15190) );
  NAND2_X1 U9877 ( .A1(n15193), .A2(n15080), .ZN(n13116) );
  INV_X1 U9878 ( .A(n12387), .ZN(n13146) );
  INV_X1 U9879 ( .A(n15176), .ZN(n15174) );
  NAND2_X1 U9880 ( .A1(n8810), .A2(n6518), .ZN(n11696) );
  INV_X1 U9881 ( .A(SI_16_), .ZN(n10383) );
  INV_X1 U9882 ( .A(SI_11_), .ZN(n10008) );
  INV_X1 U9883 ( .A(n13170), .ZN(n12293) );
  NAND2_X1 U9884 ( .A1(n10418), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14870) );
  INV_X1 U9885 ( .A(n14860), .ZN(n13269) );
  OR2_X1 U9886 ( .A1(n9270), .A2(n9269), .ZN(n9271) );
  INV_X1 U9887 ( .A(n13484), .ZN(n13297) );
  OAI21_X1 U9888 ( .B1(n13202), .B2(n8247), .A(n7686), .ZN(n13577) );
  INV_X1 U9889 ( .A(n14939), .ZN(n14874) );
  OR2_X1 U9890 ( .A1(n14964), .A2(n6864), .ZN(n14958) );
  OR2_X1 U9891 ( .A1(n14964), .A2(n11000), .ZN(n13646) );
  INV_X1 U9892 ( .A(n15027), .ZN(n15025) );
  AND2_X2 U9893 ( .A1(n10632), .A2(n10631), .ZN(n15027) );
  INV_X1 U9894 ( .A(n13419), .ZN(n13779) );
  AND3_X1 U9895 ( .A1(n14998), .A2(n14997), .A3(n14996), .ZN(n15023) );
  OR2_X1 U9896 ( .A1(n10630), .A2(n10624), .ZN(n15017) );
  NOR2_X1 U9897 ( .A1(n14970), .A2(n14965), .ZN(n14966) );
  INV_X1 U9898 ( .A(n14966), .ZN(n14967) );
  INV_X1 U9899 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n12251) );
  INV_X1 U9900 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11173) );
  INV_X1 U9901 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10001) );
  NAND2_X1 U9902 ( .A1(n11098), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15204) );
  INV_X1 U9903 ( .A(n14193), .ZN(n14361) );
  INV_X1 U9904 ( .A(n15197), .ZN(n14707) );
  INV_X1 U9905 ( .A(n12139), .ZN(n14621) );
  OR2_X1 U9906 ( .A1(n10158), .A2(n10156), .ZN(n11995) );
  INV_X1 U9907 ( .A(n14604), .ZN(n14300) );
  AND2_X1 U9908 ( .A1(n14171), .A2(n11040), .ZN(n14286) );
  INV_X1 U9909 ( .A(n14388), .ZN(n14853) );
  NAND2_X1 U9910 ( .A1(n14845), .A2(n14828), .ZN(n14446) );
  OR2_X1 U9911 ( .A1(n10946), .A2(n10598), .ZN(n14843) );
  INV_X2 U9912 ( .A(n14843), .ZN(n14845) );
  AND2_X1 U9913 ( .A1(n9973), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9994) );
  NAND2_X1 U9914 ( .A1(n9906), .A2(n9905), .ZN(n14469) );
  INV_X1 U9915 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11765) );
  INV_X1 U9916 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10613) );
  INV_X2 U9917 ( .A(n12703), .ZN(P3_U3897) );
  AND2_X1 U9918 ( .A1(n10541), .A2(n9994), .ZN(P1_U4016) );
  AND2_X1 U9919 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n7569) );
  NAND2_X1 U9920 ( .A1(n9975), .A2(n7569), .ZN(n9352) );
  AND2_X1 U9921 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7570) );
  NAND2_X1 U9922 ( .A1(n7580), .A2(n7570), .ZN(n7712) );
  NAND2_X1 U9923 ( .A1(n9352), .A2(n7712), .ZN(n7707) );
  INV_X1 U9924 ( .A(SI_1_), .ZN(n10011) );
  NOR2_X1 U9925 ( .A1(n7571), .A2(n10011), .ZN(n7572) );
  INV_X1 U9926 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9944) );
  MUX2_X1 U9927 ( .A(n9944), .B(n9956), .S(n7580), .Z(n7573) );
  INV_X1 U9928 ( .A(n7573), .ZN(n7574) );
  NAND2_X1 U9929 ( .A1(n7574), .A2(SI_2_), .ZN(n7575) );
  MUX2_X1 U9930 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n7580), .Z(n7577) );
  XNOR2_X1 U9931 ( .A(n7577), .B(SI_3_), .ZN(n7751) );
  INV_X1 U9932 ( .A(n7751), .ZN(n7576) );
  NAND2_X1 U9933 ( .A1(n7577), .A2(SI_3_), .ZN(n7578) );
  NAND2_X1 U9934 ( .A1(n7579), .A2(n7578), .ZN(n7765) );
  INV_X2 U9935 ( .A(n7580), .ZN(n9975) );
  MUX2_X1 U9936 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n7580), .Z(n7582) );
  XNOR2_X1 U9937 ( .A(n7582), .B(SI_4_), .ZN(n7766) );
  INV_X1 U9938 ( .A(n7766), .ZN(n7581) );
  NAND2_X1 U9939 ( .A1(n7765), .A2(n7581), .ZN(n7584) );
  NAND2_X1 U9940 ( .A1(n7582), .A2(SI_4_), .ZN(n7583) );
  INV_X1 U9941 ( .A(n7786), .ZN(n7585) );
  NAND2_X1 U9942 ( .A1(n7785), .A2(n7585), .ZN(n7588) );
  NAND2_X1 U9943 ( .A1(n7586), .A2(SI_5_), .ZN(n7587) );
  NAND2_X1 U9944 ( .A1(n7588), .A2(n7587), .ZN(n7801) );
  MUX2_X1 U9945 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9945), .Z(n7590) );
  XNOR2_X1 U9946 ( .A(n7590), .B(SI_6_), .ZN(n7802) );
  INV_X1 U9947 ( .A(n7802), .ZN(n7589) );
  NAND2_X1 U9948 ( .A1(n7801), .A2(n7589), .ZN(n7592) );
  NAND2_X1 U9949 ( .A1(n7590), .A2(SI_6_), .ZN(n7591) );
  MUX2_X1 U9950 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9945), .Z(n7594) );
  XNOR2_X1 U9951 ( .A(n7594), .B(SI_7_), .ZN(n7824) );
  INV_X1 U9952 ( .A(n7824), .ZN(n7593) );
  NAND2_X1 U9953 ( .A1(n7594), .A2(SI_7_), .ZN(n7595) );
  MUX2_X1 U9954 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9945), .Z(n7843) );
  INV_X1 U9955 ( .A(n7843), .ZN(n7597) );
  MUX2_X1 U9956 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9945), .Z(n7598) );
  NAND2_X1 U9957 ( .A1(n7598), .A2(SI_9_), .ZN(n7599) );
  OAI21_X1 U9958 ( .B1(n7598), .B2(SI_9_), .A(n7599), .ZN(n7862) );
  MUX2_X1 U9959 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9945), .Z(n7600) );
  NAND2_X1 U9960 ( .A1(n7600), .A2(SI_10_), .ZN(n7602) );
  OAI21_X1 U9961 ( .B1(n7600), .B2(SI_10_), .A(n7602), .ZN(n7601) );
  INV_X1 U9962 ( .A(n7601), .ZN(n7883) );
  MUX2_X1 U9963 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n9945), .Z(n7603) );
  XNOR2_X1 U9964 ( .A(n7603), .B(SI_11_), .ZN(n7902) );
  INV_X1 U9965 ( .A(n7603), .ZN(n7604) );
  NAND2_X1 U9966 ( .A1(n7604), .A2(n10008), .ZN(n7605) );
  MUX2_X1 U9967 ( .A(n8496), .B(n10504), .S(n9945), .Z(n7606) );
  XNOR2_X1 U9968 ( .A(n7606), .B(SI_12_), .ZN(n7920) );
  MUX2_X1 U9969 ( .A(n10613), .B(n10615), .S(n9945), .Z(n7607) );
  NAND2_X1 U9970 ( .A1(n7939), .A2(n7938), .ZN(n7609) );
  NAND2_X1 U9971 ( .A1(n7607), .A2(n10115), .ZN(n7608) );
  NAND2_X1 U9972 ( .A1(n7610), .A2(n10129), .ZN(n7611) );
  MUX2_X1 U9973 ( .A(n8524), .B(n10791), .S(n9945), .Z(n7958) );
  MUX2_X1 U9974 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n9945), .Z(n7612) );
  INV_X1 U9975 ( .A(n7612), .ZN(n7613) );
  NAND2_X1 U9976 ( .A1(n7613), .A2(n15360), .ZN(n7614) );
  MUX2_X1 U9977 ( .A(n11171), .B(n11173), .S(n9945), .Z(n7615) );
  NAND2_X1 U9978 ( .A1(n7615), .A2(n10383), .ZN(n7618) );
  INV_X1 U9979 ( .A(n8010), .ZN(n7616) );
  NAND2_X1 U9980 ( .A1(n7616), .A2(SI_17_), .ZN(n7622) );
  MUX2_X1 U9981 ( .A(n11346), .B(n11348), .S(n9945), .Z(n8008) );
  INV_X1 U9982 ( .A(n8008), .ZN(n7617) );
  AND2_X1 U9983 ( .A1(n7618), .A2(n7617), .ZN(n7619) );
  MUX2_X1 U9984 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9945), .Z(n7688) );
  MUX2_X1 U9985 ( .A(n11765), .B(n12285), .S(n9945), .Z(n7624) );
  INV_X1 U9986 ( .A(SI_19_), .ZN(n12262) );
  INV_X1 U9987 ( .A(n7624), .ZN(n7625) );
  NAND2_X1 U9988 ( .A1(n7625), .A2(SI_19_), .ZN(n7626) );
  INV_X1 U9989 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11940) );
  MUX2_X1 U9990 ( .A(n11902), .B(n11940), .S(n9945), .Z(n8055) );
  INV_X1 U9991 ( .A(n8055), .ZN(n8054) );
  NAND2_X1 U9992 ( .A1(n8045), .A2(n8054), .ZN(n7630) );
  INV_X1 U9993 ( .A(n8061), .ZN(n7628) );
  NAND2_X1 U9994 ( .A1(n7628), .A2(SI_20_), .ZN(n7629) );
  NAND2_X1 U9995 ( .A1(n7630), .A2(n7629), .ZN(n7632) );
  MUX2_X1 U9996 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9945), .Z(n8056) );
  XNOR2_X1 U9997 ( .A(n8056), .B(SI_21_), .ZN(n7631) );
  NOR2_X1 U9998 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n7636) );
  NAND4_X1 U9999 ( .A1(n7655), .A2(n6764), .A3(n8199), .A4(n7638), .ZN(n8201)
         );
  NOR2_X1 U10000 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .ZN(n7639) );
  NAND2_X1 U10001 ( .A1(n11980), .A2(n9209), .ZN(n7643) );
  INV_X1 U10002 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11985) );
  OR2_X1 U10003 ( .A1(n9207), .A2(n11985), .ZN(n7642) );
  NAND2_X1 U10004 ( .A1(n8202), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7645) );
  INV_X1 U10005 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7647) );
  AND2_X1 U10006 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n7648) );
  NAND2_X1 U10007 ( .A1(n7963), .A2(n7648), .ZN(n7654) );
  INV_X1 U10008 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7649) );
  NAND2_X1 U10009 ( .A1(n7649), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n7651) );
  XNOR2_X1 U10010 ( .A(P2_IR_REG_20__SCAN_IN), .B(P2_IR_REG_31__SCAN_IN), .ZN(
        n7650) );
  OAI21_X1 U10011 ( .B1(n7652), .B2(n7651), .A(n7650), .ZN(n7653) );
  XNOR2_X1 U10012 ( .A(n8993), .B(n9923), .ZN(n7668) );
  INV_X1 U10013 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7982) );
  AND3_X1 U10014 ( .A1(n7657), .A2(n7656), .A3(n7982), .ZN(n7658) );
  INV_X1 U10015 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7660) );
  NAND2_X1 U10016 ( .A1(n7662), .A2(n7660), .ZN(n7667) );
  AND2_X1 U10017 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n7665) );
  INV_X1 U10018 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7661) );
  NAND3_X1 U10019 ( .A1(n7662), .A2(n7661), .A3(P2_IR_REG_19__SCAN_IN), .ZN(
        n7664) );
  XNOR2_X1 U10020 ( .A(P2_IR_REG_19__SCAN_IN), .B(P2_IR_REG_31__SCAN_IN), .ZN(
        n7663) );
  XNOR2_X1 U10021 ( .A(n13568), .B(n6809), .ZN(n8051) );
  NAND2_X1 U10022 ( .A1(n7792), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7811) );
  NOR2_X1 U10023 ( .A1(n7811), .A2(n7810), .ZN(n7832) );
  NAND2_X1 U10024 ( .A1(n7832), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7852) );
  INV_X1 U10025 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7925) );
  INV_X1 U10026 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11807) );
  NAND2_X1 U10027 ( .A1(n7987), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8002) );
  INV_X1 U10028 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n13232) );
  OR2_X1 U10029 ( .A1(n8039), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n7669) );
  AND2_X1 U10030 ( .A1(n7669), .A2(n8064), .ZN(n13569) );
  XNOR2_X2 U10031 ( .A(n7670), .B(n7671), .ZN(n7720) );
  INV_X1 U10033 ( .A(n8247), .ZN(n7947) );
  NAND2_X1 U10034 ( .A1(n13569), .A2(n7947), .ZN(n7677) );
  INV_X1 U10035 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13707) );
  NAND2_X1 U10036 ( .A1(n7701), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7674) );
  NAND2_X1 U10037 ( .A1(n7702), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7673) );
  OAI211_X1 U10038 ( .C1(n7736), .C2(n13707), .A(n7674), .B(n7673), .ZN(n7675)
         );
  INV_X1 U10039 ( .A(n7675), .ZN(n7676) );
  NAND2_X1 U10040 ( .A1(n7677), .A2(n7676), .ZN(n13579) );
  NAND2_X1 U10041 ( .A1(n13579), .A2(n11080), .ZN(n8052) );
  XNOR2_X1 U10042 ( .A(n7679), .B(n7678), .ZN(n11764) );
  NAND2_X1 U10043 ( .A1(n11764), .A2(n9209), .ZN(n7681) );
  INV_X4 U10044 ( .A(n10069), .ZN(n8015) );
  AOI22_X1 U10045 ( .A1(n8016), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8015), 
        .B2(n6864), .ZN(n7680) );
  XNOR2_X1 U10046 ( .A(n13603), .B(n6809), .ZN(n8035) );
  NOR2_X1 U10047 ( .A1(n7695), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n7682) );
  OR2_X1 U10048 ( .A1(n8037), .A2(n7682), .ZN(n13202) );
  INV_X1 U10049 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13718) );
  NAND2_X1 U10050 ( .A1(n7701), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n7684) );
  NAND2_X1 U10051 ( .A1(n7702), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n7683) );
  OAI211_X1 U10052 ( .C1(n7736), .C2(n13718), .A(n7684), .B(n7683), .ZN(n7685)
         );
  INV_X1 U10053 ( .A(n7685), .ZN(n7686) );
  NAND2_X1 U10054 ( .A1(n13577), .A2(n11080), .ZN(n8036) );
  XNOR2_X1 U10055 ( .A(n8035), .B(n8036), .ZN(n13200) );
  NAND2_X1 U10056 ( .A1(n7687), .A2(n7688), .ZN(n7689) );
  NAND2_X1 U10057 ( .A1(n7690), .A2(n7689), .ZN(n11547) );
  NAND2_X1 U10058 ( .A1(n11547), .A2(n9209), .ZN(n7693) );
  NAND2_X1 U10059 ( .A1(n8013), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7691) );
  XNOR2_X1 U10060 ( .A(n7691), .B(P2_IR_REG_18__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U10061 ( .A1(n8016), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8015), 
        .B2(n12060), .ZN(n7692) );
  XNOR2_X1 U10062 ( .A(n13625), .B(n6809), .ZN(n8030) );
  NOR2_X1 U10063 ( .A1(n8021), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7694) );
  OR2_X1 U10064 ( .A1(n7695), .A2(n7694), .ZN(n13619) );
  INV_X1 U10065 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7698) );
  NAND2_X1 U10066 ( .A1(n7702), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7697) );
  INV_X1 U10067 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13620) );
  OR2_X1 U10068 ( .A1(n8248), .A2(n13620), .ZN(n7696) );
  OAI211_X1 U10069 ( .C1(n7736), .C2(n7698), .A(n7697), .B(n7696), .ZN(n7699)
         );
  INV_X1 U10070 ( .A(n7699), .ZN(n7700) );
  OAI21_X1 U10071 ( .B1(n13619), .B2(n8247), .A(n7700), .ZN(n13396) );
  AND2_X1 U10072 ( .A1(n13396), .A2(n11080), .ZN(n8031) );
  NAND2_X1 U10073 ( .A1(n8030), .A2(n8031), .ZN(n8034) );
  INV_X1 U10074 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10429) );
  INV_X1 U10075 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10075) );
  OR2_X1 U10076 ( .A1(n7736), .A2(n10075), .ZN(n7703) );
  NAND2_X1 U10077 ( .A1(n9002), .A2(n11080), .ZN(n7734) );
  XNOR2_X1 U10078 ( .A(n7708), .B(n7707), .ZN(n9947) );
  NAND2_X1 U10079 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n7709) );
  XNOR2_X1 U10080 ( .A(n7709), .B(P2_IR_REG_1__SCAN_IN), .ZN(n10150) );
  NAND2_X1 U10081 ( .A1(n8015), .A2(n10150), .ZN(n7710) );
  INV_X1 U10082 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10145) );
  NAND2_X1 U10083 ( .A1(n9945), .A2(SI_0_), .ZN(n7711) );
  NAND2_X1 U10084 ( .A1(n7711), .A2(n8285), .ZN(n7713) );
  NAND2_X1 U10085 ( .A1(n7713), .A2(n7712), .ZN(n13808) );
  AOI22_X1 U10086 ( .A1(n7722), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_IR_REG_30__SCAN_IN), .B2(P2_REG0_REG_0__SCAN_IN), .ZN(n7719) );
  INV_X1 U10087 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7716) );
  NAND2_X1 U10088 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n7715) );
  OAI21_X1 U10089 ( .B1(n7716), .B2(P2_IR_REG_30__SCAN_IN), .A(n7715), .ZN(
        n7717) );
  NAND2_X1 U10090 ( .A1(n7714), .A2(n7717), .ZN(n7718) );
  OAI21_X1 U10091 ( .B1(n7714), .B2(n7719), .A(n7718), .ZN(n7721) );
  NAND2_X1 U10092 ( .A1(n7721), .A2(n7720), .ZN(n7731) );
  AOI22_X1 U10093 ( .A1(n7722), .A2(P2_REG3_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(P2_IR_REG_30__SCAN_IN), .ZN(n7727) );
  INV_X1 U10094 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7724) );
  NAND2_X1 U10095 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(P2_REG3_REG_0__SCAN_IN), 
        .ZN(n7723) );
  OAI21_X1 U10096 ( .B1(n7724), .B2(P2_IR_REG_30__SCAN_IN), .A(n7723), .ZN(
        n7725) );
  NAND2_X1 U10097 ( .A1(n7714), .A2(n7725), .ZN(n7726) );
  OAI21_X1 U10098 ( .B1(n7714), .B2(n7727), .A(n7726), .ZN(n7729) );
  NAND2_X1 U10099 ( .A1(n7729), .A2(n7728), .ZN(n7730) );
  NAND2_X1 U10100 ( .A1(n10421), .A2(n10323), .ZN(n9917) );
  OR2_X1 U10101 ( .A1(n9917), .A2(n11674), .ZN(n10419) );
  NAND2_X1 U10102 ( .A1(n8159), .A2(n8994), .ZN(n7732) );
  INV_X1 U10103 ( .A(n10434), .ZN(n7733) );
  NAND2_X1 U10104 ( .A1(n7734), .A2(n7733), .ZN(n7735) );
  NAND2_X1 U10105 ( .A1(n7702), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7740) );
  INV_X1 U10106 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10440) );
  OR2_X1 U10107 ( .A1(n8247), .A2(n10440), .ZN(n7739) );
  INV_X1 U10108 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10061) );
  OR2_X1 U10109 ( .A1(n8248), .A2(n10061), .ZN(n7738) );
  INV_X1 U10110 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10074) );
  OR2_X1 U10111 ( .A1(n7736), .A2(n10074), .ZN(n7737) );
  NAND2_X1 U10112 ( .A1(n13311), .A2(n11080), .ZN(n7749) );
  XNOR2_X1 U10113 ( .A(n7742), .B(n7741), .ZN(n9942) );
  NAND2_X1 U10114 ( .A1(n9942), .A2(n7753), .ZN(n7746) );
  INV_X1 U10115 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13786) );
  OR2_X1 U10116 ( .A1(n7743), .A2(n13786), .ZN(n7744) );
  XNOR2_X1 U10117 ( .A(n7744), .B(P2_IR_REG_2__SCAN_IN), .ZN(n13323) );
  NAND2_X1 U10118 ( .A1(n8015), .A2(n13323), .ZN(n7745) );
  XNOR2_X1 U10119 ( .A(n10915), .B(n8181), .ZN(n7747) );
  XNOR2_X1 U10120 ( .A(n7749), .B(n7747), .ZN(n10436) );
  INV_X1 U10121 ( .A(n7747), .ZN(n7748) );
  NAND2_X1 U10122 ( .A1(n7749), .A2(n7748), .ZN(n7750) );
  XNOR2_X1 U10123 ( .A(n7752), .B(n7751), .ZN(n9948) );
  NAND2_X1 U10124 ( .A1(n9948), .A2(n9209), .ZN(n7756) );
  OR2_X1 U10125 ( .A1(n7768), .A2(n13786), .ZN(n7754) );
  XNOR2_X1 U10126 ( .A(n7754), .B(P2_IR_REG_3__SCAN_IN), .ZN(n10081) );
  XNOR2_X1 U10127 ( .A(n10953), .B(n8181), .ZN(n7761) );
  NAND2_X1 U10128 ( .A1(n7702), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7760) );
  OR2_X1 U10129 ( .A1(n8247), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7759) );
  INV_X1 U10130 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10063) );
  OR2_X1 U10131 ( .A1(n8248), .A2(n10063), .ZN(n7758) );
  INV_X1 U10132 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10073) );
  OR2_X1 U10133 ( .A1(n7736), .A2(n10073), .ZN(n7757) );
  NAND4_X1 U10134 ( .A1(n7760), .A2(n7759), .A3(n7758), .A4(n7757), .ZN(n13310) );
  AND2_X1 U10135 ( .A1(n13310), .A2(n11080), .ZN(n7762) );
  NAND2_X1 U10136 ( .A1(n7761), .A2(n7762), .ZN(n7781) );
  INV_X1 U10137 ( .A(n7761), .ZN(n10528) );
  INV_X1 U10138 ( .A(n7762), .ZN(n7763) );
  NAND2_X1 U10139 ( .A1(n10528), .A2(n7763), .ZN(n7764) );
  NAND2_X1 U10140 ( .A1(n7781), .A2(n7764), .ZN(n10588) );
  XNOR2_X1 U10141 ( .A(n7765), .B(n7766), .ZN(n9953) );
  NAND2_X1 U10142 ( .A1(n9953), .A2(n9209), .ZN(n7771) );
  NAND2_X1 U10143 ( .A1(n7768), .A2(n7767), .ZN(n7787) );
  NAND2_X1 U10144 ( .A1(n7787), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7769) );
  XNOR2_X1 U10145 ( .A(n7769), .B(P2_IR_REG_4__SCAN_IN), .ZN(n10126) );
  AOI22_X1 U10146 ( .A1(n8016), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8015), .B2(
        n10126), .ZN(n7770) );
  XNOR2_X1 U10147 ( .A(n14984), .B(n8181), .ZN(n7783) );
  NAND2_X1 U10148 ( .A1(n9210), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7780) );
  INV_X1 U10149 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7772) );
  OR2_X1 U10150 ( .A1(n8246), .A2(n7772), .ZN(n7779) );
  INV_X1 U10151 ( .A(n7792), .ZN(n7776) );
  INV_X1 U10152 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7774) );
  INV_X1 U10153 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7773) );
  NAND2_X1 U10154 ( .A1(n7774), .A2(n7773), .ZN(n7775) );
  NAND2_X1 U10155 ( .A1(n7776), .A2(n7775), .ZN(n11011) );
  OR2_X1 U10156 ( .A1(n8247), .A2(n11011), .ZN(n7778) );
  INV_X1 U10157 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11007) );
  OR2_X1 U10158 ( .A1(n8248), .A2(n11007), .ZN(n7777) );
  NAND2_X1 U10159 ( .A1(n13309), .A2(n11080), .ZN(n7784) );
  XNOR2_X1 U10160 ( .A(n7783), .B(n7784), .ZN(n10527) );
  INV_X1 U10161 ( .A(n7783), .ZN(n10656) );
  XNOR2_X1 U10162 ( .A(n7785), .B(n7786), .ZN(n9951) );
  NAND2_X1 U10163 ( .A1(n9951), .A2(n9209), .ZN(n7790) );
  NAND2_X1 U10164 ( .A1(n7803), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7788) );
  XNOR2_X1 U10165 ( .A(n7788), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U10166 ( .A1(n8016), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8015), .B2(
        n10332), .ZN(n7789) );
  NAND2_X1 U10167 ( .A1(n7790), .A2(n7789), .ZN(n11071) );
  XNOR2_X1 U10168 ( .A(n11071), .B(n8181), .ZN(n7797) );
  NAND2_X1 U10169 ( .A1(n9210), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7796) );
  INV_X1 U10170 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7791) );
  OR2_X1 U10171 ( .A1(n8246), .A2(n7791), .ZN(n7795) );
  OAI21_X1 U10172 ( .B1(n7792), .B2(P2_REG3_REG_5__SCAN_IN), .A(n7811), .ZN(
        n11060) );
  OR2_X1 U10173 ( .A1(n8247), .A2(n11060), .ZN(n7794) );
  INV_X1 U10174 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11059) );
  OR2_X1 U10175 ( .A1(n8248), .A2(n11059), .ZN(n7793) );
  NAND4_X1 U10176 ( .A1(n7796), .A2(n7795), .A3(n7794), .A4(n7793), .ZN(n13308) );
  NAND2_X1 U10177 ( .A1(n13308), .A2(n11080), .ZN(n7798) );
  XNOR2_X1 U10178 ( .A(n7797), .B(n7798), .ZN(n10657) );
  INV_X1 U10179 ( .A(n7797), .ZN(n7799) );
  NAND2_X1 U10180 ( .A1(n7799), .A2(n7798), .ZN(n7800) );
  XNOR2_X1 U10181 ( .A(n7801), .B(n7802), .ZN(n9964) );
  NAND2_X1 U10182 ( .A1(n9964), .A2(n9209), .ZN(n7808) );
  INV_X1 U10183 ( .A(n7803), .ZN(n7805) );
  NAND2_X1 U10184 ( .A1(n7805), .A2(n7804), .ZN(n7825) );
  NAND2_X1 U10185 ( .A1(n7825), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7806) );
  XNOR2_X1 U10186 ( .A(n7806), .B(P2_IR_REG_6__SCAN_IN), .ZN(n13335) );
  AOI22_X1 U10187 ( .A1(n8016), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8015), .B2(
        n13335), .ZN(n7807) );
  NAND2_X1 U10188 ( .A1(n7808), .A2(n7807), .ZN(n14991) );
  XNOR2_X1 U10189 ( .A(n14991), .B(n8181), .ZN(n7817) );
  NAND2_X1 U10190 ( .A1(n9210), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7816) );
  INV_X1 U10191 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7809) );
  OR2_X1 U10192 ( .A1(n8246), .A2(n7809), .ZN(n7815) );
  AND2_X1 U10193 ( .A1(n7811), .A2(n7810), .ZN(n7812) );
  OR2_X1 U10194 ( .A1(n7812), .A2(n7832), .ZN(n11083) );
  OR2_X1 U10195 ( .A1(n8247), .A2(n11083), .ZN(n7814) );
  INV_X1 U10196 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11078) );
  OR2_X1 U10197 ( .A1(n8248), .A2(n11078), .ZN(n7813) );
  NAND4_X1 U10198 ( .A1(n7816), .A2(n7815), .A3(n7814), .A4(n7813), .ZN(n13307) );
  AND2_X1 U10199 ( .A1(n13307), .A2(n11080), .ZN(n7818) );
  NAND2_X1 U10200 ( .A1(n7817), .A2(n7818), .ZN(n7822) );
  INV_X1 U10201 ( .A(n7817), .ZN(n10877) );
  INV_X1 U10202 ( .A(n7818), .ZN(n7819) );
  NAND2_X1 U10203 ( .A1(n10877), .A2(n7819), .ZN(n7820) );
  NAND2_X1 U10204 ( .A1(n7822), .A2(n7820), .ZN(n10792) );
  INV_X1 U10205 ( .A(n10792), .ZN(n7821) );
  NAND2_X1 U10206 ( .A1(n10876), .A2(n7822), .ZN(n7838) );
  NAND2_X1 U10207 ( .A1(n9969), .A2(n9209), .ZN(n7830) );
  INV_X1 U10208 ( .A(n7825), .ZN(n7827) );
  INV_X1 U10209 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7826) );
  NAND2_X1 U10210 ( .A1(n7827), .A2(n7826), .ZN(n7846) );
  NAND2_X1 U10211 ( .A1(n7846), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7828) );
  XNOR2_X1 U10212 ( .A(n7828), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10134) );
  AOI22_X1 U10213 ( .A1(n8016), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8015), .B2(
        n10134), .ZN(n7829) );
  NAND2_X1 U10214 ( .A1(n7830), .A2(n7829), .ZN(n14954) );
  XNOR2_X1 U10215 ( .A(n14954), .B(n6809), .ZN(n7841) );
  NAND2_X1 U10216 ( .A1(n9210), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7837) );
  INV_X1 U10217 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7831) );
  OR2_X1 U10218 ( .A1(n8246), .A2(n7831), .ZN(n7836) );
  OR2_X1 U10219 ( .A1(n7832), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7833) );
  NAND2_X1 U10220 ( .A1(n7852), .A2(n7833), .ZN(n14951) );
  OR2_X1 U10221 ( .A1(n8247), .A2(n14951), .ZN(n7835) );
  OR2_X1 U10222 ( .A1(n8248), .A2(n10064), .ZN(n7834) );
  NAND4_X1 U10223 ( .A1(n7837), .A2(n7836), .A3(n7835), .A4(n7834), .ZN(n13306) );
  NAND2_X1 U10224 ( .A1(n13306), .A2(n11080), .ZN(n7839) );
  XNOR2_X1 U10225 ( .A(n7841), .B(n7839), .ZN(n10874) );
  NAND2_X1 U10226 ( .A1(n7838), .A2(n10874), .ZN(n10878) );
  INV_X1 U10227 ( .A(n7839), .ZN(n7840) );
  NAND2_X1 U10228 ( .A1(n7841), .A2(n7840), .ZN(n7842) );
  XNOR2_X1 U10229 ( .A(n7843), .B(SI_8_), .ZN(n7844) );
  XNOR2_X1 U10230 ( .A(n7845), .B(n7844), .ZN(n10000) );
  NAND2_X1 U10231 ( .A1(n10000), .A2(n9209), .ZN(n7849) );
  NAND2_X1 U10232 ( .A1(n7865), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7847) );
  XNOR2_X1 U10233 ( .A(n7847), .B(P2_IR_REG_8__SCAN_IN), .ZN(n13352) );
  AOI22_X1 U10234 ( .A1(n8016), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8015), .B2(
        n13352), .ZN(n7848) );
  NAND2_X1 U10235 ( .A1(n7849), .A2(n7848), .ZN(n11437) );
  XNOR2_X1 U10236 ( .A(n11437), .B(n8159), .ZN(n11214) );
  NAND2_X1 U10237 ( .A1(n9210), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7857) );
  INV_X1 U10238 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7850) );
  OR2_X1 U10239 ( .A1(n8246), .A2(n7850), .ZN(n7856) );
  NAND2_X1 U10240 ( .A1(n7852), .A2(n7851), .ZN(n7853) );
  NAND2_X1 U10241 ( .A1(n7874), .A2(n7853), .ZN(n11257) );
  OR2_X1 U10242 ( .A1(n8247), .A2(n11257), .ZN(n7855) );
  INV_X1 U10243 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11253) );
  OR2_X1 U10244 ( .A1(n8248), .A2(n11253), .ZN(n7854) );
  NAND4_X1 U10245 ( .A1(n7857), .A2(n7856), .A3(n7855), .A4(n7854), .ZN(n13305) );
  NAND2_X1 U10246 ( .A1(n13305), .A2(n11080), .ZN(n7859) );
  NAND2_X1 U10247 ( .A1(n11214), .A2(n7859), .ZN(n7858) );
  NAND2_X1 U10248 ( .A1(n11220), .A2(n7858), .ZN(n11219) );
  INV_X1 U10249 ( .A(n11214), .ZN(n7861) );
  INV_X1 U10250 ( .A(n7859), .ZN(n7860) );
  NAND2_X1 U10251 ( .A1(n7861), .A2(n7860), .ZN(n11222) );
  INV_X1 U10252 ( .A(n7862), .ZN(n7863) );
  XNOR2_X1 U10253 ( .A(n7864), .B(n7863), .ZN(n10056) );
  NAND2_X1 U10254 ( .A1(n10056), .A2(n9209), .ZN(n7872) );
  INV_X1 U10255 ( .A(n7865), .ZN(n7867) );
  INV_X1 U10256 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7866) );
  NAND2_X1 U10257 ( .A1(n7867), .A2(n7866), .ZN(n7869) );
  NAND2_X1 U10258 ( .A1(n7869), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7868) );
  MUX2_X1 U10259 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7868), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n7870) );
  AOI22_X1 U10260 ( .A1(n10108), .A2(n8015), .B1(n8016), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n7871) );
  XNOR2_X1 U10261 ( .A(n11554), .B(n8159), .ZN(n7881) );
  NAND2_X1 U10262 ( .A1(n9210), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7879) );
  INV_X1 U10263 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7873) );
  OR2_X1 U10264 ( .A1(n8246), .A2(n7873), .ZN(n7878) );
  AND2_X1 U10265 ( .A1(n7874), .A2(n11266), .ZN(n7875) );
  OR2_X1 U10266 ( .A1(n7875), .A2(n7890), .ZN(n11397) );
  OR2_X1 U10267 ( .A1(n8247), .A2(n11397), .ZN(n7877) );
  INV_X1 U10268 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11398) );
  OR2_X1 U10269 ( .A1(n8248), .A2(n11398), .ZN(n7876) );
  NAND4_X1 U10270 ( .A1(n7879), .A2(n7878), .A3(n7877), .A4(n7876), .ZN(n13304) );
  NAND2_X1 U10271 ( .A1(n13304), .A2(n11080), .ZN(n7880) );
  XNOR2_X1 U10272 ( .A(n7881), .B(n7880), .ZN(n11263) );
  NAND2_X1 U10273 ( .A1(n7881), .A2(n7880), .ZN(n7882) );
  OR2_X1 U10274 ( .A1(n7884), .A2(n7883), .ZN(n7885) );
  NAND2_X1 U10275 ( .A1(n10221), .A2(n9209), .ZN(n7889) );
  NAND2_X1 U10276 ( .A1(n7904), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7887) );
  XNOR2_X1 U10277 ( .A(n7887), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10365) );
  AOI22_X1 U10278 ( .A1(n10365), .A2(n8015), .B1(n8016), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n7888) );
  XNOR2_X1 U10279 ( .A(n11663), .B(n6809), .ZN(n7896) );
  NAND2_X1 U10280 ( .A1(n7702), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7895) );
  INV_X1 U10281 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10364) );
  OR2_X1 U10282 ( .A1(n7736), .A2(n10364), .ZN(n7894) );
  NOR2_X1 U10283 ( .A1(n7890), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7891) );
  OR2_X1 U10284 ( .A1(n7909), .A2(n7891), .ZN(n11525) );
  OR2_X1 U10285 ( .A1(n8247), .A2(n11525), .ZN(n7893) );
  INV_X1 U10286 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10356) );
  OR2_X1 U10287 ( .A1(n8248), .A2(n10356), .ZN(n7892) );
  NAND4_X1 U10288 ( .A1(n7895), .A2(n7894), .A3(n7893), .A4(n7892), .ZN(n13303) );
  AND2_X1 U10289 ( .A1(n13303), .A2(n11080), .ZN(n7897) );
  NAND2_X1 U10290 ( .A1(n7896), .A2(n7897), .ZN(n7901) );
  INV_X1 U10291 ( .A(n7896), .ZN(n11502) );
  INV_X1 U10292 ( .A(n7897), .ZN(n7898) );
  NAND2_X1 U10293 ( .A1(n11502), .A2(n7898), .ZN(n7899) );
  NAND2_X1 U10294 ( .A1(n7901), .A2(n7899), .ZN(n11409) );
  NAND2_X1 U10295 ( .A1(n10375), .A2(n9209), .ZN(n7907) );
  OAI21_X1 U10296 ( .B1(n7904), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7905) );
  XNOR2_X1 U10297 ( .A(n7905), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10702) );
  AOI22_X1 U10298 ( .A1(n10702), .A2(n8015), .B1(n8016), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n7906) );
  XNOR2_X1 U10299 ( .A(n11816), .B(n6809), .ZN(n7915) );
  NAND2_X1 U10300 ( .A1(n9210), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7914) );
  INV_X1 U10301 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7908) );
  OR2_X1 U10302 ( .A1(n8246), .A2(n7908), .ZN(n7913) );
  OR2_X1 U10303 ( .A1(n7909), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7910) );
  NAND2_X1 U10304 ( .A1(n7926), .A2(n7910), .ZN(n11676) );
  OR2_X1 U10305 ( .A1(n8247), .A2(n11676), .ZN(n7912) );
  INV_X1 U10306 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11677) );
  OR2_X1 U10307 ( .A1(n8248), .A2(n11677), .ZN(n7911) );
  NAND4_X1 U10308 ( .A1(n7914), .A2(n7913), .A3(n7912), .A4(n7911), .ZN(n13302) );
  AND2_X1 U10309 ( .A1(n13302), .A2(n11080), .ZN(n7916) );
  NAND2_X1 U10310 ( .A1(n7915), .A2(n7916), .ZN(n7932) );
  INV_X1 U10311 ( .A(n7915), .ZN(n13222) );
  INV_X1 U10312 ( .A(n7916), .ZN(n7917) );
  NAND2_X1 U10313 ( .A1(n13222), .A2(n7917), .ZN(n7918) );
  AND2_X1 U10314 ( .A1(n7932), .A2(n7918), .ZN(n11498) );
  NAND2_X1 U10315 ( .A1(n7919), .A2(n11498), .ZN(n11503) );
  XNOR2_X1 U10316 ( .A(n7921), .B(n7920), .ZN(n10424) );
  NAND2_X1 U10317 ( .A1(n10424), .A2(n9209), .ZN(n7924) );
  XNOR2_X1 U10318 ( .A(n7922), .B(P2_IR_REG_12__SCAN_IN), .ZN(n13370) );
  AOI22_X1 U10319 ( .A1(n8016), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8015), 
        .B2(n13370), .ZN(n7923) );
  XNOR2_X1 U10320 ( .A(n13221), .B(n6809), .ZN(n7934) );
  NAND2_X1 U10321 ( .A1(n7702), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7931) );
  NAND2_X1 U10322 ( .A1(n7926), .A2(n7925), .ZN(n7927) );
  NAND2_X1 U10323 ( .A1(n7944), .A2(n7927), .ZN(n13219) );
  OR2_X1 U10324 ( .A1(n8247), .A2(n13219), .ZN(n7930) );
  OR2_X1 U10325 ( .A1(n8248), .A2(n11824), .ZN(n7929) );
  INV_X1 U10326 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10703) );
  OR2_X1 U10327 ( .A1(n7736), .A2(n10703), .ZN(n7928) );
  NAND4_X1 U10328 ( .A1(n7931), .A2(n7930), .A3(n7929), .A4(n7928), .ZN(n13301) );
  NAND2_X1 U10329 ( .A1(n13301), .A2(n11080), .ZN(n7935) );
  XNOR2_X1 U10330 ( .A(n7934), .B(n7935), .ZN(n13223) );
  AND2_X1 U10331 ( .A1(n13223), .A2(n7932), .ZN(n7933) );
  INV_X1 U10332 ( .A(n7934), .ZN(n7936) );
  NAND2_X1 U10333 ( .A1(n7936), .A2(n7935), .ZN(n7937) );
  XNOR2_X1 U10334 ( .A(n7939), .B(n7938), .ZN(n10612) );
  NAND2_X1 U10335 ( .A1(n10612), .A2(n9209), .ZN(n7942) );
  NAND2_X1 U10336 ( .A1(n7963), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7940) );
  XNOR2_X1 U10337 ( .A(n7940), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U10338 ( .A1(n8016), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8015), 
        .B2(n11700), .ZN(n7941) );
  XNOR2_X1 U10339 ( .A(n14868), .B(n6809), .ZN(n11801) );
  NAND2_X1 U10340 ( .A1(n7944), .A2(n7943), .ZN(n7945) );
  NAND2_X1 U10341 ( .A1(n7967), .A2(n7945), .ZN(n14871) );
  INV_X1 U10342 ( .A(n14871), .ZN(n7946) );
  NAND2_X1 U10343 ( .A1(n7947), .A2(n7946), .ZN(n7953) );
  INV_X1 U10344 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7948) );
  OR2_X1 U10345 ( .A1(n8246), .A2(n7948), .ZN(n7952) );
  INV_X1 U10346 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7949) );
  OR2_X1 U10347 ( .A1(n8248), .A2(n7949), .ZN(n7951) );
  INV_X1 U10348 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11711) );
  OR2_X1 U10349 ( .A1(n7736), .A2(n11711), .ZN(n7950) );
  NAND4_X1 U10350 ( .A1(n7953), .A2(n7952), .A3(n7951), .A4(n7950), .ZN(n13300) );
  AND2_X1 U10351 ( .A1(n13300), .A2(n11080), .ZN(n7954) );
  NAND2_X1 U10352 ( .A1(n11801), .A2(n7954), .ZN(n7973) );
  INV_X1 U10353 ( .A(n11801), .ZN(n7956) );
  INV_X1 U10354 ( .A(n7954), .ZN(n7955) );
  NAND2_X1 U10355 ( .A1(n7956), .A2(n7955), .ZN(n7957) );
  AND2_X1 U10356 ( .A1(n7973), .A2(n7957), .ZN(n14863) );
  NAND2_X1 U10357 ( .A1(n7959), .A2(n7958), .ZN(n7960) );
  NAND2_X1 U10358 ( .A1(n7961), .A2(n7960), .ZN(n10790) );
  OR2_X1 U10359 ( .A1(n10790), .A2(n7962), .ZN(n7966) );
  NAND2_X1 U10360 ( .A1(n7981), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7964) );
  XNOR2_X1 U10361 ( .A(n7964), .B(P2_IR_REG_14__SCAN_IN), .ZN(n14905) );
  AOI22_X1 U10362 ( .A1(n8016), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8015), 
        .B2(n14905), .ZN(n7965) );
  XNOR2_X1 U10363 ( .A(n13744), .B(n6809), .ZN(n7975) );
  AND2_X1 U10364 ( .A1(n7967), .A2(n11807), .ZN(n7968) );
  OR2_X1 U10365 ( .A1(n7968), .A2(n7987), .ZN(n12022) );
  INV_X1 U10366 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11712) );
  OR2_X1 U10367 ( .A1(n7736), .A2(n11712), .ZN(n7970) );
  INV_X1 U10368 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n12197) );
  OR2_X1 U10369 ( .A1(n8246), .A2(n12197), .ZN(n7969) );
  AND2_X1 U10370 ( .A1(n7970), .A2(n7969), .ZN(n7972) );
  NAND2_X1 U10371 ( .A1(n7701), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7971) );
  OAI211_X1 U10372 ( .C1(n12022), .C2(n8247), .A(n7972), .B(n7971), .ZN(n13299) );
  NAND2_X1 U10373 ( .A1(n13299), .A2(n11080), .ZN(n7976) );
  XNOR2_X1 U10374 ( .A(n7975), .B(n7976), .ZN(n11803) );
  INV_X1 U10375 ( .A(n7975), .ZN(n7977) );
  NAND2_X1 U10376 ( .A1(n7977), .A2(n7976), .ZN(n7978) );
  NAND2_X1 U10377 ( .A1(n11812), .A2(n7978), .ZN(n7994) );
  XNOR2_X1 U10378 ( .A(n7980), .B(n7979), .ZN(n10949) );
  NAND2_X1 U10379 ( .A1(n10949), .A2(n9209), .ZN(n7986) );
  INV_X1 U10380 ( .A(n7981), .ZN(n7983) );
  NAND2_X1 U10381 ( .A1(n7983), .A2(n7982), .ZN(n7998) );
  NAND2_X1 U10382 ( .A1(n7998), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7984) );
  XNOR2_X1 U10383 ( .A(n7984), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14915) );
  AOI22_X1 U10384 ( .A1(n8016), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n14915), 
        .B2(n8015), .ZN(n7985) );
  XNOR2_X1 U10385 ( .A(n13782), .B(n6809), .ZN(n7992) );
  OR2_X1 U10386 ( .A1(n7987), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7988) );
  NAND2_X1 U10387 ( .A1(n8002), .A2(n7988), .ZN(n12170) );
  AOI22_X1 U10388 ( .A1(n9210), .A2(P2_REG1_REG_15__SCAN_IN), .B1(n7702), .B2(
        P2_REG0_REG_15__SCAN_IN), .ZN(n7990) );
  INV_X1 U10389 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n12175) );
  OR2_X1 U10390 ( .A1(n8248), .A2(n12175), .ZN(n7989) );
  OAI211_X1 U10391 ( .C1(n12170), .C2(n8247), .A(n7990), .B(n7989), .ZN(n13298) );
  AND2_X1 U10392 ( .A1(n13298), .A2(n11080), .ZN(n7991) );
  INV_X1 U10393 ( .A(n7992), .ZN(n7993) );
  OR2_X1 U10394 ( .A1(n7994), .A2(n7993), .ZN(n7995) );
  XNOR2_X1 U10395 ( .A(n7997), .B(n7996), .ZN(n11170) );
  NAND2_X1 U10396 ( .A1(n11170), .A2(n9209), .ZN(n8001) );
  OAI21_X1 U10397 ( .B1(n7998), .B2(P2_IR_REG_15__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7999) );
  XNOR2_X1 U10398 ( .A(n7999), .B(P2_IR_REG_16__SCAN_IN), .ZN(n14924) );
  AOI22_X1 U10399 ( .A1(n8016), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n14924), 
        .B2(n8015), .ZN(n8000) );
  XNOR2_X1 U10400 ( .A(n13419), .B(n8159), .ZN(n13242) );
  NAND2_X1 U10401 ( .A1(n8002), .A2(n13232), .ZN(n8003) );
  NAND2_X1 U10402 ( .A1(n8020), .A2(n8003), .ZN(n13231) );
  AOI22_X1 U10403 ( .A1(n9210), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n7702), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n8005) );
  INV_X1 U10404 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12207) );
  OR2_X1 U10405 ( .A1(n8248), .A2(n12207), .ZN(n8004) );
  OAI211_X1 U10406 ( .C1(n13231), .C2(n8247), .A(n8005), .B(n8004), .ZN(n13391) );
  NAND2_X1 U10407 ( .A1(n13391), .A2(n11080), .ZN(n8006) );
  XNOR2_X1 U10408 ( .A(n13242), .B(n8006), .ZN(n13230) );
  NAND2_X1 U10409 ( .A1(n13242), .A2(n8006), .ZN(n8007) );
  NAND2_X1 U10410 ( .A1(n13245), .A2(n8007), .ZN(n8025) );
  XNOR2_X1 U10411 ( .A(n8008), .B(SI_17_), .ZN(n8009) );
  XNOR2_X1 U10412 ( .A(n8010), .B(n8009), .ZN(n11345) );
  NAND2_X1 U10413 ( .A1(n11345), .A2(n9209), .ZN(n8018) );
  NAND2_X1 U10414 ( .A1(n8011), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8012) );
  MUX2_X1 U10415 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8012), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8014) );
  AOI22_X1 U10416 ( .A1(n8016), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8015), 
        .B2(n14937), .ZN(n8017) );
  XNOR2_X1 U10417 ( .A(n13727), .B(n6809), .ZN(n8026) );
  AND2_X1 U10418 ( .A1(n8020), .A2(n8019), .ZN(n8022) );
  OR2_X1 U10419 ( .A1(n8022), .A2(n8021), .ZN(n13636) );
  AOI22_X1 U10420 ( .A1(n7702), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n7701), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n8024) );
  INV_X1 U10421 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11718) );
  OR2_X1 U10422 ( .A1(n7736), .A2(n11718), .ZN(n8023) );
  OAI211_X1 U10423 ( .C1(n13636), .C2(n8247), .A(n8024), .B(n8023), .ZN(n13394) );
  NAND2_X1 U10424 ( .A1(n13394), .A2(n11080), .ZN(n8027) );
  XNOR2_X1 U10425 ( .A(n8026), .B(n8027), .ZN(n13241) );
  INV_X1 U10426 ( .A(n8026), .ZN(n8028) );
  NAND2_X1 U10427 ( .A1(n8028), .A2(n8027), .ZN(n8029) );
  INV_X1 U10428 ( .A(n8030), .ZN(n13199) );
  INV_X1 U10429 ( .A(n8031), .ZN(n8032) );
  NAND2_X1 U10430 ( .A1(n13199), .A2(n8032), .ZN(n8033) );
  NAND2_X1 U10431 ( .A1(n8034), .A2(n8033), .ZN(n13270) );
  INV_X1 U10432 ( .A(n8035), .ZN(n13262) );
  NAND2_X1 U10433 ( .A1(n13262), .A2(n8036), .ZN(n8047) );
  NOR2_X1 U10434 ( .A1(n8037), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8038) );
  OR2_X1 U10435 ( .A1(n8039), .A2(n8038), .ZN(n13582) );
  INV_X1 U10436 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n15371) );
  NAND2_X1 U10437 ( .A1(n9210), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8042) );
  INV_X1 U10438 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8040) );
  OR2_X1 U10439 ( .A1(n8248), .A2(n8040), .ZN(n8041) );
  OAI211_X1 U10440 ( .C1(n8246), .C2(n15371), .A(n8042), .B(n8041), .ZN(n8043)
         );
  INV_X1 U10441 ( .A(n8043), .ZN(n8044) );
  OAI21_X1 U10442 ( .B1(n13582), .B2(n8247), .A(n8044), .ZN(n13401) );
  NAND2_X1 U10443 ( .A1(n13401), .A2(n11080), .ZN(n8049) );
  OR2_X1 U10444 ( .A1(n9207), .A2(n11940), .ZN(n8046) );
  INV_X1 U10445 ( .A(n8048), .ZN(n8050) );
  XNOR2_X1 U10446 ( .A(n8051), .B(n8052), .ZN(n13211) );
  INV_X1 U10447 ( .A(n8056), .ZN(n8053) );
  NAND2_X1 U10448 ( .A1(n8053), .A2(n15362), .ZN(n8057) );
  OAI21_X1 U10449 ( .B1(SI_20_), .B2(n8054), .A(n8057), .ZN(n8060) );
  INV_X1 U10450 ( .A(SI_20_), .ZN(n10891) );
  NOR2_X1 U10451 ( .A1(n8055), .A2(n10891), .ZN(n8058) );
  AOI22_X1 U10452 ( .A1(n8058), .A2(n8057), .B1(n8056), .B2(SI_21_), .ZN(n8059) );
  MUX2_X1 U10453 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9945), .Z(n8075) );
  XNOR2_X1 U10454 ( .A(n9682), .B(n8075), .ZN(n12369) );
  NAND2_X1 U10455 ( .A1(n12369), .A2(n9209), .ZN(n8063) );
  INV_X1 U10456 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12371) );
  OR2_X1 U10457 ( .A1(n9207), .A2(n12371), .ZN(n8062) );
  NAND2_X2 U10458 ( .A1(n8063), .A2(n8062), .ZN(n13548) );
  XNOR2_X1 U10459 ( .A(n13548), .B(n6809), .ZN(n8073) );
  XNOR2_X1 U10460 ( .A(n8072), .B(n8073), .ZN(n12295) );
  NAND2_X1 U10461 ( .A1(n7702), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8070) );
  INV_X1 U10462 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n13702) );
  OR2_X1 U10463 ( .A1(n7736), .A2(n13702), .ZN(n8069) );
  INV_X1 U10464 ( .A(n8064), .ZN(n8066) );
  INV_X1 U10465 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n12297) );
  INV_X1 U10466 ( .A(n8084), .ZN(n8065) );
  OAI21_X1 U10467 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(n8066), .A(n8065), .ZN(
        n13549) );
  OR2_X1 U10468 ( .A1(n8247), .A2(n13549), .ZN(n8068) );
  INV_X1 U10469 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13550) );
  OR2_X1 U10470 ( .A1(n8248), .A2(n13550), .ZN(n8067) );
  NAND4_X1 U10471 ( .A1(n8070), .A2(n8069), .A3(n8068), .A4(n8067), .ZN(n13406) );
  INV_X1 U10472 ( .A(n13406), .ZN(n13563) );
  OR2_X1 U10473 ( .A1(n13563), .A2(n11674), .ZN(n8071) );
  AND2_X1 U10474 ( .A1(n8073), .A2(n8072), .ZN(n8074) );
  INV_X1 U10475 ( .A(n8075), .ZN(n8078) );
  NAND2_X1 U10476 ( .A1(n8076), .A2(SI_22_), .ZN(n8077) );
  OAI21_X2 U10477 ( .B1(n8079), .B2(n8078), .A(n8077), .ZN(n8093) );
  MUX2_X1 U10478 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9945), .Z(n8092) );
  XNOR2_X1 U10479 ( .A(n8091), .B(SI_23_), .ZN(n12248) );
  NAND2_X1 U10480 ( .A1(n12248), .A2(n9209), .ZN(n8081) );
  OR2_X1 U10481 ( .A1(n9207), .A2(n12251), .ZN(n8080) );
  XNOR2_X1 U10482 ( .A(n13536), .B(n6809), .ZN(n8089) );
  INV_X1 U10483 ( .A(n8089), .ZN(n8082) );
  NAND2_X1 U10484 ( .A1(n9210), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8088) );
  INV_X1 U10485 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8083) );
  OR2_X1 U10486 ( .A1(n8246), .A2(n8083), .ZN(n8087) );
  NAND2_X1 U10487 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(n8084), .ZN(n8098) );
  OAI21_X1 U10488 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(n8084), .A(n8098), .ZN(
        n13542) );
  OR2_X1 U10489 ( .A1(n8247), .A2(n13542), .ZN(n8086) );
  INV_X1 U10490 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13535) );
  OR2_X1 U10491 ( .A1(n8248), .A2(n13535), .ZN(n8085) );
  NAND2_X1 U10492 ( .A1(n8093), .A2(n8092), .ZN(n8094) );
  MUX2_X1 U10493 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9945), .Z(n8125) );
  NAND2_X1 U10494 ( .A1(n9715), .A2(n9209), .ZN(n8096) );
  INV_X1 U10495 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13806) );
  OR2_X1 U10496 ( .A1(n9207), .A2(n13806), .ZN(n8095) );
  XNOR2_X1 U10497 ( .A(n13688), .B(n8159), .ZN(n12268) );
  NAND2_X1 U10498 ( .A1(n7702), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8104) );
  INV_X1 U10499 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8097) );
  OR2_X1 U10500 ( .A1(n7736), .A2(n8097), .ZN(n8103) );
  OAI21_X1 U10501 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n8099), .A(n8138), .ZN(
        n13252) );
  OR2_X1 U10502 ( .A1(n8247), .A2(n13252), .ZN(n8102) );
  INV_X1 U10503 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8100) );
  OR2_X1 U10504 ( .A1(n8248), .A2(n8100), .ZN(n8101) );
  NAND4_X1 U10505 ( .A1(n8104), .A2(n8103), .A3(n8102), .A4(n8101), .ZN(n13412) );
  NAND2_X1 U10506 ( .A1(n13412), .A2(n11080), .ZN(n8105) );
  NOR2_X1 U10507 ( .A1(n12268), .A2(n8105), .ZN(n8123) );
  AOI21_X1 U10508 ( .B1(n12268), .B2(n8105), .A(n8123), .ZN(n13251) );
  NAND2_X1 U10509 ( .A1(n8106), .A2(n8125), .ZN(n8108) );
  NAND2_X1 U10510 ( .A1(n8132), .A2(SI_24_), .ZN(n8107) );
  MUX2_X1 U10511 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n9945), .Z(n8109) );
  NAND2_X1 U10512 ( .A1(n8109), .A2(SI_25_), .ZN(n8128) );
  INV_X1 U10513 ( .A(n8109), .ZN(n8110) );
  INV_X1 U10514 ( .A(SI_25_), .ZN(n11695) );
  NAND2_X1 U10515 ( .A1(n8110), .A2(n11695), .ZN(n8126) );
  NAND2_X1 U10516 ( .A1(n8128), .A2(n8126), .ZN(n8111) );
  INV_X1 U10517 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13803) );
  OR2_X1 U10518 ( .A1(n9207), .A2(n13803), .ZN(n8113) );
  XNOR2_X1 U10519 ( .A(n13512), .B(n8159), .ZN(n8119) );
  NAND2_X1 U10520 ( .A1(n9210), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8118) );
  INV_X1 U10521 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8114) );
  OR2_X1 U10522 ( .A1(n8246), .A2(n8114), .ZN(n8117) );
  INV_X1 U10523 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n12274) );
  XNOR2_X1 U10524 ( .A(n8138), .B(n12274), .ZN(n13506) );
  OR2_X1 U10525 ( .A1(n8247), .A2(n13506), .ZN(n8116) );
  INV_X1 U10526 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13511) );
  OR2_X1 U10527 ( .A1(n8248), .A2(n13511), .ZN(n8115) );
  NOR2_X1 U10528 ( .A1(n13485), .A2(n11674), .ZN(n8120) );
  NAND2_X1 U10529 ( .A1(n8119), .A2(n8120), .ZN(n8146) );
  INV_X1 U10530 ( .A(n8119), .ZN(n13288) );
  INV_X1 U10531 ( .A(n8120), .ZN(n8121) );
  NAND2_X1 U10532 ( .A1(n13288), .A2(n8121), .ZN(n8122) );
  INV_X1 U10533 ( .A(SI_24_), .ZN(n11605) );
  INV_X1 U10534 ( .A(n8125), .ZN(n8124) );
  OAI21_X1 U10535 ( .B1(n11605), .B2(n8124), .A(n8128), .ZN(n8131) );
  NOR2_X1 U10536 ( .A1(n8125), .A2(SI_24_), .ZN(n8129) );
  INV_X1 U10537 ( .A(n8126), .ZN(n8127) );
  AOI21_X1 U10538 ( .B1(n8129), .B2(n8128), .A(n8127), .ZN(n8130) );
  OAI21_X2 U10539 ( .B1(n8132), .B2(n8131), .A(n8130), .ZN(n8152) );
  INV_X1 U10540 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14462) );
  INV_X1 U10541 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13799) );
  MUX2_X1 U10542 ( .A(n14462), .B(n13799), .S(n9945), .Z(n8151) );
  XNOR2_X1 U10543 ( .A(n8151), .B(SI_26_), .ZN(n8133) );
  XNOR2_X1 U10544 ( .A(n8152), .B(n8133), .ZN(n13798) );
  NAND2_X1 U10545 ( .A1(n13798), .A2(n9209), .ZN(n8135) );
  OR2_X1 U10546 ( .A1(n9207), .A2(n13799), .ZN(n8134) );
  XNOR2_X1 U10547 ( .A(n13495), .B(n6809), .ZN(n8149) );
  NAND2_X1 U10548 ( .A1(n9210), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8145) );
  INV_X1 U10549 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8136) );
  OR2_X1 U10550 ( .A1(n8246), .A2(n8136), .ZN(n8144) );
  INV_X1 U10551 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8137) );
  OAI21_X1 U10552 ( .B1(n8138), .B2(n12274), .A(n8137), .ZN(n8141) );
  INV_X1 U10553 ( .A(n8138), .ZN(n8140) );
  AND2_X1 U10554 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n8139) );
  NAND2_X1 U10555 ( .A1(n8140), .A2(n8139), .ZN(n8163) );
  NAND2_X1 U10556 ( .A1(n8141), .A2(n8163), .ZN(n13492) );
  OR2_X1 U10557 ( .A1(n8247), .A2(n13492), .ZN(n8143) );
  INV_X1 U10558 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13493) );
  OR2_X1 U10559 ( .A1(n8248), .A2(n13493), .ZN(n8142) );
  NAND4_X1 U10560 ( .A1(n8145), .A2(n8144), .A3(n8143), .A4(n8142), .ZN(n13438) );
  NAND2_X1 U10561 ( .A1(n13438), .A2(n11080), .ZN(n8147) );
  XNOR2_X1 U10562 ( .A(n8149), .B(n8147), .ZN(n13287) );
  INV_X1 U10563 ( .A(n8147), .ZN(n8148) );
  INV_X1 U10564 ( .A(SI_26_), .ZN(n11798) );
  NAND2_X1 U10565 ( .A1(n8152), .A2(n11798), .ZN(n8153) );
  NAND2_X1 U10566 ( .A1(n8154), .A2(n8153), .ZN(n8173) );
  MUX2_X1 U10567 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n9945), .Z(n8174) );
  INV_X1 U10568 ( .A(n8174), .ZN(n8155) );
  XNOR2_X1 U10569 ( .A(n8155), .B(SI_27_), .ZN(n8156) );
  XNOR2_X1 U10570 ( .A(n8173), .B(n8156), .ZN(n13795) );
  NAND2_X1 U10571 ( .A1(n13795), .A2(n9209), .ZN(n8158) );
  INV_X1 U10572 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13797) );
  OR2_X1 U10573 ( .A1(n9207), .A2(n13797), .ZN(n8157) );
  XNOR2_X1 U10574 ( .A(n13416), .B(n8159), .ZN(n8170) );
  NAND2_X1 U10575 ( .A1(n9210), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8168) );
  INV_X1 U10576 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8160) );
  OR2_X1 U10577 ( .A1(n8246), .A2(n8160), .ZN(n8167) );
  INV_X1 U10578 ( .A(n8163), .ZN(n8161) );
  NAND2_X1 U10579 ( .A1(n8161), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8183) );
  INV_X1 U10580 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8162) );
  NAND2_X1 U10581 ( .A1(n8163), .A2(n8162), .ZN(n8164) );
  NAND2_X1 U10582 ( .A1(n8183), .A2(n8164), .ZN(n13472) );
  OR2_X1 U10583 ( .A1(n8247), .A2(n13472), .ZN(n8166) );
  INV_X1 U10584 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13473) );
  OR2_X1 U10585 ( .A1(n8248), .A2(n13473), .ZN(n8165) );
  NOR2_X1 U10586 ( .A1(n13484), .A2(n11674), .ZN(n8169) );
  NAND2_X1 U10587 ( .A1(n8170), .A2(n8169), .ZN(n8171) );
  OAI21_X1 U10588 ( .B1(n8170), .B2(n8169), .A(n8171), .ZN(n13179) );
  NOR2_X1 U10589 ( .A1(n8174), .A2(SI_27_), .ZN(n8172) );
  NAND2_X1 U10590 ( .A1(n8174), .A2(SI_27_), .ZN(n8175) );
  INV_X1 U10591 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14458) );
  INV_X1 U10592 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8842) );
  MUX2_X1 U10593 ( .A(n14458), .B(n8842), .S(n9945), .Z(n8176) );
  INV_X1 U10594 ( .A(SI_28_), .ZN(n11978) );
  NAND2_X1 U10595 ( .A1(n8176), .A2(n11978), .ZN(n9174) );
  INV_X1 U10596 ( .A(n8176), .ZN(n8177) );
  NAND2_X1 U10597 ( .A1(n8177), .A2(SI_28_), .ZN(n8178) );
  NAND2_X1 U10598 ( .A1(n9174), .A2(n8178), .ZN(n9172) );
  NAND2_X1 U10599 ( .A1(n13790), .A2(n9209), .ZN(n8180) );
  OR2_X1 U10600 ( .A1(n9207), .A2(n8842), .ZN(n8179) );
  NAND2_X1 U10601 ( .A1(n7702), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8189) );
  INV_X1 U10602 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8182) );
  OR2_X1 U10603 ( .A1(n7736), .A2(n8182), .ZN(n8188) );
  INV_X1 U10604 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8254) );
  NAND2_X1 U10605 ( .A1(n8183), .A2(n8254), .ZN(n8184) );
  NAND2_X1 U10606 ( .A1(n13447), .A2(n8184), .ZN(n13460) );
  OR2_X1 U10607 ( .A1(n8247), .A2(n13460), .ZN(n8187) );
  INV_X1 U10608 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8185) );
  OR2_X1 U10609 ( .A1(n8248), .A2(n8185), .ZN(n8186) );
  NOR4_X1 U10610 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8193) );
  NOR4_X1 U10611 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8192) );
  NOR4_X1 U10612 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8191) );
  NOR4_X1 U10613 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8190) );
  NAND4_X1 U10614 ( .A1(n8193), .A2(n8192), .A3(n8191), .A4(n8190), .ZN(n8217)
         );
  NOR2_X1 U10615 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .ZN(
        n8197) );
  NOR4_X1 U10616 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n8196) );
  NOR4_X1 U10617 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8195) );
  NOR4_X1 U10618 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8194) );
  NAND4_X1 U10619 ( .A1(n8197), .A2(n8196), .A3(n8195), .A4(n8194), .ZN(n8216)
         );
  NAND2_X1 U10620 ( .A1(n8227), .A2(n8199), .ZN(n8230) );
  NAND2_X1 U10621 ( .A1(n8230), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8200) );
  MUX2_X1 U10622 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8200), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8203) );
  INV_X1 U10623 ( .A(P2_B_REG_SCAN_IN), .ZN(n8204) );
  XNOR2_X1 U10624 ( .A(n8226), .B(n8204), .ZN(n8210) );
  NAND2_X1 U10625 ( .A1(n8206), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8205) );
  MUX2_X1 U10626 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8205), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8209) );
  INV_X1 U10627 ( .A(n8206), .ZN(n8208) );
  NAND2_X1 U10628 ( .A1(n8208), .A2(n8207), .ZN(n8211) );
  NAND2_X1 U10629 ( .A1(n8209), .A2(n8211), .ZN(n13802) );
  NAND2_X1 U10630 ( .A1(n8210), .A2(n13802), .ZN(n8215) );
  NAND2_X1 U10631 ( .A1(n8211), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8212) );
  MUX2_X1 U10632 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8212), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8213) );
  INV_X1 U10633 ( .A(n13800), .ZN(n8214) );
  OAI21_X1 U10634 ( .B1(n8217), .B2(n8216), .A(n14965), .ZN(n10623) );
  INV_X1 U10635 ( .A(n10623), .ZN(n8220) );
  INV_X1 U10636 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14971) );
  NAND2_X1 U10637 ( .A1(n14965), .A2(n14971), .ZN(n8219) );
  NAND2_X1 U10638 ( .A1(n13800), .A2(n13802), .ZN(n8218) );
  NAND2_X1 U10639 ( .A1(n8219), .A2(n8218), .ZN(n14972) );
  INV_X1 U10640 ( .A(n9211), .ZN(n9267) );
  AND2_X1 U10641 ( .A1(n10616), .A2(n8221), .ZN(n10067) );
  OR2_X1 U10642 ( .A1(n14990), .A2(n10067), .ZN(n8222) );
  NOR2_X1 U10643 ( .A1(n8242), .A2(n8222), .ZN(n8232) );
  INV_X1 U10644 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14969) );
  NAND2_X1 U10645 ( .A1(n14965), .A2(n14969), .ZN(n8224) );
  INV_X1 U10646 ( .A(n8226), .ZN(n13804) );
  NAND2_X1 U10647 ( .A1(n13804), .A2(n13800), .ZN(n8223) );
  NAND2_X1 U10648 ( .A1(n8224), .A2(n8223), .ZN(n9931) );
  NOR2_X1 U10649 ( .A1(n13800), .A2(n13802), .ZN(n8225) );
  NAND2_X1 U10650 ( .A1(n8226), .A2(n8225), .ZN(n9915) );
  INV_X1 U10651 ( .A(n8227), .ZN(n8228) );
  NAND2_X1 U10652 ( .A1(n8228), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8229) );
  MUX2_X1 U10653 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8229), .S(
        P2_IR_REG_23__SCAN_IN), .Z(n8231) );
  NAND2_X1 U10654 ( .A1(n8231), .A2(n8230), .ZN(n10068) );
  INV_X1 U10655 ( .A(n14973), .ZN(n14970) );
  OR2_X1 U10656 ( .A1(n9931), .A2(n14970), .ZN(n14968) );
  INV_X1 U10657 ( .A(n14968), .ZN(n10631) );
  OAI21_X1 U10658 ( .B1(n11674), .B2(n13444), .A(n14860), .ZN(n8258) );
  INV_X1 U10659 ( .A(n8242), .ZN(n9933) );
  AND2_X1 U10660 ( .A1(n8236), .A2(n9924), .ZN(n9936) );
  NAND3_X1 U10661 ( .A1(n9933), .A2(n10631), .A3(n9936), .ZN(n8238) );
  INV_X1 U10662 ( .A(n10637), .ZN(n9257) );
  NAND2_X1 U10663 ( .A1(n8236), .A2(n9257), .ZN(n10622) );
  INV_X1 U10664 ( .A(n10622), .ZN(n8237) );
  OAI21_X1 U10665 ( .B1(n8242), .B2(n9931), .A(n10622), .ZN(n8241) );
  INV_X1 U10666 ( .A(n10629), .ZN(n9930) );
  AND2_X1 U10667 ( .A1(n8239), .A2(n9930), .ZN(n8240) );
  NAND2_X1 U10668 ( .A1(n8241), .A2(n8240), .ZN(n10418) );
  NOR2_X1 U10669 ( .A1(n14870), .A2(n13460), .ZN(n8256) );
  NOR2_X1 U10670 ( .A1(n8242), .A2(n9267), .ZN(n8243) );
  NAND2_X1 U10671 ( .A1(n8243), .A2(n10631), .ZN(n14859) );
  NAND2_X1 U10672 ( .A1(n9210), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8252) );
  INV_X1 U10673 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8245) );
  OR2_X1 U10674 ( .A1(n8246), .A2(n8245), .ZN(n8251) );
  OR2_X1 U10675 ( .A1(n8247), .A2(n13447), .ZN(n8250) );
  INV_X1 U10676 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n13448) );
  OR2_X1 U10677 ( .A1(n8248), .A2(n13448), .ZN(n8249) );
  AND4_X1 U10678 ( .A1(n8252), .A2(n8251), .A3(n8250), .A4(n8249), .ZN(n9176)
         );
  INV_X1 U10679 ( .A(n8244), .ZN(n8253) );
  NAND2_X1 U10680 ( .A1(n10067), .A2(n8253), .ZN(n13594) );
  AOI22_X1 U10681 ( .A1(n15413), .A2(n13295), .B1(n13297), .B2(n13576), .ZN(
        n13456) );
  OAI22_X1 U10682 ( .A1(n14859), .A2(n13456), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8254), .ZN(n8255) );
  AOI211_X1 U10683 ( .C1(n13668), .C2(n14867), .A(n8256), .B(n8255), .ZN(n8257) );
  INV_X1 U10684 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n8836) );
  NAND4_X1 U10685 ( .A1(n8267), .A2(n7471), .A3(n8833), .A4(n8805), .ZN(n8268)
         );
  INV_X1 U10686 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10226) );
  NAND2_X1 U10687 ( .A1(n8299), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8278) );
  AND2_X4 U10688 ( .A1(n13176), .A2(n12294), .ZN(n8313) );
  NAND2_X1 U10689 ( .A1(n8313), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8277) );
  NAND2_X1 U10690 ( .A1(n8282), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8283) );
  XNOR2_X1 U10691 ( .A(n8305), .B(n8303), .ZN(n10012) );
  XNOR2_X1 U10692 ( .A(P3_IR_REG_1__SCAN_IN), .B(n8286), .ZN(n10416) );
  INV_X1 U10693 ( .A(n8887), .ZN(n15104) );
  NAND2_X1 U10694 ( .A1(n8534), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8292) );
  NAND2_X1 U10695 ( .A1(n8299), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8291) );
  NAND2_X1 U10696 ( .A1(n8313), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8289) );
  NAND4_X2 U10697 ( .A1(n8292), .A2(n8291), .A3(n8290), .A4(n8289), .ZN(n15108) );
  NAND2_X1 U10698 ( .A1(n8371), .A2(SI_0_), .ZN(n8297) );
  INV_X1 U10699 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9350) );
  NAND2_X1 U10700 ( .A1(n9350), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8293) );
  NAND2_X1 U10701 ( .A1(n8303), .A2(n8293), .ZN(n9997) );
  INV_X1 U10702 ( .A(n9997), .ZN(n8294) );
  NAND2_X1 U10703 ( .A1(n8601), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n8295) );
  AND3_X2 U10704 ( .A1(n8297), .A2(n8296), .A3(n8295), .ZN(n10698) );
  INV_X1 U10705 ( .A(n10698), .ZN(n10583) );
  NAND2_X1 U10706 ( .A1(n10522), .A2(n15104), .ZN(n8884) );
  NAND2_X1 U10707 ( .A1(n8313), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8301) );
  NAND2_X1 U10708 ( .A1(n8534), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8300) );
  INV_X1 U10709 ( .A(n8303), .ZN(n8304) );
  NAND2_X1 U10710 ( .A1(n9946), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8306) );
  NAND2_X1 U10711 ( .A1(n9956), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U10712 ( .A1(n9944), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8307) );
  AND2_X1 U10713 ( .A1(n8318), .A2(n8307), .ZN(n8316) );
  XNOR2_X1 U10714 ( .A(n8317), .B(n8316), .ZN(n9978) );
  NOR2_X1 U10715 ( .A1(n8552), .A2(SI_2_), .ZN(n8310) );
  INV_X1 U10716 ( .A(n8892), .ZN(n15088) );
  NAND2_X1 U10717 ( .A1(n10894), .A2(n15088), .ZN(n8312) );
  NAND2_X1 U10718 ( .A1(n8747), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8315) );
  NAND2_X1 U10719 ( .A1(n8313), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8314) );
  NAND2_X1 U10720 ( .A1(n9960), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8334) );
  INV_X1 U10721 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9950) );
  NAND2_X1 U10722 ( .A1(n9950), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8319) );
  NAND2_X1 U10723 ( .A1(n8334), .A2(n8319), .ZN(n8331) );
  XNOR2_X1 U10724 ( .A(n8333), .B(n8331), .ZN(n10004) );
  NAND2_X1 U10725 ( .A1(n12487), .A2(n10004), .ZN(n8323) );
  OR2_X1 U10726 ( .A1(n8320), .A2(n8273), .ZN(n8321) );
  XNOR2_X1 U10727 ( .A(n8321), .B(n8337), .ZN(n10501) );
  NAND2_X1 U10728 ( .A1(n8601), .A2(n10501), .ZN(n8322) );
  OAI211_X1 U10729 ( .C1(SI_3_), .C2(n8552), .A(n8323), .B(n8322), .ZN(n10901)
         );
  NAND2_X1 U10730 ( .A1(n12712), .A2(n10901), .ZN(n12545) );
  NAND2_X1 U10731 ( .A1(n12712), .A2(n8324), .ZN(n8325) );
  NAND2_X1 U10732 ( .A1(n8747), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8330) );
  NAND2_X1 U10733 ( .A1(n8299), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8329) );
  AND2_X1 U10734 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8326) );
  NOR2_X1 U10735 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8344) );
  OR2_X1 U10736 ( .A1(n8326), .A2(n8344), .ZN(n10943) );
  NAND2_X1 U10737 ( .A1(n8765), .A2(n10943), .ZN(n8328) );
  NAND2_X1 U10738 ( .A1(n8313), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8327) );
  INV_X1 U10739 ( .A(n8331), .ZN(n8332) );
  NAND2_X1 U10740 ( .A1(n8333), .A2(n8332), .ZN(n8335) );
  NAND2_X1 U10741 ( .A1(n9963), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8353) );
  NAND2_X1 U10742 ( .A1(n9954), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8336) );
  XNOR2_X1 U10743 ( .A(n8352), .B(n8351), .ZN(n9976) );
  NAND2_X1 U10744 ( .A1(n8320), .A2(n8337), .ZN(n8339) );
  NAND2_X1 U10745 ( .A1(n8339), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8338) );
  MUX2_X1 U10746 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8338), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n8340) );
  OAI22_X1 U10747 ( .A1(n8412), .A2(n9976), .B1(n10390), .B2(n10243), .ZN(
        n8342) );
  NOR2_X1 U10748 ( .A1(n8552), .A2(SI_4_), .ZN(n8341) );
  NOR2_X1 U10749 ( .A1(n8342), .A2(n8341), .ZN(n8900) );
  INV_X1 U10750 ( .A(n8900), .ZN(n10942) );
  NAND2_X1 U10751 ( .A1(n10942), .A2(n15074), .ZN(n12553) );
  NAND2_X1 U10752 ( .A1(n15074), .A2(n8900), .ZN(n8343) );
  NAND2_X1 U10753 ( .A1(n8747), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8350) );
  NAND2_X1 U10754 ( .A1(n12489), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8349) );
  NAND2_X1 U10755 ( .A1(n8344), .A2(n8345), .ZN(n8361) );
  OR2_X1 U10756 ( .A1(n8345), .A2(n8344), .ZN(n8346) );
  NAND2_X1 U10757 ( .A1(n8361), .A2(n8346), .ZN(n15082) );
  NAND2_X1 U10758 ( .A1(n8765), .A2(n15082), .ZN(n8348) );
  NAND2_X1 U10759 ( .A1(n8313), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8347) );
  NAND2_X1 U10760 ( .A1(n9958), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8369) );
  NAND2_X1 U10761 ( .A1(n9952), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8354) );
  XNOR2_X1 U10762 ( .A(n8368), .B(n8367), .ZN(n9983) );
  NAND2_X1 U10763 ( .A1(n8372), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8355) );
  OAI22_X1 U10764 ( .A1(n8412), .A2(n9983), .B1(n10400), .B2(n10243), .ZN(
        n8357) );
  NOR2_X1 U10765 ( .A1(n8552), .A2(SI_5_), .ZN(n8356) );
  NOR2_X1 U10766 ( .A1(n8357), .A2(n8356), .ZN(n15081) );
  NAND2_X1 U10767 ( .A1(n11092), .A2(n15081), .ZN(n12555) );
  INV_X1 U10768 ( .A(n15081), .ZN(n10908) );
  NAND2_X1 U10769 ( .A1(n10908), .A2(n12711), .ZN(n12551) );
  NAND2_X1 U10770 ( .A1(n11092), .A2(n10908), .ZN(n8360) );
  NAND2_X1 U10771 ( .A1(n8747), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8366) );
  NAND2_X1 U10772 ( .A1(n12489), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8365) );
  NAND2_X1 U10773 ( .A1(n8361), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8362) );
  NAND2_X1 U10774 ( .A1(n8377), .A2(n8362), .ZN(n11316) );
  NAND2_X1 U10775 ( .A1(n8765), .A2(n11316), .ZN(n8364) );
  NAND2_X1 U10776 ( .A1(n8313), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8363) );
  INV_X1 U10777 ( .A(n15073), .ZN(n11208) );
  XNOR2_X1 U10778 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8370) );
  XNOR2_X1 U10779 ( .A(n8387), .B(n8370), .ZN(n10013) );
  NAND2_X1 U10780 ( .A1(n12487), .A2(n10013), .ZN(n8376) );
  NAND2_X1 U10781 ( .A1(n12479), .A2(SI_6_), .ZN(n8375) );
  OR2_X1 U10782 ( .A1(n8384), .A2(n8273), .ZN(n8373) );
  INV_X1 U10783 ( .A(n11028), .ZN(n10845) );
  NAND2_X1 U10784 ( .A1(n8601), .A2(n10845), .ZN(n8374) );
  INV_X1 U10785 ( .A(n15147), .ZN(n11317) );
  NAND2_X1 U10786 ( .A1(n15073), .A2(n15147), .ZN(n12556) );
  NAND2_X1 U10787 ( .A1(n12564), .A2(n12556), .ZN(n11309) );
  NAND2_X1 U10788 ( .A1(n8747), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U10789 ( .A1(n12489), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8381) );
  AND2_X1 U10790 ( .A1(n8377), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8378) );
  OR2_X1 U10791 ( .A1(n8378), .A2(n8426), .ZN(n11237) );
  NAND2_X1 U10792 ( .A1(n8765), .A2(n11237), .ZN(n8380) );
  NAND2_X1 U10793 ( .A1(n8313), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8379) );
  NAND4_X1 U10794 ( .A1(n8382), .A2(n8381), .A3(n8380), .A4(n8379), .ZN(n12710) );
  OR2_X1 U10795 ( .A1(n8408), .A2(n8273), .ZN(n8385) );
  XNOR2_X1 U10796 ( .A(n8385), .B(P3_IR_REG_7__SCAN_IN), .ZN(n11292) );
  OAI22_X1 U10797 ( .A1(n8552), .A2(SI_7_), .B1(n11292), .B2(n10243), .ZN(
        n8395) );
  NAND2_X1 U10798 ( .A1(n9965), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8386) );
  NAND2_X1 U10799 ( .A1(n9968), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8388) );
  NAND2_X1 U10800 ( .A1(n9972), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8401) );
  NAND2_X1 U10801 ( .A1(n9970), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8390) );
  NAND2_X1 U10802 ( .A1(n8401), .A2(n8390), .ZN(n8391) );
  NAND2_X1 U10803 ( .A1(n8392), .A2(n8391), .ZN(n8393) );
  AND2_X1 U10804 ( .A1(n8402), .A2(n8393), .ZN(n9985) );
  NOR2_X1 U10805 ( .A1(n8412), .A2(n9985), .ZN(n8394) );
  NOR2_X1 U10806 ( .A1(n8395), .A2(n8394), .ZN(n11236) );
  XNOR2_X1 U10807 ( .A(n12710), .B(n11236), .ZN(n12562) );
  INV_X1 U10808 ( .A(n12562), .ZN(n11231) );
  NAND2_X1 U10809 ( .A1(n12710), .A2(n11236), .ZN(n8396) );
  NAND2_X1 U10810 ( .A1(n8747), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8400) );
  NAND2_X1 U10811 ( .A1(n12489), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8399) );
  INV_X1 U10812 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n8425) );
  XNOR2_X1 U10813 ( .A(n8426), .B(n8425), .ZN(n11576) );
  NAND2_X1 U10814 ( .A1(n8765), .A2(n11576), .ZN(n8398) );
  NAND2_X1 U10815 ( .A1(n8313), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8397) );
  NAND4_X1 U10816 ( .A1(n8400), .A2(n8399), .A3(n8398), .A4(n8397), .ZN(n12709) );
  INV_X1 U10817 ( .A(n12709), .ZN(n11560) );
  NAND2_X1 U10818 ( .A1(n10003), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8415) );
  NAND2_X1 U10819 ( .A1(n10001), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8403) );
  OR2_X1 U10820 ( .A1(n8405), .A2(n8404), .ZN(n8406) );
  NAND2_X1 U10821 ( .A1(n8416), .A2(n8406), .ZN(n10006) );
  INV_X1 U10822 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8407) );
  INV_X1 U10823 ( .A(n11286), .ZN(n15035) );
  NAND2_X1 U10824 ( .A1(n8601), .A2(n15035), .ZN(n8411) );
  NAND2_X1 U10825 ( .A1(n12479), .A2(SI_8_), .ZN(n8410) );
  OAI211_X1 U10826 ( .C1(n10006), .C2(n8412), .A(n8411), .B(n8410), .ZN(n11575) );
  NAND2_X1 U10827 ( .A1(n11560), .A2(n11575), .ZN(n12573) );
  INV_X1 U10828 ( .A(n11575), .ZN(n11360) );
  NAND2_X1 U10829 ( .A1(n12709), .A2(n11360), .ZN(n12572) );
  NAND2_X1 U10830 ( .A1(n11560), .A2(n11360), .ZN(n8414) );
  NAND2_X1 U10831 ( .A1(n10057), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8442) );
  NAND2_X1 U10832 ( .A1(n10059), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8417) );
  XNOR2_X1 U10833 ( .A(n6885), .B(n8440), .ZN(n10017) );
  NAND2_X1 U10834 ( .A1(n10017), .A2(n12487), .ZN(n8422) );
  NAND2_X1 U10835 ( .A1(n8418), .A2(n7369), .ZN(n8447) );
  NAND2_X1 U10836 ( .A1(n8447), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8419) );
  OAI22_X1 U10837 ( .A1(n8552), .A2(SI_9_), .B1(n15053), .B2(n10243), .ZN(
        n8420) );
  INV_X1 U10838 ( .A(n8420), .ZN(n8421) );
  NAND2_X1 U10839 ( .A1(n8422), .A2(n8421), .ZN(n11624) );
  INV_X1 U10840 ( .A(n11624), .ZN(n12577) );
  NAND2_X1 U10841 ( .A1(n12489), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8431) );
  NAND2_X1 U10842 ( .A1(n8313), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8430) );
  NOR2_X1 U10843 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_REG3_REG_9__SCAN_IN), 
        .ZN(n8423) );
  INV_X1 U10844 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8424) );
  AOI21_X1 U10845 ( .B1(n8426), .B2(n8425), .A(n8424), .ZN(n8427) );
  OR2_X1 U10846 ( .A1(n8434), .A2(n8427), .ZN(n11625) );
  NAND2_X1 U10847 ( .A1(n8765), .A2(n11625), .ZN(n8429) );
  NAND2_X1 U10848 ( .A1(n8747), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8428) );
  NAND4_X1 U10849 ( .A1(n8431), .A2(n8430), .A3(n8429), .A4(n8428), .ZN(n12708) );
  NAND2_X1 U10850 ( .A1(n12577), .A2(n12708), .ZN(n12578) );
  INV_X1 U10851 ( .A(n12708), .ZN(n11655) );
  NAND2_X1 U10852 ( .A1(n11655), .A2(n11624), .ZN(n8432) );
  NAND2_X1 U10853 ( .A1(n12489), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8439) );
  OR2_X1 U10854 ( .A1(n8434), .A2(n8433), .ZN(n8435) );
  NAND2_X1 U10855 ( .A1(n8477), .A2(n8435), .ZN(n11650) );
  NAND2_X1 U10856 ( .A1(n8765), .A2(n11650), .ZN(n8438) );
  NAND2_X1 U10857 ( .A1(n8313), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8437) );
  INV_X1 U10858 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11689) );
  OR2_X1 U10859 ( .A1(n12493), .A2(n11689), .ZN(n8436) );
  NAND2_X1 U10860 ( .A1(n10224), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8459) );
  NAND2_X1 U10861 ( .A1(n10222), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8443) );
  OR2_X1 U10862 ( .A1(n8445), .A2(n8444), .ZN(n8446) );
  NAND2_X1 U10863 ( .A1(n8460), .A2(n8446), .ZN(n10009) );
  NAND2_X1 U10864 ( .A1(n10009), .A2(n12487), .ZN(n8451) );
  INV_X1 U10865 ( .A(SI_10_), .ZN(n10010) );
  NAND2_X1 U10866 ( .A1(n8462), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8449) );
  INV_X1 U10867 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8448) );
  AOI22_X1 U10868 ( .A1(n12479), .A2(n10010), .B1(n11842), .B2(n8601), .ZN(
        n8450) );
  NAND2_X1 U10869 ( .A1(n8451), .A2(n8450), .ZN(n15168) );
  XNOR2_X1 U10870 ( .A(n12707), .B(n15168), .ZN(n12508) );
  NAND2_X1 U10871 ( .A1(n11685), .A2(n12508), .ZN(n11684) );
  OR2_X1 U10872 ( .A1(n14674), .A2(n15168), .ZN(n8452) );
  NAND2_X1 U10873 ( .A1(n11684), .A2(n8452), .ZN(n14672) );
  NAND2_X1 U10874 ( .A1(n12489), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8458) );
  XNOR2_X1 U10875 ( .A(n8477), .B(P3_REG3_REG_11__SCAN_IN), .ZN(n14678) );
  NAND2_X1 U10876 ( .A1(n8765), .A2(n14678), .ZN(n8457) );
  INV_X1 U10877 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n8453) );
  OR2_X1 U10878 ( .A1(n8750), .A2(n8453), .ZN(n8456) );
  INV_X1 U10879 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n8454) );
  OR2_X1 U10880 ( .A1(n12493), .A2(n8454), .ZN(n8455) );
  XNOR2_X1 U10881 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8461) );
  XNOR2_X1 U10882 ( .A(n8470), .B(n8461), .ZN(n10007) );
  NAND2_X1 U10883 ( .A1(n10007), .A2(n12487), .ZN(n8466) );
  OAI21_X1 U10884 ( .B1(n8462), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8464) );
  INV_X1 U10885 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8463) );
  XNOR2_X1 U10886 ( .A(n8464), .B(n8463), .ZN(n11949) );
  AOI22_X1 U10887 ( .A1(n11949), .A2(n8601), .B1(n12479), .B2(n10008), .ZN(
        n8465) );
  NAND2_X1 U10888 ( .A1(n8466), .A2(n8465), .ZN(n14677) );
  INV_X1 U10889 ( .A(n14677), .ZN(n8467) );
  NAND2_X1 U10890 ( .A1(n14672), .A2(n14657), .ZN(n8468) );
  NAND2_X1 U10891 ( .A1(n10380), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8469) );
  NAND2_X1 U10892 ( .A1(n8470), .A2(n8469), .ZN(n8472) );
  NAND2_X1 U10893 ( .A1(n10377), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8471) );
  XNOR2_X1 U10894 ( .A(n10504), .B(P2_DATAO_REG_12__SCAN_IN), .ZN(n8493) );
  XNOR2_X1 U10895 ( .A(n8495), .B(n8493), .ZN(n9980) );
  XNOR2_X1 U10896 ( .A(n8474), .B(P3_IR_REG_12__SCAN_IN), .ZN(n11964) );
  OAI22_X1 U10897 ( .A1(n8552), .A2(n9982), .B1(n10243), .B2(n12726), .ZN(
        n8475) );
  AOI21_X1 U10898 ( .B1(n9980), .B2(n12487), .A(n8475), .ZN(n14663) );
  NAND2_X1 U10899 ( .A1(n12489), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8482) );
  NAND2_X1 U10900 ( .A1(n8747), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8481) );
  OAI21_X1 U10901 ( .B1(n8477), .B2(P3_REG3_REG_11__SCAN_IN), .A(
        P3_REG3_REG_12__SCAN_IN), .ZN(n8478) );
  NAND2_X1 U10902 ( .A1(n8478), .A2(n8486), .ZN(n14660) );
  NAND2_X1 U10903 ( .A1(n8765), .A2(n14660), .ZN(n8480) );
  NAND2_X1 U10904 ( .A1(n8313), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8479) );
  NAND4_X1 U10905 ( .A1(n8482), .A2(n8481), .A3(n8480), .A4(n8479), .ZN(n12706) );
  OR2_X1 U10906 ( .A1(n14663), .A2(n12706), .ZN(n12593) );
  NAND2_X1 U10907 ( .A1(n14663), .A2(n12706), .ZN(n12594) );
  NAND2_X1 U10908 ( .A1(n12593), .A2(n12594), .ZN(n8783) );
  INV_X1 U10909 ( .A(n12706), .ZN(n14675) );
  OR2_X1 U10910 ( .A1(n14663), .A2(n14675), .ZN(n8483) );
  NAND2_X1 U10911 ( .A1(n12489), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8492) );
  INV_X1 U10912 ( .A(n8486), .ZN(n8485) );
  NAND2_X1 U10913 ( .A1(n8486), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8487) );
  AND2_X1 U10914 ( .A1(n8514), .A2(n8487), .ZN(n14648) );
  INV_X1 U10915 ( .A(n14648), .ZN(n8488) );
  NAND2_X1 U10916 ( .A1(n8765), .A2(n8488), .ZN(n8491) );
  NAND2_X1 U10917 ( .A1(n8313), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8490) );
  INV_X1 U10918 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12716) );
  OR2_X1 U10919 ( .A1(n12493), .A2(n12716), .ZN(n8489) );
  INV_X1 U10920 ( .A(n8493), .ZN(n8494) );
  NAND2_X1 U10921 ( .A1(n8495), .A2(n8494), .ZN(n8498) );
  NAND2_X1 U10922 ( .A1(n8496), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8497) );
  XNOR2_X1 U10923 ( .A(n8505), .B(n10615), .ZN(n10113) );
  NAND2_X1 U10924 ( .A1(n10113), .A2(n12487), .ZN(n8504) );
  NAND2_X1 U10925 ( .A1(n8500), .A2(n8499), .ZN(n8508) );
  NAND2_X1 U10926 ( .A1(n8508), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8501) );
  XNOR2_X1 U10927 ( .A(n8501), .B(P3_IR_REG_13__SCAN_IN), .ZN(n12745) );
  INV_X1 U10928 ( .A(n12745), .ZN(n12717) );
  OAI22_X1 U10929 ( .A1(n8552), .A2(n10115), .B1(n10243), .B2(n12717), .ZN(
        n8502) );
  INV_X1 U10930 ( .A(n8502), .ZN(n8503) );
  NAND2_X1 U10931 ( .A1(n8504), .A2(n8503), .ZN(n12036) );
  INV_X1 U10932 ( .A(n12036), .ZN(n14651) );
  NAND2_X1 U10933 ( .A1(n8506), .A2(n10613), .ZN(n8507) );
  XNOR2_X1 U10934 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8522) );
  XNOR2_X1 U10935 ( .A(n8523), .B(n8522), .ZN(n10128) );
  NAND2_X1 U10936 ( .A1(n10128), .A2(n12487), .ZN(n8512) );
  OR2_X1 U10937 ( .A1(n8527), .A2(n8273), .ZN(n8509) );
  XNOR2_X1 U10938 ( .A(n8509), .B(n8526), .ZN(n12766) );
  INV_X1 U10939 ( .A(n12766), .ZN(n12753) );
  OAI22_X1 U10940 ( .A1(n8552), .A2(SI_14_), .B1(n12753), .B2(n10243), .ZN(
        n8510) );
  INV_X1 U10941 ( .A(n8510), .ZN(n8511) );
  NAND2_X1 U10942 ( .A1(n8747), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8519) );
  NAND2_X1 U10943 ( .A1(n12489), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8518) );
  INV_X1 U10944 ( .A(n8514), .ZN(n8513) );
  NAND2_X1 U10945 ( .A1(n8514), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8515) );
  NAND2_X1 U10946 ( .A1(n8532), .A2(n8515), .ZN(n12131) );
  NAND2_X1 U10947 ( .A1(n8765), .A2(n12131), .ZN(n8517) );
  NAND2_X1 U10948 ( .A1(n8313), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8516) );
  NAND4_X1 U10949 ( .A1(n8519), .A2(n8518), .A3(n8517), .A4(n8516), .ZN(n12705) );
  NAND2_X1 U10950 ( .A1(n12243), .A2(n12705), .ZN(n12604) );
  INV_X1 U10951 ( .A(n12705), .ZN(n14647) );
  OR2_X1 U10952 ( .A1(n12243), .A2(n14647), .ZN(n8521) );
  NAND2_X1 U10953 ( .A1(n8524), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8525) );
  XNOR2_X1 U10954 ( .A(n10950), .B(P1_DATAO_REG_15__SCAN_IN), .ZN(n8540) );
  XNOR2_X1 U10955 ( .A(n8542), .B(n8540), .ZN(n10325) );
  NAND2_X1 U10956 ( .A1(n10325), .A2(n12487), .ZN(n8531) );
  OR2_X1 U10957 ( .A1(n8546), .A2(n8273), .ZN(n8528) );
  XNOR2_X1 U10958 ( .A(n8528), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12788) );
  INV_X1 U10959 ( .A(n12788), .ZN(n12782) );
  OAI22_X1 U10960 ( .A1(n8552), .A2(n15360), .B1(n10243), .B2(n12782), .ZN(
        n8529) );
  INV_X1 U10961 ( .A(n8529), .ZN(n8530) );
  NAND2_X1 U10962 ( .A1(n8747), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U10963 ( .A1(n12489), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8537) );
  NAND2_X1 U10964 ( .A1(n8532), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U10965 ( .A1(n8554), .A2(n8533), .ZN(n12187) );
  NAND2_X1 U10966 ( .A1(n8765), .A2(n12187), .ZN(n8536) );
  NAND2_X1 U10967 ( .A1(n8313), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8535) );
  NAND4_X1 U10968 ( .A1(n8538), .A2(n8537), .A3(n8536), .A4(n8535), .ZN(n12704) );
  OR2_X1 U10969 ( .A1(n12152), .A2(n12412), .ZN(n12608) );
  NAND2_X1 U10970 ( .A1(n12152), .A2(n12412), .ZN(n12613) );
  NAND2_X1 U10971 ( .A1(n12608), .A2(n12613), .ZN(n12182) );
  NAND2_X1 U10972 ( .A1(n12152), .A2(n12704), .ZN(n8539) );
  INV_X1 U10973 ( .A(n8540), .ZN(n8541) );
  NAND2_X1 U10974 ( .A1(n10950), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8543) );
  XNOR2_X1 U10975 ( .A(n11173), .B(P2_DATAO_REG_16__SCAN_IN), .ZN(n8561) );
  XNOR2_X1 U10976 ( .A(n8563), .B(n8561), .ZN(n10381) );
  NOR2_X1 U10977 ( .A1(n8550), .A2(n8273), .ZN(n8547) );
  MUX2_X1 U10978 ( .A(n8273), .B(n8547), .S(P3_IR_REG_16__SCAN_IN), .Z(n8548)
         );
  INV_X1 U10979 ( .A(n8548), .ZN(n8551) );
  NAND2_X1 U10980 ( .A1(n8551), .A2(n8581), .ZN(n12802) );
  OAI22_X1 U10981 ( .A1(n8552), .A2(n10383), .B1(n12802), .B2(n10243), .ZN(
        n8553) );
  NAND2_X1 U10982 ( .A1(n8747), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8559) );
  NAND2_X1 U10983 ( .A1(n12489), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8558) );
  INV_X1 U10984 ( .A(n8569), .ZN(n8570) );
  NAND2_X1 U10985 ( .A1(n8554), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8555) );
  NAND2_X1 U10986 ( .A1(n8570), .A2(n8555), .ZN(n12415) );
  NAND2_X1 U10987 ( .A1(n8765), .A2(n12415), .ZN(n8557) );
  NAND2_X1 U10988 ( .A1(n8313), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8556) );
  NAND4_X1 U10989 ( .A1(n8559), .A2(n8558), .A3(n8557), .A4(n8556), .ZN(n13035) );
  NAND2_X1 U10990 ( .A1(n13158), .A2(n13035), .ZN(n12615) );
  NAND2_X1 U10991 ( .A1(n12614), .A2(n12615), .ZN(n12253) );
  INV_X1 U10992 ( .A(n13035), .ZN(n12424) );
  OR2_X1 U10993 ( .A1(n13158), .A2(n12424), .ZN(n8560) );
  INV_X1 U10994 ( .A(n8561), .ZN(n8562) );
  NAND2_X1 U10995 ( .A1(n11171), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8564) );
  XNOR2_X1 U10996 ( .A(n11346), .B(P1_DATAO_REG_17__SCAN_IN), .ZN(n8577) );
  XNOR2_X1 U10997 ( .A(n8579), .B(n8577), .ZN(n10516) );
  NAND2_X1 U10998 ( .A1(n10516), .A2(n12487), .ZN(n8567) );
  NAND2_X1 U10999 ( .A1(n8581), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8565) );
  XNOR2_X1 U11000 ( .A(n8565), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12831) );
  AOI22_X1 U11001 ( .A1(n12479), .A2(SI_17_), .B1(n8601), .B2(n12831), .ZN(
        n8566) );
  INV_X1 U11002 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8568) );
  INV_X1 U11003 ( .A(n8586), .ZN(n8587) );
  NAND2_X1 U11004 ( .A1(n8570), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8571) );
  NAND2_X1 U11005 ( .A1(n8587), .A2(n8571), .ZN(n13042) );
  NAND2_X1 U11006 ( .A1(n13042), .A2(n8765), .ZN(n8575) );
  NAND2_X1 U11007 ( .A1(n8747), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8574) );
  NAND2_X1 U11008 ( .A1(n12489), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8573) );
  INV_X1 U11009 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n15334) );
  OR2_X1 U11010 ( .A1(n8750), .A2(n15334), .ZN(n8572) );
  OR2_X1 U11011 ( .A1(n13041), .A2(n12418), .ZN(n12619) );
  NAND2_X1 U11012 ( .A1(n13041), .A2(n12418), .ZN(n12618) );
  NAND2_X1 U11013 ( .A1(n12619), .A2(n12618), .ZN(n13033) );
  NAND2_X1 U11014 ( .A1(n13041), .A2(n13021), .ZN(n8576) );
  INV_X1 U11015 ( .A(n8577), .ZN(n8578) );
  NAND2_X1 U11016 ( .A1(n11346), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8580) );
  XNOR2_X1 U11017 ( .A(n8595), .B(P1_DATAO_REG_18__SCAN_IN), .ZN(n8592) );
  XNOR2_X1 U11018 ( .A(n8594), .B(n8592), .ZN(n10643) );
  NAND2_X1 U11019 ( .A1(n10643), .A2(n12487), .ZN(n8584) );
  NAND2_X1 U11020 ( .A1(n8598), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8582) );
  XNOR2_X1 U11021 ( .A(n8582), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12839) );
  AOI22_X1 U11022 ( .A1(SI_18_), .A2(n12479), .B1(n12839), .B2(n8601), .ZN(
        n8583) );
  INV_X1 U11023 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n8591) );
  INV_X1 U11024 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n8585) );
  NAND2_X1 U11025 ( .A1(n8587), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U11026 ( .A1(n8604), .A2(n8588), .ZN(n13024) );
  NAND2_X1 U11027 ( .A1(n13024), .A2(n8765), .ZN(n8590) );
  AOI22_X1 U11028 ( .A1(n8747), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n12489), 
        .B2(P3_REG1_REG_18__SCAN_IN), .ZN(n8589) );
  OAI211_X1 U11029 ( .C1(n8750), .C2(n8591), .A(n8590), .B(n8589), .ZN(n13036)
         );
  INV_X1 U11030 ( .A(n13036), .ZN(n8931) );
  NAND2_X1 U11031 ( .A1(n13098), .A2(n8931), .ZN(n12625) );
  INV_X1 U11032 ( .A(n8592), .ZN(n8593) );
  NAND2_X1 U11033 ( .A1(n8595), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8596) );
  XNOR2_X1 U11034 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .ZN(n8608) );
  XNOR2_X1 U11035 ( .A(n8609), .B(n8608), .ZN(n12263) );
  NAND2_X1 U11036 ( .A1(n12263), .A2(n12487), .ZN(n8603) );
  XNOR2_X1 U11037 ( .A(n8600), .B(n8599), .ZN(n8880) );
  AOI22_X1 U11038 ( .A1(n12859), .A2(n8601), .B1(n12479), .B2(n12262), .ZN(
        n8602) );
  INV_X1 U11039 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13149) );
  NAND2_X1 U11040 ( .A1(n8604), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8605) );
  NAND2_X1 U11041 ( .A1(n8613), .A2(n8605), .ZN(n13013) );
  NAND2_X1 U11042 ( .A1(n13013), .A2(n8765), .ZN(n8607) );
  AOI22_X1 U11043 ( .A1(n8747), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n12489), 
        .B2(P3_REG1_REG_19__SCAN_IN), .ZN(n8606) );
  OAI211_X1 U11044 ( .C1(n8750), .C2(n13149), .A(n8607), .B(n8606), .ZN(n13022) );
  INV_X1 U11045 ( .A(n13022), .ZN(n12457) );
  NAND2_X1 U11046 ( .A1(n11765), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8610) );
  XNOR2_X1 U11047 ( .A(n8620), .B(n11902), .ZN(n10889) );
  NAND2_X1 U11048 ( .A1(n10889), .A2(n12487), .ZN(n8612) );
  NAND2_X1 U11049 ( .A1(n12479), .A2(SI_20_), .ZN(n8611) );
  INV_X1 U11050 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n8617) );
  INV_X1 U11051 ( .A(n8628), .ZN(n8629) );
  NAND2_X1 U11052 ( .A1(n8613), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8614) );
  NAND2_X1 U11053 ( .A1(n8629), .A2(n8614), .ZN(n12995) );
  NAND2_X1 U11054 ( .A1(n12995), .A2(n8765), .ZN(n8616) );
  AOI22_X1 U11055 ( .A1(n8747), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n12489), 
        .B2(P3_REG1_REG_20__SCAN_IN), .ZN(n8615) );
  OAI211_X1 U11056 ( .C1(n8750), .C2(n8617), .A(n8616), .B(n8615), .ZN(n13004)
         );
  INV_X1 U11057 ( .A(n13004), .ZN(n12974) );
  NAND2_X1 U11058 ( .A1(n13090), .A2(n12974), .ZN(n12635) );
  NAND2_X1 U11059 ( .A1(n12634), .A2(n12635), .ZN(n12991) );
  OR2_X1 U11060 ( .A1(n13151), .A2(n13022), .ZN(n12630) );
  NAND2_X1 U11061 ( .A1(n13151), .A2(n13022), .ZN(n12631) );
  NAND2_X1 U11062 ( .A1(n12630), .A2(n12631), .ZN(n13008) );
  OR2_X1 U11063 ( .A1(n13098), .A2(n13036), .ZN(n13003) );
  NAND2_X1 U11064 ( .A1(n13008), .A2(n13003), .ZN(n12984) );
  NAND2_X1 U11065 ( .A1(n12984), .A2(n6497), .ZN(n8618) );
  AND2_X1 U11066 ( .A1(n12991), .A2(n8618), .ZN(n8619) );
  NAND2_X1 U11067 ( .A1(n8621), .A2(n11902), .ZN(n8624) );
  NAND2_X1 U11068 ( .A1(n8622), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8623) );
  INV_X1 U11069 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11982) );
  XNOR2_X1 U11070 ( .A(n11982), .B(P1_DATAO_REG_21__SCAN_IN), .ZN(n8637) );
  XNOR2_X1 U11071 ( .A(n8639), .B(n8637), .ZN(n11066) );
  NAND2_X1 U11072 ( .A1(n11066), .A2(n12487), .ZN(n8626) );
  NAND2_X1 U11073 ( .A1(n12479), .A2(SI_21_), .ZN(n8625) );
  INV_X1 U11074 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U11075 ( .A1(n8629), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8630) );
  NAND2_X1 U11076 ( .A1(n8647), .A2(n8630), .ZN(n12978) );
  NAND2_X1 U11077 ( .A1(n12978), .A2(n8765), .ZN(n8636) );
  INV_X1 U11078 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n8633) );
  NAND2_X1 U11079 ( .A1(n8313), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8632) );
  NAND2_X1 U11080 ( .A1(n12489), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8631) );
  OAI211_X1 U11081 ( .C1(n12493), .C2(n8633), .A(n8632), .B(n8631), .ZN(n8634)
         );
  INV_X1 U11082 ( .A(n8634), .ZN(n8635) );
  AND2_X1 U11083 ( .A1(n12387), .A2(n12988), .ZN(n12515) );
  OR2_X1 U11084 ( .A1(n12387), .A2(n12988), .ZN(n12514) );
  INV_X1 U11085 ( .A(n8637), .ZN(n8638) );
  NAND2_X1 U11086 ( .A1(n11982), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8640) );
  NAND2_X1 U11087 ( .A1(n12371), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U11088 ( .A1(n15226), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8641) );
  NAND2_X1 U11089 ( .A1(n8658), .A2(n8641), .ZN(n8642) );
  NAND2_X1 U11090 ( .A1(n8643), .A2(n8642), .ZN(n8644) );
  NAND2_X1 U11091 ( .A1(n8659), .A2(n8644), .ZN(n11146) );
  NAND2_X1 U11092 ( .A1(n11146), .A2(n12487), .ZN(n8646) );
  NAND2_X1 U11093 ( .A1(n12479), .A2(SI_22_), .ZN(n8645) );
  NAND2_X1 U11094 ( .A1(n8647), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8648) );
  NAND2_X1 U11095 ( .A1(n8666), .A2(n8648), .ZN(n12967) );
  NAND2_X1 U11096 ( .A1(n12967), .A2(n8765), .ZN(n8654) );
  INV_X1 U11097 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U11098 ( .A1(n8313), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8650) );
  NAND2_X1 U11099 ( .A1(n12489), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8649) );
  OAI211_X1 U11100 ( .C1(n12493), .C2(n8651), .A(n8650), .B(n8649), .ZN(n8652)
         );
  INV_X1 U11101 ( .A(n8652), .ZN(n8653) );
  NAND2_X1 U11102 ( .A1(n8654), .A2(n8653), .ZN(n12702) );
  NAND2_X1 U11103 ( .A1(n12966), .A2(n12702), .ZN(n8655) );
  NAND2_X1 U11104 ( .A1(n12960), .A2(n8655), .ZN(n8657) );
  OR2_X1 U11105 ( .A1(n12966), .A2(n12702), .ZN(n8656) );
  NAND2_X1 U11106 ( .A1(n8657), .A2(n8656), .ZN(n12947) );
  NAND2_X1 U11107 ( .A1(n12251), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8676) );
  INV_X1 U11108 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n15248) );
  NAND2_X1 U11109 ( .A1(n15248), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8660) );
  NAND2_X1 U11110 ( .A1(n8677), .A2(n8663), .ZN(n11272) );
  NAND2_X1 U11111 ( .A1(n11272), .A2(n12487), .ZN(n8665) );
  NAND2_X1 U11112 ( .A1(n12479), .A2(SI_23_), .ZN(n8664) );
  NAND2_X1 U11113 ( .A1(n8666), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U11114 ( .A1(n8680), .A2(n8667), .ZN(n12955) );
  NAND2_X1 U11115 ( .A1(n12955), .A2(n8765), .ZN(n8674) );
  INV_X1 U11116 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n8670) );
  NAND2_X1 U11117 ( .A1(n8747), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8669) );
  NAND2_X1 U11118 ( .A1(n8313), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8668) );
  OAI211_X1 U11119 ( .C1(n8671), .C2(n8670), .A(n8669), .B(n8668), .ZN(n8672)
         );
  INV_X1 U11120 ( .A(n8672), .ZN(n8673) );
  NAND2_X1 U11121 ( .A1(n8674), .A2(n8673), .ZN(n12701) );
  NAND2_X1 U11122 ( .A1(n12952), .A2(n12701), .ZN(n8675) );
  XNOR2_X1 U11123 ( .A(n8687), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n11604) );
  NAND2_X1 U11124 ( .A1(n11604), .A2(n12487), .ZN(n8679) );
  NAND2_X1 U11125 ( .A1(n12479), .A2(SI_24_), .ZN(n8678) );
  INV_X1 U11126 ( .A(n8695), .ZN(n8696) );
  NAND2_X1 U11127 ( .A1(n8680), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8681) );
  NAND2_X1 U11128 ( .A1(n8696), .A2(n8681), .ZN(n12940) );
  INV_X1 U11129 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n8684) );
  NAND2_X1 U11130 ( .A1(n8313), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8683) );
  NAND2_X1 U11131 ( .A1(n12489), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8682) );
  OAI211_X1 U11132 ( .C1(n12493), .C2(n8684), .A(n8683), .B(n8682), .ZN(n8685)
         );
  AOI21_X1 U11133 ( .B1(n12940), .B2(n8765), .A(n8685), .ZN(n12948) );
  OR2_X1 U11134 ( .A1(n12941), .A2(n12948), .ZN(n12650) );
  NAND2_X1 U11135 ( .A1(n12941), .A2(n12948), .ZN(n12653) );
  NAND2_X1 U11136 ( .A1(n12650), .A2(n12653), .ZN(n12933) );
  INV_X1 U11137 ( .A(n12948), .ZN(n12920) );
  OR2_X1 U11138 ( .A1(n12941), .A2(n12920), .ZN(n8686) );
  INV_X1 U11139 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n14473) );
  XNOR2_X1 U11140 ( .A(n13803), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8691) );
  XNOR2_X1 U11141 ( .A(n8706), .B(n8691), .ZN(n11693) );
  NAND2_X1 U11142 ( .A1(n11693), .A2(n12487), .ZN(n8693) );
  NAND2_X1 U11143 ( .A1(n12479), .A2(SI_25_), .ZN(n8692) );
  INV_X1 U11144 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8694) );
  INV_X1 U11145 ( .A(n8713), .ZN(n8714) );
  NAND2_X1 U11146 ( .A1(n8696), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8697) );
  NAND2_X1 U11147 ( .A1(n8714), .A2(n8697), .ZN(n12924) );
  NAND2_X1 U11148 ( .A1(n12924), .A2(n8765), .ZN(n8703) );
  INV_X1 U11149 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n8700) );
  NAND2_X1 U11150 ( .A1(n8313), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8699) );
  NAND2_X1 U11151 ( .A1(n12489), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8698) );
  OAI211_X1 U11152 ( .C1(n12493), .C2(n8700), .A(n8699), .B(n8698), .ZN(n8701)
         );
  INV_X1 U11153 ( .A(n8701), .ZN(n8702) );
  OR2_X1 U11154 ( .A1(n13066), .A2(n12936), .ZN(n12658) );
  NAND2_X1 U11155 ( .A1(n13066), .A2(n12936), .ZN(n12659) );
  NAND2_X1 U11156 ( .A1(n12658), .A2(n12659), .ZN(n12918) );
  NAND2_X1 U11157 ( .A1(n13066), .A2(n12904), .ZN(n8704) );
  NOR2_X1 U11158 ( .A1(n13803), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8705) );
  NAND2_X1 U11159 ( .A1(n13803), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8707) );
  XNOR2_X1 U11160 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .ZN(n8709) );
  XNOR2_X1 U11161 ( .A(n8724), .B(n8709), .ZN(n11797) );
  NAND2_X1 U11162 ( .A1(n11797), .A2(n12487), .ZN(n8711) );
  NAND2_X1 U11163 ( .A1(n12479), .A2(SI_26_), .ZN(n8710) );
  INV_X1 U11164 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n8712) );
  NAND2_X1 U11165 ( .A1(n8714), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8715) );
  NAND2_X1 U11166 ( .A1(n8729), .A2(n8715), .ZN(n12911) );
  NAND2_X1 U11167 ( .A1(n12911), .A2(n8765), .ZN(n8721) );
  INV_X1 U11168 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n8718) );
  NAND2_X1 U11169 ( .A1(n12489), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8717) );
  NAND2_X1 U11170 ( .A1(n8313), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8716) );
  OAI211_X1 U11171 ( .C1(n8718), .C2(n12493), .A(n8717), .B(n8716), .ZN(n8719)
         );
  INV_X1 U11172 ( .A(n8719), .ZN(n8720) );
  NAND2_X1 U11173 ( .A1(n12464), .A2(n12921), .ZN(n8722) );
  AND2_X1 U11174 ( .A1(n13799), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U11175 ( .A1(n14462), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8725) );
  XNOR2_X1 U11176 ( .A(n13797), .B(P2_DATAO_REG_27__SCAN_IN), .ZN(n8726) );
  XNOR2_X1 U11177 ( .A(n8739), .B(n8726), .ZN(n11875) );
  NAND2_X1 U11178 ( .A1(n11875), .A2(n12487), .ZN(n8728) );
  NAND2_X1 U11179 ( .A1(n12479), .A2(SI_27_), .ZN(n8727) );
  NAND2_X1 U11180 ( .A1(n8729), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8730) );
  NAND2_X1 U11181 ( .A1(n8745), .A2(n8730), .ZN(n12897) );
  NAND2_X1 U11182 ( .A1(n12897), .A2(n8765), .ZN(n8736) );
  INV_X1 U11183 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n8733) );
  NAND2_X1 U11184 ( .A1(n12489), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8732) );
  NAND2_X1 U11185 ( .A1(n8313), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8731) );
  OAI211_X1 U11186 ( .C1(n8733), .C2(n12493), .A(n8732), .B(n8731), .ZN(n8734)
         );
  INV_X1 U11187 ( .A(n8734), .ZN(n8735) );
  INV_X1 U11188 ( .A(n12890), .ZN(n8737) );
  OR2_X1 U11189 ( .A1(n12667), .A2(n12905), .ZN(n8738) );
  NAND2_X1 U11190 ( .A1(n13797), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8740) );
  AOI22_X1 U11191 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n8842), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n14458), .ZN(n8742) );
  XNOR2_X1 U11192 ( .A(n8843), .B(n8742), .ZN(n11976) );
  NAND2_X1 U11193 ( .A1(n11976), .A2(n12487), .ZN(n8744) );
  NAND2_X1 U11194 ( .A1(n12479), .A2(SI_28_), .ZN(n8743) );
  AND2_X1 U11195 ( .A1(n8745), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8746) );
  NAND2_X1 U11196 ( .A1(n12880), .A2(n8765), .ZN(n8753) );
  NAND2_X1 U11197 ( .A1(n12489), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8749) );
  NAND2_X1 U11198 ( .A1(n8747), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8748) );
  OAI211_X1 U11199 ( .C1(n8750), .C2(n8836), .A(n8749), .B(n8748), .ZN(n8751)
         );
  INV_X1 U11200 ( .A(n8751), .ZN(n8752) );
  NAND2_X1 U11201 ( .A1(n8840), .A2(n8848), .ZN(n8859) );
  NAND2_X1 U11202 ( .A1(n12671), .A2(n8859), .ZN(n12676) );
  NAND2_X1 U11203 ( .A1(n8764), .A2(n12670), .ZN(n8763) );
  NAND2_X1 U11204 ( .A1(n6514), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8754) );
  NAND2_X1 U11205 ( .A1(n12501), .A2(n12695), .ZN(n8827) );
  INV_X1 U11206 ( .A(n8527), .ZN(n8757) );
  INV_X1 U11207 ( .A(n8755), .ZN(n8756) );
  NAND2_X1 U11208 ( .A1(n8760), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8761) );
  MUX2_X1 U11209 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8761), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n8762) );
  NAND2_X1 U11210 ( .A1(n8868), .A2(n12524), .ZN(n12690) );
  NAND2_X1 U11211 ( .A1(n8763), .A2(n15112), .ZN(n8773) );
  NAND2_X1 U11212 ( .A1(n12872), .A2(n8765), .ZN(n12496) );
  INV_X1 U11213 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n8768) );
  NAND2_X1 U11214 ( .A1(n12489), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8767) );
  NAND2_X1 U11215 ( .A1(n8313), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8766) );
  OAI211_X1 U11216 ( .C1(n8768), .C2(n12493), .A(n8767), .B(n8766), .ZN(n8769)
         );
  INV_X1 U11217 ( .A(n8769), .ZN(n8770) );
  NAND2_X1 U11218 ( .A1(n12496), .A2(n8770), .ZN(n12700) );
  INV_X1 U11219 ( .A(n6870), .ZN(n12692) );
  INV_X1 U11220 ( .A(n8771), .ZN(n12846) );
  NAND2_X1 U11221 ( .A1(n12692), .A2(n12846), .ZN(n10250) );
  NAND2_X1 U11222 ( .A1(n10250), .A2(n10243), .ZN(n8968) );
  INV_X1 U11223 ( .A(n8968), .ZN(n8969) );
  AOI22_X1 U11224 ( .A1(n12700), .A2(n15106), .B1(n15109), .B2(n12905), .ZN(
        n8772) );
  OAI21_X2 U11225 ( .B1(n8773), .B2(n8841), .A(n8772), .ZN(n12883) );
  NAND2_X1 U11226 ( .A1(n15105), .A2(n12532), .ZN(n8890) );
  NAND2_X1 U11227 ( .A1(n8890), .A2(n8883), .ZN(n15087) );
  NAND2_X1 U11228 ( .A1(n8774), .A2(n12541), .ZN(n10893) );
  NAND2_X1 U11229 ( .A1(n10893), .A2(n12505), .ZN(n8775) );
  INV_X1 U11230 ( .A(n12547), .ZN(n8776) );
  NAND2_X1 U11231 ( .A1(n10935), .A2(n8776), .ZN(n8777) );
  NAND2_X1 U11232 ( .A1(n8777), .A2(n12550), .ZN(n15068) );
  NAND2_X1 U11233 ( .A1(n15068), .A2(n15072), .ZN(n8778) );
  NAND2_X1 U11234 ( .A1(n8778), .A2(n12555), .ZN(n11307) );
  INV_X1 U11235 ( .A(n11309), .ZN(n12504) );
  NAND2_X1 U11236 ( .A1(n11307), .A2(n12504), .ZN(n8779) );
  NAND2_X1 U11237 ( .A1(n8779), .A2(n12564), .ZN(n11229) );
  NAND2_X1 U11238 ( .A1(n11229), .A2(n12562), .ZN(n8780) );
  INV_X1 U11239 ( .A(n12710), .ZN(n11361) );
  NAND2_X1 U11240 ( .A1(n11361), .A2(n11236), .ZN(n12567) );
  NOR2_X1 U11241 ( .A1(n12708), .A2(n11624), .ZN(n8781) );
  INV_X1 U11242 ( .A(n12508), .ZN(n12587) );
  NAND2_X1 U11243 ( .A1(n11683), .A2(n12587), .ZN(n8782) );
  NAND2_X1 U11244 ( .A1(n12707), .A2(n15168), .ZN(n12584) );
  NAND2_X1 U11245 ( .A1(n14677), .A2(n14657), .ZN(n12589) );
  NAND2_X1 U11246 ( .A1(n12590), .A2(n12589), .ZN(n14671) );
  INV_X1 U11247 ( .A(n14650), .ZN(n8784) );
  OR2_X1 U11248 ( .A1(n12036), .A2(n8921), .ZN(n12599) );
  INV_X1 U11249 ( .A(n12253), .ZN(n12512) );
  NAND2_X1 U11250 ( .A1(n12257), .A2(n12512), .ZN(n8786) );
  NAND2_X1 U11251 ( .A1(n8786), .A2(n12614), .ZN(n13040) );
  NAND2_X1 U11252 ( .A1(n13040), .A2(n13039), .ZN(n8787) );
  NAND2_X1 U11253 ( .A1(n8787), .A2(n12618), .ZN(n13029) );
  OR2_X2 U11254 ( .A1(n13029), .A2(n13028), .ZN(n13100) );
  INV_X1 U11255 ( .A(n12622), .ZN(n13009) );
  NOR2_X1 U11256 ( .A1(n13008), .A2(n13009), .ZN(n8788) );
  INV_X1 U11257 ( .A(n12988), .ZN(n12963) );
  NAND2_X1 U11258 ( .A1(n12387), .A2(n12963), .ZN(n12639) );
  NAND2_X1 U11259 ( .A1(n12977), .A2(n12639), .ZN(n8789) );
  OR2_X1 U11260 ( .A1(n12387), .A2(n12963), .ZN(n12638) );
  NAND2_X1 U11261 ( .A1(n8789), .A2(n12638), .ZN(n12965) );
  NAND2_X1 U11262 ( .A1(n12966), .A2(n12975), .ZN(n12642) );
  NAND2_X1 U11263 ( .A1(n12965), .A2(n12642), .ZN(n8790) );
  NAND2_X1 U11264 ( .A1(n8790), .A2(n12643), .ZN(n12954) );
  INV_X1 U11265 ( .A(n12701), .ZN(n12962) );
  OR2_X1 U11266 ( .A1(n12952), .A2(n12962), .ZN(n12649) );
  NAND2_X1 U11267 ( .A1(n12931), .A2(n12653), .ZN(n12916) );
  INV_X1 U11268 ( .A(n12918), .ZN(n12655) );
  NAND2_X1 U11269 ( .A1(n12916), .A2(n12655), .ZN(n8791) );
  NAND2_X1 U11270 ( .A1(n8791), .A2(n12659), .ZN(n12907) );
  INV_X1 U11271 ( .A(n12921), .ZN(n12404) );
  OR2_X1 U11272 ( .A1(n12464), .A2(n12404), .ZN(n12662) );
  NAND2_X1 U11273 ( .A1(n12907), .A2(n12662), .ZN(n8792) );
  NAND2_X1 U11274 ( .A1(n12464), .A2(n12404), .ZN(n12663) );
  NAND2_X1 U11275 ( .A1(n8792), .A2(n12663), .ZN(n12891) );
  AND2_X2 U11276 ( .A1(n12891), .A2(n12890), .ZN(n12893) );
  INV_X1 U11277 ( .A(n12905), .ZN(n12668) );
  NAND2_X1 U11278 ( .A1(n12667), .A2(n12668), .ZN(n8858) );
  INV_X1 U11279 ( .A(n8858), .ZN(n8793) );
  XNOR2_X1 U11280 ( .A(n8794), .B(n12670), .ZN(n12879) );
  NAND2_X1 U11281 ( .A1(n10890), .A2(n12695), .ZN(n8795) );
  AOI21_X1 U11282 ( .B1(n12501), .B2(n8795), .A(n12524), .ZN(n8797) );
  AOI21_X1 U11283 ( .B1(n10890), .B2(n12529), .A(n12695), .ZN(n8796) );
  OR2_X1 U11284 ( .A1(n8797), .A2(n8796), .ZN(n8971) );
  AND2_X1 U11285 ( .A1(n12859), .A2(n10890), .ZN(n12687) );
  INV_X1 U11286 ( .A(n12695), .ZN(n8798) );
  NAND3_X1 U11287 ( .A1(n8971), .A2(n12687), .A3(n15169), .ZN(n8800) );
  AND2_X1 U11288 ( .A1(n8868), .A2(n12695), .ZN(n8799) );
  NAND2_X1 U11289 ( .A1(n12859), .A2(n8799), .ZN(n8871) );
  OR2_X1 U11290 ( .A1(n15117), .A2(n12695), .ZN(n15148) );
  AND2_X1 U11291 ( .A1(n12879), .A2(n14692), .ZN(n8801) );
  NOR2_X1 U11292 ( .A1(n12883), .A2(n8801), .ZN(n13053) );
  NAND2_X1 U11293 ( .A1(n8804), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8803) );
  INV_X1 U11294 ( .A(n8804), .ZN(n8806) );
  XNOR2_X1 U11295 ( .A(n11607), .B(P3_B_REG_SCAN_IN), .ZN(n8811) );
  NAND2_X1 U11296 ( .A1(n8808), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8809) );
  NAND2_X1 U11297 ( .A1(n6518), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8812) );
  OAI22_X1 U11298 ( .A1(n8815), .A2(P3_D_REG_1__SCAN_IN), .B1(n8813), .B2(
        n8831), .ZN(n10577) );
  INV_X1 U11299 ( .A(n8813), .ZN(n11800) );
  NAND2_X1 U11300 ( .A1(n11607), .A2(n11800), .ZN(n8814) );
  OR2_X1 U11301 ( .A1(n10577), .A2(n8878), .ZN(n8867) );
  INV_X1 U11302 ( .A(n8867), .ZN(n8826) );
  NOR2_X1 U11303 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_4__SCAN_IN), .ZN(
        n8819) );
  NOR4_X1 U11304 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n8818) );
  NOR4_X1 U11305 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8817) );
  NOR4_X1 U11306 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n8816) );
  NAND4_X1 U11307 ( .A1(n8819), .A2(n8818), .A3(n8817), .A4(n8816), .ZN(n8825)
         );
  NOR4_X1 U11308 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n8823) );
  NOR4_X1 U11309 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_21__SCAN_IN), .ZN(n8822) );
  NOR4_X1 U11310 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8821) );
  NOR4_X1 U11311 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n8820) );
  NAND4_X1 U11312 ( .A1(n8823), .A2(n8822), .A3(n8821), .A4(n8820), .ZN(n8824)
         );
  INV_X1 U11313 ( .A(n8815), .ZN(n10028) );
  OAI21_X1 U11314 ( .B1(n8825), .B2(n8824), .A(n10028), .ZN(n8865) );
  NAND2_X1 U11315 ( .A1(n8826), .A2(n8865), .ZN(n8972) );
  NAND2_X1 U11316 ( .A1(n8868), .A2(n12529), .ZN(n12521) );
  OR2_X1 U11317 ( .A1(n8827), .A2(n12521), .ZN(n8958) );
  INV_X1 U11318 ( .A(n8958), .ZN(n8975) );
  AND2_X1 U11319 ( .A1(n12687), .A2(n12657), .ZN(n10519) );
  NOR2_X1 U11320 ( .A1(n8975), .A2(n10519), .ZN(n8829) );
  INV_X1 U11321 ( .A(n8971), .ZN(n8828) );
  NAND3_X1 U11322 ( .A1(n10577), .A2(n8878), .A3(n8865), .ZN(n8980) );
  OAI22_X1 U11323 ( .A1(n8972), .A2(n8829), .B1(n8828), .B2(n8980), .ZN(n8835)
         );
  NOR2_X1 U11324 ( .A1(n11607), .A2(n11800), .ZN(n8830) );
  NAND2_X1 U11325 ( .A1(n8831), .A2(n8830), .ZN(n9916) );
  NAND2_X1 U11326 ( .A1(n8832), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8834) );
  MUX2_X1 U11327 ( .A(n8836), .B(n13053), .S(n15176), .Z(n8839) );
  NAND2_X1 U11328 ( .A1(n8840), .A2(n8837), .ZN(n8838) );
  NAND2_X1 U11329 ( .A1(n8839), .A2(n8838), .ZN(P3_U3455) );
  NAND2_X1 U11330 ( .A1(n14458), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8844) );
  INV_X1 U11331 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n12282) );
  XNOR2_X1 U11332 ( .A(n12282), .B(P2_DATAO_REG_29__SCAN_IN), .ZN(n12286) );
  XNOR2_X1 U11333 ( .A(n12288), .B(n12286), .ZN(n13173) );
  NAND2_X1 U11334 ( .A1(n13173), .A2(n12487), .ZN(n8846) );
  NAND2_X1 U11335 ( .A1(n12479), .A2(SI_29_), .ZN(n8845) );
  NAND2_X1 U11336 ( .A1(n8846), .A2(n8845), .ZN(n8860) );
  INV_X1 U11337 ( .A(n12700), .ZN(n8847) );
  NAND2_X1 U11338 ( .A1(n8860), .A2(n8847), .ZN(n12678) );
  NAND2_X1 U11339 ( .A1(n12682), .A2(n12678), .ZN(n12502) );
  INV_X1 U11340 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n8851) );
  NAND2_X1 U11341 ( .A1(n8313), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8850) );
  NAND2_X1 U11342 ( .A1(n12489), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8849) );
  OAI211_X1 U11343 ( .C1(n12493), .C2(n8851), .A(n8850), .B(n8849), .ZN(n8852)
         );
  INV_X1 U11344 ( .A(n8852), .ZN(n8853) );
  AND2_X1 U11345 ( .A1(n12496), .A2(n8853), .ZN(n12498) );
  INV_X1 U11346 ( .A(P3_B_REG_SCAN_IN), .ZN(n8854) );
  OAI21_X1 U11347 ( .B1(n6870), .B2(n8854), .A(n15106), .ZN(n12865) );
  NOR2_X1 U11348 ( .A1(n12498), .A2(n12865), .ZN(n8855) );
  NAND2_X1 U11349 ( .A1(n8859), .A2(n8858), .ZN(n12673) );
  OAI21_X2 U11350 ( .B1(n12893), .B2(n12673), .A(n12671), .ZN(n12497) );
  XNOR2_X1 U11351 ( .A(n12497), .B(n12502), .ZN(n12876) );
  INV_X1 U11352 ( .A(n8860), .ZN(n12874) );
  INV_X1 U11353 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8861) );
  OAI21_X1 U11354 ( .B1(n8877), .B2(n15174), .A(n8863), .ZN(P3_U3456) );
  INV_X1 U11355 ( .A(n12687), .ZN(n8864) );
  NAND2_X1 U11356 ( .A1(n8864), .A2(n12657), .ZN(n8973) );
  AND3_X1 U11357 ( .A1(n8973), .A2(n8865), .A3(n8967), .ZN(n8866) );
  NOR2_X1 U11358 ( .A1(n15169), .A2(n8868), .ZN(n8869) );
  AOI21_X1 U11359 ( .B1(n12859), .B2(n12695), .A(n8869), .ZN(n8870) );
  OAI21_X1 U11360 ( .B1(n8870), .B2(n12687), .A(n12675), .ZN(n8872) );
  OAI22_X1 U11361 ( .A1(n8872), .A2(n8878), .B1(n10578), .B2(n10577), .ZN(
        n8873) );
  INV_X1 U11362 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n15348) );
  OR2_X1 U11363 ( .A1(n15193), .A2(n15348), .ZN(n8874) );
  OAI21_X1 U11364 ( .B1(n8877), .B2(n15190), .A(n8876), .ZN(P3_U3488) );
  INV_X1 U11365 ( .A(n12521), .ZN(n8879) );
  NAND2_X1 U11366 ( .A1(n13166), .A2(n8879), .ZN(n8882) );
  OAI21_X1 U11367 ( .B1(n8880), .B2(n12524), .A(n10890), .ZN(n8881) );
  NAND2_X2 U11368 ( .A1(n8882), .A2(n8881), .ZN(n8893) );
  XNOR2_X1 U11369 ( .A(n13158), .B(n8957), .ZN(n8926) );
  INV_X1 U11370 ( .A(n8926), .ZN(n8927) );
  XNOR2_X1 U11371 ( .A(n12152), .B(n10646), .ZN(n8925) );
  NAND2_X1 U11372 ( .A1(n8883), .A2(n8957), .ZN(n8886) );
  NAND2_X1 U11373 ( .A1(n8884), .A2(n8956), .ZN(n8885) );
  NAND2_X1 U11374 ( .A1(n8886), .A2(n8885), .ZN(n8891) );
  NAND3_X1 U11375 ( .A1(n8956), .A2(n10730), .A3(n8887), .ZN(n8888) );
  NAND2_X1 U11376 ( .A1(n8956), .A2(n15110), .ZN(n8889) );
  XNOR2_X1 U11377 ( .A(n8892), .B(n8893), .ZN(n8894) );
  XNOR2_X1 U11378 ( .A(n15107), .B(n8894), .ZN(n10729) );
  NAND2_X1 U11379 ( .A1(n8894), .A2(n10894), .ZN(n8895) );
  NAND2_X1 U11380 ( .A1(n8896), .A2(n8895), .ZN(n10686) );
  INV_X1 U11381 ( .A(n10686), .ZN(n8897) );
  XNOR2_X1 U11382 ( .A(n8893), .B(n10901), .ZN(n8898) );
  XNOR2_X1 U11383 ( .A(n8898), .B(n12712), .ZN(n10687) );
  NAND2_X1 U11384 ( .A1(n8898), .A2(n12712), .ZN(n8899) );
  XNOR2_X1 U11385 ( .A(n8893), .B(n8900), .ZN(n8901) );
  XNOR2_X1 U11386 ( .A(n8901), .B(n15074), .ZN(n10816) );
  NAND2_X1 U11387 ( .A1(n8901), .A2(n10909), .ZN(n8902) );
  XNOR2_X1 U11388 ( .A(n8957), .B(n15081), .ZN(n8903) );
  XNOR2_X1 U11389 ( .A(n8903), .B(n12711), .ZN(n10906) );
  NAND2_X1 U11390 ( .A1(n8903), .A2(n11092), .ZN(n8904) );
  XNOR2_X1 U11391 ( .A(n8957), .B(n15147), .ZN(n8905) );
  XNOR2_X1 U11392 ( .A(n8905), .B(n15073), .ZN(n11089) );
  NAND2_X1 U11393 ( .A1(n8905), .A2(n15073), .ZN(n8906) );
  XNOR2_X1 U11394 ( .A(n12562), .B(n8957), .ZN(n11206) );
  INV_X1 U11395 ( .A(n11206), .ZN(n8907) );
  NAND2_X1 U11396 ( .A1(n8907), .A2(n12710), .ZN(n8908) );
  XNOR2_X1 U11397 ( .A(n8957), .B(n11575), .ZN(n8909) );
  XNOR2_X1 U11398 ( .A(n8909), .B(n12709), .ZN(n11358) );
  INV_X1 U11399 ( .A(n8909), .ZN(n8910) );
  NAND2_X1 U11400 ( .A1(n8910), .A2(n12709), .ZN(n8911) );
  XNOR2_X1 U11401 ( .A(n8957), .B(n11624), .ZN(n8912) );
  XNOR2_X1 U11402 ( .A(n8912), .B(n12708), .ZN(n11559) );
  INV_X1 U11403 ( .A(n8912), .ZN(n8913) );
  XNOR2_X1 U11404 ( .A(n15168), .B(n10646), .ZN(n8914) );
  XNOR2_X1 U11405 ( .A(n8914), .B(n14674), .ZN(n11652) );
  NAND2_X1 U11406 ( .A1(n8914), .A2(n12707), .ZN(n8915) );
  XNOR2_X1 U11407 ( .A(n14677), .B(n10646), .ZN(n8916) );
  NAND2_X1 U11408 ( .A1(n8917), .A2(n8916), .ZN(n11879) );
  INV_X1 U11409 ( .A(n11892), .ZN(n8920) );
  XNOR2_X1 U11410 ( .A(n14663), .B(n10646), .ZN(n11890) );
  OAI21_X1 U11411 ( .B1(n11892), .B2(n12706), .A(n11890), .ZN(n8919) );
  XNOR2_X1 U11412 ( .A(n12036), .B(n10646), .ZN(n8922) );
  NOR2_X1 U11413 ( .A1(n8922), .A2(n8921), .ZN(n12029) );
  XNOR2_X1 U11414 ( .A(n12243), .B(n10646), .ZN(n8923) );
  XOR2_X1 U11415 ( .A(n12705), .B(n8923), .Z(n12120) );
  INV_X1 U11416 ( .A(n8923), .ZN(n8924) );
  XNOR2_X1 U11417 ( .A(n8925), .B(n12704), .ZN(n12154) );
  XNOR2_X1 U11418 ( .A(n8926), .B(n13035), .ZN(n12410) );
  XOR2_X1 U11419 ( .A(n8957), .B(n13041), .Z(n12419) );
  INV_X1 U11420 ( .A(n12419), .ZN(n8928) );
  NAND2_X1 U11421 ( .A1(n8928), .A2(n12418), .ZN(n8929) );
  XNOR2_X1 U11422 ( .A(n13098), .B(n10646), .ZN(n8930) );
  XOR2_X1 U11423 ( .A(n13036), .B(n8930), .Z(n12454) );
  XNOR2_X1 U11424 ( .A(n13151), .B(n10646), .ZN(n8932) );
  XOR2_X1 U11425 ( .A(n13022), .B(n8932), .Z(n12380) );
  XNOR2_X1 U11426 ( .A(n13090), .B(n8956), .ZN(n8933) );
  NOR2_X1 U11427 ( .A1(n8933), .A2(n13004), .ZN(n12390) );
  AOI21_X1 U11428 ( .B1(n8933), .B2(n13004), .A(n12390), .ZN(n12435) );
  XNOR2_X1 U11429 ( .A(n12387), .B(n8957), .ZN(n8934) );
  XNOR2_X1 U11430 ( .A(n8934), .B(n12988), .ZN(n12389) );
  NAND2_X1 U11431 ( .A1(n12388), .A2(n8935), .ZN(n8937) );
  XNOR2_X1 U11432 ( .A(n12966), .B(n10646), .ZN(n8936) );
  NAND2_X1 U11433 ( .A1(n12447), .A2(n8938), .ZN(n8942) );
  INV_X1 U11434 ( .A(n8942), .ZN(n8940) );
  INV_X1 U11435 ( .A(n8941), .ZN(n8939) );
  NAND2_X1 U11436 ( .A1(n8940), .A2(n8939), .ZN(n8943) );
  NAND2_X1 U11437 ( .A1(n8943), .A2(n12429), .ZN(n12372) );
  INV_X1 U11438 ( .A(n12372), .ZN(n8944) );
  XNOR2_X1 U11439 ( .A(n12941), .B(n10646), .ZN(n8945) );
  NAND2_X1 U11440 ( .A1(n8945), .A2(n12948), .ZN(n8948) );
  INV_X1 U11441 ( .A(n8945), .ZN(n8946) );
  NAND2_X1 U11442 ( .A1(n8946), .A2(n12920), .ZN(n8947) );
  NAND2_X1 U11443 ( .A1(n8948), .A2(n8947), .ZN(n12428) );
  INV_X1 U11444 ( .A(n8948), .ZN(n12400) );
  XNOR2_X1 U11445 ( .A(n13066), .B(n10646), .ZN(n8949) );
  NAND2_X1 U11446 ( .A1(n8949), .A2(n12936), .ZN(n8952) );
  INV_X1 U11447 ( .A(n8949), .ZN(n8950) );
  NAND2_X1 U11448 ( .A1(n8950), .A2(n12904), .ZN(n8951) );
  XNOR2_X1 U11449 ( .A(n12464), .B(n8956), .ZN(n8953) );
  NOR2_X1 U11450 ( .A1(n8953), .A2(n12921), .ZN(n8954) );
  AOI21_X1 U11451 ( .B1(n8953), .B2(n12921), .A(n8954), .ZN(n12467) );
  INV_X1 U11452 ( .A(n8954), .ZN(n8955) );
  XNOR2_X1 U11453 ( .A(n12667), .B(n8956), .ZN(n8964) );
  NOR2_X1 U11454 ( .A1(n8964), .A2(n12905), .ZN(n8961) );
  AOI21_X1 U11455 ( .B1(n8964), .B2(n12905), .A(n8961), .ZN(n9274) );
  XNOR2_X1 U11456 ( .A(n12676), .B(n8957), .ZN(n8965) );
  INV_X1 U11457 ( .A(n8965), .ZN(n8962) );
  NAND2_X1 U11458 ( .A1(n8971), .A2(n15169), .ZN(n8959) );
  OAI22_X1 U11459 ( .A1(n8972), .A2(n8959), .B1(n8958), .B2(n8980), .ZN(n8960)
         );
  NAND2_X1 U11460 ( .A1(n8962), .A2(n12468), .ZN(n8989) );
  NOR3_X1 U11461 ( .A1(n8962), .A2(n8961), .A3(n12462), .ZN(n8963) );
  NOR4_X1 U11462 ( .A1(n8965), .A2(n8964), .A3(n12462), .A4(n12905), .ZN(n8986) );
  NAND2_X1 U11463 ( .A1(n8972), .A2(n15117), .ZN(n8966) );
  INV_X1 U11464 ( .A(n8967), .ZN(n10240) );
  NOR2_X1 U11465 ( .A1(n10240), .A2(n15169), .ZN(n10581) );
  NAND2_X2 U11466 ( .A1(n8966), .A2(n10581), .ZN(n12477) );
  NAND2_X1 U11467 ( .A1(n10519), .A2(n8967), .ZN(n8979) );
  OR2_X1 U11468 ( .A1(n8979), .A2(n8980), .ZN(n8970) );
  NOR2_X2 U11469 ( .A1(n8970), .A2(n8968), .ZN(n12470) );
  AOI22_X1 U11470 ( .A1(n12905), .A2(n12470), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n8984) );
  NOR2_X2 U11471 ( .A1(n8970), .A2(n8969), .ZN(n12439) );
  NAND2_X1 U11472 ( .A1(n8972), .A2(n8971), .ZN(n8977) );
  NAND3_X1 U11473 ( .A1(n8973), .A2(n9916), .A3(n10241), .ZN(n8974) );
  AOI21_X1 U11474 ( .B1(n8980), .B2(n8975), .A(n8974), .ZN(n8976) );
  NAND2_X1 U11475 ( .A1(n8977), .A2(n8976), .ZN(n8978) );
  NAND2_X1 U11476 ( .A1(n8978), .A2(P3_STATE_REG_SCAN_IN), .ZN(n8982) );
  INV_X1 U11477 ( .A(n8979), .ZN(n12693) );
  NAND2_X1 U11478 ( .A1(n12693), .A2(n8980), .ZN(n8981) );
  AOI22_X1 U11479 ( .A1(n12700), .A2(n12439), .B1(n12880), .B2(n12474), .ZN(
        n8983) );
  OAI211_X1 U11480 ( .C1(n13056), .C2(n12477), .A(n8984), .B(n8983), .ZN(n8985) );
  OAI211_X1 U11481 ( .C1(n9272), .C2(n8989), .A(n8988), .B(n8987), .ZN(
        P3_U3160) );
  INV_X2 U11482 ( .A(n8996), .ZN(n9017) );
  NAND2_X1 U11483 ( .A1(n9002), .A2(n9168), .ZN(n8991) );
  NAND2_X1 U11484 ( .A1(n8991), .A2(n8990), .ZN(n9006) );
  NAND2_X1 U11485 ( .A1(n9923), .A2(n6864), .ZN(n8992) );
  NAND2_X1 U11486 ( .A1(n8993), .A2(n8992), .ZN(n8997) );
  OAI21_X1 U11487 ( .B1(n10323), .B2(n8997), .A(n8994), .ZN(n8995) );
  INV_X1 U11488 ( .A(n8995), .ZN(n9001) );
  NAND2_X1 U11489 ( .A1(n10421), .A2(n8996), .ZN(n8999) );
  NAND3_X1 U11490 ( .A1(n10323), .A2(n6472), .A3(n8997), .ZN(n8998) );
  INV_X1 U11491 ( .A(n8996), .ZN(n9152) );
  NAND2_X1 U11492 ( .A1(n9002), .A2(n9213), .ZN(n9003) );
  NAND2_X1 U11493 ( .A1(n9004), .A2(n9003), .ZN(n9005) );
  INV_X1 U11494 ( .A(n9006), .ZN(n9009) );
  INV_X1 U11495 ( .A(n9007), .ZN(n9008) );
  NAND2_X1 U11496 ( .A1(n9009), .A2(n9008), .ZN(n9010) );
  NAND2_X1 U11497 ( .A1(n13311), .A2(n9213), .ZN(n9013) );
  NAND2_X1 U11498 ( .A1(n10915), .A2(n9168), .ZN(n9012) );
  NAND2_X1 U11499 ( .A1(n9013), .A2(n9012), .ZN(n9015) );
  AOI22_X1 U11500 ( .A1(n13311), .A2(n9214), .B1(n10915), .B2(n6473), .ZN(
        n9014) );
  NAND2_X1 U11501 ( .A1(n13310), .A2(n9214), .ZN(n9019) );
  NAND2_X1 U11502 ( .A1(n10953), .A2(n9152), .ZN(n9018) );
  NAND2_X1 U11503 ( .A1(n9019), .A2(n9018), .ZN(n9020) );
  AOI22_X1 U11504 ( .A1(n13310), .A2(n9152), .B1(n10953), .B2(n9168), .ZN(
        n9022) );
  NAND2_X1 U11505 ( .A1(n14984), .A2(n9214), .ZN(n9026) );
  NAND2_X1 U11506 ( .A1(n13309), .A2(n9213), .ZN(n9025) );
  NAND2_X1 U11507 ( .A1(n9026), .A2(n9025), .ZN(n9028) );
  AOI22_X1 U11508 ( .A1(n14984), .A2(n9152), .B1(n9214), .B2(n13309), .ZN(
        n9027) );
  NAND2_X1 U11509 ( .A1(n11071), .A2(n9213), .ZN(n9031) );
  NAND2_X1 U11510 ( .A1(n13308), .A2(n9214), .ZN(n9030) );
  NAND2_X1 U11511 ( .A1(n9031), .A2(n9030), .ZN(n9033) );
  AOI22_X1 U11512 ( .A1(n11071), .A2(n9214), .B1(n13308), .B2(n9152), .ZN(
        n9032) );
  NAND2_X1 U11513 ( .A1(n14991), .A2(n9214), .ZN(n9036) );
  NAND2_X1 U11514 ( .A1(n13307), .A2(n9213), .ZN(n9035) );
  NAND2_X1 U11515 ( .A1(n9036), .A2(n9035), .ZN(n9040) );
  INV_X1 U11516 ( .A(n13307), .ZN(n11156) );
  NAND2_X1 U11517 ( .A1(n14991), .A2(n9213), .ZN(n9037) );
  OAI21_X1 U11518 ( .B1(n11156), .B2(n9213), .A(n9037), .ZN(n9038) );
  INV_X1 U11519 ( .A(n9040), .ZN(n9041) );
  NAND2_X1 U11520 ( .A1(n14954), .A2(n9213), .ZN(n9043) );
  NAND2_X1 U11521 ( .A1(n13306), .A2(n9214), .ZN(n9042) );
  NAND2_X1 U11522 ( .A1(n9043), .A2(n9042), .ZN(n9045) );
  AOI22_X1 U11523 ( .A1(n14954), .A2(n9214), .B1(n13306), .B2(n9152), .ZN(
        n9044) );
  NAND2_X1 U11524 ( .A1(n11437), .A2(n9168), .ZN(n9048) );
  NAND2_X1 U11525 ( .A1(n13305), .A2(n9213), .ZN(n9047) );
  NAND2_X1 U11526 ( .A1(n9048), .A2(n9047), .ZN(n9053) );
  INV_X1 U11527 ( .A(n13305), .ZN(n11401) );
  NAND2_X1 U11528 ( .A1(n11437), .A2(n9213), .ZN(n9049) );
  NAND2_X1 U11529 ( .A1(n9051), .A2(n9050), .ZN(n9057) );
  INV_X1 U11530 ( .A(n9052), .ZN(n9055) );
  NAND2_X1 U11531 ( .A1(n9055), .A2(n9054), .ZN(n9056) );
  NAND2_X1 U11532 ( .A1(n11554), .A2(n9152), .ZN(n9059) );
  NAND2_X1 U11533 ( .A1(n13304), .A2(n9214), .ZN(n9058) );
  NAND2_X1 U11534 ( .A1(n9059), .A2(n9058), .ZN(n9062) );
  AOI22_X1 U11535 ( .A1(n11554), .A2(n9168), .B1(n13304), .B2(n9152), .ZN(
        n9060) );
  INV_X1 U11536 ( .A(n9060), .ZN(n9061) );
  NAND2_X1 U11537 ( .A1(n11663), .A2(n9168), .ZN(n9064) );
  NAND2_X1 U11538 ( .A1(n13303), .A2(n9152), .ZN(n9063) );
  NAND2_X1 U11539 ( .A1(n9064), .A2(n9063), .ZN(n9067) );
  AOI22_X1 U11540 ( .A1(n11663), .A2(n9152), .B1(n9214), .B2(n13303), .ZN(
        n9065) );
  NAND2_X1 U11541 ( .A1(n11816), .A2(n9152), .ZN(n9070) );
  NAND2_X1 U11542 ( .A1(n13302), .A2(n9168), .ZN(n9069) );
  NAND2_X1 U11543 ( .A1(n9070), .A2(n9069), .ZN(n9075) );
  INV_X1 U11544 ( .A(n13302), .ZN(n11815) );
  NAND2_X1 U11545 ( .A1(n11816), .A2(n9214), .ZN(n9071) );
  OAI21_X1 U11546 ( .B1(n11815), .B2(n9214), .A(n9071), .ZN(n9072) );
  NAND2_X1 U11547 ( .A1(n9073), .A2(n9072), .ZN(n9079) );
  INV_X1 U11548 ( .A(n9074), .ZN(n9077) );
  INV_X1 U11549 ( .A(n9075), .ZN(n9076) );
  NAND2_X1 U11550 ( .A1(n9077), .A2(n9076), .ZN(n9078) );
  NAND2_X1 U11551 ( .A1(n13221), .A2(n9168), .ZN(n9081) );
  NAND2_X1 U11552 ( .A1(n13301), .A2(n9213), .ZN(n9080) );
  NAND2_X1 U11553 ( .A1(n9081), .A2(n9080), .ZN(n9083) );
  AOI22_X1 U11554 ( .A1(n13221), .A2(n9152), .B1(n9214), .B2(n13301), .ZN(
        n9082) );
  NAND2_X1 U11555 ( .A1(n14868), .A2(n9152), .ZN(n9086) );
  NAND2_X1 U11556 ( .A1(n13300), .A2(n9168), .ZN(n9085) );
  NAND2_X1 U11557 ( .A1(n9086), .A2(n9085), .ZN(n9088) );
  AOI22_X1 U11558 ( .A1(n14868), .A2(n9214), .B1(n13300), .B2(n6473), .ZN(
        n9087) );
  AND2_X1 U11559 ( .A1(n13299), .A2(n9214), .ZN(n9089) );
  AOI21_X1 U11560 ( .B1(n13744), .B2(n9152), .A(n9089), .ZN(n9102) );
  NAND2_X1 U11561 ( .A1(n13744), .A2(n9168), .ZN(n9091) );
  NAND2_X1 U11562 ( .A1(n13299), .A2(n9152), .ZN(n9090) );
  NAND2_X1 U11563 ( .A1(n9091), .A2(n9090), .ZN(n9101) );
  AND2_X1 U11564 ( .A1(n13394), .A2(n9214), .ZN(n9092) );
  AOI21_X1 U11565 ( .B1(n13727), .B2(n9152), .A(n9092), .ZN(n9115) );
  NAND2_X1 U11566 ( .A1(n13727), .A2(n9168), .ZN(n9094) );
  NAND2_X1 U11567 ( .A1(n13394), .A2(n9152), .ZN(n9093) );
  NAND2_X1 U11568 ( .A1(n9094), .A2(n9093), .ZN(n9113) );
  AND2_X1 U11569 ( .A1(n13391), .A2(n9214), .ZN(n9095) );
  AOI21_X1 U11570 ( .B1(n13419), .B2(n9152), .A(n9095), .ZN(n9110) );
  NAND2_X1 U11571 ( .A1(n13419), .A2(n9214), .ZN(n9097) );
  NAND2_X1 U11572 ( .A1(n13391), .A2(n9152), .ZN(n9096) );
  NAND2_X1 U11573 ( .A1(n9097), .A2(n9096), .ZN(n9109) );
  AOI22_X1 U11574 ( .A1(n9115), .A2(n9113), .B1(n9110), .B2(n9109), .ZN(n9105)
         );
  AND2_X1 U11575 ( .A1(n13298), .A2(n9214), .ZN(n9098) );
  AOI21_X1 U11576 ( .B1(n13782), .B2(n9017), .A(n9098), .ZN(n9107) );
  NAND2_X1 U11577 ( .A1(n13782), .A2(n9168), .ZN(n9100) );
  NAND2_X1 U11578 ( .A1(n13298), .A2(n9017), .ZN(n9099) );
  NAND2_X1 U11579 ( .A1(n9100), .A2(n9099), .ZN(n9106) );
  AOI22_X1 U11580 ( .A1(n9107), .A2(n9106), .B1(n9102), .B2(n9101), .ZN(n9103)
         );
  INV_X1 U11581 ( .A(n9105), .ZN(n9108) );
  INV_X1 U11582 ( .A(n9109), .ZN(n9112) );
  INV_X1 U11583 ( .A(n9110), .ZN(n9111) );
  NAND2_X1 U11584 ( .A1(n9112), .A2(n9111), .ZN(n9114) );
  INV_X1 U11585 ( .A(n13394), .ZN(n13423) );
  INV_X1 U11586 ( .A(n13727), .ZN(n13641) );
  NAND3_X1 U11587 ( .A1(n9114), .A2(n13423), .A3(n13641), .ZN(n9119) );
  INV_X1 U11588 ( .A(n9113), .ZN(n9118) );
  INV_X1 U11589 ( .A(n9114), .ZN(n9117) );
  INV_X1 U11590 ( .A(n9115), .ZN(n9116) );
  AOI22_X1 U11591 ( .A1(n9119), .A2(n9118), .B1(n9117), .B2(n9116), .ZN(n9120)
         );
  AND2_X1 U11592 ( .A1(n9121), .A2(n9120), .ZN(n9122) );
  AND2_X1 U11593 ( .A1(n13396), .A2(n9152), .ZN(n9124) );
  AOI21_X1 U11594 ( .B1(n13625), .B2(n9214), .A(n9124), .ZN(n9128) );
  NAND2_X1 U11595 ( .A1(n13625), .A2(n9213), .ZN(n9126) );
  NAND2_X1 U11596 ( .A1(n13396), .A2(n9168), .ZN(n9125) );
  NAND2_X1 U11597 ( .A1(n9126), .A2(n9125), .ZN(n9127) );
  NAND2_X1 U11598 ( .A1(n9129), .A2(n9128), .ZN(n9130) );
  NAND2_X1 U11599 ( .A1(n13603), .A2(n9017), .ZN(n9133) );
  NAND2_X1 U11600 ( .A1(n13577), .A2(n9168), .ZN(n9132) );
  NAND2_X1 U11601 ( .A1(n9133), .A2(n9132), .ZN(n9135) );
  AOI22_X1 U11602 ( .A1(n13603), .A2(n9168), .B1(n13577), .B2(n9213), .ZN(
        n9134) );
  NAND2_X1 U11603 ( .A1(n13710), .A2(n9168), .ZN(n9137) );
  NAND2_X1 U11604 ( .A1(n13401), .A2(n9017), .ZN(n9136) );
  NAND2_X1 U11605 ( .A1(n9137), .A2(n9136), .ZN(n9139) );
  AOI22_X1 U11606 ( .A1(n13710), .A2(n9152), .B1(n9214), .B2(n13401), .ZN(
        n9138) );
  NAND2_X1 U11607 ( .A1(n13568), .A2(n6473), .ZN(n9141) );
  NAND2_X1 U11608 ( .A1(n13579), .A2(n9168), .ZN(n9140) );
  NAND2_X1 U11609 ( .A1(n9141), .A2(n9140), .ZN(n9144) );
  AOI22_X1 U11610 ( .A1(n13568), .A2(n9168), .B1(n13579), .B2(n6473), .ZN(
        n9142) );
  NAND2_X1 U11611 ( .A1(n13548), .A2(n9214), .ZN(n9146) );
  NAND2_X1 U11612 ( .A1(n13406), .A2(n9017), .ZN(n9145) );
  NAND2_X1 U11613 ( .A1(n9146), .A2(n9145), .ZN(n9149) );
  AOI22_X1 U11614 ( .A1(n13548), .A2(n9017), .B1(n9214), .B2(n13406), .ZN(
        n9147) );
  OAI22_X1 U11615 ( .A1(n13536), .A2(n9214), .B1(n13555), .B2(n9213), .ZN(
        n9151) );
  AOI22_X1 U11616 ( .A1(n13695), .A2(n9168), .B1(n13520), .B2(n6473), .ZN(
        n9150) );
  AOI22_X1 U11617 ( .A1(n13688), .A2(n9168), .B1(n13412), .B2(n6473), .ZN(
        n9154) );
  AOI22_X1 U11618 ( .A1(n13688), .A2(n9152), .B1(n9214), .B2(n13412), .ZN(
        n9153) );
  OAI22_X1 U11619 ( .A1(n13512), .A2(n9214), .B1(n13485), .B2(n9213), .ZN(
        n9157) );
  INV_X1 U11620 ( .A(n9157), .ZN(n9160) );
  AOI22_X1 U11621 ( .A1(n13684), .A2(n9168), .B1(n6840), .B2(n6473), .ZN(n9158) );
  INV_X1 U11622 ( .A(n9164), .ZN(n9167) );
  AOI22_X1 U11623 ( .A1(n13495), .A2(n9168), .B1(n13438), .B2(n6473), .ZN(
        n9163) );
  INV_X1 U11624 ( .A(n9163), .ZN(n9166) );
  AOI22_X1 U11625 ( .A1(n13495), .A2(n6473), .B1(n9214), .B2(n13438), .ZN(
        n9161) );
  OAI21_X1 U11626 ( .B1(n9167), .B2(n9166), .A(n9165), .ZN(n9171) );
  OAI22_X1 U11627 ( .A1(n13416), .A2(n9214), .B1(n13484), .B2(n9017), .ZN(
        n9170) );
  AOI22_X1 U11628 ( .A1(n13668), .A2(n9168), .B1(n13296), .B2(n6473), .ZN(
        n9179) );
  OAI22_X1 U11629 ( .A1(n7097), .A2(n9214), .B1(n13444), .B2(n6473), .ZN(n9178) );
  AOI22_X1 U11630 ( .A1(n7100), .A2(n9168), .B1(n13297), .B2(n6473), .ZN(n9169) );
  INV_X1 U11631 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14455) );
  MUX2_X1 U11632 ( .A(n14455), .B(n12282), .S(n9945), .Z(n9186) );
  XNOR2_X1 U11633 ( .A(n9186), .B(SI_29_), .ZN(n9180) );
  NOR2_X1 U11634 ( .A1(n9207), .A2(n12282), .ZN(n9175) );
  OAI22_X1 U11635 ( .A1(n13446), .A2(n9214), .B1(n9176), .B2(n9213), .ZN(n9216) );
  AOI22_X1 U11636 ( .A1(n13659), .A2(n9214), .B1(n13295), .B2(n6473), .ZN(
        n9217) );
  AOI22_X1 U11637 ( .A1(n9216), .A2(n9217), .B1(n9179), .B2(n9178), .ZN(n9200)
         );
  MUX2_X1 U11638 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9945), .Z(n9183) );
  INV_X1 U11639 ( .A(SI_31_), .ZN(n9182) );
  XNOR2_X1 U11640 ( .A(n9183), .B(n9182), .ZN(n9188) );
  INV_X1 U11641 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12482) );
  INV_X1 U11642 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12290) );
  MUX2_X1 U11643 ( .A(n12482), .B(n12290), .S(n9945), .Z(n9185) );
  INV_X1 U11644 ( .A(n9185), .ZN(n9184) );
  NAND2_X1 U11645 ( .A1(n9184), .A2(SI_30_), .ZN(n9204) );
  NAND2_X1 U11646 ( .A1(n9188), .A2(n9204), .ZN(n9194) );
  INV_X1 U11647 ( .A(SI_30_), .ZN(n12292) );
  NAND2_X1 U11648 ( .A1(n9185), .A2(n12292), .ZN(n9203) );
  INV_X1 U11649 ( .A(SI_29_), .ZN(n13177) );
  NAND2_X1 U11650 ( .A1(n9186), .A2(n13177), .ZN(n9201) );
  NAND2_X1 U11651 ( .A1(n9203), .A2(n9201), .ZN(n9190) );
  NOR2_X1 U11652 ( .A1(n9190), .A2(n9188), .ZN(n9187) );
  NAND2_X1 U11653 ( .A1(n9202), .A2(n9187), .ZN(n9193) );
  INV_X1 U11654 ( .A(n9188), .ZN(n9191) );
  XNOR2_X1 U11655 ( .A(n9188), .B(n9204), .ZN(n9189) );
  OAI21_X1 U11656 ( .B1(n9191), .B2(n9190), .A(n9189), .ZN(n9192) );
  NAND2_X1 U11657 ( .A1(n13785), .A2(n9209), .ZN(n9197) );
  INV_X1 U11658 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9195) );
  OR2_X1 U11659 ( .A1(n9207), .A2(n9195), .ZN(n9196) );
  INV_X1 U11660 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13652) );
  NAND2_X1 U11661 ( .A1(n7701), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9199) );
  NAND2_X1 U11662 ( .A1(n7702), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9198) );
  OAI211_X1 U11663 ( .C1(n7736), .C2(n13652), .A(n9199), .B(n9198), .ZN(n13384) );
  XNOR2_X1 U11664 ( .A(n13380), .B(n13384), .ZN(n9220) );
  AND2_X1 U11665 ( .A1(n9204), .A2(n9203), .ZN(n9205) );
  NOR2_X1 U11666 ( .A1(n9207), .A2(n12290), .ZN(n9208) );
  AOI222_X1 U11667 ( .A1(n9210), .A2(P2_REG1_REG_30__SCAN_IN), .B1(n7702), 
        .B2(P2_REG0_REG_30__SCAN_IN), .C1(n7701), .C2(P2_REG2_REG_30__SCAN_IN), 
        .ZN(n13441) );
  AND2_X1 U11668 ( .A1(n13384), .A2(n9017), .ZN(n9225) );
  NOR2_X1 U11669 ( .A1(n10637), .A2(n9923), .ZN(n9262) );
  NOR4_X1 U11670 ( .A1(n9225), .A2(n9262), .A3(n9211), .A4(n11983), .ZN(n9212)
         );
  OAI22_X1 U11671 ( .A1(n13754), .A2(n9152), .B1(n13441), .B2(n9212), .ZN(
        n9223) );
  INV_X1 U11672 ( .A(n13754), .ZN(n9215) );
  INV_X1 U11673 ( .A(n13441), .ZN(n13294) );
  AOI22_X1 U11674 ( .A1(n9215), .A2(n9213), .B1(n9214), .B2(n13294), .ZN(n9222) );
  INV_X1 U11675 ( .A(n9216), .ZN(n9219) );
  INV_X1 U11676 ( .A(n9217), .ZN(n9218) );
  AOI22_X1 U11677 ( .A1(n9223), .A2(n9222), .B1(n9219), .B2(n9218), .ZN(n9221)
         );
  INV_X1 U11678 ( .A(n9220), .ZN(n9253) );
  NAND2_X1 U11679 ( .A1(n13384), .A2(n9214), .ZN(n9228) );
  INV_X1 U11680 ( .A(n9225), .ZN(n9226) );
  NAND2_X1 U11681 ( .A1(n9226), .A2(n9017), .ZN(n9227) );
  MUX2_X1 U11682 ( .A(n9228), .B(n9227), .S(n13380), .Z(n9229) );
  NAND2_X1 U11683 ( .A1(n13668), .A2(n13296), .ZN(n13417) );
  XNOR2_X1 U11684 ( .A(n13568), .B(n13579), .ZN(n13564) );
  INV_X1 U11685 ( .A(n13396), .ZN(n13595) );
  XNOR2_X1 U11686 ( .A(n13625), .B(n13595), .ZN(n13614) );
  XNOR2_X1 U11687 ( .A(n13727), .B(n13423), .ZN(n13642) );
  INV_X1 U11688 ( .A(n13391), .ZN(n13418) );
  XNOR2_X1 U11689 ( .A(n13419), .B(n13418), .ZN(n12212) );
  INV_X1 U11690 ( .A(n13298), .ZN(n9232) );
  OR2_X1 U11691 ( .A1(n13782), .A2(n9232), .ZN(n12210) );
  NAND2_X1 U11692 ( .A1(n13782), .A2(n9232), .ZN(n9233) );
  NAND2_X1 U11693 ( .A1(n12210), .A2(n9233), .ZN(n12200) );
  XNOR2_X1 U11694 ( .A(n13744), .B(n13299), .ZN(n12011) );
  INV_X1 U11695 ( .A(n13301), .ZN(n9234) );
  OR2_X1 U11696 ( .A1(n13221), .A2(n9234), .ZN(n11905) );
  NAND2_X1 U11697 ( .A1(n13221), .A2(n9234), .ZN(n9235) );
  NAND2_X1 U11698 ( .A1(n11905), .A2(n9235), .ZN(n11903) );
  XNOR2_X1 U11699 ( .A(n11816), .B(n11815), .ZN(n11668) );
  XNOR2_X1 U11700 ( .A(n11663), .B(n13303), .ZN(n11660) );
  XNOR2_X1 U11701 ( .A(n11437), .B(n11401), .ZN(n11249) );
  XNOR2_X1 U11702 ( .A(n14954), .B(n13306), .ZN(n11159) );
  NAND2_X1 U11703 ( .A1(n13311), .A2(n14978), .ZN(n9238) );
  INV_X1 U11704 ( .A(n10323), .ZN(n10428) );
  NAND2_X1 U11705 ( .A1(n10428), .A2(n10421), .ZN(n9921) );
  NAND2_X1 U11706 ( .A1(n8994), .A2(n10323), .ZN(n9239) );
  NAND2_X1 U11707 ( .A1(n9921), .A2(n9239), .ZN(n14976) );
  INV_X1 U11708 ( .A(n13309), .ZN(n10965) );
  NOR2_X1 U11709 ( .A1(n9240), .A2(n10964), .ZN(n9241) );
  XNOR2_X1 U11710 ( .A(n14991), .B(n13307), .ZN(n11149) );
  XNOR2_X1 U11711 ( .A(n11071), .B(n13308), .ZN(n10967) );
  NAND4_X1 U11712 ( .A1(n11159), .A2(n9241), .A3(n11149), .A4(n10967), .ZN(
        n9242) );
  NOR2_X1 U11713 ( .A1(n11249), .A2(n9242), .ZN(n9243) );
  XNOR2_X1 U11714 ( .A(n11554), .B(n13304), .ZN(n11513) );
  NAND3_X1 U11715 ( .A1(n11660), .A2(n9243), .A3(n11513), .ZN(n9244) );
  NOR3_X1 U11716 ( .A1(n11903), .A2(n11668), .A3(n9244), .ZN(n9245) );
  XNOR2_X1 U11717 ( .A(n14868), .B(n13300), .ZN(n11907) );
  NAND3_X1 U11718 ( .A1(n12011), .A2(n9245), .A3(n11907), .ZN(n9246) );
  OR4_X1 U11719 ( .A1(n13642), .A2(n12212), .A3(n12200), .A4(n9246), .ZN(n9247) );
  NOR2_X1 U11720 ( .A1(n13614), .A2(n9247), .ZN(n9248) );
  XNOR2_X1 U11721 ( .A(n13710), .B(n13401), .ZN(n13586) );
  OR2_X1 U11722 ( .A1(n13603), .A2(n13577), .ZN(n13398) );
  NAND2_X1 U11723 ( .A1(n13603), .A2(n13577), .ZN(n13397) );
  NAND2_X1 U11724 ( .A1(n13398), .A2(n13397), .ZN(n13592) );
  NAND4_X1 U11725 ( .A1(n13564), .A2(n9248), .A3(n13586), .A4(n13592), .ZN(
        n9249) );
  XNOR2_X1 U11726 ( .A(n13548), .B(n13563), .ZN(n13431) );
  NOR2_X1 U11727 ( .A1(n9249), .A2(n13431), .ZN(n9250) );
  XNOR2_X1 U11728 ( .A(n13695), .B(n13520), .ZN(n13538) );
  XNOR2_X1 U11729 ( .A(n13495), .B(n13438), .ZN(n13489) );
  NAND4_X1 U11730 ( .A1(n13454), .A2(n9250), .A3(n13538), .A4(n13489), .ZN(
        n9252) );
  XNOR2_X1 U11731 ( .A(n7100), .B(n13297), .ZN(n13468) );
  NAND2_X1 U11732 ( .A1(n13468), .A2(n13517), .ZN(n9251) );
  XNOR2_X1 U11733 ( .A(n13659), .B(n13295), .ZN(n13439) );
  XNOR2_X1 U11734 ( .A(n13754), .B(n13441), .ZN(n9254) );
  NAND3_X1 U11735 ( .A1(n9255), .A2(n13439), .A3(n9254), .ZN(n9256) );
  NAND2_X1 U11736 ( .A1(n8221), .A2(n12284), .ZN(n9258) );
  OAI211_X1 U11737 ( .C1(n9259), .C2(n10616), .A(n9267), .B(n9258), .ZN(n9260)
         );
  NAND2_X1 U11738 ( .A1(n6864), .A2(n9924), .ZN(n9264) );
  INV_X1 U11739 ( .A(n9262), .ZN(n9263) );
  OAI21_X1 U11740 ( .B1(n9264), .B2(n11983), .A(n9263), .ZN(n9265) );
  NOR2_X1 U11741 ( .A1(n10068), .A2(P2_U3088), .ZN(n9268) );
  NOR4_X1 U11742 ( .A1(n14970), .A2(n13796), .A3(n9267), .A4(n13594), .ZN(
        n9270) );
  INV_X1 U11743 ( .A(n9268), .ZN(n12249) );
  OAI21_X1 U11744 ( .B1(n12249), .B2(n10616), .A(P2_B_REG_SCAN_IN), .ZN(n9269)
         );
  OAI21_X1 U11745 ( .B1(n9274), .B2(n9273), .A(n9272), .ZN(n9275) );
  NAND2_X1 U11746 ( .A1(n9275), .A2(n12468), .ZN(n9282) );
  INV_X1 U11747 ( .A(n12897), .ZN(n9277) );
  AOI22_X1 U11748 ( .A1(n12921), .A2(n12470), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9276) );
  OAI21_X1 U11749 ( .B1(n9277), .B2(n12034), .A(n9276), .ZN(n9278) );
  AOI21_X1 U11750 ( .B1(n12889), .B2(n12439), .A(n9278), .ZN(n9279) );
  INV_X1 U11751 ( .A(n9280), .ZN(n9281) );
  NAND2_X1 U11752 ( .A1(n9282), .A2(n9281), .ZN(P3_U3154) );
  NAND2_X1 U11753 ( .A1(n9424), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9459) );
  NAND2_X1 U11754 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n9283) );
  NOR2_X1 U11755 ( .A1(n9459), .A2(n9283), .ZN(n9476) );
  NAND2_X1 U11756 ( .A1(n9476), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9508) );
  INV_X1 U11757 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10296) );
  INV_X1 U11758 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n12050) );
  NAND2_X1 U11759 ( .A1(n9591), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9592) );
  INV_X1 U11760 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9284) );
  NAND2_X1 U11761 ( .A1(n9592), .A2(n9284), .ZN(n9285) );
  NAND2_X1 U11762 ( .A1(n9614), .A2(n9285), .ZN(n14724) );
  INV_X1 U11763 ( .A(n14724), .ZN(n9297) );
  INV_X1 U11764 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9292) );
  XNOR2_X2 U11765 ( .A(n9294), .B(n9293), .ZN(n12265) );
  NAND2_X1 U11766 ( .A1(n9297), .A2(n9331), .ZN(n9303) );
  NAND2_X1 U11767 ( .A1(n9386), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9302) );
  INV_X1 U11768 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14295) );
  OR2_X1 U11769 ( .A1(n6475), .A2(n14295), .ZN(n9301) );
  NAND2_X1 U11770 ( .A1(n9791), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9300) );
  NAND4_X1 U11771 ( .A1(n9303), .A2(n9302), .A3(n9301), .A4(n9300), .ZN(n14028) );
  NAND2_X1 U11772 ( .A1(n11170), .A2(n9825), .ZN(n9310) );
  NAND2_X1 U11773 ( .A1(n9431), .A2(n9305), .ZN(n9325) );
  NAND2_X1 U11774 ( .A1(n9325), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9307) );
  XNOR2_X1 U11775 ( .A(n9307), .B(n9306), .ZN(n14079) );
  OAI22_X1 U11776 ( .A1(n9633), .A2(n11171), .B1(n6853), .B2(n14079), .ZN(
        n9308) );
  INV_X1 U11777 ( .A(n9308), .ZN(n9309) );
  INV_X1 U11778 ( .A(n9311), .ZN(n9327) );
  NAND2_X1 U11779 ( .A1(n9327), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9312) );
  XNOR2_X1 U11780 ( .A(n9312), .B(P1_IR_REG_20__SCAN_IN), .ZN(n9833) );
  NAND2_X1 U11781 ( .A1(n9316), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9315) );
  MUX2_X1 U11782 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9317), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n9321) );
  NAND2_X1 U11783 ( .A1(n9321), .A2(n9891), .ZN(n9829) );
  INV_X1 U11784 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9322) );
  AND3_X1 U11785 ( .A1(n9323), .A2(n9322), .A3(P1_IR_REG_19__SCAN_IN), .ZN(
        n9329) );
  INV_X1 U11786 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9324) );
  XNOR2_X1 U11787 ( .A(n9324), .B(P1_IR_REG_31__SCAN_IN), .ZN(n9328) );
  NOR2_X2 U11788 ( .A1(n9330), .A2(n10599), .ZN(n9399) );
  INV_X1 U11789 ( .A(n9399), .ZN(n9492) );
  MUX2_X1 U11790 ( .A(n14028), .B(n14721), .S(n9821), .Z(n9606) );
  INV_X1 U11791 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10173) );
  INV_X1 U11792 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9332) );
  OR2_X1 U11793 ( .A1(n9387), .A2(n9332), .ZN(n9334) );
  NAND2_X1 U11794 ( .A1(n9409), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9333) );
  NAND2_X1 U11795 ( .A1(n9338), .A2(n9942), .ZN(n9344) );
  OR2_X1 U11796 ( .A1(n9340), .A2(n9292), .ZN(n9341) );
  XNOR2_X1 U11797 ( .A(n9341), .B(P1_IR_REG_2__SCAN_IN), .ZN(n10750) );
  NAND2_X1 U11798 ( .A1(n9627), .A2(n10750), .ZN(n9342) );
  INV_X1 U11799 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11349) );
  INV_X1 U11800 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9345) );
  OR2_X1 U11801 ( .A1(n9387), .A2(n9345), .ZN(n9347) );
  NAND2_X1 U11802 ( .A1(n9409), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9346) );
  INV_X1 U11803 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9349) );
  INV_X1 U11804 ( .A(SI_0_), .ZN(n9999) );
  OAI21_X1 U11805 ( .B1(n9945), .B2(n9999), .A(n9350), .ZN(n9351) );
  AND2_X1 U11806 ( .A1(n9352), .A2(n9351), .ZN(n14477) );
  MUX2_X1 U11807 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14477), .S(n9339), .Z(n11045)
         );
  NAND2_X1 U11808 ( .A1(n14041), .A2(n11351), .ZN(n9857) );
  NAND2_X1 U11809 ( .A1(n9857), .A2(n10599), .ZN(n9363) );
  NAND2_X1 U11810 ( .A1(n9409), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9358) );
  INV_X1 U11811 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9353) );
  INV_X1 U11812 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9355) );
  OR2_X1 U11813 ( .A1(n9387), .A2(n9355), .ZN(n9356) );
  INV_X1 U11814 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10153) );
  NAND2_X1 U11815 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9361) );
  XNOR2_X1 U11816 ( .A(n9361), .B(P1_IR_REG_1__SCAN_IN), .ZN(n10189) );
  NAND3_X1 U11817 ( .A1(n9363), .A2(n10850), .A3(n10849), .ZN(n9364) );
  NAND2_X1 U11818 ( .A1(n9364), .A2(n7555), .ZN(n9367) );
  OAI211_X1 U11819 ( .C1(n10849), .C2(n9365), .A(n9399), .B(n10850), .ZN(n9366) );
  NAND2_X1 U11820 ( .A1(n9367), .A2(n9366), .ZN(n9368) );
  OAI21_X1 U11821 ( .B1(n9370), .B2(n9369), .A(n9368), .ZN(n9372) );
  NAND2_X1 U11822 ( .A1(n9372), .A2(n9371), .ZN(n9382) );
  OR2_X1 U11823 ( .A1(n9354), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9376) );
  NAND2_X1 U11824 ( .A1(n9386), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9375) );
  NAND2_X1 U11825 ( .A1(n9791), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9374) );
  INV_X1 U11826 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n14305) );
  OR2_X1 U11827 ( .A1(n9812), .A2(n14305), .ZN(n9373) );
  NAND4_X1 U11828 ( .A1(n9376), .A2(n9375), .A3(n9374), .A4(n9373), .ZN(n14037) );
  NAND2_X1 U11829 ( .A1(n9338), .A2(n9948), .ZN(n9381) );
  NAND2_X1 U11830 ( .A1(n9377), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9378) );
  MUX2_X1 U11831 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9378), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9379) );
  AND2_X1 U11832 ( .A1(n9393), .A2(n9379), .ZN(n14052) );
  NAND2_X1 U11833 ( .A1(n9627), .A2(n14052), .ZN(n9380) );
  OAI211_X1 U11834 ( .C1(n9633), .C2(n9950), .A(n9381), .B(n9380), .ZN(n11119)
         );
  XNOR2_X1 U11835 ( .A(n14037), .B(n11119), .ZN(n10989) );
  NAND2_X1 U11836 ( .A1(n9382), .A2(n10989), .ZN(n9385) );
  INV_X1 U11837 ( .A(n14037), .ZN(n11200) );
  MUX2_X1 U11838 ( .A(n11200), .B(n14306), .S(n9399), .Z(n9383) );
  NAND2_X1 U11839 ( .A1(n11200), .A2(n14306), .ZN(n11117) );
  NAND2_X1 U11840 ( .A1(n9383), .A2(n11117), .ZN(n9384) );
  NAND2_X1 U11841 ( .A1(n9385), .A2(n9384), .ZN(n9402) );
  NAND2_X1 U11842 ( .A1(n9386), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9392) );
  INV_X1 U11843 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9388) );
  OR2_X1 U11844 ( .A1(n9387), .A2(n9388), .ZN(n9391) );
  XNOR2_X1 U11845 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n11197) );
  OR2_X1 U11846 ( .A1(n9354), .A2(n11197), .ZN(n9390) );
  INV_X1 U11847 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10178) );
  OR2_X1 U11848 ( .A1(n9812), .A2(n10178), .ZN(n9389) );
  NAND2_X1 U11849 ( .A1(n9953), .A2(n9338), .ZN(n9398) );
  NAND2_X1 U11850 ( .A1(n9393), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9395) );
  INV_X1 U11851 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9394) );
  XNOR2_X1 U11852 ( .A(n9395), .B(n9394), .ZN(n10786) );
  OAI22_X1 U11853 ( .A1(n9633), .A2(n9954), .B1(n9339), .B2(n10786), .ZN(n9396) );
  INV_X1 U11854 ( .A(n9396), .ZN(n9397) );
  AND2_X2 U11855 ( .A1(n9398), .A2(n9397), .ZN(n11193) );
  MUX2_X1 U11856 ( .A(n11194), .B(n11193), .S(n9399), .Z(n9401) );
  INV_X2 U11857 ( .A(n11194), .ZN(n14036) );
  MUX2_X1 U11858 ( .A(n14809), .B(n14036), .S(n9830), .Z(n9400) );
  OAI21_X1 U11859 ( .B1(n9402), .B2(n9401), .A(n9400), .ZN(n9404) );
  NAND2_X1 U11860 ( .A1(n9402), .A2(n9401), .ZN(n9403) );
  NAND2_X1 U11861 ( .A1(n9404), .A2(n9403), .ZN(n9418) );
  NAND2_X1 U11862 ( .A1(n9951), .A2(n9338), .ZN(n9408) );
  OR2_X1 U11863 ( .A1(n9431), .A2(n9292), .ZN(n9405) );
  XNOR2_X1 U11864 ( .A(n9405), .B(n9430), .ZN(n10198) );
  OAI22_X1 U11865 ( .A1(n9633), .A2(n9952), .B1(n9339), .B2(n10198), .ZN(n9406) );
  INV_X1 U11866 ( .A(n9406), .ZN(n9407) );
  NAND2_X1 U11867 ( .A1(n9408), .A2(n9407), .ZN(n14813) );
  NAND2_X1 U11868 ( .A1(n9386), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9415) );
  AOI21_X1 U11869 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9410) );
  NOR2_X1 U11870 ( .A1(n9410), .A2(n9424), .ZN(n11440) );
  NAND2_X1 U11871 ( .A1(n9331), .A2(n11440), .ZN(n9414) );
  INV_X1 U11872 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9411) );
  OR2_X1 U11873 ( .A1(n9814), .A2(n9411), .ZN(n9413) );
  INV_X1 U11874 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11137) );
  OR2_X1 U11875 ( .A1(n6475), .A2(n11137), .ZN(n9412) );
  NAND4_X1 U11876 ( .A1(n9415), .A2(n9414), .A3(n9413), .A4(n9412), .ZN(n14035) );
  MUX2_X1 U11877 ( .A(n14813), .B(n14035), .S(n9802), .Z(n9419) );
  NAND2_X1 U11878 ( .A1(n9418), .A2(n9419), .ZN(n9417) );
  MUX2_X1 U11879 ( .A(n14035), .B(n14813), .S(n9802), .Z(n9416) );
  NAND2_X1 U11880 ( .A1(n9417), .A2(n9416), .ZN(n9423) );
  INV_X1 U11881 ( .A(n9418), .ZN(n9421) );
  INV_X1 U11882 ( .A(n9419), .ZN(n9420) );
  NAND2_X1 U11883 ( .A1(n9421), .A2(n9420), .ZN(n9422) );
  NAND2_X1 U11884 ( .A1(n9423), .A2(n9422), .ZN(n9439) );
  INV_X2 U11885 ( .A(n9331), .ZN(n9709) );
  OAI21_X1 U11886 ( .B1(n9424), .B2(P1_REG3_REG_6__SCAN_IN), .A(n9459), .ZN(
        n11610) );
  OR2_X1 U11887 ( .A1(n9709), .A2(n11610), .ZN(n9429) );
  NAND2_X1 U11888 ( .A1(n9791), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9428) );
  NAND2_X1 U11889 ( .A1(n9386), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9427) );
  INV_X1 U11890 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9425) );
  OR2_X1 U11891 ( .A1(n6475), .A2(n9425), .ZN(n9426) );
  NAND2_X1 U11892 ( .A1(n9964), .A2(n9825), .ZN(n9436) );
  NAND2_X1 U11893 ( .A1(n9431), .A2(n9430), .ZN(n9450) );
  NAND2_X1 U11894 ( .A1(n9450), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9433) );
  XNOR2_X1 U11895 ( .A(n9433), .B(n9432), .ZN(n14057) );
  OAI22_X1 U11896 ( .A1(n9633), .A2(n9965), .B1(n6853), .B2(n14057), .ZN(n9434) );
  INV_X1 U11897 ( .A(n9434), .ZN(n9435) );
  NAND2_X1 U11898 ( .A1(n9436), .A2(n9435), .ZN(n11617) );
  INV_X2 U11899 ( .A(n9492), .ZN(n9830) );
  MUX2_X1 U11900 ( .A(n14034), .B(n11617), .S(n9830), .Z(n9440) );
  NAND2_X1 U11901 ( .A1(n9439), .A2(n9440), .ZN(n9438) );
  MUX2_X1 U11902 ( .A(n14034), .B(n11617), .S(n9821), .Z(n9437) );
  NAND2_X1 U11903 ( .A1(n9438), .A2(n9437), .ZN(n9444) );
  INV_X1 U11904 ( .A(n9439), .ZN(n9442) );
  INV_X1 U11905 ( .A(n9440), .ZN(n9441) );
  NAND2_X1 U11906 ( .A1(n9442), .A2(n9441), .ZN(n9443) );
  NAND2_X1 U11907 ( .A1(n9386), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9449) );
  XNOR2_X1 U11908 ( .A(n9459), .B(P1_REG3_REG_7__SCAN_IN), .ZN(n11535) );
  NAND2_X1 U11909 ( .A1(n9331), .A2(n11535), .ZN(n9448) );
  INV_X1 U11910 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9445) );
  OR2_X1 U11911 ( .A1(n9814), .A2(n9445), .ZN(n9447) );
  INV_X1 U11912 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10179) );
  OR2_X1 U11913 ( .A1(n6475), .A2(n10179), .ZN(n9446) );
  NAND4_X1 U11914 ( .A1(n9449), .A2(n9448), .A3(n9447), .A4(n9446), .ZN(n14033) );
  NAND2_X1 U11915 ( .A1(n9969), .A2(n9825), .ZN(n9455) );
  NAND2_X1 U11916 ( .A1(n9466), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9452) );
  XNOR2_X1 U11917 ( .A(n9452), .B(n9451), .ZN(n10220) );
  OAI22_X1 U11918 ( .A1(n9633), .A2(n9972), .B1(n6853), .B2(n10220), .ZN(n9453) );
  INV_X1 U11919 ( .A(n9453), .ZN(n9454) );
  MUX2_X1 U11920 ( .A(n14033), .B(n11536), .S(n9821), .Z(n9458) );
  MUX2_X1 U11921 ( .A(n14033), .B(n11536), .S(n9830), .Z(n9456) );
  INV_X1 U11922 ( .A(n9459), .ZN(n9460) );
  AOI21_X1 U11923 ( .B1(n9460), .B2(P1_REG3_REG_7__SCAN_IN), .A(
        P1_REG3_REG_8__SCAN_IN), .ZN(n9461) );
  OR2_X1 U11924 ( .A1(n9461), .A2(n9476), .ZN(n15203) );
  OR2_X1 U11925 ( .A1(n9709), .A2(n15203), .ZN(n9465) );
  NAND2_X1 U11926 ( .A1(n9791), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9464) );
  NAND2_X1 U11927 ( .A1(n9386), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9463) );
  INV_X1 U11928 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11383) );
  OR2_X1 U11929 ( .A1(n6475), .A2(n11383), .ZN(n9462) );
  NAND4_X1 U11930 ( .A1(n9465), .A2(n9464), .A3(n9463), .A4(n9462), .ZN(n14032) );
  NAND2_X1 U11931 ( .A1(n10000), .A2(n9825), .ZN(n9470) );
  NAND2_X1 U11932 ( .A1(n9587), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9467) );
  XNOR2_X1 U11933 ( .A(n9467), .B(n9482), .ZN(n10281) );
  OAI22_X1 U11934 ( .A1(n9633), .A2(n10003), .B1(n6853), .B2(n10281), .ZN(
        n9468) );
  INV_X1 U11935 ( .A(n9468), .ZN(n9469) );
  MUX2_X1 U11936 ( .A(n14032), .B(n15198), .S(n9830), .Z(n9473) );
  MUX2_X1 U11937 ( .A(n14032), .B(n15198), .S(n9821), .Z(n9471) );
  NAND2_X1 U11938 ( .A1(n9472), .A2(n9471), .ZN(n9475) );
  OR2_X1 U11939 ( .A1(n9476), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9477) );
  NAND2_X1 U11940 ( .A1(n9508), .A2(n9477), .ZN(n11789) );
  OR2_X1 U11941 ( .A1(n9709), .A2(n11789), .ZN(n9481) );
  NAND2_X1 U11942 ( .A1(n9791), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9480) );
  NAND2_X1 U11943 ( .A1(n9386), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9479) );
  INV_X1 U11944 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11601) );
  OR2_X1 U11945 ( .A1(n6475), .A2(n11601), .ZN(n9478) );
  NAND4_X1 U11946 ( .A1(n9481), .A2(n9480), .A3(n9479), .A4(n9478), .ZN(n14031) );
  NAND2_X1 U11947 ( .A1(n10056), .A2(n9825), .ZN(n9491) );
  INV_X1 U11948 ( .A(n9587), .ZN(n9483) );
  NAND2_X1 U11949 ( .A1(n9483), .A2(n9482), .ZN(n9485) );
  NAND2_X1 U11950 ( .A1(n9485), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9484) );
  MUX2_X1 U11951 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9484), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n9488) );
  INV_X1 U11952 ( .A(n9485), .ZN(n9487) );
  INV_X1 U11953 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9486) );
  NAND2_X1 U11954 ( .A1(n9487), .A2(n9486), .ZN(n9502) );
  NAND2_X1 U11955 ( .A1(n9488), .A2(n9502), .ZN(n10300) );
  OAI22_X1 U11956 ( .A1(n9633), .A2(n10057), .B1(n10300), .B2(n6853), .ZN(
        n9489) );
  INV_X1 U11957 ( .A(n9489), .ZN(n9490) );
  MUX2_X1 U11958 ( .A(n14031), .B(n11767), .S(n9821), .Z(n9496) );
  NAND2_X1 U11959 ( .A1(n9495), .A2(n9496), .ZN(n9494) );
  MUX2_X1 U11960 ( .A(n14031), .B(n11767), .S(n9830), .Z(n9493) );
  NAND2_X1 U11961 ( .A1(n9494), .A2(n9493), .ZN(n9500) );
  INV_X1 U11962 ( .A(n9495), .ZN(n9498) );
  INV_X1 U11963 ( .A(n9496), .ZN(n9497) );
  NAND2_X1 U11964 ( .A1(n9498), .A2(n9497), .ZN(n9499) );
  NAND2_X1 U11965 ( .A1(n9500), .A2(n9499), .ZN(n9517) );
  NAND2_X1 U11966 ( .A1(n10221), .A2(n9825), .ZN(n9506) );
  NAND2_X1 U11967 ( .A1(n9502), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9501) );
  MUX2_X1 U11968 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9501), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n9503) );
  NAND2_X1 U11969 ( .A1(n9503), .A2(n9544), .ZN(n10303) );
  OAI22_X1 U11970 ( .A1(n10303), .A2(n6853), .B1(n9633), .B2(n10224), .ZN(
        n9504) );
  INV_X1 U11971 ( .A(n9504), .ZN(n9505) );
  NAND2_X1 U11972 ( .A1(n9506), .A2(n9505), .ZN(n11853) );
  NAND2_X1 U11973 ( .A1(n9508), .A2(n9507), .ZN(n9509) );
  NAND2_X1 U11974 ( .A1(n9523), .A2(n9509), .ZN(n11644) );
  OR2_X1 U11975 ( .A1(n9709), .A2(n11644), .ZN(n9514) );
  NAND2_X1 U11976 ( .A1(n9791), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n9513) );
  NAND2_X1 U11977 ( .A1(n9409), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9512) );
  INV_X1 U11978 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9510) );
  OR2_X1 U11979 ( .A1(n6475), .A2(n9510), .ZN(n9511) );
  NAND4_X1 U11980 ( .A1(n9514), .A2(n9513), .A3(n9512), .A4(n9511), .ZN(n14030) );
  MUX2_X1 U11981 ( .A(n11853), .B(n14030), .S(n9821), .Z(n9518) );
  NAND2_X1 U11982 ( .A1(n9517), .A2(n9518), .ZN(n9516) );
  MUX2_X1 U11983 ( .A(n11853), .B(n14030), .S(n9830), .Z(n9515) );
  NAND2_X1 U11984 ( .A1(n9516), .A2(n9515), .ZN(n9522) );
  INV_X1 U11985 ( .A(n9517), .ZN(n9520) );
  INV_X1 U11986 ( .A(n9518), .ZN(n9519) );
  NAND2_X1 U11987 ( .A1(n9520), .A2(n9519), .ZN(n9521) );
  NAND2_X1 U11988 ( .A1(n9523), .A2(n10296), .ZN(n9524) );
  NAND2_X1 U11989 ( .A1(n9536), .A2(n9524), .ZN(n11929) );
  OR2_X1 U11990 ( .A1(n9709), .A2(n11929), .ZN(n9529) );
  NAND2_X1 U11991 ( .A1(n9409), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9528) );
  NAND2_X1 U11992 ( .A1(n9790), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9527) );
  INV_X1 U11993 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9525) );
  OR2_X1 U11994 ( .A1(n9814), .A2(n9525), .ZN(n9526) );
  NAND4_X1 U11995 ( .A1(n9529), .A2(n9528), .A3(n9527), .A4(n9526), .ZN(n14029) );
  NAND2_X1 U11996 ( .A1(n10375), .A2(n9825), .ZN(n9532) );
  NAND2_X1 U11997 ( .A1(n9544), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9530) );
  XNOR2_X1 U11998 ( .A(n9530), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10450) );
  AOI22_X1 U11999 ( .A1(n10450), .A2(n9627), .B1(n9826), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n9531) );
  MUX2_X1 U12000 ( .A(n14029), .B(n12087), .S(n9821), .Z(n9534) );
  MUX2_X1 U12001 ( .A(n14029), .B(n12087), .S(n9830), .Z(n9533) );
  INV_X1 U12002 ( .A(n9534), .ZN(n9535) );
  NAND2_X1 U12003 ( .A1(n9386), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9543) );
  AND2_X1 U12004 ( .A1(n9536), .A2(n12050), .ZN(n9537) );
  NOR2_X1 U12005 ( .A1(n9556), .A2(n9537), .ZN(n14600) );
  NAND2_X1 U12006 ( .A1(n9331), .A2(n14600), .ZN(n9542) );
  INV_X1 U12007 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9538) );
  OR2_X1 U12008 ( .A1(n9814), .A2(n9538), .ZN(n9541) );
  INV_X1 U12009 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9539) );
  OR2_X1 U12010 ( .A1(n6475), .A2(n9539), .ZN(n9540) );
  NAND4_X1 U12011 ( .A1(n9543), .A2(n9542), .A3(n9541), .A4(n9540), .ZN(n14618) );
  NAND2_X1 U12012 ( .A1(n10424), .A2(n9825), .ZN(n9546) );
  OAI21_X1 U12013 ( .B1(n9544), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9563) );
  XNOR2_X1 U12014 ( .A(n9563), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10676) );
  AOI22_X1 U12015 ( .A1(n10676), .A2(n9627), .B1(n9826), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n9545) );
  MUX2_X1 U12016 ( .A(n14618), .B(n14602), .S(n9830), .Z(n9550) );
  MUX2_X1 U12017 ( .A(n14618), .B(n14602), .S(n9821), .Z(n9547) );
  NAND2_X1 U12018 ( .A1(n9548), .A2(n9547), .ZN(n9554) );
  INV_X1 U12019 ( .A(n9549), .ZN(n9552) );
  INV_X1 U12020 ( .A(n9550), .ZN(n9551) );
  NAND2_X1 U12021 ( .A1(n9552), .A2(n9551), .ZN(n9553) );
  NAND2_X1 U12022 ( .A1(n9554), .A2(n9553), .ZN(n9569) );
  NAND2_X1 U12023 ( .A1(n9386), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9561) );
  INV_X1 U12024 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9555) );
  OR2_X1 U12025 ( .A1(n9814), .A2(n9555), .ZN(n9560) );
  NOR2_X1 U12026 ( .A1(n9556), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9557) );
  OR2_X1 U12027 ( .A1(n9579), .A2(n9557), .ZN(n14612) );
  OR2_X1 U12028 ( .A1(n9709), .A2(n14612), .ZN(n9559) );
  INV_X1 U12029 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10671) );
  OR2_X1 U12030 ( .A1(n6475), .A2(n10671), .ZN(n9558) );
  NAND2_X1 U12031 ( .A1(n10612), .A2(n9825), .ZN(n9566) );
  NAND2_X1 U12032 ( .A1(n9563), .A2(n9562), .ZN(n9564) );
  NAND2_X1 U12033 ( .A1(n9564), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9574) );
  XNOR2_X1 U12034 ( .A(n9574), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10756) );
  AOI22_X1 U12035 ( .A1(n10756), .A2(n9627), .B1(n9826), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n9565) );
  MUX2_X1 U12036 ( .A(n12224), .B(n14745), .S(n9830), .Z(n9568) );
  INV_X1 U12037 ( .A(n12224), .ZN(n14704) );
  MUX2_X1 U12038 ( .A(n14704), .B(n12234), .S(n9821), .Z(n9567) );
  AOI21_X1 U12039 ( .B1(n9569), .B2(n9568), .A(n9567), .ZN(n9571) );
  NOR2_X1 U12040 ( .A1(n9569), .A2(n9568), .ZN(n9570) );
  OR2_X1 U12041 ( .A1(n10790), .A2(n9572), .ZN(n9578) );
  INV_X1 U12042 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9573) );
  NAND2_X1 U12043 ( .A1(n9574), .A2(n9573), .ZN(n9575) );
  NAND2_X1 U12044 ( .A1(n9575), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9576) );
  AOI22_X1 U12045 ( .A1(n11476), .A2(n9627), .B1(n9826), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9577) );
  NAND2_X1 U12046 ( .A1(n9409), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9585) );
  NOR2_X1 U12047 ( .A1(n9579), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9580) );
  OR2_X1 U12048 ( .A1(n9591), .A2(n9580), .ZN(n14712) );
  OR2_X1 U12049 ( .A1(n9709), .A2(n14712), .ZN(n9584) );
  INV_X1 U12050 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n12097) );
  OR2_X1 U12051 ( .A1(n6475), .A2(n12097), .ZN(n9583) );
  INV_X1 U12052 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9581) );
  OR2_X1 U12053 ( .A1(n9814), .A2(n9581), .ZN(n9582) );
  NAND2_X1 U12054 ( .A1(n13820), .A2(n12139), .ZN(n9599) );
  NAND2_X1 U12055 ( .A1(n10949), .A2(n9825), .ZN(n9590) );
  OAI21_X1 U12056 ( .B1(n9587), .B2(n9586), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9588) );
  XNOR2_X1 U12057 ( .A(n9588), .B(P1_IR_REG_15__SCAN_IN), .ZN(n14783) );
  AOI22_X1 U12058 ( .A1(n9826), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9627), 
        .B2(n14783), .ZN(n9589) );
  NAND2_X1 U12059 ( .A1(n9386), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9598) );
  OR2_X1 U12060 ( .A1(n9591), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9593) );
  AND2_X1 U12061 ( .A1(n9593), .A2(n9592), .ZN(n14019) );
  NAND2_X1 U12062 ( .A1(n9331), .A2(n14019), .ZN(n9597) );
  INV_X1 U12063 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9594) );
  OR2_X1 U12064 ( .A1(n9814), .A2(n9594), .ZN(n9596) );
  INV_X1 U12065 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n12142) );
  OR2_X1 U12066 ( .A1(n6475), .A2(n12142), .ZN(n9595) );
  NAND4_X1 U12067 ( .A1(n9598), .A2(n9597), .A3(n9596), .A4(n9595), .ZN(n14702) );
  INV_X1 U12068 ( .A(n14702), .ZN(n14713) );
  NAND2_X1 U12069 ( .A1(n13828), .A2(n14713), .ZN(n9855) );
  NAND2_X1 U12070 ( .A1(n9855), .A2(n9599), .ZN(n9601) );
  NAND2_X1 U12071 ( .A1(n12305), .A2(n12136), .ZN(n9600) );
  MUX2_X1 U12072 ( .A(n9601), .B(n9600), .S(n9821), .Z(n9602) );
  MUX2_X1 U12073 ( .A(n9855), .B(n12305), .S(n9830), .Z(n9604) );
  MUX2_X1 U12074 ( .A(n14028), .B(n14721), .S(n9830), .Z(n9605) );
  NAND2_X1 U12075 ( .A1(n11345), .A2(n9825), .ZN(n9612) );
  NAND2_X1 U12076 ( .A1(n9608), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9607) );
  MUX2_X1 U12077 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9607), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n9609) );
  OR2_X1 U12078 ( .A1(n9608), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n9625) );
  NAND2_X1 U12079 ( .A1(n9609), .A2(n9625), .ZN(n11729) );
  OAI22_X1 U12080 ( .A1(n9633), .A2(n11346), .B1(n6853), .B2(n11729), .ZN(
        n9610) );
  INV_X1 U12081 ( .A(n9610), .ZN(n9611) );
  INV_X1 U12082 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9613) );
  AND2_X1 U12083 ( .A1(n9614), .A2(n9613), .ZN(n9615) );
  OR2_X1 U12084 ( .A1(n9615), .A2(n9621), .ZN(n14738) );
  AOI22_X1 U12085 ( .A1(n9386), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n9791), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n9617) );
  INV_X1 U12086 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14278) );
  OR2_X1 U12087 ( .A1(n6475), .A2(n14278), .ZN(n9616) );
  OAI211_X1 U12088 ( .C1(n14738), .C2(n9709), .A(n9617), .B(n9616), .ZN(n14296) );
  NAND2_X1 U12089 ( .A1(n14735), .A2(n14296), .ZN(n12333) );
  NOR2_X1 U12090 ( .A1(n14735), .A2(n14296), .ZN(n12334) );
  MUX2_X1 U12091 ( .A(n14296), .B(n14735), .S(n9802), .Z(n9618) );
  INV_X1 U12092 ( .A(n9619), .ZN(n9620) );
  NOR2_X1 U12093 ( .A1(n9621), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9622) );
  OR2_X1 U12094 ( .A1(n9637), .A2(n9622), .ZN(n14264) );
  AOI22_X1 U12095 ( .A1(n9386), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9791), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n9624) );
  INV_X1 U12096 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14265) );
  OR2_X1 U12097 ( .A1(n6475), .A2(n14265), .ZN(n9623) );
  OAI211_X1 U12098 ( .C1(n14264), .C2(n9709), .A(n9624), .B(n9623), .ZN(n14027) );
  XNOR2_X1 U12099 ( .A(n14027), .B(n9830), .ZN(n9631) );
  NAND2_X1 U12100 ( .A1(n11547), .A2(n9825), .ZN(n9629) );
  NAND2_X1 U12101 ( .A1(n9625), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9626) );
  XNOR2_X1 U12102 ( .A(n9626), .B(P1_IR_REG_18__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U12103 ( .A1(n9826), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9627), 
        .B2(n11991), .ZN(n9628) );
  XNOR2_X1 U12104 ( .A(n14385), .B(n9821), .ZN(n9630) );
  OAI21_X1 U12105 ( .B1(n9632), .B2(n9631), .A(n9630), .ZN(n9645) );
  NAND2_X1 U12106 ( .A1(n9632), .A2(n9631), .ZN(n9644) );
  NAND2_X1 U12107 ( .A1(n11764), .A2(n9825), .ZN(n9636) );
  OAI22_X1 U12108 ( .A1(n9633), .A2(n11765), .B1(n14626), .B2(n6853), .ZN(
        n9634) );
  INV_X1 U12109 ( .A(n9634), .ZN(n9635) );
  OR2_X1 U12110 ( .A1(n9637), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9638) );
  AND2_X1 U12111 ( .A1(n9650), .A2(n9638), .ZN(n14249) );
  NAND2_X1 U12112 ( .A1(n14249), .A2(n9331), .ZN(n9643) );
  INV_X1 U12113 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n14439) );
  NAND2_X1 U12114 ( .A1(n9790), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9640) );
  NAND2_X1 U12115 ( .A1(n9409), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n9639) );
  OAI211_X1 U12116 ( .C1(n9814), .C2(n14439), .A(n9640), .B(n9639), .ZN(n9641)
         );
  INV_X1 U12117 ( .A(n9641), .ZN(n9642) );
  NAND2_X1 U12118 ( .A1(n9643), .A2(n9642), .ZN(n14259) );
  NAND3_X1 U12119 ( .A1(n9645), .A2(n9644), .A3(n14247), .ZN(n9649) );
  NAND2_X1 U12120 ( .A1(n14259), .A2(n9821), .ZN(n9647) );
  INV_X1 U12121 ( .A(n14259), .ZN(n12312) );
  NAND2_X1 U12122 ( .A1(n12312), .A2(n9802), .ZN(n9646) );
  MUX2_X1 U12123 ( .A(n9647), .B(n9646), .S(n14237), .Z(n9648) );
  INV_X1 U12124 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13983) );
  NAND2_X1 U12125 ( .A1(n9650), .A2(n13983), .ZN(n9652) );
  INV_X1 U12126 ( .A(n9662), .ZN(n9651) );
  NAND2_X1 U12127 ( .A1(n9652), .A2(n9651), .ZN(n13981) );
  OR2_X1 U12128 ( .A1(n13981), .A2(n9709), .ZN(n9657) );
  INV_X1 U12129 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n14376) );
  NAND2_X1 U12130 ( .A1(n9791), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9654) );
  NAND2_X1 U12131 ( .A1(n9790), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9653) );
  OAI211_X1 U12132 ( .C1(n6476), .C2(n14376), .A(n9654), .B(n9653), .ZN(n9655)
         );
  INV_X1 U12133 ( .A(n9655), .ZN(n9656) );
  NAND2_X1 U12134 ( .A1(n11900), .A2(n9825), .ZN(n9659) );
  NAND2_X1 U12135 ( .A1(n9826), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9658) );
  MUX2_X1 U12136 ( .A(n13956), .B(n14437), .S(n9821), .Z(n9661) );
  INV_X1 U12137 ( .A(n13956), .ZN(n14026) );
  MUX2_X1 U12138 ( .A(n14026), .B(n14231), .S(n9830), .Z(n9660) );
  NAND2_X1 U12139 ( .A1(n9662), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9675) );
  OAI21_X1 U12140 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n9662), .A(n9675), .ZN(
        n14215) );
  OR2_X1 U12141 ( .A1(n9709), .A2(n14215), .ZN(n9667) );
  NAND2_X1 U12142 ( .A1(n9791), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9666) );
  NAND2_X1 U12143 ( .A1(n9386), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9665) );
  INV_X1 U12144 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9663) );
  OR2_X1 U12145 ( .A1(n6475), .A2(n9663), .ZN(n9664) );
  NAND4_X1 U12146 ( .A1(n9667), .A2(n9666), .A3(n9665), .A4(n9664), .ZN(n14197) );
  NAND2_X1 U12147 ( .A1(n11980), .A2(n9825), .ZN(n9669) );
  NAND2_X1 U12148 ( .A1(n9826), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9668) );
  MUX2_X1 U12149 ( .A(n14197), .B(n14431), .S(n9802), .Z(n9672) );
  MUX2_X1 U12150 ( .A(n14197), .B(n14431), .S(n9821), .Z(n9670) );
  NAND2_X1 U12151 ( .A1(n9671), .A2(n9670), .ZN(n9674) );
  NAND2_X1 U12152 ( .A1(n9674), .A2(n9673), .ZN(n9686) );
  NAND2_X1 U12153 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n9676), .ZN(n9694) );
  OAI21_X1 U12154 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n9676), .A(n9694), .ZN(
        n13991) );
  OR2_X1 U12155 ( .A1(n9709), .A2(n13991), .ZN(n9681) );
  NAND2_X1 U12156 ( .A1(n9791), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9680) );
  NAND2_X1 U12157 ( .A1(n9409), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n9679) );
  INV_X1 U12158 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9677) );
  OR2_X1 U12159 ( .A1(n6475), .A2(n9677), .ZN(n9678) );
  NAND4_X1 U12160 ( .A1(n9681), .A2(n9680), .A3(n9679), .A4(n9678), .ZN(n14025) );
  NOR2_X1 U12161 ( .A1(n9682), .A2(n9945), .ZN(n9683) );
  XNOR2_X1 U12162 ( .A(n9683), .B(n15226), .ZN(n14476) );
  MUX2_X1 U12163 ( .A(n14025), .B(n14193), .S(n9821), .Z(n9687) );
  NAND2_X1 U12164 ( .A1(n9686), .A2(n9687), .ZN(n9685) );
  MUX2_X1 U12165 ( .A(n14025), .B(n14193), .S(n9830), .Z(n9684) );
  NAND2_X1 U12166 ( .A1(n9685), .A2(n9684), .ZN(n9691) );
  INV_X1 U12167 ( .A(n9686), .ZN(n9689) );
  INV_X1 U12168 ( .A(n9687), .ZN(n9688) );
  NAND2_X1 U12169 ( .A1(n9689), .A2(n9688), .ZN(n9690) );
  INV_X1 U12170 ( .A(n9694), .ZN(n9692) );
  NAND2_X1 U12171 ( .A1(n9692), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9707) );
  INV_X1 U12172 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9693) );
  NAND2_X1 U12173 ( .A1(n9694), .A2(n9693), .ZN(n9695) );
  NAND2_X1 U12174 ( .A1(n9707), .A2(n9695), .ZN(n14179) );
  OR2_X1 U12175 ( .A1(n9709), .A2(n14179), .ZN(n9699) );
  NAND2_X1 U12176 ( .A1(n9409), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9698) );
  NAND2_X1 U12177 ( .A1(n9790), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9697) );
  INV_X1 U12178 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n15335) );
  OR2_X1 U12179 ( .A1(n9814), .A2(n15335), .ZN(n9696) );
  NAND4_X1 U12180 ( .A1(n9699), .A2(n9698), .A3(n9697), .A4(n9696), .ZN(n14196) );
  NAND2_X1 U12181 ( .A1(n12248), .A2(n9825), .ZN(n9701) );
  NAND2_X1 U12182 ( .A1(n9826), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9700) );
  MUX2_X1 U12183 ( .A(n14196), .B(n14356), .S(n9802), .Z(n9703) );
  MUX2_X1 U12184 ( .A(n14196), .B(n14356), .S(n9821), .Z(n9702) );
  INV_X1 U12185 ( .A(n9703), .ZN(n9704) );
  INV_X1 U12186 ( .A(n9707), .ZN(n9705) );
  NAND2_X1 U12187 ( .A1(n9705), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9728) );
  INV_X1 U12188 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9706) );
  NAND2_X1 U12189 ( .A1(n9707), .A2(n9706), .ZN(n9708) );
  NAND2_X1 U12190 ( .A1(n9728), .A2(n9708), .ZN(n14167) );
  OR2_X1 U12191 ( .A1(n9709), .A2(n14167), .ZN(n9714) );
  NAND2_X1 U12192 ( .A1(n9409), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9713) );
  NAND2_X1 U12193 ( .A1(n9790), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9712) );
  INV_X1 U12194 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9710) );
  OR2_X1 U12195 ( .A1(n9814), .A2(n9710), .ZN(n9711) );
  NAND4_X1 U12196 ( .A1(n9714), .A2(n9713), .A3(n9712), .A4(n9711), .ZN(n14142) );
  NAND2_X1 U12197 ( .A1(n9826), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9716) );
  MUX2_X1 U12198 ( .A(n14142), .B(n14351), .S(n9821), .Z(n9721) );
  NAND2_X1 U12199 ( .A1(n9720), .A2(n9721), .ZN(n9719) );
  MUX2_X1 U12200 ( .A(n14142), .B(n14351), .S(n9802), .Z(n9718) );
  NAND2_X1 U12201 ( .A1(n9719), .A2(n9718), .ZN(n9725) );
  INV_X1 U12202 ( .A(n9720), .ZN(n9723) );
  INV_X1 U12203 ( .A(n9721), .ZN(n9722) );
  NAND2_X1 U12204 ( .A1(n9723), .A2(n9722), .ZN(n9724) );
  NAND2_X1 U12205 ( .A1(n9409), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9735) );
  INV_X1 U12206 ( .A(n9728), .ZN(n9726) );
  NAND2_X1 U12207 ( .A1(n9726), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9742) );
  INV_X1 U12208 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9727) );
  NAND2_X1 U12209 ( .A1(n9728), .A2(n9727), .ZN(n9729) );
  AND2_X1 U12210 ( .A1(n9742), .A2(n9729), .ZN(n14137) );
  NAND2_X1 U12211 ( .A1(n9331), .A2(n14137), .ZN(n9734) );
  INV_X1 U12212 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9730) );
  OR2_X1 U12213 ( .A1(n9814), .A2(n9730), .ZN(n9733) );
  INV_X1 U12214 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9731) );
  OR2_X1 U12215 ( .A1(n6475), .A2(n9731), .ZN(n9732) );
  NAND4_X1 U12216 ( .A1(n9735), .A2(n9734), .A3(n9733), .A4(n9732), .ZN(n14159) );
  NAND2_X1 U12217 ( .A1(n13801), .A2(n9825), .ZN(n9737) );
  NAND2_X1 U12218 ( .A1(n9826), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9736) );
  MUX2_X1 U12219 ( .A(n14159), .B(n14346), .S(n9830), .Z(n9739) );
  MUX2_X1 U12220 ( .A(n14159), .B(n14346), .S(n9821), .Z(n9738) );
  INV_X1 U12221 ( .A(n9739), .ZN(n9740) );
  NAND2_X1 U12222 ( .A1(n9409), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9748) );
  INV_X1 U12223 ( .A(n9742), .ZN(n9741) );
  NAND2_X1 U12224 ( .A1(n9741), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9761) );
  INV_X1 U12225 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14007) );
  NAND2_X1 U12226 ( .A1(n9742), .A2(n14007), .ZN(n9743) );
  AND2_X1 U12227 ( .A1(n9761), .A2(n9743), .ZN(n14131) );
  NAND2_X1 U12228 ( .A1(n9331), .A2(n14131), .ZN(n9747) );
  INV_X1 U12229 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n14422) );
  OR2_X1 U12230 ( .A1(n9814), .A2(n14422), .ZN(n9746) );
  INV_X1 U12231 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9744) );
  OR2_X1 U12232 ( .A1(n6475), .A2(n9744), .ZN(n9745) );
  NAND4_X1 U12233 ( .A1(n9748), .A2(n9747), .A3(n9746), .A4(n9745), .ZN(n14143) );
  NAND2_X1 U12234 ( .A1(n13798), .A2(n9825), .ZN(n9750) );
  NAND2_X1 U12235 ( .A1(n9826), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9749) );
  MUX2_X1 U12236 ( .A(n14143), .B(n14130), .S(n9821), .Z(n9754) );
  NAND2_X1 U12237 ( .A1(n9753), .A2(n9754), .ZN(n9752) );
  MUX2_X1 U12238 ( .A(n14143), .B(n14130), .S(n9830), .Z(n9751) );
  NAND2_X1 U12239 ( .A1(n9752), .A2(n9751), .ZN(n9758) );
  INV_X1 U12240 ( .A(n9753), .ZN(n9756) );
  INV_X1 U12241 ( .A(n9754), .ZN(n9755) );
  NAND2_X1 U12242 ( .A1(n9756), .A2(n9755), .ZN(n9757) );
  NAND2_X1 U12243 ( .A1(n9409), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9768) );
  INV_X1 U12244 ( .A(n9761), .ZN(n9759) );
  NAND2_X1 U12245 ( .A1(n9759), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9810) );
  INV_X1 U12246 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9760) );
  NAND2_X1 U12247 ( .A1(n9761), .A2(n9760), .ZN(n9762) );
  NAND2_X1 U12248 ( .A1(n9331), .A2(n14116), .ZN(n9767) );
  INV_X1 U12249 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9763) );
  OR2_X1 U12250 ( .A1(n9814), .A2(n9763), .ZN(n9766) );
  INV_X1 U12251 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9764) );
  OR2_X1 U12252 ( .A1(n6475), .A2(n9764), .ZN(n9765) );
  NAND4_X1 U12253 ( .A1(n9768), .A2(n9767), .A3(n9766), .A4(n9765), .ZN(n14024) );
  NAND2_X1 U12254 ( .A1(n13795), .A2(n9825), .ZN(n9770) );
  NAND2_X1 U12255 ( .A1(n9826), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9769) );
  MUX2_X1 U12256 ( .A(n14024), .B(n14337), .S(n9830), .Z(n9772) );
  MUX2_X1 U12257 ( .A(n14024), .B(n14337), .S(n9821), .Z(n9771) );
  INV_X1 U12258 ( .A(n9772), .ZN(n9773) );
  NAND2_X1 U12259 ( .A1(n9409), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9779) );
  XNOR2_X1 U12260 ( .A(n9810), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n13945) );
  NAND2_X1 U12261 ( .A1(n9331), .A2(n13945), .ZN(n9778) );
  INV_X1 U12262 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9774) );
  OR2_X1 U12263 ( .A1(n9814), .A2(n9774), .ZN(n9777) );
  INV_X1 U12264 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9775) );
  OR2_X1 U12265 ( .A1(n6475), .A2(n9775), .ZN(n9776) );
  NAND4_X1 U12266 ( .A1(n9779), .A2(n9778), .A3(n9777), .A4(n9776), .ZN(n14107) );
  NAND2_X1 U12267 ( .A1(n13790), .A2(n9825), .ZN(n9781) );
  NAND2_X1 U12268 ( .A1(n9826), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9780) );
  MUX2_X1 U12269 ( .A(n14107), .B(n14330), .S(n9821), .Z(n9783) );
  NAND2_X1 U12270 ( .A1(n9782), .A2(n9783), .ZN(n9787) );
  MUX2_X1 U12271 ( .A(n14330), .B(n14107), .S(n9821), .Z(n9786) );
  INV_X1 U12272 ( .A(n9782), .ZN(n9785) );
  INV_X1 U12273 ( .A(n9783), .ZN(n9784) );
  INV_X1 U12274 ( .A(n9890), .ZN(n9887) );
  NAND2_X1 U12275 ( .A1(n12264), .A2(n9825), .ZN(n9789) );
  NAND2_X1 U12276 ( .A1(n9826), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9788) );
  INV_X1 U12277 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14317) );
  NAND2_X1 U12278 ( .A1(n9790), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9793) );
  NAND2_X1 U12279 ( .A1(n9791), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9792) );
  OAI211_X1 U12280 ( .C1(n6476), .C2(n14317), .A(n9793), .B(n9792), .ZN(n14092) );
  NAND2_X1 U12281 ( .A1(n9409), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9797) );
  INV_X1 U12282 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9794) );
  OR2_X1 U12283 ( .A1(n6475), .A2(n9794), .ZN(n9796) );
  INV_X1 U12284 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14415) );
  OR2_X1 U12285 ( .A1(n9814), .A2(n14415), .ZN(n9795) );
  AND3_X1 U12286 ( .A1(n9797), .A2(n9796), .A3(n9795), .ZN(n9805) );
  INV_X1 U12287 ( .A(n9805), .ZN(n14022) );
  OAI21_X1 U12288 ( .B1(n14092), .B2(n11901), .A(n14022), .ZN(n9798) );
  NAND2_X1 U12289 ( .A1(n9802), .A2(n14092), .ZN(n9831) );
  INV_X1 U12290 ( .A(n9803), .ZN(n9804) );
  NAND2_X1 U12291 ( .A1(n9804), .A2(n11981), .ZN(n9806) );
  AOI21_X1 U12292 ( .B1(n9831), .B2(n9806), .A(n9805), .ZN(n9807) );
  AOI21_X1 U12293 ( .B1(n9851), .B2(n9821), .A(n9807), .ZN(n9843) );
  NAND2_X1 U12294 ( .A1(n9409), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9818) );
  INV_X1 U12295 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9809) );
  NOR2_X1 U12296 ( .A1(n9810), .A2(n9809), .ZN(n12356) );
  NAND2_X1 U12297 ( .A1(n9331), .A2(n12356), .ZN(n9817) );
  INV_X1 U12298 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9811) );
  OR2_X1 U12299 ( .A1(n6475), .A2(n9811), .ZN(n9816) );
  INV_X1 U12300 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9813) );
  OR2_X1 U12301 ( .A1(n9814), .A2(n9813), .ZN(n9815) );
  NAND4_X1 U12302 ( .A1(n9818), .A2(n9817), .A3(n9816), .A4(n9815), .ZN(n14023) );
  NAND2_X1 U12303 ( .A1(n12281), .A2(n9825), .ZN(n9820) );
  NAND2_X1 U12304 ( .A1(n9826), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9819) );
  MUX2_X1 U12305 ( .A(n14023), .B(n14327), .S(n9821), .Z(n9838) );
  INV_X1 U12306 ( .A(n9838), .ZN(n9822) );
  MUX2_X1 U12307 ( .A(n14327), .B(n14023), .S(n9821), .Z(n9837) );
  NAND2_X1 U12308 ( .A1(n9822), .A2(n9837), .ZN(n9823) );
  NAND2_X1 U12309 ( .A1(n9824), .A2(n9823), .ZN(n9835) );
  NAND2_X1 U12310 ( .A1(n13785), .A2(n9825), .ZN(n9828) );
  NAND2_X1 U12311 ( .A1(n9826), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n9827) );
  XNOR2_X1 U12312 ( .A(n14089), .B(n14092), .ZN(n9876) );
  NAND2_X1 U12313 ( .A1(n9829), .A2(n11901), .ZN(n10538) );
  INV_X1 U12314 ( .A(n10538), .ZN(n10603) );
  OR2_X1 U12315 ( .A1(n10600), .A2(n14626), .ZN(n11037) );
  OAI21_X1 U12316 ( .B1(n10564), .B2(n10603), .A(n11037), .ZN(n9834) );
  INV_X1 U12317 ( .A(n9834), .ZN(n9880) );
  NAND2_X1 U12318 ( .A1(n9876), .A2(n9880), .ZN(n9848) );
  MUX2_X1 U12319 ( .A(n14092), .B(n9830), .S(n14089), .Z(n9832) );
  NAND2_X1 U12320 ( .A1(n9832), .A2(n9831), .ZN(n9879) );
  NAND2_X1 U12321 ( .A1(n11981), .A2(n9833), .ZN(n10565) );
  AND2_X1 U12322 ( .A1(n9834), .A2(n10565), .ZN(n9875) );
  NAND2_X1 U12323 ( .A1(n9879), .A2(n9875), .ZN(n9888) );
  INV_X1 U12324 ( .A(n9888), .ZN(n9836) );
  NAND2_X1 U12325 ( .A1(n9836), .A2(n9835), .ZN(n9849) );
  INV_X1 U12326 ( .A(n9837), .ZN(n9839) );
  NAND2_X1 U12327 ( .A1(n9839), .A2(n9838), .ZN(n9842) );
  NAND2_X1 U12328 ( .A1(n9842), .A2(n9843), .ZN(n9841) );
  NAND2_X1 U12329 ( .A1(n9841), .A2(n9840), .ZN(n9847) );
  INV_X1 U12330 ( .A(n9842), .ZN(n9845) );
  INV_X1 U12331 ( .A(n9843), .ZN(n9844) );
  NAND2_X1 U12332 ( .A1(n9845), .A2(n9844), .ZN(n9846) );
  NAND2_X1 U12333 ( .A1(n9847), .A2(n9846), .ZN(n9889) );
  MUX2_X1 U12334 ( .A(n9849), .B(n9848), .S(n9889), .Z(n9850) );
  INV_X1 U12335 ( .A(n9850), .ZN(n9884) );
  XNOR2_X1 U12336 ( .A(n9851), .B(n14022), .ZN(n9873) );
  NAND2_X1 U12337 ( .A1(n14330), .A2(n13937), .ZN(n12363) );
  OR2_X1 U12338 ( .A1(n14330), .A2(n13937), .ZN(n9852) );
  NAND2_X1 U12339 ( .A1(n14337), .A2(n13948), .ZN(n12322) );
  OR2_X1 U12340 ( .A1(n14337), .A2(n13948), .ZN(n9853) );
  NAND2_X1 U12341 ( .A1(n12322), .A2(n9853), .ZN(n14100) );
  XNOR2_X1 U12342 ( .A(n14130), .B(n14143), .ZN(n14127) );
  XNOR2_X1 U12343 ( .A(n14361), .B(n14025), .ZN(n14191) );
  XNOR2_X1 U12344 ( .A(n14431), .B(n14197), .ZN(n14207) );
  NAND2_X1 U12345 ( .A1(n14231), .A2(n13956), .ZN(n9854) );
  INV_X1 U12346 ( .A(n14027), .ZN(n14727) );
  XNOR2_X1 U12347 ( .A(n14385), .B(n14727), .ZN(n12310) );
  XNOR2_X1 U12348 ( .A(n14735), .B(n14296), .ZN(n14270) );
  XNOR2_X1 U12349 ( .A(n12234), .B(n12224), .ZN(n14628) );
  XNOR2_X1 U12350 ( .A(n14602), .B(n14618), .ZN(n12109) );
  NAND2_X1 U12351 ( .A1(n14838), .A2(n14030), .ZN(n11755) );
  INV_X1 U12352 ( .A(n14030), .ZN(n11925) );
  NAND2_X1 U12353 ( .A1(n11853), .A2(n11925), .ZN(n9856) );
  INV_X1 U12354 ( .A(n14031), .ZN(n11766) );
  XNOR2_X1 U12355 ( .A(n11767), .B(n11766), .ZN(n11595) );
  INV_X1 U12356 ( .A(n14032), .ZN(n11592) );
  XNOR2_X1 U12357 ( .A(n15198), .B(n11592), .ZN(n11380) );
  XNOR2_X1 U12358 ( .A(n11536), .B(n14033), .ZN(n11539) );
  AND2_X1 U12359 ( .A1(n10849), .A2(n9857), .ZN(n11356) );
  NAND2_X1 U12360 ( .A1(n14038), .A2(n11339), .ZN(n9858) );
  NAND4_X1 U12361 ( .A1(n10851), .A2(n11356), .A3(n10989), .A4(n11048), .ZN(
        n9859) );
  INV_X1 U12362 ( .A(n14035), .ZN(n11447) );
  XNOR2_X1 U12363 ( .A(n14813), .B(n11447), .ZN(n11135) );
  XNOR2_X1 U12364 ( .A(n11193), .B(n14036), .ZN(n11121) );
  NOR3_X1 U12365 ( .A1(n9859), .A2(n11135), .A3(n11121), .ZN(n9860) );
  XNOR2_X1 U12366 ( .A(n11617), .B(n14034), .ZN(n11369) );
  NAND3_X1 U12367 ( .A1(n11539), .A2(n9860), .A3(n11369), .ZN(n9861) );
  NOR4_X1 U12368 ( .A1(n11638), .A2(n11595), .A3(n11380), .A4(n9861), .ZN(
        n9862) );
  NAND3_X1 U12369 ( .A1(n12109), .A2(n9862), .A3(n11757), .ZN(n9863) );
  NOR3_X1 U12370 ( .A1(n7513), .A2(n14628), .A3(n9863), .ZN(n9864) );
  XNOR2_X1 U12371 ( .A(n14721), .B(n14028), .ZN(n12307) );
  NAND4_X1 U12372 ( .A1(n14270), .A2(n12330), .A3(n9864), .A4(n12307), .ZN(
        n9865) );
  NOR2_X1 U12373 ( .A1(n12310), .A2(n9865), .ZN(n9866) );
  NAND4_X1 U12374 ( .A1(n14207), .A2(n14225), .A3(n9866), .A4(n14247), .ZN(
        n9867) );
  NOR2_X1 U12375 ( .A1(n14191), .A2(n9867), .ZN(n9868) );
  XNOR2_X1 U12376 ( .A(n14356), .B(n14196), .ZN(n14176) );
  NAND3_X1 U12377 ( .A1(n14127), .A2(n9868), .A3(n14176), .ZN(n9869) );
  NOR2_X1 U12378 ( .A1(n14100), .A2(n9869), .ZN(n9871) );
  XNOR2_X1 U12379 ( .A(n14351), .B(n14142), .ZN(n14162) );
  NAND2_X1 U12380 ( .A1(n14346), .A2(n14159), .ZN(n12340) );
  OR2_X1 U12381 ( .A1(n14346), .A2(n14159), .ZN(n9870) );
  NAND2_X1 U12382 ( .A1(n12340), .A2(n9870), .ZN(n14140) );
  AND4_X1 U12383 ( .A1(n12341), .A2(n9871), .A3(n14162), .A4(n14140), .ZN(
        n9872) );
  XNOR2_X1 U12384 ( .A(n14327), .B(n14023), .ZN(n12365) );
  NAND4_X1 U12385 ( .A1(n9876), .A2(n9873), .A3(n9872), .A4(n12365), .ZN(n9874) );
  XNOR2_X1 U12386 ( .A(n9874), .B(n14626), .ZN(n9882) );
  INV_X1 U12387 ( .A(n9875), .ZN(n9877) );
  OAI21_X1 U12388 ( .B1(n9877), .B2(n9876), .A(n9879), .ZN(n9878) );
  OAI21_X1 U12389 ( .B1(n9880), .B2(n9879), .A(n9878), .ZN(n9881) );
  OAI21_X1 U12390 ( .B1(n9882), .B2(n10565), .A(n9881), .ZN(n9883) );
  NOR2_X1 U12391 ( .A1(n9884), .A2(n9883), .ZN(n9885) );
  NAND2_X1 U12392 ( .A1(n9891), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9892) );
  MUX2_X1 U12393 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9892), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n9894) );
  NAND2_X1 U12394 ( .A1(n9894), .A2(n9903), .ZN(n9973) );
  INV_X1 U12395 ( .A(n9973), .ZN(n9895) );
  NAND2_X1 U12396 ( .A1(n9895), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12245) );
  OAI21_X1 U12397 ( .B1(n9898), .B2(n9897), .A(n9896), .ZN(n9913) );
  INV_X1 U12398 ( .A(n9829), .ZN(n14475) );
  NAND2_X1 U12399 ( .A1(n14626), .A2(n11901), .ZN(n10560) );
  NAND2_X1 U12400 ( .A1(n10564), .A2(n10560), .ZN(n9910) );
  NAND2_X1 U12401 ( .A1(n9905), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9899) );
  MUX2_X1 U12402 ( .A(n9899), .B(P1_IR_REG_31__SCAN_IN), .S(n9900), .Z(n9902)
         );
  NAND2_X1 U12403 ( .A1(n9902), .A2(n9907), .ZN(n14466) );
  NAND2_X1 U12404 ( .A1(n9903), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9904) );
  MUX2_X1 U12405 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9904), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9906) );
  NOR2_X1 U12406 ( .A1(n14466), .A2(n14469), .ZN(n9909) );
  NAND3_X1 U12407 ( .A1(n9910), .A2(n10539), .A3(n9973), .ZN(n10572) );
  INV_X1 U12408 ( .A(n14459), .ZN(n12354) );
  INV_X1 U12409 ( .A(n14456), .ZN(n10156) );
  AND2_X2 U12410 ( .A1(n10564), .A2(n10156), .ZN(n14619) );
  NAND3_X1 U12411 ( .A1(n10595), .A2(n12354), .A3(n14619), .ZN(n9911) );
  OAI211_X1 U12412 ( .C1(n14475), .C2(n12245), .A(n9911), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9912) );
  NAND2_X1 U12413 ( .A1(n9913), .A2(n9912), .ZN(P1_U3242) );
  INV_X1 U12414 ( .A(n10539), .ZN(n10541) );
  INV_X1 U12415 ( .A(n10068), .ZN(n9914) );
  NAND2_X1 U12416 ( .A1(n9918), .A2(n9917), .ZN(n10858) );
  INV_X1 U12417 ( .A(n10858), .ZN(n9919) );
  AOI22_X1 U12418 ( .A1(n13311), .A2(n15413), .B1(n13576), .B2(n10323), .ZN(
        n9929) );
  INV_X1 U12419 ( .A(n9921), .ZN(n9922) );
  OR2_X1 U12420 ( .A1(n9923), .A2(n12284), .ZN(n9926) );
  NAND2_X1 U12421 ( .A1(n8221), .A2(n9924), .ZN(n9925) );
  INV_X2 U12422 ( .A(n13562), .ZN(n13631) );
  NAND2_X1 U12423 ( .A1(n9927), .A2(n13631), .ZN(n9928) );
  OAI211_X1 U12424 ( .C1(n10617), .C2(n9920), .A(n9929), .B(n9928), .ZN(n10619) );
  NAND3_X1 U12425 ( .A1(n9931), .A2(n14973), .A3(n9930), .ZN(n10624) );
  INV_X1 U12426 ( .A(n10624), .ZN(n9932) );
  NAND2_X1 U12427 ( .A1(n9933), .A2(n9932), .ZN(n9934) );
  MUX2_X1 U12428 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10619), .S(n14952), .Z(
        n9940) );
  INV_X1 U12429 ( .A(n9935), .ZN(n10999) );
  OR2_X1 U12430 ( .A1(n14964), .A2(n10999), .ZN(n13609) );
  OAI211_X1 U12431 ( .C1(n10626), .C2(n8994), .A(n11674), .B(n10868), .ZN(
        n10618) );
  OAI22_X1 U12432 ( .A1(n10617), .A2(n13609), .B1(n14958), .B2(n10618), .ZN(
        n9939) );
  INV_X1 U12433 ( .A(n9936), .ZN(n9937) );
  OR2_X2 U12434 ( .A1(n14964), .A2(n9937), .ZN(n13640) );
  OAI22_X1 U12435 ( .A1(n13640), .A2(n10626), .B1(n10429), .B2(n14950), .ZN(
        n9938) );
  OR3_X1 U12436 ( .A1(n9940), .A2(n9939), .A3(n9938), .ZN(P2_U3264) );
  NAND2_X1 U12437 ( .A1(n9975), .A2(P1_U3086), .ZN(n14472) );
  INV_X1 U12438 ( .A(n9942), .ZN(n9955) );
  INV_X1 U12439 ( .A(n10750), .ZN(n9943) );
  OAI222_X1 U12440 ( .A1(n14474), .A2(n9944), .B1(n14472), .B2(n9955), .C1(
        P1_U3086), .C2(n9943), .ZN(P1_U3353) );
  AND2_X1 U12441 ( .A1(n9975), .A2(P2_U3088), .ZN(n13792) );
  INV_X2 U12442 ( .A(n13792), .ZN(n13807) );
  NAND2_X1 U12443 ( .A1(n9945), .A2(P2_U3088), .ZN(n13805) );
  INV_X1 U12444 ( .A(n10150), .ZN(n10060) );
  OAI222_X1 U12445 ( .A1(n13807), .A2(n9946), .B1(n13805), .B2(n9947), .C1(
        P2_U3088), .C2(n10060), .ZN(P2_U3326) );
  INV_X1 U12446 ( .A(n14472), .ZN(n12244) );
  INV_X1 U12447 ( .A(n12244), .ZN(n14464) );
  INV_X1 U12448 ( .A(n10189), .ZN(n10171) );
  OAI222_X1 U12449 ( .A1(n14474), .A2(n7406), .B1(n14464), .B2(n9947), .C1(
        P1_U3086), .C2(n10171), .ZN(P1_U3354) );
  INV_X1 U12450 ( .A(n9948), .ZN(n9959) );
  INV_X1 U12451 ( .A(n14052), .ZN(n9949) );
  OAI222_X1 U12452 ( .A1(n14474), .A2(n9950), .B1(n14464), .B2(n9959), .C1(
        P1_U3086), .C2(n9949), .ZN(P1_U3352) );
  INV_X1 U12453 ( .A(n9951), .ZN(n9957) );
  OAI222_X1 U12454 ( .A1(n14474), .A2(n9952), .B1(n14472), .B2(n9957), .C1(
        P1_U3086), .C2(n10198), .ZN(P1_U3350) );
  INV_X1 U12455 ( .A(n9953), .ZN(n9962) );
  OAI222_X1 U12456 ( .A1(n14474), .A2(n9954), .B1(n14472), .B2(n9962), .C1(
        P1_U3086), .C2(n10786), .ZN(P1_U3351) );
  INV_X1 U12457 ( .A(n13805), .ZN(n12247) );
  INV_X1 U12458 ( .A(n12247), .ZN(n13794) );
  INV_X1 U12459 ( .A(n13323), .ZN(n10062) );
  OAI222_X1 U12460 ( .A1(n13807), .A2(n9956), .B1(n13794), .B2(n9955), .C1(
        P2_U3088), .C2(n10062), .ZN(P2_U3325) );
  INV_X1 U12461 ( .A(n10332), .ZN(n10339) );
  OAI222_X1 U12462 ( .A1(n13807), .A2(n9958), .B1(n13794), .B2(n9957), .C1(
        P2_U3088), .C2(n10339), .ZN(P2_U3322) );
  INV_X1 U12463 ( .A(n10081), .ZN(n14879) );
  OAI222_X1 U12464 ( .A1(n13807), .A2(n9960), .B1(n13794), .B2(n9959), .C1(
        P2_U3088), .C2(n14879), .ZN(P2_U3324) );
  INV_X1 U12465 ( .A(n10126), .ZN(n9961) );
  OAI222_X1 U12466 ( .A1(n13807), .A2(n9963), .B1(n13794), .B2(n9962), .C1(
        P2_U3088), .C2(n9961), .ZN(P2_U3323) );
  INV_X1 U12467 ( .A(n9964), .ZN(n9967) );
  OAI222_X1 U12468 ( .A1(n14474), .A2(n9965), .B1(n14472), .B2(n9967), .C1(
        P1_U3086), .C2(n14057), .ZN(P1_U3349) );
  INV_X1 U12469 ( .A(n13335), .ZN(n9966) );
  OAI222_X1 U12470 ( .A1(n13807), .A2(n9968), .B1(n13794), .B2(n9967), .C1(
        P2_U3088), .C2(n9966), .ZN(P2_U3321) );
  INV_X1 U12471 ( .A(n9969), .ZN(n9971) );
  INV_X1 U12472 ( .A(n10134), .ZN(n10065) );
  OAI222_X1 U12473 ( .A1(n13807), .A2(n9970), .B1(n13794), .B2(n9971), .C1(
        P2_U3088), .C2(n10065), .ZN(P2_U3320) );
  OAI222_X1 U12474 ( .A1(n14474), .A2(n9972), .B1(n14464), .B2(n9971), .C1(
        P1_U3086), .C2(n10220), .ZN(P1_U3348) );
  INV_X1 U12475 ( .A(n10568), .ZN(n10559) );
  NAND2_X1 U12476 ( .A1(n10559), .A2(n12245), .ZN(n10020) );
  NAND2_X1 U12477 ( .A1(n10564), .A2(n9973), .ZN(n9974) );
  NAND2_X1 U12478 ( .A1(n9974), .A2(n6853), .ZN(n10018) );
  AND2_X1 U12479 ( .A1(n10020), .A2(n10018), .ZN(n14080) );
  NOR2_X1 U12480 ( .A1(n14080), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12481 ( .A(n13175), .ZN(n11271) );
  NAND2_X1 U12482 ( .A1(n9945), .A2(P3_U3151), .ZN(n13178) );
  INV_X1 U12483 ( .A(n13178), .ZN(n13170) );
  AOI222_X1 U12484 ( .A1(n9976), .A2(n11271), .B1(n10390), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_4_), .C2(n13170), .ZN(n9977) );
  INV_X1 U12485 ( .A(n9977), .ZN(P3_U3291) );
  AOI222_X1 U12486 ( .A1(n9978), .A2(n11271), .B1(n13170), .B2(SI_2_), .C1(
        n10259), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9979) );
  INV_X1 U12487 ( .A(n9979), .ZN(P3_U3293) );
  INV_X1 U12488 ( .A(n9980), .ZN(n9981) );
  OAI222_X1 U12489 ( .A1(n13178), .A2(n9982), .B1(n13175), .B2(n9981), .C1(
        n12726), .C2(P3_U3151), .ZN(P3_U3283) );
  AOI222_X1 U12490 ( .A1(n9983), .A2(n11271), .B1(SI_5_), .B2(n13170), .C1(
        n10400), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9984) );
  INV_X1 U12491 ( .A(n9984), .ZN(P3_U3290) );
  AOI222_X1 U12492 ( .A1(n9985), .A2(n11271), .B1(SI_7_), .B2(n13170), .C1(
        n11292), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9986) );
  INV_X1 U12493 ( .A(n9986), .ZN(P3_U3288) );
  NAND2_X1 U12494 ( .A1(n14466), .A2(P1_B_REG_SCAN_IN), .ZN(n9987) );
  MUX2_X1 U12495 ( .A(P1_B_REG_SCAN_IN), .B(n9987), .S(n14469), .Z(n9988) );
  INV_X1 U12496 ( .A(n9988), .ZN(n9989) );
  INV_X1 U12497 ( .A(n10556), .ZN(n10547) );
  NAND2_X1 U12498 ( .A1(n10547), .A2(n10568), .ZN(n14794) );
  INV_X1 U12499 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9991) );
  NAND2_X1 U12500 ( .A1(n14465), .A2(n14466), .ZN(n10546) );
  INV_X1 U12501 ( .A(n10546), .ZN(n9990) );
  AOI22_X1 U12502 ( .A1(n6644), .A2(n9991), .B1(n9990), .B2(n9994), .ZN(
        P1_U3446) );
  INV_X1 U12503 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9996) );
  INV_X1 U12504 ( .A(n14469), .ZN(n9992) );
  INV_X1 U12505 ( .A(n10545), .ZN(n9995) );
  AOI22_X1 U12506 ( .A1(n6644), .A2(n9996), .B1(n9995), .B2(n9994), .ZN(
        P1_U3445) );
  AOI22_X1 U12507 ( .A1(n11271), .A2(n9997), .B1(P3_IR_REG_0__SCAN_IN), .B2(
        P3_STATE_REG_SCAN_IN), .ZN(n9998) );
  OAI21_X1 U12508 ( .B1(n9999), .B2(n12293), .A(n9998), .ZN(P3_U3295) );
  INV_X1 U12509 ( .A(n10000), .ZN(n10002) );
  INV_X1 U12510 ( .A(n13352), .ZN(n13349) );
  OAI222_X1 U12511 ( .A1(n13807), .A2(n10001), .B1(n13794), .B2(n10002), .C1(
        P2_U3088), .C2(n13349), .ZN(P2_U3319) );
  OAI222_X1 U12512 ( .A1(n14474), .A2(n10003), .B1(n14472), .B2(n10002), .C1(
        P1_U3086), .C2(n10281), .ZN(P1_U3347) );
  INV_X1 U12513 ( .A(SI_3_), .ZN(n10005) );
  OAI222_X1 U12514 ( .A1(P3_U3151), .A2(n10501), .B1(n12293), .B2(n10005), 
        .C1(n13175), .C2(n10004), .ZN(P3_U3292) );
  OAI222_X1 U12515 ( .A1(P3_U3151), .A2(n11286), .B1(n12293), .B2(n7426), .C1(
        n13175), .C2(n10006), .ZN(P3_U3287) );
  OAI222_X1 U12516 ( .A1(P3_U3151), .A2(n11949), .B1(n12293), .B2(n10008), 
        .C1(n13175), .C2(n10007), .ZN(P3_U3284) );
  OAI222_X1 U12517 ( .A1(P3_U3151), .A2(n11842), .B1(n12293), .B2(n10010), 
        .C1(n13175), .C2(n10009), .ZN(P3_U3285) );
  INV_X1 U12518 ( .A(n10416), .ZN(n10256) );
  OAI222_X1 U12519 ( .A1(n13175), .A2(n10012), .B1(n12293), .B2(n10011), .C1(
        P3_U3151), .C2(n10256), .ZN(P3_U3294) );
  INV_X1 U12520 ( .A(n10013), .ZN(n10015) );
  INV_X1 U12521 ( .A(SI_6_), .ZN(n10014) );
  OAI222_X1 U12522 ( .A1(n11028), .A2(P3_U3151), .B1(n13175), .B2(n10015), 
        .C1(n10014), .C2(n12293), .ZN(P3_U3289) );
  INV_X1 U12523 ( .A(SI_9_), .ZN(n10016) );
  OAI222_X1 U12524 ( .A1(n6905), .A2(P3_U3151), .B1(n13175), .B2(n10017), .C1(
        n10016), .C2(n12293), .ZN(P3_U3286) );
  INV_X1 U12525 ( .A(n14080), .ZN(n14792) );
  INV_X1 U12526 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10026) );
  INV_X1 U12527 ( .A(n10018), .ZN(n10019) );
  NAND2_X1 U12528 ( .A1(n10020), .A2(n10019), .ZN(n10158) );
  INV_X1 U12529 ( .A(n10158), .ZN(n10161) );
  INV_X1 U12530 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10022) );
  NAND2_X1 U12531 ( .A1(n12354), .A2(n9349), .ZN(n10021) );
  NAND2_X1 U12532 ( .A1(n10156), .A2(n10021), .ZN(n10740) );
  AOI21_X1 U12533 ( .B1(n14459), .B2(n10022), .A(n10740), .ZN(n10023) );
  INV_X1 U12534 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10741) );
  XNOR2_X1 U12535 ( .A(n10023), .B(n10741), .ZN(n10024) );
  AOI22_X1 U12536 ( .A1(n10161), .A2(n10024), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10025) );
  OAI21_X1 U12537 ( .B1(n14792), .B2(n10026), .A(n10025), .ZN(P1_U3243) );
  NOR2_X1 U12538 ( .A1(n10028), .A2(n10027), .ZN(n10032) );
  INV_X1 U12539 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10029) );
  NOR2_X1 U12540 ( .A1(n10054), .A2(n10029), .ZN(P3_U3237) );
  INV_X1 U12541 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10030) );
  NOR2_X1 U12542 ( .A1(n10032), .A2(n10030), .ZN(P3_U3239) );
  INV_X1 U12543 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10031) );
  NOR2_X1 U12544 ( .A1(n10032), .A2(n10031), .ZN(P3_U3238) );
  INV_X1 U12545 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n15224) );
  NOR2_X1 U12546 ( .A1(n10032), .A2(n15224), .ZN(P3_U3234) );
  CLKBUF_X1 U12547 ( .A(n10032), .Z(n10054) );
  INV_X1 U12548 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10033) );
  NOR2_X1 U12549 ( .A1(n10054), .A2(n10033), .ZN(P3_U3251) );
  INV_X1 U12550 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n15378) );
  NOR2_X1 U12551 ( .A1(n10054), .A2(n15378), .ZN(P3_U3253) );
  INV_X1 U12552 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10034) );
  NOR2_X1 U12553 ( .A1(n10054), .A2(n10034), .ZN(P3_U3252) );
  INV_X1 U12554 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10035) );
  NOR2_X1 U12555 ( .A1(n10054), .A2(n10035), .ZN(P3_U3255) );
  INV_X1 U12556 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10036) );
  NOR2_X1 U12557 ( .A1(n10032), .A2(n10036), .ZN(P3_U3240) );
  INV_X1 U12558 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10037) );
  NOR2_X1 U12559 ( .A1(n10032), .A2(n10037), .ZN(P3_U3262) );
  INV_X1 U12560 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n15246) );
  NOR2_X1 U12561 ( .A1(n10054), .A2(n15246), .ZN(P3_U3261) );
  INV_X1 U12562 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10038) );
  NOR2_X1 U12563 ( .A1(n10032), .A2(n10038), .ZN(P3_U3260) );
  INV_X1 U12564 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n15233) );
  NOR2_X1 U12565 ( .A1(n10054), .A2(n15233), .ZN(P3_U3259) );
  INV_X1 U12566 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10039) );
  NOR2_X1 U12567 ( .A1(n10032), .A2(n10039), .ZN(P3_U3258) );
  INV_X1 U12568 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10040) );
  NOR2_X1 U12569 ( .A1(n10054), .A2(n10040), .ZN(P3_U3257) );
  INV_X1 U12570 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10041) );
  NOR2_X1 U12571 ( .A1(n10054), .A2(n10041), .ZN(P3_U3263) );
  INV_X1 U12572 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10042) );
  NOR2_X1 U12573 ( .A1(n10054), .A2(n10042), .ZN(P3_U3248) );
  INV_X1 U12574 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10043) );
  NOR2_X1 U12575 ( .A1(n10054), .A2(n10043), .ZN(P3_U3254) );
  INV_X1 U12576 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10044) );
  NOR2_X1 U12577 ( .A1(n10054), .A2(n10044), .ZN(P3_U3246) );
  INV_X1 U12578 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10045) );
  NOR2_X1 U12579 ( .A1(n10032), .A2(n10045), .ZN(P3_U3236) );
  INV_X1 U12580 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10046) );
  NOR2_X1 U12581 ( .A1(n10032), .A2(n10046), .ZN(P3_U3235) );
  INV_X1 U12582 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10047) );
  NOR2_X1 U12583 ( .A1(n10054), .A2(n10047), .ZN(P3_U3250) );
  INV_X1 U12584 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10048) );
  NOR2_X1 U12585 ( .A1(n10054), .A2(n10048), .ZN(P3_U3256) );
  INV_X1 U12586 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10049) );
  NOR2_X1 U12587 ( .A1(n10032), .A2(n10049), .ZN(P3_U3241) );
  INV_X1 U12588 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n15359) );
  NOR2_X1 U12589 ( .A1(n10054), .A2(n15359), .ZN(P3_U3247) );
  INV_X1 U12590 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10050) );
  NOR2_X1 U12591 ( .A1(n10032), .A2(n10050), .ZN(P3_U3243) );
  INV_X1 U12592 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10051) );
  NOR2_X1 U12593 ( .A1(n10054), .A2(n10051), .ZN(P3_U3245) );
  INV_X1 U12594 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10052) );
  NOR2_X1 U12595 ( .A1(n10054), .A2(n10052), .ZN(P3_U3244) );
  INV_X1 U12596 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10053) );
  NOR2_X1 U12597 ( .A1(n10054), .A2(n10053), .ZN(P3_U3249) );
  INV_X1 U12598 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10055) );
  NOR2_X1 U12599 ( .A1(n10054), .A2(n10055), .ZN(P3_U3242) );
  INV_X1 U12600 ( .A(n10056), .ZN(n10058) );
  OAI222_X1 U12601 ( .A1(n14474), .A2(n10057), .B1(n14464), .B2(n10058), .C1(
        n10300), .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U12602 ( .A(n10108), .ZN(n10361) );
  OAI222_X1 U12603 ( .A1(n13807), .A2(n10059), .B1(n13794), .B2(n10058), .C1(
        n10361), .C2(P2_U3088), .ZN(P2_U3318) );
  NOR2_X1 U12604 ( .A1(n10108), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10354) );
  INV_X1 U12605 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n15374) );
  MUX2_X1 U12606 ( .A(n15374), .B(P2_REG2_REG_1__SCAN_IN), .S(n10150), .Z(
        n10142) );
  INV_X1 U12607 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10141) );
  NOR3_X1 U12608 ( .A1(n10142), .A2(n10141), .A3(n10145), .ZN(n13319) );
  NOR2_X1 U12609 ( .A1(n10060), .A2(n15374), .ZN(n13318) );
  MUX2_X1 U12610 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10061), .S(n13323), .Z(
        n13320) );
  OAI21_X1 U12611 ( .B1(n13319), .B2(n13318), .A(n13320), .ZN(n13322) );
  OAI21_X1 U12612 ( .B1(n10061), .B2(n10062), .A(n13322), .ZN(n14884) );
  MUX2_X1 U12613 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10063), .S(n10081), .Z(
        n14883) );
  NAND2_X1 U12614 ( .A1(n14884), .A2(n14883), .ZN(n14882) );
  NAND2_X1 U12615 ( .A1(n10081), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10121) );
  MUX2_X1 U12616 ( .A(n11007), .B(P2_REG2_REG_4__SCAN_IN), .S(n10126), .Z(
        n10120) );
  AOI21_X1 U12617 ( .B1(n14882), .B2(n10121), .A(n10120), .ZN(n10123) );
  AOI21_X1 U12618 ( .B1(n10126), .B2(P2_REG2_REG_4__SCAN_IN), .A(n10123), .ZN(
        n10328) );
  MUX2_X1 U12619 ( .A(n11059), .B(P2_REG2_REG_5__SCAN_IN), .S(n10332), .Z(
        n10327) );
  NOR2_X1 U12620 ( .A1(n10328), .A2(n10327), .ZN(n13332) );
  NOR2_X1 U12621 ( .A1(n10339), .A2(n11059), .ZN(n13331) );
  MUX2_X1 U12622 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11078), .S(n13335), .Z(
        n13330) );
  OAI21_X1 U12623 ( .B1(n13332), .B2(n13331), .A(n13330), .ZN(n13334) );
  NAND2_X1 U12624 ( .A1(n13335), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10131) );
  INV_X1 U12625 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10064) );
  MUX2_X1 U12626 ( .A(n10064), .B(P2_REG2_REG_7__SCAN_IN), .S(n10134), .Z(
        n10130) );
  AOI21_X1 U12627 ( .B1(n13334), .B2(n10131), .A(n10130), .ZN(n13346) );
  NOR2_X1 U12628 ( .A1(n10065), .A2(n10064), .ZN(n13345) );
  MUX2_X1 U12629 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11253), .S(n13352), .Z(
        n13344) );
  OAI21_X1 U12630 ( .B1(n13346), .B2(n13345), .A(n13344), .ZN(n13348) );
  OAI21_X1 U12631 ( .B1(n11253), .B2(n13349), .A(n13348), .ZN(n10103) );
  MUX2_X1 U12632 ( .A(n11398), .B(P2_REG2_REG_9__SCAN_IN), .S(n10108), .Z(
        n10066) );
  NOR2_X1 U12633 ( .A1(n10103), .A2(n10066), .ZN(n10355) );
  AOI21_X1 U12634 ( .B1(n10354), .B2(n10103), .A(n10355), .ZN(n10112) );
  NAND2_X1 U12635 ( .A1(n10068), .A2(n10067), .ZN(n10070) );
  NAND2_X1 U12636 ( .A1(n10070), .A2(n10069), .ZN(n10071) );
  NAND2_X1 U12637 ( .A1(n10072), .A2(n10071), .ZN(n10104) );
  NOR2_X1 U12638 ( .A1(n8244), .A2(P2_U3088), .ZN(n13791) );
  AND2_X1 U12639 ( .A1(n10104), .A2(n13791), .ZN(n10099) );
  INV_X1 U12640 ( .A(n13796), .ZN(n13381) );
  AND2_X1 U12641 ( .A1(n10099), .A2(n13381), .ZN(n14939) );
  NOR2_X2 U12642 ( .A1(n10104), .A2(P2_U3088), .ZN(n14935) );
  AND2_X1 U12643 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10102) );
  MUX2_X1 U12644 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10073), .S(n10081), .Z(
        n14886) );
  MUX2_X1 U12645 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10074), .S(n13323), .Z(
        n10079) );
  MUX2_X1 U12646 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n10075), .S(n10150), .Z(
        n10077) );
  AND2_X1 U12647 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10076) );
  NAND2_X1 U12648 ( .A1(n10077), .A2(n10076), .ZN(n13313) );
  NAND2_X1 U12649 ( .A1(n10150), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n13312) );
  NAND2_X1 U12650 ( .A1(n13313), .A2(n13312), .ZN(n10078) );
  NAND2_X1 U12651 ( .A1(n10079), .A2(n10078), .ZN(n13316) );
  NAND2_X1 U12652 ( .A1(n13323), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10080) );
  NAND2_X1 U12653 ( .A1(n13316), .A2(n10080), .ZN(n14887) );
  NAND2_X1 U12654 ( .A1(n14886), .A2(n14887), .ZN(n14885) );
  NAND2_X1 U12655 ( .A1(n10081), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10117) );
  NAND2_X1 U12656 ( .A1(n14885), .A2(n10117), .ZN(n10083) );
  INV_X1 U12657 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n15021) );
  MUX2_X1 U12658 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n15021), .S(n10126), .Z(
        n10082) );
  NAND2_X1 U12659 ( .A1(n10083), .A2(n10082), .ZN(n10335) );
  NAND2_X1 U12660 ( .A1(n10126), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10334) );
  NAND2_X1 U12661 ( .A1(n10335), .A2(n10334), .ZN(n10086) );
  INV_X1 U12662 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10084) );
  MUX2_X1 U12663 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10084), .S(n10332), .Z(
        n10085) );
  NAND2_X1 U12664 ( .A1(n10086), .A2(n10085), .ZN(n13338) );
  NAND2_X1 U12665 ( .A1(n10332), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n13337) );
  NAND2_X1 U12666 ( .A1(n13338), .A2(n13337), .ZN(n10089) );
  INV_X1 U12667 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10087) );
  MUX2_X1 U12668 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10087), .S(n13335), .Z(
        n10088) );
  NAND2_X1 U12669 ( .A1(n10089), .A2(n10088), .ZN(n13340) );
  NAND2_X1 U12670 ( .A1(n13335), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10136) );
  NAND2_X1 U12671 ( .A1(n13340), .A2(n10136), .ZN(n10092) );
  INV_X1 U12672 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10090) );
  MUX2_X1 U12673 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10090), .S(n10134), .Z(
        n10091) );
  NAND2_X1 U12674 ( .A1(n10092), .A2(n10091), .ZN(n13355) );
  NAND2_X1 U12675 ( .A1(n10134), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n13354) );
  NAND2_X1 U12676 ( .A1(n13355), .A2(n13354), .ZN(n10095) );
  INV_X1 U12677 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10093) );
  MUX2_X1 U12678 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10093), .S(n13352), .Z(
        n10094) );
  NAND2_X1 U12679 ( .A1(n10095), .A2(n10094), .ZN(n13357) );
  NAND2_X1 U12680 ( .A1(n13352), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10096) );
  NAND2_X1 U12681 ( .A1(n13357), .A2(n10096), .ZN(n10105) );
  INV_X1 U12682 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10098) );
  MUX2_X1 U12683 ( .A(n10098), .B(P2_REG1_REG_9__SCAN_IN), .S(n10108), .Z(
        n10097) );
  OR2_X1 U12684 ( .A1(n10105), .A2(n10097), .ZN(n10363) );
  NAND3_X1 U12685 ( .A1(n10105), .A2(n10361), .A3(n10098), .ZN(n10100) );
  NAND2_X1 U12686 ( .A1(n10099), .A2(n13796), .ZN(n14873) );
  AOI21_X1 U12687 ( .B1(n10363), .B2(n10100), .A(n14873), .ZN(n10101) );
  AOI211_X1 U12688 ( .C1(n14935), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n10102), .B(
        n10101), .ZN(n10111) );
  NAND3_X1 U12689 ( .A1(n10103), .A2(n14939), .A3(P2_REG2_REG_9__SCAN_IN), 
        .ZN(n10107) );
  AND2_X1 U12690 ( .A1(n10104), .A2(n8244), .ZN(n14891) );
  AND2_X1 U12691 ( .A1(n14891), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14936) );
  INV_X1 U12692 ( .A(n14936), .ZN(n14880) );
  NAND3_X1 U12693 ( .A1(n14943), .A2(P2_REG1_REG_9__SCAN_IN), .A3(n10105), 
        .ZN(n10106) );
  NAND3_X1 U12694 ( .A1(n10107), .A2(n14880), .A3(n10106), .ZN(n10109) );
  NAND2_X1 U12695 ( .A1(n10109), .A2(n10108), .ZN(n10110) );
  OAI211_X1 U12696 ( .C1(n10112), .C2(n14874), .A(n10111), .B(n10110), .ZN(
        P2_U3223) );
  INV_X1 U12697 ( .A(n10113), .ZN(n10114) );
  OAI222_X1 U12698 ( .A1(n13178), .A2(n10115), .B1(n13175), .B2(n10114), .C1(
        n12717), .C2(P3_U3151), .ZN(P3_U3282) );
  INV_X1 U12699 ( .A(n14935), .ZN(n13368) );
  INV_X1 U12700 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14532) );
  MUX2_X1 U12701 ( .A(n15021), .B(P2_REG1_REG_4__SCAN_IN), .S(n10126), .Z(
        n10116) );
  NAND3_X1 U12702 ( .A1(n14885), .A2(n10117), .A3(n10116), .ZN(n10118) );
  NAND3_X1 U12703 ( .A1(n14943), .A2(n10335), .A3(n10118), .ZN(n10119) );
  NAND2_X1 U12704 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10530) );
  OAI211_X1 U12705 ( .C1(n13368), .C2(n14532), .A(n10119), .B(n10530), .ZN(
        n10125) );
  AND3_X1 U12706 ( .A1(n14882), .A2(n10121), .A3(n10120), .ZN(n10122) );
  NOR3_X1 U12707 ( .A1(n14874), .A2(n10123), .A3(n10122), .ZN(n10124) );
  AOI211_X1 U12708 ( .C1(n14936), .C2(n10126), .A(n10125), .B(n10124), .ZN(
        n10127) );
  INV_X1 U12709 ( .A(n10127), .ZN(P2_U3218) );
  OAI222_X1 U12710 ( .A1(P3_U3151), .A2(n12766), .B1(n12293), .B2(n10129), 
        .C1(n13175), .C2(n10128), .ZN(P3_U3281) );
  NAND3_X1 U12711 ( .A1(n13334), .A2(n10131), .A3(n10130), .ZN(n10132) );
  NAND2_X1 U12712 ( .A1(n10132), .A2(n14939), .ZN(n10140) );
  NAND2_X1 U12713 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10883) );
  OAI21_X1 U12714 ( .B1(n13368), .B2(n14543), .A(n10883), .ZN(n10133) );
  AOI21_X1 U12715 ( .B1(n10134), .B2(n14936), .A(n10133), .ZN(n10139) );
  MUX2_X1 U12716 ( .A(n10090), .B(P2_REG1_REG_7__SCAN_IN), .S(n10134), .Z(
        n10135) );
  NAND3_X1 U12717 ( .A1(n13340), .A2(n10136), .A3(n10135), .ZN(n10137) );
  NAND3_X1 U12718 ( .A1(n14943), .A2(n13355), .A3(n10137), .ZN(n10138) );
  OAI211_X1 U12719 ( .C1(n13346), .C2(n10140), .A(n10139), .B(n10138), .ZN(
        P2_U3221) );
  NOR2_X1 U12720 ( .A1(n14874), .A2(n10141), .ZN(n14872) );
  INV_X1 U12721 ( .A(n10142), .ZN(n10143) );
  AOI22_X1 U12722 ( .A1(n14872), .A2(P2_IR_REG_0__SCAN_IN), .B1(n14939), .B2(
        n10143), .ZN(n10152) );
  MUX2_X1 U12723 ( .A(n10075), .B(P2_REG1_REG_1__SCAN_IN), .S(n10150), .Z(
        n10144) );
  OAI21_X1 U12724 ( .B1(n7724), .B2(n10145), .A(n10144), .ZN(n10146) );
  AND3_X1 U12725 ( .A1(n14943), .A2(n13313), .A3(n10146), .ZN(n10149) );
  INV_X1 U12726 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10147) );
  OAI22_X1 U12727 ( .A1(n13368), .A2(n10147), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10429), .ZN(n10148) );
  AOI211_X1 U12728 ( .C1(n14936), .C2(n10150), .A(n10149), .B(n10148), .ZN(
        n10151) );
  OAI21_X1 U12729 ( .B1(n13319), .B2(n10152), .A(n10151), .ZN(P2_U3215) );
  AND2_X1 U12730 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10154) );
  INV_X1 U12731 ( .A(n10154), .ZN(n10737) );
  MUX2_X1 U12732 ( .A(n10153), .B(P1_REG2_REG_1__SCAN_IN), .S(n10189), .Z(
        n10160) );
  MUX2_X1 U12733 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n10153), .S(n10189), .Z(
        n10155) );
  NAND2_X1 U12734 ( .A1(n10155), .A2(n10154), .ZN(n10747) );
  INV_X1 U12735 ( .A(n10747), .ZN(n10159) );
  NAND2_X1 U12736 ( .A1(n10156), .A2(n12354), .ZN(n10157) );
  AOI211_X1 U12737 ( .C1(n10737), .C2(n10160), .A(n10159), .B(n14781), .ZN(
        n10168) );
  INV_X1 U12738 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10162) );
  MUX2_X1 U12739 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10162), .S(n10189), .Z(
        n10164) );
  AND2_X1 U12740 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10163) );
  NAND2_X1 U12741 ( .A1(n10164), .A2(n10163), .ZN(n10743) );
  MUX2_X1 U12742 ( .A(n10162), .B(P1_REG1_REG_1__SCAN_IN), .S(n10189), .Z(
        n10165) );
  OAI21_X1 U12743 ( .B1(n10022), .B2(n10741), .A(n10165), .ZN(n10166) );
  AND3_X1 U12744 ( .A1(n14083), .A2(n10743), .A3(n10166), .ZN(n10167) );
  NOR2_X1 U12745 ( .A1(n10168), .A2(n10167), .ZN(n10170) );
  AOI22_X1 U12746 ( .A1(n14080), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n10169) );
  OAI211_X1 U12747 ( .C1(n10171), .C2(n11995), .A(n10170), .B(n10169), .ZN(
        P1_U3244) );
  INV_X1 U12748 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n15216) );
  NAND2_X1 U12749 ( .A1(n14657), .A2(P3_U3897), .ZN(n10172) );
  OAI21_X1 U12750 ( .B1(P3_U3897), .B2(n15216), .A(n10172), .ZN(P3_U3502) );
  MUX2_X1 U12751 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n14305), .S(n14052), .Z(
        n10177) );
  MUX2_X1 U12752 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10173), .S(n10750), .Z(
        n10175) );
  NAND2_X1 U12753 ( .A1(n10189), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10746) );
  NAND2_X1 U12754 ( .A1(n10747), .A2(n10746), .ZN(n10174) );
  NAND2_X1 U12755 ( .A1(n10175), .A2(n10174), .ZN(n14043) );
  NAND2_X1 U12756 ( .A1(n10750), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14042) );
  NAND2_X1 U12757 ( .A1(n14043), .A2(n14042), .ZN(n10176) );
  NAND2_X1 U12758 ( .A1(n10177), .A2(n10176), .ZN(n14046) );
  NAND2_X1 U12759 ( .A1(n14052), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n10782) );
  MUX2_X1 U12760 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10178), .S(n10786), .Z(
        n10781) );
  AOI21_X1 U12761 ( .B1(n14046), .B2(n10782), .A(n10781), .ZN(n10780) );
  NOR2_X1 U12762 ( .A1(n10786), .A2(n10178), .ZN(n10343) );
  MUX2_X1 U12763 ( .A(n11137), .B(P1_REG2_REG_5__SCAN_IN), .S(n10198), .Z(
        n10344) );
  OAI21_X1 U12764 ( .B1(n10780), .B2(n10343), .A(n10344), .ZN(n14064) );
  INV_X1 U12765 ( .A(n10198), .ZN(n10347) );
  NAND2_X1 U12766 ( .A1(n10347), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n14063) );
  MUX2_X1 U12767 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9425), .S(n14057), .Z(
        n14062) );
  AOI21_X1 U12768 ( .B1(n14064), .B2(n14063), .A(n14062), .ZN(n14061) );
  NOR2_X1 U12769 ( .A1(n14057), .A2(n9425), .ZN(n10210) );
  MUX2_X1 U12770 ( .A(n10179), .B(P1_REG2_REG_7__SCAN_IN), .S(n10220), .Z(
        n10209) );
  OAI21_X1 U12771 ( .B1(n14061), .B2(n10210), .A(n10209), .ZN(n10212) );
  INV_X1 U12772 ( .A(n10220), .ZN(n10180) );
  NAND2_X1 U12773 ( .A1(n10180), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10182) );
  MUX2_X1 U12774 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11383), .S(n10281), .Z(
        n10181) );
  AOI21_X1 U12775 ( .B1(n10212), .B2(n10182), .A(n10181), .ZN(n10275) );
  NAND3_X1 U12776 ( .A1(n10212), .A2(n10182), .A3(n10181), .ZN(n10183) );
  NAND2_X1 U12777 ( .A1(n14074), .A2(n10183), .ZN(n10208) );
  INV_X1 U12778 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10184) );
  NOR2_X1 U12779 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10184), .ZN(n10186) );
  NOR2_X1 U12780 ( .A1(n11995), .A2(n10281), .ZN(n10185) );
  AOI211_X1 U12781 ( .C1(n14080), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10186), .B(
        n10185), .ZN(n10207) );
  INV_X1 U12782 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n14851) );
  MUX2_X1 U12783 ( .A(n14851), .B(P1_REG1_REG_8__SCAN_IN), .S(n10281), .Z(
        n10204) );
  INV_X1 U12784 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10187) );
  MUX2_X1 U12785 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10187), .S(n14052), .Z(
        n10193) );
  INV_X1 U12786 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10188) );
  MUX2_X1 U12787 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10188), .S(n10750), .Z(
        n10191) );
  NAND2_X1 U12788 ( .A1(n10189), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10742) );
  NAND2_X1 U12789 ( .A1(n10743), .A2(n10742), .ZN(n10190) );
  NAND2_X1 U12790 ( .A1(n10191), .A2(n10190), .ZN(n14048) );
  NAND2_X1 U12791 ( .A1(n10750), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14047) );
  NAND2_X1 U12792 ( .A1(n14048), .A2(n14047), .ZN(n10192) );
  NAND2_X1 U12793 ( .A1(n10193), .A2(n10192), .ZN(n14051) );
  NAND2_X1 U12794 ( .A1(n14052), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10775) );
  NAND2_X1 U12795 ( .A1(n14051), .A2(n10775), .ZN(n10195) );
  INV_X1 U12796 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10196) );
  MUX2_X1 U12797 ( .A(n10196), .B(P1_REG1_REG_4__SCAN_IN), .S(n10786), .Z(
        n10194) );
  NAND2_X1 U12798 ( .A1(n10195), .A2(n10194), .ZN(n10777) );
  OR2_X1 U12799 ( .A1(n10786), .A2(n10196), .ZN(n10197) );
  AND2_X1 U12800 ( .A1(n10777), .A2(n10197), .ZN(n10341) );
  INV_X1 U12801 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14848) );
  MUX2_X1 U12802 ( .A(n14848), .B(P1_REG1_REG_5__SCAN_IN), .S(n10198), .Z(
        n10342) );
  NAND2_X1 U12803 ( .A1(n10341), .A2(n10342), .ZN(n10340) );
  NAND2_X1 U12804 ( .A1(n10198), .A2(n14848), .ZN(n10199) );
  NAND2_X1 U12805 ( .A1(n10340), .A2(n10199), .ZN(n14068) );
  INV_X1 U12806 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n11329) );
  MUX2_X1 U12807 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n11329), .S(n14057), .Z(
        n14067) );
  OR2_X1 U12808 ( .A1(n14068), .A2(n14067), .ZN(n14070) );
  OR2_X1 U12809 ( .A1(n14057), .A2(n11329), .ZN(n10200) );
  NAND2_X1 U12810 ( .A1(n14070), .A2(n10200), .ZN(n10215) );
  INV_X1 U12811 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10201) );
  MUX2_X1 U12812 ( .A(n10201), .B(P1_REG1_REG_7__SCAN_IN), .S(n10220), .Z(
        n10214) );
  NAND2_X1 U12813 ( .A1(n10215), .A2(n10214), .ZN(n10213) );
  OR2_X1 U12814 ( .A1(n10220), .A2(n10201), .ZN(n10202) );
  AND2_X1 U12815 ( .A1(n10213), .A2(n10202), .ZN(n10203) );
  NAND2_X1 U12816 ( .A1(n10203), .A2(n10204), .ZN(n10286) );
  OAI21_X1 U12817 ( .B1(n10204), .B2(n10203), .A(n10286), .ZN(n10205) );
  NAND2_X1 U12818 ( .A1(n14083), .A2(n10205), .ZN(n10206) );
  OAI211_X1 U12819 ( .C1(n10275), .C2(n10208), .A(n10207), .B(n10206), .ZN(
        P1_U3251) );
  OR3_X1 U12820 ( .A1(n14061), .A2(n10210), .A3(n10209), .ZN(n10211) );
  NAND3_X1 U12821 ( .A1(n14074), .A2(n10212), .A3(n10211), .ZN(n10219) );
  NAND2_X1 U12822 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11471) );
  OAI211_X1 U12823 ( .C1(n10215), .C2(n10214), .A(n14083), .B(n10213), .ZN(
        n10216) );
  NAND2_X1 U12824 ( .A1(n11471), .A2(n10216), .ZN(n10217) );
  AOI21_X1 U12825 ( .B1(n14080), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n10217), .ZN(
        n10218) );
  OAI211_X1 U12826 ( .C1(n11995), .C2(n10220), .A(n10219), .B(n10218), .ZN(
        P1_U3250) );
  INV_X1 U12827 ( .A(n10221), .ZN(n10223) );
  INV_X1 U12828 ( .A(n10365), .ZN(n14892) );
  OAI222_X1 U12829 ( .A1(n13807), .A2(n10222), .B1(n13794), .B2(n10223), .C1(
        n14892), .C2(P2_U3088), .ZN(P2_U3317) );
  OAI222_X1 U12830 ( .A1(n14474), .A2(n10224), .B1(n14464), .B2(n10223), .C1(
        n10303), .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U12831 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10225) );
  INV_X1 U12832 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10227) );
  MUX2_X1 U12833 ( .A(n10227), .B(n10694), .S(n12824), .Z(n10510) );
  NAND2_X1 U12834 ( .A1(n10510), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10514) );
  NOR2_X1 U12835 ( .A1(n10411), .A2(n10514), .ZN(n10478) );
  INV_X1 U12836 ( .A(n10228), .ZN(n10477) );
  INV_X1 U12837 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10248) );
  INV_X1 U12838 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10258) );
  MUX2_X1 U12839 ( .A(n10248), .B(n10258), .S(n12824), .Z(n10229) );
  NAND2_X1 U12840 ( .A1(n10229), .A2(n10259), .ZN(n10495) );
  INV_X1 U12841 ( .A(n10229), .ZN(n10230) );
  INV_X1 U12842 ( .A(n10259), .ZN(n10483) );
  NAND2_X1 U12843 ( .A1(n10230), .A2(n10483), .ZN(n10231) );
  AND2_X1 U12844 ( .A1(n10495), .A2(n10231), .ZN(n10476) );
  OAI21_X1 U12845 ( .B1(n10478), .B2(n10477), .A(n10476), .ZN(n10496) );
  INV_X1 U12846 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10900) );
  INV_X1 U12847 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10232) );
  MUX2_X1 U12848 ( .A(n10900), .B(n10232), .S(n12824), .Z(n10233) );
  NAND2_X1 U12849 ( .A1(n10233), .A2(n10260), .ZN(n10236) );
  INV_X1 U12850 ( .A(n10233), .ZN(n10234) );
  NAND2_X1 U12851 ( .A1(n10234), .A2(n10501), .ZN(n10235) );
  NAND2_X1 U12852 ( .A1(n10236), .A2(n10235), .ZN(n10494) );
  AOI21_X1 U12853 ( .B1(n10496), .B2(n10495), .A(n10494), .ZN(n10498) );
  INV_X1 U12854 ( .A(n10236), .ZN(n10237) );
  NOR2_X1 U12855 ( .A1(n10498), .A2(n10237), .ZN(n10239) );
  MUX2_X1 U12856 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12824), .Z(n10384) );
  XOR2_X1 U12857 ( .A(n10390), .B(n10384), .Z(n10238) );
  NOR2_X1 U12858 ( .A1(n10239), .A2(n10238), .ZN(n10385) );
  AOI21_X1 U12859 ( .B1(n10239), .B2(n10238), .A(n10385), .ZN(n10273) );
  NAND2_X1 U12860 ( .A1(P3_U3897), .A2(n6870), .ZN(n12855) );
  OR2_X1 U12861 ( .A1(n10241), .A2(P3_U3151), .ZN(n12697) );
  NAND2_X1 U12862 ( .A1(n10240), .A2(n12697), .ZN(n10254) );
  NAND2_X1 U12863 ( .A1(n12657), .A2(n10241), .ZN(n10242) );
  NAND2_X1 U12864 ( .A1(n10243), .A2(n10242), .ZN(n10253) );
  INV_X1 U12865 ( .A(n10253), .ZN(n10244) );
  INV_X1 U12866 ( .A(n10266), .ZN(n10245) );
  MUX2_X1 U12867 ( .A(n12703), .B(n10245), .S(n6870), .Z(n12860) );
  NOR2_X1 U12868 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10227), .ZN(n10509) );
  NAND2_X1 U12869 ( .A1(n6891), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10247) );
  OAI21_X1 U12870 ( .B1(n10256), .B2(n10509), .A(n10247), .ZN(n10410) );
  NOR2_X1 U12871 ( .A1(n10410), .A2(n10226), .ZN(n10409) );
  INV_X1 U12872 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10941) );
  XNOR2_X1 U12873 ( .A(n10390), .B(n10941), .ZN(n10249) );
  AND3_X1 U12874 ( .A1(n10484), .A2(n10249), .A3(n7286), .ZN(n10252) );
  INV_X1 U12875 ( .A(n10250), .ZN(n10251) );
  AND2_X1 U12876 ( .A1(n10266), .A2(n10251), .ZN(n11289) );
  OAI21_X1 U12877 ( .B1(n10397), .B2(n10252), .A(n11289), .ZN(n10270) );
  AND2_X1 U12878 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n10819) );
  AOI21_X1 U12879 ( .B1(n15028), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n10819), .ZN(
        n10269) );
  INV_X1 U12880 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10694) );
  NOR2_X1 U12881 ( .A1(n10694), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10255) );
  INV_X1 U12882 ( .A(n10255), .ZN(n10506) );
  NOR2_X1 U12883 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10506), .ZN(n10257) );
  AOI21_X1 U12884 ( .B1(n10261), .B2(n10260), .A(n10262), .ZN(n10486) );
  INV_X1 U12885 ( .A(n10262), .ZN(n10264) );
  INV_X1 U12886 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10263) );
  XNOR2_X1 U12887 ( .A(n10390), .B(n10263), .ZN(n10265) );
  AND3_X1 U12888 ( .A1(n10487), .A2(n10265), .A3(n10264), .ZN(n10267) );
  AND2_X1 U12889 ( .A1(n10266), .A2(n12824), .ZN(n12862) );
  OAI21_X1 U12890 ( .B1(n10392), .B2(n10267), .A(n12862), .ZN(n10268) );
  NAND3_X1 U12891 ( .A1(n10270), .A2(n10269), .A3(n10268), .ZN(n10271) );
  AOI21_X1 U12892 ( .B1(n10390), .B2(n15054), .A(n10271), .ZN(n10272) );
  OAI21_X1 U12893 ( .B1(n10273), .B2(n12855), .A(n10272), .ZN(P3_U3186) );
  NOR2_X1 U12894 ( .A1(n10281), .A2(n11383), .ZN(n10274) );
  MUX2_X1 U12895 ( .A(n11601), .B(P1_REG2_REG_9__SCAN_IN), .S(n10300), .Z(
        n10276) );
  OAI21_X1 U12896 ( .B1(n10275), .B2(n10274), .A(n10276), .ZN(n10290) );
  OR3_X1 U12897 ( .A1(n10276), .A2(n10275), .A3(n10274), .ZN(n10277) );
  NAND3_X1 U12898 ( .A1(n10290), .A2(n10277), .A3(n14074), .ZN(n10280) );
  INV_X1 U12899 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10278) );
  NOR2_X1 U12900 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10278), .ZN(n11790) );
  AOI21_X1 U12901 ( .B1(n14080), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n11790), .ZN(
        n10279) );
  OAI211_X1 U12902 ( .C1(n11995), .C2(n10300), .A(n10280), .B(n10279), .ZN(
        n10289) );
  NAND2_X1 U12903 ( .A1(n10281), .A2(n14851), .ZN(n10284) );
  NAND2_X1 U12904 ( .A1(n10286), .A2(n10284), .ZN(n10282) );
  INV_X1 U12905 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10299) );
  MUX2_X1 U12906 ( .A(n10299), .B(P1_REG1_REG_9__SCAN_IN), .S(n10300), .Z(
        n10283) );
  NAND2_X1 U12907 ( .A1(n10282), .A2(n10283), .ZN(n10302) );
  INV_X1 U12908 ( .A(n10283), .ZN(n10285) );
  NAND3_X1 U12909 ( .A1(n10286), .A2(n10285), .A3(n10284), .ZN(n10287) );
  INV_X1 U12910 ( .A(n14083), .ZN(n14787) );
  AOI21_X1 U12911 ( .B1(n10302), .B2(n10287), .A(n14787), .ZN(n10288) );
  OR2_X1 U12912 ( .A1(n10289), .A2(n10288), .ZN(P1_U3252) );
  OAI21_X1 U12913 ( .B1(n11601), .B2(n10300), .A(n10290), .ZN(n10313) );
  MUX2_X1 U12914 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n9510), .S(n10303), .Z(
        n10291) );
  INV_X1 U12915 ( .A(n10291), .ZN(n10312) );
  NAND2_X1 U12916 ( .A1(n10313), .A2(n10312), .ZN(n10311) );
  INV_X1 U12917 ( .A(n10303), .ZN(n10318) );
  NAND2_X1 U12918 ( .A1(n10318), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10294) );
  INV_X1 U12919 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10292) );
  MUX2_X1 U12920 ( .A(n10292), .B(P1_REG2_REG_11__SCAN_IN), .S(n10450), .Z(
        n10293) );
  AOI21_X1 U12921 ( .B1(n10311), .B2(n10294), .A(n10293), .ZN(n10447) );
  NAND3_X1 U12922 ( .A1(n10311), .A2(n10294), .A3(n10293), .ZN(n10295) );
  NAND2_X1 U12923 ( .A1(n10295), .A2(n14074), .ZN(n10310) );
  NOR2_X1 U12924 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10296), .ZN(n11927) );
  INV_X1 U12925 ( .A(n10450), .ZN(n10376) );
  NOR2_X1 U12926 ( .A1(n11995), .A2(n10376), .ZN(n10297) );
  AOI211_X1 U12927 ( .C1(n14080), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n11927), 
        .B(n10297), .ZN(n10309) );
  INV_X1 U12928 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10298) );
  MUX2_X1 U12929 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10298), .S(n10450), .Z(
        n10306) );
  NAND2_X1 U12930 ( .A1(n10300), .A2(n10299), .ZN(n10301) );
  NAND2_X1 U12931 ( .A1(n10302), .A2(n10301), .ZN(n10317) );
  INV_X1 U12932 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14854) );
  MUX2_X1 U12933 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n14854), .S(n10303), .Z(
        n10316) );
  OR2_X1 U12934 ( .A1(n10317), .A2(n10316), .ZN(n10319) );
  NAND2_X1 U12935 ( .A1(n10318), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10304) );
  AND2_X1 U12936 ( .A1(n10319), .A2(n10304), .ZN(n10305) );
  NAND2_X1 U12937 ( .A1(n10305), .A2(n10306), .ZN(n10456) );
  OAI21_X1 U12938 ( .B1(n10306), .B2(n10305), .A(n10456), .ZN(n10307) );
  NAND2_X1 U12939 ( .A1(n10307), .A2(n14083), .ZN(n10308) );
  OAI211_X1 U12940 ( .C1(n10447), .C2(n10310), .A(n10309), .B(n10308), .ZN(
        P1_U3254) );
  AND2_X1 U12941 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11862) );
  OAI211_X1 U12942 ( .C1(n10313), .C2(n10312), .A(n10311), .B(n14074), .ZN(
        n10314) );
  OAI21_X1 U12943 ( .B1(n14517), .B2(n14792), .A(n10314), .ZN(n10315) );
  NOR2_X1 U12944 ( .A1(n11862), .A2(n10315), .ZN(n10322) );
  AOI21_X1 U12945 ( .B1(n10317), .B2(n10316), .A(n14787), .ZN(n10320) );
  INV_X1 U12946 ( .A(n11995), .ZN(n14784) );
  AOI22_X1 U12947 ( .A1(n10320), .A2(n10319), .B1(n10318), .B2(n14784), .ZN(
        n10321) );
  NAND2_X1 U12948 ( .A1(n10322), .A2(n10321), .ZN(P1_U3253) );
  CLKBUF_X2 U12949 ( .A(P2_U3947), .Z(n14856) );
  NAND2_X1 U12950 ( .A1(n14856), .A2(n10323), .ZN(n10324) );
  OAI21_X1 U12951 ( .B1(n14856), .B2(n9350), .A(n10324), .ZN(P2_U3531) );
  INV_X1 U12952 ( .A(n10325), .ZN(n10326) );
  OAI222_X1 U12953 ( .A1(n13178), .A2(n15360), .B1(n13175), .B2(n10326), .C1(
        n12782), .C2(P3_U3151), .ZN(P3_U3280) );
  NAND2_X1 U12954 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10661) );
  AOI211_X1 U12955 ( .C1(n10328), .C2(n10327), .A(n13332), .B(n14874), .ZN(
        n10329) );
  INV_X1 U12956 ( .A(n10329), .ZN(n10330) );
  NAND2_X1 U12957 ( .A1(n10661), .A2(n10330), .ZN(n10331) );
  AOI21_X1 U12958 ( .B1(n14935), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n10331), .ZN(
        n10338) );
  MUX2_X1 U12959 ( .A(n10084), .B(P2_REG1_REG_5__SCAN_IN), .S(n10332), .Z(
        n10333) );
  NAND3_X1 U12960 ( .A1(n10335), .A2(n10334), .A3(n10333), .ZN(n10336) );
  NAND3_X1 U12961 ( .A1(n14943), .A2(n13338), .A3(n10336), .ZN(n10337) );
  OAI211_X1 U12962 ( .C1(n14880), .C2(n10339), .A(n10338), .B(n10337), .ZN(
        P2_U3219) );
  OAI21_X1 U12963 ( .B1(n10342), .B2(n10341), .A(n10340), .ZN(n10352) );
  INV_X1 U12964 ( .A(n14064), .ZN(n10346) );
  NOR3_X1 U12965 ( .A1(n10780), .A2(n10344), .A3(n10343), .ZN(n10345) );
  NOR3_X1 U12966 ( .A1(n14781), .A2(n10346), .A3(n10345), .ZN(n10351) );
  INV_X1 U12967 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10349) );
  NAND2_X1 U12968 ( .A1(n14784), .A2(n10347), .ZN(n10348) );
  NAND2_X1 U12969 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n11442) );
  OAI211_X1 U12970 ( .C1(n10349), .C2(n14792), .A(n10348), .B(n11442), .ZN(
        n10350) );
  AOI211_X1 U12971 ( .C1(n14083), .C2(n10352), .A(n10351), .B(n10350), .ZN(
        n10353) );
  INV_X1 U12972 ( .A(n10353), .ZN(P1_U3248) );
  NOR2_X1 U12973 ( .A1(n10355), .A2(n10354), .ZN(n14897) );
  MUX2_X1 U12974 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n10356), .S(n10365), .Z(
        n14896) );
  NAND2_X1 U12975 ( .A1(n14897), .A2(n14896), .ZN(n14895) );
  OAI21_X1 U12976 ( .B1(n10356), .B2(n14892), .A(n14895), .ZN(n10358) );
  MUX2_X1 U12977 ( .A(n11677), .B(P2_REG2_REG_11__SCAN_IN), .S(n10702), .Z(
        n10357) );
  NOR2_X1 U12978 ( .A1(n10358), .A2(n10357), .ZN(n13364) );
  AOI21_X1 U12979 ( .B1(n10358), .B2(n10357), .A(n13364), .ZN(n10374) );
  INV_X1 U12980 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n11508) );
  NOR2_X1 U12981 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11508), .ZN(n10360) );
  INV_X1 U12982 ( .A(n10702), .ZN(n10378) );
  NOR2_X1 U12983 ( .A1(n14880), .A2(n10378), .ZN(n10359) );
  AOI211_X1 U12984 ( .C1(n14935), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n10360), 
        .B(n10359), .ZN(n10373) );
  NAND2_X1 U12985 ( .A1(n10361), .A2(n10098), .ZN(n10362) );
  AND2_X1 U12986 ( .A1(n10363), .A2(n10362), .ZN(n14900) );
  MUX2_X1 U12987 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n10364), .S(n10365), .Z(
        n14899) );
  NAND2_X1 U12988 ( .A1(n14900), .A2(n14899), .ZN(n14898) );
  NAND2_X1 U12989 ( .A1(n10365), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10370) );
  NAND2_X1 U12990 ( .A1(n14898), .A2(n10370), .ZN(n10368) );
  INV_X1 U12991 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10366) );
  MUX2_X1 U12992 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10366), .S(n10702), .Z(
        n10367) );
  NAND2_X1 U12993 ( .A1(n10368), .A2(n10367), .ZN(n13373) );
  MUX2_X1 U12994 ( .A(n10366), .B(P2_REG1_REG_11__SCAN_IN), .S(n10702), .Z(
        n10369) );
  NAND3_X1 U12995 ( .A1(n14898), .A2(n10370), .A3(n10369), .ZN(n10371) );
  NAND3_X1 U12996 ( .A1(n13373), .A2(n14943), .A3(n10371), .ZN(n10372) );
  OAI211_X1 U12997 ( .C1(n10374), .C2(n14874), .A(n10373), .B(n10372), .ZN(
        P2_U3225) );
  INV_X1 U12998 ( .A(n10375), .ZN(n10379) );
  OAI222_X1 U12999 ( .A1(n14474), .A2(n10377), .B1(n14464), .B2(n10379), .C1(
        P1_U3086), .C2(n10376), .ZN(P1_U3344) );
  OAI222_X1 U13000 ( .A1(n13807), .A2(n10380), .B1(n13794), .B2(n10379), .C1(
        P2_U3088), .C2(n10378), .ZN(P2_U3316) );
  INV_X1 U13001 ( .A(n10381), .ZN(n10382) );
  OAI222_X1 U13002 ( .A1(n13178), .A2(n10383), .B1(n13175), .B2(n10382), .C1(
        n12802), .C2(P3_U3151), .ZN(P3_U3279) );
  INV_X1 U13003 ( .A(n10384), .ZN(n10386) );
  AOI21_X1 U13004 ( .B1(n10390), .B2(n10386), .A(n10385), .ZN(n10829) );
  MUX2_X1 U13005 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12824), .Z(n10387) );
  OR2_X1 U13006 ( .A1(n10387), .A2(n6961), .ZN(n10828) );
  INV_X1 U13007 ( .A(n10828), .ZN(n10388) );
  AND2_X1 U13008 ( .A1(n10387), .A2(n6961), .ZN(n10830) );
  NOR2_X1 U13009 ( .A1(n10388), .A2(n10830), .ZN(n10389) );
  XNOR2_X1 U13010 ( .A(n10829), .B(n10389), .ZN(n10404) );
  NOR2_X1 U13011 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8345), .ZN(n10911) );
  INV_X1 U13012 ( .A(n10390), .ZN(n10398) );
  INV_X1 U13013 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15181) );
  AOI21_X1 U13014 ( .B1(n10394), .B2(n15181), .A(n10824), .ZN(n10395) );
  NOR2_X1 U13015 ( .A1(n10395), .A2(n15060), .ZN(n10396) );
  AOI211_X1 U13016 ( .C1(n15028), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n10911), .B(
        n10396), .ZN(n10403) );
  INV_X1 U13017 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15085) );
  OAI21_X1 U13018 ( .B1(n6512), .B2(P3_REG2_REG_5__SCAN_IN), .A(n6640), .ZN(
        n10401) );
  AOI22_X1 U13019 ( .A1(n10401), .A2(n11289), .B1(n10400), .B2(n15054), .ZN(
        n10402) );
  OAI211_X1 U13020 ( .C1(n12855), .C2(n10404), .A(n10403), .B(n10402), .ZN(
        P3_U3187) );
  AOI21_X1 U13021 ( .B1(n10406), .B2(n10225), .A(n10405), .ZN(n10408) );
  AOI22_X1 U13022 ( .A1(n15028), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10407) );
  OAI21_X1 U13023 ( .B1(n15060), .B2(n10408), .A(n10407), .ZN(n10415) );
  AOI21_X1 U13024 ( .B1(n10226), .B2(n10410), .A(n10409), .ZN(n10413) );
  AOI21_X1 U13025 ( .B1(n10514), .B2(n10411), .A(n10478), .ZN(n10412) );
  OAI22_X1 U13026 ( .A1(n15056), .A2(n10413), .B1(n10412), .B2(n12855), .ZN(
        n10414) );
  AOI211_X1 U13027 ( .C1(n10416), .C2(n15054), .A(n10415), .B(n10414), .ZN(
        n10417) );
  INV_X1 U13028 ( .A(n10417), .ZN(P3_U3183) );
  NOR2_X1 U13029 ( .A1(n10418), .A2(P2_U3088), .ZN(n10441) );
  INV_X1 U13030 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10638) );
  OAI22_X1 U13031 ( .A1(n8233), .A2(n10428), .B1(n8994), .B2(n13269), .ZN(
        n10420) );
  NAND2_X1 U13032 ( .A1(n10420), .A2(n10419), .ZN(n10423) );
  INV_X1 U13033 ( .A(n13578), .ZN(n13596) );
  OR2_X1 U13034 ( .A1(n14859), .A2(n13596), .ZN(n13254) );
  AOI22_X1 U13035 ( .A1(n13284), .A2(n9002), .B1(n10421), .B2(n14867), .ZN(
        n10422) );
  OAI211_X1 U13036 ( .C1(n10441), .C2(n10638), .A(n10423), .B(n10422), .ZN(
        P2_U3204) );
  INV_X1 U13037 ( .A(n10424), .ZN(n10503) );
  INV_X1 U13038 ( .A(n14474), .ZN(n14450) );
  AOI22_X1 U13039 ( .A1(n10676), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n14450), .ZN(n10425) );
  OAI21_X1 U13040 ( .B1(n10503), .B2(n14472), .A(n10425), .ZN(P1_U3343) );
  OAI21_X1 U13041 ( .B1(n10427), .B2(n10426), .A(n10435), .ZN(n10432) );
  INV_X1 U13042 ( .A(n14867), .ZN(n13281) );
  OR2_X1 U13043 ( .A1(n14859), .A2(n13594), .ZN(n12298) );
  OAI22_X1 U13044 ( .A1(n10626), .A2(n13281), .B1(n12298), .B2(n10428), .ZN(
        n10431) );
  OAI22_X1 U13045 ( .A1(n10441), .A2(n10429), .B1(n6836), .B2(n13254), .ZN(
        n10430) );
  AOI211_X1 U13046 ( .C1(n14860), .C2(n10432), .A(n10431), .B(n10430), .ZN(
        n10433) );
  INV_X1 U13047 ( .A(n10433), .ZN(P2_U3194) );
  AOI22_X1 U13048 ( .A1(n13189), .A2(n9002), .B1(n14860), .B2(n10434), .ZN(
        n10438) );
  INV_X1 U13049 ( .A(n10435), .ZN(n10437) );
  NOR3_X1 U13050 ( .A1(n10438), .A2(n10437), .A3(n10436), .ZN(n10444) );
  OAI22_X1 U13051 ( .A1(n14978), .A2(n13281), .B1(n12298), .B2(n9236), .ZN(
        n10443) );
  INV_X1 U13052 ( .A(n13310), .ZN(n10439) );
  OAI22_X1 U13053 ( .A1(n10441), .A2(n10440), .B1(n10439), .B2(n13254), .ZN(
        n10442) );
  NOR3_X1 U13054 ( .A1(n10444), .A2(n10443), .A3(n10442), .ZN(n10445) );
  OAI21_X1 U13055 ( .B1(n10446), .B2(n13269), .A(n10445), .ZN(P2_U3209) );
  MUX2_X1 U13056 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n9539), .S(n10676), .Z(
        n10449) );
  AOI21_X1 U13057 ( .B1(n10450), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10447), 
        .ZN(n10448) );
  NAND2_X1 U13058 ( .A1(n10448), .A2(n10449), .ZN(n10670) );
  OAI21_X1 U13059 ( .B1(n10449), .B2(n10448), .A(n10670), .ZN(n10463) );
  OR2_X1 U13060 ( .A1(n10450), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10454) );
  NAND2_X1 U13061 ( .A1(n10456), .A2(n10454), .ZN(n10452) );
  INV_X1 U13062 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10451) );
  MUX2_X1 U13063 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10451), .S(n10676), .Z(
        n10453) );
  NAND2_X1 U13064 ( .A1(n10452), .A2(n10453), .ZN(n10678) );
  INV_X1 U13065 ( .A(n10453), .ZN(n10455) );
  NAND3_X1 U13066 ( .A1(n10456), .A2(n10455), .A3(n10454), .ZN(n10457) );
  AOI21_X1 U13067 ( .B1(n10678), .B2(n10457), .A(n14787), .ZN(n10462) );
  INV_X1 U13068 ( .A(n10676), .ZN(n10460) );
  AND2_X1 U13069 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10458) );
  AOI21_X1 U13070 ( .B1(n14080), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n10458), 
        .ZN(n10459) );
  OAI21_X1 U13071 ( .B1(n10460), .B2(n11995), .A(n10459), .ZN(n10461) );
  AOI211_X1 U13072 ( .C1(n10463), .C2(n14074), .A(n10462), .B(n10461), .ZN(
        n10464) );
  INV_X1 U13073 ( .A(n10464), .ZN(P1_U3255) );
  AOI21_X1 U13074 ( .B1(n10467), .B2(n10466), .A(n10465), .ZN(n10468) );
  NOR2_X1 U13075 ( .A1(n15056), .A2(n10468), .ZN(n10475) );
  AOI21_X1 U13076 ( .B1(n10471), .B2(n10470), .A(n10469), .ZN(n10473) );
  AOI22_X1 U13077 ( .A1(n15028), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10472) );
  OAI21_X1 U13078 ( .B1(n15060), .B2(n10473), .A(n10472), .ZN(n10474) );
  NOR2_X1 U13079 ( .A1(n10475), .A2(n10474), .ZN(n10482) );
  INV_X1 U13080 ( .A(n10496), .ZN(n10480) );
  NOR3_X1 U13081 ( .A1(n10478), .A2(n10477), .A3(n10476), .ZN(n10479) );
  OAI21_X1 U13082 ( .B1(n10480), .B2(n10479), .A(n15052), .ZN(n10481) );
  OAI211_X1 U13083 ( .C1(n12860), .C2(n10483), .A(n10482), .B(n10481), .ZN(
        P3_U3184) );
  OAI21_X1 U13084 ( .B1(n10485), .B2(P3_REG2_REG_3__SCAN_IN), .A(n10484), .ZN(
        n10493) );
  INV_X1 U13085 ( .A(n10486), .ZN(n10489) );
  INV_X1 U13086 ( .A(n10487), .ZN(n10488) );
  AOI21_X1 U13087 ( .B1(n10232), .B2(n10489), .A(n10488), .ZN(n10491) );
  INV_X1 U13088 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10902) );
  NOR2_X1 U13089 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10902), .ZN(n10691) );
  AOI21_X1 U13090 ( .B1(n15028), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10691), .ZN(
        n10490) );
  OAI21_X1 U13091 ( .B1(n10491), .B2(n15060), .A(n10490), .ZN(n10492) );
  AOI21_X1 U13092 ( .B1(n11289), .B2(n10493), .A(n10492), .ZN(n10500) );
  AND3_X1 U13093 ( .A1(n10496), .A2(n10495), .A3(n10494), .ZN(n10497) );
  OAI21_X1 U13094 ( .B1(n10498), .B2(n10497), .A(n15052), .ZN(n10499) );
  OAI211_X1 U13095 ( .C1(n12860), .C2(n10501), .A(n10500), .B(n10499), .ZN(
        P3_U3185) );
  INV_X1 U13096 ( .A(n13370), .ZN(n10502) );
  OAI222_X1 U13097 ( .A1(n13807), .A2(n10504), .B1(n13794), .B2(n10503), .C1(
        n10502), .C2(P2_U3088), .ZN(P2_U3315) );
  NOR3_X1 U13098 ( .A1(n11289), .A2(n12862), .A3(n15052), .ZN(n10515) );
  INV_X1 U13099 ( .A(n15028), .ZN(n15066) );
  INV_X1 U13100 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n10505) );
  INV_X1 U13101 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10611) );
  OAI22_X1 U13102 ( .A1(n15066), .A2(n10505), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10611), .ZN(n10508) );
  NOR2_X1 U13103 ( .A1(n15060), .A2(n10506), .ZN(n10507) );
  AOI211_X1 U13104 ( .C1(n10509), .C2(n11289), .A(n10508), .B(n10507), .ZN(
        n10513) );
  OR2_X1 U13105 ( .A1(n12855), .A2(n10510), .ZN(n10511) );
  MUX2_X1 U13106 ( .A(n10511), .B(n12860), .S(P3_IR_REG_0__SCAN_IN), .Z(n10512) );
  OAI211_X1 U13107 ( .C1(n10515), .C2(n10514), .A(n10513), .B(n10512), .ZN(
        P3_U3182) );
  INV_X1 U13108 ( .A(n12831), .ZN(n12817) );
  INV_X1 U13109 ( .A(n10516), .ZN(n10517) );
  OAI222_X1 U13110 ( .A1(P3_U3151), .A2(n12817), .B1(n12293), .B2(n10518), 
        .C1(n13175), .C2(n10517), .ZN(P3_U3278) );
  AND2_X1 U13111 ( .A1(n15108), .A2(n10698), .ZN(n12523) );
  NOR2_X1 U13112 ( .A1(n12523), .A2(n15105), .ZN(n12503) );
  INV_X1 U13113 ( .A(n10519), .ZN(n10520) );
  NAND2_X1 U13114 ( .A1(n10520), .A2(n15169), .ZN(n10523) );
  CLKBUF_X1 U13115 ( .A(n10521), .Z(n10522) );
  INV_X1 U13116 ( .A(n15106), .ZN(n15095) );
  OAI22_X1 U13117 ( .A1(n12503), .A2(n10523), .B1(n10522), .B2(n15095), .ZN(
        n10696) );
  INV_X1 U13118 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10524) );
  NOR2_X1 U13119 ( .A1(n15176), .A2(n10524), .ZN(n10525) );
  AOI21_X1 U13120 ( .B1(n15176), .B2(n10696), .A(n10525), .ZN(n10526) );
  OAI21_X1 U13121 ( .B1(n10698), .B2(n13162), .A(n10526), .ZN(P3_U3390) );
  OAI21_X1 U13122 ( .B1(n10586), .B2(n10527), .A(n10659), .ZN(n10535) );
  NOR3_X1 U13123 ( .A1(n8233), .A2(n10528), .A3(n10527), .ZN(n10529) );
  INV_X1 U13124 ( .A(n12298), .ZN(n13289) );
  OAI21_X1 U13125 ( .B1(n10529), .B2(n13289), .A(n13310), .ZN(n10533) );
  INV_X1 U13126 ( .A(n13308), .ZN(n11070) );
  OAI21_X1 U13127 ( .B1(n13254), .B2(n11070), .A(n10530), .ZN(n10531) );
  AOI21_X1 U13128 ( .B1(n14984), .B2(n14867), .A(n10531), .ZN(n10532) );
  OAI211_X1 U13129 ( .C1(n14870), .C2(n11011), .A(n10533), .B(n10532), .ZN(
        n10534) );
  AOI21_X1 U13130 ( .B1(n14860), .B2(n10535), .A(n10534), .ZN(n10536) );
  INV_X1 U13131 ( .A(n10536), .ZN(P2_U3202) );
  NAND2_X2 U13132 ( .A1(n10539), .A2(n10600), .ZN(n13936) );
  NOR2_X4 U13133 ( .A1(n10538), .A2(n10537), .ZN(n14814) );
  NAND2_X2 U13134 ( .A1(n10539), .A2(n10599), .ZN(n13938) );
  OAI22_X1 U13135 ( .A1(n11351), .A2(n13938), .B1(n10741), .B2(n10539), .ZN(
        n10540) );
  AOI22_X1 U13136 ( .A1(n11045), .A2(n13902), .B1(P1_REG1_REG_0__SCAN_IN), 
        .B2(n10541), .ZN(n10542) );
  OAI21_X1 U13137 ( .B1(n11054), .B2(n13938), .A(n10542), .ZN(n10719) );
  NAND2_X1 U13138 ( .A1(n10543), .A2(n10719), .ZN(n10720) );
  OR2_X1 U13139 ( .A1(n10543), .A2(n10719), .ZN(n10544) );
  NAND2_X1 U13140 ( .A1(n10720), .A2(n10544), .ZN(n10736) );
  OAI21_X1 U13141 ( .B1(n10547), .B2(P1_D_REG_1__SCAN_IN), .A(n10546), .ZN(
        n10596) );
  INV_X1 U13142 ( .A(n10596), .ZN(n10563) );
  NOR2_X1 U13143 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n10551) );
  NOR4_X1 U13144 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n10550) );
  NOR4_X1 U13145 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n10549) );
  NOR4_X1 U13146 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n10548) );
  NAND4_X1 U13147 ( .A1(n10551), .A2(n10550), .A3(n10549), .A4(n10548), .ZN(
        n10558) );
  NOR4_X1 U13148 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n10555) );
  NOR4_X1 U13149 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n10554) );
  NOR4_X1 U13150 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n10553) );
  NOR4_X1 U13151 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n10552) );
  NAND4_X1 U13152 ( .A1(n10555), .A2(n10554), .A3(n10553), .A4(n10552), .ZN(
        n10557) );
  OAI21_X1 U13153 ( .B1(n10558), .B2(n10557), .A(n10556), .ZN(n10597) );
  NAND3_X1 U13154 ( .A1(n10598), .A2(n10563), .A3(n10597), .ZN(n10571) );
  AND2_X1 U13155 ( .A1(n10560), .A2(n11981), .ZN(n10561) );
  NAND2_X1 U13156 ( .A1(n9829), .A2(n10561), .ZN(n14837) );
  NOR2_X1 U13157 ( .A1(n10564), .A2(n14828), .ZN(n10562) );
  AND3_X1 U13158 ( .A1(n10563), .A2(n10597), .A3(n10595), .ZN(n11036) );
  NAND2_X1 U13159 ( .A1(n11036), .A2(n10598), .ZN(n14015) );
  AND2_X2 U13160 ( .A1(n10564), .A2(n14456), .ZN(n14620) );
  INV_X1 U13161 ( .A(n14620), .ZN(n14274) );
  AOI22_X1 U13162 ( .A1(n10736), .A2(n15206), .B1(n14703), .B2(n14040), .ZN(
        n10576) );
  INV_X1 U13163 ( .A(n10565), .ZN(n10566) );
  NAND2_X1 U13164 ( .A1(n9829), .A2(n10566), .ZN(n14613) );
  INV_X1 U13165 ( .A(n14613), .ZN(n11042) );
  NAND2_X1 U13166 ( .A1(n10567), .A2(n11042), .ZN(n10570) );
  INV_X1 U13167 ( .A(n10594), .ZN(n10569) );
  NAND2_X1 U13168 ( .A1(n10571), .A2(n10594), .ZN(n10574) );
  INV_X1 U13169 ( .A(n10572), .ZN(n10573) );
  NAND2_X1 U13170 ( .A1(n10574), .A2(n10573), .ZN(n11098) );
  OR2_X1 U13171 ( .A1(n11098), .A2(P1_U3086), .ZN(n10811) );
  AOI22_X1 U13172 ( .A1(n15197), .A2(n11045), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n10811), .ZN(n10575) );
  NAND2_X1 U13173 ( .A1(n10576), .A2(n10575), .ZN(P1_U3232) );
  INV_X1 U13174 ( .A(n10577), .ZN(n13164) );
  MUX2_X1 U13175 ( .A(n13166), .B(n13164), .S(n10578), .Z(n10580) );
  INV_X2 U13176 ( .A(n15089), .ZN(n15119) );
  AOI22_X1 U13177 ( .A1(n10696), .A2(n15122), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(n15119), .ZN(n10585) );
  INV_X1 U13178 ( .A(n13044), .ZN(n13027) );
  NAND2_X1 U13179 ( .A1(n13027), .A2(n10583), .ZN(n10584) );
  OAI211_X1 U13180 ( .C1(n10227), .C2(n15122), .A(n10585), .B(n10584), .ZN(
        P3_U3233) );
  INV_X1 U13181 ( .A(n10586), .ZN(n10587) );
  AOI211_X1 U13182 ( .C1(n10589), .C2(n10588), .A(n13269), .B(n10587), .ZN(
        n10593) );
  AOI22_X1 U13183 ( .A1(n13289), .A2(n13311), .B1(n13284), .B2(n13309), .ZN(
        n10591) );
  AOI22_X1 U13184 ( .A1(n14867), .A2(n10953), .B1(P2_U3088), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n10590) );
  OAI211_X1 U13185 ( .C1(n14870), .C2(P2_REG3_REG_3__SCAN_IN), .A(n10591), .B(
        n10590), .ZN(n10592) );
  OR2_X1 U13186 ( .A1(n10593), .A2(n10592), .ZN(P2_U3190) );
  NAND4_X1 U13187 ( .A1(n10597), .A2(n10596), .A3(n10595), .A4(n10594), .ZN(
        n10946) );
  AOI21_X1 U13188 ( .B1(n14475), .B2(n10599), .A(n11043), .ZN(n10602) );
  OAI21_X1 U13189 ( .B1(n9829), .B2(n11043), .A(n10600), .ZN(n10601) );
  NAND2_X1 U13190 ( .A1(n10602), .A2(n13940), .ZN(n14797) );
  NAND2_X1 U13191 ( .A1(n10603), .A2(n11043), .ZN(n14796) );
  OR2_X1 U13192 ( .A1(n11981), .A2(n11901), .ZN(n10604) );
  OAI21_X1 U13193 ( .B1(n9829), .B2(n14626), .A(n10604), .ZN(n14614) );
  NOR2_X1 U13194 ( .A1(n14842), .A2(n14255), .ZN(n10606) );
  NAND3_X1 U13195 ( .A1(n11045), .A2(n11981), .A3(n9829), .ZN(n10605) );
  NAND2_X1 U13196 ( .A1(n14040), .A2(n14620), .ZN(n11350) );
  OAI211_X1 U13197 ( .C1(n11356), .C2(n10606), .A(n10605), .B(n11350), .ZN(
        n10947) );
  NAND2_X1 U13198 ( .A1(n10947), .A2(n14845), .ZN(n10607) );
  OAI21_X1 U13199 ( .B1(n14845), .B2(n9345), .A(n10607), .ZN(P1_U3459) );
  NOR2_X1 U13200 ( .A1(n12474), .A2(P3_U3151), .ZN(n10731) );
  INV_X1 U13201 ( .A(n12503), .ZN(n10609) );
  OAI22_X1 U13202 ( .A1(n12472), .A2(n10522), .B1(n10698), .B2(n12477), .ZN(
        n10608) );
  AOI21_X1 U13203 ( .B1(n12468), .B2(n10609), .A(n10608), .ZN(n10610) );
  OAI21_X1 U13204 ( .B1(n10731), .B2(n10611), .A(n10610), .ZN(P3_U3172) );
  INV_X1 U13205 ( .A(n10612), .ZN(n10614) );
  INV_X1 U13206 ( .A(n10756), .ZN(n10762) );
  OAI222_X1 U13207 ( .A1(n14474), .A2(n10613), .B1(n14464), .B2(n10614), .C1(
        n10762), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U13208 ( .A(n11700), .ZN(n11710) );
  OAI222_X1 U13209 ( .A1(n13807), .A2(n10615), .B1(n13805), .B2(n10614), .C1(
        n11710), .C2(P2_U3088), .ZN(P2_U3314) );
  NOR2_X1 U13210 ( .A1(n10637), .A2(n10616), .ZN(n15000) );
  INV_X1 U13211 ( .A(n10617), .ZN(n10621) );
  INV_X1 U13212 ( .A(n10618), .ZN(n10620) );
  AOI211_X1 U13213 ( .C1(n15000), .C2(n10621), .A(n10620), .B(n10619), .ZN(
        n10634) );
  NAND3_X1 U13214 ( .A1(n14972), .A2(n10623), .A3(n10622), .ZN(n10630) );
  NAND2_X1 U13215 ( .A1(n15018), .A2(n14990), .ZN(n13778) );
  INV_X1 U13216 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10625) );
  OAI22_X1 U13217 ( .A1(n13778), .A2(n10626), .B1(n15018), .B2(n10625), .ZN(
        n10627) );
  INV_X1 U13218 ( .A(n10627), .ZN(n10628) );
  OAI21_X1 U13219 ( .B1(n10634), .B2(n15017), .A(n10628), .ZN(P2_U3433) );
  NOR2_X1 U13220 ( .A1(n10630), .A2(n10629), .ZN(n10632) );
  NAND2_X1 U13221 ( .A1(n15027), .A2(n14990), .ZN(n13736) );
  INV_X1 U13222 ( .A(n13736), .ZN(n13745) );
  AOI22_X1 U13223 ( .A1(n13745), .A2(n7233), .B1(n15025), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n10633) );
  OAI21_X1 U13224 ( .B1(n10634), .B2(n15025), .A(n10633), .ZN(P2_U3500) );
  INV_X1 U13225 ( .A(n14976), .ZN(n10642) );
  NOR2_X1 U13226 ( .A1(n8994), .A2(n10635), .ZN(n14975) );
  INV_X1 U13227 ( .A(n9920), .ZN(n14999) );
  OAI21_X1 U13228 ( .B1(n14999), .B2(n13631), .A(n14976), .ZN(n10636) );
  OAI21_X1 U13229 ( .B1(n9236), .B2(n13596), .A(n10636), .ZN(n14974) );
  AOI21_X1 U13230 ( .B1(n14975), .B2(n10637), .A(n14974), .ZN(n10639) );
  OAI22_X1 U13231 ( .A1(n14964), .A2(n10639), .B1(n10638), .B2(n14950), .ZN(
        n10640) );
  AOI21_X1 U13232 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n14964), .A(n10640), .ZN(
        n10641) );
  OAI21_X1 U13233 ( .B1(n10642), .B2(n13609), .A(n10641), .ZN(P2_U3265) );
  INV_X1 U13234 ( .A(n12839), .ZN(n12850) );
  INV_X1 U13235 ( .A(n10643), .ZN(n10644) );
  OAI222_X1 U13236 ( .A1(P3_U3151), .A2(n12850), .B1(n13178), .B2(n7434), .C1(
        n13175), .C2(n10644), .ZN(P3_U3277) );
  INV_X1 U13237 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10654) );
  OAI22_X1 U13238 ( .A1(n12472), .A2(n10894), .B1(n15104), .B2(n12477), .ZN(
        n10645) );
  AOI21_X1 U13239 ( .B1(n12470), .B2(n15108), .A(n10645), .ZN(n10653) );
  INV_X1 U13240 ( .A(n15105), .ZN(n10647) );
  NAND3_X1 U13241 ( .A1(n10647), .A2(n15111), .A3(n10646), .ZN(n10648) );
  OAI211_X1 U13242 ( .C1(n10650), .C2(n15110), .A(n10649), .B(n10648), .ZN(
        n10651) );
  NAND2_X1 U13243 ( .A1(n10651), .A2(n12468), .ZN(n10652) );
  OAI211_X1 U13244 ( .C1(n10731), .C2(n10654), .A(n10653), .B(n10652), .ZN(
        P3_U3162) );
  NAND2_X1 U13245 ( .A1(n13189), .A2(n13309), .ZN(n10655) );
  OAI21_X1 U13246 ( .B1(n10656), .B2(n13269), .A(n10655), .ZN(n10660) );
  INV_X1 U13247 ( .A(n10657), .ZN(n10658) );
  NAND3_X1 U13248 ( .A1(n10660), .A2(n10659), .A3(n10658), .ZN(n10667) );
  OAI21_X1 U13249 ( .B1(n13254), .B2(n11156), .A(n10661), .ZN(n10663) );
  NOR2_X1 U13250 ( .A1(n12298), .A2(n10965), .ZN(n10662) );
  NOR2_X1 U13251 ( .A1(n10663), .A2(n10662), .ZN(n10666) );
  NAND2_X1 U13252 ( .A1(n14867), .A2(n11071), .ZN(n10665) );
  OR2_X1 U13253 ( .A1(n14870), .A2(n11060), .ZN(n10664) );
  AND4_X1 U13254 ( .A1(n10667), .A2(n10666), .A3(n10665), .A4(n10664), .ZN(
        n10668) );
  OAI21_X1 U13255 ( .B1(n10669), .B2(n13269), .A(n10668), .ZN(P2_U3199) );
  OAI21_X1 U13256 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n10676), .A(n10670), 
        .ZN(n10673) );
  INV_X1 U13257 ( .A(n10673), .ZN(n10675) );
  MUX2_X1 U13258 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n10671), .S(n10756), .Z(
        n10674) );
  MUX2_X1 U13259 ( .A(n10671), .B(P1_REG2_REG_13__SCAN_IN), .S(n10756), .Z(
        n10672) );
  NOR2_X1 U13260 ( .A1(n10673), .A2(n10672), .ZN(n10764) );
  INV_X1 U13261 ( .A(n10764), .ZN(n10768) );
  OAI211_X1 U13262 ( .C1(n10675), .C2(n10674), .A(n10768), .B(n14074), .ZN(
        n10685) );
  NAND2_X1 U13263 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n12220)
         );
  INV_X1 U13264 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n14751) );
  MUX2_X1 U13265 ( .A(n14751), .B(P1_REG1_REG_13__SCAN_IN), .S(n10756), .Z(
        n10679) );
  OR2_X1 U13266 ( .A1(n10676), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10677) );
  NAND2_X1 U13267 ( .A1(n10678), .A2(n10677), .ZN(n10680) );
  AOI21_X1 U13268 ( .B1(n10679), .B2(n10680), .A(n14787), .ZN(n10681) );
  NAND2_X1 U13269 ( .A1(n10681), .A2(n10758), .ZN(n10682) );
  NAND2_X1 U13270 ( .A1(n12220), .A2(n10682), .ZN(n10683) );
  AOI21_X1 U13271 ( .B1(n14080), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10683), 
        .ZN(n10684) );
  OAI211_X1 U13272 ( .C1(n11995), .C2(n10762), .A(n10685), .B(n10684), .ZN(
        P1_U3256) );
  AOI21_X1 U13273 ( .B1(n10686), .B2(n10687), .A(n12462), .ZN(n10689) );
  NAND2_X1 U13274 ( .A1(n10689), .A2(n10688), .ZN(n10693) );
  INV_X1 U13275 ( .A(n12470), .ZN(n12441) );
  OAI22_X1 U13276 ( .A1(n12441), .A2(n10894), .B1(n10901), .B2(n12477), .ZN(
        n10690) );
  AOI211_X1 U13277 ( .C1(n12439), .C2(n15074), .A(n10691), .B(n10690), .ZN(
        n10692) );
  OAI211_X1 U13278 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12034), .A(n10693), .B(
        n10692), .ZN(P3_U3158) );
  NOR2_X1 U13279 ( .A1(n15193), .A2(n10694), .ZN(n10695) );
  AOI21_X1 U13280 ( .B1(n10696), .B2(n15193), .A(n10695), .ZN(n10697) );
  OAI21_X1 U13281 ( .B1(n10698), .B2(n13116), .A(n10697), .ZN(P3_U3459) );
  NOR2_X1 U13282 ( .A1(n10702), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n13363) );
  INV_X1 U13283 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11824) );
  NAND2_X1 U13284 ( .A1(n13370), .A2(n11824), .ZN(n10699) );
  OAI21_X1 U13285 ( .B1(n13370), .B2(n11824), .A(n10699), .ZN(n13362) );
  OAI21_X1 U13286 ( .B1(n13364), .B2(n13363), .A(n13362), .ZN(n13361) );
  OAI21_X1 U13287 ( .B1(n13370), .B2(P2_REG2_REG_12__SCAN_IN), .A(n13361), 
        .ZN(n10701) );
  MUX2_X1 U13288 ( .A(n7949), .B(P2_REG2_REG_13__SCAN_IN), .S(n11700), .Z(
        n10700) );
  NOR2_X1 U13289 ( .A1(n10701), .A2(n10700), .ZN(n11699) );
  AOI211_X1 U13290 ( .C1(n10701), .C2(n10700), .A(n14874), .B(n11699), .ZN(
        n10713) );
  XNOR2_X1 U13291 ( .A(n11700), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n10709) );
  NAND2_X1 U13292 ( .A1(n10702), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n13372) );
  XNOR2_X1 U13293 ( .A(n13370), .B(n10703), .ZN(n13371) );
  AND2_X1 U13294 ( .A1(n13372), .A2(n13371), .ZN(n10704) );
  INV_X1 U13295 ( .A(n13374), .ZN(n10706) );
  NOR2_X1 U13296 ( .A1(n13370), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10707) );
  INV_X1 U13297 ( .A(n10707), .ZN(n10705) );
  NAND2_X1 U13298 ( .A1(n10706), .A2(n10705), .ZN(n10708) );
  NOR3_X1 U13299 ( .A1(n13374), .A2(n10707), .A3(n10709), .ZN(n11708) );
  AOI211_X1 U13300 ( .C1(n10709), .C2(n10708), .A(n14873), .B(n11708), .ZN(
        n10712) );
  NAND2_X1 U13301 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n14857)
         );
  NAND2_X1 U13302 ( .A1(n14935), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n10710) );
  OAI211_X1 U13303 ( .C1(n14880), .C2(n11710), .A(n14857), .B(n10710), .ZN(
        n10711) );
  OR3_X1 U13304 ( .A1(n10713), .A2(n10712), .A3(n10711), .ZN(P2_U3227) );
  AOI22_X1 U13305 ( .A1(n11476), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n14450), .ZN(n10714) );
  OAI21_X1 U13306 ( .B1(n10790), .B2(n14472), .A(n10714), .ZN(P1_U3341) );
  OAI22_X1 U13307 ( .A1(n10810), .A2(n13938), .B1(n14802), .B2(n13936), .ZN(
        n10715) );
  XNOR2_X1 U13308 ( .A(n10715), .B(n10601), .ZN(n10717) );
  OAI22_X1 U13309 ( .A1(n10810), .A2(n10801), .B1(n14802), .B2(n13938), .ZN(
        n10716) );
  NOR2_X1 U13310 ( .A1(n10717), .A2(n10716), .ZN(n10803) );
  NAND2_X1 U13311 ( .A1(n10720), .A2(n7563), .ZN(n10721) );
  NAND2_X1 U13312 ( .A1(n10722), .A2(n10721), .ZN(n10805) );
  OAI21_X1 U13313 ( .B1(n10722), .B2(n10721), .A(n10805), .ZN(n10723) );
  NAND2_X1 U13314 ( .A1(n10723), .A2(n15206), .ZN(n10727) );
  NAND2_X1 U13315 ( .A1(n15200), .A2(n14619), .ZN(n14725) );
  OAI22_X1 U13316 ( .A1(n14728), .A2(n10724), .B1(n11054), .B2(n14725), .ZN(
        n10725) );
  AOI21_X1 U13317 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n10811), .A(n10725), .ZN(
        n10726) );
  OAI211_X1 U13318 ( .C1(n14802), .C2(n14707), .A(n10727), .B(n10726), .ZN(
        P1_U3222) );
  XOR2_X1 U13319 ( .A(n10729), .B(n10728), .Z(n10735) );
  OAI22_X1 U13320 ( .A1(n12472), .A2(n15096), .B1(n12477), .B2(n15088), .ZN(
        n10733) );
  INV_X1 U13321 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15227) );
  NOR2_X1 U13322 ( .A1(n10731), .A2(n15227), .ZN(n10732) );
  AOI211_X1 U13323 ( .C1(n12470), .C2(n10730), .A(n10733), .B(n10732), .ZN(
        n10734) );
  OAI21_X1 U13324 ( .B1(n12462), .B2(n10735), .A(n10734), .ZN(P3_U3177) );
  INV_X2 U13325 ( .A(P1_U4016), .ZN(n14039) );
  MUX2_X1 U13326 ( .A(n10737), .B(n10736), .S(n14459), .Z(n10738) );
  NOR2_X1 U13327 ( .A1(n10738), .A2(n14456), .ZN(n10739) );
  AOI211_X1 U13328 ( .C1(n10741), .C2(n10740), .A(n14039), .B(n10739), .ZN(
        n10789) );
  MUX2_X1 U13329 ( .A(n10188), .B(P1_REG1_REG_2__SCAN_IN), .S(n10750), .Z(
        n10744) );
  NAND3_X1 U13330 ( .A1(n10744), .A2(n10743), .A3(n10742), .ZN(n10745) );
  NAND3_X1 U13331 ( .A1(n14083), .A2(n14048), .A3(n10745), .ZN(n10754) );
  MUX2_X1 U13332 ( .A(n10173), .B(P1_REG2_REG_2__SCAN_IN), .S(n10750), .Z(
        n10748) );
  NAND3_X1 U13333 ( .A1(n10748), .A2(n10747), .A3(n10746), .ZN(n10749) );
  NAND3_X1 U13334 ( .A1(n14074), .A2(n14043), .A3(n10749), .ZN(n10753) );
  NAND2_X1 U13335 ( .A1(n14784), .A2(n10750), .ZN(n10752) );
  AOI22_X1 U13336 ( .A1(n14080), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10751) );
  NAND4_X1 U13337 ( .A1(n10754), .A2(n10753), .A3(n10752), .A4(n10751), .ZN(
        n10755) );
  OR2_X1 U13338 ( .A1(n10789), .A2(n10755), .ZN(P1_U3245) );
  INV_X1 U13339 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14743) );
  MUX2_X1 U13340 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n14743), .S(n11476), .Z(
        n10760) );
  NAND2_X1 U13341 ( .A1(n10756), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10757) );
  AND2_X1 U13342 ( .A1(n10758), .A2(n10757), .ZN(n10759) );
  NAND2_X1 U13343 ( .A1(n10759), .A2(n10760), .ZN(n11478) );
  OAI21_X1 U13344 ( .B1(n10760), .B2(n10759), .A(n11478), .ZN(n10772) );
  INV_X1 U13345 ( .A(n11476), .ZN(n11488) );
  NAND2_X1 U13346 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14710)
         );
  NAND2_X1 U13347 ( .A1(n14080), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n10761) );
  OAI211_X1 U13348 ( .C1(n11488), .C2(n11995), .A(n14710), .B(n10761), .ZN(
        n10771) );
  NOR2_X1 U13349 ( .A1(n10762), .A2(n10671), .ZN(n10765) );
  MUX2_X1 U13350 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n12097), .S(n11476), .Z(
        n10763) );
  NOR3_X1 U13351 ( .A1(n10764), .A2(n10765), .A3(n10763), .ZN(n10769) );
  INV_X1 U13352 ( .A(n10765), .ZN(n10767) );
  MUX2_X1 U13353 ( .A(n12097), .B(P1_REG2_REG_14__SCAN_IN), .S(n11476), .Z(
        n10766) );
  AOI21_X1 U13354 ( .B1(n10768), .B2(n10767), .A(n10766), .ZN(n11486) );
  NOR3_X1 U13355 ( .A1(n10769), .A2(n11486), .A3(n14781), .ZN(n10770) );
  AOI211_X1 U13356 ( .C1(n14083), .C2(n10772), .A(n10771), .B(n10770), .ZN(
        n10773) );
  INV_X1 U13357 ( .A(n10773), .ZN(P1_U3257) );
  INV_X1 U13358 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10779) );
  MUX2_X1 U13359 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10196), .S(n10786), .Z(
        n10774) );
  NAND3_X1 U13360 ( .A1(n14051), .A2(n10775), .A3(n10774), .ZN(n10776) );
  NAND3_X1 U13361 ( .A1(n14083), .A2(n10777), .A3(n10776), .ZN(n10778) );
  NAND2_X1 U13362 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n11198) );
  OAI211_X1 U13363 ( .C1(n10779), .C2(n14792), .A(n10778), .B(n11198), .ZN(
        n10788) );
  INV_X1 U13364 ( .A(n10780), .ZN(n10784) );
  NAND3_X1 U13365 ( .A1(n14046), .A2(n10782), .A3(n10781), .ZN(n10783) );
  NAND2_X1 U13366 ( .A1(n10784), .A2(n10783), .ZN(n10785) );
  OAI22_X1 U13367 ( .A1(n10786), .A2(n11995), .B1(n14781), .B2(n10785), .ZN(
        n10787) );
  OR3_X1 U13368 ( .A1(n10789), .A2(n10788), .A3(n10787), .ZN(P1_U3247) );
  INV_X1 U13369 ( .A(n14905), .ZN(n11713) );
  OAI222_X1 U13370 ( .A1(n13807), .A2(n10791), .B1(n13805), .B2(n10790), .C1(
        n11713), .C2(P2_U3088), .ZN(P2_U3313) );
  INV_X1 U13371 ( .A(n14991), .ZN(n11084) );
  AOI21_X1 U13372 ( .B1(n10793), .B2(n10792), .A(n13269), .ZN(n10794) );
  NAND2_X1 U13373 ( .A1(n10794), .A2(n10876), .ZN(n10798) );
  NOR2_X1 U13374 ( .A1(n14870), .A2(n11083), .ZN(n10796) );
  NAND2_X1 U13375 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n13328) );
  OAI21_X1 U13376 ( .B1(n12298), .B2(n11070), .A(n13328), .ZN(n10795) );
  AOI211_X1 U13377 ( .C1(n13284), .C2(n13306), .A(n10796), .B(n10795), .ZN(
        n10797) );
  OAI211_X1 U13378 ( .C1(n11084), .C2(n13281), .A(n10798), .B(n10797), .ZN(
        P2_U3211) );
  NAND2_X1 U13379 ( .A1(n14038), .A2(n11103), .ZN(n10799) );
  OAI21_X1 U13380 ( .B1(n11339), .B2(n13936), .A(n10799), .ZN(n10800) );
  XNOR2_X1 U13381 ( .A(n10800), .B(n13940), .ZN(n11107) );
  OAI22_X1 U13382 ( .A1(n10724), .A2(n10801), .B1(n11339), .B2(n13938), .ZN(
        n11108) );
  INV_X1 U13383 ( .A(n10803), .ZN(n10804) );
  NAND2_X1 U13384 ( .A1(n10805), .A2(n10804), .ZN(n10806) );
  NAND2_X1 U13385 ( .A1(n10806), .A2(n10807), .ZN(n11111) );
  OAI21_X1 U13386 ( .B1(n10807), .B2(n10806), .A(n11111), .ZN(n10808) );
  NAND2_X1 U13387 ( .A1(n10808), .A2(n15206), .ZN(n10813) );
  INV_X1 U13388 ( .A(n14619), .ZN(n14273) );
  NAND2_X1 U13389 ( .A1(n14037), .A2(n14620), .ZN(n10809) );
  OAI21_X1 U13390 ( .B1(n10810), .B2(n14273), .A(n10809), .ZN(n11336) );
  AOI22_X1 U13391 ( .A1(n10811), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n15200), 
        .B2(n11336), .ZN(n10812) );
  OAI211_X1 U13392 ( .C1(n11339), .C2(n14707), .A(n10813), .B(n10812), .ZN(
        P1_U3237) );
  INV_X1 U13393 ( .A(n10943), .ZN(n10822) );
  OAI21_X1 U13394 ( .B1(n10816), .B2(n10815), .A(n10814), .ZN(n10817) );
  NAND2_X1 U13395 ( .A1(n10817), .A2(n12468), .ZN(n10821) );
  OAI22_X1 U13396 ( .A1(n12441), .A2(n15096), .B1(n10942), .B2(n12477), .ZN(
        n10818) );
  AOI211_X1 U13397 ( .C1(n12439), .C2(n12711), .A(n10819), .B(n10818), .ZN(
        n10820) );
  OAI211_X1 U13398 ( .C1(n10822), .C2(n12034), .A(n10821), .B(n10820), .ZN(
        P3_U3170) );
  NAND2_X1 U13399 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n11028), .ZN(n10825) );
  OAI21_X1 U13400 ( .B1(P3_REG1_REG_6__SCAN_IN), .B2(n11028), .A(n10825), .ZN(
        n10826) );
  AOI21_X1 U13401 ( .B1(n10827), .B2(n10826), .A(n11016), .ZN(n10847) );
  INV_X1 U13402 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n10837) );
  MUX2_X1 U13403 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12824), .Z(n11018) );
  XNOR2_X1 U13404 ( .A(n11018), .B(n10845), .ZN(n10832) );
  OAI21_X1 U13405 ( .B1(n10832), .B2(n10831), .A(n11019), .ZN(n10833) );
  NAND2_X1 U13406 ( .A1(n15052), .A2(n10833), .ZN(n10836) );
  INV_X1 U13407 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10834) );
  NOR2_X1 U13408 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10834), .ZN(n11094) );
  INV_X1 U13409 ( .A(n11094), .ZN(n10835) );
  OAI211_X1 U13410 ( .C1(n15066), .C2(n10837), .A(n10836), .B(n10835), .ZN(
        n10844) );
  NAND2_X1 U13411 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n11028), .ZN(n10839) );
  OAI21_X1 U13412 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n11028), .A(n10839), .ZN(
        n10840) );
  AOI21_X1 U13413 ( .B1(n10841), .B2(n10840), .A(n11027), .ZN(n10842) );
  NOR2_X1 U13414 ( .A1(n10842), .A2(n15056), .ZN(n10843) );
  AOI211_X1 U13415 ( .C1(n15054), .C2(n10845), .A(n10844), .B(n10843), .ZN(
        n10846) );
  OAI21_X1 U13416 ( .B1(n10847), .B2(n15060), .A(n10846), .ZN(P3_U3188) );
  XNOR2_X1 U13417 ( .A(n10851), .B(n10985), .ZN(n11344) );
  OAI21_X1 U13418 ( .B1(n10852), .B2(n10851), .A(n10988), .ZN(n11342) );
  INV_X1 U13419 ( .A(n11044), .ZN(n10853) );
  AOI211_X1 U13420 ( .C1(n10982), .C2(n10853), .A(n14822), .B(n10994), .ZN(
        n11337) );
  AOI211_X1 U13421 ( .C1(n14614), .C2(n11342), .A(n11336), .B(n11337), .ZN(
        n10854) );
  OAI21_X1 U13422 ( .B1(n14819), .B2(n11344), .A(n10854), .ZN(n11175) );
  OAI22_X1 U13423 ( .A1(n14446), .A2(n11339), .B1(n14845), .B2(n9332), .ZN(
        n10855) );
  AOI21_X1 U13424 ( .B1(n11175), .B2(n14845), .A(n10855), .ZN(n10856) );
  INV_X1 U13425 ( .A(n10856), .ZN(P1_U3465) );
  OR2_X1 U13426 ( .A1(n9002), .A2(n7233), .ZN(n10857) );
  NAND2_X1 U13427 ( .A1(n10858), .A2(n10857), .ZN(n10859) );
  NAND2_X1 U13428 ( .A1(n10859), .A2(n6718), .ZN(n10917) );
  OAI21_X1 U13429 ( .B1(n10859), .B2(n6718), .A(n10917), .ZN(n14981) );
  INV_X1 U13430 ( .A(n14981), .ZN(n10870) );
  AOI22_X1 U13431 ( .A1(n13576), .A2(n9002), .B1(n13310), .B2(n15413), .ZN(
        n10866) );
  OAI21_X1 U13432 ( .B1(n10863), .B2(n10862), .A(n10921), .ZN(n10864) );
  NAND2_X1 U13433 ( .A1(n10864), .A2(n13631), .ZN(n10865) );
  OAI211_X1 U13434 ( .C1(n10870), .C2(n9920), .A(n10866), .B(n10865), .ZN(
        n14979) );
  INV_X1 U13435 ( .A(n14950), .ZN(n13637) );
  AOI22_X1 U13436 ( .A1(n14964), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n13637), .ZN(n10867) );
  OAI21_X1 U13437 ( .B1(n13640), .B2(n14978), .A(n10867), .ZN(n10872) );
  AOI21_X1 U13438 ( .B1(n10868), .B2(n10915), .A(n11080), .ZN(n10869) );
  NAND2_X1 U13439 ( .A1(n10869), .A2(n10926), .ZN(n14977) );
  OAI22_X1 U13440 ( .A1(n10870), .A2(n13609), .B1(n14958), .B2(n14977), .ZN(
        n10871) );
  AOI211_X1 U13441 ( .C1(n14952), .C2(n14979), .A(n10872), .B(n10871), .ZN(
        n10873) );
  INV_X1 U13442 ( .A(n10873), .ZN(P2_U3263) );
  INV_X1 U13443 ( .A(n14954), .ZN(n11166) );
  INV_X1 U13444 ( .A(n10874), .ZN(n10875) );
  AOI21_X1 U13445 ( .B1(n10876), .B2(n10875), .A(n13269), .ZN(n10880) );
  NOR3_X1 U13446 ( .A1(n8233), .A2(n10877), .A3(n11156), .ZN(n10879) );
  OAI21_X1 U13447 ( .B1(n10880), .B2(n10879), .A(n10878), .ZN(n10888) );
  INV_X1 U13448 ( .A(n14870), .ZN(n13277) );
  INV_X1 U13449 ( .A(n14951), .ZN(n10886) );
  NAND2_X1 U13450 ( .A1(n13307), .A2(n13576), .ZN(n10882) );
  NAND2_X1 U13451 ( .A1(n13305), .A2(n15413), .ZN(n10881) );
  NAND2_X1 U13452 ( .A1(n10882), .A2(n10881), .ZN(n11160) );
  INV_X1 U13453 ( .A(n11160), .ZN(n10884) );
  OAI21_X1 U13454 ( .B1(n14859), .B2(n10884), .A(n10883), .ZN(n10885) );
  AOI21_X1 U13455 ( .B1(n13277), .B2(n10886), .A(n10885), .ZN(n10887) );
  OAI211_X1 U13456 ( .C1(n11166), .C2(n13281), .A(n10888), .B(n10887), .ZN(
        P2_U3185) );
  INV_X1 U13457 ( .A(n10889), .ZN(n10892) );
  OAI222_X1 U13458 ( .A1(n13175), .A2(n10892), .B1(n12293), .B2(n10891), .C1(
        P3_U3151), .C2(n10890), .ZN(P3_U3275) );
  XNOR2_X1 U13459 ( .A(n10893), .B(n12505), .ZN(n15136) );
  INV_X1 U13460 ( .A(n15136), .ZN(n10905) );
  NOR2_X1 U13461 ( .A1(n15117), .A2(n12529), .ZN(n15102) );
  OAI22_X1 U13462 ( .A1(n10894), .A2(n15094), .B1(n10909), .B2(n15095), .ZN(
        n10899) );
  INV_X1 U13463 ( .A(n10895), .ZN(n10896) );
  AOI211_X1 U13464 ( .C1(n12505), .C2(n10897), .A(n15078), .B(n10896), .ZN(
        n10898) );
  AOI211_X1 U13465 ( .C1(n15136), .C2(n15075), .A(n10899), .B(n10898), .ZN(
        n15133) );
  MUX2_X1 U13466 ( .A(n10900), .B(n15133), .S(n15122), .Z(n10904) );
  NOR2_X1 U13467 ( .A1(n10901), .A2(n15169), .ZN(n15135) );
  AOI22_X1 U13468 ( .A1(n15083), .A2(n15135), .B1(n15119), .B2(n10902), .ZN(
        n10903) );
  OAI211_X1 U13469 ( .C1(n10905), .C2(n12944), .A(n10904), .B(n10903), .ZN(
        P3_U3230) );
  XOR2_X1 U13470 ( .A(n10907), .B(n10906), .Z(n10914) );
  OAI22_X1 U13471 ( .A1(n12441), .A2(n10909), .B1(n10908), .B2(n12477), .ZN(
        n10910) );
  AOI211_X1 U13472 ( .C1(n12439), .C2(n15073), .A(n10911), .B(n10910), .ZN(
        n10913) );
  NAND2_X1 U13473 ( .A1(n12474), .A2(n15082), .ZN(n10912) );
  OAI211_X1 U13474 ( .C1(n10914), .C2(n12462), .A(n10913), .B(n10912), .ZN(
        P3_U3167) );
  INV_X1 U13475 ( .A(n15000), .ZN(n13692) );
  OR2_X1 U13476 ( .A1(n13311), .A2(n10915), .ZN(n10916) );
  NAND2_X1 U13477 ( .A1(n10917), .A2(n10916), .ZN(n10919) );
  INV_X1 U13478 ( .A(n10922), .ZN(n10918) );
  NAND2_X1 U13479 ( .A1(n10919), .A2(n10918), .ZN(n10955) );
  OAI21_X1 U13480 ( .B1(n10919), .B2(n10918), .A(n10955), .ZN(n11183) );
  INV_X1 U13481 ( .A(n11183), .ZN(n10928) );
  NAND2_X1 U13482 ( .A1(n10921), .A2(n10920), .ZN(n10923) );
  OAI21_X1 U13483 ( .B1(n10923), .B2(n10922), .A(n10963), .ZN(n10924) );
  AOI222_X1 U13484 ( .A1(n13631), .A2(n10924), .B1(n13309), .B2(n13578), .C1(
        n13311), .C2(n13576), .ZN(n11179) );
  NAND2_X1 U13485 ( .A1(n10926), .A2(n10953), .ZN(n10925) );
  NAND2_X1 U13486 ( .A1(n10925), .A2(n11674), .ZN(n10927) );
  NOR2_X1 U13487 ( .A1(n10926), .A2(n10953), .ZN(n11008) );
  OR2_X1 U13488 ( .A1(n10927), .A2(n11008), .ZN(n11177) );
  OAI211_X1 U13489 ( .C1(n14994), .C2(n10928), .A(n11179), .B(n11177), .ZN(
        n10933) );
  INV_X1 U13490 ( .A(n10953), .ZN(n11178) );
  OAI22_X1 U13491 ( .A1(n13736), .A2(n11178), .B1(n15027), .B2(n10073), .ZN(
        n10929) );
  AOI21_X1 U13492 ( .B1(n10933), .B2(n15027), .A(n10929), .ZN(n10930) );
  INV_X1 U13493 ( .A(n10930), .ZN(P2_U3502) );
  INV_X1 U13494 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10931) );
  OAI22_X1 U13495 ( .A1(n13778), .A2(n11178), .B1(n15018), .B2(n10931), .ZN(
        n10932) );
  AOI21_X1 U13496 ( .B1(n10933), .B2(n15018), .A(n10932), .ZN(n10934) );
  INV_X1 U13497 ( .A(n10934), .ZN(P2_U3439) );
  XNOR2_X1 U13498 ( .A(n10935), .B(n12547), .ZN(n15138) );
  AOI22_X1 U13499 ( .A1(n15109), .A2(n12712), .B1(n12711), .B2(n15106), .ZN(
        n10939) );
  OAI211_X1 U13500 ( .C1(n10937), .C2(n12547), .A(n10936), .B(n15112), .ZN(
        n10938) );
  OAI211_X1 U13501 ( .C1(n15138), .C2(n15116), .A(n10939), .B(n10938), .ZN(
        n15139) );
  INV_X1 U13502 ( .A(n15139), .ZN(n10940) );
  MUX2_X1 U13503 ( .A(n10941), .B(n10940), .S(n15122), .Z(n10945) );
  NOR2_X1 U13504 ( .A1(n10942), .A2(n15169), .ZN(n15140) );
  AOI22_X1 U13505 ( .A1(n15083), .A2(n15140), .B1(n15119), .B2(n10943), .ZN(
        n10944) );
  OAI211_X1 U13506 ( .C1(n15138), .C2(n12944), .A(n10945), .B(n10944), .ZN(
        P3_U3229) );
  NOR2_X4 U13507 ( .A1(n10946), .A2(n11035), .ZN(n14388) );
  NAND2_X1 U13508 ( .A1(n10947), .A2(n14388), .ZN(n10948) );
  OAI21_X1 U13509 ( .B1(n14388), .B2(n10022), .A(n10948), .ZN(P1_U3528) );
  INV_X1 U13510 ( .A(n10949), .ZN(n10951) );
  INV_X1 U13511 ( .A(n14783), .ZN(n11489) );
  OAI222_X1 U13512 ( .A1(n14474), .A2(n10950), .B1(n14464), .B2(n10951), .C1(
        P1_U3086), .C2(n11489), .ZN(P1_U3340) );
  INV_X1 U13513 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10952) );
  INV_X1 U13514 ( .A(n14915), .ZN(n11715) );
  OAI222_X1 U13515 ( .A1(n13807), .A2(n10952), .B1(n13805), .B2(n10951), .C1(
        P2_U3088), .C2(n11715), .ZN(P2_U3312) );
  OR2_X1 U13516 ( .A1(n13310), .A2(n10953), .ZN(n10954) );
  NAND2_X1 U13517 ( .A1(n10955), .A2(n10954), .ZN(n11001) );
  NAND2_X1 U13518 ( .A1(n11001), .A2(n10964), .ZN(n10957) );
  OR2_X1 U13519 ( .A1(n14984), .A2(n13309), .ZN(n10956) );
  NAND2_X1 U13520 ( .A1(n10957), .A2(n10956), .ZN(n10959) );
  INV_X1 U13521 ( .A(n10967), .ZN(n10958) );
  NAND2_X1 U13522 ( .A1(n10959), .A2(n10958), .ZN(n11069) );
  OR2_X1 U13523 ( .A1(n10959), .A2(n10958), .ZN(n10960) );
  NAND2_X1 U13524 ( .A1(n11069), .A2(n10960), .ZN(n10961) );
  INV_X1 U13525 ( .A(n10961), .ZN(n11065) );
  NAND2_X1 U13526 ( .A1(n10961), .A2(n14999), .ZN(n10974) );
  OR2_X1 U13527 ( .A1(n11178), .A2(n13310), .ZN(n10962) );
  NAND2_X1 U13528 ( .A1(n14984), .A2(n10965), .ZN(n10966) );
  NAND2_X1 U13529 ( .A1(n10968), .A2(n10967), .ZN(n11073) );
  OAI21_X1 U13530 ( .B1(n10968), .B2(n10967), .A(n11073), .ZN(n10972) );
  NAND2_X1 U13531 ( .A1(n13309), .A2(n13576), .ZN(n10970) );
  NAND2_X1 U13532 ( .A1(n13307), .A2(n15413), .ZN(n10969) );
  NAND2_X1 U13533 ( .A1(n10970), .A2(n10969), .ZN(n10971) );
  AOI21_X1 U13534 ( .B1(n10972), .B2(n13631), .A(n10971), .ZN(n10973) );
  AND2_X1 U13535 ( .A1(n10974), .A2(n10973), .ZN(n11058) );
  NAND2_X1 U13536 ( .A1(n11008), .A2(n6696), .ZN(n11010) );
  INV_X1 U13537 ( .A(n11079), .ZN(n10975) );
  AOI211_X1 U13538 ( .C1(n11071), .C2(n11010), .A(n11080), .B(n10975), .ZN(
        n11062) );
  INV_X1 U13539 ( .A(n11062), .ZN(n10976) );
  OAI211_X1 U13540 ( .C1(n11065), .C2(n13692), .A(n11058), .B(n10976), .ZN(
        n10980) );
  OAI22_X1 U13541 ( .A1(n13778), .A2(n7105), .B1(n15018), .B2(n7791), .ZN(
        n10977) );
  AOI21_X1 U13542 ( .B1(n10980), .B2(n15018), .A(n10977), .ZN(n10978) );
  INV_X1 U13543 ( .A(n10978), .ZN(P2_U3445) );
  OAI22_X1 U13544 ( .A1(n13736), .A2(n7105), .B1(n15027), .B2(n10084), .ZN(
        n10979) );
  AOI21_X1 U13545 ( .B1(n10980), .B2(n15027), .A(n10979), .ZN(n10981) );
  INV_X1 U13546 ( .A(n10981), .ZN(P2_U3504) );
  NOR2_X1 U13547 ( .A1(n10982), .A2(n14038), .ZN(n10984) );
  NAND2_X1 U13548 ( .A1(n10982), .A2(n14038), .ZN(n10983) );
  INV_X1 U13549 ( .A(n10989), .ZN(n10986) );
  OAI21_X1 U13550 ( .B1(n10987), .B2(n10986), .A(n11118), .ZN(n14309) );
  INV_X1 U13551 ( .A(n14309), .ZN(n10995) );
  INV_X1 U13552 ( .A(n14797), .ZN(n14112) );
  OAI22_X1 U13553 ( .A1(n10724), .A2(n14273), .B1(n11194), .B2(n14274), .ZN(
        n10993) );
  AND2_X1 U13554 ( .A1(n10991), .A2(n14255), .ZN(n10992) );
  AOI211_X1 U13555 ( .C1(n14112), .C2(n14309), .A(n10993), .B(n10992), .ZN(
        n14304) );
  OAI211_X1 U13556 ( .C1(n10994), .C2(n14306), .A(n14814), .B(n11127), .ZN(
        n14310) );
  OAI211_X1 U13557 ( .C1(n10995), .C2(n14796), .A(n14304), .B(n14310), .ZN(
        n11186) );
  INV_X1 U13558 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10996) );
  OAI22_X1 U13559 ( .A1(n14446), .A2(n14306), .B1(n14845), .B2(n10996), .ZN(
        n10997) );
  AOI21_X1 U13560 ( .B1(n11186), .B2(n14845), .A(n10997), .ZN(n10998) );
  INV_X1 U13561 ( .A(n10998), .ZN(P1_U3468) );
  AND2_X1 U13562 ( .A1(n9920), .A2(n10999), .ZN(n11000) );
  XNOR2_X1 U13563 ( .A(n11001), .B(n11003), .ZN(n14983) );
  NAND2_X1 U13564 ( .A1(n11004), .A2(n13631), .ZN(n11006) );
  AOI22_X1 U13565 ( .A1(n13576), .A2(n13310), .B1(n13308), .B2(n15413), .ZN(
        n11005) );
  AND2_X1 U13566 ( .A1(n11006), .A2(n11005), .ZN(n14989) );
  MUX2_X1 U13567 ( .A(n14989), .B(n11007), .S(n14964), .Z(n11014) );
  OR2_X1 U13568 ( .A1(n11008), .A2(n6696), .ZN(n11009) );
  AND3_X1 U13569 ( .A1(n11010), .A2(n11674), .A3(n11009), .ZN(n14986) );
  OAI22_X1 U13570 ( .A1(n13640), .A2(n6696), .B1(n11011), .B2(n14950), .ZN(
        n11012) );
  AOI21_X1 U13571 ( .B1(n13649), .B2(n14986), .A(n11012), .ZN(n11013) );
  OAI211_X1 U13572 ( .C1(n13646), .C2(n14983), .A(n11014), .B(n11013), .ZN(
        P2_U3261) );
  INV_X1 U13573 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15185) );
  AOI21_X1 U13574 ( .B1(n15185), .B2(n11017), .A(n11275), .ZN(n11034) );
  INV_X1 U13575 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n11026) );
  MUX2_X1 U13576 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12824), .Z(n11295) );
  XNOR2_X1 U13577 ( .A(n11295), .B(n11292), .ZN(n11022) );
  OR2_X1 U13578 ( .A1(n11018), .A2(n11028), .ZN(n11020) );
  OAI21_X1 U13579 ( .B1(n11022), .B2(n11021), .A(n11293), .ZN(n11023) );
  NAND2_X1 U13580 ( .A1(n15052), .A2(n11023), .ZN(n11025) );
  AND2_X1 U13581 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11210) );
  INV_X1 U13582 ( .A(n11210), .ZN(n11024) );
  OAI211_X1 U13583 ( .C1(n15066), .C2(n11026), .A(n11025), .B(n11024), .ZN(
        n11032) );
  INV_X1 U13584 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11239) );
  AOI21_X1 U13585 ( .B1(n11239), .B2(n11029), .A(n6517), .ZN(n11030) );
  NOR2_X1 U13586 ( .A1(n11030), .A2(n15056), .ZN(n11031) );
  AOI211_X1 U13587 ( .C1(n15054), .C2(n11292), .A(n11032), .B(n11031), .ZN(
        n11033) );
  OAI21_X1 U13588 ( .B1(n11034), .B2(n15060), .A(n11033), .ZN(P3_U3189) );
  NAND2_X1 U13589 ( .A1(n11036), .A2(n11035), .ZN(n12358) );
  INV_X2 U13590 ( .A(n14630), .ZN(n14279) );
  INV_X1 U13591 ( .A(n11037), .ZN(n11038) );
  NAND2_X1 U13592 ( .A1(n14279), .A2(n11038), .ZN(n14171) );
  INV_X1 U13593 ( .A(n12358), .ZN(n11039) );
  NAND2_X1 U13594 ( .A1(n11039), .A2(n14112), .ZN(n11040) );
  XOR2_X1 U13595 ( .A(n11048), .B(n11041), .Z(n14795) );
  NOR2_X2 U13596 ( .A1(n12358), .A2(n11043), .ZN(n14604) );
  AOI21_X1 U13597 ( .B1(n11045), .B2(n11053), .A(n11044), .ZN(n11050) );
  INV_X1 U13598 ( .A(n11050), .ZN(n11046) );
  NOR2_X1 U13599 ( .A1(n11046), .A2(n14822), .ZN(n14800) );
  INV_X1 U13600 ( .A(n14611), .ZN(n14599) );
  AOI22_X1 U13601 ( .A1(n14604), .A2(n14800), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n14599), .ZN(n11047) );
  OAI21_X1 U13602 ( .B1(n10153), .B2(n14279), .A(n11047), .ZN(n11052) );
  NAND2_X1 U13603 ( .A1(n14279), .A2(n14255), .ZN(n14303) );
  AOI21_X1 U13604 ( .B1(n11048), .B2(n14041), .A(n14831), .ZN(n11049) );
  NOR2_X1 U13605 ( .A1(n11049), .A2(n14619), .ZN(n14799) );
  XNOR2_X1 U13606 ( .A(n11050), .B(n14040), .ZN(n14798) );
  NOR3_X1 U13607 ( .A1(n14303), .A2(n14799), .A3(n14798), .ZN(n11051) );
  AOI211_X1 U13608 ( .C1(n14601), .C2(n11053), .A(n11052), .B(n11051), .ZN(
        n11056) );
  OAI22_X1 U13609 ( .A1(n14799), .A2(n11054), .B1(n10724), .B2(n14274), .ZN(
        n14804) );
  NAND2_X1 U13610 ( .A1(n14804), .A2(n14279), .ZN(n11055) );
  OAI211_X1 U13611 ( .C1(n14286), .C2(n14795), .A(n11056), .B(n11055), .ZN(
        P1_U3292) );
  NAND2_X1 U13612 ( .A1(n12703), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n11057) );
  OAI21_X1 U13613 ( .B1(n12498), .B2(n12703), .A(n11057), .ZN(P3_U3521) );
  MUX2_X1 U13614 ( .A(n11059), .B(n11058), .S(n14952), .Z(n11064) );
  OAI22_X1 U13615 ( .A1(n13640), .A2(n7105), .B1(n14950), .B2(n11060), .ZN(
        n11061) );
  AOI21_X1 U13616 ( .B1(n11062), .B2(n13649), .A(n11061), .ZN(n11063) );
  OAI211_X1 U13617 ( .C1(n11065), .C2(n13609), .A(n11064), .B(n11063), .ZN(
        P2_U3260) );
  INV_X1 U13618 ( .A(n11066), .ZN(n11067) );
  OAI222_X1 U13619 ( .A1(n13175), .A2(n11067), .B1(n13178), .B2(n15362), .C1(
        P3_U3151), .C2(n12529), .ZN(P3_U3274) );
  OR2_X1 U13620 ( .A1(n11071), .A2(n13308), .ZN(n11068) );
  NAND2_X1 U13621 ( .A1(n11069), .A2(n11068), .ZN(n11151) );
  XNOR2_X1 U13622 ( .A(n11151), .B(n11149), .ZN(n14995) );
  NAND2_X1 U13623 ( .A1(n11071), .A2(n11070), .ZN(n11072) );
  OAI21_X1 U13624 ( .B1(n11074), .B2(n11149), .A(n11158), .ZN(n11075) );
  NAND2_X1 U13625 ( .A1(n11075), .A2(n13631), .ZN(n11077) );
  AOI22_X1 U13626 ( .A1(n15413), .A2(n13306), .B1(n13308), .B2(n13576), .ZN(
        n11076) );
  AND2_X1 U13627 ( .A1(n11077), .A2(n11076), .ZN(n14998) );
  MUX2_X1 U13628 ( .A(n11078), .B(n14998), .S(n14952), .Z(n11087) );
  NAND2_X1 U13629 ( .A1(n11079), .A2(n14991), .ZN(n11081) );
  NAND2_X1 U13630 ( .A1(n11081), .A2(n11674), .ZN(n11082) );
  NOR2_X1 U13631 ( .A1(n11162), .A2(n11082), .ZN(n14993) );
  OAI22_X1 U13632 ( .A1(n13640), .A2(n11084), .B1(n14950), .B2(n11083), .ZN(
        n11085) );
  AOI21_X1 U13633 ( .B1(n13649), .B2(n14993), .A(n11085), .ZN(n11086) );
  OAI211_X1 U13634 ( .C1(n13646), .C2(n14995), .A(n11087), .B(n11086), .ZN(
        P2_U3259) );
  INV_X1 U13635 ( .A(n11316), .ZN(n11097) );
  AOI21_X1 U13636 ( .B1(n11088), .B2(n11089), .A(n12462), .ZN(n11091) );
  NAND2_X1 U13637 ( .A1(n11091), .A2(n11090), .ZN(n11096) );
  OAI22_X1 U13638 ( .A1(n12441), .A2(n11092), .B1(n15147), .B2(n12477), .ZN(
        n11093) );
  AOI211_X1 U13639 ( .C1(n12439), .C2(n12710), .A(n11094), .B(n11093), .ZN(
        n11095) );
  OAI211_X1 U13640 ( .C1(n11097), .C2(n12034), .A(n11096), .B(n11095), .ZN(
        P3_U3179) );
  INV_X1 U13641 ( .A(n15204), .ZN(n14018) );
  INV_X1 U13642 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n15357) );
  INV_X1 U13643 ( .A(n14725), .ZN(n14705) );
  NAND2_X1 U13644 ( .A1(n14705), .A2(n14038), .ZN(n11102) );
  NAND2_X1 U13645 ( .A1(n15197), .A2(n11119), .ZN(n11101) );
  NAND2_X1 U13646 ( .A1(n14703), .A2(n14036), .ZN(n11100) );
  NAND2_X1 U13647 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n11099) );
  NAND4_X1 U13648 ( .A1(n11102), .A2(n11101), .A3(n11100), .A4(n11099), .ZN(
        n11115) );
  AOI22_X1 U13649 ( .A1(n14037), .A2(n13906), .B1(n11103), .B2(n11119), .ZN(
        n11189) );
  NAND2_X1 U13650 ( .A1(n14037), .A2(n11103), .ZN(n11105) );
  NAND2_X1 U13651 ( .A1(n11119), .A2(n13902), .ZN(n11104) );
  NAND2_X1 U13652 ( .A1(n11105), .A2(n11104), .ZN(n11106) );
  XNOR2_X1 U13653 ( .A(n11106), .B(n10601), .ZN(n11188) );
  XOR2_X1 U13654 ( .A(n11189), .B(n11188), .Z(n11113) );
  INV_X1 U13655 ( .A(n11107), .ZN(n11109) );
  NAND2_X1 U13656 ( .A1(n11109), .A2(n10802), .ZN(n11110) );
  AOI211_X1 U13657 ( .C1(n11113), .C2(n11112), .A(n14731), .B(n11192), .ZN(
        n11114) );
  AOI211_X1 U13658 ( .C1(n14018), .C2(n15357), .A(n11115), .B(n11114), .ZN(
        n11116) );
  INV_X1 U13659 ( .A(n11116), .ZN(P1_U3218) );
  XNOR2_X1 U13660 ( .A(n11132), .B(n11131), .ZN(n14811) );
  NAND2_X1 U13661 ( .A1(n11200), .A2(n11119), .ZN(n11120) );
  NAND2_X1 U13662 ( .A1(n11122), .A2(n11121), .ZN(n11123) );
  NAND3_X1 U13663 ( .A1(n11134), .A2(n14255), .A3(n11123), .ZN(n11125) );
  AOI22_X1 U13664 ( .A1(n14619), .A2(n14037), .B1(n14035), .B2(n14620), .ZN(
        n11124) );
  NAND2_X1 U13665 ( .A1(n11125), .A2(n11124), .ZN(n14807) );
  MUX2_X1 U13666 ( .A(n14807), .B(P1_REG2_REG_4__SCAN_IN), .S(n14630), .Z(
        n11126) );
  INV_X1 U13667 ( .A(n11126), .ZN(n11130) );
  AOI211_X1 U13668 ( .C1(n14809), .C2(n11127), .A(n14822), .B(n11138), .ZN(
        n14808) );
  OAI22_X1 U13669 ( .A1(n14307), .A2(n11193), .B1(n11197), .B2(n14611), .ZN(
        n11128) );
  AOI21_X1 U13670 ( .B1(n14808), .B2(n14604), .A(n11128), .ZN(n11129) );
  OAI211_X1 U13671 ( .C1(n14286), .C2(n14811), .A(n11130), .B(n11129), .ZN(
        P1_U3289) );
  XNOR2_X1 U13672 ( .A(n11323), .B(n11135), .ZN(n14818) );
  NAND2_X1 U13673 ( .A1(n14036), .A2(n11193), .ZN(n11133) );
  XNOR2_X1 U13674 ( .A(n11321), .B(n11135), .ZN(n11136) );
  AOI222_X1 U13675 ( .A1(n14614), .A2(n11136), .B1(n14034), .B2(n14620), .C1(
        n14036), .C2(n14619), .ZN(n14817) );
  MUX2_X1 U13676 ( .A(n11137), .B(n14817), .S(n14279), .Z(n11145) );
  INV_X1 U13677 ( .A(n11138), .ZN(n11140) );
  INV_X1 U13678 ( .A(n14813), .ZN(n11448) );
  INV_X1 U13679 ( .A(n11324), .ZN(n11139) );
  AOI21_X1 U13680 ( .B1(n14813), .B2(n11140), .A(n11139), .ZN(n14815) );
  NOR2_X1 U13681 ( .A1(n14630), .A2(n11141), .ZN(n14186) );
  INV_X1 U13682 ( .A(n11440), .ZN(n11142) );
  OAI22_X1 U13683 ( .A1(n14307), .A2(n11448), .B1(n14611), .B2(n11142), .ZN(
        n11143) );
  AOI21_X1 U13684 ( .B1(n14815), .B2(n14186), .A(n11143), .ZN(n11144) );
  OAI211_X1 U13685 ( .C1(n14286), .C2(n14818), .A(n11145), .B(n11144), .ZN(
        P1_U3288) );
  INV_X1 U13686 ( .A(n11146), .ZN(n11148) );
  OAI22_X1 U13687 ( .A1(n12695), .A2(P3_U3151), .B1(SI_22_), .B2(n12293), .ZN(
        n11147) );
  AOI21_X1 U13688 ( .B1(n11148), .B2(n11271), .A(n11147), .ZN(P3_U3273) );
  INV_X1 U13689 ( .A(n11149), .ZN(n11150) );
  NAND2_X1 U13690 ( .A1(n11151), .A2(n11150), .ZN(n11153) );
  OR2_X1 U13691 ( .A1(n14991), .A2(n13307), .ZN(n11152) );
  NAND2_X1 U13692 ( .A1(n11153), .A2(n11152), .ZN(n11155) );
  INV_X1 U13693 ( .A(n11159), .ZN(n11154) );
  NAND2_X1 U13694 ( .A1(n11155), .A2(n11154), .ZN(n11244) );
  OAI21_X1 U13695 ( .B1(n11155), .B2(n11154), .A(n11244), .ZN(n14961) );
  INV_X1 U13696 ( .A(n14961), .ZN(n11163) );
  NAND2_X1 U13697 ( .A1(n14991), .A2(n11156), .ZN(n11157) );
  XNOR2_X1 U13698 ( .A(n11246), .B(n11159), .ZN(n11161) );
  AOI21_X1 U13699 ( .B1(n11161), .B2(n13631), .A(n11160), .ZN(n14963) );
  INV_X1 U13700 ( .A(n11254), .ZN(n11256) );
  OAI211_X1 U13701 ( .C1(n11166), .C2(n11162), .A(n11256), .B(n11674), .ZN(
        n14957) );
  OAI211_X1 U13702 ( .C1(n11163), .C2(n14994), .A(n14963), .B(n14957), .ZN(
        n11168) );
  OAI22_X1 U13703 ( .A1(n11166), .A2(n13778), .B1(n15018), .B2(n7831), .ZN(
        n11164) );
  AOI21_X1 U13704 ( .B1(n11168), .B2(n15018), .A(n11164), .ZN(n11165) );
  INV_X1 U13705 ( .A(n11165), .ZN(P2_U3451) );
  OAI22_X1 U13706 ( .A1(n13736), .A2(n11166), .B1(n15027), .B2(n10090), .ZN(
        n11167) );
  AOI21_X1 U13707 ( .B1(n11168), .B2(n15027), .A(n11167), .ZN(n11169) );
  INV_X1 U13708 ( .A(n11169), .ZN(P2_U3506) );
  INV_X1 U13709 ( .A(n11170), .ZN(n11172) );
  OAI222_X1 U13710 ( .A1(n14474), .A2(n11171), .B1(n14464), .B2(n11172), .C1(
        n14079), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U13711 ( .A(n14924), .ZN(n11717) );
  OAI222_X1 U13712 ( .A1(n13807), .A2(n11173), .B1(n13805), .B2(n11172), .C1(
        n11717), .C2(P2_U3088), .ZN(P2_U3311) );
  NAND2_X1 U13713 ( .A1(n14388), .A2(n14828), .ZN(n14409) );
  OAI22_X1 U13714 ( .A1(n14409), .A2(n11339), .B1(n14388), .B2(n10188), .ZN(
        n11174) );
  AOI21_X1 U13715 ( .B1(n11175), .B2(n14388), .A(n11174), .ZN(n11176) );
  INV_X1 U13716 ( .A(n11176), .ZN(P1_U3530) );
  INV_X1 U13717 ( .A(n13646), .ZN(n14960) );
  OAI22_X1 U13718 ( .A1(n11178), .A2(n13640), .B1(n14958), .B2(n11177), .ZN(
        n11182) );
  OAI21_X1 U13719 ( .B1(n14950), .B2(P2_REG3_REG_3__SCAN_IN), .A(n11179), .ZN(
        n11180) );
  MUX2_X1 U13720 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11180), .S(n14952), .Z(
        n11181) );
  AOI211_X1 U13721 ( .C1(n14960), .C2(n11183), .A(n11182), .B(n11181), .ZN(
        n11184) );
  INV_X1 U13722 ( .A(n11184), .ZN(P2_U3262) );
  OAI22_X1 U13723 ( .A1(n14409), .A2(n14306), .B1(n14388), .B2(n10187), .ZN(
        n11185) );
  AOI21_X1 U13724 ( .B1(n11186), .B2(n14388), .A(n11185), .ZN(n11187) );
  INV_X1 U13725 ( .A(n11187), .ZN(P1_U3531) );
  INV_X1 U13726 ( .A(n11188), .ZN(n11190) );
  OAI22_X1 U13727 ( .A1(n11194), .A2(n10801), .B1(n11193), .B2(n13938), .ZN(
        n11191) );
  NAND2_X1 U13728 ( .A1(n6631), .A2(n11445), .ZN(n11196) );
  OAI22_X1 U13729 ( .A1(n11194), .A2(n13938), .B1(n11193), .B2(n13936), .ZN(
        n11195) );
  XOR2_X1 U13730 ( .A(n13940), .B(n11195), .Z(n11446) );
  XNOR2_X1 U13731 ( .A(n11196), .B(n11446), .ZN(n11204) );
  NOR2_X1 U13732 ( .A1(n15204), .A2(n11197), .ZN(n11202) );
  NAND2_X1 U13733 ( .A1(n14703), .A2(n14035), .ZN(n11199) );
  OAI211_X1 U13734 ( .C1(n11200), .C2(n14725), .A(n11199), .B(n11198), .ZN(
        n11201) );
  AOI211_X1 U13735 ( .C1(n14809), .C2(n15197), .A(n11202), .B(n11201), .ZN(
        n11203) );
  OAI21_X1 U13736 ( .B1(n11204), .B2(n14731), .A(n11203), .ZN(P1_U3230) );
  INV_X1 U13737 ( .A(n11237), .ZN(n11213) );
  OAI211_X1 U13738 ( .C1(n11207), .C2(n11206), .A(n11205), .B(n12468), .ZN(
        n11212) );
  INV_X1 U13739 ( .A(n11236), .ZN(n12565) );
  OAI22_X1 U13740 ( .A1(n12441), .A2(n11208), .B1(n12565), .B2(n12477), .ZN(
        n11209) );
  AOI211_X1 U13741 ( .C1(n12439), .C2(n12709), .A(n11210), .B(n11209), .ZN(
        n11211) );
  OAI211_X1 U13742 ( .C1(n11213), .C2(n12034), .A(n11212), .B(n11211), .ZN(
        P3_U3153) );
  OAI22_X1 U13743 ( .A1(n11214), .A2(n13269), .B1(n11401), .B2(n8233), .ZN(
        n11226) );
  INV_X1 U13744 ( .A(n14859), .ZN(n13238) );
  NAND2_X1 U13745 ( .A1(n13306), .A2(n13576), .ZN(n11216) );
  NAND2_X1 U13746 ( .A1(n13304), .A2(n15413), .ZN(n11215) );
  NAND2_X1 U13747 ( .A1(n11216), .A2(n11215), .ZN(n11251) );
  AND2_X1 U13748 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n13351) );
  AOI21_X1 U13749 ( .B1(n13238), .B2(n11251), .A(n13351), .ZN(n11218) );
  NAND2_X1 U13750 ( .A1(n11437), .A2(n14867), .ZN(n11217) );
  OAI211_X1 U13751 ( .C1(n14870), .C2(n11257), .A(n11218), .B(n11217), .ZN(
        n11225) );
  INV_X1 U13752 ( .A(n11219), .ZN(n11223) );
  INV_X1 U13753 ( .A(n11220), .ZN(n11221) );
  AOI211_X1 U13754 ( .C1(n11223), .C2(n11222), .A(n13269), .B(n11221), .ZN(
        n11224) );
  AOI211_X1 U13755 ( .C1(n11227), .C2(n11226), .A(n11225), .B(n11224), .ZN(
        n11228) );
  INV_X1 U13756 ( .A(n11228), .ZN(P2_U3193) );
  XNOR2_X1 U13757 ( .A(n11231), .B(n11229), .ZN(n11235) );
  OAI211_X1 U13758 ( .C1(n11232), .C2(n11231), .A(n11230), .B(n15112), .ZN(
        n11234) );
  AOI22_X1 U13759 ( .A1(n15109), .A2(n15073), .B1(n12709), .B2(n15106), .ZN(
        n11233) );
  OAI211_X1 U13760 ( .C1(n15116), .C2(n11235), .A(n11234), .B(n11233), .ZN(
        n15153) );
  INV_X1 U13761 ( .A(n15153), .ZN(n11242) );
  INV_X1 U13762 ( .A(n11235), .ZN(n15155) );
  AND2_X1 U13763 ( .A1(n11236), .A2(n15080), .ZN(n15154) );
  AOI22_X1 U13764 ( .A1(n15083), .A2(n15154), .B1(n15119), .B2(n11237), .ZN(
        n11238) );
  OAI21_X1 U13765 ( .B1(n11239), .B2(n15122), .A(n11238), .ZN(n11240) );
  AOI21_X1 U13766 ( .B1(n15155), .B2(n15120), .A(n11240), .ZN(n11241) );
  OAI21_X1 U13767 ( .B1(n11242), .B2(n15124), .A(n11241), .ZN(P3_U3226) );
  OR2_X1 U13768 ( .A1(n14954), .A2(n13306), .ZN(n11243) );
  OAI21_X1 U13769 ( .B1(n7566), .B2(n11249), .A(n11393), .ZN(n11429) );
  INV_X1 U13770 ( .A(n13306), .ZN(n11247) );
  OR2_X1 U13771 ( .A1(n14954), .A2(n11247), .ZN(n11245) );
  NAND2_X1 U13772 ( .A1(n14954), .A2(n11247), .ZN(n11248) );
  AOI21_X1 U13773 ( .B1(n11250), .B2(n11249), .A(n13562), .ZN(n11252) );
  AOI21_X1 U13774 ( .B1(n11252), .B2(n11402), .A(n11251), .ZN(n11430) );
  MUX2_X1 U13775 ( .A(n11253), .B(n11430), .S(n14952), .Z(n11260) );
  INV_X1 U13776 ( .A(n11437), .ZN(n11434) );
  INV_X1 U13777 ( .A(n11395), .ZN(n11255) );
  AOI211_X1 U13778 ( .C1(n11437), .C2(n11256), .A(n11080), .B(n11255), .ZN(
        n11432) );
  OAI22_X1 U13779 ( .A1(n11434), .A2(n13640), .B1(n14950), .B2(n11257), .ZN(
        n11258) );
  AOI21_X1 U13780 ( .B1(n11432), .B2(n13649), .A(n11258), .ZN(n11259) );
  OAI211_X1 U13781 ( .C1(n13646), .C2(n11429), .A(n11260), .B(n11259), .ZN(
        P2_U3257) );
  INV_X1 U13782 ( .A(n11261), .ZN(n11262) );
  AOI21_X1 U13783 ( .B1(n11263), .B2(n6756), .A(n11262), .ZN(n11270) );
  NAND2_X1 U13784 ( .A1(n13305), .A2(n13576), .ZN(n11265) );
  NAND2_X1 U13785 ( .A1(n13303), .A2(n15413), .ZN(n11264) );
  AND2_X1 U13786 ( .A1(n11265), .A2(n11264), .ZN(n11404) );
  OAI22_X1 U13787 ( .A1(n14859), .A2(n11404), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11266), .ZN(n11268) );
  NOR2_X1 U13788 ( .A1(n14870), .A2(n11397), .ZN(n11267) );
  AOI211_X1 U13789 ( .C1(n11554), .C2(n14867), .A(n11268), .B(n11267), .ZN(
        n11269) );
  OAI21_X1 U13790 ( .B1(n11270), .B2(n13269), .A(n11269), .ZN(P2_U3203) );
  NAND2_X1 U13791 ( .A1(n11272), .A2(n11271), .ZN(n11273) );
  OAI211_X1 U13792 ( .C1(n7405), .C2(n12293), .A(n11273), .B(n12697), .ZN(
        P3_U3272) );
  NOR2_X1 U13793 ( .A1(n11292), .A2(n11274), .ZN(n11276) );
  NAND2_X1 U13794 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n11286), .ZN(n11277) );
  OAI21_X1 U13795 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n11286), .A(n11277), .ZN(
        n15039) );
  NOR2_X1 U13796 ( .A1(n15053), .A2(n11278), .ZN(n11279) );
  INV_X1 U13797 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15188) );
  NAND2_X1 U13798 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11842), .ZN(n11280) );
  OAI21_X1 U13799 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(n11842), .A(n11280), 
        .ZN(n11281) );
  AOI21_X1 U13800 ( .B1(n11282), .B2(n11281), .A(n11841), .ZN(n11306) );
  NOR2_X1 U13801 ( .A1(n11292), .A2(n11283), .ZN(n11284) );
  NAND2_X1 U13802 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n11286), .ZN(n11285) );
  OAI21_X1 U13803 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n11286), .A(n11285), .ZN(
        n15030) );
  NOR2_X1 U13804 ( .A1(n15053), .A2(n6601), .ZN(n11287) );
  INV_X1 U13805 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15048) );
  NOR2_X1 U13806 ( .A1(n11287), .A2(n15046), .ZN(n11291) );
  NAND2_X1 U13807 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n11842), .ZN(n11288) );
  OAI21_X1 U13808 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11842), .A(n11288), 
        .ZN(n11290) );
  OAI221_X1 U13809 ( .B1(n11830), .B2(n11291), .C1(n11830), .C2(n11290), .A(
        n11289), .ZN(n11305) );
  MUX2_X1 U13810 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12824), .Z(n11296) );
  XNOR2_X1 U13811 ( .A(n11296), .B(n15035), .ZN(n15033) );
  INV_X1 U13812 ( .A(n11292), .ZN(n11294) );
  OAI21_X1 U13813 ( .B1(n11295), .B2(n11294), .A(n11293), .ZN(n15032) );
  INV_X1 U13814 ( .A(n11296), .ZN(n11297) );
  MUX2_X1 U13815 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n12824), .Z(n11298) );
  XOR2_X1 U13816 ( .A(n15053), .B(n11298), .Z(n15049) );
  OAI22_X1 U13817 ( .A1(n15050), .A2(n15049), .B1(n11298), .B2(n6905), .ZN(
        n11300) );
  MUX2_X1 U13818 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12824), .Z(n11832) );
  XOR2_X1 U13819 ( .A(n11832), .B(n11842), .Z(n11299) );
  NAND2_X1 U13820 ( .A1(n11300), .A2(n11299), .ZN(n11833) );
  OAI21_X1 U13821 ( .B1(n11300), .B2(n11299), .A(n11833), .ZN(n11303) );
  INV_X1 U13822 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14495) );
  NAND2_X1 U13823 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n11654)
         );
  OAI21_X1 U13824 ( .B1(n15066), .B2(n14495), .A(n11654), .ZN(n11302) );
  NOR2_X1 U13825 ( .A1(n12860), .A2(n11842), .ZN(n11301) );
  AOI211_X1 U13826 ( .C1(n15052), .C2(n11303), .A(n11302), .B(n11301), .ZN(
        n11304) );
  OAI211_X1 U13827 ( .C1(n11306), .C2(n15060), .A(n11305), .B(n11304), .ZN(
        P3_U3192) );
  XNOR2_X1 U13828 ( .A(n11307), .B(n12504), .ZN(n11311) );
  INV_X1 U13829 ( .A(n11311), .ZN(n15149) );
  OAI211_X1 U13830 ( .C1(n11310), .C2(n11309), .A(n11308), .B(n15112), .ZN(
        n11314) );
  AOI22_X1 U13831 ( .A1(n15109), .A2(n12711), .B1(n12710), .B2(n15106), .ZN(
        n11313) );
  NAND2_X1 U13832 ( .A1(n11311), .A2(n15075), .ZN(n11312) );
  NAND3_X1 U13833 ( .A1(n11314), .A2(n11313), .A3(n11312), .ZN(n15151) );
  MUX2_X1 U13834 ( .A(n15151), .B(P3_REG2_REG_6__SCAN_IN), .S(n15124), .Z(
        n11315) );
  INV_X1 U13835 ( .A(n11315), .ZN(n11319) );
  AOI22_X1 U13836 ( .A1(n13027), .A2(n11317), .B1(n15119), .B2(n11316), .ZN(
        n11318) );
  OAI211_X1 U13837 ( .C1(n15149), .C2(n12944), .A(n11319), .B(n11318), .ZN(
        P3_U3227) );
  OR2_X1 U13838 ( .A1(n14035), .A2(n14813), .ZN(n11322) );
  XNOR2_X1 U13839 ( .A(n11375), .B(n11374), .ZN(n11426) );
  AOI21_X1 U13840 ( .B1(n11324), .B2(n11617), .A(n14822), .ZN(n11325) );
  OR2_X1 U13841 ( .A1(n11324), .A2(n11617), .ZN(n11532) );
  AND2_X1 U13842 ( .A1(n11325), .A2(n11532), .ZN(n11421) );
  NAND2_X1 U13843 ( .A1(n14035), .A2(n14619), .ZN(n11327) );
  NAND2_X1 U13844 ( .A1(n14033), .A2(n14620), .ZN(n11326) );
  NAND2_X1 U13845 ( .A1(n11327), .A2(n11326), .ZN(n11608) );
  AOI211_X1 U13846 ( .C1(n11426), .C2(n14842), .A(n11421), .B(n11608), .ZN(
        n11328) );
  OAI21_X1 U13847 ( .B1(n14831), .B2(n11428), .A(n11328), .ZN(n11334) );
  INV_X1 U13848 ( .A(n11617), .ZN(n11424) );
  OAI22_X1 U13849 ( .A1(n14409), .A2(n11424), .B1(n14388), .B2(n11329), .ZN(
        n11330) );
  AOI21_X1 U13850 ( .B1(n11334), .B2(n14388), .A(n11330), .ZN(n11331) );
  INV_X1 U13851 ( .A(n11331), .ZN(P1_U3534) );
  INV_X1 U13852 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n11332) );
  OAI22_X1 U13853 ( .A1(n14446), .A2(n11424), .B1(n14845), .B2(n11332), .ZN(
        n11333) );
  AOI21_X1 U13854 ( .B1(n11334), .B2(n14845), .A(n11333), .ZN(n11335) );
  INV_X1 U13855 ( .A(n11335), .ZN(P1_U3477) );
  INV_X1 U13856 ( .A(n14303), .ZN(n14283) );
  MUX2_X1 U13857 ( .A(n11336), .B(P1_REG2_REG_2__SCAN_IN), .S(n14630), .Z(
        n11341) );
  AOI22_X1 U13858 ( .A1(n11337), .A2(n14604), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n14599), .ZN(n11338) );
  OAI21_X1 U13859 ( .B1(n11339), .B2(n14307), .A(n11338), .ZN(n11340) );
  AOI211_X1 U13860 ( .C1(n14283), .C2(n11342), .A(n11341), .B(n11340), .ZN(
        n11343) );
  OAI21_X1 U13861 ( .B1(n14286), .B2(n11344), .A(n11343), .ZN(P1_U3291) );
  INV_X1 U13862 ( .A(n11345), .ZN(n11347) );
  OAI222_X1 U13863 ( .A1(n14474), .A2(n11346), .B1(n14464), .B2(n11347), .C1(
        n11729), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U13864 ( .A(n14937), .ZN(n11719) );
  OAI222_X1 U13865 ( .A1(n13807), .A2(n11348), .B1(n13805), .B2(n11347), .C1(
        n11719), .C2(P2_U3088), .ZN(P2_U3310) );
  NOR2_X1 U13866 ( .A1(n14631), .A2(n14283), .ZN(n11355) );
  OAI22_X1 U13867 ( .A1(n14630), .A2(n11350), .B1(n11349), .B2(n14611), .ZN(
        n11353) );
  INV_X1 U13868 ( .A(n14186), .ZN(n12100) );
  AOI21_X1 U13869 ( .B1(n12100), .B2(n14307), .A(n11351), .ZN(n11352) );
  AOI211_X1 U13870 ( .C1(n14630), .C2(P1_REG2_REG_0__SCAN_IN), .A(n11353), .B(
        n11352), .ZN(n11354) );
  OAI21_X1 U13871 ( .B1(n11356), .B2(n11355), .A(n11354), .ZN(P1_U3293) );
  INV_X1 U13872 ( .A(n11576), .ZN(n11366) );
  OAI211_X1 U13873 ( .C1(n11359), .C2(n11358), .A(n11357), .B(n12468), .ZN(
        n11365) );
  NAND2_X1 U13874 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n15043) );
  INV_X1 U13875 ( .A(n15043), .ZN(n11363) );
  OAI22_X1 U13876 ( .A1(n12441), .A2(n11361), .B1(n11360), .B2(n12477), .ZN(
        n11362) );
  AOI211_X1 U13877 ( .C1(n12439), .C2(n12708), .A(n11363), .B(n11362), .ZN(
        n11364) );
  OAI211_X1 U13878 ( .C1(n12034), .C2(n11366), .A(n11365), .B(n11364), .ZN(
        P3_U3161) );
  INV_X1 U13879 ( .A(n14034), .ZN(n11367) );
  AND2_X1 U13880 ( .A1(n11617), .A2(n11367), .ZN(n11368) );
  NAND2_X1 U13881 ( .A1(n11540), .A2(n11539), .ZN(n11538) );
  INV_X1 U13882 ( .A(n14033), .ZN(n11370) );
  OR2_X1 U13883 ( .A1(n11536), .A2(n11370), .ZN(n11371) );
  INV_X1 U13884 ( .A(n11380), .ZN(n11372) );
  OAI21_X1 U13885 ( .B1(n11373), .B2(n11372), .A(n11594), .ZN(n14832) );
  OR2_X1 U13886 ( .A1(n11617), .A2(n14034), .ZN(n11376) );
  INV_X1 U13887 ( .A(n11539), .ZN(n11378) );
  OR2_X1 U13888 ( .A1(n11536), .A2(n14033), .ZN(n11379) );
  XNOR2_X1 U13889 ( .A(n11582), .B(n11380), .ZN(n14834) );
  NAND2_X1 U13890 ( .A1(n14834), .A2(n14631), .ZN(n11391) );
  NAND2_X1 U13891 ( .A1(n14031), .A2(n14620), .ZN(n11382) );
  NAND2_X1 U13892 ( .A1(n14033), .A2(n14619), .ZN(n11381) );
  NAND2_X1 U13893 ( .A1(n11382), .A2(n11381), .ZN(n15199) );
  INV_X1 U13894 ( .A(n15199), .ZN(n11384) );
  MUX2_X1 U13895 ( .A(n11384), .B(n11383), .S(n14630), .Z(n11385) );
  OAI21_X1 U13896 ( .B1(n14611), .B2(n15203), .A(n11385), .ZN(n11389) );
  OR2_X1 U13897 ( .A1(n11532), .A2(n11536), .ZN(n11533) );
  NAND2_X1 U13898 ( .A1(n11533), .A2(n15198), .ZN(n11386) );
  NAND2_X1 U13899 ( .A1(n11386), .A2(n14814), .ZN(n11387) );
  OR2_X1 U13900 ( .A1(n11387), .A2(n11589), .ZN(n14829) );
  NOR2_X1 U13901 ( .A1(n14829), .A2(n14300), .ZN(n11388) );
  AOI211_X1 U13902 ( .C1(n14601), .C2(n15198), .A(n11389), .B(n11388), .ZN(
        n11390) );
  OAI211_X1 U13903 ( .C1(n14832), .C2(n14303), .A(n11391), .B(n11390), .ZN(
        P1_U3285) );
  NAND2_X1 U13904 ( .A1(n11437), .A2(n13305), .ZN(n11392) );
  XNOR2_X1 U13905 ( .A(n11515), .B(n11513), .ZN(n11551) );
  INV_X1 U13906 ( .A(n11551), .ZN(n11408) );
  INV_X1 U13907 ( .A(n11522), .ZN(n11394) );
  AOI211_X1 U13908 ( .C1(n11554), .C2(n11395), .A(n11080), .B(n11394), .ZN(
        n11550) );
  INV_X1 U13909 ( .A(n11554), .ZN(n11396) );
  NOR2_X1 U13910 ( .A1(n11396), .A2(n13640), .ZN(n11400) );
  OAI22_X1 U13911 ( .A1(n14952), .A2(n11398), .B1(n11397), .B2(n14950), .ZN(
        n11399) );
  AOI211_X1 U13912 ( .C1(n11550), .C2(n13649), .A(n11400), .B(n11399), .ZN(
        n11407) );
  OAI211_X1 U13913 ( .C1(n11403), .C2(n11513), .A(n11518), .B(n13631), .ZN(
        n11405) );
  NAND2_X1 U13914 ( .A1(n11405), .A2(n11404), .ZN(n11549) );
  NAND2_X1 U13915 ( .A1(n11549), .A2(n14952), .ZN(n11406) );
  OAI211_X1 U13916 ( .C1(n11408), .C2(n13646), .A(n11407), .B(n11406), .ZN(
        P2_U3256) );
  INV_X1 U13917 ( .A(n11663), .ZN(n15003) );
  AOI21_X1 U13918 ( .B1(n11410), .B2(n11409), .A(n13269), .ZN(n11411) );
  NAND2_X1 U13919 ( .A1(n11411), .A2(n11500), .ZN(n11418) );
  INV_X1 U13920 ( .A(n11525), .ZN(n11416) );
  NAND2_X1 U13921 ( .A1(n13304), .A2(n13576), .ZN(n11413) );
  NAND2_X1 U13922 ( .A1(n13302), .A2(n15413), .ZN(n11412) );
  AND2_X1 U13923 ( .A1(n11413), .A2(n11412), .ZN(n11520) );
  INV_X1 U13924 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n11414) );
  OAI22_X1 U13925 ( .A1(n14859), .A2(n11520), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11414), .ZN(n11415) );
  AOI21_X1 U13926 ( .B1(n13277), .B2(n11416), .A(n11415), .ZN(n11417) );
  OAI211_X1 U13927 ( .C1(n15003), .C2(n13281), .A(n11418), .B(n11417), .ZN(
        P2_U3189) );
  INV_X1 U13928 ( .A(n11610), .ZN(n11420) );
  MUX2_X1 U13929 ( .A(n11608), .B(P1_REG2_REG_6__SCAN_IN), .S(n14630), .Z(
        n11419) );
  AOI21_X1 U13930 ( .B1(n14599), .B2(n11420), .A(n11419), .ZN(n11423) );
  NAND2_X1 U13931 ( .A1(n11421), .A2(n14604), .ZN(n11422) );
  OAI211_X1 U13932 ( .C1(n11424), .C2(n14307), .A(n11423), .B(n11422), .ZN(
        n11425) );
  AOI21_X1 U13933 ( .B1(n11426), .B2(n14631), .A(n11425), .ZN(n11427) );
  OAI21_X1 U13934 ( .B1(n11428), .B2(n14303), .A(n11427), .ZN(P1_U3287) );
  INV_X1 U13935 ( .A(n11429), .ZN(n11433) );
  INV_X1 U13936 ( .A(n11430), .ZN(n11431) );
  AOI211_X1 U13937 ( .C1(n11433), .C2(n15009), .A(n11432), .B(n11431), .ZN(
        n11439) );
  OAI22_X1 U13938 ( .A1(n11434), .A2(n13778), .B1(n15018), .B2(n7850), .ZN(
        n11435) );
  INV_X1 U13939 ( .A(n11435), .ZN(n11436) );
  OAI21_X1 U13940 ( .B1(n11439), .B2(n15017), .A(n11436), .ZN(P2_U3454) );
  AOI22_X1 U13941 ( .A1(n13745), .A2(n11437), .B1(n15025), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n11438) );
  OAI21_X1 U13942 ( .B1(n11439), .B2(n15025), .A(n11438), .ZN(P2_U3507) );
  NAND2_X1 U13943 ( .A1(n14705), .A2(n14036), .ZN(n11444) );
  NAND2_X1 U13944 ( .A1(n14018), .A2(n11440), .ZN(n11443) );
  NAND2_X1 U13945 ( .A1(n14703), .A2(n14034), .ZN(n11441) );
  NAND4_X1 U13946 ( .A1(n11444), .A2(n11443), .A3(n11442), .A4(n11441), .ZN(
        n11456) );
  OAI22_X1 U13947 ( .A1(n11448), .A2(n13936), .B1(n11447), .B2(n13938), .ZN(
        n11449) );
  XOR2_X1 U13948 ( .A(n13940), .B(n11449), .Z(n11451) );
  AOI22_X1 U13949 ( .A1(n14813), .A2(n11103), .B1(n13906), .B2(n14035), .ZN(
        n11450) );
  NOR2_X1 U13950 ( .A1(n11451), .A2(n11450), .ZN(n11459) );
  NAND2_X1 U13951 ( .A1(n11451), .A2(n11450), .ZN(n11458) );
  INV_X1 U13952 ( .A(n11458), .ZN(n11452) );
  NOR2_X1 U13953 ( .A1(n11459), .A2(n11452), .ZN(n11453) );
  XNOR2_X1 U13954 ( .A(n11460), .B(n11453), .ZN(n11454) );
  NOR2_X1 U13955 ( .A1(n11454), .A2(n14731), .ZN(n11455) );
  AOI211_X1 U13956 ( .C1(n14813), .C2(n15197), .A(n11456), .B(n11455), .ZN(
        n11457) );
  INV_X1 U13957 ( .A(n11457), .ZN(P1_U3227) );
  NAND2_X1 U13958 ( .A1(n11617), .A2(n13902), .ZN(n11462) );
  NAND2_X1 U13959 ( .A1(n14034), .A2(n11103), .ZN(n11461) );
  NAND2_X1 U13960 ( .A1(n11462), .A2(n11461), .ZN(n11463) );
  XNOR2_X1 U13961 ( .A(n11463), .B(n10601), .ZN(n11467) );
  NAND2_X1 U13962 ( .A1(n11617), .A2(n11103), .ZN(n11465) );
  NAND2_X1 U13963 ( .A1(n14034), .A2(n13906), .ZN(n11464) );
  NAND2_X1 U13964 ( .A1(n11465), .A2(n11464), .ZN(n11466) );
  NAND2_X1 U13965 ( .A1(n11467), .A2(n11466), .ZN(n11611) );
  AOI22_X1 U13966 ( .A1(n11536), .A2(n11103), .B1(n13906), .B2(n14033), .ZN(
        n11771) );
  AOI22_X1 U13967 ( .A1(n11536), .A2(n13902), .B1(n11103), .B2(n14033), .ZN(
        n11468) );
  XNOR2_X1 U13968 ( .A(n11468), .B(n10601), .ZN(n11772) );
  XOR2_X1 U13969 ( .A(n11771), .B(n11772), .Z(n11775) );
  XNOR2_X1 U13970 ( .A(n11776), .B(n11775), .ZN(n11475) );
  NAND2_X1 U13971 ( .A1(n14034), .A2(n14619), .ZN(n11470) );
  NAND2_X1 U13972 ( .A1(n14032), .A2(n14620), .ZN(n11469) );
  AND2_X1 U13973 ( .A1(n11470), .A2(n11469), .ZN(n11542) );
  OAI21_X1 U13974 ( .B1(n14015), .B2(n11542), .A(n11471), .ZN(n11472) );
  AOI21_X1 U13975 ( .B1(n14018), .B2(n11535), .A(n11472), .ZN(n11474) );
  NAND2_X1 U13976 ( .A1(n15197), .A2(n11536), .ZN(n11473) );
  OAI211_X1 U13977 ( .C1(n11475), .C2(n14731), .A(n11474), .B(n11473), .ZN(
        P1_U3213) );
  NAND2_X1 U13978 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3086), .ZN(n14736)
         );
  XNOR2_X1 U13979 ( .A(n11729), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n11482) );
  INV_X1 U13980 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11480) );
  XNOR2_X1 U13981 ( .A(n14079), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n14084) );
  OR2_X1 U13982 ( .A1(n11476), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11477) );
  NAND2_X1 U13983 ( .A1(n11478), .A2(n11477), .ZN(n11479) );
  XNOR2_X1 U13984 ( .A(n11479), .B(n11489), .ZN(n14778) );
  NOR2_X1 U13985 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14778), .ZN(n14777) );
  AOI21_X1 U13986 ( .B1(n11479), .B2(n11489), .A(n14777), .ZN(n14085) );
  NAND2_X1 U13987 ( .A1(n14084), .A2(n14085), .ZN(n14082) );
  OAI21_X1 U13988 ( .B1(n14079), .B2(n11480), .A(n14082), .ZN(n11481) );
  NAND2_X1 U13989 ( .A1(n11482), .A2(n11481), .ZN(n11728) );
  OAI211_X1 U13990 ( .C1(n11482), .C2(n11481), .A(n14083), .B(n11728), .ZN(
        n11483) );
  NAND2_X1 U13991 ( .A1(n14736), .A2(n11483), .ZN(n11497) );
  NOR2_X1 U13992 ( .A1(n11729), .A2(n14278), .ZN(n11484) );
  AOI21_X1 U13993 ( .B1(n14278), .B2(n11729), .A(n11484), .ZN(n11493) );
  NOR2_X1 U13994 ( .A1(n14079), .A2(n14295), .ZN(n11485) );
  AOI21_X1 U13995 ( .B1(n14295), .B2(n14079), .A(n11485), .ZN(n14076) );
  INV_X1 U13996 ( .A(n11486), .ZN(n11487) );
  OAI21_X1 U13997 ( .B1(n11488), .B2(n12097), .A(n11487), .ZN(n11490) );
  NOR2_X1 U13998 ( .A1(n14783), .A2(n11490), .ZN(n11491) );
  XOR2_X1 U13999 ( .A(n11490), .B(n11489), .Z(n14780) );
  NOR2_X1 U14000 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14780), .ZN(n14779) );
  NOR2_X1 U14001 ( .A1(n11491), .A2(n14779), .ZN(n14077) );
  NAND2_X1 U14002 ( .A1(n14076), .A2(n14077), .ZN(n14075) );
  OAI21_X1 U14003 ( .B1(n14079), .B2(n14295), .A(n14075), .ZN(n11492) );
  NAND2_X1 U14004 ( .A1(n11493), .A2(n11492), .ZN(n11726) );
  OAI211_X1 U14005 ( .C1(n11493), .C2(n11492), .A(n14074), .B(n11726), .ZN(
        n11495) );
  NAND2_X1 U14006 ( .A1(n14080), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n11494) );
  OAI211_X1 U14007 ( .C1(n11995), .C2(n11729), .A(n11495), .B(n11494), .ZN(
        n11496) );
  OR2_X1 U14008 ( .A1(n11497), .A2(n11496), .ZN(P1_U3260) );
  INV_X1 U14009 ( .A(n11816), .ZN(n15013) );
  INV_X1 U14010 ( .A(n11498), .ZN(n11499) );
  AOI21_X1 U14011 ( .B1(n11500), .B2(n11499), .A(n13269), .ZN(n11505) );
  INV_X1 U14012 ( .A(n13303), .ZN(n11501) );
  NOR3_X1 U14013 ( .A1(n11502), .A2(n11501), .A3(n8233), .ZN(n11504) );
  OAI21_X1 U14014 ( .B1(n11505), .B2(n11504), .A(n11503), .ZN(n11512) );
  INV_X1 U14015 ( .A(n11676), .ZN(n11510) );
  NAND2_X1 U14016 ( .A1(n13303), .A2(n13576), .ZN(n11507) );
  NAND2_X1 U14017 ( .A1(n13301), .A2(n15413), .ZN(n11506) );
  AND2_X1 U14018 ( .A1(n11507), .A2(n11506), .ZN(n11672) );
  OAI22_X1 U14019 ( .A1(n14859), .A2(n11672), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11508), .ZN(n11509) );
  AOI21_X1 U14020 ( .B1(n13277), .B2(n11510), .A(n11509), .ZN(n11511) );
  OAI211_X1 U14021 ( .C1(n15013), .C2(n13281), .A(n11512), .B(n11511), .ZN(
        P2_U3208) );
  INV_X1 U14022 ( .A(n11513), .ZN(n11514) );
  XNOR2_X1 U14023 ( .A(n11662), .B(n11660), .ZN(n15001) );
  INV_X1 U14024 ( .A(n15001), .ZN(n11530) );
  INV_X1 U14025 ( .A(n13304), .ZN(n11516) );
  OR2_X1 U14026 ( .A1(n11554), .A2(n11516), .ZN(n11517) );
  OAI211_X1 U14027 ( .C1(n11519), .C2(n11660), .A(n11667), .B(n13631), .ZN(
        n11521) );
  NAND2_X1 U14028 ( .A1(n11521), .A2(n11520), .ZN(n15005) );
  NOR2_X2 U14029 ( .A1(n11663), .A2(n11522), .ZN(n11675) );
  NAND2_X1 U14030 ( .A1(n11663), .A2(n11522), .ZN(n11523) );
  NAND2_X1 U14031 ( .A1(n11523), .A2(n11674), .ZN(n11524) );
  OR2_X1 U14032 ( .A1(n11675), .A2(n11524), .ZN(n15002) );
  INV_X1 U14033 ( .A(n13640), .ZN(n14955) );
  OAI22_X1 U14034 ( .A1(n14952), .A2(n10356), .B1(n11525), .B2(n14950), .ZN(
        n11526) );
  AOI21_X1 U14035 ( .B1(n11663), .B2(n14955), .A(n11526), .ZN(n11527) );
  OAI21_X1 U14036 ( .B1(n15002), .B2(n14958), .A(n11527), .ZN(n11528) );
  AOI21_X1 U14037 ( .B1(n15005), .B2(n14952), .A(n11528), .ZN(n11529) );
  OAI21_X1 U14038 ( .B1(n11530), .B2(n13646), .A(n11529), .ZN(P2_U3255) );
  XNOR2_X1 U14039 ( .A(n11531), .B(n11539), .ZN(n11543) );
  INV_X1 U14040 ( .A(n11543), .ZN(n14826) );
  INV_X1 U14041 ( .A(n14171), .ZN(n14605) );
  INV_X1 U14042 ( .A(n11532), .ZN(n11534) );
  INV_X1 U14043 ( .A(n11536), .ZN(n14821) );
  OAI21_X1 U14044 ( .B1(n11534), .B2(n14821), .A(n11533), .ZN(n14823) );
  AOI22_X1 U14045 ( .A1(n14601), .A2(n11536), .B1(n11535), .B2(n14599), .ZN(
        n11537) );
  OAI21_X1 U14046 ( .B1(n14823), .B2(n12100), .A(n11537), .ZN(n11545) );
  OAI211_X1 U14047 ( .C1(n11540), .C2(n11539), .A(n11538), .B(n14255), .ZN(
        n11541) );
  OAI211_X1 U14048 ( .C1(n11543), .C2(n14797), .A(n11542), .B(n11541), .ZN(
        n14824) );
  MUX2_X1 U14049 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n14824), .S(n14279), .Z(
        n11544) );
  AOI211_X1 U14050 ( .C1(n14826), .C2(n14605), .A(n11545), .B(n11544), .ZN(
        n11546) );
  INV_X1 U14051 ( .A(n11546), .ZN(P1_U3286) );
  INV_X1 U14052 ( .A(n11547), .ZN(n11580) );
  AOI22_X1 U14053 ( .A1(n11991), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n14450), .ZN(n11548) );
  OAI21_X1 U14054 ( .B1(n11580), .B2(n14472), .A(n11548), .ZN(P1_U3337) );
  AOI211_X1 U14055 ( .C1(n15009), .C2(n11551), .A(n11550), .B(n11549), .ZN(
        n11556) );
  INV_X1 U14056 ( .A(n13778), .ZN(n13783) );
  NOR2_X1 U14057 ( .A1(n15018), .A2(n7873), .ZN(n11552) );
  AOI21_X1 U14058 ( .B1(n11554), .B2(n13783), .A(n11552), .ZN(n11553) );
  OAI21_X1 U14059 ( .B1(n11556), .B2(n15017), .A(n11553), .ZN(P2_U3457) );
  AOI22_X1 U14060 ( .A1(n11554), .A2(n13745), .B1(n15025), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11555) );
  OAI21_X1 U14061 ( .B1(n11556), .B2(n15025), .A(n11555), .ZN(P2_U3508) );
  AOI21_X1 U14062 ( .B1(n11559), .B2(n11558), .A(n11557), .ZN(n11565) );
  NAND2_X1 U14063 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n15064) );
  INV_X1 U14064 ( .A(n15064), .ZN(n11562) );
  OAI22_X1 U14065 ( .A1(n12441), .A2(n11560), .B1(n11624), .B2(n12477), .ZN(
        n11561) );
  AOI211_X1 U14066 ( .C1(n12439), .C2(n12707), .A(n11562), .B(n11561), .ZN(
        n11564) );
  NAND2_X1 U14067 ( .A1(n12474), .A2(n11625), .ZN(n11563) );
  OAI211_X1 U14068 ( .C1(n11565), .C2(n12462), .A(n11564), .B(n11563), .ZN(
        P3_U3171) );
  INV_X1 U14069 ( .A(n12569), .ZN(n11566) );
  XNOR2_X1 U14070 ( .A(n11567), .B(n11566), .ZN(n15157) );
  NAND2_X1 U14071 ( .A1(n11568), .A2(n12569), .ZN(n11569) );
  NAND2_X1 U14072 ( .A1(n11570), .A2(n11569), .ZN(n11571) );
  NAND2_X1 U14073 ( .A1(n11571), .A2(n15112), .ZN(n11573) );
  AOI22_X1 U14074 ( .A1(n15109), .A2(n12710), .B1(n12708), .B2(n15106), .ZN(
        n11572) );
  OAI211_X1 U14075 ( .C1(n15116), .C2(n15157), .A(n11573), .B(n11572), .ZN(
        n15158) );
  MUX2_X1 U14076 ( .A(n15158), .B(P3_REG2_REG_8__SCAN_IN), .S(n15124), .Z(
        n11574) );
  INV_X1 U14077 ( .A(n11574), .ZN(n11578) );
  AND2_X1 U14078 ( .A1(n11575), .A2(n15080), .ZN(n15159) );
  AOI22_X1 U14079 ( .A1(n15083), .A2(n15159), .B1(n11576), .B2(n15119), .ZN(
        n11577) );
  OAI211_X1 U14080 ( .C1(n15157), .C2(n12944), .A(n11578), .B(n11577), .ZN(
        P3_U3225) );
  INV_X1 U14081 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11581) );
  INV_X1 U14082 ( .A(n12060), .ZN(n11579) );
  OAI222_X1 U14083 ( .A1(n13807), .A2(n11581), .B1(n13805), .B2(n11580), .C1(
        P2_U3088), .C2(n11579), .ZN(P2_U3309) );
  INV_X1 U14084 ( .A(n11595), .ZN(n11588) );
  NAND2_X1 U14085 ( .A1(n15198), .A2(n14032), .ZN(n11583) );
  NAND2_X1 U14086 ( .A1(n11584), .A2(n11583), .ZN(n11587) );
  INV_X1 U14087 ( .A(n11587), .ZN(n11585) );
  INV_X1 U14088 ( .A(n11637), .ZN(n11586) );
  AOI21_X1 U14089 ( .B1(n11588), .B2(n11587), .A(n11586), .ZN(n11737) );
  INV_X1 U14090 ( .A(n11589), .ZN(n11590) );
  AOI211_X1 U14091 ( .C1(n11767), .C2(n11590), .A(n14822), .B(n11640), .ZN(
        n11740) );
  OAI22_X1 U14092 ( .A1(n11796), .A2(n14307), .B1(n14611), .B2(n11789), .ZN(
        n11591) );
  AOI21_X1 U14093 ( .B1(n11740), .B2(n14604), .A(n11591), .ZN(n11603) );
  OR2_X1 U14094 ( .A1(n15198), .A2(n11592), .ZN(n11593) );
  NAND2_X1 U14095 ( .A1(n11596), .A2(n11595), .ZN(n11597) );
  NAND2_X1 U14096 ( .A1(n11631), .A2(n11597), .ZN(n11598) );
  NAND2_X1 U14097 ( .A1(n11598), .A2(n14255), .ZN(n11600) );
  AOI22_X1 U14098 ( .A1(n14619), .A2(n14032), .B1(n14030), .B2(n14620), .ZN(
        n11599) );
  AND2_X1 U14099 ( .A1(n11600), .A2(n11599), .ZN(n11738) );
  MUX2_X1 U14100 ( .A(n11601), .B(n11738), .S(n14279), .Z(n11602) );
  OAI211_X1 U14101 ( .C1(n11737), .C2(n14286), .A(n11603), .B(n11602), .ZN(
        P1_U3284) );
  INV_X1 U14102 ( .A(n11604), .ZN(n11606) );
  OAI222_X1 U14103 ( .A1(n11607), .A2(P3_U3151), .B1(n13175), .B2(n11606), 
        .C1(n11605), .C2(n13178), .ZN(P3_U3271) );
  NAND2_X1 U14104 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n14058) );
  NAND2_X1 U14105 ( .A1(n15200), .A2(n11608), .ZN(n11609) );
  OAI211_X1 U14106 ( .C1(n15204), .C2(n11610), .A(n14058), .B(n11609), .ZN(
        n11616) );
  NAND2_X1 U14107 ( .A1(n6628), .A2(n11611), .ZN(n11612) );
  XNOR2_X1 U14108 ( .A(n11613), .B(n11612), .ZN(n11614) );
  NOR2_X1 U14109 ( .A1(n11614), .A2(n14731), .ZN(n11615) );
  AOI211_X1 U14110 ( .C1(n11617), .C2(n15197), .A(n11616), .B(n11615), .ZN(
        n11618) );
  INV_X1 U14111 ( .A(n11618), .ZN(P1_U3239) );
  XNOR2_X1 U14112 ( .A(n11619), .B(n12571), .ZN(n15162) );
  OAI211_X1 U14113 ( .C1(n11621), .C2(n12571), .A(n11620), .B(n15112), .ZN(
        n11623) );
  AOI22_X1 U14114 ( .A1(n12707), .A2(n15106), .B1(n15109), .B2(n12709), .ZN(
        n11622) );
  OAI211_X1 U14115 ( .C1(n15116), .C2(n15162), .A(n11623), .B(n11622), .ZN(
        n15163) );
  NAND2_X1 U14116 ( .A1(n15163), .A2(n15122), .ZN(n11629) );
  NOR2_X1 U14117 ( .A1(n11624), .A2(n15169), .ZN(n15164) );
  INV_X1 U14118 ( .A(n11625), .ZN(n11626) );
  OAI22_X1 U14119 ( .A1(n15122), .A2(n15048), .B1(n11626), .B2(n15089), .ZN(
        n11627) );
  AOI21_X1 U14120 ( .B1(n15083), .B2(n15164), .A(n11627), .ZN(n11628) );
  OAI211_X1 U14121 ( .C1(n15162), .C2(n12944), .A(n11629), .B(n11628), .ZN(
        P3_U3224) );
  NAND2_X1 U14122 ( .A1(n11767), .A2(n11766), .ZN(n11630) );
  NAND2_X1 U14123 ( .A1(n11632), .A2(n11638), .ZN(n11633) );
  NAND3_X1 U14124 ( .A1(n11756), .A2(n14614), .A3(n11633), .ZN(n11635) );
  NAND2_X1 U14125 ( .A1(n14031), .A2(n14619), .ZN(n11634) );
  NAND2_X1 U14126 ( .A1(n11635), .A2(n11634), .ZN(n14839) );
  INV_X1 U14127 ( .A(n14839), .ZN(n11649) );
  OR2_X1 U14128 ( .A1(n11767), .A2(n14031), .ZN(n11636) );
  NAND2_X1 U14129 ( .A1(n11637), .A2(n11636), .ZN(n11639) );
  NAND2_X1 U14130 ( .A1(n11639), .A2(n11638), .ZN(n11748) );
  OAI21_X1 U14131 ( .B1(n11639), .B2(n11638), .A(n11748), .ZN(n14841) );
  OAI21_X1 U14132 ( .B1(n11640), .B2(n14838), .A(n14814), .ZN(n11641) );
  OR2_X1 U14133 ( .A1(n11750), .A2(n11641), .ZN(n11643) );
  NAND2_X1 U14134 ( .A1(n14029), .A2(n14620), .ZN(n11642) );
  AND2_X1 U14135 ( .A1(n11643), .A2(n11642), .ZN(n14836) );
  INV_X1 U14136 ( .A(n11644), .ZN(n11865) );
  AOI22_X1 U14137 ( .A1(n14630), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n11865), 
        .B2(n14599), .ZN(n11646) );
  NAND2_X1 U14138 ( .A1(n11853), .A2(n14601), .ZN(n11645) );
  OAI211_X1 U14139 ( .C1(n14836), .C2(n14300), .A(n11646), .B(n11645), .ZN(
        n11647) );
  AOI21_X1 U14140 ( .B1(n14841), .B2(n14631), .A(n11647), .ZN(n11648) );
  OAI21_X1 U14141 ( .B1(n11649), .B2(n14630), .A(n11648), .ZN(P1_U3283) );
  INV_X1 U14142 ( .A(n11650), .ZN(n11688) );
  OAI211_X1 U14143 ( .C1(n11653), .C2(n11652), .A(n11651), .B(n12468), .ZN(
        n11659) );
  INV_X1 U14144 ( .A(n11654), .ZN(n11657) );
  OAI22_X1 U14145 ( .A1(n12441), .A2(n11655), .B1(n15168), .B2(n12477), .ZN(
        n11656) );
  AOI211_X1 U14146 ( .C1(n12439), .C2(n14657), .A(n11657), .B(n11656), .ZN(
        n11658) );
  OAI211_X1 U14147 ( .C1(n11688), .C2(n12034), .A(n11659), .B(n11658), .ZN(
        P3_U3157) );
  INV_X1 U14148 ( .A(n11660), .ZN(n11661) );
  NAND2_X1 U14149 ( .A1(n11662), .A2(n11661), .ZN(n11665) );
  NAND2_X1 U14150 ( .A1(n11663), .A2(n13303), .ZN(n11664) );
  XNOR2_X1 U14151 ( .A(n11813), .B(n6837), .ZN(n15010) );
  INV_X1 U14152 ( .A(n15010), .ZN(n11682) );
  NAND2_X1 U14153 ( .A1(n15003), .A2(n13303), .ZN(n11666) );
  NAND2_X1 U14154 ( .A1(n11669), .A2(n11668), .ZN(n11670) );
  NAND2_X1 U14155 ( .A1(n11818), .A2(n11670), .ZN(n11671) );
  NAND2_X1 U14156 ( .A1(n11671), .A2(n13631), .ZN(n11673) );
  NAND2_X1 U14157 ( .A1(n11673), .A2(n11672), .ZN(n15015) );
  NAND2_X1 U14158 ( .A1(n15013), .A2(n11675), .ZN(n11822) );
  OAI211_X1 U14159 ( .C1(n15013), .C2(n11675), .A(n11674), .B(n11822), .ZN(
        n15011) );
  OAI22_X1 U14160 ( .A1(n14952), .A2(n11677), .B1(n11676), .B2(n14950), .ZN(
        n11678) );
  AOI21_X1 U14161 ( .B1(n11816), .B2(n14955), .A(n11678), .ZN(n11679) );
  OAI21_X1 U14162 ( .B1(n15011), .B2(n14958), .A(n11679), .ZN(n11680) );
  AOI21_X1 U14163 ( .B1(n15015), .B2(n14952), .A(n11680), .ZN(n11681) );
  OAI21_X1 U14164 ( .B1(n11682), .B2(n13646), .A(n11681), .ZN(P2_U3254) );
  XNOR2_X1 U14165 ( .A(n11683), .B(n12587), .ZN(n15171) );
  OR2_X1 U14166 ( .A1(n15075), .A2(n15102), .ZN(n14676) );
  INV_X1 U14167 ( .A(n14664), .ZN(n12998) );
  OAI211_X1 U14168 ( .C1(n11685), .C2(n12508), .A(n11684), .B(n15112), .ZN(
        n11687) );
  AOI22_X1 U14169 ( .A1(n14657), .A2(n15106), .B1(n15109), .B2(n12708), .ZN(
        n11686) );
  NAND2_X1 U14170 ( .A1(n11687), .A2(n11686), .ZN(n15173) );
  NAND2_X1 U14171 ( .A1(n15173), .A2(n15122), .ZN(n11692) );
  INV_X1 U14172 ( .A(n15168), .ZN(n12582) );
  OAI22_X1 U14173 ( .A1(n15122), .A2(n11689), .B1(n11688), .B2(n15089), .ZN(
        n11690) );
  AOI21_X1 U14174 ( .B1(n13027), .B2(n12582), .A(n11690), .ZN(n11691) );
  OAI211_X1 U14175 ( .C1(n15171), .C2(n12998), .A(n11692), .B(n11691), .ZN(
        P3_U3223) );
  INV_X1 U14176 ( .A(n11693), .ZN(n11694) );
  OAI222_X1 U14177 ( .A1(P3_U3151), .A2(n11696), .B1(n13178), .B2(n11695), 
        .C1(n13175), .C2(n11694), .ZN(P3_U3270) );
  NAND2_X1 U14178 ( .A1(n14937), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11705) );
  INV_X1 U14179 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11697) );
  NAND2_X1 U14180 ( .A1(n11719), .A2(n11697), .ZN(n11698) );
  AND2_X1 U14181 ( .A1(n11698), .A2(n11705), .ZN(n14941) );
  MUX2_X1 U14182 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n12207), .S(n14924), .Z(
        n14926) );
  AOI21_X1 U14183 ( .B1(n11700), .B2(P2_REG2_REG_13__SCAN_IN), .A(n11699), 
        .ZN(n11701) );
  OR2_X1 U14184 ( .A1(n11701), .A2(n11713), .ZN(n11702) );
  XNOR2_X1 U14185 ( .A(n11701), .B(n14905), .ZN(n14910) );
  NAND2_X1 U14186 ( .A1(n14910), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n14909) );
  NAND2_X1 U14187 ( .A1(n11702), .A2(n14909), .ZN(n11703) );
  NAND2_X1 U14188 ( .A1(n14915), .A2(n11703), .ZN(n11704) );
  XNOR2_X1 U14189 ( .A(n11715), .B(n11703), .ZN(n14917) );
  NAND2_X1 U14190 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14917), .ZN(n14916) );
  NAND2_X1 U14191 ( .A1(n11704), .A2(n14916), .ZN(n14927) );
  NAND2_X1 U14192 ( .A1(n14926), .A2(n14927), .ZN(n14925) );
  OAI21_X1 U14193 ( .B1(n11717), .B2(n12207), .A(n14925), .ZN(n14940) );
  NAND2_X1 U14194 ( .A1(n14941), .A2(n14940), .ZN(n14938) );
  NAND2_X1 U14195 ( .A1(n11705), .A2(n14938), .ZN(n12055) );
  XNOR2_X1 U14196 ( .A(n12060), .B(n12055), .ZN(n11706) );
  NOR2_X1 U14197 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n11706), .ZN(n12057) );
  AOI21_X1 U14198 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n11706), .A(n12057), 
        .ZN(n11725) );
  INV_X1 U14199 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n11707) );
  NAND2_X1 U14200 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13275)
         );
  OAI21_X1 U14201 ( .B1(n13368), .B2(n11707), .A(n13275), .ZN(n11723) );
  XNOR2_X1 U14202 ( .A(n11719), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14945) );
  INV_X1 U14203 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n13734) );
  XNOR2_X1 U14204 ( .A(n14924), .B(n13734), .ZN(n14929) );
  INV_X1 U14205 ( .A(n11708), .ZN(n11709) );
  OAI21_X1 U14206 ( .B1(n11711), .B2(n11710), .A(n11709), .ZN(n14908) );
  XNOR2_X1 U14207 ( .A(n11713), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n14907) );
  NAND2_X1 U14208 ( .A1(n14908), .A2(n14907), .ZN(n14906) );
  OAI21_X1 U14209 ( .B1(n11713), .B2(n11712), .A(n14906), .ZN(n11714) );
  NAND2_X1 U14210 ( .A1(n14915), .A2(n11714), .ZN(n11716) );
  XNOR2_X1 U14211 ( .A(n11715), .B(n11714), .ZN(n14919) );
  NAND2_X1 U14212 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n14919), .ZN(n14918) );
  NAND2_X1 U14213 ( .A1(n11716), .A2(n14918), .ZN(n14930) );
  NAND2_X1 U14214 ( .A1(n14929), .A2(n14930), .ZN(n14928) );
  OAI21_X1 U14215 ( .B1(n11717), .B2(n13734), .A(n14928), .ZN(n14944) );
  NAND2_X1 U14216 ( .A1(n14945), .A2(n14944), .ZN(n14942) );
  OAI21_X1 U14217 ( .B1(n11719), .B2(n11718), .A(n14942), .ZN(n12059) );
  XOR2_X1 U14218 ( .A(n12060), .B(n12059), .Z(n11720) );
  NAND2_X1 U14219 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n11720), .ZN(n12062) );
  OAI21_X1 U14220 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n11720), .A(n12062), 
        .ZN(n11721) );
  NOR2_X1 U14221 ( .A1(n11721), .A2(n14873), .ZN(n11722) );
  AOI211_X1 U14222 ( .C1(n14936), .C2(n12060), .A(n11723), .B(n11722), .ZN(
        n11724) );
  OAI21_X1 U14223 ( .B1(n11725), .B2(n14874), .A(n11724), .ZN(P2_U3232) );
  INV_X1 U14224 ( .A(n11991), .ZN(n11736) );
  OAI21_X1 U14225 ( .B1(n14278), .B2(n11729), .A(n11726), .ZN(n11990) );
  XOR2_X1 U14226 ( .A(n11990), .B(n11991), .Z(n11727) );
  NAND2_X1 U14227 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n11727), .ZN(n11993) );
  OAI211_X1 U14228 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n11727), .A(n14074), 
        .B(n11993), .ZN(n11735) );
  NAND2_X1 U14229 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13999)
         );
  INV_X1 U14230 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n11730) );
  OAI21_X1 U14231 ( .B1(n11730), .B2(n11729), .A(n11728), .ZN(n11986) );
  XNOR2_X1 U14232 ( .A(n11986), .B(n11736), .ZN(n11731) );
  NAND2_X1 U14233 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n11731), .ZN(n11988) );
  OAI211_X1 U14234 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n11731), .A(n14083), 
        .B(n11988), .ZN(n11732) );
  NAND2_X1 U14235 ( .A1(n13999), .A2(n11732), .ZN(n11733) );
  AOI21_X1 U14236 ( .B1(n14080), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n11733), 
        .ZN(n11734) );
  OAI211_X1 U14237 ( .C1(n11995), .C2(n11736), .A(n11735), .B(n11734), .ZN(
        P1_U3261) );
  INV_X1 U14238 ( .A(n11737), .ZN(n11741) );
  INV_X1 U14239 ( .A(n11738), .ZN(n11739) );
  AOI211_X1 U14240 ( .C1(n11741), .C2(n14842), .A(n11740), .B(n11739), .ZN(
        n11746) );
  INV_X1 U14241 ( .A(n14409), .ZN(n14371) );
  AOI22_X1 U14242 ( .A1(n11767), .A2(n14371), .B1(n14853), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n11742) );
  OAI21_X1 U14243 ( .B1(n11746), .B2(n14853), .A(n11742), .ZN(P1_U3537) );
  INV_X1 U14244 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11743) );
  OAI22_X1 U14245 ( .A1(n11796), .A2(n14446), .B1(n14845), .B2(n11743), .ZN(
        n11744) );
  INV_X1 U14246 ( .A(n11744), .ZN(n11745) );
  OAI21_X1 U14247 ( .B1(n11746), .B2(n14843), .A(n11745), .ZN(P1_U3486) );
  NAND2_X1 U14248 ( .A1(n14838), .A2(n11925), .ZN(n11747) );
  NAND2_X1 U14249 ( .A1(n11748), .A2(n11747), .ZN(n11749) );
  NAND2_X1 U14250 ( .A1(n11749), .A2(n7323), .ZN(n12089) );
  OAI21_X1 U14251 ( .B1(n11749), .B2(n7323), .A(n12089), .ZN(n11870) );
  INV_X1 U14252 ( .A(n11870), .ZN(n11763) );
  INV_X1 U14253 ( .A(n11750), .ZN(n11752) );
  INV_X1 U14254 ( .A(n12107), .ZN(n11751) );
  AOI211_X1 U14255 ( .C1(n12087), .C2(n11752), .A(n14822), .B(n11751), .ZN(
        n11869) );
  NOR2_X1 U14256 ( .A1(n11919), .A2(n14307), .ZN(n11754) );
  OAI22_X1 U14257 ( .A1(n14279), .A2(n10292), .B1(n11929), .B2(n14611), .ZN(
        n11753) );
  AOI211_X1 U14258 ( .C1(n11869), .C2(n14604), .A(n11754), .B(n11753), .ZN(
        n11762) );
  OAI211_X1 U14259 ( .C1(n11758), .C2(n11757), .A(n12081), .B(n14255), .ZN(
        n11760) );
  AOI22_X1 U14260 ( .A1(n14619), .A2(n14030), .B1(n14618), .B2(n14620), .ZN(
        n11759) );
  NAND2_X1 U14261 ( .A1(n11760), .A2(n11759), .ZN(n11868) );
  NAND2_X1 U14262 ( .A1(n11868), .A2(n14279), .ZN(n11761) );
  OAI211_X1 U14263 ( .C1(n11763), .C2(n14286), .A(n11762), .B(n11761), .ZN(
        P1_U3282) );
  INV_X1 U14264 ( .A(n11764), .ZN(n12283) );
  OAI222_X1 U14265 ( .A1(n14474), .A2(n11765), .B1(n14464), .B2(n12283), .C1(
        n14626), .C2(P1_U3086), .ZN(P1_U3336) );
  OAI22_X1 U14266 ( .A1(n11796), .A2(n13938), .B1(n11766), .B2(n10801), .ZN(
        n11850) );
  NAND2_X1 U14267 ( .A1(n11767), .A2(n13902), .ZN(n11769) );
  NAND2_X1 U14268 ( .A1(n14031), .A2(n11103), .ZN(n11768) );
  NAND2_X1 U14269 ( .A1(n11769), .A2(n11768), .ZN(n11770) );
  XNOR2_X1 U14270 ( .A(n11770), .B(n10601), .ZN(n11849) );
  XOR2_X1 U14271 ( .A(n11850), .B(n11849), .Z(n11787) );
  INV_X1 U14272 ( .A(n11771), .ZN(n11774) );
  INV_X1 U14273 ( .A(n11772), .ZN(n11773) );
  NAND2_X1 U14274 ( .A1(n15198), .A2(n13902), .ZN(n11778) );
  NAND2_X1 U14275 ( .A1(n14032), .A2(n11103), .ZN(n11777) );
  NAND2_X1 U14276 ( .A1(n11778), .A2(n11777), .ZN(n11779) );
  XNOR2_X1 U14277 ( .A(n11779), .B(n10601), .ZN(n11783) );
  NAND2_X1 U14278 ( .A1(n15198), .A2(n11103), .ZN(n11781) );
  NAND2_X1 U14279 ( .A1(n14032), .A2(n13906), .ZN(n11780) );
  NAND2_X1 U14280 ( .A1(n11781), .A2(n11780), .ZN(n11782) );
  NOR2_X1 U14281 ( .A1(n11783), .A2(n11782), .ZN(n11784) );
  AOI21_X1 U14282 ( .B1(n11783), .B2(n11782), .A(n11784), .ZN(n15195) );
  INV_X1 U14283 ( .A(n11784), .ZN(n11785) );
  OAI21_X1 U14284 ( .B1(n11787), .B2(n11786), .A(n11859), .ZN(n11788) );
  NAND2_X1 U14285 ( .A1(n11788), .A2(n15206), .ZN(n11795) );
  INV_X1 U14286 ( .A(n11789), .ZN(n11793) );
  AOI21_X1 U14287 ( .B1(n14705), .B2(n14032), .A(n11790), .ZN(n11791) );
  OAI21_X1 U14288 ( .B1(n11925), .B2(n14728), .A(n11791), .ZN(n11792) );
  AOI21_X1 U14289 ( .B1(n11793), .B2(n14018), .A(n11792), .ZN(n11794) );
  OAI211_X1 U14290 ( .C1(n11796), .C2(n14707), .A(n11795), .B(n11794), .ZN(
        P1_U3231) );
  INV_X1 U14291 ( .A(n11797), .ZN(n11799) );
  OAI222_X1 U14292 ( .A1(n11800), .A2(P3_U3151), .B1(n13175), .B2(n11799), 
        .C1(n11798), .C2(n12293), .ZN(P3_U3269) );
  NAND3_X1 U14293 ( .A1(n11801), .A2(n13189), .A3(n13300), .ZN(n11802) );
  OAI21_X1 U14294 ( .B1(n14861), .B2(n13269), .A(n11802), .ZN(n11805) );
  INV_X1 U14295 ( .A(n11803), .ZN(n11804) );
  NAND2_X1 U14296 ( .A1(n11805), .A2(n11804), .ZN(n11811) );
  NOR2_X1 U14297 ( .A1(n14870), .A2(n12022), .ZN(n11809) );
  AND2_X1 U14298 ( .A1(n13300), .A2(n13576), .ZN(n11806) );
  AOI21_X1 U14299 ( .B1(n13298), .B2(n13578), .A(n11806), .ZN(n12016) );
  OAI22_X1 U14300 ( .A1(n14859), .A2(n12016), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11807), .ZN(n11808) );
  AOI211_X1 U14301 ( .C1(n13744), .C2(n14867), .A(n11809), .B(n11808), .ZN(
        n11810) );
  OAI211_X1 U14302 ( .C1(n11812), .C2(n13269), .A(n11811), .B(n11810), .ZN(
        P2_U3187) );
  OR2_X1 U14303 ( .A1(n11816), .A2(n13302), .ZN(n11814) );
  XNOR2_X1 U14304 ( .A(n11904), .B(n11903), .ZN(n11935) );
  INV_X1 U14305 ( .A(n11935), .ZN(n11829) );
  NAND2_X1 U14306 ( .A1(n11816), .A2(n11815), .ZN(n11817) );
  INV_X1 U14307 ( .A(n11903), .ZN(n11819) );
  OAI211_X1 U14308 ( .C1(n6625), .C2(n11819), .A(n11906), .B(n13631), .ZN(
        n11821) );
  AOI22_X1 U14309 ( .A1(n13576), .A2(n13302), .B1(n13300), .B2(n15413), .ZN(
        n11820) );
  NAND2_X1 U14310 ( .A1(n11821), .A2(n11820), .ZN(n11933) );
  NAND2_X1 U14311 ( .A1(n11933), .A2(n14952), .ZN(n11828) );
  AOI211_X1 U14312 ( .C1(n13221), .C2(n11822), .A(n11080), .B(n7103), .ZN(
        n11934) );
  INV_X1 U14313 ( .A(n13221), .ZN(n11823) );
  NOR2_X1 U14314 ( .A1(n11823), .A2(n13640), .ZN(n11826) );
  OAI22_X1 U14315 ( .A1(n14952), .A2(n11824), .B1(n13219), .B2(n14950), .ZN(
        n11825) );
  AOI211_X1 U14316 ( .C1(n11934), .C2(n13649), .A(n11826), .B(n11825), .ZN(
        n11827) );
  OAI211_X1 U14317 ( .C1(n11829), .C2(n13646), .A(n11828), .B(n11827), .ZN(
        P2_U3253) );
  AOI21_X1 U14318 ( .B1(n11831), .B2(n8454), .A(n11941), .ZN(n11848) );
  MUX2_X1 U14319 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12824), .Z(n11948) );
  XNOR2_X1 U14320 ( .A(n7231), .B(n11948), .ZN(n11836) );
  OR2_X1 U14321 ( .A1(n11832), .A2(n11842), .ZN(n11834) );
  NAND2_X1 U14322 ( .A1(n11834), .A2(n11833), .ZN(n11835) );
  OAI21_X1 U14323 ( .B1(n11836), .B2(n11835), .A(n11950), .ZN(n11837) );
  NAND2_X1 U14324 ( .A1(n11837), .A2(n15052), .ZN(n11840) );
  INV_X1 U14325 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11838) );
  NOR2_X1 U14326 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11838), .ZN(n11882) );
  INV_X1 U14327 ( .A(n11882), .ZN(n11839) );
  OAI211_X1 U14328 ( .C1(n15066), .C2(n14497), .A(n11840), .B(n11839), .ZN(
        n11846) );
  INV_X1 U14329 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14693) );
  AOI21_X1 U14330 ( .B1(n14693), .B2(n11843), .A(n6511), .ZN(n11844) );
  NOR2_X1 U14331 ( .A1(n11844), .A2(n15060), .ZN(n11845) );
  AOI211_X1 U14332 ( .C1(n15054), .C2(n7231), .A(n11846), .B(n11845), .ZN(
        n11847) );
  OAI21_X1 U14333 ( .B1(n11848), .B2(n15056), .A(n11847), .ZN(P3_U3193) );
  INV_X1 U14334 ( .A(n11849), .ZN(n11852) );
  INV_X1 U14335 ( .A(n11850), .ZN(n11851) );
  NAND2_X1 U14336 ( .A1(n11852), .A2(n11851), .ZN(n11857) );
  AND2_X1 U14337 ( .A1(n11859), .A2(n11857), .ZN(n11861) );
  OAI22_X1 U14338 ( .A1(n14838), .A2(n13938), .B1(n11925), .B2(n10801), .ZN(
        n11920) );
  NAND2_X1 U14339 ( .A1(n11853), .A2(n13902), .ZN(n11855) );
  NAND2_X1 U14340 ( .A1(n14030), .A2(n11103), .ZN(n11854) );
  NAND2_X1 U14341 ( .A1(n11855), .A2(n11854), .ZN(n11856) );
  XNOR2_X1 U14342 ( .A(n11856), .B(n10601), .ZN(n11921) );
  XOR2_X1 U14343 ( .A(n11920), .B(n11921), .Z(n11860) );
  OAI211_X1 U14344 ( .C1(n11861), .C2(n11860), .A(n15206), .B(n11922), .ZN(
        n11867) );
  INV_X1 U14345 ( .A(n14029), .ZN(n12079) );
  AOI21_X1 U14346 ( .B1(n14705), .B2(n14031), .A(n11862), .ZN(n11863) );
  OAI21_X1 U14347 ( .B1(n12079), .B2(n14728), .A(n11863), .ZN(n11864) );
  AOI21_X1 U14348 ( .B1(n11865), .B2(n14018), .A(n11864), .ZN(n11866) );
  OAI211_X1 U14349 ( .C1(n14838), .C2(n14707), .A(n11867), .B(n11866), .ZN(
        P1_U3217) );
  AOI211_X1 U14350 ( .C1(n14842), .C2(n11870), .A(n11869), .B(n11868), .ZN(
        n11874) );
  AOI22_X1 U14351 ( .A1(n12087), .A2(n14371), .B1(n14853), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n11871) );
  OAI21_X1 U14352 ( .B1(n11874), .B2(n14853), .A(n11871), .ZN(P1_U3539) );
  OAI22_X1 U14353 ( .A1(n11919), .A2(n14446), .B1(n14845), .B2(n9525), .ZN(
        n11872) );
  INV_X1 U14354 ( .A(n11872), .ZN(n11873) );
  OAI21_X1 U14355 ( .B1(n11874), .B2(n14843), .A(n11873), .ZN(P1_U3492) );
  INV_X1 U14356 ( .A(n11875), .ZN(n11877) );
  INV_X1 U14357 ( .A(SI_27_), .ZN(n11876) );
  OAI222_X1 U14358 ( .A1(n13175), .A2(n11877), .B1(n13178), .B2(n11876), .C1(
        P3_U3151), .C2(n12824), .ZN(P3_U3268) );
  INV_X1 U14359 ( .A(n11878), .ZN(n11880) );
  NAND2_X1 U14360 ( .A1(n11880), .A2(n11879), .ZN(n11881) );
  XNOR2_X1 U14361 ( .A(n11881), .B(n14657), .ZN(n11888) );
  NOR2_X1 U14362 ( .A1(n12477), .A2(n14677), .ZN(n11887) );
  INV_X1 U14363 ( .A(n14678), .ZN(n11885) );
  AOI21_X1 U14364 ( .B1(n12439), .B2(n12706), .A(n11882), .ZN(n11884) );
  NAND2_X1 U14365 ( .A1(n12470), .A2(n12707), .ZN(n11883) );
  OAI211_X1 U14366 ( .C1(n12034), .C2(n11885), .A(n11884), .B(n11883), .ZN(
        n11886) );
  AOI211_X1 U14367 ( .C1(n11888), .C2(n12468), .A(n11887), .B(n11886), .ZN(
        n11889) );
  INV_X1 U14368 ( .A(n11889), .ZN(P3_U3176) );
  XNOR2_X1 U14369 ( .A(n11890), .B(n12706), .ZN(n11891) );
  XNOR2_X1 U14370 ( .A(n11892), .B(n11891), .ZN(n11893) );
  NAND2_X1 U14371 ( .A1(n11893), .A2(n12468), .ZN(n11899) );
  NAND2_X1 U14372 ( .A1(n12470), .A2(n14657), .ZN(n11896) );
  NAND2_X1 U14373 ( .A1(n12439), .A2(n14658), .ZN(n11895) );
  INV_X1 U14374 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11894) );
  OR2_X1 U14375 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11894), .ZN(n11955) );
  NAND3_X1 U14376 ( .A1(n11896), .A2(n11895), .A3(n11955), .ZN(n11897) );
  AOI21_X1 U14377 ( .B1(n12474), .B2(n14660), .A(n11897), .ZN(n11898) );
  OAI211_X1 U14378 ( .C1(n14663), .C2(n12477), .A(n11899), .B(n11898), .ZN(
        P3_U3164) );
  INV_X1 U14379 ( .A(n11900), .ZN(n11939) );
  OAI222_X1 U14380 ( .A1(n14474), .A2(n11902), .B1(n14472), .B2(n11939), .C1(
        n11901), .C2(P1_U3086), .ZN(P1_U3335) );
  XNOR2_X1 U14381 ( .A(n12005), .B(n11907), .ZN(n12075) );
  INV_X1 U14382 ( .A(n12075), .ZN(n11917) );
  OAI211_X1 U14383 ( .C1(n11908), .C2(n11907), .A(n12010), .B(n13631), .ZN(
        n11909) );
  AOI22_X1 U14384 ( .A1(n13299), .A2(n15413), .B1(n13576), .B2(n13301), .ZN(
        n14858) );
  NAND2_X1 U14385 ( .A1(n11909), .A2(n14858), .ZN(n12073) );
  AOI21_X1 U14386 ( .B1(n14868), .B2(n11910), .A(n11080), .ZN(n11911) );
  NAND2_X1 U14387 ( .A1(n11911), .A2(n12018), .ZN(n12071) );
  NAND2_X1 U14388 ( .A1(n14964), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11912) );
  OAI21_X1 U14389 ( .B1(n14950), .B2(n14871), .A(n11912), .ZN(n11913) );
  AOI21_X1 U14390 ( .B1(n14868), .B2(n14955), .A(n11913), .ZN(n11914) );
  OAI21_X1 U14391 ( .B1(n12071), .B2(n14958), .A(n11914), .ZN(n11915) );
  AOI21_X1 U14392 ( .B1(n12073), .B2(n14952), .A(n11915), .ZN(n11916) );
  OAI21_X1 U14393 ( .B1(n13646), .B2(n11917), .A(n11916), .ZN(P2_U3252) );
  OAI22_X1 U14394 ( .A1(n11919), .A2(n13936), .B1(n12079), .B2(n13938), .ZN(
        n11918) );
  XNOR2_X1 U14395 ( .A(n11918), .B(n13940), .ZN(n12039) );
  OAI22_X1 U14396 ( .A1(n11919), .A2(n13938), .B1(n12079), .B2(n10801), .ZN(
        n12040) );
  XNOR2_X1 U14397 ( .A(n12039), .B(n12040), .ZN(n11924) );
  AOI21_X1 U14398 ( .B1(n11924), .B2(n11923), .A(n6615), .ZN(n11932) );
  NOR2_X1 U14399 ( .A1(n14725), .A2(n11925), .ZN(n11926) );
  AOI211_X1 U14400 ( .C1(n14703), .C2(n14618), .A(n11927), .B(n11926), .ZN(
        n11928) );
  OAI21_X1 U14401 ( .B1(n11929), .B2(n15204), .A(n11928), .ZN(n11930) );
  AOI21_X1 U14402 ( .B1(n12087), .B2(n15197), .A(n11930), .ZN(n11931) );
  OAI21_X1 U14403 ( .B1(n11932), .B2(n14731), .A(n11931), .ZN(P1_U3236) );
  AOI211_X1 U14404 ( .C1(n15009), .C2(n11935), .A(n11934), .B(n11933), .ZN(
        n11938) );
  AOI22_X1 U14405 ( .A1(n13221), .A2(n13745), .B1(P2_REG1_REG_12__SCAN_IN), 
        .B2(n15025), .ZN(n11936) );
  OAI21_X1 U14406 ( .B1(n11938), .B2(n15025), .A(n11936), .ZN(P2_U3511) );
  AOI22_X1 U14407 ( .A1(n13221), .A2(n13783), .B1(P2_REG0_REG_12__SCAN_IN), 
        .B2(n15017), .ZN(n11937) );
  OAI21_X1 U14408 ( .B1(n11938), .B2(n15017), .A(n11937), .ZN(P2_U3466) );
  OAI222_X1 U14409 ( .A1(n13807), .A2(n11940), .B1(P2_U3088), .B2(n6863), .C1(
        n13794), .C2(n11939), .ZN(P2_U3307) );
  NOR2_X1 U14410 ( .A1(n7231), .A2(n6596), .ZN(n11942) );
  NOR2_X1 U14411 ( .A1(n11942), .A2(n11941), .ZN(n11945) );
  INV_X1 U14412 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U14413 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n11964), .B1(n12726), 
        .B2(n11943), .ZN(n11944) );
  NOR2_X1 U14414 ( .A1(n11945), .A2(n11944), .ZN(n12713) );
  AOI21_X1 U14415 ( .B1(n11945), .B2(n11944), .A(n12713), .ZN(n11966) );
  INV_X1 U14416 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14499) );
  MUX2_X1 U14417 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12824), .Z(n11946) );
  AND2_X1 U14418 ( .A1(n11946), .A2(n12726), .ZN(n12719) );
  NOR2_X1 U14419 ( .A1(n11946), .A2(n12726), .ZN(n11947) );
  NOR2_X1 U14420 ( .A1(n12719), .A2(n11947), .ZN(n11954) );
  OR2_X1 U14421 ( .A1(n11949), .A2(n11948), .ZN(n11951) );
  INV_X1 U14422 ( .A(n12718), .ZN(n11952) );
  OAI211_X1 U14423 ( .C1(n11954), .C2(n11953), .A(n11952), .B(n15052), .ZN(
        n11956) );
  OAI211_X1 U14424 ( .C1(n15066), .C2(n14499), .A(n11956), .B(n11955), .ZN(
        n11963) );
  NOR2_X1 U14425 ( .A1(n7231), .A2(n11957), .ZN(n11958) );
  INV_X1 U14426 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14688) );
  AOI22_X1 U14427 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n11964), .B1(n12726), 
        .B2(n14688), .ZN(n11959) );
  AOI21_X1 U14428 ( .B1(n11960), .B2(n11959), .A(n12725), .ZN(n11961) );
  NOR2_X1 U14429 ( .A1(n11961), .A2(n15060), .ZN(n11962) );
  AOI211_X1 U14430 ( .C1(n15054), .C2(n11964), .A(n11963), .B(n11962), .ZN(
        n11965) );
  OAI21_X1 U14431 ( .B1(n11966), .B2(n15056), .A(n11965), .ZN(P3_U3194) );
  AOI22_X1 U14432 ( .A1(n11967), .A2(n14860), .B1(n13189), .B2(n13298), .ZN(
        n11975) );
  INV_X1 U14433 ( .A(n11968), .ZN(n11974) );
  AND2_X1 U14434 ( .A1(n13299), .A2(n13576), .ZN(n11969) );
  AOI21_X1 U14435 ( .B1(n13391), .B2(n15413), .A(n11969), .ZN(n12168) );
  INV_X1 U14436 ( .A(n12168), .ZN(n11970) );
  AOI22_X1 U14437 ( .A1(n13238), .A2(n11970), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11971) );
  OAI21_X1 U14438 ( .B1(n12170), .B2(n14870), .A(n11971), .ZN(n11972) );
  AOI21_X1 U14439 ( .B1(n13782), .B2(n14867), .A(n11972), .ZN(n11973) );
  OAI21_X1 U14440 ( .B1(n11975), .B2(n11974), .A(n11973), .ZN(P2_U3213) );
  INV_X1 U14441 ( .A(n11976), .ZN(n11979) );
  OAI222_X1 U14442 ( .A1(n13175), .A2(n11979), .B1(n13178), .B2(n11978), .C1(
        P3_U3151), .C2(n6870), .ZN(P3_U3267) );
  INV_X1 U14443 ( .A(n11980), .ZN(n11984) );
  OAI222_X1 U14444 ( .A1(n14474), .A2(n11982), .B1(n14472), .B2(n11984), .C1(
        P1_U3086), .C2(n11981), .ZN(P1_U3334) );
  OAI222_X1 U14445 ( .A1(n13807), .A2(n11985), .B1(n13805), .B2(n11984), .C1(
        n11983), .C2(P2_U3088), .ZN(P2_U3306) );
  NAND2_X1 U14446 ( .A1(n11991), .A2(n11986), .ZN(n11987) );
  NAND2_X1 U14447 ( .A1(n11988), .A2(n11987), .ZN(n11989) );
  XOR2_X1 U14448 ( .A(n11989), .B(P1_REG1_REG_19__SCAN_IN), .Z(n11999) );
  INV_X1 U14449 ( .A(n11999), .ZN(n11997) );
  NAND2_X1 U14450 ( .A1(n11991), .A2(n11990), .ZN(n11992) );
  NAND2_X1 U14451 ( .A1(n11993), .A2(n11992), .ZN(n11994) );
  XOR2_X1 U14452 ( .A(n11994), .B(P1_REG2_REG_19__SCAN_IN), .Z(n11998) );
  OAI21_X1 U14453 ( .B1(n11998), .B2(n14781), .A(n11995), .ZN(n11996) );
  AOI21_X1 U14454 ( .B1(n14083), .B2(n11997), .A(n11996), .ZN(n12001) );
  AOI22_X1 U14455 ( .A1(n11999), .A2(n14083), .B1(n11998), .B2(n14074), .ZN(
        n12000) );
  MUX2_X1 U14456 ( .A(n12001), .B(n12000), .S(n14626), .Z(n12002) );
  NAND2_X1 U14457 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13927)
         );
  OAI211_X1 U14458 ( .C1(n12003), .C2(n14792), .A(n12002), .B(n13927), .ZN(
        P1_U3262) );
  OR2_X1 U14459 ( .A1(n14868), .A2(n13300), .ZN(n12004) );
  NAND2_X1 U14460 ( .A1(n14868), .A2(n13300), .ZN(n12006) );
  NAND2_X1 U14461 ( .A1(n12007), .A2(n12006), .ZN(n12161) );
  XNOR2_X1 U14462 ( .A(n12161), .B(n12011), .ZN(n12192) );
  INV_X1 U14463 ( .A(n12192), .ZN(n12028) );
  INV_X1 U14464 ( .A(n13300), .ZN(n12008) );
  OR2_X1 U14465 ( .A1(n14868), .A2(n12008), .ZN(n12009) );
  INV_X1 U14466 ( .A(n12011), .ZN(n12012) );
  NAND2_X1 U14467 ( .A1(n12013), .A2(n12012), .ZN(n12014) );
  NAND2_X1 U14468 ( .A1(n12165), .A2(n12014), .ZN(n12015) );
  NAND2_X1 U14469 ( .A1(n12015), .A2(n13631), .ZN(n12017) );
  NAND2_X1 U14470 ( .A1(n12017), .A2(n12016), .ZN(n12195) );
  NAND2_X1 U14471 ( .A1(n12195), .A2(n14952), .ZN(n12027) );
  AOI21_X1 U14472 ( .B1(n13744), .B2(n12018), .A(n11080), .ZN(n12021) );
  AND2_X1 U14473 ( .A1(n12021), .A2(n12172), .ZN(n12193) );
  INV_X1 U14474 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n12023) );
  OAI22_X1 U14475 ( .A1(n14952), .A2(n12023), .B1(n12022), .B2(n14950), .ZN(
        n12025) );
  NOR2_X1 U14476 ( .A1(n12019), .A2(n13640), .ZN(n12024) );
  AOI211_X1 U14477 ( .C1(n12193), .C2(n13649), .A(n12025), .B(n12024), .ZN(
        n12026) );
  OAI211_X1 U14478 ( .C1(n12028), .C2(n13646), .A(n12027), .B(n12026), .ZN(
        P2_U3251) );
  NOR2_X1 U14479 ( .A1(n12029), .A2(n6636), .ZN(n12030) );
  XNOR2_X1 U14480 ( .A(n12031), .B(n12030), .ZN(n12038) );
  INV_X1 U14481 ( .A(n12477), .ZN(n12459) );
  NAND2_X1 U14482 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12723)
         );
  OAI21_X1 U14483 ( .B1(n12472), .B2(n14647), .A(n12723), .ZN(n12032) );
  AOI21_X1 U14484 ( .B1(n12470), .B2(n12706), .A(n12032), .ZN(n12033) );
  OAI21_X1 U14485 ( .B1(n14648), .B2(n12034), .A(n12033), .ZN(n12035) );
  AOI21_X1 U14486 ( .B1(n12459), .B2(n12036), .A(n12035), .ZN(n12037) );
  OAI21_X1 U14487 ( .B1(n12038), .B2(n12462), .A(n12037), .ZN(P3_U3174) );
  INV_X1 U14488 ( .A(n12039), .ZN(n12042) );
  INV_X1 U14489 ( .A(n12040), .ZN(n12041) );
  NAND2_X1 U14490 ( .A1(n14602), .A2(n13902), .ZN(n12044) );
  NAND2_X1 U14491 ( .A1(n14618), .A2(n11103), .ZN(n12043) );
  NAND2_X1 U14492 ( .A1(n12044), .A2(n12043), .ZN(n12045) );
  XNOR2_X1 U14493 ( .A(n12045), .B(n13812), .ZN(n12048) );
  AND2_X1 U14494 ( .A1(n14618), .A2(n13906), .ZN(n12046) );
  AOI21_X1 U14495 ( .B1(n14602), .B2(n11103), .A(n12046), .ZN(n12047) );
  NOR2_X1 U14496 ( .A1(n12048), .A2(n12047), .ZN(n12228) );
  NOR2_X1 U14497 ( .A1(n12228), .A2(n6629), .ZN(n12049) );
  XNOR2_X1 U14498 ( .A(n12229), .B(n12049), .ZN(n12054) );
  AOI22_X1 U14499 ( .A1(n14704), .A2(n14620), .B1(n14619), .B2(n14029), .ZN(
        n12111) );
  OAI22_X1 U14500 ( .A1(n12111), .A2(n14015), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12050), .ZN(n12051) );
  AOI21_X1 U14501 ( .B1(n14600), .B2(n14018), .A(n12051), .ZN(n12053) );
  NAND2_X1 U14502 ( .A1(n14602), .A2(n15197), .ZN(n12052) );
  OAI211_X1 U14503 ( .C1(n12054), .C2(n14731), .A(n12053), .B(n12052), .ZN(
        P1_U3224) );
  INV_X1 U14504 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n15373) );
  NOR2_X1 U14505 ( .A1(n12060), .A2(n12055), .ZN(n12056) );
  NOR2_X1 U14506 ( .A1(n12057), .A2(n12056), .ZN(n12058) );
  XOR2_X1 U14507 ( .A(n12058), .B(P2_REG2_REG_19__SCAN_IN), .Z(n12067) );
  INV_X1 U14508 ( .A(n12067), .ZN(n12065) );
  NAND2_X1 U14509 ( .A1(n12060), .A2(n12059), .ZN(n12061) );
  NAND2_X1 U14510 ( .A1(n12062), .A2(n12061), .ZN(n12063) );
  XOR2_X1 U14511 ( .A(n12063), .B(P2_REG1_REG_19__SCAN_IN), .Z(n12066) );
  NOR2_X1 U14512 ( .A1(n12066), .A2(n14873), .ZN(n12064) );
  AOI211_X1 U14513 ( .C1(n12065), .C2(n14939), .A(n14936), .B(n12064), .ZN(
        n12069) );
  AOI22_X1 U14514 ( .A1(n12067), .A2(n14939), .B1(n14943), .B2(n12066), .ZN(
        n12068) );
  MUX2_X1 U14515 ( .A(n12069), .B(n12068), .S(n12284), .Z(n12070) );
  NAND2_X1 U14516 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13203)
         );
  OAI211_X1 U14517 ( .C1(n15373), .C2(n13368), .A(n12070), .B(n13203), .ZN(
        P2_U3233) );
  INV_X1 U14518 ( .A(n14868), .ZN(n12072) );
  INV_X1 U14519 ( .A(n14990), .ZN(n15012) );
  OAI21_X1 U14520 ( .B1(n12072), .B2(n15012), .A(n12071), .ZN(n12074) );
  AOI211_X1 U14521 ( .C1(n12075), .C2(n15009), .A(n12074), .B(n12073), .ZN(
        n12078) );
  NAND2_X1 U14522 ( .A1(n15017), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n12076) );
  OAI21_X1 U14523 ( .B1(n12078), .B2(n15017), .A(n12076), .ZN(P2_U3469) );
  NAND2_X1 U14524 ( .A1(n15025), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n12077) );
  OAI21_X1 U14525 ( .B1(n12078), .B2(n15025), .A(n12077), .ZN(P2_U3512) );
  OR2_X1 U14526 ( .A1(n12087), .A2(n12079), .ZN(n12080) );
  INV_X1 U14527 ( .A(n14618), .ZN(n12221) );
  OR2_X1 U14528 ( .A1(n14602), .A2(n12221), .ZN(n12082) );
  INV_X1 U14529 ( .A(n14628), .ZN(n14616) );
  NAND2_X1 U14530 ( .A1(n14745), .A2(n14704), .ZN(n12083) );
  OAI211_X1 U14531 ( .C1(n12084), .C2(n12095), .A(n12137), .B(n14614), .ZN(
        n12086) );
  AOI22_X1 U14532 ( .A1(n14704), .A2(n14619), .B1(n14620), .B2(n14702), .ZN(
        n12085) );
  NAND2_X1 U14533 ( .A1(n12086), .A2(n12085), .ZN(n14740) );
  INV_X1 U14534 ( .A(n14740), .ZN(n12103) );
  OR2_X1 U14535 ( .A1(n12087), .A2(n14029), .ZN(n12088) );
  NAND2_X1 U14536 ( .A1(n12089), .A2(n12088), .ZN(n12106) );
  INV_X1 U14537 ( .A(n12109), .ZN(n12105) );
  NAND2_X1 U14538 ( .A1(n12106), .A2(n12105), .ZN(n12104) );
  OR2_X1 U14539 ( .A1(n14602), .A2(n14618), .ZN(n12090) );
  NAND2_X1 U14540 ( .A1(n12104), .A2(n12090), .ZN(n14629) );
  NAND2_X1 U14541 ( .A1(n14629), .A2(n14628), .ZN(n12092) );
  NAND2_X1 U14542 ( .A1(n14745), .A2(n12224), .ZN(n12091) );
  NAND2_X1 U14543 ( .A1(n12092), .A2(n12091), .ZN(n12094) );
  INV_X1 U14544 ( .A(n12149), .ZN(n12093) );
  AOI21_X1 U14545 ( .B1(n12095), .B2(n12094), .A(n12093), .ZN(n14742) );
  INV_X1 U14546 ( .A(n14610), .ZN(n12096) );
  OAI21_X1 U14547 ( .B1(n7008), .B2(n12096), .A(n12143), .ZN(n14739) );
  OAI22_X1 U14548 ( .A1(n14279), .A2(n12097), .B1(n14712), .B2(n14611), .ZN(
        n12098) );
  AOI21_X1 U14549 ( .B1(n13820), .B2(n14601), .A(n12098), .ZN(n12099) );
  OAI21_X1 U14550 ( .B1(n14739), .B2(n12100), .A(n12099), .ZN(n12101) );
  AOI21_X1 U14551 ( .B1(n14742), .B2(n14631), .A(n12101), .ZN(n12102) );
  OAI21_X1 U14552 ( .B1(n14630), .B2(n12103), .A(n12102), .ZN(P1_U3279) );
  INV_X1 U14553 ( .A(n14796), .ZN(n14827) );
  OAI21_X1 U14554 ( .B1(n12106), .B2(n12105), .A(n12104), .ZN(n14606) );
  AOI211_X1 U14555 ( .C1(n14602), .C2(n12107), .A(n14822), .B(n6627), .ZN(
        n14603) );
  OAI211_X1 U14556 ( .C1(n12110), .C2(n12109), .A(n12108), .B(n14255), .ZN(
        n12112) );
  NAND2_X1 U14557 ( .A1(n12112), .A2(n12111), .ZN(n12113) );
  AOI21_X1 U14558 ( .B1(n14112), .B2(n14606), .A(n12113), .ZN(n14609) );
  INV_X1 U14559 ( .A(n14609), .ZN(n12114) );
  AOI211_X1 U14560 ( .C1(n14827), .C2(n14606), .A(n14603), .B(n12114), .ZN(
        n12118) );
  INV_X1 U14561 ( .A(n14446), .ZN(n14432) );
  NOR2_X1 U14562 ( .A1(n14845), .A2(n9538), .ZN(n12115) );
  AOI21_X1 U14563 ( .B1(n14602), .B2(n14432), .A(n12115), .ZN(n12116) );
  OAI21_X1 U14564 ( .B1(n12118), .B2(n14843), .A(n12116), .ZN(P1_U3495) );
  AOI22_X1 U14565 ( .A1(n14602), .A2(n14371), .B1(n14853), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n12117) );
  OAI21_X1 U14566 ( .B1(n12118), .B2(n14853), .A(n12117), .ZN(P1_U3540) );
  XOR2_X1 U14567 ( .A(n12120), .B(n12119), .Z(n12125) );
  NAND2_X1 U14568 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(P3_U3151), .ZN(n12743)
         );
  NAND2_X1 U14569 ( .A1(n12470), .A2(n14658), .ZN(n12121) );
  OAI211_X1 U14570 ( .C1(n12472), .C2(n12412), .A(n12743), .B(n12121), .ZN(
        n12123) );
  NOR2_X1 U14571 ( .A1(n12243), .A2(n12477), .ZN(n12122) );
  AOI211_X1 U14572 ( .C1(n12131), .C2(n12474), .A(n12123), .B(n12122), .ZN(
        n12124) );
  OAI21_X1 U14573 ( .B1(n12125), .B2(n12462), .A(n12124), .ZN(P3_U3155) );
  OAI211_X1 U14574 ( .C1(n12127), .C2(n8520), .A(n15112), .B(n12126), .ZN(
        n12129) );
  AOI22_X1 U14575 ( .A1(n14658), .A2(n15109), .B1(n15106), .B2(n12704), .ZN(
        n12128) );
  NAND2_X1 U14576 ( .A1(n12129), .A2(n12128), .ZN(n12236) );
  INV_X1 U14577 ( .A(n12236), .ZN(n12135) );
  XNOR2_X1 U14578 ( .A(n12130), .B(n8520), .ZN(n12237) );
  AOI22_X1 U14579 ( .A1(n15124), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15119), 
        .B2(n12131), .ZN(n12132) );
  OAI21_X1 U14580 ( .B1(n12243), .B2(n13044), .A(n12132), .ZN(n12133) );
  AOI21_X1 U14581 ( .B1(n12237), .B2(n14664), .A(n12133), .ZN(n12134) );
  OAI21_X1 U14582 ( .B1(n12135), .B2(n15124), .A(n12134), .ZN(P3_U3219) );
  OAI211_X1 U14583 ( .C1(n12138), .C2(n12330), .A(n12306), .B(n14255), .ZN(
        n12140) );
  AOI22_X1 U14584 ( .A1(n14621), .A2(n14619), .B1(n14620), .B2(n14028), .ZN(
        n14016) );
  AND2_X1 U14585 ( .A1(n12140), .A2(n14016), .ZN(n14406) );
  INV_X1 U14586 ( .A(n14019), .ZN(n12141) );
  OAI22_X1 U14587 ( .A1(n14279), .A2(n12142), .B1(n12141), .B2(n14611), .ZN(
        n12147) );
  NAND2_X1 U14588 ( .A1(n13828), .A2(n12143), .ZN(n12144) );
  NAND2_X1 U14589 ( .A1(n12144), .A2(n14814), .ZN(n12145) );
  OR2_X1 U14590 ( .A1(n14294), .A2(n12145), .ZN(n14404) );
  NOR2_X1 U14591 ( .A1(n14404), .A2(n14300), .ZN(n12146) );
  AOI211_X1 U14592 ( .C1(n14601), .C2(n13828), .A(n12147), .B(n12146), .ZN(
        n12151) );
  NAND2_X1 U14593 ( .A1(n13820), .A2(n14621), .ZN(n12148) );
  XNOR2_X1 U14594 ( .A(n12329), .B(n12330), .ZN(n14403) );
  NAND2_X1 U14595 ( .A1(n14403), .A2(n14631), .ZN(n12150) );
  OAI211_X1 U14596 ( .C1(n14406), .C2(n14630), .A(n12151), .B(n12150), .ZN(
        P1_U3278) );
  INV_X1 U14597 ( .A(n12152), .ZN(n13163) );
  OAI211_X1 U14598 ( .C1(n12155), .C2(n12154), .A(n12153), .B(n12468), .ZN(
        n12159) );
  AND2_X1 U14599 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12763) );
  AOI21_X1 U14600 ( .B1(n12470), .B2(n12705), .A(n12763), .ZN(n12156) );
  OAI21_X1 U14601 ( .B1(n12472), .B2(n12424), .A(n12156), .ZN(n12157) );
  AOI21_X1 U14602 ( .B1(n12187), .B2(n12474), .A(n12157), .ZN(n12158) );
  OAI211_X1 U14603 ( .C1(n13163), .C2(n12477), .A(n12159), .B(n12158), .ZN(
        P3_U3181) );
  AND2_X1 U14604 ( .A1(n13744), .A2(n13299), .ZN(n12160) );
  OR2_X1 U14605 ( .A1(n13744), .A2(n13299), .ZN(n12162) );
  XNOR2_X1 U14606 ( .A(n12201), .B(n7137), .ZN(n13739) );
  INV_X1 U14607 ( .A(n13299), .ZN(n12163) );
  NAND2_X1 U14608 ( .A1(n13744), .A2(n12163), .ZN(n12164) );
  NAND2_X1 U14609 ( .A1(n12166), .A2(n12200), .ZN(n12167) );
  NAND3_X1 U14610 ( .A1(n12211), .A2(n13631), .A3(n12167), .ZN(n12169) );
  AND2_X1 U14611 ( .A1(n12169), .A2(n12168), .ZN(n13738) );
  OAI21_X1 U14612 ( .B1(n12170), .B2(n14950), .A(n13738), .ZN(n12171) );
  NAND2_X1 U14613 ( .A1(n12171), .A2(n14952), .ZN(n12180) );
  NAND2_X1 U14614 ( .A1(n13782), .A2(n12172), .ZN(n12173) );
  NAND2_X1 U14615 ( .A1(n12173), .A2(n11674), .ZN(n12174) );
  OR2_X1 U14616 ( .A1(n12204), .A2(n12174), .ZN(n13737) );
  INV_X1 U14617 ( .A(n13737), .ZN(n12178) );
  INV_X1 U14618 ( .A(n13782), .ZN(n12176) );
  OAI22_X1 U14619 ( .A1(n12176), .A2(n13640), .B1(n14952), .B2(n12175), .ZN(
        n12177) );
  AOI21_X1 U14620 ( .B1(n12178), .B2(n13649), .A(n12177), .ZN(n12179) );
  OAI211_X1 U14621 ( .C1(n13739), .C2(n13646), .A(n12180), .B(n12179), .ZN(
        P2_U3250) );
  OAI211_X1 U14622 ( .C1(n12183), .C2(n12182), .A(n12181), .B(n15112), .ZN(
        n12185) );
  AOI22_X1 U14623 ( .A1(n15109), .A2(n12705), .B1(n13035), .B2(n15106), .ZN(
        n12184) );
  NAND2_X1 U14624 ( .A1(n12185), .A2(n12184), .ZN(n13112) );
  INV_X1 U14625 ( .A(n13112), .ZN(n12191) );
  XNOR2_X1 U14626 ( .A(n12186), .B(n12606), .ZN(n13113) );
  AOI22_X1 U14627 ( .A1(n15124), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15119), 
        .B2(n12187), .ZN(n12188) );
  OAI21_X1 U14628 ( .B1(n13163), .B2(n13044), .A(n12188), .ZN(n12189) );
  AOI21_X1 U14629 ( .B1(n13113), .B2(n14664), .A(n12189), .ZN(n12190) );
  OAI21_X1 U14630 ( .B1(n12191), .B2(n15124), .A(n12190), .ZN(P3_U3218) );
  AND2_X1 U14631 ( .A1(n12192), .A2(n15009), .ZN(n12194) );
  INV_X1 U14632 ( .A(n13742), .ZN(n12196) );
  MUX2_X1 U14633 ( .A(n12197), .B(n12196), .S(n15018), .Z(n12198) );
  OAI21_X1 U14634 ( .B1(n12019), .B2(n13778), .A(n12198), .ZN(P2_U3472) );
  NOR2_X1 U14635 ( .A1(n13782), .A2(n13298), .ZN(n12199) );
  OR2_X1 U14636 ( .A1(n12202), .A2(n12212), .ZN(n12203) );
  INV_X1 U14637 ( .A(n13733), .ZN(n12219) );
  INV_X1 U14638 ( .A(n12204), .ZN(n12206) );
  NAND2_X1 U14639 ( .A1(n13779), .A2(n12204), .ZN(n13635) );
  INV_X1 U14640 ( .A(n13635), .ZN(n12205) );
  AOI211_X1 U14641 ( .C1(n13419), .C2(n12206), .A(n11080), .B(n12205), .ZN(
        n13732) );
  NOR2_X1 U14642 ( .A1(n13779), .A2(n13640), .ZN(n12209) );
  OAI22_X1 U14643 ( .A1(n14952), .A2(n12207), .B1(n13231), .B2(n14950), .ZN(
        n12208) );
  AOI211_X1 U14644 ( .C1(n13732), .C2(n13649), .A(n12209), .B(n12208), .ZN(
        n12218) );
  INV_X1 U14645 ( .A(n12212), .ZN(n12213) );
  OAI211_X1 U14646 ( .C1(n12214), .C2(n12213), .A(n13421), .B(n13631), .ZN(
        n12216) );
  AND2_X1 U14647 ( .A1(n13298), .A2(n13576), .ZN(n12215) );
  AOI21_X1 U14648 ( .B1(n13394), .B2(n15413), .A(n12215), .ZN(n13233) );
  NAND2_X1 U14649 ( .A1(n12216), .A2(n13233), .ZN(n13731) );
  NAND2_X1 U14650 ( .A1(n13731), .A2(n14952), .ZN(n12217) );
  OAI211_X1 U14651 ( .C1(n12219), .C2(n13646), .A(n12218), .B(n12217), .ZN(
        P2_U3249) );
  OAI21_X1 U14652 ( .B1(n14725), .B2(n12221), .A(n12220), .ZN(n12222) );
  AOI21_X1 U14653 ( .B1(n14703), .B2(n14621), .A(n12222), .ZN(n12223) );
  OAI21_X1 U14654 ( .B1(n14612), .B2(n15204), .A(n12223), .ZN(n12233) );
  OAI22_X1 U14655 ( .A1(n14745), .A2(n13936), .B1(n12224), .B2(n13938), .ZN(
        n12225) );
  XNOR2_X1 U14656 ( .A(n12225), .B(n13940), .ZN(n13815) );
  OR2_X1 U14657 ( .A1(n14745), .A2(n13938), .ZN(n12227) );
  NAND2_X1 U14658 ( .A1(n14704), .A2(n13906), .ZN(n12226) );
  NAND2_X1 U14659 ( .A1(n12227), .A2(n12226), .ZN(n13816) );
  XNOR2_X1 U14660 ( .A(n13815), .B(n13816), .ZN(n12231) );
  AOI211_X1 U14661 ( .C1(n12231), .C2(n12230), .A(n14731), .B(n13814), .ZN(
        n12232) );
  AOI211_X1 U14662 ( .C1(n12234), .C2(n15197), .A(n12233), .B(n12232), .ZN(
        n12235) );
  INV_X1 U14663 ( .A(n12235), .ZN(P1_U3234) );
  INV_X1 U14664 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12238) );
  AOI21_X1 U14665 ( .B1(n14692), .B2(n12237), .A(n12236), .ZN(n12240) );
  MUX2_X1 U14666 ( .A(n12238), .B(n12240), .S(n15193), .Z(n12239) );
  OAI21_X1 U14667 ( .B1(n13116), .B2(n12243), .A(n12239), .ZN(P3_U3473) );
  INV_X1 U14668 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12241) );
  MUX2_X1 U14669 ( .A(n12241), .B(n12240), .S(n15176), .Z(n12242) );
  OAI21_X1 U14670 ( .B1(n13162), .B2(n12243), .A(n12242), .ZN(P3_U3432) );
  NAND2_X1 U14671 ( .A1(n12248), .A2(n12244), .ZN(n12246) );
  OAI211_X1 U14672 ( .C1(n15248), .C2(n14474), .A(n12246), .B(n12245), .ZN(
        P1_U3332) );
  NAND2_X1 U14673 ( .A1(n12248), .A2(n12247), .ZN(n12250) );
  OAI211_X1 U14674 ( .C1(n12251), .C2(n13807), .A(n12250), .B(n12249), .ZN(
        P2_U3304) );
  OAI211_X1 U14675 ( .C1(n12254), .C2(n12253), .A(n12252), .B(n15112), .ZN(
        n12256) );
  AOI22_X1 U14676 ( .A1(n13021), .A2(n15106), .B1(n15109), .B2(n12704), .ZN(
        n12255) );
  NAND2_X1 U14677 ( .A1(n12256), .A2(n12255), .ZN(n13108) );
  INV_X1 U14678 ( .A(n13108), .ZN(n12261) );
  XNOR2_X1 U14679 ( .A(n12257), .B(n12512), .ZN(n13109) );
  AOI22_X1 U14680 ( .A1(n15124), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15119), 
        .B2(n12415), .ZN(n12258) );
  OAI21_X1 U14681 ( .B1(n13158), .B2(n13044), .A(n12258), .ZN(n12259) );
  AOI21_X1 U14682 ( .B1(n13109), .B2(n14664), .A(n12259), .ZN(n12260) );
  OAI21_X1 U14683 ( .B1(n12261), .B2(n15124), .A(n12260), .ZN(P3_U3217) );
  OAI222_X1 U14684 ( .A1(n13175), .A2(n12263), .B1(n12293), .B2(n12262), .C1(
        P3_U3151), .C2(n12859), .ZN(P3_U3276) );
  INV_X1 U14685 ( .A(n12264), .ZN(n12280) );
  INV_X1 U14686 ( .A(n12266), .ZN(n13249) );
  AOI21_X1 U14687 ( .B1(n13249), .B2(n7084), .A(n13269), .ZN(n12271) );
  INV_X1 U14688 ( .A(n13412), .ZN(n13434) );
  NOR3_X1 U14689 ( .A1(n12268), .A2(n13434), .A3(n8233), .ZN(n12270) );
  OAI21_X1 U14690 ( .B1(n12271), .B2(n12270), .A(n12269), .ZN(n12278) );
  INV_X1 U14691 ( .A(n13506), .ZN(n12276) );
  NAND2_X1 U14692 ( .A1(n13438), .A2(n15413), .ZN(n12273) );
  NAND2_X1 U14693 ( .A1(n13412), .A2(n13576), .ZN(n12272) );
  AND2_X1 U14694 ( .A1(n12273), .A2(n12272), .ZN(n13504) );
  OAI22_X1 U14695 ( .A1(n14859), .A2(n13504), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12274), .ZN(n12275) );
  AOI21_X1 U14696 ( .B1(n13277), .B2(n12276), .A(n12275), .ZN(n12277) );
  OAI211_X1 U14697 ( .C1(n13512), .C2(n13281), .A(n12278), .B(n12277), .ZN(
        P2_U3197) );
  OAI222_X1 U14698 ( .A1(n13805), .A2(n12280), .B1(P2_U3088), .B2(n12279), 
        .C1(n12290), .C2(n13807), .ZN(P2_U3297) );
  INV_X1 U14699 ( .A(n12281), .ZN(n14454) );
  OAI222_X1 U14700 ( .A1(n13805), .A2(n14454), .B1(P2_U3088), .B2(n7720), .C1(
        n12282), .C2(n13807), .ZN(P2_U3298) );
  OAI222_X1 U14701 ( .A1(n13807), .A2(n12285), .B1(P2_U3088), .B2(n12284), 
        .C1(n13805), .C2(n12283), .ZN(P2_U3308) );
  INV_X1 U14702 ( .A(n12286), .ZN(n12287) );
  NAND2_X1 U14703 ( .A1(n14455), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12289) );
  XNOR2_X1 U14704 ( .A(n12290), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n12483) );
  XNOR2_X1 U14705 ( .A(n12484), .B(n12483), .ZN(n12478) );
  INV_X1 U14706 ( .A(n12478), .ZN(n12291) );
  OAI222_X1 U14707 ( .A1(n12294), .A2(P3_U3151), .B1(n12293), .B2(n12292), 
        .C1(n13175), .C2(n12291), .ZN(P3_U3265) );
  INV_X1 U14708 ( .A(n12295), .ZN(n12296) );
  AOI22_X1 U14709 ( .A1(n12296), .A2(n14860), .B1(n13189), .B2(n13406), .ZN(
        n12303) );
  INV_X1 U14710 ( .A(n13579), .ZN(n13556) );
  OAI22_X1 U14711 ( .A1(n13556), .A2(n12298), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12297), .ZN(n12299) );
  AOI21_X1 U14712 ( .B1(n13284), .B2(n13520), .A(n12299), .ZN(n12300) );
  OAI21_X1 U14713 ( .B1(n13549), .B2(n14870), .A(n12300), .ZN(n12301) );
  AOI21_X1 U14714 ( .B1(n13548), .B2(n14867), .A(n12301), .ZN(n12302) );
  OAI21_X1 U14715 ( .B1(n12304), .B2(n12303), .A(n12302), .ZN(P2_U3207) );
  INV_X1 U14716 ( .A(n14028), .ZN(n14726) );
  NAND2_X1 U14717 ( .A1(n14721), .A2(n14726), .ZN(n12308) );
  INV_X1 U14718 ( .A(n14270), .ZN(n14281) );
  INV_X1 U14719 ( .A(n14296), .ZN(n14714) );
  OR2_X1 U14720 ( .A1(n14735), .A2(n14714), .ZN(n12309) );
  OR2_X1 U14721 ( .A1(n14385), .A2(n14727), .ZN(n12311) );
  INV_X1 U14722 ( .A(n14247), .ZN(n14244) );
  NAND2_X1 U14723 ( .A1(n14237), .A2(n12312), .ZN(n12313) );
  INV_X1 U14724 ( .A(n14197), .ZN(n12315) );
  OR2_X1 U14725 ( .A1(n14431), .A2(n12315), .ZN(n12316) );
  INV_X1 U14726 ( .A(n14025), .ZN(n13919) );
  INV_X1 U14727 ( .A(n14196), .ZN(n13993) );
  AND2_X1 U14728 ( .A1(n14356), .A2(n13993), .ZN(n12317) );
  INV_X1 U14729 ( .A(n14142), .ZN(n13918) );
  OR2_X1 U14730 ( .A1(n14351), .A2(n13918), .ZN(n12318) );
  INV_X1 U14731 ( .A(n14159), .ZN(n12319) );
  INV_X1 U14732 ( .A(n14143), .ZN(n13967) );
  OR2_X1 U14733 ( .A1(n14130), .A2(n13967), .ZN(n12321) );
  INV_X1 U14734 ( .A(n14100), .ZN(n14106) );
  NAND2_X1 U14735 ( .A1(n12364), .A2(n12324), .ZN(n12328) );
  NAND2_X1 U14736 ( .A1(n14023), .A2(n14620), .ZN(n12326) );
  NAND2_X1 U14737 ( .A1(n14024), .A2(n14619), .ZN(n12325) );
  OR2_X1 U14738 ( .A1(n13828), .A2(n14702), .ZN(n12331) );
  NAND2_X1 U14739 ( .A1(n14292), .A2(n14291), .ZN(n14290) );
  OR2_X1 U14740 ( .A1(n14721), .A2(n14028), .ZN(n12332) );
  NAND2_X1 U14741 ( .A1(n14385), .A2(n14027), .ZN(n12335) );
  NAND2_X1 U14742 ( .A1(n14192), .A2(n14191), .ZN(n14190) );
  OR2_X1 U14743 ( .A1(n14193), .A2(n14025), .ZN(n12336) );
  NAND2_X1 U14744 ( .A1(n14356), .A2(n14196), .ZN(n12338) );
  OR2_X1 U14745 ( .A1(n14351), .A2(n14142), .ZN(n12339) );
  NAND2_X1 U14746 ( .A1(n14148), .A2(n14147), .ZN(n14146) );
  OAI21_X1 U14747 ( .B1(n12343), .B2(n12342), .A(n12352), .ZN(n14332) );
  INV_X1 U14748 ( .A(n14332), .ZN(n12350) );
  INV_X1 U14749 ( .A(n14330), .ZN(n13939) );
  INV_X1 U14750 ( .A(n14721), .ZN(n14398) );
  NAND2_X1 U14751 ( .A1(n14437), .A2(n14240), .ZN(n14228) );
  OR2_X1 U14752 ( .A1(n14228), .A2(n14431), .ZN(n14212) );
  AOI21_X1 U14753 ( .B1(n14114), .B2(n14330), .A(n14822), .ZN(n12346) );
  NAND2_X1 U14754 ( .A1(n14329), .A2(n14604), .ZN(n12348) );
  AOI22_X1 U14755 ( .A1(n14630), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n13945), 
        .B2(n14599), .ZN(n12347) );
  OAI211_X1 U14756 ( .C1(n13939), .C2(n14307), .A(n12348), .B(n12347), .ZN(
        n12349) );
  AOI21_X1 U14757 ( .B1(n12350), .B2(n14631), .A(n12349), .ZN(n12351) );
  OAI21_X1 U14758 ( .B1(n14335), .B2(n14630), .A(n12351), .ZN(P1_U3265) );
  INV_X1 U14759 ( .A(n14327), .ZN(n12361) );
  NAND2_X1 U14760 ( .A1(n12354), .A2(P1_B_REG_SCAN_IN), .ZN(n12355) );
  AND2_X1 U14761 ( .A1(n14620), .A2(n12355), .ZN(n14091) );
  NAND2_X1 U14762 ( .A1(n14022), .A2(n14091), .ZN(n14324) );
  INV_X1 U14763 ( .A(n12356), .ZN(n12357) );
  OAI22_X1 U14764 ( .A1(n12358), .A2(n14324), .B1(n12357), .B2(n14611), .ZN(
        n12359) );
  AOI21_X1 U14765 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n14630), .A(n12359), 
        .ZN(n12360) );
  OAI21_X1 U14766 ( .B1(n12361), .B2(n14307), .A(n12360), .ZN(n12362) );
  AOI21_X1 U14767 ( .B1(n14325), .B2(n14604), .A(n12362), .ZN(n12368) );
  NAND2_X1 U14768 ( .A1(n12364), .A2(n12363), .ZN(n12366) );
  XNOR2_X1 U14769 ( .A(n12366), .B(n12365), .ZN(n12367) );
  NAND2_X1 U14770 ( .A1(n14107), .A2(n14619), .ZN(n14323) );
  INV_X1 U14771 ( .A(n12369), .ZN(n12370) );
  OAI222_X1 U14772 ( .A1(n13807), .A2(n12371), .B1(n13805), .B2(n12370), .C1(
        n9923), .C2(P2_U3088), .ZN(P2_U3305) );
  INV_X1 U14773 ( .A(n12373), .ZN(n12374) );
  AOI21_X1 U14774 ( .B1(n12701), .B2(n12372), .A(n12374), .ZN(n12379) );
  AOI22_X1 U14775 ( .A1(n12702), .A2(n12470), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12376) );
  NAND2_X1 U14776 ( .A1(n12474), .A2(n12955), .ZN(n12375) );
  OAI211_X1 U14777 ( .C1(n12948), .C2(n12472), .A(n12376), .B(n12375), .ZN(
        n12377) );
  AOI21_X1 U14778 ( .B1(n12952), .B2(n12459), .A(n12377), .ZN(n12378) );
  OAI21_X1 U14779 ( .B1(n12379), .B2(n12462), .A(n12378), .ZN(P3_U3156) );
  XNOR2_X1 U14780 ( .A(n12381), .B(n12380), .ZN(n12386) );
  NAND2_X1 U14781 ( .A1(n12470), .A2(n13036), .ZN(n12382) );
  NAND2_X1 U14782 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12858)
         );
  OAI211_X1 U14783 ( .C1(n12472), .C2(n12974), .A(n12382), .B(n12858), .ZN(
        n12384) );
  NOR2_X1 U14784 ( .A1(n13151), .A2(n12477), .ZN(n12383) );
  AOI211_X1 U14785 ( .C1(n13013), .C2(n12474), .A(n12384), .B(n12383), .ZN(
        n12385) );
  OAI21_X1 U14786 ( .B1(n12386), .B2(n12462), .A(n12385), .ZN(P3_U3159) );
  INV_X1 U14787 ( .A(n12388), .ZN(n12392) );
  NOR3_X1 U14788 ( .A1(n12437), .A2(n12390), .A3(n12389), .ZN(n12391) );
  OAI21_X1 U14789 ( .B1(n12392), .B2(n12391), .A(n12468), .ZN(n12396) );
  AOI22_X1 U14790 ( .A1(n12470), .A2(n13004), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12393) );
  OAI21_X1 U14791 ( .B1(n12975), .B2(n12472), .A(n12393), .ZN(n12394) );
  AOI21_X1 U14792 ( .B1(n12978), .B2(n12474), .A(n12394), .ZN(n12395) );
  OAI211_X1 U14793 ( .C1(n13146), .C2(n12477), .A(n12396), .B(n12395), .ZN(
        P3_U3163) );
  INV_X1 U14794 ( .A(n13066), .ZN(n12926) );
  INV_X1 U14795 ( .A(n12397), .ZN(n12402) );
  NOR3_X1 U14796 ( .A1(n12398), .A2(n12400), .A3(n12399), .ZN(n12401) );
  OAI21_X1 U14797 ( .B1(n12402), .B2(n12401), .A(n12468), .ZN(n12407) );
  AOI22_X1 U14798 ( .A1(n12920), .A2(n12470), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12403) );
  OAI21_X1 U14799 ( .B1(n12404), .B2(n12472), .A(n12403), .ZN(n12405) );
  AOI21_X1 U14800 ( .B1(n12924), .B2(n12474), .A(n12405), .ZN(n12406) );
  OAI211_X1 U14801 ( .C1(n12926), .C2(n12477), .A(n12407), .B(n12406), .ZN(
        P3_U3165) );
  AOI21_X1 U14802 ( .B1(n12410), .B2(n12409), .A(n12408), .ZN(n12417) );
  AOI22_X1 U14803 ( .A1(n12439), .A2(n13021), .B1(P3_REG3_REG_16__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12411) );
  OAI21_X1 U14804 ( .B1(n12412), .B2(n12441), .A(n12411), .ZN(n12414) );
  NOR2_X1 U14805 ( .A1(n13158), .A2(n12477), .ZN(n12413) );
  AOI211_X1 U14806 ( .C1(n12415), .C2(n12474), .A(n12414), .B(n12413), .ZN(
        n12416) );
  OAI21_X1 U14807 ( .B1(n12417), .B2(n12462), .A(n12416), .ZN(P3_U3166) );
  XNOR2_X1 U14808 ( .A(n12419), .B(n12418), .ZN(n12420) );
  XNOR2_X1 U14809 ( .A(n12421), .B(n12420), .ZN(n12427) );
  NAND2_X1 U14810 ( .A1(n12474), .A2(n13042), .ZN(n12423) );
  AND2_X1 U14811 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12806) );
  AOI21_X1 U14812 ( .B1(n12439), .B2(n13036), .A(n12806), .ZN(n12422) );
  OAI211_X1 U14813 ( .C1(n12424), .C2(n12441), .A(n12423), .B(n12422), .ZN(
        n12425) );
  AOI21_X1 U14814 ( .B1(n13041), .B2(n12459), .A(n12425), .ZN(n12426) );
  OAI21_X1 U14815 ( .B1(n12427), .B2(n12462), .A(n12426), .ZN(P3_U3168) );
  INV_X1 U14816 ( .A(n12941), .ZN(n13072) );
  AND3_X1 U14817 ( .A1(n12373), .A2(n12429), .A3(n12428), .ZN(n12430) );
  OAI21_X1 U14818 ( .B1(n12398), .B2(n12430), .A(n12468), .ZN(n12434) );
  AOI22_X1 U14819 ( .A1(n12904), .A2(n12439), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12431) );
  OAI21_X1 U14820 ( .B1(n12962), .B2(n12441), .A(n12431), .ZN(n12432) );
  AOI21_X1 U14821 ( .B1(n12940), .B2(n12474), .A(n12432), .ZN(n12433) );
  OAI211_X1 U14822 ( .C1(n13072), .C2(n12477), .A(n12434), .B(n12433), .ZN(
        P3_U3169) );
  INV_X1 U14823 ( .A(n13090), .ZN(n12445) );
  NOR2_X1 U14824 ( .A1(n12436), .A2(n12435), .ZN(n12438) );
  OAI21_X1 U14825 ( .B1(n12438), .B2(n12437), .A(n12468), .ZN(n12444) );
  AOI22_X1 U14826 ( .A1(n12988), .A2(n12439), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12440) );
  OAI21_X1 U14827 ( .B1(n12457), .B2(n12441), .A(n12440), .ZN(n12442) );
  AOI21_X1 U14828 ( .B1(n12995), .B2(n12474), .A(n12442), .ZN(n12443) );
  OAI211_X1 U14829 ( .C1(n12445), .C2(n12477), .A(n12444), .B(n12443), .ZN(
        P3_U3173) );
  INV_X1 U14830 ( .A(n12447), .ZN(n12448) );
  AOI21_X1 U14831 ( .B1(n12702), .B2(n12446), .A(n12448), .ZN(n12453) );
  AOI22_X1 U14832 ( .A1(n12988), .A2(n12470), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12450) );
  NAND2_X1 U14833 ( .A1(n12474), .A2(n12967), .ZN(n12449) );
  OAI211_X1 U14834 ( .C1(n12962), .C2(n12472), .A(n12450), .B(n12449), .ZN(
        n12451) );
  AOI21_X1 U14835 ( .B1(n12966), .B2(n12459), .A(n12451), .ZN(n12452) );
  OAI21_X1 U14836 ( .B1(n12453), .B2(n12462), .A(n12452), .ZN(P3_U3175) );
  XNOR2_X1 U14837 ( .A(n12455), .B(n12454), .ZN(n12463) );
  NAND2_X1 U14838 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(P3_U3151), .ZN(n12828)
         );
  NAND2_X1 U14839 ( .A1(n12470), .A2(n13021), .ZN(n12456) );
  OAI211_X1 U14840 ( .C1(n12472), .C2(n12457), .A(n12828), .B(n12456), .ZN(
        n12458) );
  AOI21_X1 U14841 ( .B1(n13024), .B2(n12474), .A(n12458), .ZN(n12461) );
  NAND2_X1 U14842 ( .A1(n13098), .A2(n12459), .ZN(n12460) );
  OAI211_X1 U14843 ( .C1(n12463), .C2(n12462), .A(n12461), .B(n12460), .ZN(
        P3_U3178) );
  OAI21_X1 U14844 ( .B1(n12467), .B2(n12465), .A(n12466), .ZN(n12469) );
  NAND2_X1 U14845 ( .A1(n12469), .A2(n12468), .ZN(n12476) );
  AOI22_X1 U14846 ( .A1(n12904), .A2(n12470), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12471) );
  OAI21_X1 U14847 ( .B1(n12668), .B2(n12472), .A(n12471), .ZN(n12473) );
  AOI21_X1 U14848 ( .B1(n12911), .B2(n12474), .A(n12473), .ZN(n12475) );
  OAI211_X1 U14849 ( .C1(n13133), .C2(n12477), .A(n12476), .B(n12475), .ZN(
        P3_U3180) );
  NAND2_X1 U14850 ( .A1(n12478), .A2(n12487), .ZN(n12481) );
  NAND2_X1 U14851 ( .A1(n12479), .A2(SI_30_), .ZN(n12480) );
  NOR2_X1 U14852 ( .A1(n13122), .A2(n12498), .ZN(n12680) );
  OAI22_X1 U14853 ( .A1(n12484), .A2(n12483), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n12482), .ZN(n12486) );
  XNOR2_X1 U14854 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12485) );
  XNOR2_X1 U14855 ( .A(n12486), .B(n12485), .ZN(n13167) );
  NAND2_X1 U14856 ( .A1(n12479), .A2(SI_31_), .ZN(n12488) );
  INV_X1 U14857 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12492) );
  NAND2_X1 U14858 ( .A1(n8313), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12491) );
  NAND2_X1 U14859 ( .A1(n12489), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12490) );
  OAI211_X1 U14860 ( .C1(n12493), .C2(n12492), .A(n12491), .B(n12490), .ZN(
        n12494) );
  INV_X1 U14861 ( .A(n12494), .ZN(n12495) );
  AND2_X1 U14862 ( .A1(n13117), .A2(n12866), .ZN(n12684) );
  NAND2_X1 U14863 ( .A1(n13122), .A2(n12498), .ZN(n12499) );
  INV_X1 U14864 ( .A(n12866), .ZN(n12699) );
  OAI21_X1 U14865 ( .B1(n13052), .B2(n12699), .A(n12678), .ZN(n12500) );
  NAND4_X1 U14866 ( .A1(n12505), .A2(n15072), .A3(n12504), .A4(n12503), .ZN(
        n12506) );
  NOR4_X1 U14867 ( .A1(n15092), .A2(n12547), .A3(n12506), .A4(n15111), .ZN(
        n12507) );
  NAND3_X1 U14868 ( .A1(n12507), .A2(n12562), .A3(n12569), .ZN(n12509) );
  NOR4_X1 U14869 ( .A1(n12571), .A2(n14671), .A3(n12509), .A4(n12508), .ZN(
        n12510) );
  AND4_X1 U14870 ( .A1(n12601), .A2(n14661), .A3(n14649), .A4(n12510), .ZN(
        n12511) );
  NAND4_X1 U14871 ( .A1(n13039), .A2(n12606), .A3(n12512), .A4(n12511), .ZN(
        n12513) );
  NOR4_X1 U14872 ( .A1(n12991), .A2(n13028), .A3(n13008), .A4(n12513), .ZN(
        n12517) );
  INV_X1 U14873 ( .A(n12514), .ZN(n12516) );
  NAND4_X1 U14874 ( .A1(n12953), .A2(n12964), .A3(n12517), .A4(n12976), .ZN(
        n12518) );
  NOR4_X1 U14875 ( .A1(n12902), .A2(n12918), .A3(n12933), .A4(n12518), .ZN(
        n12519) );
  XNOR2_X1 U14876 ( .A(n12520), .B(n12859), .ZN(n12689) );
  INV_X1 U14877 ( .A(n12902), .ZN(n12906) );
  INV_X1 U14878 ( .A(n12523), .ZN(n12525) );
  NAND2_X1 U14879 ( .A1(n12525), .A2(n12695), .ZN(n12528) );
  NAND2_X1 U14880 ( .A1(n12525), .A2(n12524), .ZN(n12526) );
  NAND3_X1 U14881 ( .A1(n8883), .A2(n12675), .A3(n12526), .ZN(n12527) );
  OAI21_X1 U14882 ( .B1(n15111), .B2(n12528), .A(n12527), .ZN(n12531) );
  NAND2_X1 U14883 ( .A1(n15105), .A2(n12529), .ZN(n12530) );
  NAND2_X1 U14884 ( .A1(n12531), .A2(n12530), .ZN(n12535) );
  MUX2_X1 U14885 ( .A(n8883), .B(n12532), .S(n12675), .Z(n12533) );
  NAND3_X1 U14886 ( .A1(n12535), .A2(n12534), .A3(n12533), .ZN(n12540) );
  NAND2_X1 U14887 ( .A1(n12536), .A2(n12545), .ZN(n12537) );
  NAND2_X1 U14888 ( .A1(n12537), .A2(n12657), .ZN(n12539) );
  INV_X1 U14889 ( .A(n12542), .ZN(n12538) );
  AOI21_X1 U14890 ( .B1(n12540), .B2(n12539), .A(n12538), .ZN(n12544) );
  AOI21_X1 U14891 ( .B1(n12542), .B2(n12541), .A(n12657), .ZN(n12543) );
  OR2_X1 U14892 ( .A1(n12544), .A2(n12543), .ZN(n12549) );
  NOR2_X1 U14893 ( .A1(n12545), .A2(n12657), .ZN(n12546) );
  NOR2_X1 U14894 ( .A1(n12547), .A2(n12546), .ZN(n12548) );
  NAND2_X1 U14895 ( .A1(n12549), .A2(n12548), .ZN(n12554) );
  NAND3_X1 U14896 ( .A1(n12554), .A2(n15072), .A3(n12550), .ZN(n12552) );
  NAND3_X1 U14897 ( .A1(n12552), .A2(n12551), .A3(n12556), .ZN(n12561) );
  NAND3_X1 U14898 ( .A1(n12554), .A2(n15072), .A3(n12553), .ZN(n12559) );
  AND2_X1 U14899 ( .A1(n12564), .A2(n12555), .ZN(n12558) );
  INV_X1 U14900 ( .A(n12556), .ZN(n12557) );
  AOI21_X1 U14901 ( .B1(n12559), .B2(n12558), .A(n12557), .ZN(n12560) );
  MUX2_X1 U14902 ( .A(n12561), .B(n12560), .S(n12657), .Z(n12563) );
  OAI211_X1 U14903 ( .C1(n12657), .C2(n12564), .A(n12563), .B(n12562), .ZN(
        n12570) );
  NAND2_X1 U14904 ( .A1(n12565), .A2(n12710), .ZN(n12566) );
  MUX2_X1 U14905 ( .A(n12567), .B(n12566), .S(n12675), .Z(n12568) );
  NAND3_X1 U14906 ( .A1(n12570), .A2(n12569), .A3(n12568), .ZN(n12576) );
  INV_X1 U14907 ( .A(n12571), .ZN(n12575) );
  MUX2_X1 U14908 ( .A(n12573), .B(n12572), .S(n12657), .Z(n12574) );
  NAND3_X1 U14909 ( .A1(n12576), .A2(n12575), .A3(n12574), .ZN(n12581) );
  MUX2_X1 U14910 ( .A(n12708), .B(n12577), .S(n12657), .Z(n12579) );
  NAND2_X1 U14911 ( .A1(n12579), .A2(n12578), .ZN(n12580) );
  NAND2_X1 U14912 ( .A1(n12581), .A2(n12580), .ZN(n12588) );
  INV_X1 U14913 ( .A(n14671), .ZN(n14669) );
  NAND2_X1 U14914 ( .A1(n12582), .A2(n14674), .ZN(n12583) );
  MUX2_X1 U14915 ( .A(n12584), .B(n12583), .S(n12657), .Z(n12585) );
  NAND2_X1 U14916 ( .A1(n14669), .A2(n12585), .ZN(n12586) );
  AOI21_X1 U14917 ( .B1(n12588), .B2(n12587), .A(n12586), .ZN(n12597) );
  NAND2_X1 U14918 ( .A1(n12594), .A2(n12589), .ZN(n12592) );
  NAND2_X1 U14919 ( .A1(n12593), .A2(n12590), .ZN(n12591) );
  MUX2_X1 U14920 ( .A(n12592), .B(n12591), .S(n12675), .Z(n12596) );
  MUX2_X1 U14921 ( .A(n12594), .B(n12593), .S(n12657), .Z(n12595) );
  OAI21_X1 U14922 ( .B1(n12597), .B2(n12596), .A(n12595), .ZN(n12598) );
  NAND2_X1 U14923 ( .A1(n12598), .A2(n14649), .ZN(n12602) );
  MUX2_X1 U14924 ( .A(n12599), .B(n6516), .S(n12657), .Z(n12600) );
  NAND3_X1 U14925 ( .A1(n12602), .A2(n12601), .A3(n12600), .ZN(n12607) );
  MUX2_X1 U14926 ( .A(n12604), .B(n12603), .S(n12675), .Z(n12605) );
  NAND3_X1 U14927 ( .A1(n12607), .A2(n12606), .A3(n12605), .ZN(n12612) );
  NAND2_X1 U14928 ( .A1(n12615), .A2(n12608), .ZN(n12609) );
  NAND2_X1 U14929 ( .A1(n12609), .A2(n12675), .ZN(n12611) );
  INV_X1 U14930 ( .A(n12614), .ZN(n12610) );
  AOI21_X1 U14931 ( .B1(n12612), .B2(n12611), .A(n12610), .ZN(n12617) );
  AOI21_X1 U14932 ( .B1(n12614), .B2(n12613), .A(n12675), .ZN(n12616) );
  OAI22_X1 U14933 ( .A1(n12617), .A2(n12616), .B1(n12615), .B2(n12675), .ZN(
        n12624) );
  INV_X1 U14934 ( .A(n12618), .ZN(n12623) );
  INV_X1 U14935 ( .A(n12619), .ZN(n12620) );
  NAND2_X1 U14936 ( .A1(n12625), .A2(n12620), .ZN(n12621) );
  NAND4_X1 U14937 ( .A1(n12631), .A2(n12657), .A3(n12622), .A4(n12621), .ZN(
        n12627) );
  AOI22_X1 U14938 ( .A1(n12624), .A2(n13039), .B1(n12623), .B2(n12627), .ZN(
        n12629) );
  NAND3_X1 U14939 ( .A1(n12630), .A2(n12625), .A3(n12675), .ZN(n12626) );
  NAND2_X1 U14940 ( .A1(n12627), .A2(n12626), .ZN(n12628) );
  OAI21_X1 U14941 ( .B1(n12629), .B2(n13028), .A(n12628), .ZN(n12633) );
  INV_X1 U14942 ( .A(n12991), .ZN(n12985) );
  MUX2_X1 U14943 ( .A(n12631), .B(n12630), .S(n12657), .Z(n12632) );
  NAND3_X1 U14944 ( .A1(n12633), .A2(n12985), .A3(n12632), .ZN(n12637) );
  MUX2_X1 U14945 ( .A(n12635), .B(n12634), .S(n12657), .Z(n12636) );
  NAND3_X1 U14946 ( .A1(n12637), .A2(n12976), .A3(n12636), .ZN(n12641) );
  MUX2_X1 U14947 ( .A(n12639), .B(n12638), .S(n12675), .Z(n12640) );
  NAND3_X1 U14948 ( .A1(n12641), .A2(n12964), .A3(n12640), .ZN(n12644) );
  NAND3_X1 U14949 ( .A1(n12644), .A2(n12642), .A3(n12953), .ZN(n12648) );
  NAND3_X1 U14950 ( .A1(n12644), .A2(n12643), .A3(n12953), .ZN(n12646) );
  NAND2_X1 U14951 ( .A1(n12952), .A2(n12962), .ZN(n12645) );
  AND2_X1 U14952 ( .A1(n12646), .A2(n12645), .ZN(n12647) );
  MUX2_X1 U14953 ( .A(n12648), .B(n12647), .S(n12657), .Z(n12656) );
  NAND2_X1 U14954 ( .A1(n12650), .A2(n12649), .ZN(n12651) );
  NAND2_X1 U14955 ( .A1(n12651), .A2(n12653), .ZN(n12652) );
  MUX2_X1 U14956 ( .A(n12653), .B(n12652), .S(n12675), .Z(n12654) );
  OAI211_X1 U14957 ( .C1(n12656), .C2(n12933), .A(n12655), .B(n12654), .ZN(
        n12661) );
  MUX2_X1 U14958 ( .A(n12659), .B(n12658), .S(n12657), .Z(n12660) );
  NAND3_X1 U14959 ( .A1(n12906), .A2(n12661), .A3(n12660), .ZN(n12665) );
  MUX2_X1 U14960 ( .A(n12663), .B(n12662), .S(n12675), .Z(n12664) );
  NAND2_X1 U14961 ( .A1(n12665), .A2(n12664), .ZN(n12666) );
  OAI21_X1 U14962 ( .B1(n12668), .B2(n12667), .A(n12674), .ZN(n12669) );
  NAND2_X1 U14963 ( .A1(n12670), .A2(n12669), .ZN(n12672) );
  OAI211_X1 U14964 ( .C1(n12673), .C2(n12675), .A(n12672), .B(n12671), .ZN(
        n12679) );
  NAND3_X1 U14965 ( .A1(n12679), .A2(n12678), .A3(n12677), .ZN(n12683) );
  INV_X1 U14966 ( .A(n12680), .ZN(n12681) );
  NAND3_X1 U14967 ( .A1(n12683), .A2(n12682), .A3(n12681), .ZN(n12685) );
  AOI21_X1 U14968 ( .B1(n6829), .B2(n12685), .A(n12684), .ZN(n12686) );
  MUX2_X1 U14969 ( .A(n15090), .B(n12687), .S(n12686), .Z(n12688) );
  NAND3_X1 U14970 ( .A1(n12693), .A2(n12692), .A3(n12824), .ZN(n12694) );
  OAI211_X1 U14971 ( .C1(n12695), .C2(n12697), .A(n12694), .B(P3_B_REG_SCAN_IN), .ZN(n12696) );
  OAI21_X1 U14972 ( .B1(n12698), .B2(n12697), .A(n12696), .ZN(P3_U3296) );
  MUX2_X1 U14973 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12699), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14974 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12700), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U14975 ( .A(n12889), .B(P3_DATAO_REG_28__SCAN_IN), .S(n12703), .Z(
        P3_U3519) );
  MUX2_X1 U14976 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12905), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14977 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12921), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14978 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12904), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14979 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12920), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14980 ( .A(n12701), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12703), .Z(
        P3_U3514) );
  MUX2_X1 U14981 ( .A(n12702), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12703), .Z(
        P3_U3513) );
  MUX2_X1 U14982 ( .A(n12988), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12703), .Z(
        P3_U3512) );
  MUX2_X1 U14983 ( .A(n13004), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12703), .Z(
        P3_U3511) );
  MUX2_X1 U14984 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n13022), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14985 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13036), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14986 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13021), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14987 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13035), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14988 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12704), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14989 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12705), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14990 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n14658), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14991 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12706), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14992 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12707), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14993 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12708), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14994 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12709), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14995 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12710), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14996 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n15073), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14997 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12711), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14998 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n15074), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14999 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12712), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15000 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n15107), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15001 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n10730), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15002 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n15108), .S(P3_U3897), .Z(
        P3_U3491) );
  AOI21_X1 U15003 ( .B1(n12714), .B2(n12716), .A(n12734), .ZN(n12732) );
  INV_X1 U15004 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12715) );
  MUX2_X1 U15005 ( .A(n12716), .B(n12715), .S(n12824), .Z(n12737) );
  XNOR2_X1 U15006 ( .A(n12737), .B(n12717), .ZN(n12721) );
  NAND2_X1 U15007 ( .A1(n12721), .A2(n12720), .ZN(n12736) );
  OAI21_X1 U15008 ( .B1(n12721), .B2(n12720), .A(n12736), .ZN(n12722) );
  NAND2_X1 U15009 ( .A1(n15052), .A2(n12722), .ZN(n12724) );
  OAI211_X1 U15010 ( .C1(n15066), .C2(n14501), .A(n12724), .B(n12723), .ZN(
        n12730) );
  AOI21_X1 U15011 ( .B1(n12715), .B2(n12727), .A(n12746), .ZN(n12728) );
  NOR2_X1 U15012 ( .A1(n12728), .A2(n15060), .ZN(n12729) );
  AOI211_X1 U15013 ( .C1(n15054), .C2(n12745), .A(n12730), .B(n12729), .ZN(
        n12731) );
  OAI21_X1 U15014 ( .B1(n12732), .B2(n15056), .A(n12731), .ZN(P3_U3195) );
  NOR2_X1 U15015 ( .A1(n12745), .A2(n12733), .ZN(n12735) );
  XNOR2_X1 U15016 ( .A(n12766), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n12738) );
  INV_X1 U15017 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14504) );
  XNOR2_X1 U15018 ( .A(n12766), .B(P3_REG1_REG_14__SCAN_IN), .ZN(n12748) );
  MUX2_X1 U15019 ( .A(n12748), .B(n12738), .S(n12846), .Z(n12739) );
  INV_X1 U15020 ( .A(n12739), .ZN(n12740) );
  OAI211_X1 U15021 ( .C1(n12741), .C2(n12740), .A(n15052), .B(n12759), .ZN(
        n12742) );
  OAI211_X1 U15022 ( .C1(n15066), .C2(n14504), .A(n12743), .B(n12742), .ZN(
        n12752) );
  NOR2_X1 U15023 ( .A1(n12745), .A2(n12744), .ZN(n12747) );
  AOI21_X1 U15024 ( .B1(n12749), .B2(n12748), .A(n12765), .ZN(n12750) );
  NOR2_X1 U15025 ( .A1(n12750), .A2(n15060), .ZN(n12751) );
  AOI211_X1 U15026 ( .C1(n15054), .C2(n12753), .A(n12752), .B(n12751), .ZN(
        n12754) );
  OAI21_X1 U15027 ( .B1(n12755), .B2(n15056), .A(n12754), .ZN(P3_U3196) );
  XNOR2_X1 U15028 ( .A(n12774), .B(n12788), .ZN(n12756) );
  INV_X1 U15029 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12760) );
  NOR2_X1 U15030 ( .A1(n12760), .A2(n12756), .ZN(n12775) );
  AOI21_X1 U15031 ( .B1(n12756), .B2(n12760), .A(n12775), .ZN(n12773) );
  MUX2_X1 U15032 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n12824), .Z(n12757) );
  NAND2_X1 U15033 ( .A1(n12757), .A2(n12766), .ZN(n12758) );
  XNOR2_X1 U15034 ( .A(n12781), .B(n12788), .ZN(n12762) );
  INV_X1 U15035 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13114) );
  MUX2_X1 U15036 ( .A(n12760), .B(n13114), .S(n12824), .Z(n12761) );
  NAND2_X1 U15037 ( .A1(n12762), .A2(n12761), .ZN(n12783) );
  OAI21_X1 U15038 ( .B1(n12762), .B2(n12761), .A(n12783), .ZN(n12771) );
  AOI21_X1 U15039 ( .B1(n15028), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n12763), 
        .ZN(n12764) );
  OAI21_X1 U15040 ( .B1(n12860), .B2(n12782), .A(n12764), .ZN(n12770) );
  AOI21_X1 U15041 ( .B1(n13114), .B2(n12767), .A(n12789), .ZN(n12768) );
  NOR2_X1 U15042 ( .A1(n12768), .A2(n15060), .ZN(n12769) );
  AOI211_X1 U15043 ( .C1(n15052), .C2(n12771), .A(n12770), .B(n12769), .ZN(
        n12772) );
  OAI21_X1 U15044 ( .B1(n12773), .B2(n15056), .A(n12772), .ZN(P3_U3197) );
  NOR2_X1 U15045 ( .A1(n12788), .A2(n12774), .ZN(n12776) );
  NAND2_X1 U15046 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12802), .ZN(n12777) );
  OAI21_X1 U15047 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n12802), .A(n12777), 
        .ZN(n12778) );
  AOI21_X1 U15048 ( .B1(n12779), .B2(n12778), .A(n12801), .ZN(n12798) );
  MUX2_X1 U15049 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12824), .Z(n12780) );
  NOR2_X1 U15050 ( .A1(n12802), .A2(n12780), .ZN(n12809) );
  AND2_X1 U15051 ( .A1(n12802), .A2(n12780), .ZN(n12808) );
  NOR2_X1 U15052 ( .A1(n12809), .A2(n12808), .ZN(n12785) );
  OR2_X1 U15053 ( .A1(n12782), .A2(n12781), .ZN(n12784) );
  XNOR2_X1 U15054 ( .A(n12785), .B(n12807), .ZN(n12796) );
  INV_X1 U15055 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n15346) );
  NOR2_X1 U15056 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15346), .ZN(n12786) );
  AOI21_X1 U15057 ( .B1(n15028), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n12786), 
        .ZN(n12787) );
  OAI21_X1 U15058 ( .B1(n12860), .B2(n12802), .A(n12787), .ZN(n12795) );
  NAND2_X1 U15059 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12802), .ZN(n12790) );
  OAI21_X1 U15060 ( .B1(P3_REG1_REG_16__SCAN_IN), .B2(n12802), .A(n12790), 
        .ZN(n12791) );
  AOI21_X1 U15061 ( .B1(n12792), .B2(n12791), .A(n12799), .ZN(n12793) );
  NOR2_X1 U15062 ( .A1(n12793), .A2(n15060), .ZN(n12794) );
  AOI211_X1 U15063 ( .C1(n15052), .C2(n12796), .A(n12795), .B(n12794), .ZN(
        n12797) );
  OAI21_X1 U15064 ( .B1(n12798), .B2(n15056), .A(n12797), .ZN(P3_U3198) );
  INV_X1 U15065 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13106) );
  AOI21_X1 U15066 ( .B1(n13106), .B2(n12800), .A(n12832), .ZN(n12812) );
  INV_X1 U15067 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12804) );
  AOI22_X1 U15068 ( .A1(n15054), .A2(n12831), .B1(n15028), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n12805) );
  MUX2_X1 U15069 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12824), .Z(n12818) );
  XOR2_X1 U15070 ( .A(n12831), .B(n12818), .Z(n12819) );
  XNOR2_X1 U15071 ( .A(n12821), .B(n12819), .ZN(n12810) );
  NAND2_X1 U15072 ( .A1(n12810), .A2(n15052), .ZN(n12811) );
  NOR2_X1 U15073 ( .A1(n12831), .A2(n12813), .ZN(n12815) );
  INV_X1 U15074 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n15345) );
  AOI22_X1 U15075 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n12839), .B1(n12850), 
        .B2(n15345), .ZN(n12816) );
  AOI21_X1 U15076 ( .B1(n6556), .B2(n12816), .A(n12843), .ZN(n12841) );
  NAND2_X1 U15077 ( .A1(n12818), .A2(n12817), .ZN(n12823) );
  INV_X1 U15078 ( .A(n12819), .ZN(n12820) );
  NAND2_X1 U15079 ( .A1(n12821), .A2(n12820), .ZN(n12822) );
  NAND2_X1 U15080 ( .A1(n12823), .A2(n12822), .ZN(n12849) );
  XNOR2_X1 U15081 ( .A(n12850), .B(n12849), .ZN(n12826) );
  MUX2_X1 U15082 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12824), .Z(n12825) );
  NOR2_X1 U15083 ( .A1(n12826), .A2(n12825), .ZN(n12852) );
  AOI21_X1 U15084 ( .B1(n12826), .B2(n12825), .A(n12852), .ZN(n12829) );
  NAND2_X1 U15085 ( .A1(n15028), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n12827) );
  OAI211_X1 U15086 ( .C1(n12829), .C2(n12855), .A(n12828), .B(n12827), .ZN(
        n12838) );
  INV_X1 U15087 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12834) );
  AOI22_X1 U15088 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n12839), .B1(n12850), 
        .B2(n12834), .ZN(n12835) );
  AOI21_X1 U15089 ( .B1(n6728), .B2(n12836), .A(n15060), .ZN(n12837) );
  AOI211_X1 U15090 ( .C1(n15054), .C2(n12839), .A(n12838), .B(n12837), .ZN(
        n12840) );
  OAI21_X1 U15091 ( .B1(n12841), .B2(n15056), .A(n12840), .ZN(P3_U3200) );
  INV_X1 U15092 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12842) );
  MUX2_X1 U15093 ( .A(n12842), .B(P3_REG2_REG_19__SCAN_IN), .S(n12859), .Z(
        n12847) );
  AOI21_X1 U15094 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n12850), .A(n12843), 
        .ZN(n12844) );
  XOR2_X1 U15095 ( .A(n12847), .B(n12844), .Z(n12864) );
  XNOR2_X1 U15096 ( .A(n12859), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12848) );
  MUX2_X1 U15097 ( .A(n12848), .B(n12847), .S(n12846), .Z(n12854) );
  NOR2_X1 U15098 ( .A1(n12850), .A2(n12849), .ZN(n12851) );
  XOR2_X1 U15099 ( .A(n12854), .B(n12853), .Z(n12856) );
  NAND2_X1 U15100 ( .A1(n15028), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12857) );
  OAI211_X1 U15101 ( .C1(n12860), .C2(n12859), .A(n12858), .B(n12857), .ZN(
        n12861) );
  OAI21_X1 U15102 ( .B1(n12864), .B2(n15056), .A(n12863), .ZN(P3_U3201) );
  INV_X1 U15103 ( .A(n13117), .ZN(n13049) );
  NAND2_X1 U15104 ( .A1(n12872), .A2(n15119), .ZN(n12867) );
  OR2_X1 U15105 ( .A1(n12866), .A2(n12865), .ZN(n13118) );
  AOI21_X1 U15106 ( .B1(n12867), .B2(n13118), .A(n15124), .ZN(n12869) );
  AOI21_X1 U15107 ( .B1(n15124), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12869), 
        .ZN(n12868) );
  OAI21_X1 U15108 ( .B1(n13049), .B2(n13044), .A(n12868), .ZN(P3_U3202) );
  AOI21_X1 U15109 ( .B1(n15124), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12869), 
        .ZN(n12870) );
  OAI21_X1 U15110 ( .B1(n13052), .B2(n13044), .A(n12870), .ZN(P3_U3203) );
  INV_X1 U15111 ( .A(n12871), .ZN(n12878) );
  AOI22_X1 U15112 ( .A1(n12872), .A2(n15119), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n15124), .ZN(n12873) );
  OAI21_X1 U15113 ( .B1(n12874), .B2(n13044), .A(n12873), .ZN(n12875) );
  AOI21_X1 U15114 ( .B1(n12876), .B2(n14664), .A(n12875), .ZN(n12877) );
  OAI21_X1 U15115 ( .B1(n12878), .B2(n15124), .A(n12877), .ZN(P3_U3204) );
  INV_X1 U15116 ( .A(n12879), .ZN(n12885) );
  AOI22_X1 U15117 ( .A1(n12880), .A2(n15119), .B1(n15124), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12881) );
  OAI21_X1 U15118 ( .B1(n13056), .B2(n13044), .A(n12881), .ZN(n12882) );
  AOI21_X1 U15119 ( .B1(n12883), .B2(n15122), .A(n12882), .ZN(n12884) );
  OAI21_X1 U15120 ( .B1(n12885), .B2(n12998), .A(n12884), .ZN(P3_U3205) );
  INV_X1 U15121 ( .A(n12886), .ZN(n12887) );
  AOI21_X1 U15122 ( .B1(n12890), .B2(n12888), .A(n12887), .ZN(n12896) );
  AOI22_X1 U15123 ( .A1(n12889), .A2(n15106), .B1(n15109), .B2(n12921), .ZN(
        n12895) );
  NOR2_X1 U15124 ( .A1(n12891), .A2(n12890), .ZN(n12892) );
  NAND2_X1 U15125 ( .A1(n13058), .A2(n15075), .ZN(n12894) );
  OAI211_X1 U15126 ( .C1(n12896), .C2(n15078), .A(n12895), .B(n12894), .ZN(
        n13057) );
  NAND2_X1 U15127 ( .A1(n13058), .A2(n15120), .ZN(n12899) );
  AOI22_X1 U15128 ( .A1(n12897), .A2(n15119), .B1(n15124), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12898) );
  OAI211_X1 U15129 ( .C1(n13129), .C2(n13044), .A(n12899), .B(n12898), .ZN(
        n12900) );
  AOI21_X1 U15130 ( .B1(n13057), .B2(n15122), .A(n12900), .ZN(n12901) );
  INV_X1 U15131 ( .A(n12901), .ZN(P3_U3206) );
  XNOR2_X1 U15132 ( .A(n12903), .B(n12902), .ZN(n12910) );
  AOI22_X1 U15133 ( .A1(n12905), .A2(n15106), .B1(n15109), .B2(n12904), .ZN(
        n12909) );
  XNOR2_X1 U15134 ( .A(n12906), .B(n12907), .ZN(n13062) );
  NAND2_X1 U15135 ( .A1(n13062), .A2(n15075), .ZN(n12908) );
  OAI211_X1 U15136 ( .C1(n12910), .C2(n15078), .A(n12909), .B(n12908), .ZN(
        n13061) );
  NAND2_X1 U15137 ( .A1(n13062), .A2(n15120), .ZN(n12913) );
  AOI22_X1 U15138 ( .A1(n12911), .A2(n15119), .B1(n15124), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12912) );
  OAI211_X1 U15139 ( .C1(n13133), .C2(n13044), .A(n12913), .B(n12912), .ZN(
        n12914) );
  AOI21_X1 U15140 ( .B1(n13061), .B2(n15122), .A(n12914), .ZN(n12915) );
  INV_X1 U15141 ( .A(n12915), .ZN(P3_U3207) );
  XNOR2_X1 U15142 ( .A(n12916), .B(n12918), .ZN(n13068) );
  OAI211_X1 U15143 ( .C1(n12919), .C2(n12918), .A(n12917), .B(n15112), .ZN(
        n12923) );
  AOI22_X1 U15144 ( .A1(n12921), .A2(n15106), .B1(n15109), .B2(n12920), .ZN(
        n12922) );
  NAND2_X1 U15145 ( .A1(n12923), .A2(n12922), .ZN(n13065) );
  AOI22_X1 U15146 ( .A1(n12924), .A2(n15119), .B1(n15124), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12925) );
  OAI21_X1 U15147 ( .B1(n12926), .B2(n13044), .A(n12925), .ZN(n12927) );
  AOI21_X1 U15148 ( .B1(n13065), .B2(n15122), .A(n12927), .ZN(n12928) );
  OAI21_X1 U15149 ( .B1(n12998), .B2(n13068), .A(n12928), .ZN(P3_U3208) );
  NAND2_X1 U15150 ( .A1(n12929), .A2(n12933), .ZN(n12930) );
  OAI21_X1 U15151 ( .B1(n12934), .B2(n12933), .A(n12932), .ZN(n12935) );
  NAND2_X1 U15152 ( .A1(n12935), .A2(n15112), .ZN(n12939) );
  OAI22_X1 U15153 ( .A1(n12936), .A2(n15095), .B1(n12962), .B2(n15094), .ZN(
        n12937) );
  INV_X1 U15154 ( .A(n12937), .ZN(n12938) );
  OAI211_X1 U15155 ( .C1(n15116), .C2(n13069), .A(n12939), .B(n12938), .ZN(
        n13074) );
  AOI22_X1 U15156 ( .A1(n12940), .A2(n15119), .B1(n15124), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12943) );
  NAND2_X1 U15157 ( .A1(n12941), .A2(n13027), .ZN(n12942) );
  OAI211_X1 U15158 ( .C1(n13069), .C2(n12944), .A(n12943), .B(n12942), .ZN(
        n12945) );
  AOI21_X1 U15159 ( .B1(n13074), .B2(n15122), .A(n12945), .ZN(n12946) );
  INV_X1 U15160 ( .A(n12946), .ZN(P3_U3209) );
  AOI21_X1 U15161 ( .B1(n12947), .B2(n12953), .A(n15078), .ZN(n12951) );
  OAI22_X1 U15162 ( .A1(n12948), .A2(n15095), .B1(n12975), .B2(n15094), .ZN(
        n12949) );
  AOI21_X1 U15163 ( .B1(n12951), .B2(n12950), .A(n12949), .ZN(n13080) );
  NOR2_X1 U15164 ( .A1(n13080), .A2(n15124), .ZN(n12959) );
  INV_X1 U15165 ( .A(n12952), .ZN(n13081) );
  OR2_X1 U15166 ( .A1(n12954), .A2(n12953), .ZN(n13078) );
  NAND3_X1 U15167 ( .A1(n13078), .A2(n13077), .A3(n14664), .ZN(n12957) );
  AOI22_X1 U15168 ( .A1(n12955), .A2(n15119), .B1(n15124), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n12956) );
  OAI211_X1 U15169 ( .C1(n13081), .C2(n13044), .A(n12957), .B(n12956), .ZN(
        n12958) );
  OR2_X1 U15170 ( .A1(n12959), .A2(n12958), .ZN(P3_U3210) );
  XNOR2_X1 U15171 ( .A(n12960), .B(n12964), .ZN(n12961) );
  OAI222_X1 U15172 ( .A1(n15094), .A2(n12963), .B1(n15095), .B2(n12962), .C1(
        n15078), .C2(n12961), .ZN(n13082) );
  INV_X1 U15173 ( .A(n13082), .ZN(n12971) );
  XOR2_X1 U15174 ( .A(n12965), .B(n12964), .Z(n13083) );
  INV_X1 U15175 ( .A(n12966), .ZN(n13142) );
  AOI22_X1 U15176 ( .A1(n15124), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n12967), 
        .B2(n15119), .ZN(n12968) );
  OAI21_X1 U15177 ( .B1(n13142), .B2(n13044), .A(n12968), .ZN(n12969) );
  AOI21_X1 U15178 ( .B1(n13083), .B2(n14664), .A(n12969), .ZN(n12970) );
  OAI21_X1 U15179 ( .B1(n12971), .B2(n15124), .A(n12970), .ZN(P3_U3211) );
  XOR2_X1 U15180 ( .A(n12972), .B(n12976), .Z(n12973) );
  OAI222_X1 U15181 ( .A1(n15095), .A2(n12975), .B1(n15094), .B2(n12974), .C1(
        n15078), .C2(n12973), .ZN(n13086) );
  INV_X1 U15182 ( .A(n13086), .ZN(n12982) );
  XOR2_X1 U15183 ( .A(n12977), .B(n12976), .Z(n13087) );
  AOI22_X1 U15184 ( .A1(n15124), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15119), 
        .B2(n12978), .ZN(n12979) );
  OAI21_X1 U15185 ( .B1(n13146), .B2(n13044), .A(n12979), .ZN(n12980) );
  AOI21_X1 U15186 ( .B1(n13087), .B2(n14664), .A(n12980), .ZN(n12981) );
  OAI21_X1 U15187 ( .B1(n12982), .B2(n15124), .A(n12981), .ZN(P3_U3212) );
  NOR2_X1 U15188 ( .A1(n13018), .A2(n12983), .ZN(n13002) );
  OR2_X1 U15189 ( .A1(n13002), .A2(n12984), .ZN(n13001) );
  NAND3_X1 U15190 ( .A1(n13001), .A2(n12985), .A3(n6497), .ZN(n12987) );
  NAND3_X1 U15191 ( .A1(n12987), .A2(n15112), .A3(n12986), .ZN(n12990) );
  AOI22_X1 U15192 ( .A1(n12988), .A2(n15106), .B1(n15109), .B2(n13022), .ZN(
        n12989) );
  AND2_X1 U15193 ( .A1(n12990), .A2(n12989), .ZN(n13092) );
  NAND2_X1 U15194 ( .A1(n12992), .A2(n12991), .ZN(n12993) );
  NAND2_X1 U15195 ( .A1(n12994), .A2(n12993), .ZN(n13093) );
  AOI22_X1 U15196 ( .A1(n15124), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15119), 
        .B2(n12995), .ZN(n12997) );
  NAND2_X1 U15197 ( .A1(n13090), .A2(n13027), .ZN(n12996) );
  OAI211_X1 U15198 ( .C1(n13093), .C2(n12998), .A(n12997), .B(n12996), .ZN(
        n12999) );
  INV_X1 U15199 ( .A(n12999), .ZN(n13000) );
  OAI21_X1 U15200 ( .B1(n13092), .B2(n15124), .A(n13000), .ZN(P3_U3213) );
  NAND2_X1 U15201 ( .A1(n13001), .A2(n15112), .ZN(n13007) );
  INV_X1 U15202 ( .A(n13002), .ZN(n13019) );
  AOI21_X1 U15203 ( .B1(n13019), .B2(n13003), .A(n13008), .ZN(n13006) );
  AOI22_X1 U15204 ( .A1(n13004), .A2(n15106), .B1(n15109), .B2(n13036), .ZN(
        n13005) );
  OAI21_X1 U15205 ( .B1(n13007), .B2(n13006), .A(n13005), .ZN(n13094) );
  INV_X1 U15206 ( .A(n13094), .ZN(n13017) );
  INV_X1 U15207 ( .A(n13100), .ZN(n13010) );
  OAI21_X1 U15208 ( .B1(n13010), .B2(n13009), .A(n13008), .ZN(n13012) );
  NAND2_X1 U15209 ( .A1(n13012), .A2(n13011), .ZN(n13095) );
  AOI22_X1 U15210 ( .A1(n15124), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15119), 
        .B2(n13013), .ZN(n13014) );
  OAI21_X1 U15211 ( .B1(n13151), .B2(n13044), .A(n13014), .ZN(n13015) );
  AOI21_X1 U15212 ( .B1(n13095), .B2(n14664), .A(n13015), .ZN(n13016) );
  OAI21_X1 U15213 ( .B1(n13017), .B2(n15124), .A(n13016), .ZN(P3_U3214) );
  INV_X1 U15214 ( .A(n13018), .ZN(n13020) );
  OAI21_X1 U15215 ( .B1(n13020), .B2(n13028), .A(n13019), .ZN(n13023) );
  AOI222_X1 U15216 ( .A1(n15112), .A2(n13023), .B1(n13022), .B2(n15106), .C1(
        n13021), .C2(n15109), .ZN(n13102) );
  INV_X1 U15217 ( .A(n13024), .ZN(n13025) );
  OAI22_X1 U15218 ( .A1(n15122), .A2(n15345), .B1(n13025), .B2(n15089), .ZN(
        n13026) );
  AOI21_X1 U15219 ( .B1(n13098), .B2(n13027), .A(n13026), .ZN(n13031) );
  NAND2_X1 U15220 ( .A1(n13029), .A2(n13028), .ZN(n13099) );
  NAND3_X1 U15221 ( .A1(n13100), .A2(n14664), .A3(n13099), .ZN(n13030) );
  OAI211_X1 U15222 ( .C1(n13102), .C2(n15124), .A(n13031), .B(n13030), .ZN(
        P3_U3215) );
  OAI211_X1 U15223 ( .C1(n13034), .C2(n13033), .A(n13032), .B(n15112), .ZN(
        n13038) );
  AOI22_X1 U15224 ( .A1(n13036), .A2(n15106), .B1(n15109), .B2(n13035), .ZN(
        n13037) );
  NAND2_X1 U15225 ( .A1(n13038), .A2(n13037), .ZN(n13104) );
  INV_X1 U15226 ( .A(n13104), .ZN(n13047) );
  XNOR2_X1 U15227 ( .A(n13040), .B(n13039), .ZN(n13105) );
  INV_X1 U15228 ( .A(n13041), .ZN(n13155) );
  AOI22_X1 U15229 ( .A1(n15124), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15119), 
        .B2(n13042), .ZN(n13043) );
  OAI21_X1 U15230 ( .B1(n13155), .B2(n13044), .A(n13043), .ZN(n13045) );
  AOI21_X1 U15231 ( .B1(n13105), .B2(n14664), .A(n13045), .ZN(n13046) );
  OAI21_X1 U15232 ( .B1(n13047), .B2(n15124), .A(n13046), .ZN(P3_U3216) );
  NOR2_X1 U15233 ( .A1(n13118), .A2(n15190), .ZN(n13050) );
  AOI21_X1 U15234 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n15190), .A(n13050), 
        .ZN(n13048) );
  OAI21_X1 U15235 ( .B1(n13049), .B2(n13116), .A(n13048), .ZN(P3_U3490) );
  AOI21_X1 U15236 ( .B1(P3_REG1_REG_30__SCAN_IN), .B2(n15190), .A(n13050), 
        .ZN(n13051) );
  OAI21_X1 U15237 ( .B1(n13052), .B2(n13116), .A(n13051), .ZN(P3_U3489) );
  INV_X1 U15238 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13054) );
  MUX2_X1 U15239 ( .A(n13054), .B(n13053), .S(n15193), .Z(n13055) );
  OAI21_X1 U15240 ( .B1(n13056), .B2(n13116), .A(n13055), .ZN(P3_U3487) );
  INV_X1 U15241 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13059) );
  AOI21_X1 U15242 ( .B1(n15166), .B2(n13058), .A(n13057), .ZN(n13126) );
  MUX2_X1 U15243 ( .A(n13059), .B(n13126), .S(n15193), .Z(n13060) );
  OAI21_X1 U15244 ( .B1(n13129), .B2(n13116), .A(n13060), .ZN(P3_U3486) );
  INV_X1 U15245 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13063) );
  AOI21_X1 U15246 ( .B1(n15166), .B2(n13062), .A(n13061), .ZN(n13130) );
  MUX2_X1 U15247 ( .A(n13063), .B(n13130), .S(n15193), .Z(n13064) );
  OAI21_X1 U15248 ( .B1(n13133), .B2(n13116), .A(n13064), .ZN(P3_U3485) );
  INV_X1 U15249 ( .A(n14692), .ZN(n15170) );
  AOI21_X1 U15250 ( .B1(n15080), .B2(n13066), .A(n13065), .ZN(n13067) );
  OAI21_X1 U15251 ( .B1(n15170), .B2(n13068), .A(n13067), .ZN(n13134) );
  MUX2_X1 U15252 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13134), .S(n15193), .Z(
        P3_U3484) );
  INV_X1 U15253 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13075) );
  INV_X1 U15254 ( .A(n13069), .ZN(n13070) );
  NAND2_X1 U15255 ( .A1(n13070), .A2(n15166), .ZN(n13071) );
  OAI21_X1 U15256 ( .B1(n13072), .B2(n15169), .A(n13071), .ZN(n13073) );
  NOR2_X1 U15257 ( .A1(n13074), .A2(n13073), .ZN(n13135) );
  MUX2_X1 U15258 ( .A(n13075), .B(n13135), .S(n15193), .Z(n13076) );
  INV_X1 U15259 ( .A(n13076), .ZN(P3_U3483) );
  NAND3_X1 U15260 ( .A1(n13078), .A2(n13077), .A3(n14692), .ZN(n13079) );
  OAI211_X1 U15261 ( .C1(n13081), .C2(n15169), .A(n13080), .B(n13079), .ZN(
        n13138) );
  MUX2_X1 U15262 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n13138), .S(n15193), .Z(
        P3_U3482) );
  INV_X1 U15263 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13084) );
  AOI21_X1 U15264 ( .B1(n14692), .B2(n13083), .A(n13082), .ZN(n13139) );
  MUX2_X1 U15265 ( .A(n13084), .B(n13139), .S(n15193), .Z(n13085) );
  OAI21_X1 U15266 ( .B1(n13142), .B2(n13116), .A(n13085), .ZN(P3_U3481) );
  INV_X1 U15267 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13088) );
  AOI21_X1 U15268 ( .B1(n13087), .B2(n14692), .A(n13086), .ZN(n13143) );
  MUX2_X1 U15269 ( .A(n13088), .B(n13143), .S(n15193), .Z(n13089) );
  OAI21_X1 U15270 ( .B1(n13146), .B2(n13116), .A(n13089), .ZN(P3_U3480) );
  NAND2_X1 U15271 ( .A1(n13090), .A2(n15080), .ZN(n13091) );
  OAI211_X1 U15272 ( .C1(n15170), .C2(n13093), .A(n13092), .B(n13091), .ZN(
        n13147) );
  MUX2_X1 U15273 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n13147), .S(n15193), .Z(
        P3_U3479) );
  INV_X1 U15274 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13096) );
  AOI21_X1 U15275 ( .B1(n14692), .B2(n13095), .A(n13094), .ZN(n13148) );
  MUX2_X1 U15276 ( .A(n13096), .B(n13148), .S(n15193), .Z(n13097) );
  OAI21_X1 U15277 ( .B1(n13116), .B2(n13151), .A(n13097), .ZN(P3_U3478) );
  INV_X1 U15278 ( .A(n13098), .ZN(n13103) );
  NAND3_X1 U15279 ( .A1(n13100), .A2(n14692), .A3(n13099), .ZN(n13101) );
  OAI211_X1 U15280 ( .C1(n13103), .C2(n15169), .A(n13102), .B(n13101), .ZN(
        n13152) );
  MUX2_X1 U15281 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n13152), .S(n15193), .Z(
        P3_U3477) );
  AOI21_X1 U15282 ( .B1(n13105), .B2(n14692), .A(n13104), .ZN(n13153) );
  MUX2_X1 U15283 ( .A(n13106), .B(n13153), .S(n15193), .Z(n13107) );
  OAI21_X1 U15284 ( .B1(n13155), .B2(n13116), .A(n13107), .ZN(P3_U3476) );
  INV_X1 U15285 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13110) );
  AOI21_X1 U15286 ( .B1(n13109), .B2(n14692), .A(n13108), .ZN(n13156) );
  MUX2_X1 U15287 ( .A(n13110), .B(n13156), .S(n15193), .Z(n13111) );
  OAI21_X1 U15288 ( .B1(n13158), .B2(n13116), .A(n13111), .ZN(P3_U3475) );
  AOI21_X1 U15289 ( .B1(n13113), .B2(n14692), .A(n13112), .ZN(n13159) );
  MUX2_X1 U15290 ( .A(n13114), .B(n13159), .S(n15193), .Z(n13115) );
  OAI21_X1 U15291 ( .B1(n13163), .B2(n13116), .A(n13115), .ZN(P3_U3474) );
  INV_X1 U15292 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n13121) );
  NAND2_X1 U15293 ( .A1(n13117), .A2(n8837), .ZN(n13120) );
  INV_X1 U15294 ( .A(n13118), .ZN(n13119) );
  NAND2_X1 U15295 ( .A1(n13119), .A2(n15176), .ZN(n13123) );
  OAI211_X1 U15296 ( .C1(n15176), .C2(n13121), .A(n13120), .B(n13123), .ZN(
        P3_U3458) );
  INV_X1 U15297 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n13125) );
  NAND2_X1 U15298 ( .A1(n13122), .A2(n8837), .ZN(n13124) );
  OAI211_X1 U15299 ( .C1(n15176), .C2(n13125), .A(n13124), .B(n13123), .ZN(
        P3_U3457) );
  INV_X1 U15300 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13127) );
  MUX2_X1 U15301 ( .A(n13127), .B(n13126), .S(n15176), .Z(n13128) );
  OAI21_X1 U15302 ( .B1(n13129), .B2(n13162), .A(n13128), .ZN(P3_U3454) );
  INV_X1 U15303 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13131) );
  MUX2_X1 U15304 ( .A(n13131), .B(n13130), .S(n15176), .Z(n13132) );
  OAI21_X1 U15305 ( .B1(n13133), .B2(n13162), .A(n13132), .ZN(P3_U3453) );
  MUX2_X1 U15306 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n13134), .S(n15176), .Z(
        P3_U3452) );
  INV_X1 U15307 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13136) );
  MUX2_X1 U15308 ( .A(n13136), .B(n13135), .S(n15176), .Z(n13137) );
  INV_X1 U15309 ( .A(n13137), .ZN(P3_U3451) );
  MUX2_X1 U15310 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n13138), .S(n15176), .Z(
        P3_U3450) );
  INV_X1 U15311 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13140) );
  MUX2_X1 U15312 ( .A(n13140), .B(n13139), .S(n15176), .Z(n13141) );
  OAI21_X1 U15313 ( .B1(n13142), .B2(n13162), .A(n13141), .ZN(P3_U3449) );
  INV_X1 U15314 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13144) );
  MUX2_X1 U15315 ( .A(n13144), .B(n13143), .S(n15176), .Z(n13145) );
  OAI21_X1 U15316 ( .B1(n13146), .B2(n13162), .A(n13145), .ZN(P3_U3448) );
  MUX2_X1 U15317 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n13147), .S(n15176), .Z(
        P3_U3447) );
  MUX2_X1 U15318 ( .A(n13149), .B(n13148), .S(n15176), .Z(n13150) );
  OAI21_X1 U15319 ( .B1(n13162), .B2(n13151), .A(n13150), .ZN(P3_U3446) );
  MUX2_X1 U15320 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n13152), .S(n15176), .Z(
        P3_U3444) );
  MUX2_X1 U15321 ( .A(n15334), .B(n13153), .S(n15176), .Z(n13154) );
  OAI21_X1 U15322 ( .B1(n13155), .B2(n13162), .A(n13154), .ZN(P3_U3441) );
  INV_X1 U15323 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n15237) );
  MUX2_X1 U15324 ( .A(n15237), .B(n13156), .S(n15176), .Z(n13157) );
  OAI21_X1 U15325 ( .B1(n13158), .B2(n13162), .A(n13157), .ZN(P3_U3438) );
  INV_X1 U15326 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13160) );
  MUX2_X1 U15327 ( .A(n13160), .B(n13159), .S(n15176), .Z(n13161) );
  OAI21_X1 U15328 ( .B1(n13163), .B2(n13162), .A(n13161), .ZN(P3_U3435) );
  MUX2_X1 U15329 ( .A(P3_D_REG_1__SCAN_IN), .B(n13164), .S(n13165), .Z(
        P3_U3377) );
  MUX2_X1 U15330 ( .A(P3_D_REG_0__SCAN_IN), .B(n13166), .S(n13165), .Z(
        P3_U3376) );
  INV_X1 U15331 ( .A(n13167), .ZN(n13172) );
  NOR4_X1 U15332 ( .A1(n13168), .A2(P3_IR_REG_30__SCAN_IN), .A3(n8273), .A4(
        P3_U3151), .ZN(n13169) );
  AOI21_X1 U15333 ( .B1(n13170), .B2(SI_31_), .A(n13169), .ZN(n13171) );
  OAI21_X1 U15334 ( .B1(n13172), .B2(n13175), .A(n13171), .ZN(P3_U3264) );
  INV_X1 U15335 ( .A(n13173), .ZN(n13174) );
  NAND2_X1 U15336 ( .A1(n13180), .A2(n13179), .ZN(n13181) );
  NAND3_X1 U15337 ( .A1(n13182), .A2(n14860), .A3(n13181), .ZN(n13188) );
  OR2_X1 U15338 ( .A1(n13444), .A2(n13596), .ZN(n13184) );
  NAND2_X1 U15339 ( .A1(n13438), .A2(n13576), .ZN(n13183) );
  NAND2_X1 U15340 ( .A1(n13184), .A2(n13183), .ZN(n13470) );
  AOI22_X1 U15341 ( .A1(n13238), .A2(n13470), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13185) );
  OAI21_X1 U15342 ( .B1(n13472), .B2(n14870), .A(n13185), .ZN(n13186) );
  AOI21_X1 U15343 ( .B1(n7100), .B2(n14867), .A(n13186), .ZN(n13187) );
  NAND2_X1 U15344 ( .A1(n13188), .A2(n13187), .ZN(P2_U3186) );
  AOI22_X1 U15345 ( .A1(n13190), .A2(n14860), .B1(n13189), .B2(n13520), .ZN(
        n13198) );
  INV_X1 U15346 ( .A(n13191), .ZN(n13197) );
  NAND2_X1 U15347 ( .A1(n13406), .A2(n13576), .ZN(n13193) );
  NAND2_X1 U15348 ( .A1(n13412), .A2(n15413), .ZN(n13192) );
  NAND2_X1 U15349 ( .A1(n13193), .A2(n13192), .ZN(n13694) );
  AOI22_X1 U15350 ( .A1(n13238), .A2(n13694), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13194) );
  OAI21_X1 U15351 ( .B1(n13542), .B2(n14870), .A(n13194), .ZN(n13195) );
  AOI21_X1 U15352 ( .B1(n13695), .B2(n14867), .A(n13195), .ZN(n13196) );
  OAI21_X1 U15353 ( .B1(n13198), .B2(n13197), .A(n13196), .ZN(P2_U3188) );
  OAI21_X1 U15354 ( .B1(n13272), .B2(n13200), .A(n13264), .ZN(n13208) );
  NOR3_X1 U15355 ( .A1(n13200), .A2(n13199), .A3(n8233), .ZN(n13201) );
  OAI21_X1 U15356 ( .B1(n13201), .B2(n13289), .A(n13396), .ZN(n13206) );
  INV_X1 U15357 ( .A(n13202), .ZN(n13604) );
  INV_X1 U15358 ( .A(n13401), .ZN(n13597) );
  OAI21_X1 U15359 ( .B1(n13597), .B2(n13254), .A(n13203), .ZN(n13204) );
  AOI21_X1 U15360 ( .B1(n13604), .B2(n13277), .A(n13204), .ZN(n13205) );
  OAI211_X1 U15361 ( .C1(n7109), .C2(n13281), .A(n13206), .B(n13205), .ZN(
        n13207) );
  AOI21_X1 U15362 ( .B1(n14860), .B2(n13208), .A(n13207), .ZN(n13209) );
  INV_X1 U15363 ( .A(n13209), .ZN(P2_U3191) );
  OAI211_X1 U15364 ( .C1(n6626), .C2(n13211), .A(n13210), .B(n14860), .ZN(
        n13215) );
  AOI22_X1 U15365 ( .A1(n13401), .A2(n13289), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13212) );
  OAI21_X1 U15366 ( .B1(n13563), .B2(n13254), .A(n13212), .ZN(n13213) );
  AOI21_X1 U15367 ( .B1(n13569), .B2(n13277), .A(n13213), .ZN(n13214) );
  OAI211_X1 U15368 ( .C1(n7107), .C2(n13281), .A(n13215), .B(n13214), .ZN(
        P2_U3195) );
  OAI21_X1 U15369 ( .B1(n11503), .B2(n13223), .A(n13216), .ZN(n13217) );
  NAND2_X1 U15370 ( .A1(n13217), .A2(n14860), .ZN(n13227) );
  AOI22_X1 U15371 ( .A1(n13284), .A2(n13300), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13218) );
  OAI21_X1 U15372 ( .B1(n13219), .B2(n14870), .A(n13218), .ZN(n13220) );
  AOI21_X1 U15373 ( .B1(n13221), .B2(n14867), .A(n13220), .ZN(n13226) );
  NOR3_X1 U15374 ( .A1(n13223), .A2(n13222), .A3(n8233), .ZN(n13224) );
  OAI21_X1 U15375 ( .B1(n13224), .B2(n13289), .A(n13302), .ZN(n13225) );
  NAND3_X1 U15376 ( .A1(n13227), .A2(n13226), .A3(n13225), .ZN(P2_U3196) );
  INV_X1 U15377 ( .A(n13245), .ZN(n13228) );
  AOI21_X1 U15378 ( .B1(n13230), .B2(n13229), .A(n13228), .ZN(n13237) );
  NOR2_X1 U15379 ( .A1(n14870), .A2(n13231), .ZN(n13235) );
  OAI22_X1 U15380 ( .A1(n13233), .A2(n14859), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13232), .ZN(n13234) );
  AOI211_X1 U15381 ( .C1(n13419), .C2(n14867), .A(n13235), .B(n13234), .ZN(
        n13236) );
  OAI21_X1 U15382 ( .B1(n13237), .B2(n13269), .A(n13236), .ZN(P2_U3198) );
  OAI22_X1 U15383 ( .A1(n13595), .A2(n13596), .B1(n13418), .B2(n13594), .ZN(
        n13630) );
  AOI22_X1 U15384 ( .A1(n13630), .A2(n13238), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13239) );
  OAI21_X1 U15385 ( .B1(n13636), .B2(n14870), .A(n13239), .ZN(n13240) );
  AOI21_X1 U15386 ( .B1(n13727), .B2(n14867), .A(n13240), .ZN(n13247) );
  INV_X1 U15387 ( .A(n13241), .ZN(n13244) );
  OAI22_X1 U15388 ( .A1(n13242), .A2(n13269), .B1(n13418), .B2(n8233), .ZN(
        n13243) );
  NAND3_X1 U15389 ( .A1(n13245), .A2(n13244), .A3(n13243), .ZN(n13246) );
  OAI211_X1 U15390 ( .C1(n13248), .C2(n13269), .A(n13247), .B(n13246), .ZN(
        P2_U3200) );
  INV_X1 U15391 ( .A(n13688), .ZN(n13527) );
  OAI211_X1 U15392 ( .C1(n13251), .C2(n13250), .A(n13249), .B(n14860), .ZN(
        n13257) );
  INV_X1 U15393 ( .A(n13252), .ZN(n13525) );
  AOI22_X1 U15394 ( .A1(n13289), .A2(n13520), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13253) );
  OAI21_X1 U15395 ( .B1(n13485), .B2(n13254), .A(n13253), .ZN(n13255) );
  AOI21_X1 U15396 ( .B1(n13525), .B2(n13277), .A(n13255), .ZN(n13256) );
  OAI211_X1 U15397 ( .C1(n13527), .C2(n13281), .A(n13257), .B(n13256), .ZN(
        P2_U3201) );
  INV_X1 U15398 ( .A(n13258), .ZN(n13268) );
  NAND2_X1 U15399 ( .A1(n13579), .A2(n13284), .ZN(n13260) );
  AOI22_X1 U15400 ( .A1(n13289), .A2(n13577), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13259) );
  OAI211_X1 U15401 ( .C1(n14870), .C2(n13582), .A(n13260), .B(n13259), .ZN(
        n13261) );
  AOI21_X1 U15402 ( .B1(n13710), .B2(n14867), .A(n13261), .ZN(n13267) );
  INV_X1 U15403 ( .A(n13577), .ZN(n13425) );
  OAI22_X1 U15404 ( .A1(n13262), .A2(n13269), .B1(n13425), .B2(n8233), .ZN(
        n13263) );
  NAND3_X1 U15405 ( .A1(n13265), .A2(n13264), .A3(n13263), .ZN(n13266) );
  OAI211_X1 U15406 ( .C1(n13268), .C2(n13269), .A(n13267), .B(n13266), .ZN(
        P2_U3205) );
  INV_X1 U15407 ( .A(n13625), .ZN(n13723) );
  AOI21_X1 U15408 ( .B1(n13271), .B2(n13270), .A(n13269), .ZN(n13273) );
  NAND2_X1 U15409 ( .A1(n13273), .A2(n13272), .ZN(n13280) );
  INV_X1 U15410 ( .A(n13619), .ZN(n13278) );
  AND2_X1 U15411 ( .A1(n13394), .A2(n13576), .ZN(n13274) );
  AOI21_X1 U15412 ( .B1(n13577), .B2(n15413), .A(n13274), .ZN(n13617) );
  OAI21_X1 U15413 ( .B1(n13617), .B2(n14859), .A(n13275), .ZN(n13276) );
  AOI21_X1 U15414 ( .B1(n13278), .B2(n13277), .A(n13276), .ZN(n13279) );
  OAI211_X1 U15415 ( .C1(n13723), .C2(n13281), .A(n13280), .B(n13279), .ZN(
        P2_U3210) );
  OAI21_X1 U15416 ( .B1(n13287), .B2(n12269), .A(n13282), .ZN(n13283) );
  NAND2_X1 U15417 ( .A1(n13283), .A2(n14860), .ZN(n13293) );
  AOI22_X1 U15418 ( .A1(n13284), .A2(n13297), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13285) );
  OAI21_X1 U15419 ( .B1(n13492), .B2(n14870), .A(n13285), .ZN(n13286) );
  AOI21_X1 U15420 ( .B1(n13495), .B2(n14867), .A(n13286), .ZN(n13292) );
  NOR3_X1 U15421 ( .A1(n13288), .A2(n13287), .A3(n8233), .ZN(n13290) );
  OAI21_X1 U15422 ( .B1(n13290), .B2(n13289), .A(n6840), .ZN(n13291) );
  NAND3_X1 U15423 ( .A1(n13293), .A2(n13292), .A3(n13291), .ZN(P2_U3212) );
  MUX2_X1 U15424 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13384), .S(n14856), .Z(
        P2_U3562) );
  MUX2_X1 U15425 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13294), .S(n14856), .Z(
        P2_U3561) );
  MUX2_X1 U15426 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13295), .S(n14856), .Z(
        P2_U3560) );
  MUX2_X1 U15427 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13296), .S(n14856), .Z(
        P2_U3559) );
  MUX2_X1 U15428 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13297), .S(n14856), .Z(
        P2_U3558) );
  MUX2_X1 U15429 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13438), .S(n14856), .Z(
        P2_U3557) );
  MUX2_X1 U15430 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n6840), .S(n14856), .Z(
        P2_U3556) );
  MUX2_X1 U15431 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13412), .S(n14856), .Z(
        P2_U3555) );
  MUX2_X1 U15432 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13520), .S(n14856), .Z(
        P2_U3554) );
  MUX2_X1 U15433 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13406), .S(n14856), .Z(
        P2_U3553) );
  MUX2_X1 U15434 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13579), .S(n14856), .Z(
        P2_U3552) );
  MUX2_X1 U15435 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13401), .S(n14856), .Z(
        P2_U3551) );
  MUX2_X1 U15436 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13577), .S(n14856), .Z(
        P2_U3550) );
  MUX2_X1 U15437 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13396), .S(n14856), .Z(
        P2_U3549) );
  MUX2_X1 U15438 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13394), .S(n14856), .Z(
        P2_U3548) );
  MUX2_X1 U15439 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13391), .S(n14856), .Z(
        P2_U3547) );
  MUX2_X1 U15440 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13298), .S(n14856), .Z(
        P2_U3546) );
  MUX2_X1 U15441 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13299), .S(n14856), .Z(
        P2_U3545) );
  MUX2_X1 U15442 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13300), .S(n14856), .Z(
        P2_U3544) );
  MUX2_X1 U15443 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13301), .S(n14856), .Z(
        P2_U3543) );
  MUX2_X1 U15444 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13302), .S(P2_U3947), .Z(
        P2_U3542) );
  MUX2_X1 U15445 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13303), .S(P2_U3947), .Z(
        P2_U3541) );
  MUX2_X1 U15446 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13304), .S(P2_U3947), .Z(
        P2_U3540) );
  MUX2_X1 U15447 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13305), .S(P2_U3947), .Z(
        P2_U3539) );
  MUX2_X1 U15448 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13306), .S(P2_U3947), .Z(
        P2_U3538) );
  MUX2_X1 U15449 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13307), .S(P2_U3947), .Z(
        P2_U3537) );
  MUX2_X1 U15450 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13308), .S(n14856), .Z(
        P2_U3536) );
  MUX2_X1 U15451 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13309), .S(P2_U3947), .Z(
        P2_U3535) );
  MUX2_X1 U15452 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13310), .S(P2_U3947), .Z(
        P2_U3534) );
  MUX2_X1 U15453 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13311), .S(P2_U3947), .Z(
        P2_U3533) );
  MUX2_X1 U15454 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n9002), .S(n14856), .Z(
        P2_U3532) );
  MUX2_X1 U15455 ( .A(n10074), .B(P2_REG1_REG_2__SCAN_IN), .S(n13323), .Z(
        n13314) );
  NAND3_X1 U15456 ( .A1(n13314), .A2(n13313), .A3(n13312), .ZN(n13315) );
  NAND3_X1 U15457 ( .A1(n14943), .A2(n13316), .A3(n13315), .ZN(n13327) );
  AOI22_X1 U15458 ( .A1(n14935), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n13326) );
  OR3_X1 U15459 ( .A1(n13320), .A2(n13319), .A3(n13318), .ZN(n13321) );
  NAND3_X1 U15460 ( .A1(n14939), .A2(n13322), .A3(n13321), .ZN(n13325) );
  NAND2_X1 U15461 ( .A1(n14936), .A2(n13323), .ZN(n13324) );
  NAND4_X1 U15462 ( .A1(n13327), .A2(n13326), .A3(n13325), .A4(n13324), .ZN(
        P2_U3216) );
  INV_X1 U15463 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n14540) );
  OAI21_X1 U15464 ( .B1(n13368), .B2(n14540), .A(n13328), .ZN(n13329) );
  AOI21_X1 U15465 ( .B1(n13335), .B2(n14936), .A(n13329), .ZN(n13343) );
  OR3_X1 U15466 ( .A1(n13332), .A2(n13331), .A3(n13330), .ZN(n13333) );
  NAND3_X1 U15467 ( .A1(n13334), .A2(n14939), .A3(n13333), .ZN(n13342) );
  MUX2_X1 U15468 ( .A(n10087), .B(P2_REG1_REG_6__SCAN_IN), .S(n13335), .Z(
        n13336) );
  NAND3_X1 U15469 ( .A1(n13338), .A2(n13337), .A3(n13336), .ZN(n13339) );
  NAND3_X1 U15470 ( .A1(n14943), .A2(n13340), .A3(n13339), .ZN(n13341) );
  NAND3_X1 U15471 ( .A1(n13343), .A2(n13342), .A3(n13341), .ZN(P2_U3220) );
  OR3_X1 U15472 ( .A1(n13346), .A2(n13345), .A3(n13344), .ZN(n13347) );
  NAND3_X1 U15473 ( .A1(n13348), .A2(n14939), .A3(n13347), .ZN(n13360) );
  NOR2_X1 U15474 ( .A1(n14880), .A2(n13349), .ZN(n13350) );
  AOI211_X1 U15475 ( .C1(n14935), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n13351), .B(
        n13350), .ZN(n13359) );
  MUX2_X1 U15476 ( .A(n10093), .B(P2_REG1_REG_8__SCAN_IN), .S(n13352), .Z(
        n13353) );
  NAND3_X1 U15477 ( .A1(n13355), .A2(n13354), .A3(n13353), .ZN(n13356) );
  NAND3_X1 U15478 ( .A1(n14943), .A2(n13357), .A3(n13356), .ZN(n13358) );
  NAND3_X1 U15479 ( .A1(n13360), .A2(n13359), .A3(n13358), .ZN(P2_U3222) );
  INV_X1 U15480 ( .A(n13361), .ZN(n13366) );
  NOR3_X1 U15481 ( .A1(n13364), .A2(n13363), .A3(n13362), .ZN(n13365) );
  OAI21_X1 U15482 ( .B1(n13366), .B2(n13365), .A(n14939), .ZN(n13378) );
  INV_X1 U15483 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14759) );
  NAND2_X1 U15484 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n13367)
         );
  OAI21_X1 U15485 ( .B1(n13368), .B2(n14759), .A(n13367), .ZN(n13369) );
  AOI21_X1 U15486 ( .B1(n13370), .B2(n14936), .A(n13369), .ZN(n13377) );
  AOI21_X1 U15487 ( .B1(n13373), .B2(n13372), .A(n13371), .ZN(n13375) );
  OAI21_X1 U15488 ( .B1(n13375), .B2(n13374), .A(n14943), .ZN(n13376) );
  NAND3_X1 U15489 ( .A1(n13378), .A2(n13377), .A3(n13376), .ZN(P2_U3226) );
  OR2_X2 U15490 ( .A1(n13635), .A2(n13727), .ZN(n13633) );
  NOR2_X2 U15491 ( .A1(n13566), .A2(n13548), .ZN(n13547) );
  NAND2_X1 U15492 ( .A1(n13536), .A2(n13547), .ZN(n13532) );
  NAND2_X1 U15493 ( .A1(n13381), .A2(P2_B_REG_SCAN_IN), .ZN(n13382) );
  NAND2_X1 U15494 ( .A1(n15413), .A2(n13382), .ZN(n13442) );
  INV_X1 U15495 ( .A(n13442), .ZN(n13383) );
  NAND2_X1 U15496 ( .A1(n13384), .A2(n13383), .ZN(n13654) );
  NOR2_X1 U15497 ( .A1(n14964), .A2(n13654), .ZN(n13389) );
  NOR2_X1 U15498 ( .A1(n13750), .A2(n13640), .ZN(n13385) );
  AOI211_X1 U15499 ( .C1(n14964), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13389), 
        .B(n13385), .ZN(n13386) );
  OAI21_X1 U15500 ( .B1(n13651), .B2(n14958), .A(n13386), .ZN(P2_U3234) );
  OAI211_X1 U15501 ( .C1(n13445), .C2(n13754), .A(n11674), .B(n13387), .ZN(
        n13655) );
  NOR2_X1 U15502 ( .A1(n13754), .A2(n13640), .ZN(n13388) );
  AOI211_X1 U15503 ( .C1(n14964), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13389), 
        .B(n13388), .ZN(n13390) );
  OAI21_X1 U15504 ( .B1(n14958), .B2(n13655), .A(n13390), .ZN(P2_U3235) );
  NAND2_X1 U15505 ( .A1(n13419), .A2(n13391), .ZN(n13392) );
  NAND2_X1 U15506 ( .A1(n13393), .A2(n13392), .ZN(n13643) );
  NAND2_X1 U15507 ( .A1(n13727), .A2(n13394), .ZN(n13395) );
  INV_X1 U15508 ( .A(n13614), .ZN(n13610) );
  NAND2_X1 U15509 ( .A1(n13591), .A2(n13397), .ZN(n13399) );
  NAND2_X1 U15510 ( .A1(n13399), .A2(n13398), .ZN(n13587) );
  NAND2_X1 U15511 ( .A1(n13710), .A2(n13401), .ZN(n13400) );
  NAND2_X1 U15512 ( .A1(n13587), .A2(n13400), .ZN(n13403) );
  OR2_X1 U15513 ( .A1(n13710), .A2(n13401), .ZN(n13402) );
  NOR2_X1 U15514 ( .A1(n13568), .A2(n13579), .ZN(n13404) );
  NAND2_X1 U15515 ( .A1(n13568), .A2(n13579), .ZN(n13405) );
  AND2_X1 U15516 ( .A1(n13548), .A2(n13406), .ZN(n13407) );
  NAND2_X1 U15517 ( .A1(n13536), .A2(n13555), .ZN(n13408) );
  INV_X1 U15518 ( .A(n13516), .ZN(n13411) );
  NAND2_X1 U15519 ( .A1(n13688), .A2(n13412), .ZN(n13413) );
  NAND2_X1 U15520 ( .A1(n13519), .A2(n13413), .ZN(n13500) );
  NAND2_X1 U15521 ( .A1(n13512), .A2(n13485), .ZN(n13415) );
  INV_X1 U15522 ( .A(n13438), .ZN(n13436) );
  INV_X1 U15523 ( .A(n13495), .ZN(n13678) );
  INV_X1 U15524 ( .A(n13468), .ZN(n13478) );
  NAND2_X1 U15525 ( .A1(n13464), .A2(n6699), .ZN(n13463) );
  OR2_X1 U15526 ( .A1(n13419), .A2(n13418), .ZN(n13420) );
  NAND2_X1 U15527 ( .A1(n13727), .A2(n13423), .ZN(n13422) );
  OR2_X1 U15528 ( .A1(n13625), .A2(n13595), .ZN(n13424) );
  NAND2_X1 U15529 ( .A1(n13603), .A2(n13425), .ZN(n13427) );
  NOR2_X1 U15530 ( .A1(n13603), .A2(n13425), .ZN(n13426) );
  OR2_X1 U15531 ( .A1(n13710), .A2(n13597), .ZN(n13428) );
  NAND2_X1 U15532 ( .A1(n13710), .A2(n13597), .ZN(n13429) );
  AND2_X1 U15533 ( .A1(n13568), .A2(n13556), .ZN(n13430) );
  OR2_X1 U15534 ( .A1(n13548), .A2(n13563), .ZN(n13432) );
  OR2_X1 U15535 ( .A1(n13512), .A2(n6840), .ZN(n13435) );
  XNOR2_X1 U15536 ( .A(n13440), .B(n13439), .ZN(n13443) );
  OAI222_X1 U15537 ( .A1(n13594), .A2(n13444), .B1(n13443), .B2(n13562), .C1(
        n13442), .C2(n13441), .ZN(n13658) );
  NAND2_X1 U15538 ( .A1(n13658), .A2(n14952), .ZN(n13452) );
  AOI211_X1 U15539 ( .C1(n13659), .C2(n13458), .A(n11080), .B(n13445), .ZN(
        n13660) );
  NOR2_X1 U15540 ( .A1(n13446), .A2(n13640), .ZN(n13450) );
  OAI22_X1 U15541 ( .A1(n14952), .A2(n13448), .B1(n13447), .B2(n14950), .ZN(
        n13449) );
  AOI211_X1 U15542 ( .C1(n13660), .C2(n13649), .A(n13450), .B(n13449), .ZN(
        n13451) );
  OAI211_X1 U15543 ( .C1(n13662), .C2(n13646), .A(n13452), .B(n13451), .ZN(
        P2_U3236) );
  OAI211_X1 U15544 ( .C1(n13455), .C2(n13454), .A(n13453), .B(n13631), .ZN(
        n13457) );
  AND2_X1 U15545 ( .A1(n13457), .A2(n13456), .ZN(n13669) );
  AOI21_X1 U15546 ( .B1(n13474), .B2(n13668), .A(n11080), .ZN(n13459) );
  NOR2_X1 U15547 ( .A1(n14950), .A2(n13460), .ZN(n13461) );
  AOI21_X1 U15548 ( .B1(n14964), .B2(P2_REG2_REG_28__SCAN_IN), .A(n13461), 
        .ZN(n13462) );
  OAI21_X1 U15549 ( .B1(n7097), .B2(n13640), .A(n13462), .ZN(n13466) );
  NOR2_X1 U15550 ( .A1(n13666), .A2(n13646), .ZN(n13465) );
  AOI211_X1 U15551 ( .C1(n13667), .C2(n13649), .A(n13466), .B(n13465), .ZN(
        n13467) );
  OAI21_X1 U15552 ( .B1(n14964), .B2(n13669), .A(n13467), .ZN(P2_U3237) );
  XNOR2_X1 U15553 ( .A(n13469), .B(n13468), .ZN(n13471) );
  AOI21_X1 U15554 ( .B1(n13471), .B2(n13631), .A(n13470), .ZN(n13675) );
  OAI22_X1 U15555 ( .A1(n14952), .A2(n13473), .B1(n13472), .B2(n14950), .ZN(
        n13477) );
  AOI21_X1 U15556 ( .B1(n6505), .B2(n7100), .A(n11080), .ZN(n13475) );
  NAND2_X1 U15557 ( .A1(n13475), .A2(n13474), .ZN(n13672) );
  NOR2_X1 U15558 ( .A1(n13672), .A2(n14958), .ZN(n13476) );
  AOI211_X1 U15559 ( .C1(n14955), .C2(n7100), .A(n13477), .B(n13476), .ZN(
        n13481) );
  OR2_X1 U15560 ( .A1(n13479), .A2(n13478), .ZN(n13671) );
  NAND3_X1 U15561 ( .A1(n13671), .A2(n13670), .A3(n14960), .ZN(n13480) );
  OAI211_X1 U15562 ( .C1(n13675), .C2(n14964), .A(n13481), .B(n13480), .ZN(
        P2_U3238) );
  XNOR2_X1 U15563 ( .A(n13482), .B(n13489), .ZN(n13483) );
  NAND2_X1 U15564 ( .A1(n13483), .A2(n13631), .ZN(n13488) );
  OAI22_X1 U15565 ( .A1(n13485), .A2(n13594), .B1(n13484), .B2(n13596), .ZN(
        n13486) );
  INV_X1 U15566 ( .A(n13486), .ZN(n13487) );
  NAND2_X1 U15567 ( .A1(n13488), .A2(n13487), .ZN(n13680) );
  INV_X1 U15568 ( .A(n13680), .ZN(n13499) );
  INV_X1 U15569 ( .A(n13489), .ZN(n13490) );
  XNOR2_X1 U15570 ( .A(n6591), .B(n13490), .ZN(n13676) );
  AOI21_X1 U15571 ( .B1(n13508), .B2(n13495), .A(n11080), .ZN(n13491) );
  NAND2_X1 U15572 ( .A1(n13491), .A2(n6505), .ZN(n13677) );
  OAI22_X1 U15573 ( .A1(n14952), .A2(n13493), .B1(n13492), .B2(n14950), .ZN(
        n13494) );
  AOI21_X1 U15574 ( .B1(n13495), .B2(n14955), .A(n13494), .ZN(n13496) );
  OAI21_X1 U15575 ( .B1(n13677), .B2(n14958), .A(n13496), .ZN(n13497) );
  AOI21_X1 U15576 ( .B1(n13676), .B2(n14960), .A(n13497), .ZN(n13498) );
  OAI21_X1 U15577 ( .B1(n13499), .B2(n14964), .A(n13498), .ZN(P2_U3239) );
  XNOR2_X1 U15578 ( .A(n13500), .B(n7267), .ZN(n13686) );
  INV_X1 U15579 ( .A(n13501), .ZN(n13502) );
  AOI21_X1 U15580 ( .B1(n13503), .B2(n7267), .A(n13502), .ZN(n13505) );
  OAI21_X1 U15581 ( .B1(n13505), .B2(n13562), .A(n13504), .ZN(n13682) );
  NOR2_X1 U15582 ( .A1(n14950), .A2(n13506), .ZN(n13507) );
  OAI21_X1 U15583 ( .B1(n13682), .B2(n13507), .A(n14952), .ZN(n13515) );
  INV_X1 U15584 ( .A(n13524), .ZN(n13510) );
  INV_X1 U15585 ( .A(n13508), .ZN(n13509) );
  AOI211_X1 U15586 ( .C1(n13684), .C2(n13510), .A(n11080), .B(n13509), .ZN(
        n13683) );
  OAI22_X1 U15587 ( .A1(n13512), .A2(n13640), .B1(n14952), .B2(n13511), .ZN(
        n13513) );
  AOI21_X1 U15588 ( .B1(n13683), .B2(n13649), .A(n13513), .ZN(n13514) );
  OAI211_X1 U15589 ( .C1(n13686), .C2(n13646), .A(n13515), .B(n13514), .ZN(
        P2_U3240) );
  XNOR2_X1 U15590 ( .A(n13517), .B(n6590), .ZN(n13523) );
  NAND2_X1 U15591 ( .A1(n13517), .A2(n13516), .ZN(n13518) );
  NAND2_X1 U15592 ( .A1(n13519), .A2(n13518), .ZN(n13691) );
  AOI22_X1 U15593 ( .A1(n15413), .A2(n6840), .B1(n13520), .B2(n13576), .ZN(
        n13521) );
  OAI21_X1 U15594 ( .B1(n13691), .B2(n9920), .A(n13521), .ZN(n13522) );
  AOI21_X1 U15595 ( .B1(n13523), .B2(n13631), .A(n13522), .ZN(n13689) );
  AOI211_X1 U15596 ( .C1(n13688), .C2(n13532), .A(n11080), .B(n13524), .ZN(
        n13687) );
  AOI22_X1 U15597 ( .A1(n14964), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13525), 
        .B2(n13637), .ZN(n13526) );
  OAI21_X1 U15598 ( .B1(n13527), .B2(n13640), .A(n13526), .ZN(n13529) );
  NOR2_X1 U15599 ( .A1(n13691), .A2(n13609), .ZN(n13528) );
  AOI211_X1 U15600 ( .C1(n13687), .C2(n13649), .A(n13529), .B(n13528), .ZN(
        n13530) );
  OAI21_X1 U15601 ( .B1(n14964), .B2(n13689), .A(n13530), .ZN(P2_U3241) );
  XNOR2_X1 U15602 ( .A(n13538), .B(n13531), .ZN(n13698) );
  INV_X1 U15603 ( .A(n13547), .ZN(n13534) );
  INV_X1 U15604 ( .A(n13532), .ZN(n13533) );
  AOI211_X1 U15605 ( .C1(n13695), .C2(n13534), .A(n11080), .B(n13533), .ZN(
        n13693) );
  OAI22_X1 U15606 ( .A1(n13536), .A2(n13640), .B1(n14952), .B2(n13535), .ZN(
        n13537) );
  AOI21_X1 U15607 ( .B1(n13693), .B2(n13649), .A(n13537), .ZN(n13545) );
  XOR2_X1 U15608 ( .A(n13539), .B(n13538), .Z(n13540) );
  NAND2_X1 U15609 ( .A1(n13540), .A2(n13631), .ZN(n13696) );
  INV_X1 U15610 ( .A(n13694), .ZN(n13541) );
  OAI211_X1 U15611 ( .C1(n14950), .C2(n13542), .A(n13696), .B(n13541), .ZN(
        n13543) );
  NAND2_X1 U15612 ( .A1(n13543), .A2(n14952), .ZN(n13544) );
  OAI211_X1 U15613 ( .C1(n13698), .C2(n13646), .A(n13545), .B(n13544), .ZN(
        P2_U3242) );
  XNOR2_X1 U15614 ( .A(n7165), .B(n13546), .ZN(n13701) );
  INV_X1 U15615 ( .A(n13701), .ZN(n13559) );
  AOI211_X1 U15616 ( .C1(n13548), .C2(n13566), .A(n11080), .B(n13547), .ZN(
        n13700) );
  INV_X1 U15617 ( .A(n13548), .ZN(n13765) );
  NOR2_X1 U15618 ( .A1(n13765), .A2(n13640), .ZN(n13552) );
  OAI22_X1 U15619 ( .A1(n14952), .A2(n13550), .B1(n13549), .B2(n14950), .ZN(
        n13551) );
  AOI211_X1 U15620 ( .C1(n13700), .C2(n13649), .A(n13552), .B(n13551), .ZN(
        n13558) );
  XNOR2_X1 U15621 ( .A(n13553), .B(n7165), .ZN(n13554) );
  OAI222_X1 U15622 ( .A1(n13594), .A2(n13556), .B1(n13596), .B2(n13555), .C1(
        n13554), .C2(n13562), .ZN(n13699) );
  NAND2_X1 U15623 ( .A1(n13699), .A2(n14952), .ZN(n13557) );
  OAI211_X1 U15624 ( .C1(n13559), .C2(n13646), .A(n13558), .B(n13557), .ZN(
        P2_U3243) );
  XOR2_X1 U15625 ( .A(n13560), .B(n13564), .Z(n13561) );
  OAI222_X1 U15626 ( .A1(n13594), .A2(n13597), .B1(n13596), .B2(n13563), .C1(
        n13562), .C2(n13561), .ZN(n13704) );
  INV_X1 U15627 ( .A(n13704), .ZN(n13574) );
  XOR2_X1 U15628 ( .A(n13565), .B(n13564), .Z(n13706) );
  INV_X1 U15629 ( .A(n13566), .ZN(n13567) );
  AOI211_X1 U15630 ( .C1(n13568), .C2(n13581), .A(n11080), .B(n13567), .ZN(
        n13705) );
  NAND2_X1 U15631 ( .A1(n13705), .A2(n13649), .ZN(n13571) );
  AOI22_X1 U15632 ( .A1(n13569), .A2(n13637), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n14964), .ZN(n13570) );
  OAI211_X1 U15633 ( .C1(n7107), .C2(n13640), .A(n13571), .B(n13570), .ZN(
        n13572) );
  AOI21_X1 U15634 ( .B1(n14960), .B2(n13706), .A(n13572), .ZN(n13573) );
  OAI21_X1 U15635 ( .B1(n14964), .B2(n13574), .A(n13573), .ZN(P2_U3244) );
  XNOR2_X1 U15636 ( .A(n13575), .B(n13586), .ZN(n13580) );
  AOI222_X1 U15637 ( .A1(n13631), .A2(n13580), .B1(n13579), .B2(n15413), .C1(
        n13577), .C2(n13576), .ZN(n13711) );
  AOI211_X1 U15638 ( .C1(n13710), .C2(n13601), .A(n11080), .B(n7108), .ZN(
        n13709) );
  INV_X1 U15639 ( .A(n13710), .ZN(n13585) );
  INV_X1 U15640 ( .A(n13582), .ZN(n13583) );
  AOI22_X1 U15641 ( .A1(n13583), .A2(n13637), .B1(P2_REG2_REG_20__SCAN_IN), 
        .B2(n14964), .ZN(n13584) );
  OAI21_X1 U15642 ( .B1(n13585), .B2(n13640), .A(n13584), .ZN(n13589) );
  XNOR2_X1 U15643 ( .A(n13587), .B(n13586), .ZN(n13713) );
  NOR2_X1 U15644 ( .A1(n13713), .A2(n13646), .ZN(n13588) );
  AOI211_X1 U15645 ( .C1(n13709), .C2(n13649), .A(n13589), .B(n13588), .ZN(
        n13590) );
  OAI21_X1 U15646 ( .B1(n14964), .B2(n13711), .A(n13590), .ZN(P2_U3245) );
  XNOR2_X1 U15647 ( .A(n13591), .B(n13592), .ZN(n13714) );
  XOR2_X1 U15648 ( .A(n13593), .B(n13592), .Z(n13599) );
  OAI22_X1 U15649 ( .A1(n13597), .A2(n13596), .B1(n13595), .B2(n13594), .ZN(
        n13598) );
  AOI21_X1 U15650 ( .B1(n13599), .B2(n13631), .A(n13598), .ZN(n13600) );
  OAI21_X1 U15651 ( .B1(n9920), .B2(n13714), .A(n13600), .ZN(n13715) );
  NAND2_X1 U15652 ( .A1(n13715), .A2(n14952), .ZN(n13608) );
  INV_X1 U15653 ( .A(n13601), .ZN(n13602) );
  AOI211_X1 U15654 ( .C1(n13603), .C2(n13621), .A(n11080), .B(n13602), .ZN(
        n13716) );
  AOI22_X1 U15655 ( .A1(n14964), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13604), 
        .B2(n13637), .ZN(n13605) );
  OAI21_X1 U15656 ( .B1(n7109), .B2(n13640), .A(n13605), .ZN(n13606) );
  AOI21_X1 U15657 ( .B1(n13716), .B2(n13649), .A(n13606), .ZN(n13607) );
  OAI211_X1 U15658 ( .C1(n13714), .C2(n13609), .A(n13608), .B(n13607), .ZN(
        P2_U3246) );
  NAND2_X1 U15659 ( .A1(n13611), .A2(n13610), .ZN(n13612) );
  NAND2_X1 U15660 ( .A1(n13613), .A2(n13612), .ZN(n13720) );
  INV_X1 U15661 ( .A(n13720), .ZN(n13628) );
  XNOR2_X1 U15662 ( .A(n13615), .B(n13614), .ZN(n13616) );
  NAND2_X1 U15663 ( .A1(n13616), .A2(n13631), .ZN(n13618) );
  NAND2_X1 U15664 ( .A1(n13618), .A2(n13617), .ZN(n13724) );
  NAND2_X1 U15665 ( .A1(n13724), .A2(n14952), .ZN(n13627) );
  OAI22_X1 U15666 ( .A1(n14952), .A2(n13620), .B1(n13619), .B2(n14950), .ZN(
        n13624) );
  AOI21_X1 U15667 ( .B1(n13625), .B2(n13633), .A(n11080), .ZN(n13622) );
  NAND2_X1 U15668 ( .A1(n13622), .A2(n13621), .ZN(n13721) );
  NOR2_X1 U15669 ( .A1(n13721), .A2(n14958), .ZN(n13623) );
  AOI211_X1 U15670 ( .C1(n14955), .C2(n13625), .A(n13624), .B(n13623), .ZN(
        n13626) );
  OAI211_X1 U15671 ( .C1(n13646), .C2(n13628), .A(n13627), .B(n13626), .ZN(
        P2_U3247) );
  XNOR2_X1 U15672 ( .A(n13629), .B(n13642), .ZN(n13632) );
  AOI21_X1 U15673 ( .B1(n13632), .B2(n13631), .A(n13630), .ZN(n13729) );
  INV_X1 U15674 ( .A(n13633), .ZN(n13634) );
  AOI211_X1 U15675 ( .C1(n13727), .C2(n13635), .A(n11080), .B(n13634), .ZN(
        n13726) );
  INV_X1 U15676 ( .A(n13636), .ZN(n13638) );
  AOI22_X1 U15677 ( .A1(n14964), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13638), 
        .B2(n13637), .ZN(n13639) );
  OAI21_X1 U15678 ( .B1(n13641), .B2(n13640), .A(n13639), .ZN(n13648) );
  OR2_X1 U15679 ( .A1(n13643), .A2(n13642), .ZN(n13644) );
  NAND2_X1 U15680 ( .A1(n13645), .A2(n13644), .ZN(n13730) );
  NOR2_X1 U15681 ( .A1(n13730), .A2(n13646), .ZN(n13647) );
  AOI211_X1 U15682 ( .C1(n13726), .C2(n13649), .A(n13648), .B(n13647), .ZN(
        n13650) );
  OAI21_X1 U15683 ( .B1(n14964), .B2(n13729), .A(n13650), .ZN(P2_U3248) );
  AND2_X1 U15684 ( .A1(n13651), .A2(n13654), .ZN(n13748) );
  MUX2_X1 U15685 ( .A(n13748), .B(n13652), .S(n15025), .Z(n13653) );
  OAI21_X1 U15686 ( .B1(n13750), .B2(n13736), .A(n13653), .ZN(P2_U3530) );
  NAND2_X1 U15687 ( .A1(n13655), .A2(n13654), .ZN(n13751) );
  MUX2_X1 U15688 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13751), .S(n15027), .Z(
        n13656) );
  INV_X1 U15689 ( .A(n13656), .ZN(n13657) );
  OAI21_X1 U15690 ( .B1(n13754), .B2(n13736), .A(n13657), .ZN(P2_U3529) );
  INV_X1 U15691 ( .A(n13663), .ZN(n13664) );
  NAND2_X1 U15692 ( .A1(n13665), .A2(n13664), .ZN(n13755) );
  MUX2_X1 U15693 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13755), .S(n15027), .Z(
        P2_U3528) );
  MUX2_X1 U15694 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13756), .S(n15027), .Z(
        P2_U3527) );
  NAND2_X1 U15695 ( .A1(n7100), .A2(n14990), .ZN(n13674) );
  NAND3_X1 U15696 ( .A1(n13671), .A2(n13670), .A3(n15009), .ZN(n13673) );
  NAND4_X1 U15697 ( .A1(n13675), .A2(n13674), .A3(n13673), .A4(n13672), .ZN(
        n13757) );
  MUX2_X1 U15698 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13757), .S(n15027), .Z(
        P2_U3526) );
  AND2_X1 U15699 ( .A1(n13676), .A2(n15009), .ZN(n13681) );
  OAI21_X1 U15700 ( .B1(n13678), .B2(n15012), .A(n13677), .ZN(n13679) );
  MUX2_X1 U15701 ( .A(n13758), .B(P2_REG1_REG_26__SCAN_IN), .S(n15025), .Z(
        P2_U3525) );
  AOI211_X1 U15702 ( .C1(n14990), .C2(n13684), .A(n13683), .B(n13682), .ZN(
        n13685) );
  OAI21_X1 U15703 ( .B1(n14994), .B2(n13686), .A(n13685), .ZN(n13759) );
  MUX2_X1 U15704 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13759), .S(n15027), .Z(
        P2_U3524) );
  AOI21_X1 U15705 ( .B1(n14990), .B2(n13688), .A(n13687), .ZN(n13690) );
  OAI211_X1 U15706 ( .C1(n13692), .C2(n13691), .A(n13690), .B(n13689), .ZN(
        n13760) );
  MUX2_X1 U15707 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13760), .S(n15027), .Z(
        P2_U3523) );
  AOI211_X1 U15708 ( .C1(n14990), .C2(n13695), .A(n13694), .B(n13693), .ZN(
        n13697) );
  OAI211_X1 U15709 ( .C1(n14994), .C2(n13698), .A(n13697), .B(n13696), .ZN(
        n13761) );
  MUX2_X1 U15710 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13761), .S(n15027), .Z(
        P2_U3522) );
  AOI211_X1 U15711 ( .C1(n15009), .C2(n13701), .A(n13700), .B(n13699), .ZN(
        n13762) );
  MUX2_X1 U15712 ( .A(n13702), .B(n13762), .S(n15027), .Z(n13703) );
  OAI21_X1 U15713 ( .B1(n13765), .B2(n13736), .A(n13703), .ZN(P2_U3521) );
  AOI211_X1 U15714 ( .C1(n13706), .C2(n15009), .A(n13705), .B(n13704), .ZN(
        n13766) );
  MUX2_X1 U15715 ( .A(n13707), .B(n13766), .S(n15027), .Z(n13708) );
  OAI21_X1 U15716 ( .B1(n7107), .B2(n13736), .A(n13708), .ZN(P2_U3520) );
  AOI21_X1 U15717 ( .B1(n14990), .B2(n13710), .A(n13709), .ZN(n13712) );
  OAI211_X1 U15718 ( .C1(n14994), .C2(n13713), .A(n13712), .B(n13711), .ZN(
        n13769) );
  MUX2_X1 U15719 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13769), .S(n15027), .Z(
        P2_U3519) );
  INV_X1 U15720 ( .A(n13714), .ZN(n13717) );
  AOI211_X1 U15721 ( .C1(n13717), .C2(n15000), .A(n13716), .B(n13715), .ZN(
        n13770) );
  MUX2_X1 U15722 ( .A(n13718), .B(n13770), .S(n15027), .Z(n13719) );
  OAI21_X1 U15723 ( .B1(n7109), .B2(n13736), .A(n13719), .ZN(P2_U3518) );
  NAND2_X1 U15724 ( .A1(n13720), .A2(n15009), .ZN(n13722) );
  OAI211_X1 U15725 ( .C1(n13723), .C2(n15012), .A(n13722), .B(n13721), .ZN(
        n13725) );
  MUX2_X1 U15726 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13773), .S(n15027), .Z(
        P2_U3517) );
  AOI21_X1 U15727 ( .B1(n14990), .B2(n13727), .A(n13726), .ZN(n13728) );
  OAI211_X1 U15728 ( .C1(n14994), .C2(n13730), .A(n13729), .B(n13728), .ZN(
        n13774) );
  MUX2_X1 U15729 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13774), .S(n15027), .Z(
        P2_U3516) );
  AOI211_X1 U15730 ( .C1(n13733), .C2(n15009), .A(n13732), .B(n13731), .ZN(
        n13775) );
  MUX2_X1 U15731 ( .A(n13734), .B(n13775), .S(n15027), .Z(n13735) );
  OAI21_X1 U15732 ( .B1(n13779), .B2(n13736), .A(n13735), .ZN(P2_U3515) );
  OAI211_X1 U15733 ( .C1(n14994), .C2(n13739), .A(n13738), .B(n13737), .ZN(
        n13780) );
  MUX2_X1 U15734 ( .A(n13780), .B(P2_REG1_REG_15__SCAN_IN), .S(n15025), .Z(
        n13740) );
  AOI21_X1 U15735 ( .B1(n13745), .B2(n13782), .A(n13740), .ZN(n13741) );
  INV_X1 U15736 ( .A(n13741), .ZN(P2_U3514) );
  MUX2_X1 U15737 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13742), .S(n15027), .Z(
        n13743) );
  AOI21_X1 U15738 ( .B1(n13745), .B2(n13744), .A(n13743), .ZN(n13746) );
  INV_X1 U15739 ( .A(n13746), .ZN(P2_U3513) );
  INV_X1 U15740 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13747) );
  MUX2_X1 U15741 ( .A(n13748), .B(n13747), .S(n15017), .Z(n13749) );
  OAI21_X1 U15742 ( .B1(n13750), .B2(n13778), .A(n13749), .ZN(P2_U3498) );
  MUX2_X1 U15743 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13751), .S(n15018), .Z(
        n13752) );
  INV_X1 U15744 ( .A(n13752), .ZN(n13753) );
  OAI21_X1 U15745 ( .B1(n13754), .B2(n13778), .A(n13753), .ZN(P2_U3497) );
  MUX2_X1 U15746 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13755), .S(n15018), .Z(
        P2_U3496) );
  MUX2_X1 U15747 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13757), .S(n15018), .Z(
        P2_U3494) );
  MUX2_X1 U15748 ( .A(n13758), .B(P2_REG0_REG_26__SCAN_IN), .S(n15017), .Z(
        P2_U3493) );
  MUX2_X1 U15749 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13759), .S(n15018), .Z(
        P2_U3492) );
  MUX2_X1 U15750 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13760), .S(n15018), .Z(
        P2_U3491) );
  MUX2_X1 U15751 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13761), .S(n15018), .Z(
        P2_U3490) );
  INV_X1 U15752 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n13763) );
  MUX2_X1 U15753 ( .A(n13763), .B(n13762), .S(n15018), .Z(n13764) );
  OAI21_X1 U15754 ( .B1(n13765), .B2(n13778), .A(n13764), .ZN(P2_U3489) );
  INV_X1 U15755 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13767) );
  MUX2_X1 U15756 ( .A(n13767), .B(n13766), .S(n15018), .Z(n13768) );
  OAI21_X1 U15757 ( .B1(n7107), .B2(n13778), .A(n13768), .ZN(P2_U3488) );
  MUX2_X1 U15758 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13769), .S(n15018), .Z(
        P2_U3487) );
  INV_X1 U15759 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n13771) );
  MUX2_X1 U15760 ( .A(n13771), .B(n13770), .S(n15018), .Z(n13772) );
  OAI21_X1 U15761 ( .B1(n7109), .B2(n13778), .A(n13772), .ZN(P2_U3486) );
  MUX2_X1 U15762 ( .A(n13773), .B(P2_REG0_REG_18__SCAN_IN), .S(n15017), .Z(
        P2_U3484) );
  MUX2_X1 U15763 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13774), .S(n15018), .Z(
        P2_U3481) );
  INV_X1 U15764 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n13776) );
  MUX2_X1 U15765 ( .A(n13776), .B(n13775), .S(n15018), .Z(n13777) );
  OAI21_X1 U15766 ( .B1(n13779), .B2(n13778), .A(n13777), .ZN(P2_U3478) );
  MUX2_X1 U15767 ( .A(n13780), .B(P2_REG0_REG_15__SCAN_IN), .S(n15017), .Z(
        n13781) );
  AOI21_X1 U15768 ( .B1(n13783), .B2(n13782), .A(n13781), .ZN(n13784) );
  INV_X1 U15769 ( .A(n13784), .ZN(P2_U3475) );
  INV_X1 U15770 ( .A(n13785), .ZN(n14452) );
  NOR4_X1 U15771 ( .A1(n13787), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13786), .A4(
        P2_U3088), .ZN(n13788) );
  AOI21_X1 U15772 ( .B1(n13792), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13788), 
        .ZN(n13789) );
  OAI21_X1 U15773 ( .B1(n14452), .B2(n13794), .A(n13789), .ZN(P2_U3296) );
  INV_X1 U15774 ( .A(n13790), .ZN(n14457) );
  AOI21_X1 U15775 ( .B1(n13792), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13791), 
        .ZN(n13793) );
  OAI21_X1 U15776 ( .B1(n14457), .B2(n13794), .A(n13793), .ZN(P2_U3299) );
  INV_X1 U15777 ( .A(n13795), .ZN(n14460) );
  OAI222_X1 U15778 ( .A1(n13807), .A2(n13797), .B1(n13805), .B2(n14460), .C1(
        n13796), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U15779 ( .A(n13798), .ZN(n14463) );
  OAI222_X1 U15780 ( .A1(n13800), .A2(P2_U3088), .B1(n13805), .B2(n14463), 
        .C1(n13799), .C2(n13807), .ZN(P2_U3301) );
  INV_X1 U15781 ( .A(n13801), .ZN(n14467) );
  OAI222_X1 U15782 ( .A1(n13807), .A2(n13803), .B1(n13805), .B2(n14467), .C1(
        n13802), .C2(P2_U3088), .ZN(P2_U3302) );
  OAI222_X1 U15783 ( .A1(n13807), .A2(n13806), .B1(n13805), .B2(n14471), .C1(
        n13804), .C2(P2_U3088), .ZN(P2_U3303) );
  INV_X1 U15784 ( .A(n13808), .ZN(n13809) );
  MUX2_X1 U15785 ( .A(n13809), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI22_X1 U15786 ( .A1(n14118), .A2(n13938), .B1(n13948), .B2(n10801), .ZN(
        n13932) );
  NAND2_X1 U15787 ( .A1(n14337), .A2(n13902), .ZN(n13811) );
  NAND2_X1 U15788 ( .A1(n14024), .A2(n11103), .ZN(n13810) );
  NAND2_X1 U15789 ( .A1(n13811), .A2(n13810), .ZN(n13813) );
  INV_X2 U15790 ( .A(n13812), .ZN(n13940) );
  XNOR2_X1 U15791 ( .A(n13813), .B(n13940), .ZN(n13931) );
  XOR2_X1 U15792 ( .A(n13932), .B(n13931), .Z(n13935) );
  NAND2_X1 U15793 ( .A1(n13820), .A2(n13902), .ZN(n13818) );
  NAND2_X1 U15794 ( .A1(n14621), .A2(n11103), .ZN(n13817) );
  NAND2_X1 U15795 ( .A1(n13818), .A2(n13817), .ZN(n13819) );
  XNOR2_X1 U15796 ( .A(n13819), .B(n13940), .ZN(n13823) );
  AOI22_X1 U15797 ( .A1(n13820), .A2(n11103), .B1(n13906), .B2(n14621), .ZN(
        n13821) );
  XNOR2_X1 U15798 ( .A(n13823), .B(n13821), .ZN(n14701) );
  INV_X1 U15799 ( .A(n13821), .ZN(n13822) );
  OR2_X1 U15800 ( .A1(n13823), .A2(n13822), .ZN(n13824) );
  NAND2_X1 U15801 ( .A1(n14699), .A2(n13824), .ZN(n13829) );
  NAND2_X1 U15802 ( .A1(n13828), .A2(n13902), .ZN(n13826) );
  NAND2_X1 U15803 ( .A1(n14702), .A2(n11103), .ZN(n13825) );
  NAND2_X1 U15804 ( .A1(n13826), .A2(n13825), .ZN(n13827) );
  XNOR2_X1 U15805 ( .A(n13827), .B(n13940), .ZN(n13830) );
  XNOR2_X1 U15806 ( .A(n13829), .B(n13830), .ZN(n14014) );
  OAI22_X1 U15807 ( .A1(n14447), .A2(n13938), .B1(n14713), .B2(n10801), .ZN(
        n14013) );
  INV_X1 U15808 ( .A(n13829), .ZN(n13831) );
  NAND2_X1 U15809 ( .A1(n14721), .A2(n13902), .ZN(n13833) );
  NAND2_X1 U15810 ( .A1(n14028), .A2(n11103), .ZN(n13832) );
  NAND2_X1 U15811 ( .A1(n13833), .A2(n13832), .ZN(n13834) );
  XNOR2_X1 U15812 ( .A(n13834), .B(n13940), .ZN(n13841) );
  AND2_X1 U15813 ( .A1(n14028), .A2(n13906), .ZN(n13835) );
  AOI21_X1 U15814 ( .B1(n14721), .B2(n11103), .A(n13835), .ZN(n13839) );
  XNOR2_X1 U15815 ( .A(n13841), .B(n13839), .ZN(n14715) );
  INV_X1 U15816 ( .A(n13839), .ZN(n13840) );
  NAND2_X1 U15817 ( .A1(n14735), .A2(n13902), .ZN(n13844) );
  NAND2_X1 U15818 ( .A1(n14296), .A2(n11103), .ZN(n13843) );
  NAND2_X1 U15819 ( .A1(n13844), .A2(n13843), .ZN(n13845) );
  XNOR2_X1 U15820 ( .A(n13845), .B(n13940), .ZN(n13848) );
  AOI22_X1 U15821 ( .A1(n14735), .A2(n11103), .B1(n13906), .B2(n14296), .ZN(
        n13846) );
  XNOR2_X1 U15822 ( .A(n13848), .B(n13846), .ZN(n14729) );
  INV_X1 U15823 ( .A(n13846), .ZN(n13847) );
  OR2_X1 U15824 ( .A1(n13848), .A2(n13847), .ZN(n13849) );
  NAND2_X1 U15825 ( .A1(n14385), .A2(n13902), .ZN(n13851) );
  NAND2_X1 U15826 ( .A1(n14027), .A2(n11103), .ZN(n13850) );
  NAND2_X1 U15827 ( .A1(n13851), .A2(n13850), .ZN(n13852) );
  XNOR2_X1 U15828 ( .A(n13852), .B(n13940), .ZN(n13855) );
  AOI22_X1 U15829 ( .A1(n14385), .A2(n11103), .B1(n13906), .B2(n14027), .ZN(
        n13853) );
  XNOR2_X1 U15830 ( .A(n13855), .B(n13853), .ZN(n13997) );
  INV_X1 U15831 ( .A(n13853), .ZN(n13854) );
  NOR2_X1 U15832 ( .A1(n13855), .A2(n13854), .ZN(n13856) );
  NAND2_X1 U15833 ( .A1(n14237), .A2(n13902), .ZN(n13858) );
  NAND2_X1 U15834 ( .A1(n14259), .A2(n11103), .ZN(n13857) );
  NAND2_X1 U15835 ( .A1(n13858), .A2(n13857), .ZN(n13859) );
  XNOR2_X1 U15836 ( .A(n13859), .B(n13940), .ZN(n13863) );
  AND2_X1 U15837 ( .A1(n14259), .A2(n13906), .ZN(n13860) );
  AOI21_X1 U15838 ( .B1(n14237), .B2(n11103), .A(n13860), .ZN(n13861) );
  XNOR2_X1 U15839 ( .A(n13863), .B(n13861), .ZN(n13925) );
  INV_X1 U15840 ( .A(n13861), .ZN(n13862) );
  NAND2_X1 U15841 ( .A1(n13863), .A2(n13862), .ZN(n13864) );
  NAND2_X1 U15842 ( .A1(n13924), .A2(n13864), .ZN(n13980) );
  OAI22_X1 U15843 ( .A1(n14437), .A2(n13938), .B1(n13956), .B2(n10801), .ZN(
        n13866) );
  OAI22_X1 U15844 ( .A1(n14437), .A2(n13936), .B1(n13956), .B2(n13938), .ZN(
        n13865) );
  XNOR2_X1 U15845 ( .A(n13865), .B(n13940), .ZN(n13867) );
  XOR2_X1 U15846 ( .A(n13866), .B(n13867), .Z(n13979) );
  NAND2_X1 U15847 ( .A1(n13867), .A2(n13866), .ZN(n13868) );
  AOI22_X1 U15848 ( .A1(n14431), .A2(n13902), .B1(n11103), .B2(n14197), .ZN(
        n13869) );
  XNOR2_X1 U15849 ( .A(n13869), .B(n13940), .ZN(n13871) );
  AOI22_X1 U15850 ( .A1(n14431), .A2(n11103), .B1(n13906), .B2(n14197), .ZN(
        n13870) );
  XNOR2_X1 U15851 ( .A(n13871), .B(n13870), .ZN(n13955) );
  NAND2_X1 U15852 ( .A1(n13871), .A2(n13870), .ZN(n13872) );
  NAND2_X1 U15853 ( .A1(n13952), .A2(n13872), .ZN(n13988) );
  OAI22_X1 U15854 ( .A1(n14361), .A2(n13936), .B1(n13919), .B2(n13938), .ZN(
        n13873) );
  XNOR2_X1 U15855 ( .A(n13873), .B(n13940), .ZN(n13875) );
  AND2_X1 U15856 ( .A1(n14025), .A2(n13906), .ZN(n13874) );
  AOI21_X1 U15857 ( .B1(n14193), .B2(n11103), .A(n13874), .ZN(n13876) );
  XNOR2_X1 U15858 ( .A(n13875), .B(n13876), .ZN(n13989) );
  NAND2_X1 U15859 ( .A1(n13988), .A2(n13989), .ZN(n13987) );
  INV_X1 U15860 ( .A(n13875), .ZN(n13877) );
  NAND2_X1 U15861 ( .A1(n13877), .A2(n13876), .ZN(n13878) );
  NAND2_X1 U15862 ( .A1(n13987), .A2(n13878), .ZN(n13917) );
  NAND2_X1 U15863 ( .A1(n14356), .A2(n13902), .ZN(n13880) );
  NAND2_X1 U15864 ( .A1(n14196), .A2(n11103), .ZN(n13879) );
  NAND2_X1 U15865 ( .A1(n13880), .A2(n13879), .ZN(n13881) );
  XNOR2_X1 U15866 ( .A(n13881), .B(n13940), .ZN(n13882) );
  AOI22_X1 U15867 ( .A1(n14356), .A2(n11103), .B1(n13906), .B2(n14196), .ZN(
        n13883) );
  XNOR2_X1 U15868 ( .A(n13882), .B(n13883), .ZN(n13916) );
  NAND2_X1 U15869 ( .A1(n13917), .A2(n13916), .ZN(n13886) );
  INV_X1 U15870 ( .A(n13882), .ZN(n13884) );
  NAND2_X1 U15871 ( .A1(n13884), .A2(n13883), .ZN(n13885) );
  NAND2_X1 U15872 ( .A1(n14351), .A2(n13902), .ZN(n13888) );
  NAND2_X1 U15873 ( .A1(n14142), .A2(n11103), .ZN(n13887) );
  NAND2_X1 U15874 ( .A1(n13888), .A2(n13887), .ZN(n13889) );
  XNOR2_X1 U15875 ( .A(n13889), .B(n13940), .ZN(n13892) );
  AOI22_X1 U15876 ( .A1(n14351), .A2(n11103), .B1(n13906), .B2(n14142), .ZN(
        n13890) );
  XNOR2_X1 U15877 ( .A(n13892), .B(n13890), .ZN(n13972) );
  INV_X1 U15878 ( .A(n13890), .ZN(n13891) );
  NAND2_X1 U15879 ( .A1(n14346), .A2(n13902), .ZN(n13895) );
  NAND2_X1 U15880 ( .A1(n14159), .A2(n11103), .ZN(n13894) );
  NAND2_X1 U15881 ( .A1(n13895), .A2(n13894), .ZN(n13896) );
  XNOR2_X1 U15882 ( .A(n13896), .B(n13940), .ZN(n13897) );
  AOI22_X1 U15883 ( .A1(n14346), .A2(n11103), .B1(n13906), .B2(n14159), .ZN(
        n13898) );
  XNOR2_X1 U15884 ( .A(n13897), .B(n13898), .ZN(n13964) );
  INV_X1 U15885 ( .A(n13897), .ZN(n13899) );
  NAND2_X1 U15886 ( .A1(n13899), .A2(n13898), .ZN(n13900) );
  NAND2_X1 U15887 ( .A1(n14130), .A2(n13902), .ZN(n13904) );
  NAND2_X1 U15888 ( .A1(n14143), .A2(n11103), .ZN(n13903) );
  NAND2_X1 U15889 ( .A1(n13904), .A2(n13903), .ZN(n13905) );
  XNOR2_X1 U15890 ( .A(n13905), .B(n13940), .ZN(n13907) );
  AOI22_X1 U15891 ( .A1(n14130), .A2(n11103), .B1(n13906), .B2(n14143), .ZN(
        n13908) );
  XNOR2_X1 U15892 ( .A(n13907), .B(n13908), .ZN(n14006) );
  INV_X1 U15893 ( .A(n13907), .ZN(n13909) );
  NAND2_X1 U15894 ( .A1(n13909), .A2(n13908), .ZN(n13910) );
  AOI22_X1 U15895 ( .A1(n14703), .A2(n14107), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13912) );
  NAND2_X1 U15896 ( .A1(n14018), .A2(n14116), .ZN(n13911) );
  OAI211_X1 U15897 ( .C1(n13967), .C2(n14725), .A(n13912), .B(n13911), .ZN(
        n13913) );
  AOI21_X1 U15898 ( .B1(n14337), .B2(n15197), .A(n13913), .ZN(n13914) );
  OAI21_X1 U15899 ( .B1(n13915), .B2(n14731), .A(n13914), .ZN(P1_U3214) );
  XOR2_X1 U15900 ( .A(n13917), .B(n13916), .Z(n13923) );
  OAI22_X1 U15901 ( .A1(n13919), .A2(n14273), .B1(n13918), .B2(n14274), .ZN(
        n14177) );
  AOI22_X1 U15902 ( .A1(n15200), .A2(n14177), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13920) );
  OAI21_X1 U15903 ( .B1(n14179), .B2(n15204), .A(n13920), .ZN(n13921) );
  AOI21_X1 U15904 ( .B1(n14356), .B2(n15197), .A(n13921), .ZN(n13922) );
  OAI21_X1 U15905 ( .B1(n13923), .B2(n14731), .A(n13922), .ZN(P1_U3216) );
  OAI211_X1 U15906 ( .C1(n13926), .C2(n13925), .A(n13924), .B(n15206), .ZN(
        n13930) );
  AOI22_X1 U15907 ( .A1(n14026), .A2(n14620), .B1(n14619), .B2(n14027), .ZN(
        n14245) );
  OAI21_X1 U15908 ( .B1(n14245), .B2(n14015), .A(n13927), .ZN(n13928) );
  AOI21_X1 U15909 ( .B1(n14249), .B2(n14018), .A(n13928), .ZN(n13929) );
  OAI211_X1 U15910 ( .C1(n7003), .C2(n14707), .A(n13930), .B(n13929), .ZN(
        P1_U3219) );
  INV_X1 U15911 ( .A(n13931), .ZN(n13934) );
  INV_X1 U15912 ( .A(n13932), .ZN(n13933) );
  OAI22_X1 U15913 ( .A1(n13939), .A2(n13936), .B1(n13937), .B2(n13938), .ZN(
        n13943) );
  OAI22_X1 U15914 ( .A1(n13939), .A2(n13938), .B1(n13937), .B2(n10801), .ZN(
        n13941) );
  XNOR2_X1 U15915 ( .A(n13941), .B(n13940), .ZN(n13942) );
  XOR2_X1 U15916 ( .A(n13943), .B(n13942), .Z(n13944) );
  AOI22_X1 U15917 ( .A1(n14703), .A2(n14023), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13947) );
  NAND2_X1 U15918 ( .A1(n14018), .A2(n13945), .ZN(n13946) );
  OAI211_X1 U15919 ( .C1(n13948), .C2(n14725), .A(n13947), .B(n13946), .ZN(
        n13949) );
  AOI21_X1 U15920 ( .B1(n14330), .B2(n15197), .A(n13949), .ZN(n13950) );
  OAI21_X1 U15921 ( .B1(n13951), .B2(n14731), .A(n13950), .ZN(P1_U3220) );
  INV_X1 U15922 ( .A(n13952), .ZN(n13953) );
  AOI21_X1 U15923 ( .B1(n13955), .B2(n13954), .A(n13953), .ZN(n13962) );
  OR2_X1 U15924 ( .A1(n13956), .A2(n14273), .ZN(n13958) );
  NAND2_X1 U15925 ( .A1(n14025), .A2(n14620), .ZN(n13957) );
  NAND2_X1 U15926 ( .A1(n13958), .A2(n13957), .ZN(n14209) );
  AOI22_X1 U15927 ( .A1(n14209), .A2(n15200), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13959) );
  OAI21_X1 U15928 ( .B1(n14215), .B2(n15204), .A(n13959), .ZN(n13960) );
  AOI21_X1 U15929 ( .B1(n14431), .B2(n15197), .A(n13960), .ZN(n13961) );
  OAI21_X1 U15930 ( .B1(n13962), .B2(n14731), .A(n13961), .ZN(P1_U3223) );
  XOR2_X1 U15931 ( .A(n13964), .B(n13963), .Z(n13970) );
  AOI22_X1 U15932 ( .A1(n14705), .A2(n14142), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13966) );
  NAND2_X1 U15933 ( .A1(n14018), .A2(n14137), .ZN(n13965) );
  OAI211_X1 U15934 ( .C1(n13967), .C2(n14728), .A(n13966), .B(n13965), .ZN(
        n13968) );
  AOI21_X1 U15935 ( .B1(n14346), .B2(n15197), .A(n13968), .ZN(n13969) );
  OAI21_X1 U15936 ( .B1(n13970), .B2(n14731), .A(n13969), .ZN(P1_U3225) );
  XOR2_X1 U15937 ( .A(n13972), .B(n13971), .Z(n13977) );
  AOI22_X1 U15938 ( .A1(n14705), .A2(n14196), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13974) );
  NAND2_X1 U15939 ( .A1(n14703), .A2(n14159), .ZN(n13973) );
  OAI211_X1 U15940 ( .C1(n15204), .C2(n14167), .A(n13974), .B(n13973), .ZN(
        n13975) );
  AOI21_X1 U15941 ( .B1(n14351), .B2(n15197), .A(n13975), .ZN(n13976) );
  OAI21_X1 U15942 ( .B1(n13977), .B2(n14731), .A(n13976), .ZN(P1_U3229) );
  OAI211_X1 U15943 ( .C1(n13980), .C2(n13979), .A(n13978), .B(n15206), .ZN(
        n13986) );
  INV_X1 U15944 ( .A(n13981), .ZN(n14224) );
  AND2_X1 U15945 ( .A1(n14197), .A2(n14620), .ZN(n13982) );
  AOI21_X1 U15946 ( .B1(n14259), .B2(n14619), .A(n13982), .ZN(n14222) );
  OAI22_X1 U15947 ( .A1(n14222), .A2(n14015), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13983), .ZN(n13984) );
  AOI21_X1 U15948 ( .B1(n14224), .B2(n14018), .A(n13984), .ZN(n13985) );
  OAI211_X1 U15949 ( .C1(n14437), .C2(n14707), .A(n13986), .B(n13985), .ZN(
        P1_U3233) );
  OAI21_X1 U15950 ( .B1(n13989), .B2(n13988), .A(n13987), .ZN(n13990) );
  NAND2_X1 U15951 ( .A1(n13990), .A2(n15206), .ZN(n13996) );
  INV_X1 U15952 ( .A(n13991), .ZN(n14200) );
  AOI22_X1 U15953 ( .A1(n14705), .A2(n14197), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13992) );
  OAI21_X1 U15954 ( .B1(n13993), .B2(n14728), .A(n13992), .ZN(n13994) );
  AOI21_X1 U15955 ( .B1(n14200), .B2(n14018), .A(n13994), .ZN(n13995) );
  OAI211_X1 U15956 ( .C1(n14707), .C2(n14361), .A(n13996), .B(n13995), .ZN(
        P1_U3235) );
  XOR2_X1 U15957 ( .A(n13998), .B(n13997), .Z(n14004) );
  OAI21_X1 U15958 ( .B1(n14725), .B2(n14714), .A(n13999), .ZN(n14000) );
  AOI21_X1 U15959 ( .B1(n14703), .B2(n14259), .A(n14000), .ZN(n14001) );
  OAI21_X1 U15960 ( .B1(n14264), .B2(n15204), .A(n14001), .ZN(n14002) );
  AOI21_X1 U15961 ( .B1(n14385), .B2(n15197), .A(n14002), .ZN(n14003) );
  OAI21_X1 U15962 ( .B1(n14004), .B2(n14731), .A(n14003), .ZN(P1_U3238) );
  XOR2_X1 U15963 ( .A(n14006), .B(n14005), .Z(n14011) );
  AOI22_X1 U15964 ( .A1(n14619), .A2(n14159), .B1(n14024), .B2(n14620), .ZN(
        n14125) );
  OAI22_X1 U15965 ( .A1(n14015), .A2(n14125), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14007), .ZN(n14008) );
  AOI21_X1 U15966 ( .B1(n14018), .B2(n14131), .A(n14008), .ZN(n14010) );
  NAND2_X1 U15967 ( .A1(n14130), .A2(n15197), .ZN(n14009) );
  OAI211_X1 U15968 ( .C1(n14011), .C2(n14731), .A(n14010), .B(n14009), .ZN(
        P1_U3240) );
  OAI211_X1 U15969 ( .C1(n14014), .C2(n14013), .A(n14012), .B(n15206), .ZN(
        n14021) );
  NAND2_X1 U15970 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14790)
         );
  OAI21_X1 U15971 ( .B1(n14016), .B2(n14015), .A(n14790), .ZN(n14017) );
  AOI21_X1 U15972 ( .B1(n14019), .B2(n14018), .A(n14017), .ZN(n14020) );
  OAI211_X1 U15973 ( .C1(n14447), .C2(n14707), .A(n14021), .B(n14020), .ZN(
        P1_U3241) );
  MUX2_X1 U15974 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14092), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15975 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14022), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15976 ( .A(n14023), .B(P1_DATAO_REG_29__SCAN_IN), .S(n14039), .Z(
        P1_U3589) );
  MUX2_X1 U15977 ( .A(n14107), .B(P1_DATAO_REG_28__SCAN_IN), .S(n14039), .Z(
        P1_U3588) );
  MUX2_X1 U15978 ( .A(n14024), .B(P1_DATAO_REG_27__SCAN_IN), .S(n14039), .Z(
        P1_U3587) );
  MUX2_X1 U15979 ( .A(n14143), .B(P1_DATAO_REG_26__SCAN_IN), .S(n14039), .Z(
        P1_U3586) );
  MUX2_X1 U15980 ( .A(n14159), .B(P1_DATAO_REG_25__SCAN_IN), .S(n14039), .Z(
        P1_U3585) );
  MUX2_X1 U15981 ( .A(n14142), .B(P1_DATAO_REG_24__SCAN_IN), .S(n14039), .Z(
        P1_U3584) );
  MUX2_X1 U15982 ( .A(n14196), .B(P1_DATAO_REG_23__SCAN_IN), .S(n14039), .Z(
        P1_U3583) );
  MUX2_X1 U15983 ( .A(n14025), .B(P1_DATAO_REG_22__SCAN_IN), .S(n14039), .Z(
        P1_U3582) );
  MUX2_X1 U15984 ( .A(n14197), .B(P1_DATAO_REG_21__SCAN_IN), .S(n14039), .Z(
        P1_U3581) );
  MUX2_X1 U15985 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14026), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15986 ( .A(n14259), .B(P1_DATAO_REG_19__SCAN_IN), .S(n14039), .Z(
        P1_U3579) );
  MUX2_X1 U15987 ( .A(n14027), .B(P1_DATAO_REG_18__SCAN_IN), .S(n14039), .Z(
        P1_U3578) );
  MUX2_X1 U15988 ( .A(n14296), .B(P1_DATAO_REG_17__SCAN_IN), .S(n14039), .Z(
        P1_U3577) );
  MUX2_X1 U15989 ( .A(n14028), .B(P1_DATAO_REG_16__SCAN_IN), .S(n14039), .Z(
        P1_U3576) );
  MUX2_X1 U15990 ( .A(n14702), .B(P1_DATAO_REG_15__SCAN_IN), .S(n14039), .Z(
        P1_U3575) );
  MUX2_X1 U15991 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14621), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15992 ( .A(n14704), .B(P1_DATAO_REG_13__SCAN_IN), .S(n14039), .Z(
        P1_U3573) );
  MUX2_X1 U15993 ( .A(n14618), .B(P1_DATAO_REG_12__SCAN_IN), .S(n14039), .Z(
        P1_U3572) );
  MUX2_X1 U15994 ( .A(n14029), .B(P1_DATAO_REG_11__SCAN_IN), .S(n14039), .Z(
        P1_U3571) );
  MUX2_X1 U15995 ( .A(n14030), .B(P1_DATAO_REG_10__SCAN_IN), .S(n14039), .Z(
        P1_U3570) );
  MUX2_X1 U15996 ( .A(n14031), .B(P1_DATAO_REG_9__SCAN_IN), .S(n14039), .Z(
        P1_U3569) );
  MUX2_X1 U15997 ( .A(n14032), .B(P1_DATAO_REG_8__SCAN_IN), .S(n14039), .Z(
        P1_U3568) );
  MUX2_X1 U15998 ( .A(n14033), .B(P1_DATAO_REG_7__SCAN_IN), .S(n14039), .Z(
        P1_U3567) );
  MUX2_X1 U15999 ( .A(n14034), .B(P1_DATAO_REG_6__SCAN_IN), .S(n14039), .Z(
        P1_U3566) );
  MUX2_X1 U16000 ( .A(n14035), .B(P1_DATAO_REG_5__SCAN_IN), .S(n14039), .Z(
        P1_U3565) );
  MUX2_X1 U16001 ( .A(n14036), .B(P1_DATAO_REG_4__SCAN_IN), .S(n14039), .Z(
        P1_U3564) );
  MUX2_X1 U16002 ( .A(n14037), .B(P1_DATAO_REG_3__SCAN_IN), .S(n14039), .Z(
        P1_U3563) );
  MUX2_X1 U16003 ( .A(n14038), .B(P1_DATAO_REG_2__SCAN_IN), .S(n14039), .Z(
        P1_U3562) );
  MUX2_X1 U16004 ( .A(n14040), .B(P1_DATAO_REG_1__SCAN_IN), .S(n14039), .Z(
        P1_U3561) );
  MUX2_X1 U16005 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14041), .S(P1_U4016), .Z(
        P1_U3560) );
  MUX2_X1 U16006 ( .A(n14305), .B(P1_REG2_REG_3__SCAN_IN), .S(n14052), .Z(
        n14044) );
  NAND3_X1 U16007 ( .A1(n14044), .A2(n14043), .A3(n14042), .ZN(n14045) );
  NAND3_X1 U16008 ( .A1(n14074), .A2(n14046), .A3(n14045), .ZN(n14056) );
  MUX2_X1 U16009 ( .A(n10187), .B(P1_REG1_REG_3__SCAN_IN), .S(n14052), .Z(
        n14049) );
  NAND3_X1 U16010 ( .A1(n14049), .A2(n14048), .A3(n14047), .ZN(n14050) );
  NAND3_X1 U16011 ( .A1(n14083), .A2(n14051), .A3(n14050), .ZN(n14055) );
  NAND2_X1 U16012 ( .A1(n14784), .A2(n14052), .ZN(n14054) );
  AOI22_X1 U16013 ( .A1(n14080), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(P1_U3086), .ZN(n14053) );
  NAND4_X1 U16014 ( .A1(n14056), .A2(n14055), .A3(n14054), .A4(n14053), .ZN(
        P1_U3246) );
  INV_X1 U16015 ( .A(n14057), .ZN(n14060) );
  OAI21_X1 U16016 ( .B1(n14792), .B2(n14537), .A(n14058), .ZN(n14059) );
  AOI21_X1 U16017 ( .B1(n14060), .B2(n14784), .A(n14059), .ZN(n14073) );
  INV_X1 U16018 ( .A(n14061), .ZN(n14066) );
  NAND3_X1 U16019 ( .A1(n14064), .A2(n14063), .A3(n14062), .ZN(n14065) );
  NAND3_X1 U16020 ( .A1(n14074), .A2(n14066), .A3(n14065), .ZN(n14072) );
  NAND2_X1 U16021 ( .A1(n14068), .A2(n14067), .ZN(n14069) );
  NAND3_X1 U16022 ( .A1(n14083), .A2(n14070), .A3(n14069), .ZN(n14071) );
  NAND3_X1 U16023 ( .A1(n14073), .A2(n14072), .A3(n14071), .ZN(P1_U3249) );
  NAND2_X1 U16024 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14722)
         );
  OAI211_X1 U16025 ( .C1(n14077), .C2(n14076), .A(n14075), .B(n14074), .ZN(
        n14078) );
  AND2_X1 U16026 ( .A1(n14722), .A2(n14078), .ZN(n14088) );
  INV_X1 U16027 ( .A(n14079), .ZN(n14081) );
  AOI22_X1 U16028 ( .A1(n14784), .A2(n14081), .B1(n14080), .B2(
        P1_ADDR_REG_16__SCAN_IN), .ZN(n14087) );
  OAI211_X1 U16029 ( .C1(n14085), .C2(n14084), .A(n14083), .B(n14082), .ZN(
        n14086) );
  NAND3_X1 U16030 ( .A1(n14088), .A2(n14087), .A3(n14086), .ZN(P1_U3259) );
  NAND2_X1 U16031 ( .A1(n14096), .A2(n14417), .ZN(n14095) );
  XNOR2_X1 U16032 ( .A(n14095), .B(n14413), .ZN(n14090) );
  NAND2_X1 U16033 ( .A1(n14090), .A2(n14814), .ZN(n14316) );
  NAND2_X1 U16034 ( .A1(n14092), .A2(n14091), .ZN(n14319) );
  NOR2_X1 U16035 ( .A1(n14630), .A2(n14319), .ZN(n14098) );
  NOR2_X1 U16036 ( .A1(n14413), .A2(n14307), .ZN(n14093) );
  AOI211_X1 U16037 ( .C1(n14630), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14098), 
        .B(n14093), .ZN(n14094) );
  OAI21_X1 U16038 ( .B1(n14316), .B2(n14300), .A(n14094), .ZN(P1_U3263) );
  OAI211_X1 U16039 ( .C1(n14096), .C2(n14417), .A(n14814), .B(n14095), .ZN(
        n14320) );
  NOR2_X1 U16040 ( .A1(n14417), .A2(n14307), .ZN(n14097) );
  AOI211_X1 U16041 ( .C1(n14630), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14098), 
        .B(n14097), .ZN(n14099) );
  OAI21_X1 U16042 ( .B1(n14300), .B2(n14320), .A(n14099), .ZN(P1_U3264) );
  NOR2_X1 U16043 ( .A1(n14101), .A2(n14100), .ZN(n14102) );
  OR2_X2 U16044 ( .A1(n14103), .A2(n14102), .ZN(n14336) );
  INV_X1 U16045 ( .A(n14336), .ZN(n14122) );
  OAI21_X1 U16046 ( .B1(n14106), .B2(n14105), .A(n14104), .ZN(n14111) );
  NAND2_X1 U16047 ( .A1(n14143), .A2(n14619), .ZN(n14109) );
  NAND2_X1 U16048 ( .A1(n14107), .A2(n14620), .ZN(n14108) );
  NAND2_X1 U16049 ( .A1(n14109), .A2(n14108), .ZN(n14110) );
  AOI21_X1 U16050 ( .B1(n14111), .B2(n14255), .A(n14110), .ZN(n14113) );
  NAND2_X1 U16051 ( .A1(n14340), .A2(n14279), .ZN(n14121) );
  OR2_X1 U16052 ( .A1(n14129), .A2(n14118), .ZN(n14115) );
  AND2_X1 U16053 ( .A1(n14115), .A2(n14114), .ZN(n14338) );
  AOI22_X1 U16054 ( .A1(n14630), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14116), 
        .B2(n14599), .ZN(n14117) );
  OAI21_X1 U16055 ( .B1(n14118), .B2(n14307), .A(n14117), .ZN(n14119) );
  AOI21_X1 U16056 ( .B1(n14338), .B2(n14186), .A(n14119), .ZN(n14120) );
  OAI211_X1 U16057 ( .C1(n14122), .C2(n14171), .A(n14121), .B(n14120), .ZN(
        P1_U3266) );
  XNOR2_X1 U16058 ( .A(n14124), .B(n14123), .ZN(n14126) );
  INV_X1 U16059 ( .A(n14341), .ZN(n14136) );
  XNOR2_X1 U16060 ( .A(n14128), .B(n14127), .ZN(n14343) );
  INV_X1 U16061 ( .A(n14130), .ZN(n14424) );
  AOI211_X1 U16062 ( .C1(n14130), .C2(n14150), .A(n14822), .B(n14129), .ZN(
        n14342) );
  NAND2_X1 U16063 ( .A1(n14342), .A2(n14604), .ZN(n14133) );
  AOI22_X1 U16064 ( .A1(n14630), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n14131), 
        .B2(n14599), .ZN(n14132) );
  OAI211_X1 U16065 ( .C1(n14424), .C2(n14307), .A(n14133), .B(n14132), .ZN(
        n14134) );
  AOI21_X1 U16066 ( .B1(n14631), .B2(n14343), .A(n14134), .ZN(n14135) );
  OAI21_X1 U16067 ( .B1(n14630), .B2(n14136), .A(n14135), .ZN(P1_U3267) );
  INV_X1 U16068 ( .A(n14137), .ZN(n14145) );
  INV_X1 U16069 ( .A(n14138), .ZN(n14141) );
  OAI21_X1 U16070 ( .B1(n14141), .B2(n14140), .A(n14139), .ZN(n14144) );
  AOI222_X1 U16071 ( .A1(n14255), .A2(n14144), .B1(n14143), .B2(n14620), .C1(
        n14142), .C2(n14619), .ZN(n14349) );
  OAI21_X1 U16072 ( .B1(n14145), .B2(n14611), .A(n14349), .ZN(n14154) );
  OAI21_X1 U16073 ( .B1(n14148), .B2(n14147), .A(n14146), .ZN(n14350) );
  AOI22_X1 U16074 ( .A1(n14346), .A2(n14601), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n14630), .ZN(n14152) );
  NAND2_X1 U16075 ( .A1(n14346), .A2(n14166), .ZN(n14149) );
  AND2_X1 U16076 ( .A1(n14150), .A2(n14149), .ZN(n14347) );
  NAND2_X1 U16077 ( .A1(n14347), .A2(n14186), .ZN(n14151) );
  OAI211_X1 U16078 ( .C1(n14350), .C2(n14286), .A(n14152), .B(n14151), .ZN(
        n14153) );
  AOI21_X1 U16079 ( .B1(n14154), .B2(n14279), .A(n14153), .ZN(n14155) );
  INV_X1 U16080 ( .A(n14155), .ZN(P1_U3268) );
  INV_X1 U16081 ( .A(n14156), .ZN(n14157) );
  AOI21_X1 U16082 ( .B1(n14162), .B2(n14158), .A(n14157), .ZN(n14355) );
  AOI22_X1 U16083 ( .A1(n14619), .A2(n14196), .B1(n14159), .B2(n14620), .ZN(
        n14164) );
  OAI211_X1 U16084 ( .C1(n14162), .C2(n14161), .A(n14160), .B(n14255), .ZN(
        n14163) );
  OAI211_X1 U16085 ( .C1(n14355), .C2(n14797), .A(n14164), .B(n14163), .ZN(
        n14165) );
  INV_X1 U16086 ( .A(n14165), .ZN(n14354) );
  AOI21_X1 U16087 ( .B1(n14351), .B2(n14182), .A(n7012), .ZN(n14352) );
  INV_X1 U16088 ( .A(n14351), .ZN(n14170) );
  INV_X1 U16089 ( .A(n14167), .ZN(n14168) );
  AOI22_X1 U16090 ( .A1(n14630), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14168), 
        .B2(n14599), .ZN(n14169) );
  OAI21_X1 U16091 ( .B1(n14170), .B2(n14307), .A(n14169), .ZN(n14173) );
  NOR2_X1 U16092 ( .A1(n14355), .A2(n14171), .ZN(n14172) );
  AOI211_X1 U16093 ( .C1(n14352), .C2(n14186), .A(n14173), .B(n14172), .ZN(
        n14174) );
  OAI21_X1 U16094 ( .B1(n14630), .B2(n14354), .A(n14174), .ZN(P1_U3269) );
  XNOR2_X1 U16095 ( .A(n14175), .B(n14176), .ZN(n14178) );
  AOI21_X1 U16096 ( .B1(n14178), .B2(n14255), .A(n14177), .ZN(n14359) );
  OAI21_X1 U16097 ( .B1(n14179), .B2(n14611), .A(n14359), .ZN(n14180) );
  NAND2_X1 U16098 ( .A1(n14180), .A2(n14279), .ZN(n14188) );
  INV_X1 U16099 ( .A(n14182), .ZN(n14183) );
  AOI21_X1 U16100 ( .B1(n14356), .B2(n14195), .A(n14183), .ZN(n14357) );
  INV_X1 U16101 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14184) );
  OAI22_X1 U16102 ( .A1(n12345), .A2(n14307), .B1(n14184), .B2(n14279), .ZN(
        n14185) );
  AOI21_X1 U16103 ( .B1(n14357), .B2(n14186), .A(n14185), .ZN(n14187) );
  OAI211_X1 U16104 ( .C1(n14286), .C2(n14360), .A(n14188), .B(n14187), .ZN(
        P1_U3270) );
  AOI21_X1 U16105 ( .B1(n14191), .B2(n14189), .A(n6552), .ZN(n14366) );
  OAI21_X1 U16106 ( .B1(n14192), .B2(n14191), .A(n14190), .ZN(n14364) );
  NAND2_X1 U16107 ( .A1(n14193), .A2(n14212), .ZN(n14194) );
  NAND3_X1 U16108 ( .A1(n14195), .A2(n14814), .A3(n14194), .ZN(n14199) );
  AOI22_X1 U16109 ( .A1(n14619), .A2(n14197), .B1(n14196), .B2(n14620), .ZN(
        n14198) );
  NAND2_X1 U16110 ( .A1(n14199), .A2(n14198), .ZN(n14362) );
  NAND3_X1 U16111 ( .A1(n14362), .A2(n14626), .A3(n14279), .ZN(n14202) );
  AOI22_X1 U16112 ( .A1(n14630), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14200), 
        .B2(n14599), .ZN(n14201) );
  OAI211_X1 U16113 ( .C1(n14307), .C2(n14361), .A(n14202), .B(n14201), .ZN(
        n14203) );
  AOI21_X1 U16114 ( .B1(n14364), .B2(n14631), .A(n14203), .ZN(n14204) );
  OAI21_X1 U16115 ( .B1(n14366), .B2(n14303), .A(n14204), .ZN(P1_U3271) );
  XNOR2_X1 U16116 ( .A(n14205), .B(n6771), .ZN(n14369) );
  OAI211_X1 U16117 ( .C1(n14208), .C2(n14207), .A(n14206), .B(n14255), .ZN(
        n14211) );
  INV_X1 U16118 ( .A(n14209), .ZN(n14210) );
  AND2_X1 U16119 ( .A1(n14211), .A2(n14210), .ZN(n14368) );
  INV_X1 U16120 ( .A(n14368), .ZN(n14219) );
  AOI21_X1 U16121 ( .B1(n14228), .B2(n14431), .A(n14822), .ZN(n14213) );
  NAND2_X1 U16122 ( .A1(n14213), .A2(n14212), .ZN(n14367) );
  NAND2_X1 U16123 ( .A1(n14630), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n14214) );
  OAI21_X1 U16124 ( .B1(n14611), .B2(n14215), .A(n14214), .ZN(n14216) );
  AOI21_X1 U16125 ( .B1(n14431), .B2(n14601), .A(n14216), .ZN(n14217) );
  OAI21_X1 U16126 ( .B1(n14367), .B2(n14300), .A(n14217), .ZN(n14218) );
  AOI21_X1 U16127 ( .B1(n14219), .B2(n14279), .A(n14218), .ZN(n14220) );
  OAI21_X1 U16128 ( .B1(n14286), .B2(n14369), .A(n14220), .ZN(P1_U3272) );
  OAI211_X1 U16129 ( .C1(n7561), .C2(n14225), .A(n14221), .B(n14255), .ZN(
        n14223) );
  NAND2_X1 U16130 ( .A1(n14223), .A2(n14222), .ZN(n14374) );
  AOI21_X1 U16131 ( .B1(n14224), .B2(n14599), .A(n14374), .ZN(n14236) );
  NAND2_X1 U16132 ( .A1(n14226), .A2(n14225), .ZN(n14227) );
  AND2_X1 U16133 ( .A1(n7562), .A2(n14227), .ZN(n14375) );
  INV_X1 U16134 ( .A(n14240), .ZN(n14230) );
  INV_X1 U16135 ( .A(n14228), .ZN(n14229) );
  AOI211_X1 U16136 ( .C1(n14231), .C2(n14230), .A(n14822), .B(n14229), .ZN(
        n14373) );
  INV_X1 U16137 ( .A(n14373), .ZN(n14233) );
  AOI22_X1 U16138 ( .A1(n14231), .A2(n14601), .B1(n14630), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n14232) );
  OAI21_X1 U16139 ( .B1(n14233), .B2(n14300), .A(n14232), .ZN(n14234) );
  AOI21_X1 U16140 ( .B1(n14375), .B2(n14631), .A(n14234), .ZN(n14235) );
  OAI21_X1 U16141 ( .B1(n14630), .B2(n14236), .A(n14235), .ZN(P1_U3273) );
  NAND2_X1 U16142 ( .A1(n14237), .A2(n14262), .ZN(n14238) );
  NAND2_X1 U16143 ( .A1(n14238), .A2(n14814), .ZN(n14239) );
  NOR2_X1 U16144 ( .A1(n14240), .A2(n14239), .ZN(n14379) );
  INV_X1 U16145 ( .A(n14241), .ZN(n14242) );
  AOI21_X1 U16146 ( .B1(n14244), .B2(n14243), .A(n14242), .ZN(n14246) );
  OAI21_X1 U16147 ( .B1(n14246), .B2(n14831), .A(n14245), .ZN(n14378) );
  AOI21_X1 U16148 ( .B1(n14379), .B2(n14626), .A(n14378), .ZN(n14253) );
  XNOR2_X1 U16149 ( .A(n14248), .B(n14247), .ZN(n14380) );
  AOI22_X1 U16150 ( .A1(n14630), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14249), 
        .B2(n14599), .ZN(n14250) );
  OAI21_X1 U16151 ( .B1(n7003), .B2(n14307), .A(n14250), .ZN(n14251) );
  AOI21_X1 U16152 ( .B1(n14380), .B2(n14631), .A(n14251), .ZN(n14252) );
  OAI21_X1 U16153 ( .B1(n14253), .B2(n14630), .A(n14252), .ZN(P1_U3274) );
  XNOR2_X1 U16154 ( .A(n6893), .B(n14258), .ZN(n14387) );
  OAI211_X1 U16155 ( .C1(n14258), .C2(n14257), .A(n14256), .B(n14255), .ZN(
        n14261) );
  AOI22_X1 U16156 ( .A1(n14259), .A2(n14620), .B1(n14619), .B2(n14296), .ZN(
        n14260) );
  NAND2_X1 U16157 ( .A1(n14261), .A2(n14260), .ZN(n14383) );
  NAND2_X1 U16158 ( .A1(n14383), .A2(n14279), .ZN(n14269) );
  AOI21_X1 U16159 ( .B1(n14385), .B2(n6617), .A(n14822), .ZN(n14263) );
  AND2_X1 U16160 ( .A1(n14263), .A2(n14262), .ZN(n14384) );
  OAI22_X1 U16161 ( .A1(n14279), .A2(n14265), .B1(n14264), .B2(n14611), .ZN(
        n14267) );
  NOR2_X1 U16162 ( .A1(n12344), .A2(n14307), .ZN(n14266) );
  AOI211_X1 U16163 ( .C1(n14384), .C2(n14604), .A(n14267), .B(n14266), .ZN(
        n14268) );
  OAI211_X1 U16164 ( .C1(n14286), .C2(n14387), .A(n14269), .B(n14268), .ZN(
        P1_U3275) );
  XNOR2_X1 U16165 ( .A(n14271), .B(n14270), .ZN(n14395) );
  AOI21_X1 U16166 ( .B1(n14293), .B2(n14735), .A(n14822), .ZN(n14272) );
  AND2_X1 U16167 ( .A1(n14272), .A2(n6617), .ZN(n14389) );
  NAND2_X1 U16168 ( .A1(n14735), .A2(n14601), .ZN(n14277) );
  OAI22_X1 U16169 ( .A1(n14727), .A2(n14274), .B1(n14726), .B2(n14273), .ZN(
        n14390) );
  INV_X1 U16170 ( .A(n14738), .ZN(n14275) );
  AOI22_X1 U16171 ( .A1(n14390), .A2(n14279), .B1(n14275), .B2(n14599), .ZN(
        n14276) );
  OAI211_X1 U16172 ( .C1(n14279), .C2(n14278), .A(n14277), .B(n14276), .ZN(
        n14280) );
  AOI21_X1 U16173 ( .B1(n14389), .B2(n14604), .A(n14280), .ZN(n14285) );
  NAND2_X1 U16174 ( .A1(n14282), .A2(n14281), .ZN(n14391) );
  NAND3_X1 U16175 ( .A1(n14392), .A2(n14391), .A3(n14283), .ZN(n14284) );
  OAI211_X1 U16176 ( .C1(n14395), .C2(n14286), .A(n14285), .B(n14284), .ZN(
        P1_U3276) );
  INV_X1 U16177 ( .A(n14287), .ZN(n14288) );
  AOI21_X1 U16178 ( .B1(n14291), .B2(n14289), .A(n14288), .ZN(n14402) );
  OAI21_X1 U16179 ( .B1(n14292), .B2(n14291), .A(n14290), .ZN(n14400) );
  OAI211_X1 U16180 ( .C1(n14398), .C2(n14294), .A(n14814), .B(n14293), .ZN(
        n14397) );
  NOR2_X1 U16181 ( .A1(n14279), .A2(n14295), .ZN(n14298) );
  AOI22_X1 U16182 ( .A1(n14296), .A2(n14620), .B1(n14619), .B2(n14702), .ZN(
        n14396) );
  OAI22_X1 U16183 ( .A1(n14630), .A2(n14396), .B1(n14724), .B2(n14611), .ZN(
        n14297) );
  AOI211_X1 U16184 ( .C1(n14721), .C2(n14601), .A(n14298), .B(n14297), .ZN(
        n14299) );
  OAI21_X1 U16185 ( .B1(n14397), .B2(n14300), .A(n14299), .ZN(n14301) );
  AOI21_X1 U16186 ( .B1(n14400), .B2(n14631), .A(n14301), .ZN(n14302) );
  OAI21_X1 U16187 ( .B1(n14402), .B2(n14303), .A(n14302), .ZN(P1_U3277) );
  MUX2_X1 U16188 ( .A(n14305), .B(n14304), .S(n14279), .Z(n14315) );
  OAI22_X1 U16189 ( .A1(n14307), .A2(n14306), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14611), .ZN(n14308) );
  INV_X1 U16190 ( .A(n14308), .ZN(n14314) );
  NAND2_X1 U16191 ( .A1(n14309), .A2(n14605), .ZN(n14313) );
  INV_X1 U16192 ( .A(n14310), .ZN(n14311) );
  NAND2_X1 U16193 ( .A1(n14604), .A2(n14311), .ZN(n14312) );
  NAND4_X1 U16194 ( .A1(n14315), .A2(n14314), .A3(n14313), .A4(n14312), .ZN(
        P1_U3290) );
  AND2_X1 U16195 ( .A1(n14316), .A2(n14319), .ZN(n14411) );
  MUX2_X1 U16196 ( .A(n14317), .B(n14411), .S(n14388), .Z(n14318) );
  OAI21_X1 U16197 ( .B1(n14413), .B2(n14409), .A(n14318), .ZN(P1_U3559) );
  INV_X1 U16198 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n14321) );
  AND2_X1 U16199 ( .A1(n14320), .A2(n14319), .ZN(n14414) );
  MUX2_X1 U16200 ( .A(n14321), .B(n14414), .S(n14388), .Z(n14322) );
  OAI21_X1 U16201 ( .B1(n14417), .B2(n14409), .A(n14322), .ZN(P1_U3558) );
  NAND2_X1 U16202 ( .A1(n14324), .A2(n14323), .ZN(n14326) );
  MUX2_X1 U16203 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14418), .S(n14388), .Z(
        P1_U3557) );
  AOI21_X1 U16204 ( .B1(n14828), .B2(n14330), .A(n14329), .ZN(n14331) );
  MUX2_X1 U16205 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14419), .S(n14388), .Z(
        P1_U3556) );
  AOI22_X1 U16206 ( .A1(n14338), .A2(n14814), .B1(n14828), .B2(n14337), .ZN(
        n14339) );
  MUX2_X1 U16207 ( .A(n14420), .B(P1_REG1_REG_27__SCAN_IN), .S(n14853), .Z(
        P1_U3555) );
  INV_X1 U16208 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n14344) );
  MUX2_X1 U16209 ( .A(n14344), .B(n14421), .S(n14388), .Z(n14345) );
  AOI22_X1 U16210 ( .A1(n14347), .A2(n14814), .B1(n14828), .B2(n14346), .ZN(
        n14348) );
  OAI211_X1 U16211 ( .C1(n14819), .C2(n14350), .A(n14349), .B(n14348), .ZN(
        n14425) );
  MUX2_X1 U16212 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14425), .S(n14388), .Z(
        P1_U3553) );
  AOI22_X1 U16213 ( .A1(n14352), .A2(n14814), .B1(n14828), .B2(n14351), .ZN(
        n14353) );
  OAI211_X1 U16214 ( .C1(n14355), .C2(n14796), .A(n14354), .B(n14353), .ZN(
        n14426) );
  MUX2_X1 U16215 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14426), .S(n14388), .Z(
        P1_U3552) );
  AOI22_X1 U16216 ( .A1(n14357), .A2(n14814), .B1(n14828), .B2(n14356), .ZN(
        n14358) );
  OAI211_X1 U16217 ( .C1(n14819), .C2(n14360), .A(n14359), .B(n14358), .ZN(
        n14427) );
  MUX2_X1 U16218 ( .A(n14427), .B(P1_REG1_REG_23__SCAN_IN), .S(n14853), .Z(
        P1_U3551) );
  NOR2_X1 U16219 ( .A1(n14361), .A2(n14837), .ZN(n14363) );
  AOI211_X1 U16220 ( .C1(n14364), .C2(n14842), .A(n14363), .B(n14362), .ZN(
        n14365) );
  OAI21_X1 U16221 ( .B1(n14366), .B2(n14831), .A(n14365), .ZN(n14428) );
  MUX2_X1 U16222 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14428), .S(n14388), .Z(
        P1_U3550) );
  OAI211_X1 U16223 ( .C1(n14819), .C2(n14369), .A(n14368), .B(n14367), .ZN(
        n14429) );
  MUX2_X1 U16224 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14429), .S(n14388), .Z(
        n14370) );
  AOI21_X1 U16225 ( .B1(n14371), .B2(n14431), .A(n14370), .ZN(n14372) );
  INV_X1 U16226 ( .A(n14372), .ZN(P1_U3549) );
  AOI211_X1 U16227 ( .C1(n14375), .C2(n14842), .A(n14374), .B(n14373), .ZN(
        n14434) );
  MUX2_X1 U16228 ( .A(n14376), .B(n14434), .S(n14388), .Z(n14377) );
  OAI21_X1 U16229 ( .B1(n14437), .B2(n14409), .A(n14377), .ZN(P1_U3548) );
  INV_X1 U16230 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14381) );
  AOI211_X1 U16231 ( .C1(n14842), .C2(n14380), .A(n14379), .B(n14378), .ZN(
        n14438) );
  MUX2_X1 U16232 ( .A(n14381), .B(n14438), .S(n14388), .Z(n14382) );
  OAI21_X1 U16233 ( .B1(n7003), .B2(n14409), .A(n14382), .ZN(P1_U3547) );
  AOI211_X1 U16234 ( .C1(n14828), .C2(n14385), .A(n14384), .B(n14383), .ZN(
        n14386) );
  OAI21_X1 U16235 ( .B1(n14819), .B2(n14387), .A(n14386), .ZN(n14441) );
  MUX2_X1 U16236 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14441), .S(n14388), .Z(
        P1_U3546) );
  AOI211_X1 U16237 ( .C1(n14828), .C2(n14735), .A(n14390), .B(n14389), .ZN(
        n14394) );
  NAND3_X1 U16238 ( .A1(n14392), .A2(n14614), .A3(n14391), .ZN(n14393) );
  OAI211_X1 U16239 ( .C1(n14395), .C2(n14819), .A(n14394), .B(n14393), .ZN(
        n14442) );
  MUX2_X1 U16240 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14442), .S(n14388), .Z(
        P1_U3545) );
  OAI211_X1 U16241 ( .C1(n14398), .C2(n14837), .A(n14397), .B(n14396), .ZN(
        n14399) );
  AOI21_X1 U16242 ( .B1(n14400), .B2(n14842), .A(n14399), .ZN(n14401) );
  OAI21_X1 U16243 ( .B1(n14402), .B2(n14831), .A(n14401), .ZN(n14443) );
  MUX2_X1 U16244 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14443), .S(n14388), .Z(
        P1_U3544) );
  INV_X1 U16245 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14407) );
  NAND2_X1 U16246 ( .A1(n14403), .A2(n14842), .ZN(n14405) );
  AND3_X1 U16247 ( .A1(n14406), .A2(n14405), .A3(n14404), .ZN(n14444) );
  MUX2_X1 U16248 ( .A(n14407), .B(n14444), .S(n14388), .Z(n14408) );
  OAI21_X1 U16249 ( .B1(n14447), .B2(n14409), .A(n14408), .ZN(P1_U3543) );
  INV_X1 U16250 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14410) );
  MUX2_X1 U16251 ( .A(n14411), .B(n14410), .S(n14843), .Z(n14412) );
  OAI21_X1 U16252 ( .B1(n14413), .B2(n14446), .A(n14412), .ZN(P1_U3527) );
  MUX2_X1 U16253 ( .A(n14415), .B(n14414), .S(n14845), .Z(n14416) );
  OAI21_X1 U16254 ( .B1(n14417), .B2(n14446), .A(n14416), .ZN(P1_U3526) );
  MUX2_X1 U16255 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14418), .S(n14845), .Z(
        P1_U3525) );
  MUX2_X1 U16256 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14419), .S(n14845), .Z(
        P1_U3524) );
  OAI21_X1 U16257 ( .B1(n14424), .B2(n14446), .A(n14423), .ZN(P1_U3522) );
  MUX2_X1 U16258 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14425), .S(n14845), .Z(
        P1_U3521) );
  MUX2_X1 U16259 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14426), .S(n14845), .Z(
        P1_U3520) );
  MUX2_X1 U16260 ( .A(n14427), .B(P1_REG0_REG_23__SCAN_IN), .S(n14843), .Z(
        P1_U3519) );
  MUX2_X1 U16261 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14428), .S(n14845), .Z(
        P1_U3518) );
  MUX2_X1 U16262 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14429), .S(n14845), .Z(
        n14430) );
  AOI21_X1 U16263 ( .B1(n14432), .B2(n14431), .A(n14430), .ZN(n14433) );
  INV_X1 U16264 ( .A(n14433), .ZN(P1_U3517) );
  INV_X1 U16265 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n14435) );
  MUX2_X1 U16266 ( .A(n14435), .B(n14434), .S(n14845), .Z(n14436) );
  OAI21_X1 U16267 ( .B1(n14437), .B2(n14446), .A(n14436), .ZN(P1_U3516) );
  MUX2_X1 U16268 ( .A(n14439), .B(n14438), .S(n14845), .Z(n14440) );
  OAI21_X1 U16269 ( .B1(n7003), .B2(n14446), .A(n14440), .ZN(P1_U3515) );
  MUX2_X1 U16270 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14441), .S(n14845), .Z(
        P1_U3513) );
  MUX2_X1 U16271 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14442), .S(n14845), .Z(
        P1_U3510) );
  MUX2_X1 U16272 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14443), .S(n14845), .Z(
        P1_U3507) );
  MUX2_X1 U16273 ( .A(n9594), .B(n14444), .S(n14845), .Z(n14445) );
  OAI21_X1 U16274 ( .B1(n14447), .B2(n14446), .A(n14445), .ZN(P1_U3504) );
  NOR4_X1 U16275 ( .A1(n14448), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9292), .A4(
        P1_U3086), .ZN(n14449) );
  AOI21_X1 U16276 ( .B1(n14450), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14449), 
        .ZN(n14451) );
  OAI21_X1 U16277 ( .B1(n14452), .B2(n14472), .A(n14451), .ZN(P1_U3324) );
  OAI222_X1 U16278 ( .A1(n14474), .A2(n14455), .B1(n14472), .B2(n14454), .C1(
        n14453), .C2(P1_U3086), .ZN(P1_U3326) );
  OAI222_X1 U16279 ( .A1(n14474), .A2(n14458), .B1(n14464), .B2(n14457), .C1(
        P1_U3086), .C2(n14456), .ZN(P1_U3327) );
  INV_X1 U16280 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14461) );
  OAI222_X1 U16281 ( .A1(n14474), .A2(n14461), .B1(n14472), .B2(n14460), .C1(
        n14459), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U16282 ( .A1(P1_U3086), .A2(n14465), .B1(n14464), .B2(n14463), 
        .C1(n14462), .C2(n14474), .ZN(P1_U3329) );
  INV_X1 U16283 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14468) );
  OAI222_X1 U16284 ( .A1(n14474), .A2(n14468), .B1(n14472), .B2(n14467), .C1(
        P1_U3086), .C2(n14466), .ZN(P1_U3330) );
  OAI222_X1 U16285 ( .A1(n14474), .A2(n14473), .B1(n14472), .B2(n14471), .C1(
        P1_U3086), .C2(n14469), .ZN(P1_U3331) );
  MUX2_X1 U16286 ( .A(n14476), .B(n14475), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U16287 ( .A(n14477), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16288 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14510) );
  INV_X1 U16289 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14508) );
  XNOR2_X1 U16290 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n14508), .ZN(n14574) );
  INV_X1 U16291 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14506) );
  INV_X1 U16292 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14793) );
  XOR2_X1 U16293 ( .A(n14793), .B(P3_ADDR_REG_15__SCAN_IN), .Z(n14571) );
  XOR2_X1 U16294 ( .A(n14501), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n14513) );
  XOR2_X1 U16295 ( .A(n14499), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n14560) );
  INV_X1 U16296 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15045) );
  NAND2_X1 U16297 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n10026), .ZN(n14527) );
  INV_X1 U16298 ( .A(n14522), .ZN(n14483) );
  NOR2_X1 U16299 ( .A1(n14484), .A2(n6898), .ZN(n14486) );
  NOR2_X1 U16300 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14537), .ZN(n14487) );
  NOR2_X1 U16301 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14488), .ZN(n14490) );
  XOR2_X1 U16302 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n14488), .Z(n14520) );
  XNOR2_X1 U16303 ( .A(n15045), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n14545) );
  XOR2_X1 U16304 ( .A(n15067), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n14550) );
  NAND2_X1 U16305 ( .A1(n14551), .A2(n14550), .ZN(n14492) );
  NAND2_X1 U16306 ( .A1(n14517), .A2(n14519), .ZN(n14494) );
  NOR2_X1 U16307 ( .A1(n14517), .A2(n14519), .ZN(n14493) );
  XOR2_X1 U16308 ( .A(n14497), .B(P1_ADDR_REG_11__SCAN_IN), .Z(n14516) );
  NAND2_X1 U16309 ( .A1(n14515), .A2(n14516), .ZN(n14496) );
  NAND2_X1 U16310 ( .A1(n14560), .A2(n14561), .ZN(n14498) );
  NAND2_X1 U16311 ( .A1(n14513), .A2(n14514), .ZN(n14500) );
  INV_X1 U16312 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14502) );
  XNOR2_X1 U16313 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n14502), .ZN(n14511) );
  NAND2_X1 U16314 ( .A1(n14571), .A2(n14570), .ZN(n14505) );
  NOR2_X1 U16315 ( .A1(n14574), .A2(n14573), .ZN(n14507) );
  AOI21_X1 U16316 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(n14508), .A(n14507), 
        .ZN(n14578) );
  XNOR2_X1 U16317 ( .A(n14510), .B(P1_ADDR_REG_17__SCAN_IN), .ZN(n14577) );
  NOR2_X1 U16318 ( .A1(n14578), .A2(n14577), .ZN(n14509) );
  AOI21_X1 U16319 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(n14510), .A(n14509), 
        .ZN(n14642) );
  INV_X1 U16320 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15356) );
  XNOR2_X1 U16321 ( .A(n15356), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(n14641) );
  XNOR2_X1 U16322 ( .A(n14512), .B(n14511), .ZN(n14766) );
  XOR2_X1 U16323 ( .A(n14514), .B(n14513), .Z(n14565) );
  XNOR2_X1 U16324 ( .A(n14517), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n14518) );
  XNOR2_X1 U16325 ( .A(n14519), .B(n14518), .ZN(n14555) );
  INV_X1 U16326 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14596) );
  XNOR2_X1 U16327 ( .A(n14520), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15401) );
  NAND2_X1 U16328 ( .A1(n14531), .A2(n14532), .ZN(n14533) );
  XOR2_X1 U16329 ( .A(n14523), .B(P1_ADDR_REG_3__SCAN_IN), .Z(n15404) );
  XOR2_X1 U16330 ( .A(n14525), .B(n14524), .Z(n14586) );
  NOR2_X1 U16331 ( .A1(n14528), .A2(n10147), .ZN(n14529) );
  OAI21_X1 U16332 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n10026), .A(n14527), .ZN(
        n15398) );
  NAND2_X1 U16333 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15398), .ZN(n15408) );
  NOR2_X1 U16334 ( .A1(n14586), .A2(n14585), .ZN(n14530) );
  NAND2_X1 U16335 ( .A1(n14586), .A2(n14585), .ZN(n14584) );
  NAND2_X1 U16336 ( .A1(n15395), .A2(n15394), .ZN(n15393) );
  NAND2_X1 U16337 ( .A1(n14534), .A2(n14535), .ZN(n14536) );
  INV_X1 U16338 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15396) );
  XOR2_X1 U16339 ( .A(n14537), .B(P3_ADDR_REG_6__SCAN_IN), .Z(n14539) );
  XNOR2_X1 U16340 ( .A(n14539), .B(n14538), .ZN(n14589) );
  NOR2_X1 U16341 ( .A1(n14541), .A2(n14540), .ZN(n14542) );
  XNOR2_X1 U16342 ( .A(n14546), .B(n14545), .ZN(n14547) );
  NAND2_X1 U16343 ( .A1(n14548), .A2(n14547), .ZN(n14549) );
  INV_X1 U16344 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14592) );
  XOR2_X1 U16345 ( .A(n14551), .B(n14550), .Z(n14553) );
  NOR2_X1 U16346 ( .A1(n14553), .A2(n14552), .ZN(n14554) );
  NAND2_X1 U16347 ( .A1(n14555), .A2(n14557), .ZN(n14558) );
  INV_X1 U16348 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15332) );
  INV_X1 U16349 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14559) );
  XOR2_X1 U16350 ( .A(n14561), .B(n14560), .Z(n14563) );
  NAND2_X1 U16351 ( .A1(n14563), .A2(n14562), .ZN(n14564) );
  NAND2_X1 U16352 ( .A1(n14565), .A2(n14567), .ZN(n14568) );
  INV_X1 U16353 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14762) );
  NAND2_X1 U16354 ( .A1(n14763), .A2(n14762), .ZN(n14761) );
  INV_X1 U16355 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14569) );
  XNOR2_X1 U16356 ( .A(n14571), .B(n14570), .ZN(n14572) );
  INV_X1 U16357 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14772) );
  INV_X1 U16358 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14575) );
  XNOR2_X1 U16359 ( .A(n14578), .B(n14577), .ZN(n14635) );
  INV_X1 U16360 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14579) );
  NAND2_X1 U16361 ( .A1(n14636), .A2(n14635), .ZN(n14634) );
  OAI21_X1 U16362 ( .B1(n14639), .B2(n14638), .A(n14640), .ZN(n14581) );
  XNOR2_X1 U16363 ( .A(n14581), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16364 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14582) );
  OAI21_X1 U16365 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14582), 
        .ZN(U28) );
  AOI21_X1 U16366 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14583) );
  OAI21_X1 U16367 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14583), 
        .ZN(U29) );
  OAI21_X1 U16368 ( .B1(n14586), .B2(n14585), .A(n14584), .ZN(n14587) );
  XNOR2_X1 U16369 ( .A(n14587), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16370 ( .B1(n14590), .B2(n14589), .A(n14588), .ZN(SUB_1596_U57) );
  OAI21_X1 U16371 ( .B1(n14593), .B2(n14592), .A(n14591), .ZN(SUB_1596_U55) );
  AOI21_X1 U16372 ( .B1(n14596), .B2(n14595), .A(n14594), .ZN(SUB_1596_U54) );
  OAI21_X1 U16373 ( .B1(n14598), .B2(n15332), .A(n14597), .ZN(SUB_1596_U70) );
  AOI222_X1 U16374 ( .A1(n14602), .A2(n14601), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n14630), .C1(n14600), .C2(n14599), .ZN(n14608) );
  AOI22_X1 U16375 ( .A1(n14606), .A2(n14605), .B1(n14604), .B2(n14603), .ZN(
        n14607) );
  OAI211_X1 U16376 ( .C1(n14630), .C2(n14609), .A(n14608), .B(n14607), .ZN(
        P1_U3281) );
  OAI211_X1 U16377 ( .C1(n14745), .C2(n6627), .A(n14814), .B(n14610), .ZN(
        n14747) );
  INV_X1 U16378 ( .A(n14747), .ZN(n14627) );
  OAI22_X1 U16379 ( .A1(n14745), .A2(n14613), .B1(n14612), .B2(n14611), .ZN(
        n14625) );
  OAI211_X1 U16380 ( .C1(n14617), .C2(n14616), .A(n14615), .B(n14614), .ZN(
        n14623) );
  AOI22_X1 U16381 ( .A1(n14621), .A2(n14620), .B1(n14619), .B2(n14618), .ZN(
        n14622) );
  AND2_X1 U16382 ( .A1(n14623), .A2(n14622), .ZN(n14750) );
  INV_X1 U16383 ( .A(n14750), .ZN(n14624) );
  AOI211_X1 U16384 ( .C1(n14627), .C2(n14626), .A(n14625), .B(n14624), .ZN(
        n14633) );
  XNOR2_X1 U16385 ( .A(n14629), .B(n14628), .ZN(n14744) );
  AOI22_X1 U16386 ( .A1(n14744), .A2(n14631), .B1(P1_REG2_REG_13__SCAN_IN), 
        .B2(n14630), .ZN(n14632) );
  OAI21_X1 U16387 ( .B1(n14630), .B2(n14633), .A(n14632), .ZN(P1_U3280) );
  OAI21_X1 U16388 ( .B1(n14636), .B2(n14635), .A(n14634), .ZN(n14637) );
  XNOR2_X1 U16389 ( .A(n14637), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  NOR2_X1 U16390 ( .A1(n14642), .A2(n14641), .ZN(n14643) );
  AOI21_X1 U16391 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15356), .A(n14643), 
        .ZN(n14644) );
  XOR2_X1 U16392 ( .A(n14645), .B(n14649), .Z(n14646) );
  OAI222_X1 U16393 ( .A1(n15095), .A2(n14647), .B1(n15094), .B2(n14675), .C1(
        n14646), .C2(n15078), .ZN(n14681) );
  OAI22_X1 U16394 ( .A1(n15122), .A2(n12716), .B1(n15089), .B2(n14648), .ZN(
        n14654) );
  XNOR2_X1 U16395 ( .A(n14650), .B(n14649), .ZN(n14683) );
  NOR2_X1 U16396 ( .A1(n14651), .A2(n15169), .ZN(n14682) );
  AOI22_X1 U16397 ( .A1(n14683), .A2(n14664), .B1(n15083), .B2(n14682), .ZN(
        n14652) );
  INV_X1 U16398 ( .A(n14652), .ZN(n14653) );
  AOI211_X1 U16399 ( .C1(n15122), .C2(n14681), .A(n14654), .B(n14653), .ZN(
        n14655) );
  INV_X1 U16400 ( .A(n14655), .ZN(P3_U3220) );
  XNOR2_X1 U16401 ( .A(n14656), .B(n14661), .ZN(n14659) );
  AOI222_X1 U16402 ( .A1(n15112), .A2(n14659), .B1(n14658), .B2(n15106), .C1(
        n14657), .C2(n15109), .ZN(n14684) );
  AOI22_X1 U16403 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n15124), .B1(n15119), 
        .B2(n14660), .ZN(n14666) );
  XNOR2_X1 U16404 ( .A(n14662), .B(n14661), .ZN(n14687) );
  NOR2_X1 U16405 ( .A1(n14663), .A2(n15169), .ZN(n14686) );
  AOI22_X1 U16406 ( .A1(n14687), .A2(n14664), .B1(n15083), .B2(n14686), .ZN(
        n14665) );
  OAI211_X1 U16407 ( .C1(n15124), .C2(n14684), .A(n14666), .B(n14665), .ZN(
        P3_U3221) );
  INV_X1 U16408 ( .A(n14667), .ZN(n14670) );
  OAI21_X1 U16409 ( .B1(n14670), .B2(n14669), .A(n14668), .ZN(n14691) );
  XNOR2_X1 U16410 ( .A(n14672), .B(n14671), .ZN(n14673) );
  OAI222_X1 U16411 ( .A1(n15095), .A2(n14675), .B1(n15094), .B2(n14674), .C1(
        n14673), .C2(n15078), .ZN(n14689) );
  AOI21_X1 U16412 ( .B1(n14676), .B2(n14691), .A(n14689), .ZN(n14680) );
  NOR2_X1 U16413 ( .A1(n14677), .A2(n15169), .ZN(n14690) );
  AOI22_X1 U16414 ( .A1(n14690), .A2(n15083), .B1(n14678), .B2(n15119), .ZN(
        n14679) );
  OAI221_X1 U16415 ( .B1(n15124), .B2(n14680), .C1(n15122), .C2(n8454), .A(
        n14679), .ZN(P3_U3222) );
  AOI211_X1 U16416 ( .C1(n14683), .C2(n14692), .A(n14682), .B(n14681), .ZN(
        n14695) );
  AOI22_X1 U16417 ( .A1(n15193), .A2(n14695), .B1(n12715), .B2(n15190), .ZN(
        P3_U3472) );
  INV_X1 U16418 ( .A(n14684), .ZN(n14685) );
  AOI211_X1 U16419 ( .C1(n14687), .C2(n14692), .A(n14686), .B(n14685), .ZN(
        n14697) );
  AOI22_X1 U16420 ( .A1(n15193), .A2(n14697), .B1(n14688), .B2(n15190), .ZN(
        P3_U3471) );
  AOI211_X1 U16421 ( .C1(n14692), .C2(n14691), .A(n14690), .B(n14689), .ZN(
        n14698) );
  AOI22_X1 U16422 ( .A1(n15193), .A2(n14698), .B1(n14693), .B2(n15190), .ZN(
        P3_U3470) );
  INV_X1 U16423 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14694) );
  AOI22_X1 U16424 ( .A1(n15176), .A2(n14695), .B1(n14694), .B2(n15174), .ZN(
        P3_U3429) );
  INV_X1 U16425 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14696) );
  AOI22_X1 U16426 ( .A1(n15176), .A2(n14697), .B1(n14696), .B2(n15174), .ZN(
        P3_U3426) );
  AOI22_X1 U16427 ( .A1(n15176), .A2(n14698), .B1(n8453), .B2(n15174), .ZN(
        P3_U3423) );
  OAI21_X1 U16428 ( .B1(n14701), .B2(n14700), .A(n14699), .ZN(n14709) );
  AOI22_X1 U16429 ( .A1(n14705), .A2(n14704), .B1(n14703), .B2(n14702), .ZN(
        n14706) );
  OAI21_X1 U16430 ( .B1(n7008), .B2(n14707), .A(n14706), .ZN(n14708) );
  AOI21_X1 U16431 ( .B1(n14709), .B2(n15206), .A(n14708), .ZN(n14711) );
  OAI211_X1 U16432 ( .C1(n15204), .C2(n14712), .A(n14711), .B(n14710), .ZN(
        P1_U3215) );
  OAI22_X1 U16433 ( .A1(n14728), .A2(n14714), .B1(n14713), .B2(n14725), .ZN(
        n14720) );
  INV_X1 U16434 ( .A(n14716), .ZN(n14718) );
  AOI21_X1 U16435 ( .B1(n14718), .B2(n14717), .A(n14731), .ZN(n14719) );
  AOI211_X1 U16436 ( .C1(n14721), .C2(n15197), .A(n14720), .B(n14719), .ZN(
        n14723) );
  OAI211_X1 U16437 ( .C1(n15204), .C2(n14724), .A(n14723), .B(n14722), .ZN(
        P1_U3226) );
  OAI22_X1 U16438 ( .A1(n14728), .A2(n14727), .B1(n14726), .B2(n14725), .ZN(
        n14734) );
  XOR2_X1 U16439 ( .A(n14730), .B(n14729), .Z(n14732) );
  NOR2_X1 U16440 ( .A1(n14732), .A2(n14731), .ZN(n14733) );
  AOI211_X1 U16441 ( .C1(n14735), .C2(n15197), .A(n14734), .B(n14733), .ZN(
        n14737) );
  OAI211_X1 U16442 ( .C1(n15204), .C2(n14738), .A(n14737), .B(n14736), .ZN(
        P1_U3228) );
  OAI22_X1 U16443 ( .A1(n14739), .A2(n14822), .B1(n7008), .B2(n14837), .ZN(
        n14741) );
  AOI211_X1 U16444 ( .C1(n14742), .C2(n14842), .A(n14741), .B(n14740), .ZN(
        n14752) );
  AOI22_X1 U16445 ( .A1(n14388), .A2(n14752), .B1(n14743), .B2(n14853), .ZN(
        P1_U3542) );
  NAND2_X1 U16446 ( .A1(n14744), .A2(n14842), .ZN(n14749) );
  OR2_X1 U16447 ( .A1(n14745), .A2(n14837), .ZN(n14746) );
  AND2_X1 U16448 ( .A1(n14747), .A2(n14746), .ZN(n14748) );
  AND3_X1 U16449 ( .A1(n14750), .A2(n14749), .A3(n14748), .ZN(n14753) );
  AOI22_X1 U16450 ( .A1(n14388), .A2(n14753), .B1(n14751), .B2(n14853), .ZN(
        P1_U3541) );
  AOI22_X1 U16451 ( .A1(n14845), .A2(n14752), .B1(n9581), .B2(n14843), .ZN(
        P1_U3501) );
  AOI22_X1 U16452 ( .A1(n14845), .A2(n14753), .B1(n9555), .B2(n14843), .ZN(
        P1_U3498) );
  OAI21_X1 U16453 ( .B1(n14756), .B2(n14755), .A(n14754), .ZN(n14757) );
  XNOR2_X1 U16454 ( .A(n14757), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI21_X1 U16455 ( .B1(n14760), .B2(n14759), .A(n14758), .ZN(SUB_1596_U68) );
  OAI21_X1 U16456 ( .B1(n14763), .B2(n14762), .A(n14761), .ZN(SUB_1596_U67) );
  OAI21_X1 U16457 ( .B1(n14766), .B2(n14765), .A(n14764), .ZN(n14767) );
  XNOR2_X1 U16458 ( .A(n14767), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI222_X1 U16459 ( .A1(n14772), .A2(n14771), .B1(n14772), .B2(n14770), .C1(
        n14769), .C2(n14768), .ZN(SUB_1596_U65) );
  OAI21_X1 U16460 ( .B1(n14775), .B2(n14774), .A(n14773), .ZN(n14776) );
  XNOR2_X1 U16461 ( .A(n14776), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  AOI21_X1 U16462 ( .B1(n14778), .B2(P1_REG1_REG_15__SCAN_IN), .A(n14777), 
        .ZN(n14788) );
  AOI21_X1 U16463 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14780), .A(n14779), 
        .ZN(n14782) );
  OR2_X1 U16464 ( .A1(n14782), .A2(n14781), .ZN(n14786) );
  NAND2_X1 U16465 ( .A1(n14784), .A2(n14783), .ZN(n14785) );
  OAI211_X1 U16466 ( .C1(n14788), .C2(n14787), .A(n14786), .B(n14785), .ZN(
        n14789) );
  INV_X1 U16467 ( .A(n14789), .ZN(n14791) );
  OAI211_X1 U16468 ( .C1(n14793), .C2(n14792), .A(n14791), .B(n14790), .ZN(
        P1_U3258) );
  AND2_X1 U16469 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14794), .ZN(P1_U3294) );
  AND2_X1 U16470 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14794), .ZN(P1_U3295) );
  AND2_X1 U16471 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14794), .ZN(P1_U3296) );
  AND2_X1 U16472 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14794), .ZN(P1_U3297) );
  AND2_X1 U16473 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14794), .ZN(P1_U3298) );
  AND2_X1 U16474 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14794), .ZN(P1_U3299) );
  AND2_X1 U16475 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14794), .ZN(P1_U3300) );
  AND2_X1 U16476 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14794), .ZN(P1_U3301) );
  AND2_X1 U16477 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14794), .ZN(P1_U3302) );
  AND2_X1 U16478 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14794), .ZN(P1_U3303) );
  AND2_X1 U16479 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14794), .ZN(P1_U3304) );
  AND2_X1 U16480 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14794), .ZN(P1_U3305) );
  AND2_X1 U16481 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14794), .ZN(P1_U3306) );
  AND2_X1 U16482 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14794), .ZN(P1_U3307) );
  AND2_X1 U16483 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14794), .ZN(P1_U3308) );
  AND2_X1 U16484 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14794), .ZN(P1_U3309) );
  AND2_X1 U16485 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n6644), .ZN(P1_U3310) );
  AND2_X1 U16486 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n6644), .ZN(P1_U3311) );
  AND2_X1 U16487 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n6644), .ZN(P1_U3312) );
  AND2_X1 U16488 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n6644), .ZN(P1_U3313) );
  AND2_X1 U16489 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n6644), .ZN(P1_U3314) );
  AND2_X1 U16490 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n6644), .ZN(P1_U3315) );
  AND2_X1 U16491 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n6644), .ZN(P1_U3316) );
  AND2_X1 U16492 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n6644), .ZN(P1_U3317) );
  AND2_X1 U16493 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n6644), .ZN(P1_U3318) );
  AND2_X1 U16494 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n6644), .ZN(P1_U3319) );
  AND2_X1 U16495 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n6644), .ZN(P1_U3320) );
  AND2_X1 U16496 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n6644), .ZN(P1_U3321) );
  AND2_X1 U16497 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n6644), .ZN(P1_U3322) );
  AND2_X1 U16498 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n6644), .ZN(P1_U3323) );
  AOI21_X1 U16499 ( .B1(n14797), .B2(n14796), .A(n14795), .ZN(n14806) );
  NOR3_X1 U16500 ( .A1(n14799), .A2(n14798), .A3(n14831), .ZN(n14805) );
  INV_X1 U16501 ( .A(n14800), .ZN(n14801) );
  OAI21_X1 U16502 ( .B1(n14802), .B2(n14837), .A(n14801), .ZN(n14803) );
  NOR4_X1 U16503 ( .A1(n14806), .A2(n14805), .A3(n14804), .A4(n14803), .ZN(
        n14846) );
  AOI22_X1 U16504 ( .A1(n14845), .A2(n14846), .B1(n9355), .B2(n14843), .ZN(
        P1_U3462) );
  AOI211_X1 U16505 ( .C1(n14828), .C2(n14809), .A(n14808), .B(n14807), .ZN(
        n14810) );
  OAI21_X1 U16506 ( .B1(n14819), .B2(n14811), .A(n14810), .ZN(n14812) );
  INV_X1 U16507 ( .A(n14812), .ZN(n14847) );
  AOI22_X1 U16508 ( .A1(n14845), .A2(n14847), .B1(n9388), .B2(n14843), .ZN(
        P1_U3471) );
  AOI22_X1 U16509 ( .A1(n14815), .A2(n14814), .B1(n14828), .B2(n14813), .ZN(
        n14816) );
  OAI211_X1 U16510 ( .C1(n14819), .C2(n14818), .A(n14817), .B(n14816), .ZN(
        n14820) );
  INV_X1 U16511 ( .A(n14820), .ZN(n14849) );
  AOI22_X1 U16512 ( .A1(n14845), .A2(n14849), .B1(n9411), .B2(n14843), .ZN(
        P1_U3474) );
  OAI22_X1 U16513 ( .A1(n14823), .A2(n14822), .B1(n14821), .B2(n14837), .ZN(
        n14825) );
  AOI211_X1 U16514 ( .C1(n14827), .C2(n14826), .A(n14825), .B(n14824), .ZN(
        n14850) );
  AOI22_X1 U16515 ( .A1(n14845), .A2(n14850), .B1(n9445), .B2(n14843), .ZN(
        P1_U3480) );
  AOI21_X1 U16516 ( .B1(n15198), .B2(n14828), .A(n15199), .ZN(n14830) );
  OAI211_X1 U16517 ( .C1(n14832), .C2(n14831), .A(n14830), .B(n14829), .ZN(
        n14833) );
  AOI21_X1 U16518 ( .B1(n14834), .B2(n14842), .A(n14833), .ZN(n14852) );
  INV_X1 U16519 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14835) );
  AOI22_X1 U16520 ( .A1(n14845), .A2(n14852), .B1(n14835), .B2(n14843), .ZN(
        P1_U3483) );
  OAI21_X1 U16521 ( .B1(n14838), .B2(n14837), .A(n14836), .ZN(n14840) );
  AOI211_X1 U16522 ( .C1(n14842), .C2(n14841), .A(n14840), .B(n14839), .ZN(
        n14855) );
  INV_X1 U16523 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14844) );
  AOI22_X1 U16524 ( .A1(n14845), .A2(n14855), .B1(n14844), .B2(n14843), .ZN(
        P1_U3489) );
  AOI22_X1 U16525 ( .A1(n14388), .A2(n14846), .B1(n10162), .B2(n14853), .ZN(
        P1_U3529) );
  AOI22_X1 U16526 ( .A1(n14388), .A2(n14847), .B1(n10196), .B2(n14853), .ZN(
        P1_U3532) );
  AOI22_X1 U16527 ( .A1(n14388), .A2(n14849), .B1(n14848), .B2(n14853), .ZN(
        P1_U3533) );
  AOI22_X1 U16528 ( .A1(n14388), .A2(n14850), .B1(n10201), .B2(n14853), .ZN(
        P1_U3535) );
  AOI22_X1 U16529 ( .A1(n14388), .A2(n14852), .B1(n14851), .B2(n14853), .ZN(
        P1_U3536) );
  AOI22_X1 U16530 ( .A1(n14388), .A2(n14855), .B1(n14854), .B2(n14853), .ZN(
        P1_U3538) );
  NOR2_X1 U16531 ( .A1(n14935), .A2(n14856), .ZN(P2_U3087) );
  OAI21_X1 U16532 ( .B1(n14859), .B2(n14858), .A(n14857), .ZN(n14866) );
  OAI211_X1 U16533 ( .C1(n14863), .C2(n14862), .A(n14861), .B(n14860), .ZN(
        n14864) );
  INV_X1 U16534 ( .A(n14864), .ZN(n14865) );
  AOI211_X1 U16535 ( .C1(n14868), .C2(n14867), .A(n14866), .B(n14865), .ZN(
        n14869) );
  OAI21_X1 U16536 ( .B1(n14871), .B2(n14870), .A(n14869), .ZN(P2_U3206) );
  AOI21_X1 U16537 ( .B1(n14943), .B2(P2_REG1_REG_0__SCAN_IN), .A(n14872), .ZN(
        n14878) );
  AOI22_X1 U16538 ( .A1(n14935), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14877) );
  OAI22_X1 U16539 ( .A1(n14874), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n14873), .ZN(n14875) );
  OAI21_X1 U16540 ( .B1(n14936), .B2(n14875), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n14876) );
  OAI211_X1 U16541 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n14878), .A(n14877), .B(
        n14876), .ZN(P2_U3214) );
  OAI22_X1 U16542 ( .A1(n14880), .A2(n14879), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7774), .ZN(n14881) );
  AOI21_X1 U16543 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n14935), .A(n14881), .ZN(
        n14890) );
  OAI211_X1 U16544 ( .C1(n14884), .C2(n14883), .A(n14939), .B(n14882), .ZN(
        n14889) );
  OAI211_X1 U16545 ( .C1(n14887), .C2(n14886), .A(n14943), .B(n14885), .ZN(
        n14888) );
  NAND3_X1 U16546 ( .A1(n14890), .A2(n14889), .A3(n14888), .ZN(P2_U3217) );
  INV_X1 U16547 ( .A(n14891), .ZN(n14893) );
  OAI21_X1 U16548 ( .B1(n14893), .B2(n14892), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14894) );
  OAI21_X1 U16549 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n14894), .ZN(n14904) );
  OAI211_X1 U16550 ( .C1(n14897), .C2(n14896), .A(n14895), .B(n14939), .ZN(
        n14903) );
  NAND2_X1 U16551 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n14935), .ZN(n14902) );
  OAI211_X1 U16552 ( .C1(n14900), .C2(n14899), .A(n14898), .B(n14943), .ZN(
        n14901) );
  NAND4_X1 U16553 ( .A1(n14904), .A2(n14903), .A3(n14902), .A4(n14901), .ZN(
        P2_U3224) );
  AOI22_X1 U16554 ( .A1(n14935), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3088), .ZN(n14914) );
  NAND2_X1 U16555 ( .A1(n14905), .A2(n14936), .ZN(n14913) );
  OAI211_X1 U16556 ( .C1(n14908), .C2(n14907), .A(n14906), .B(n14943), .ZN(
        n14912) );
  OAI211_X1 U16557 ( .C1(n14910), .C2(P2_REG2_REG_14__SCAN_IN), .A(n14909), 
        .B(n14939), .ZN(n14911) );
  NAND4_X1 U16558 ( .A1(n14914), .A2(n14913), .A3(n14912), .A4(n14911), .ZN(
        P2_U3228) );
  AOI22_X1 U16559 ( .A1(n14935), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14923) );
  NAND2_X1 U16560 ( .A1(n14936), .A2(n14915), .ZN(n14922) );
  OAI211_X1 U16561 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n14917), .A(n14939), 
        .B(n14916), .ZN(n14921) );
  OAI211_X1 U16562 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n14919), .A(n14943), 
        .B(n14918), .ZN(n14920) );
  NAND4_X1 U16563 ( .A1(n14923), .A2(n14922), .A3(n14921), .A4(n14920), .ZN(
        P2_U3229) );
  AOI22_X1 U16564 ( .A1(n14935), .A2(P2_ADDR_REG_16__SCAN_IN), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(P2_U3088), .ZN(n14934) );
  NAND2_X1 U16565 ( .A1(n14936), .A2(n14924), .ZN(n14933) );
  OAI211_X1 U16566 ( .C1(n14927), .C2(n14926), .A(n14939), .B(n14925), .ZN(
        n14932) );
  OAI211_X1 U16567 ( .C1(n14930), .C2(n14929), .A(n14943), .B(n14928), .ZN(
        n14931) );
  NAND4_X1 U16568 ( .A1(n14934), .A2(n14933), .A3(n14932), .A4(n14931), .ZN(
        P2_U3230) );
  AOI22_X1 U16569 ( .A1(n14935), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3088), .ZN(n14949) );
  NAND2_X1 U16570 ( .A1(n14937), .A2(n14936), .ZN(n14948) );
  OAI211_X1 U16571 ( .C1(n14941), .C2(n14940), .A(n14939), .B(n14938), .ZN(
        n14947) );
  OAI211_X1 U16572 ( .C1(n14945), .C2(n14944), .A(n14943), .B(n14942), .ZN(
        n14946) );
  NAND4_X1 U16573 ( .A1(n14949), .A2(n14948), .A3(n14947), .A4(n14946), .ZN(
        P2_U3231) );
  OAI22_X1 U16574 ( .A1(n14952), .A2(n10064), .B1(n14951), .B2(n14950), .ZN(
        n14953) );
  AOI21_X1 U16575 ( .B1(n14955), .B2(n14954), .A(n14953), .ZN(n14956) );
  OAI21_X1 U16576 ( .B1(n14958), .B2(n14957), .A(n14956), .ZN(n14959) );
  AOI21_X1 U16577 ( .B1(n14961), .B2(n14960), .A(n14959), .ZN(n14962) );
  OAI21_X1 U16578 ( .B1(n14964), .B2(n14963), .A(n14962), .ZN(P2_U3258) );
  AND2_X1 U16579 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14967), .ZN(P2_U3266) );
  AND2_X1 U16580 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14967), .ZN(P2_U3267) );
  AND2_X1 U16581 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14967), .ZN(P2_U3268) );
  AND2_X1 U16582 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14967), .ZN(P2_U3269) );
  AND2_X1 U16583 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14967), .ZN(P2_U3270) );
  AND2_X1 U16584 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14967), .ZN(P2_U3271) );
  AND2_X1 U16585 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14967), .ZN(P2_U3272) );
  AND2_X1 U16586 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14967), .ZN(P2_U3273) );
  AND2_X1 U16587 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14967), .ZN(P2_U3274) );
  AND2_X1 U16588 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14967), .ZN(P2_U3275) );
  AND2_X1 U16589 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14967), .ZN(P2_U3276) );
  AND2_X1 U16590 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14967), .ZN(P2_U3277) );
  AND2_X1 U16591 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14967), .ZN(P2_U3278) );
  AND2_X1 U16592 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14967), .ZN(P2_U3279) );
  AND2_X1 U16593 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14967), .ZN(P2_U3280) );
  AND2_X1 U16594 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14967), .ZN(P2_U3281) );
  AND2_X1 U16595 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14967), .ZN(P2_U3282) );
  AND2_X1 U16596 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14967), .ZN(P2_U3283) );
  AND2_X1 U16597 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14967), .ZN(P2_U3284) );
  AND2_X1 U16598 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14967), .ZN(P2_U3285) );
  AND2_X1 U16599 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14967), .ZN(P2_U3286) );
  AND2_X1 U16600 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14967), .ZN(P2_U3287) );
  AND2_X1 U16601 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14967), .ZN(P2_U3288) );
  INV_X1 U16602 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15235) );
  NOR2_X1 U16603 ( .A1(n14966), .A2(n15235), .ZN(P2_U3289) );
  AND2_X1 U16604 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14967), .ZN(P2_U3290) );
  AND2_X1 U16605 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14967), .ZN(P2_U3291) );
  AND2_X1 U16606 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14967), .ZN(P2_U3292) );
  AND2_X1 U16607 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14967), .ZN(P2_U3293) );
  AND2_X1 U16608 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14967), .ZN(P2_U3294) );
  AND2_X1 U16609 ( .A1(n14967), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3295) );
  OAI21_X1 U16610 ( .B1(n14973), .B2(n14969), .A(n14968), .ZN(P2_U3416) );
  AOI22_X1 U16611 ( .A1(n14973), .A2(n14972), .B1(n14971), .B2(n14970), .ZN(
        P2_U3417) );
  AOI211_X1 U16612 ( .C1(n15000), .C2(n14976), .A(n14975), .B(n14974), .ZN(
        n15019) );
  AOI22_X1 U16613 ( .A1(n15018), .A2(n15019), .B1(n7716), .B2(n15017), .ZN(
        P2_U3430) );
  OAI21_X1 U16614 ( .B1(n14978), .B2(n15012), .A(n14977), .ZN(n14980) );
  AOI211_X1 U16615 ( .C1(n15000), .C2(n14981), .A(n14980), .B(n14979), .ZN(
        n15020) );
  INV_X1 U16616 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14982) );
  AOI22_X1 U16617 ( .A1(n15018), .A2(n15020), .B1(n14982), .B2(n15017), .ZN(
        P2_U3436) );
  OR2_X1 U16618 ( .A1(n14983), .A2(n14994), .ZN(n14988) );
  AND2_X1 U16619 ( .A1(n14984), .A2(n14990), .ZN(n14985) );
  NOR2_X1 U16620 ( .A1(n14986), .A2(n14985), .ZN(n14987) );
  AND3_X1 U16621 ( .A1(n14989), .A2(n14988), .A3(n14987), .ZN(n15022) );
  AOI22_X1 U16622 ( .A1(n15018), .A2(n15022), .B1(n7772), .B2(n15017), .ZN(
        P2_U3442) );
  AND2_X1 U16623 ( .A1(n14991), .A2(n14990), .ZN(n14992) );
  NOR2_X1 U16624 ( .A1(n14993), .A2(n14992), .ZN(n14997) );
  OR2_X1 U16625 ( .A1(n14995), .A2(n14994), .ZN(n14996) );
  AOI22_X1 U16626 ( .A1(n15018), .A2(n15023), .B1(n7809), .B2(n15017), .ZN(
        P2_U3448) );
  AND2_X1 U16627 ( .A1(n15001), .A2(n14999), .ZN(n15007) );
  AND2_X1 U16628 ( .A1(n15001), .A2(n15000), .ZN(n15006) );
  OAI21_X1 U16629 ( .B1(n15003), .B2(n15012), .A(n15002), .ZN(n15004) );
  NOR4_X1 U16630 ( .A1(n15007), .A2(n15006), .A3(n15005), .A4(n15004), .ZN(
        n15024) );
  INV_X1 U16631 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15008) );
  AOI22_X1 U16632 ( .A1(n15018), .A2(n15024), .B1(n15008), .B2(n15017), .ZN(
        P2_U3460) );
  AND2_X1 U16633 ( .A1(n15010), .A2(n15009), .ZN(n15016) );
  OAI21_X1 U16634 ( .B1(n15013), .B2(n15012), .A(n15011), .ZN(n15014) );
  NOR3_X1 U16635 ( .A1(n15016), .A2(n15015), .A3(n15014), .ZN(n15026) );
  AOI22_X1 U16636 ( .A1(n15018), .A2(n15026), .B1(n7908), .B2(n15017), .ZN(
        P2_U3463) );
  AOI22_X1 U16637 ( .A1(n15027), .A2(n15019), .B1(n7724), .B2(n15025), .ZN(
        P2_U3499) );
  AOI22_X1 U16638 ( .A1(n15027), .A2(n15020), .B1(n10074), .B2(n15025), .ZN(
        P2_U3501) );
  AOI22_X1 U16639 ( .A1(n15027), .A2(n15022), .B1(n15021), .B2(n15025), .ZN(
        P2_U3503) );
  AOI22_X1 U16640 ( .A1(n15027), .A2(n15023), .B1(n10087), .B2(n15025), .ZN(
        P2_U3505) );
  AOI22_X1 U16641 ( .A1(n15027), .A2(n15024), .B1(n10364), .B2(n15025), .ZN(
        P2_U3509) );
  AOI22_X1 U16642 ( .A1(n15027), .A2(n15026), .B1(n10366), .B2(n15025), .ZN(
        P2_U3510) );
  NOR2_X1 U16643 ( .A1(P3_U3897), .A2(n15028), .ZN(P3_U3150) );
  AOI21_X1 U16644 ( .B1(n15031), .B2(n15030), .A(n15029), .ZN(n15037) );
  XNOR2_X1 U16645 ( .A(n15033), .B(n15032), .ZN(n15034) );
  AOI22_X1 U16646 ( .A1(n15054), .A2(n15035), .B1(n15052), .B2(n15034), .ZN(
        n15036) );
  OAI21_X1 U16647 ( .B1(n15037), .B2(n15056), .A(n15036), .ZN(n15042) );
  AOI21_X1 U16648 ( .B1(n6641), .B2(n15039), .A(n15038), .ZN(n15040) );
  NOR2_X1 U16649 ( .A1(n15040), .A2(n15060), .ZN(n15041) );
  NOR2_X1 U16650 ( .A1(n15042), .A2(n15041), .ZN(n15044) );
  OAI211_X1 U16651 ( .C1(n15045), .C2(n15066), .A(n15044), .B(n15043), .ZN(
        P3_U3190) );
  AOI21_X1 U16652 ( .B1(n15048), .B2(n15047), .A(n15046), .ZN(n15057) );
  XNOR2_X1 U16653 ( .A(n15050), .B(n15049), .ZN(n15051) );
  AOI22_X1 U16654 ( .A1(n15054), .A2(n15053), .B1(n15052), .B2(n15051), .ZN(
        n15055) );
  OAI21_X1 U16655 ( .B1(n15057), .B2(n15056), .A(n15055), .ZN(n15063) );
  AOI21_X1 U16656 ( .B1(n15188), .B2(n15059), .A(n15058), .ZN(n15061) );
  NOR2_X1 U16657 ( .A1(n15061), .A2(n15060), .ZN(n15062) );
  NOR2_X1 U16658 ( .A1(n15063), .A2(n15062), .ZN(n15065) );
  OAI211_X1 U16659 ( .C1(n15067), .C2(n15066), .A(n15065), .B(n15064), .ZN(
        P3_U3191) );
  XNOR2_X1 U16660 ( .A(n15068), .B(n15072), .ZN(n15145) );
  INV_X1 U16661 ( .A(n15069), .ZN(n15070) );
  AOI21_X1 U16662 ( .B1(n15072), .B2(n15071), .A(n15070), .ZN(n15079) );
  AOI22_X1 U16663 ( .A1(n15109), .A2(n15074), .B1(n15073), .B2(n15106), .ZN(
        n15077) );
  NAND2_X1 U16664 ( .A1(n15145), .A2(n15075), .ZN(n15076) );
  OAI211_X1 U16665 ( .C1(n15079), .C2(n15078), .A(n15077), .B(n15076), .ZN(
        n15143) );
  AOI21_X1 U16666 ( .B1(n15102), .B2(n15145), .A(n15143), .ZN(n15086) );
  AND2_X1 U16667 ( .A1(n15081), .A2(n15080), .ZN(n15144) );
  AOI22_X1 U16668 ( .A1(n15083), .A2(n15144), .B1(n15119), .B2(n15082), .ZN(
        n15084) );
  OAI221_X1 U16669 ( .B1(n15124), .B2(n15086), .C1(n15122), .C2(n15085), .A(
        n15084), .ZN(P3_U3228) );
  XNOR2_X1 U16670 ( .A(n15092), .B(n15087), .ZN(n15100) );
  INV_X1 U16671 ( .A(n15100), .ZN(n15131) );
  NOR2_X1 U16672 ( .A1(n15088), .A2(n15169), .ZN(n15130) );
  INV_X1 U16673 ( .A(n15130), .ZN(n15091) );
  OAI22_X1 U16674 ( .A1(n15091), .A2(n15090), .B1(n15089), .B2(n15227), .ZN(
        n15101) );
  XNOR2_X1 U16675 ( .A(n15093), .B(n15092), .ZN(n15098) );
  OAI22_X1 U16676 ( .A1(n15096), .A2(n15095), .B1(n10522), .B2(n15094), .ZN(
        n15097) );
  AOI21_X1 U16677 ( .B1(n15098), .B2(n15112), .A(n15097), .ZN(n15099) );
  OAI21_X1 U16678 ( .B1(n15116), .B2(n15100), .A(n15099), .ZN(n15129) );
  AOI211_X1 U16679 ( .C1(n15102), .C2(n15131), .A(n15101), .B(n15129), .ZN(
        n15103) );
  AOI22_X1 U16680 ( .A1(n15124), .A2(n10248), .B1(n15103), .B2(n15122), .ZN(
        P3_U3231) );
  NOR2_X1 U16681 ( .A1(n15104), .A2(n15169), .ZN(n15126) );
  XNOR2_X1 U16682 ( .A(n15111), .B(n15105), .ZN(n15118) );
  AOI22_X1 U16683 ( .A1(n15109), .A2(n15108), .B1(n15107), .B2(n15106), .ZN(
        n15115) );
  XNOR2_X1 U16684 ( .A(n15110), .B(n15111), .ZN(n15113) );
  NAND2_X1 U16685 ( .A1(n15113), .A2(n15112), .ZN(n15114) );
  OAI211_X1 U16686 ( .C1(n15118), .C2(n15116), .A(n15115), .B(n15114), .ZN(
        n15125) );
  AOI21_X1 U16687 ( .B1(n15126), .B2(n15117), .A(n15125), .ZN(n15123) );
  INV_X1 U16688 ( .A(n15118), .ZN(n15127) );
  AOI22_X1 U16689 ( .A1(n15127), .A2(n15120), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15119), .ZN(n15121) );
  OAI221_X1 U16690 ( .B1(n15124), .B2(n15123), .C1(n15122), .C2(n10226), .A(
        n15121), .ZN(P3_U3232) );
  AOI211_X1 U16691 ( .C1(n15166), .C2(n15127), .A(n15126), .B(n15125), .ZN(
        n15177) );
  INV_X1 U16692 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15128) );
  AOI22_X1 U16693 ( .A1(n15176), .A2(n15177), .B1(n15128), .B2(n15174), .ZN(
        P3_U3393) );
  AOI211_X1 U16694 ( .C1(n15131), .C2(n15166), .A(n15130), .B(n15129), .ZN(
        n15178) );
  INV_X1 U16695 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15132) );
  AOI22_X1 U16696 ( .A1(n15176), .A2(n15178), .B1(n15132), .B2(n15174), .ZN(
        P3_U3396) );
  INV_X1 U16697 ( .A(n15133), .ZN(n15134) );
  AOI211_X1 U16698 ( .C1(n15136), .C2(n15166), .A(n15135), .B(n15134), .ZN(
        n15179) );
  INV_X1 U16699 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15137) );
  AOI22_X1 U16700 ( .A1(n15176), .A2(n15179), .B1(n15137), .B2(n15174), .ZN(
        P3_U3399) );
  INV_X1 U16701 ( .A(n15138), .ZN(n15141) );
  AOI211_X1 U16702 ( .C1(n15141), .C2(n15166), .A(n15140), .B(n15139), .ZN(
        n15180) );
  INV_X1 U16703 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15142) );
  AOI22_X1 U16704 ( .A1(n15176), .A2(n15180), .B1(n15142), .B2(n15174), .ZN(
        P3_U3402) );
  AOI211_X1 U16705 ( .C1(n15145), .C2(n15166), .A(n15144), .B(n15143), .ZN(
        n15182) );
  INV_X1 U16706 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15146) );
  AOI22_X1 U16707 ( .A1(n15176), .A2(n15182), .B1(n15146), .B2(n15174), .ZN(
        P3_U3405) );
  OAI22_X1 U16708 ( .A1(n15149), .A2(n15148), .B1(n15147), .B2(n15169), .ZN(
        n15150) );
  NOR2_X1 U16709 ( .A1(n15151), .A2(n15150), .ZN(n15184) );
  INV_X1 U16710 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15152) );
  AOI22_X1 U16711 ( .A1(n15176), .A2(n15184), .B1(n15152), .B2(n15174), .ZN(
        P3_U3408) );
  AOI211_X1 U16712 ( .C1(n15155), .C2(n15166), .A(n15154), .B(n15153), .ZN(
        n15186) );
  INV_X1 U16713 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15156) );
  AOI22_X1 U16714 ( .A1(n15176), .A2(n15186), .B1(n15156), .B2(n15174), .ZN(
        P3_U3411) );
  INV_X1 U16715 ( .A(n15157), .ZN(n15160) );
  AOI211_X1 U16716 ( .C1(n15160), .C2(n15166), .A(n15159), .B(n15158), .ZN(
        n15187) );
  INV_X1 U16717 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15161) );
  AOI22_X1 U16718 ( .A1(n15176), .A2(n15187), .B1(n15161), .B2(n15174), .ZN(
        P3_U3414) );
  INV_X1 U16719 ( .A(n15162), .ZN(n15165) );
  AOI211_X1 U16720 ( .C1(n15166), .C2(n15165), .A(n15164), .B(n15163), .ZN(
        n15189) );
  INV_X1 U16721 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15167) );
  AOI22_X1 U16722 ( .A1(n15176), .A2(n15189), .B1(n15167), .B2(n15174), .ZN(
        P3_U3417) );
  OAI22_X1 U16723 ( .A1(n15171), .A2(n15170), .B1(n15169), .B2(n15168), .ZN(
        n15172) );
  NOR2_X1 U16724 ( .A1(n15173), .A2(n15172), .ZN(n15192) );
  INV_X1 U16725 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15175) );
  AOI22_X1 U16726 ( .A1(n15176), .A2(n15192), .B1(n15175), .B2(n15174), .ZN(
        P3_U3420) );
  AOI22_X1 U16727 ( .A1(n15193), .A2(n15177), .B1(n10225), .B2(n15190), .ZN(
        P3_U3460) );
  AOI22_X1 U16728 ( .A1(n15193), .A2(n15178), .B1(n10258), .B2(n15190), .ZN(
        P3_U3461) );
  AOI22_X1 U16729 ( .A1(n15193), .A2(n15179), .B1(n10232), .B2(n15190), .ZN(
        P3_U3462) );
  AOI22_X1 U16730 ( .A1(n15193), .A2(n15180), .B1(n10263), .B2(n15190), .ZN(
        P3_U3463) );
  AOI22_X1 U16731 ( .A1(n15193), .A2(n15182), .B1(n15181), .B2(n15190), .ZN(
        P3_U3464) );
  INV_X1 U16732 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15183) );
  AOI22_X1 U16733 ( .A1(n15193), .A2(n15184), .B1(n15183), .B2(n15190), .ZN(
        P3_U3465) );
  AOI22_X1 U16734 ( .A1(n15193), .A2(n15186), .B1(n15185), .B2(n15190), .ZN(
        P3_U3466) );
  INV_X1 U16735 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15209) );
  AOI22_X1 U16736 ( .A1(n15193), .A2(n15187), .B1(n15209), .B2(n15190), .ZN(
        P3_U3467) );
  AOI22_X1 U16737 ( .A1(n15193), .A2(n15189), .B1(n15188), .B2(n15190), .ZN(
        P3_U3468) );
  INV_X1 U16738 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15191) );
  AOI22_X1 U16739 ( .A1(n15193), .A2(n15192), .B1(n15191), .B2(n15190), .ZN(
        P3_U3469) );
  OAI21_X1 U16740 ( .B1(n15196), .B2(n15195), .A(n15194), .ZN(n15207) );
  NAND2_X1 U16741 ( .A1(n15198), .A2(n15197), .ZN(n15202) );
  AOI22_X1 U16742 ( .A1(n15200), .A2(n15199), .B1(P1_U3086), .B2(
        P1_REG3_REG_8__SCAN_IN), .ZN(n15201) );
  OAI211_X1 U16743 ( .C1(n15204), .C2(n15203), .A(n15202), .B(n15201), .ZN(
        n15205) );
  AOI21_X1 U16744 ( .B1(n15207), .B2(n15206), .A(n15205), .ZN(n15392) );
  AOI22_X1 U16745 ( .A1(n15373), .A2(keyinput112), .B1(keyinput72), .B2(n15209), .ZN(n15208) );
  OAI221_X1 U16746 ( .B1(n15373), .B2(keyinput112), .C1(n15209), .C2(
        keyinput72), .A(n15208), .ZN(n15219) );
  XNOR2_X1 U16747 ( .A(n7568), .B(keyinput80), .ZN(n15211) );
  XNOR2_X1 U16748 ( .A(n15345), .B(keyinput67), .ZN(n15210) );
  NOR2_X1 U16749 ( .A1(n15211), .A2(n15210), .ZN(n15215) );
  XNOR2_X1 U16750 ( .A(keyinput96), .B(P3_ADDR_REG_18__SCAN_IN), .ZN(n15214)
         );
  XNOR2_X1 U16751 ( .A(P2_IR_REG_30__SCAN_IN), .B(keyinput126), .ZN(n15213) );
  XNOR2_X1 U16752 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput106), .ZN(n15212)
         );
  NAND4_X1 U16753 ( .A1(n15215), .A2(n15214), .A3(n15213), .A4(n15212), .ZN(
        n15218) );
  XNOR2_X1 U16754 ( .A(n15216), .B(keyinput124), .ZN(n15217) );
  NOR3_X1 U16755 ( .A1(n15219), .A2(n15218), .A3(n15217), .ZN(n15258) );
  AOI22_X1 U16756 ( .A1(P3_REG2_REG_11__SCAN_IN), .A2(keyinput86), .B1(
        P2_REG0_REG_4__SCAN_IN), .B2(keyinput97), .ZN(n15220) );
  OAI221_X1 U16757 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(keyinput86), .C1(
        P2_REG0_REG_4__SCAN_IN), .C2(keyinput97), .A(n15220), .ZN(n15231) );
  AOI22_X1 U16758 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(keyinput98), .B1(
        P3_D_REG_18__SCAN_IN), .B2(keyinput83), .ZN(n15221) );
  OAI221_X1 U16759 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(keyinput98), .C1(
        P3_D_REG_18__SCAN_IN), .C2(keyinput83), .A(n15221), .ZN(n15230) );
  INV_X1 U16760 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n15223) );
  AOI22_X1 U16761 ( .A1(n15224), .A2(keyinput123), .B1(n15223), .B2(keyinput85), .ZN(n15222) );
  OAI221_X1 U16762 ( .B1(n15224), .B2(keyinput123), .C1(n15223), .C2(
        keyinput85), .A(n15222), .ZN(n15229) );
  AOI22_X1 U16763 ( .A1(n15227), .A2(keyinput116), .B1(n15226), .B2(
        keyinput101), .ZN(n15225) );
  OAI221_X1 U16764 ( .B1(n15227), .B2(keyinput116), .C1(n15226), .C2(
        keyinput101), .A(n15225), .ZN(n15228) );
  NOR4_X1 U16765 ( .A1(n15231), .A2(n15230), .A3(n15229), .A4(n15228), .ZN(
        n15257) );
  AOI22_X1 U16766 ( .A1(n8040), .A2(keyinput77), .B1(keyinput122), .B2(n15233), 
        .ZN(n15232) );
  OAI221_X1 U16767 ( .B1(n8040), .B2(keyinput77), .C1(n15233), .C2(keyinput122), .A(n15232), .ZN(n15243) );
  AOI22_X1 U16768 ( .A1(n15235), .A2(keyinput111), .B1(keyinput70), .B2(n15346), .ZN(n15234) );
  OAI221_X1 U16769 ( .B1(n15235), .B2(keyinput111), .C1(n15346), .C2(
        keyinput70), .A(n15234), .ZN(n15242) );
  AOI22_X1 U16770 ( .A1(n8453), .A2(keyinput87), .B1(keyinput65), .B2(n15237), 
        .ZN(n15236) );
  OAI221_X1 U16771 ( .B1(n8453), .B2(keyinput87), .C1(n15237), .C2(keyinput65), 
        .A(n15236), .ZN(n15241) );
  XNOR2_X1 U16772 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput66), .ZN(n15239) );
  XNOR2_X1 U16773 ( .A(P3_REG3_REG_8__SCAN_IN), .B(keyinput90), .ZN(n15238) );
  NAND2_X1 U16774 ( .A1(n15239), .A2(n15238), .ZN(n15240) );
  NOR4_X1 U16775 ( .A1(n15243), .A2(n15242), .A3(n15241), .A4(n15240), .ZN(
        n15256) );
  AOI22_X1 U16776 ( .A1(n15378), .A2(keyinput110), .B1(n15348), .B2(
        keyinput113), .ZN(n15244) );
  OAI221_X1 U16777 ( .B1(n15378), .B2(keyinput110), .C1(n15348), .C2(
        keyinput113), .A(n15244), .ZN(n15254) );
  AOI22_X1 U16778 ( .A1(P1_U3086), .A2(keyinput88), .B1(n15246), .B2(
        keyinput76), .ZN(n15245) );
  OAI221_X1 U16779 ( .B1(P1_U3086), .B2(keyinput88), .C1(n15246), .C2(
        keyinput76), .A(n15245), .ZN(n15253) );
  AOI22_X1 U16780 ( .A1(n15248), .A2(keyinput69), .B1(keyinput89), .B2(n15371), 
        .ZN(n15247) );
  OAI221_X1 U16781 ( .B1(n15248), .B2(keyinput69), .C1(n15371), .C2(keyinput89), .A(n15247), .ZN(n15252) );
  XNOR2_X1 U16782 ( .A(P3_IR_REG_24__SCAN_IN), .B(keyinput71), .ZN(n15250) );
  XNOR2_X1 U16783 ( .A(keyinput99), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n15249) );
  NAND2_X1 U16784 ( .A1(n15250), .A2(n15249), .ZN(n15251) );
  NOR4_X1 U16785 ( .A1(n15254), .A2(n15253), .A3(n15252), .A4(n15251), .ZN(
        n15255) );
  AND4_X1 U16786 ( .A1(n15258), .A2(n15257), .A3(n15256), .A4(n15255), .ZN(
        n15390) );
  OAI22_X1 U16787 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(keyinput74), .B1(keyinput91), .B2(P3_REG1_REG_23__SCAN_IN), .ZN(n15259) );
  AOI221_X1 U16788 ( .B1(P3_IR_REG_5__SCAN_IN), .B2(keyinput74), .C1(
        P3_REG1_REG_23__SCAN_IN), .C2(keyinput91), .A(n15259), .ZN(n15266) );
  OAI22_X1 U16789 ( .A1(P1_REG2_REG_29__SCAN_IN), .A2(keyinput109), .B1(
        keyinput104), .B2(P1_REG3_REG_3__SCAN_IN), .ZN(n15260) );
  AOI221_X1 U16790 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(keyinput109), .C1(
        P1_REG3_REG_3__SCAN_IN), .C2(keyinput104), .A(n15260), .ZN(n15265) );
  OAI22_X1 U16791 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(keyinput115), .B1(
        keyinput82), .B2(P1_REG1_REG_3__SCAN_IN), .ZN(n15261) );
  AOI221_X1 U16792 ( .B1(P1_IR_REG_25__SCAN_IN), .B2(keyinput115), .C1(
        P1_REG1_REG_3__SCAN_IN), .C2(keyinput82), .A(n15261), .ZN(n15264) );
  OAI22_X1 U16793 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(keyinput114), .B1(
        keyinput102), .B2(P3_REG0_REG_17__SCAN_IN), .ZN(n15262) );
  AOI221_X1 U16794 ( .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput114), .C1(
        P3_REG0_REG_17__SCAN_IN), .C2(keyinput102), .A(n15262), .ZN(n15263) );
  NAND4_X1 U16795 ( .A1(n15266), .A2(n15265), .A3(n15264), .A4(n15263), .ZN(
        n15294) );
  OAI22_X1 U16796 ( .A1(P2_D_REG_2__SCAN_IN), .A2(keyinput107), .B1(
        P3_REG2_REG_10__SCAN_IN), .B2(keyinput100), .ZN(n15267) );
  AOI221_X1 U16797 ( .B1(P2_D_REG_2__SCAN_IN), .B2(keyinput107), .C1(
        keyinput100), .C2(P3_REG2_REG_10__SCAN_IN), .A(n15267), .ZN(n15274) );
  OAI22_X1 U16798 ( .A1(P2_REG1_REG_30__SCAN_IN), .A2(keyinput73), .B1(
        P1_REG0_REG_23__SCAN_IN), .B2(keyinput84), .ZN(n15268) );
  AOI221_X1 U16799 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(keyinput73), .C1(
        keyinput84), .C2(P1_REG0_REG_23__SCAN_IN), .A(n15268), .ZN(n15273) );
  OAI22_X1 U16800 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(keyinput105), .B1(
        P3_REG1_REG_18__SCAN_IN), .B2(keyinput103), .ZN(n15269) );
  AOI221_X1 U16801 ( .B1(P1_DATAO_REG_26__SCAN_IN), .B2(keyinput105), .C1(
        keyinput103), .C2(P3_REG1_REG_18__SCAN_IN), .A(n15269), .ZN(n15272) );
  OAI22_X1 U16802 ( .A1(SI_21_), .A2(keyinput78), .B1(keyinput93), .B2(
        P2_REG2_REG_10__SCAN_IN), .ZN(n15270) );
  AOI221_X1 U16803 ( .B1(SI_21_), .B2(keyinput78), .C1(P2_REG2_REG_10__SCAN_IN), .C2(keyinput93), .A(n15270), .ZN(n15271) );
  NAND4_X1 U16804 ( .A1(n15274), .A2(n15273), .A3(n15272), .A4(n15271), .ZN(
        n15293) );
  OAI22_X1 U16805 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(keyinput75), .B1(
        P2_ADDR_REG_10__SCAN_IN), .B2(keyinput117), .ZN(n15275) );
  AOI221_X1 U16806 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(keyinput75), .C1(
        keyinput117), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n15275), .ZN(n15282) );
  OAI22_X1 U16807 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(keyinput127), .B1(
        keyinput64), .B2(P3_ADDR_REG_9__SCAN_IN), .ZN(n15276) );
  AOI221_X1 U16808 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(keyinput127), .C1(
        P3_ADDR_REG_9__SCAN_IN), .C2(keyinput64), .A(n15276), .ZN(n15281) );
  OAI22_X1 U16809 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(keyinput125), .B1(
        keyinput94), .B2(P3_REG0_REG_28__SCAN_IN), .ZN(n15277) );
  AOI221_X1 U16810 ( .B1(P1_DATAO_REG_17__SCAN_IN), .B2(keyinput125), .C1(
        P3_REG0_REG_28__SCAN_IN), .C2(keyinput94), .A(n15277), .ZN(n15280) );
  OAI22_X1 U16811 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(keyinput79), .B1(
        P1_REG0_REG_30__SCAN_IN), .B2(keyinput121), .ZN(n15278) );
  AOI221_X1 U16812 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(keyinput79), .C1(
        keyinput121), .C2(P1_REG0_REG_30__SCAN_IN), .A(n15278), .ZN(n15279) );
  NAND4_X1 U16813 ( .A1(n15282), .A2(n15281), .A3(n15280), .A4(n15279), .ZN(
        n15292) );
  OAI22_X1 U16814 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(keyinput81), .B1(
        keyinput92), .B2(P3_REG3_REG_21__SCAN_IN), .ZN(n15283) );
  AOI221_X1 U16815 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(keyinput81), .C1(
        P3_REG3_REG_21__SCAN_IN), .C2(keyinput92), .A(n15283), .ZN(n15290) );
  OAI22_X1 U16816 ( .A1(SI_15_), .A2(keyinput120), .B1(P1_IR_REG_29__SCAN_IN), 
        .B2(keyinput108), .ZN(n15284) );
  AOI221_X1 U16817 ( .B1(SI_15_), .B2(keyinput120), .C1(keyinput108), .C2(
        P1_IR_REG_29__SCAN_IN), .A(n15284), .ZN(n15289) );
  OAI22_X1 U16818 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(keyinput68), .B1(
        keyinput118), .B2(P1_REG0_REG_19__SCAN_IN), .ZN(n15285) );
  AOI221_X1 U16819 ( .B1(P3_REG3_REG_5__SCAN_IN), .B2(keyinput68), .C1(
        P1_REG0_REG_19__SCAN_IN), .C2(keyinput118), .A(n15285), .ZN(n15288) );
  OAI22_X1 U16820 ( .A1(P2_REG2_REG_1__SCAN_IN), .A2(keyinput119), .B1(
        keyinput95), .B2(P1_IR_REG_23__SCAN_IN), .ZN(n15286) );
  AOI221_X1 U16821 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(keyinput119), .C1(
        P1_IR_REG_23__SCAN_IN), .C2(keyinput95), .A(n15286), .ZN(n15287) );
  NAND4_X1 U16822 ( .A1(n15290), .A2(n15289), .A3(n15288), .A4(n15287), .ZN(
        n15291) );
  NOR4_X1 U16823 ( .A1(n15294), .A2(n15293), .A3(n15292), .A4(n15291), .ZN(
        n15389) );
  AOI22_X1 U16824 ( .A1(P3_D_REG_6__SCAN_IN), .A2(keyinput58), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(keyinput42), .ZN(n15295) );
  OAI221_X1 U16825 ( .B1(P3_D_REG_6__SCAN_IN), .B2(keyinput58), .C1(
        P1_DATAO_REG_5__SCAN_IN), .C2(keyinput42), .A(n15295), .ZN(n15302) );
  AOI22_X1 U16826 ( .A1(P1_REG0_REG_19__SCAN_IN), .A2(keyinput54), .B1(
        P3_REG3_REG_21__SCAN_IN), .B2(keyinput28), .ZN(n15296) );
  OAI221_X1 U16827 ( .B1(P1_REG0_REG_19__SCAN_IN), .B2(keyinput54), .C1(
        P3_REG3_REG_21__SCAN_IN), .C2(keyinput28), .A(n15296), .ZN(n15301) );
  AOI22_X1 U16828 ( .A1(P3_ADDR_REG_9__SCAN_IN), .A2(keyinput0), .B1(
        P3_REG1_REG_23__SCAN_IN), .B2(keyinput27), .ZN(n15297) );
  OAI221_X1 U16829 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(keyinput0), .C1(
        P3_REG1_REG_23__SCAN_IN), .C2(keyinput27), .A(n15297), .ZN(n15300) );
  AOI22_X1 U16830 ( .A1(P3_REG0_REG_28__SCAN_IN), .A2(keyinput30), .B1(
        P2_RD_REG_SCAN_IN), .B2(keyinput16), .ZN(n15298) );
  OAI221_X1 U16831 ( .B1(P3_REG0_REG_28__SCAN_IN), .B2(keyinput30), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput16), .A(n15298), .ZN(n15299) );
  NOR4_X1 U16832 ( .A1(n15302), .A2(n15301), .A3(n15300), .A4(n15299), .ZN(
        n15330) );
  AOI22_X1 U16833 ( .A1(P1_REG0_REG_30__SCAN_IN), .A2(keyinput57), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(keyinput61), .ZN(n15303) );
  OAI221_X1 U16834 ( .B1(P1_REG0_REG_30__SCAN_IN), .B2(keyinput57), .C1(
        P1_DATAO_REG_17__SCAN_IN), .C2(keyinput61), .A(n15303), .ZN(n15310) );
  AOI22_X1 U16835 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(keyinput18), .B1(
        P3_REG1_REG_18__SCAN_IN), .B2(keyinput39), .ZN(n15304) );
  OAI221_X1 U16836 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(keyinput18), .C1(
        P3_REG1_REG_18__SCAN_IN), .C2(keyinput39), .A(n15304), .ZN(n15309) );
  AOI22_X1 U16837 ( .A1(P3_DATAO_REG_11__SCAN_IN), .A2(keyinput60), .B1(
        P2_REG2_REG_10__SCAN_IN), .B2(keyinput29), .ZN(n15305) );
  OAI221_X1 U16838 ( .B1(P3_DATAO_REG_11__SCAN_IN), .B2(keyinput60), .C1(
        P2_REG2_REG_10__SCAN_IN), .C2(keyinput29), .A(n15305), .ZN(n15308) );
  AOI22_X1 U16839 ( .A1(P3_D_REG_4__SCAN_IN), .A2(keyinput12), .B1(
        P2_REG1_REG_6__SCAN_IN), .B2(keyinput17), .ZN(n15306) );
  OAI221_X1 U16840 ( .B1(P3_D_REG_4__SCAN_IN), .B2(keyinput12), .C1(
        P2_REG1_REG_6__SCAN_IN), .C2(keyinput17), .A(n15306), .ZN(n15307) );
  NOR4_X1 U16841 ( .A1(n15310), .A2(n15309), .A3(n15308), .A4(n15307), .ZN(
        n15329) );
  AOI22_X1 U16842 ( .A1(P3_REG0_REG_11__SCAN_IN), .A2(keyinput23), .B1(
        P2_D_REG_2__SCAN_IN), .B2(keyinput43), .ZN(n15311) );
  OAI221_X1 U16843 ( .B1(P3_REG0_REG_11__SCAN_IN), .B2(keyinput23), .C1(
        P2_D_REG_2__SCAN_IN), .C2(keyinput43), .A(n15311), .ZN(n15318) );
  AOI22_X1 U16844 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(keyinput37), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(keyinput41), .ZN(n15312) );
  OAI221_X1 U16845 ( .B1(P2_DATAO_REG_22__SCAN_IN), .B2(keyinput37), .C1(
        P1_DATAO_REG_26__SCAN_IN), .C2(keyinput41), .A(n15312), .ZN(n15317) );
  AOI22_X1 U16846 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(keyinput10), .B1(
        P2_REG2_REG_20__SCAN_IN), .B2(keyinput13), .ZN(n15313) );
  OAI221_X1 U16847 ( .B1(P3_IR_REG_5__SCAN_IN), .B2(keyinput10), .C1(
        P2_REG2_REG_20__SCAN_IN), .C2(keyinput13), .A(n15313), .ZN(n15316) );
  AOI22_X1 U16848 ( .A1(P3_REG2_REG_11__SCAN_IN), .A2(keyinput22), .B1(
        P2_REG1_REG_4__SCAN_IN), .B2(keyinput35), .ZN(n15314) );
  OAI221_X1 U16849 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(keyinput22), .C1(
        P2_REG1_REG_4__SCAN_IN), .C2(keyinput35), .A(n15314), .ZN(n15315) );
  NOR4_X1 U16850 ( .A1(n15318), .A2(n15317), .A3(n15316), .A4(n15315), .ZN(
        n15328) );
  AOI22_X1 U16851 ( .A1(P1_STATE_REG_SCAN_IN), .A2(keyinput24), .B1(
        P2_D_REG_8__SCAN_IN), .B2(keyinput47), .ZN(n15319) );
  OAI221_X1 U16852 ( .B1(P1_STATE_REG_SCAN_IN), .B2(keyinput24), .C1(
        P2_D_REG_8__SCAN_IN), .C2(keyinput47), .A(n15319), .ZN(n15326) );
  AOI22_X1 U16853 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(keyinput11), .B1(
        P2_REG1_REG_8__SCAN_IN), .B2(keyinput15), .ZN(n15320) );
  OAI221_X1 U16854 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(keyinput11), .C1(
        P2_REG1_REG_8__SCAN_IN), .C2(keyinput15), .A(n15320), .ZN(n15325) );
  AOI22_X1 U16855 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(keyinput8), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(keyinput5), .ZN(n15321) );
  OAI221_X1 U16856 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(keyinput8), .C1(
        P2_DATAO_REG_23__SCAN_IN), .C2(keyinput5), .A(n15321), .ZN(n15324) );
  AOI22_X1 U16857 ( .A1(P2_REG0_REG_4__SCAN_IN), .A2(keyinput33), .B1(
        P2_REG2_REG_14__SCAN_IN), .B2(keyinput63), .ZN(n15322) );
  OAI221_X1 U16858 ( .B1(P2_REG0_REG_4__SCAN_IN), .B2(keyinput33), .C1(
        P2_REG2_REG_14__SCAN_IN), .C2(keyinput63), .A(n15322), .ZN(n15323) );
  NOR4_X1 U16859 ( .A1(n15326), .A2(n15325), .A3(n15324), .A4(n15323), .ZN(
        n15327) );
  NAND4_X1 U16860 ( .A1(n15330), .A2(n15329), .A3(n15328), .A4(n15327), .ZN(
        n15388) );
  AOI22_X1 U16861 ( .A1(n11689), .A2(keyinput36), .B1(keyinput53), .B2(n15332), 
        .ZN(n15331) );
  OAI221_X1 U16862 ( .B1(n11689), .B2(keyinput36), .C1(n15332), .C2(keyinput53), .A(n15331), .ZN(n15342) );
  AOI22_X1 U16863 ( .A1(n15335), .A2(keyinput20), .B1(n15334), .B2(keyinput38), 
        .ZN(n15333) );
  OAI221_X1 U16864 ( .B1(n15335), .B2(keyinput20), .C1(n15334), .C2(keyinput38), .A(n15333), .ZN(n15341) );
  XNOR2_X1 U16865 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput31), .ZN(n15339) );
  XNOR2_X1 U16866 ( .A(P3_IR_REG_24__SCAN_IN), .B(keyinput7), .ZN(n15338) );
  XNOR2_X1 U16867 ( .A(P3_REG0_REG_16__SCAN_IN), .B(keyinput1), .ZN(n15337) );
  XNOR2_X1 U16868 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput51), .ZN(n15336) );
  NAND4_X1 U16869 ( .A1(n15339), .A2(n15338), .A3(n15337), .A4(n15336), .ZN(
        n15340) );
  NOR3_X1 U16870 ( .A1(n15342), .A2(n15341), .A3(n15340), .ZN(n15386) );
  AOI22_X1 U16871 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(keyinput44), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(keyinput52), .ZN(n15343) );
  OAI221_X1 U16872 ( .B1(P1_IR_REG_29__SCAN_IN), .B2(keyinput44), .C1(
        P3_REG3_REG_2__SCAN_IN), .C2(keyinput52), .A(n15343), .ZN(n15354) );
  AOI22_X1 U16873 ( .A1(n15346), .A2(keyinput6), .B1(keyinput3), .B2(n15345), 
        .ZN(n15344) );
  OAI221_X1 U16874 ( .B1(n15346), .B2(keyinput6), .C1(n15345), .C2(keyinput3), 
        .A(n15344), .ZN(n15353) );
  AOI22_X1 U16875 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(keyinput26), .B1(
        P3_D_REG_31__SCAN_IN), .B2(keyinput59), .ZN(n15347) );
  OAI221_X1 U16876 ( .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput26), .C1(
        P3_D_REG_31__SCAN_IN), .C2(keyinput59), .A(n15347), .ZN(n15352) );
  XNOR2_X1 U16877 ( .A(n15348), .B(keyinput49), .ZN(n15350) );
  XNOR2_X1 U16878 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput2), .ZN(n15349) );
  NAND2_X1 U16879 ( .A1(n15350), .A2(n15349), .ZN(n15351) );
  NOR4_X1 U16880 ( .A1(n15354), .A2(n15353), .A3(n15352), .A4(n15351), .ZN(
        n15385) );
  AOI22_X1 U16881 ( .A1(n15357), .A2(keyinput40), .B1(keyinput32), .B2(n15356), 
        .ZN(n15355) );
  OAI221_X1 U16882 ( .B1(n15357), .B2(keyinput40), .C1(n15356), .C2(keyinput32), .A(n15355), .ZN(n15369) );
  AOI22_X1 U16883 ( .A1(n15360), .A2(keyinput56), .B1(keyinput19), .B2(n15359), 
        .ZN(n15358) );
  OAI221_X1 U16884 ( .B1(n15360), .B2(keyinput56), .C1(n15359), .C2(keyinput19), .A(n15358), .ZN(n15368) );
  INV_X1 U16885 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n15363) );
  AOI22_X1 U16886 ( .A1(n15363), .A2(keyinput9), .B1(n15362), .B2(keyinput14), 
        .ZN(n15361) );
  OAI221_X1 U16887 ( .B1(n15363), .B2(keyinput9), .C1(n15362), .C2(keyinput14), 
        .A(n15361), .ZN(n15367) );
  XNOR2_X1 U16888 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput21), .ZN(n15365)
         );
  XNOR2_X1 U16889 ( .A(P2_IR_REG_30__SCAN_IN), .B(keyinput62), .ZN(n15364) );
  NAND2_X1 U16890 ( .A1(n15365), .A2(n15364), .ZN(n15366) );
  NOR4_X1 U16891 ( .A1(n15369), .A2(n15368), .A3(n15367), .A4(n15366), .ZN(
        n15384) );
  AOI22_X1 U16892 ( .A1(n15371), .A2(keyinput25), .B1(keyinput45), .B2(n9811), 
        .ZN(n15370) );
  OAI221_X1 U16893 ( .B1(n15371), .B2(keyinput25), .C1(n9811), .C2(keyinput45), 
        .A(n15370), .ZN(n15382) );
  AOI22_X1 U16894 ( .A1(n15374), .A2(keyinput55), .B1(n15373), .B2(keyinput48), 
        .ZN(n15372) );
  OAI221_X1 U16895 ( .B1(n15374), .B2(keyinput55), .C1(n15373), .C2(keyinput48), .A(n15372), .ZN(n15381) );
  AOI22_X1 U16896 ( .A1(n15376), .A2(keyinput50), .B1(keyinput34), .B2(n14278), 
        .ZN(n15375) );
  OAI221_X1 U16897 ( .B1(n15376), .B2(keyinput50), .C1(n14278), .C2(keyinput34), .A(n15375), .ZN(n15380) );
  AOI22_X1 U16898 ( .A1(n8345), .A2(keyinput4), .B1(n15378), .B2(keyinput46), 
        .ZN(n15377) );
  OAI221_X1 U16899 ( .B1(n8345), .B2(keyinput4), .C1(n15378), .C2(keyinput46), 
        .A(n15377), .ZN(n15379) );
  NOR4_X1 U16900 ( .A1(n15382), .A2(n15381), .A3(n15380), .A4(n15379), .ZN(
        n15383) );
  NAND4_X1 U16901 ( .A1(n15386), .A2(n15385), .A3(n15384), .A4(n15383), .ZN(
        n15387) );
  AOI211_X1 U16902 ( .C1(n15390), .C2(n15389), .A(n15388), .B(n15387), .ZN(
        n15391) );
  XNOR2_X1 U16903 ( .A(n15392), .B(n15391), .ZN(P1_U3221) );
  OAI21_X1 U16904 ( .B1(n15395), .B2(n15394), .A(n15393), .ZN(SUB_1596_U59) );
  XOR2_X1 U16905 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15398), .Z(SUB_1596_U53) );
  AOI21_X1 U16906 ( .B1(n15401), .B2(n15400), .A(n15399), .ZN(SUB_1596_U56) );
  AOI21_X1 U16907 ( .B1(n15404), .B2(n15403), .A(n15402), .ZN(n15405) );
  XOR2_X1 U16908 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15405), .Z(SUB_1596_U60) );
  AOI21_X1 U16909 ( .B1(n15408), .B2(n15407), .A(n15406), .ZN(SUB_1596_U5) );
  CLKBUF_X1 U7236 ( .A(n9177), .Z(n6473) );
  CLKBUF_X1 U7240 ( .A(n8181), .Z(n6809) );
  INV_X2 U7291 ( .A(n10243), .ZN(n8601) );
  NAND2_X1 U7297 ( .A1(n7756), .A2(n7755), .ZN(n10953) );
  AND2_X1 U7312 ( .A1(n7096), .A2(n13524), .ZN(n13379) );
  CLKBUF_X1 U7338 ( .A(n9339), .Z(n6853) );
  NAND2_X1 U7471 ( .A1(n13168), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8272) );
  NAND2_X2 U7557 ( .A1(n8096), .A2(n8095), .ZN(n13688) );
  XNOR2_X1 U7701 ( .A(n7714), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7672) );
  INV_X4 U8015 ( .A(n9975), .ZN(n9945) );
  NOR2_X2 U8299 ( .A1(n13633), .A2(n13625), .ZN(n7110) );
  NOR2_X4 U9371 ( .A1(n13688), .A2(n13532), .ZN(n13524) );
  AOI22_X1 U9382 ( .A1(n8016), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8015), .B2(
        n10081), .ZN(n7755) );
  XNOR2_X2 U9421 ( .A(n6670), .B(n7641), .ZN(n8244) );
  AND2_X1 U10032 ( .A1(n10067), .A2(n8244), .ZN(n15413) );
endmodule

