

module b14_C_SARLock_k_64_5 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4742;

  OR2_X1 U2269 ( .A1(n3314), .A2(n2815), .ZN(n2817) );
  NAND2_X1 U2270 ( .A1(n2770), .A2(n2837), .ZN(n2729) );
  AND4_X1 U2271 ( .A1(n2346), .A2(n2345), .A3(n2344), .A4(n2343), .ZN(n2802)
         );
  NAND2_X2 U2273 ( .A1(n2260), .A2(n2261), .ZN(n2360) );
  NOR2_X1 U2274 ( .A1(n2322), .A2(n2323), .ZN(n4518) );
  AOI211_X1 U2275 ( .C1(n3714), .C2(n3713), .A(n3712), .B(n3711), .ZN(n3720)
         );
  INV_X2 U2276 ( .A(n2026), .ZN(n2711) );
  INV_X2 U2277 ( .A(n2731), .ZN(n2718) );
  OR2_X1 U2278 ( .A1(n3909), .A2(n2834), .ZN(n2070) );
  INV_X1 U2279 ( .A(n2729), .ZN(n2714) );
  INV_X1 U2280 ( .A(n2360), .ZN(n2304) );
  INV_X1 U2282 ( .A(IR_REG_31__SCAN_IN), .ZN(n2774) );
  NOR2_X2 U2283 ( .A1(n2508), .A2(n2507), .ZN(n2527) );
  AOI21_X2 U2284 ( .B1(n3984), .B2(n2829), .A(n2828), .ZN(n3973) );
  AOI21_X2 U2285 ( .B1(n2393), .B2(n2392), .A(n2233), .ZN(n3440) );
  AOI21_X2 U2286 ( .B1(n3938), .B2(n2833), .A(n2832), .ZN(n3942) );
  NOR2_X2 U2287 ( .A1(n3973), .A2(n3668), .ZN(n3938) );
  NAND2_X1 U2288 ( .A1(n4733), .A2(n4346), .ZN(n4511) );
  NAND4_X1 U2289 ( .A1(n2335), .A2(n2334), .A3(n2333), .A4(n2332), .ZN(n3745)
         );
  NAND2_X1 U2290 ( .A1(n2294), .A2(n2837), .ZN(n2728) );
  CLKBUF_X2 U2291 ( .A(n2564), .Z(n2709) );
  NAND3_X2 U2292 ( .A1(n2290), .A2(n2289), .A3(n2288), .ZN(n3651) );
  NOR2_X1 U2293 ( .A1(n3430), .A2(n3429), .ZN(n2796) );
  INV_X1 U2294 ( .A(n2069), .ZN(n3876) );
  OAI21_X1 U2295 ( .B1(n3898), .B2(n2165), .A(n2164), .ZN(n2069) );
  NAND2_X1 U2296 ( .A1(n2070), .A2(n2046), .ZN(n3898) );
  OAI21_X1 U2297 ( .B1(n3372), .B2(n2174), .A(n2173), .ZN(n2819) );
  NAND2_X1 U2298 ( .A1(n3918), .A2(n3904), .ZN(n2164) );
  AND2_X1 U2299 ( .A1(n3880), .A2(n4319), .ZN(n2165) );
  CLKBUF_X1 U2300 ( .A(n4523), .Z(n3569) );
  CLKBUF_X1 U2301 ( .A(n3570), .Z(n4525) );
  NAND2_X1 U2302 ( .A1(n4739), .A2(n4346), .ZN(n4440) );
  AND4_X1 U2303 ( .A1(n2400), .A2(n2399), .A3(n2398), .A4(n2397), .ZN(n2812)
         );
  INV_X1 U2304 ( .A(n2802), .ZN(n2806) );
  OR2_X2 U2305 ( .A1(n2728), .A2(n4346), .ZN(n2731) );
  BUF_X1 U2306 ( .A(n2798), .Z(n2799) );
  INV_X1 U2307 ( .A(n3084), .ZN(n3746) );
  NAND4_X1 U2308 ( .A1(n2268), .A2(n2267), .A3(n2266), .A4(n2265), .ZN(n3748)
         );
  AND4_X1 U2309 ( .A1(n2317), .A2(n2316), .A3(n2315), .A4(n2314), .ZN(n3084)
         );
  BUF_X2 U2310 ( .A(n2728), .Z(n2026) );
  OR2_X1 U2311 ( .A1(n2544), .A2(n4528), .ZN(n2562) );
  INV_X1 U2312 ( .A(n2261), .ZN(n2939) );
  AND2_X1 U2313 ( .A1(n2286), .A2(n2253), .ZN(n2777) );
  NAND2_X1 U2314 ( .A1(n2140), .A2(IR_REG_31__SCAN_IN), .ZN(n2286) );
  AND3_X1 U2315 ( .A1(n2035), .A2(n2474), .A3(n2183), .ZN(n2775) );
  AND2_X1 U2316 ( .A1(n2472), .A2(n2139), .ZN(n2138) );
  AND2_X1 U2317 ( .A1(n2225), .A2(n2224), .ZN(n2223) );
  NOR2_X1 U2318 ( .A1(n2248), .A2(IR_REG_14__SCAN_IN), .ZN(n2225) );
  INV_X1 U2319 ( .A(IR_REG_3__SCAN_IN), .ZN(n4239) );
  INV_X1 U2320 ( .A(IR_REG_29__SCAN_IN), .ZN(n2255) );
  NAND2_X1 U2321 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_28__SCAN_IN), .ZN(n2254) );
  INV_X1 U2322 ( .A(n2260), .ZN(n2262) );
  NAND2_X1 U2323 ( .A1(n2806), .A2(n3265), .ZN(n3600) );
  NAND2_X1 U2324 ( .A1(n3593), .A2(n3590), .ZN(n2844) );
  AND2_X1 U2325 ( .A1(n4724), .A2(n2764), .ZN(n2885) );
  AND2_X1 U2326 ( .A1(n2031), .A2(n2244), .ZN(n2139) );
  AND2_X1 U2327 ( .A1(n2250), .A2(n2251), .ZN(n2229) );
  INV_X1 U2328 ( .A(IR_REG_22__SCAN_IN), .ZN(n2251) );
  INV_X1 U2329 ( .A(IR_REG_21__SCAN_IN), .ZN(n2250) );
  INV_X1 U2330 ( .A(IR_REG_20__SCAN_IN), .ZN(n4247) );
  INV_X1 U2331 ( .A(n2454), .ZN(n2201) );
  XNOR2_X1 U2332 ( .A(n3236), .B(n2084), .ZN(n4592) );
  AND2_X1 U2333 ( .A1(n4639), .A2(n2102), .ZN(n2101) );
  INV_X1 U2334 ( .A(n3786), .ZN(n2102) );
  OAI21_X1 U2335 ( .B1(n3857), .B2(n2168), .A(n2166), .ZN(n2899) );
  AOI21_X1 U2336 ( .B1(n2169), .B2(n2167), .A(n2052), .ZN(n2166) );
  INV_X1 U2337 ( .A(n2169), .ZN(n2168) );
  INV_X1 U2338 ( .A(n3679), .ZN(n2167) );
  INV_X1 U2339 ( .A(n2071), .ZN(n4005) );
  OAI211_X1 U2340 ( .C1(n2161), .C2(n2160), .A(n2072), .B(n2051), .ZN(n2071)
         );
  INV_X1 U2341 ( .A(n2826), .ZN(n2160) );
  AOI21_X1 U2342 ( .B1(n2178), .B2(n2176), .A(n2048), .ZN(n2175) );
  INV_X1 U2343 ( .A(n2037), .ZN(n2176) );
  AND2_X1 U2344 ( .A1(n4105), .A2(n4107), .ZN(n4410) );
  NAND2_X1 U2345 ( .A1(n3600), .A2(n3596), .ZN(n2804) );
  AND4_X1 U2346 ( .A1(n2365), .A2(n2364), .A3(n2363), .A4(n2362), .ZN(n3276)
         );
  OR2_X1 U2347 ( .A1(n3745), .A2(n3475), .ZN(n2803) );
  AND2_X1 U2348 ( .A1(n2727), .A2(n2726), .ZN(n4305) );
  OR2_X1 U2349 ( .A1(n3829), .A2(n2564), .ZN(n2727) );
  AND2_X1 U2350 ( .A1(n3065), .A2(n2778), .ZN(n4346) );
  NAND2_X1 U2351 ( .A1(n2928), .A2(IR_REG_31__SCAN_IN), .ZN(n2142) );
  INV_X1 U2352 ( .A(n4305), .ZN(n3848) );
  AND2_X1 U2353 ( .A1(n4410), .A2(n2066), .ZN(n2144) );
  AOI21_X1 U2354 ( .B1(n2116), .B2(n2879), .A(n2114), .ZN(n2113) );
  INV_X1 U2355 ( .A(n3650), .ZN(n2114) );
  INV_X1 U2356 ( .A(n2113), .ZN(n2111) );
  INV_X1 U2357 ( .A(n2175), .ZN(n2174) );
  AND2_X1 U2358 ( .A1(n3462), .A2(n3463), .ZN(n3461) );
  AND2_X1 U2359 ( .A1(n2526), .A2(n2525), .ZN(n2540) );
  OR2_X1 U2360 ( .A1(n3455), .A2(n3451), .ZN(n2526) );
  INV_X1 U2361 ( .A(n2984), .ZN(n2096) );
  NOR2_X1 U2362 ( .A1(n3664), .A2(n2124), .ZN(n2123) );
  NAND2_X1 U2363 ( .A1(n3894), .A2(n3709), .ZN(n2125) );
  INV_X1 U2364 ( .A(n4118), .ZN(n2163) );
  NAND2_X1 U2365 ( .A1(n4055), .A2(n4044), .ZN(n2820) );
  OR2_X1 U2366 ( .A1(n3627), .A2(n4088), .ZN(n2120) );
  NAND2_X1 U2367 ( .A1(n4411), .A2(n3624), .ZN(n2859) );
  NAND2_X1 U2368 ( .A1(n2146), .A2(n2032), .ZN(n2151) );
  OR2_X1 U2369 ( .A1(n2153), .A2(n2028), .ZN(n2146) );
  NOR2_X1 U2370 ( .A1(n2111), .A2(n2902), .ZN(n2109) );
  OAI22_X1 U2371 ( .A1(n2112), .A2(n2111), .B1(n2902), .B2(n2113), .ZN(n2110)
         );
  NOR2_X1 U2372 ( .A1(n2116), .A2(n2902), .ZN(n2112) );
  NAND2_X1 U2373 ( .A1(n2889), .A2(n4016), .ZN(n2080) );
  OR2_X1 U2374 ( .A1(n4542), .A2(n2709), .ZN(n2550) );
  INV_X1 U2375 ( .A(n3258), .ZN(n3265) );
  INV_X1 U2376 ( .A(IR_REG_17__SCAN_IN), .ZN(n2224) );
  INV_X1 U2377 ( .A(IR_REG_23__SCAN_IN), .ZN(n4246) );
  OR3_X1 U2378 ( .A1(n2430), .A2(IR_REG_8__SCAN_IN), .A3(IR_REG_7__SCAN_IN), 
        .ZN(n2443) );
  OR3_X1 U2379 ( .A1(n3414), .A2(n2501), .A3(n2500), .ZN(n2521) );
  INV_X1 U2380 ( .A(n2216), .ZN(n2211) );
  OR2_X1 U2381 ( .A1(n2450), .A2(n2201), .ZN(n2200) );
  OR2_X1 U2382 ( .A1(n2055), .A2(n2191), .ZN(n2190) );
  INV_X1 U2383 ( .A(n3302), .ZN(n2191) );
  NAND2_X1 U2384 ( .A1(n2451), .A2(n2453), .ZN(n2454) );
  INV_X1 U2385 ( .A(n2195), .ZN(n2194) );
  OAI21_X1 U2386 ( .B1(n2354), .B2(n2196), .A(n3118), .ZN(n2195) );
  INV_X1 U2387 ( .A(n2358), .ZN(n2196) );
  INV_X1 U2388 ( .A(n2207), .ZN(n2206) );
  OAI21_X1 U2389 ( .B1(n2209), .B2(n2208), .A(n3497), .ZN(n2207) );
  INV_X1 U2390 ( .A(n2038), .ZN(n2208) );
  OR2_X1 U2391 ( .A1(n2773), .A2(n2946), .ZN(n2780) );
  OR2_X1 U2392 ( .A1(n2704), .A2(n2719), .ZN(n3431) );
  NAND2_X1 U2393 ( .A1(n2278), .A2(n2277), .ZN(n2294) );
  AND2_X1 U2394 ( .A1(n2934), .A2(n2931), .ZN(n2278) );
  INV_X1 U2395 ( .A(n2734), .ZN(n2277) );
  NAND2_X1 U2396 ( .A1(n2097), .A2(n2098), .ZN(n3032) );
  OAI21_X1 U2397 ( .B1(n2322), .B2(n2323), .A(REG1_REG_2__SCAN_IN), .ZN(n2097)
         );
  INV_X1 U2398 ( .A(n2323), .ZN(n2099) );
  OAI21_X1 U2399 ( .B1(n2991), .B2(n3770), .A(n3773), .ZN(n3005) );
  XNOR2_X1 U2400 ( .A(n3212), .B(n4712), .ZN(n4549) );
  NAND2_X1 U2401 ( .A1(n4549), .A2(REG1_REG_8__SCAN_IN), .ZN(n4548) );
  NAND2_X1 U2402 ( .A1(n4560), .A2(n3232), .ZN(n3233) );
  NAND2_X1 U2403 ( .A1(n4596), .A2(n3218), .ZN(n3220) );
  NAND2_X1 U2404 ( .A1(n3220), .A2(n3219), .ZN(n3326) );
  NAND2_X1 U2405 ( .A1(n4581), .A2(n3235), .ZN(n3236) );
  NAND2_X1 U2406 ( .A1(n4592), .A2(REG2_REG_12__SCAN_IN), .ZN(n4590) );
  OR2_X1 U2407 ( .A1(n3343), .A2(n3342), .ZN(n3793) );
  AND2_X1 U2408 ( .A1(n3793), .A2(n3792), .ZN(n3795) );
  OR2_X1 U2409 ( .A1(n2672), .A2(n3501), .ZN(n2683) );
  OR2_X1 U2410 ( .A1(n2286), .A2(IR_REG_27__SCAN_IN), .ZN(n2290) );
  NAND2_X1 U2411 ( .A1(n2286), .A2(IR_REG_28__SCAN_IN), .ZN(n2289) );
  AND4_X1 U2412 ( .A1(n2627), .A2(n2626), .A3(n2625), .A4(n2624), .ZN(n3935)
         );
  NAND2_X1 U2413 ( .A1(n2030), .A2(n2049), .ZN(n2161) );
  OAI21_X1 U2414 ( .B1(n3312), .B2(n2135), .A(n2132), .ZN(n4411) );
  AOI21_X1 U2415 ( .B1(n2136), .B2(n2134), .A(n2133), .ZN(n2132) );
  INV_X1 U2416 ( .A(n2136), .ZN(n2135) );
  INV_X1 U2417 ( .A(n3621), .ZN(n2133) );
  INV_X1 U2418 ( .A(n3372), .ZN(n2181) );
  INV_X1 U2419 ( .A(n4410), .ZN(n2179) );
  OR2_X1 U2420 ( .A1(n3318), .A2(n4427), .ZN(n2182) );
  OAI21_X1 U2421 ( .B1(n3289), .B2(n2849), .A(n3612), .ZN(n3360) );
  NOR2_X1 U2422 ( .A1(n3743), .A2(n3274), .ZN(n2155) );
  NAND2_X1 U2423 ( .A1(n2157), .A2(n2028), .ZN(n2156) );
  INV_X1 U2424 ( .A(n3272), .ZN(n2157) );
  OAI21_X1 U2425 ( .B1(n3172), .B2(n3171), .A(n3613), .ZN(n3273) );
  INV_X1 U2426 ( .A(n2804), .ZN(n2145) );
  AND2_X1 U2427 ( .A1(n2804), .A2(n3251), .ZN(n2805) );
  NAND2_X1 U2428 ( .A1(n2804), .A2(n2143), .ZN(n3254) );
  INV_X1 U2429 ( .A(n3252), .ZN(n2143) );
  NAND2_X1 U2430 ( .A1(n2838), .A2(n3802), .ZN(n4419) );
  NAND2_X1 U2431 ( .A1(n2881), .A2(n2880), .ZN(n4421) );
  INV_X1 U2432 ( .A(n3736), .ZN(n2763) );
  NAND2_X1 U2433 ( .A1(n3846), .A2(n3833), .ZN(n2910) );
  NOR2_X1 U2434 ( .A1(n3884), .A2(n2076), .ZN(n3846) );
  OR2_X1 U2435 ( .A1(n2027), .A2(n3945), .ZN(n3947) );
  NAND2_X1 U2436 ( .A1(n3266), .A2(n3265), .ZN(n3264) );
  NAND2_X1 U2437 ( .A1(n4246), .A2(n2275), .ZN(n2270) );
  OR2_X1 U2438 ( .A1(n2269), .A2(n2774), .ZN(n2751) );
  NAND2_X1 U2439 ( .A1(n2294), .A2(n4695), .ZN(n2946) );
  NAND2_X1 U2440 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2253) );
  AND2_X1 U2441 ( .A1(n4241), .A2(n4247), .ZN(n2031) );
  AND2_X1 U2442 ( .A1(n2252), .A2(n2229), .ZN(n2228) );
  NOR2_X1 U2443 ( .A1(n2270), .A2(IR_REG_25__SCAN_IN), .ZN(n2252) );
  INV_X1 U2444 ( .A(IR_REG_24__SCAN_IN), .ZN(n2275) );
  NAND2_X1 U2445 ( .A1(n2751), .A2(n4246), .ZN(n2750) );
  OAI21_X1 U2446 ( .B1(n2751), .B2(n4246), .A(n2750), .ZN(n2944) );
  NAND2_X1 U2447 ( .A1(n2282), .A2(n2036), .ZN(n2764) );
  XNOR2_X1 U2448 ( .A(n2285), .B(n4247), .ZN(n2778) );
  NAND2_X1 U2449 ( .A1(n2284), .A2(IR_REG_31__SCAN_IN), .ZN(n2285) );
  INV_X1 U2450 ( .A(IR_REG_19__SCAN_IN), .ZN(n4241) );
  NAND2_X1 U2451 ( .A1(n2702), .A2(n3564), .ZN(n3430) );
  OR2_X1 U2452 ( .A1(n3349), .A2(n3350), .ZN(n3386) );
  NAND2_X1 U2453 ( .A1(n3471), .A2(n3472), .ZN(n3470) );
  AOI21_X1 U2454 ( .B1(n2221), .B2(n2219), .A(n2063), .ZN(n2218) );
  INV_X1 U2455 ( .A(n2221), .ZN(n2220) );
  INV_X1 U2456 ( .A(n3530), .ZN(n2219) );
  INV_X1 U2457 ( .A(n4543), .ZN(n3574) );
  INV_X1 U2458 ( .A(n3802), .ZN(n3732) );
  NAND2_X1 U2459 ( .A1(n2690), .A2(n2689), .ZN(n4303) );
  INV_X1 U2460 ( .A(n4323), .ZN(n3900) );
  XNOR2_X1 U2461 ( .A(n3233), .B(n2083), .ZN(n4572) );
  NAND2_X1 U2462 ( .A1(n4572), .A2(REG2_REG_10__SCAN_IN), .ZN(n4571) );
  XNOR2_X1 U2463 ( .A(n3795), .B(n3794), .ZN(n4612) );
  NAND2_X1 U2464 ( .A1(n4612), .A2(n4610), .ZN(n4611) );
  NAND2_X1 U2465 ( .A1(n4619), .A2(n4621), .ZN(n4620) );
  NAND2_X1 U2466 ( .A1(n4632), .A2(n4633), .ZN(n2089) );
  NOR2_X1 U2467 ( .A1(n4626), .A2(n3786), .ZN(n4638) );
  NAND2_X1 U2468 ( .A1(n3760), .A2(n3797), .ZN(n2085) );
  AOI21_X1 U2469 ( .B1(n4635), .B2(ADDR_REG_18__SCAN_IN), .A(n4634), .ZN(n2086) );
  NOR2_X1 U2470 ( .A1(n4632), .A2(n4633), .ZN(n4631) );
  XNOR2_X1 U2471 ( .A(n2899), .B(n3693), .ZN(n3839) );
  XNOR2_X1 U2472 ( .A(n3257), .B(n2804), .ZN(n3263) );
  NAND2_X1 U2473 ( .A1(n3818), .A2(n2129), .ZN(n2128) );
  AOI21_X1 U2474 ( .B1(n3813), .B2(n4726), .A(n2130), .ZN(n2129) );
  OAI21_X1 U2475 ( .B1(n3657), .B2(n4428), .A(n2908), .ZN(n2130) );
  INV_X1 U2476 ( .A(n2128), .ZN(n2913) );
  INV_X1 U2477 ( .A(n3977), .ZN(n2889) );
  AND2_X1 U2478 ( .A1(n2144), .A2(n3685), .ZN(n3689) );
  OAI21_X1 U2479 ( .B1(n4186), .B2(n4710), .A(n4557), .ZN(n3214) );
  NOR2_X1 U2480 ( .A1(n2836), .A2(n2170), .ZN(n2169) );
  INV_X1 U2481 ( .A(n3680), .ZN(n2170) );
  NOR2_X1 U2482 ( .A1(n2703), .A2(n3432), .ZN(n2719) );
  INV_X1 U2483 ( .A(n2123), .ZN(n2122) );
  OR2_X1 U2484 ( .A1(n2122), .A2(n3709), .ZN(n2121) );
  AND2_X1 U2485 ( .A1(n2234), .A2(n2230), .ZN(n2131) );
  INV_X1 U2486 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2561) );
  INV_X1 U2487 ( .A(IR_REG_10__SCAN_IN), .ZN(n4240) );
  OR2_X1 U2488 ( .A1(n2486), .A2(n2466), .ZN(n2508) );
  INV_X1 U2489 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2483) );
  OR2_X1 U2490 ( .A1(n2484), .A2(n2483), .ZN(n2486) );
  INV_X1 U2491 ( .A(n3623), .ZN(n2137) );
  INV_X1 U2492 ( .A(n3606), .ZN(n2134) );
  INV_X1 U2493 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2423) );
  NOR2_X1 U2494 ( .A1(n2424), .A2(n2423), .ZN(n2437) );
  AND2_X1 U2495 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2361) );
  NAND2_X1 U2496 ( .A1(n3727), .A2(n2778), .ZN(n2837) );
  NAND2_X1 U2497 ( .A1(n3852), .A2(n3869), .ZN(n2076) );
  NAND2_X1 U2498 ( .A1(n2865), .A2(n2230), .ZN(n3986) );
  OR3_X1 U2499 ( .A1(n4381), .A2(n3676), .A3(n4372), .ZN(n2074) );
  AND2_X1 U2500 ( .A1(n2162), .A2(n2039), .ZN(n4084) );
  NAND2_X1 U2501 ( .A1(n2158), .A2(n2232), .ZN(n2162) );
  AOI21_X1 U2502 ( .B1(n2175), .B2(n2177), .A(n2042), .ZN(n2173) );
  AND2_X1 U2503 ( .A1(n2059), .A2(n2851), .ZN(n2082) );
  OR2_X1 U2504 ( .A1(n3264), .A2(n3242), .ZN(n3177) );
  NAND2_X1 U2505 ( .A1(n2141), .A2(REG0_REG_4__SCAN_IN), .ZN(n2344) );
  OR2_X1 U2506 ( .A1(n2946), .A2(n2884), .ZN(n3055) );
  AND2_X1 U2507 ( .A1(n2474), .A2(n2223), .ZN(n2584) );
  INV_X1 U2508 ( .A(IR_REG_6__SCAN_IN), .ZN(n2401) );
  CLKBUF_X1 U2509 ( .A(n2320), .Z(n2321) );
  INV_X1 U2510 ( .A(n3422), .ZN(n2214) );
  OR2_X1 U2511 ( .A1(n2664), .A2(n2671), .ZN(n2209) );
  INV_X1 U2512 ( .A(n3745), .ZN(n3193) );
  NAND2_X1 U2513 ( .A1(n3529), .A2(n3530), .ZN(n3528) );
  NOR2_X1 U2514 ( .A1(n2631), .A2(n2222), .ZN(n2221) );
  INV_X1 U2515 ( .A(n3532), .ZN(n2222) );
  NAND2_X1 U2516 ( .A1(n3386), .A2(n2450), .ZN(n3383) );
  INV_X1 U2517 ( .A(n3099), .ZN(n2328) );
  NOR2_X1 U2518 ( .A1(n2574), .A2(n2217), .ZN(n2216) );
  NAND2_X1 U2519 ( .A1(n2543), .A2(n2542), .ZN(n4533) );
  OR2_X1 U2520 ( .A1(n2773), .A2(n3734), .ZN(n2787) );
  AND3_X1 U2521 ( .A1(n3655), .A2(n3654), .A3(n3653), .ZN(n3722) );
  NAND2_X1 U2522 ( .A1(n3032), .A2(n2096), .ZN(n2095) );
  NAND2_X1 U2523 ( .A1(n3004), .A2(n2107), .ZN(n2106) );
  OR2_X1 U2524 ( .A1(n3227), .A2(n2090), .ZN(n3230) );
  NOR2_X1 U2525 ( .A1(n3228), .A2(n3295), .ZN(n2090) );
  NAND2_X1 U2526 ( .A1(n4548), .A2(n3213), .ZN(n4558) );
  NAND2_X1 U2527 ( .A1(n4558), .A2(n4559), .ZN(n4557) );
  XOR2_X1 U2528 ( .A(n3214), .B(n4568), .Z(n4570) );
  NAND2_X1 U2529 ( .A1(n3326), .A2(n3327), .ZN(n3329) );
  NAND2_X1 U2530 ( .A1(n3782), .A2(n3783), .ZN(n3784) );
  NAND2_X1 U2531 ( .A1(n2100), .A2(n2104), .ZN(n2103) );
  INV_X1 U2532 ( .A(n4624), .ZN(n2104) );
  NAND2_X1 U2533 ( .A1(n2125), .A2(n2123), .ZN(n3859) );
  NAND2_X1 U2534 ( .A1(n2125), .A2(n3667), .ZN(n3878) );
  AND2_X1 U2535 ( .A1(n3667), .A2(n3666), .ZN(n3897) );
  AND2_X1 U2536 ( .A1(n3913), .A2(n3912), .ZN(n3931) );
  AND2_X1 U2537 ( .A1(n3669), .A2(n3936), .ZN(n3972) );
  AND4_X1 U2538 ( .A1(n2583), .A2(n2582), .A3(n2581), .A4(n2580), .ZN(n3997)
         );
  NOR2_X1 U2539 ( .A1(n2562), .A2(n2561), .ZN(n2578) );
  INV_X1 U2540 ( .A(n2820), .ZN(n2823) );
  INV_X1 U2541 ( .A(n4055), .ZN(n4046) );
  NAND2_X1 U2542 ( .A1(n3701), .A2(n3699), .ZN(n4055) );
  AOI21_X1 U2543 ( .B1(n2040), .B2(n4088), .A(n2119), .ZN(n2118) );
  INV_X1 U2544 ( .A(n3609), .ZN(n2119) );
  AND4_X1 U2545 ( .A1(n2568), .A2(n2567), .A3(n2566), .A4(n2565), .ZN(n4059)
         );
  NAND2_X1 U2546 ( .A1(n4085), .A2(n2860), .ZN(n4086) );
  NAND2_X1 U2547 ( .A1(n2859), .A2(n3627), .ZN(n4085) );
  AND2_X1 U2548 ( .A1(n2437), .A2(REG3_REG_10__SCAN_IN), .ZN(n2455) );
  NAND2_X1 U2549 ( .A1(n3360), .A2(n3605), .ZN(n2850) );
  NAND2_X1 U2550 ( .A1(n2395), .A2(REG3_REG_7__SCAN_IN), .ZN(n2408) );
  OR2_X1 U2551 ( .A1(n2408), .A2(n3306), .ZN(n2424) );
  NAND2_X1 U2552 ( .A1(n2148), .A2(n2152), .ZN(n3359) );
  NAND2_X1 U2553 ( .A1(n3272), .A2(n2149), .ZN(n2148) );
  INV_X1 U2554 ( .A(n3442), .ZN(n3293) );
  NAND2_X1 U2555 ( .A1(n2847), .A2(n3601), .ZN(n3289) );
  OAI21_X1 U2556 ( .B1(n3257), .B2(n2845), .A(n3600), .ZN(n3172) );
  AND2_X1 U2557 ( .A1(n2807), .A2(n3254), .ZN(n2808) );
  NAND2_X1 U2558 ( .A1(n3146), .A2(n3595), .ZN(n3257) );
  INV_X1 U2559 ( .A(n4421), .ZN(n4115) );
  INV_X1 U2560 ( .A(n2844), .ZN(n3684) );
  NAND4_X1 U2561 ( .A1(n2309), .A2(n2308), .A3(n2307), .A4(n2306), .ZN(n2798)
         );
  OR2_X1 U2562 ( .A1(n2564), .A2(n3124), .ZN(n2307) );
  OR2_X1 U2563 ( .A1(n3652), .A2(n2305), .ZN(n2308) );
  INV_X1 U2564 ( .A(n3152), .ZN(n3137) );
  OR2_X1 U2565 ( .A1(n2842), .A2(n3078), .ZN(n3079) );
  AOI22_X1 U2566 ( .A1(n2907), .A2(n4421), .B1(n3808), .B2(n3741), .ZN(n3818)
         );
  NOR2_X1 U2567 ( .A1(n2029), .A2(n4296), .ZN(n4295) );
  NOR2_X1 U2568 ( .A1(n3884), .A2(n3863), .ZN(n3867) );
  INV_X1 U2569 ( .A(n3879), .ZN(n3885) );
  OR2_X1 U2570 ( .A1(n3899), .A2(n3879), .ZN(n3884) );
  AND3_X1 U2571 ( .A1(n2676), .A2(n2675), .A3(n2674), .ZN(n4323) );
  INV_X1 U2572 ( .A(n3917), .ZN(n3922) );
  NOR2_X1 U2573 ( .A1(n3947), .A2(n3922), .ZN(n3923) );
  NAND2_X1 U2574 ( .A1(n2079), .A2(n3998), .ZN(n2078) );
  NOR2_X1 U2575 ( .A1(n2080), .A2(n4336), .ZN(n2079) );
  NOR2_X1 U2576 ( .A1(n4029), .A2(n4009), .ZN(n4014) );
  OR2_X1 U2577 ( .A1(n4052), .A2(n4359), .ZN(n4029) );
  AND4_X1 U2578 ( .A1(n2551), .A2(n2550), .A3(n2549), .A4(n2548), .ZN(n4363)
         );
  NOR2_X1 U2579 ( .A1(n4275), .A2(n2074), .ZN(n4071) );
  AND4_X1 U2580 ( .A1(n2513), .A2(n2512), .A3(n2511), .A4(n2510), .ZN(n4376)
         );
  NOR3_X1 U2581 ( .A1(n4275), .A2(n4381), .A3(n3676), .ZN(n4091) );
  INV_X1 U2582 ( .A(n4413), .ZN(n4407) );
  NOR2_X1 U2583 ( .A1(n4404), .A2(n4413), .ZN(n4405) );
  NAND2_X1 U2584 ( .A1(n4720), .A2(n2081), .ZN(n4404) );
  AND2_X1 U2585 ( .A1(n2082), .A2(n4427), .ZN(n2081) );
  AND4_X1 U2586 ( .A1(n2460), .A2(n2459), .A3(n2458), .A4(n2457), .ZN(n4430)
         );
  NAND2_X1 U2587 ( .A1(n4720), .A2(n2082), .ZN(n3375) );
  AND4_X1 U2588 ( .A1(n2415), .A2(n2414), .A3(n2413), .A4(n2412), .ZN(n3398)
         );
  NAND2_X1 U2589 ( .A1(n4720), .A2(n2059), .ZN(n3356) );
  AND2_X1 U2590 ( .A1(n4720), .A2(n3293), .ZN(n3358) );
  NOR2_X1 U2591 ( .A1(n3177), .A2(n3274), .ZN(n4720) );
  NOR2_X1 U2592 ( .A1(n3153), .A2(n2045), .ZN(n3266) );
  INV_X1 U2593 ( .A(n3475), .ZN(n3200) );
  NAND2_X1 U2594 ( .A1(n4419), .A2(n4350), .ZN(n4726) );
  INV_X1 U2595 ( .A(n4428), .ZN(n4412) );
  INV_X1 U2596 ( .A(n4434), .ZN(n4397) );
  INV_X1 U2597 ( .A(n3126), .ZN(n3083) );
  NAND2_X1 U2598 ( .A1(n3065), .A2(n4514), .ZN(n4428) );
  AND2_X1 U2599 ( .A1(n2763), .A2(n2762), .ZN(n4724) );
  AND2_X1 U2600 ( .A1(n2228), .A2(n2184), .ZN(n2183) );
  AND2_X1 U2601 ( .A1(n2031), .A2(n2057), .ZN(n2184) );
  AND2_X1 U2602 ( .A1(n2228), .A2(n2227), .ZN(n2226) );
  INV_X1 U2603 ( .A(IR_REG_26__SCAN_IN), .ZN(n2227) );
  NAND2_X1 U2604 ( .A1(n2247), .A2(n2246), .ZN(n2248) );
  INV_X1 U2605 ( .A(IR_REG_16__SCAN_IN), .ZN(n2246) );
  INV_X1 U2606 ( .A(IR_REG_4__SCAN_IN), .ZN(n2237) );
  OAI21_X1 U2607 ( .B1(n2319), .B2(n2093), .A(n2091), .ZN(n2323) );
  NAND2_X1 U2608 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2093)
         );
  NAND2_X1 U2609 ( .A1(n2774), .A2(n2092), .ZN(n2091) );
  NAND2_X1 U2610 ( .A1(n3440), .A2(n3439), .ZN(n3438) );
  INV_X1 U2611 ( .A(n4527), .ZN(n3572) );
  OAI21_X1 U2612 ( .B1(n2560), .B2(n2212), .A(n2210), .ZN(n3480) );
  INV_X1 U2613 ( .A(n2213), .ZN(n2212) );
  AOI21_X1 U2614 ( .B1(n2213), .B2(n2211), .A(n2065), .ZN(n2210) );
  AND2_X1 U2615 ( .A1(n2577), .A2(n2214), .ZN(n2213) );
  NAND2_X1 U2616 ( .A1(n3438), .A2(n2407), .ZN(n3305) );
  NAND2_X1 U2617 ( .A1(n3528), .A2(n3532), .ZN(n3490) );
  AOI21_X1 U2618 ( .B1(n2041), .B2(n2201), .A(n2199), .ZN(n2198) );
  INV_X1 U2619 ( .A(n3406), .ZN(n2199) );
  NAND2_X1 U2620 ( .A1(n2205), .A2(n2038), .ZN(n3499) );
  NAND2_X1 U2621 ( .A1(n3554), .A2(n2209), .ZN(n2205) );
  NAND2_X1 U2622 ( .A1(n3188), .A2(n2358), .ZN(n3119) );
  INV_X1 U2623 ( .A(n2846), .ZN(n3242) );
  AOI21_X1 U2624 ( .B1(n3554), .B2(n2664), .A(n2236), .ZN(n3515) );
  NAND2_X1 U2625 ( .A1(n3470), .A2(n2354), .ZN(n3188) );
  NOR2_X1 U2626 ( .A1(n2780), .A2(n2754), .ZN(n4538) );
  AND2_X1 U2627 ( .A1(n2190), .A2(n2188), .ZN(n2187) );
  OR2_X1 U2628 ( .A1(n2407), .A2(n2189), .ZN(n2188) );
  NAND2_X1 U2629 ( .A1(n2293), .A2(n2292), .ZN(n3093) );
  NAND2_X1 U2630 ( .A1(n3383), .A2(n2454), .ZN(n3408) );
  NAND2_X1 U2631 ( .A1(n2215), .A2(n2577), .ZN(n3424) );
  NAND2_X1 U2632 ( .A1(n2560), .A2(n2216), .ZN(n2215) );
  AOI21_X1 U2633 ( .B1(n2194), .B2(n2196), .A(n2047), .ZN(n2193) );
  NAND2_X1 U2634 ( .A1(n2204), .A2(n2202), .ZN(n3568) );
  AOI21_X1 U2635 ( .B1(n2206), .B2(n2208), .A(n2203), .ZN(n2202) );
  INV_X1 U2636 ( .A(n3498), .ZN(n2203) );
  NOR2_X1 U2637 ( .A1(n2787), .A2(n3020), .ZN(n3570) );
  OAI21_X1 U2638 ( .B1(n2780), .B2(n4428), .A(n4647), .ZN(n4523) );
  NOR2_X2 U2639 ( .A1(n2787), .A2(n4521), .ZN(n4527) );
  INV_X1 U2640 ( .A(n3722), .ZN(n3809) );
  OAI211_X1 U2641 ( .C1(n3521), .C2(n2564), .A(n2658), .B(n2657), .ZN(n3880)
         );
  OAI211_X1 U2642 ( .C1(n3948), .C2(n2709), .A(n2639), .B(n2638), .ZN(n4337)
         );
  INV_X1 U2643 ( .A(n4059), .ZN(n4524) );
  INV_X1 U2644 ( .A(n4363), .ZN(n4373) );
  INV_X1 U2645 ( .A(n4376), .ZN(n4073) );
  INV_X1 U2646 ( .A(n3398), .ZN(n3441) );
  INV_X1 U2647 ( .A(n3276), .ZN(n3744) );
  OR2_X1 U2648 ( .A1(n2294), .A2(n2917), .ZN(n3747) );
  NAND2_X1 U2649 ( .A1(n3754), .A2(n3753), .ZN(n3752) );
  NAND2_X1 U2650 ( .A1(n3031), .A2(n3032), .ZN(n3030) );
  NAND2_X1 U2651 ( .A1(n3752), .A2(n2984), .ZN(n3031) );
  XNOR2_X1 U2652 ( .A(n2987), .B(n2986), .ZN(n3762) );
  XNOR2_X1 U2653 ( .A(n3230), .B(n4712), .ZN(n4551) );
  NAND2_X1 U2654 ( .A1(n4551), .A2(REG2_REG_8__SCAN_IN), .ZN(n4550) );
  NAND2_X1 U2655 ( .A1(n4571), .A2(n3234), .ZN(n4582) );
  NAND2_X1 U2656 ( .A1(n4590), .A2(n3237), .ZN(n3336) );
  XNOR2_X1 U2657 ( .A(n3329), .B(n4704), .ZN(n4607) );
  XNOR2_X1 U2658 ( .A(n3784), .B(n3794), .ZN(n4615) );
  NOR2_X1 U2659 ( .A1(n4615), .A2(REG1_REG_16__SCAN_IN), .ZN(n4616) );
  NAND2_X1 U2660 ( .A1(n4611), .A2(n3796), .ZN(n4619) );
  INV_X1 U2661 ( .A(n2103), .ZN(n4626) );
  AND2_X1 U2662 ( .A1(n2980), .A2(n3021), .ZN(n4637) );
  AOI22_X1 U2663 ( .A1(n2899), .A2(n3693), .B1(n2898), .B2(n3848), .ZN(n2900)
         );
  NAND2_X1 U2664 ( .A1(n2171), .A2(n3680), .ZN(n3840) );
  NAND2_X1 U2665 ( .A1(n2158), .A2(n2033), .ZN(n2159) );
  NAND2_X1 U2666 ( .A1(n2545), .A2(n2562), .ZN(n4542) );
  NAND2_X1 U2667 ( .A1(n2172), .A2(n2175), .ZN(n4272) );
  NAND2_X1 U2668 ( .A1(n3372), .A2(n2178), .ZN(n2172) );
  NAND2_X1 U2669 ( .A1(n2180), .A2(n2182), .ZN(n4409) );
  NAND2_X1 U2670 ( .A1(n2181), .A2(n2037), .ZN(n2180) );
  INV_X1 U2671 ( .A(n4430), .ZN(n4281) );
  INV_X1 U2672 ( .A(n4647), .ZN(n4653) );
  NAND2_X1 U2673 ( .A1(n2156), .A2(n2154), .ZN(n3299) );
  INV_X1 U2674 ( .A(n2155), .ZN(n2154) );
  NAND2_X1 U2675 ( .A1(n2156), .A2(n2149), .ZN(n4728) );
  AOI21_X1 U2676 ( .B1(n3256), .B2(n2145), .A(n2064), .ZN(n4718) );
  NAND2_X1 U2677 ( .A1(n4022), .A2(n3176), .ZN(n4064) );
  INV_X1 U2678 ( .A(n3815), .ZN(n4282) );
  OR2_X1 U2679 ( .A1(n2946), .A2(n2779), .ZN(n4647) );
  INV_X1 U2680 ( .A(n3093), .ZN(n3073) );
  AND2_X1 U2681 ( .A1(n2763), .A2(n2764), .ZN(n3065) );
  AND2_X1 U2682 ( .A1(n4022), .A2(n4412), .ZN(n4279) );
  AND2_X2 U2683 ( .A1(n2893), .A2(n2892), .ZN(n4739) );
  AND2_X2 U2684 ( .A1(n2893), .A2(n3063), .ZN(n4733) );
  XNOR2_X1 U2685 ( .A(n2272), .B(IR_REG_25__SCAN_IN), .ZN(n2949) );
  XNOR2_X1 U2686 ( .A(n2286), .B(IR_REG_27__SCAN_IN), .ZN(n4513) );
  XNOR2_X1 U2687 ( .A(n2274), .B(IR_REG_26__SCAN_IN), .ZN(n2931) );
  INV_X1 U2688 ( .A(n2949), .ZN(n2934) );
  NAND2_X1 U2689 ( .A1(n2750), .A2(IR_REG_31__SCAN_IN), .ZN(n2276) );
  XNOR2_X1 U2690 ( .A(n2298), .B(IR_REG_22__SCAN_IN), .ZN(n3736) );
  INV_X1 U2691 ( .A(n2764), .ZN(n3727) );
  XNOR2_X1 U2692 ( .A(n2302), .B(n4241), .ZN(n3802) );
  AND2_X1 U2693 ( .A1(n2552), .A2(n2534), .ZN(n3339) );
  XNOR2_X1 U2694 ( .A(n2105), .B(IR_REG_1__SCAN_IN), .ZN(n4519) );
  NAND2_X1 U2695 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2105)
         );
  INV_X2 U2696 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  AND2_X1 U2697 ( .A1(n3436), .A2(n3435), .ZN(n2185) );
  NAND2_X1 U2698 ( .A1(n2087), .A2(n2043), .ZN(U3258) );
  OR2_X1 U2699 ( .A1(n2088), .A2(n4631), .ZN(n2087) );
  NAND2_X1 U2700 ( .A1(n2089), .A2(n4591), .ZN(n2088) );
  NAND2_X1 U2701 ( .A1(n2912), .A2(n2126), .ZN(U3547) );
  OR2_X1 U2702 ( .A1(n3820), .A2(n4440), .ZN(n2912) );
  AOI21_X1 U2703 ( .B1(n2128), .B2(n4739), .A(n2127), .ZN(n2126) );
  NOR2_X1 U2704 ( .A1(n4739), .A2(n2909), .ZN(n2127) );
  OR2_X1 U2705 ( .A1(n3826), .A2(n4440), .ZN(n2890) );
  OR2_X1 U2706 ( .A1(n3820), .A2(n4511), .ZN(n2915) );
  OR2_X1 U2707 ( .A1(n3826), .A2(n4511), .ZN(n2896) );
  NAND2_X2 U2708 ( .A1(n2294), .A2(n3066), .ZN(n2318) );
  CLKBUF_X3 U2709 ( .A(n4742), .Z(n2781) );
  OR2_X1 U2711 ( .A1(n4029), .A2(n2078), .ZN(n2027) );
  NAND2_X1 U2712 ( .A1(n3743), .A2(n3274), .ZN(n2028) );
  OR3_X1 U2713 ( .A1(n3884), .A2(n2076), .A3(n2067), .ZN(n2029) );
  OR2_X1 U2714 ( .A1(n2824), .A2(n4039), .ZN(n2030) );
  NAND2_X1 U2715 ( .A1(n3742), .A2(n3442), .ZN(n2032) );
  AND2_X1 U2716 ( .A1(n2030), .A2(n2232), .ZN(n2033) );
  OR3_X1 U2717 ( .A1(n4029), .A2(n3993), .A3(n4009), .ZN(n2034) );
  MUX2_X1 U2718 ( .A(n3328), .B(DATAI_14_), .S(n3651), .Z(n4381) );
  INV_X1 U2719 ( .A(n2318), .ZN(n2716) );
  INV_X1 U2720 ( .A(n2318), .ZN(n2710) );
  AND2_X1 U2721 ( .A1(n2223), .A2(n2249), .ZN(n2035) );
  NAND2_X1 U2722 ( .A1(n2279), .A2(n2250), .ZN(n2036) );
  NAND2_X1 U2723 ( .A1(n2474), .A2(n2245), .ZN(n2515) );
  OR2_X1 U2724 ( .A1(n4416), .A2(n3387), .ZN(n2037) );
  NOR2_X1 U2725 ( .A1(n2235), .A2(n2236), .ZN(n2038) );
  NAND2_X1 U2726 ( .A1(n2035), .A2(n2474), .ZN(n2283) );
  NAND2_X1 U2727 ( .A1(n4395), .A2(n3676), .ZN(n2039) );
  AND2_X1 U2728 ( .A1(n2120), .A2(n2863), .ZN(n2040) );
  AND2_X1 U2729 ( .A1(n2200), .A2(n3407), .ZN(n2041) );
  INV_X1 U2730 ( .A(n3716), .ZN(n3842) );
  AND2_X1 U2731 ( .A1(n4415), .A2(n4394), .ZN(n2042) );
  INV_X1 U2732 ( .A(n2798), .ZN(n2797) );
  INV_X1 U2733 ( .A(n3303), .ZN(n2189) );
  AND3_X1 U2734 ( .A1(n4640), .A2(n2086), .A3(n2085), .ZN(n2043) );
  OR2_X1 U2735 ( .A1(n3302), .A2(n3303), .ZN(n2044) );
  OR2_X1 U2736 ( .A1(n3475), .A2(n3152), .ZN(n2045) );
  OR2_X1 U2737 ( .A1(n3523), .A2(n3917), .ZN(n2046) );
  INV_X1 U2738 ( .A(n2116), .ZN(n2115) );
  AOI21_X1 U2739 ( .B1(n3842), .B2(n3649), .A(n2901), .ZN(n2116) );
  INV_X1 U2740 ( .A(n3649), .ZN(n2879) );
  AND2_X1 U2741 ( .A1(n2373), .A2(n2372), .ZN(n2047) );
  AND2_X1 U2742 ( .A1(n4430), .A2(n4407), .ZN(n2048) );
  NAND2_X1 U2743 ( .A1(n2825), .A2(n2039), .ZN(n2049) );
  AND2_X1 U2744 ( .A1(n3398), .A2(n3357), .ZN(n2050) );
  AND2_X1 U2745 ( .A1(n2035), .A2(n2138), .ZN(n2279) );
  NAND2_X1 U2746 ( .A1(n4524), .A2(n4359), .ZN(n2051) );
  INV_X1 U2747 ( .A(IR_REG_14__SCAN_IN), .ZN(n2245) );
  NOR2_X1 U2748 ( .A1(n3866), .A2(n3852), .ZN(n2052) );
  NOR2_X1 U2749 ( .A1(n3841), .A2(n2879), .ZN(n2053) );
  AND2_X1 U2750 ( .A1(n2044), .A2(n3439), .ZN(n2054) );
  AND2_X1 U2751 ( .A1(n2407), .A2(n2189), .ZN(n2055) );
  AND2_X1 U2752 ( .A1(n2121), .A2(n3719), .ZN(n2056) );
  NOR2_X1 U2753 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2057)
         );
  INV_X1 U2754 ( .A(IR_REG_2__SCAN_IN), .ZN(n2092) );
  OR2_X1 U2755 ( .A1(n2115), .A2(n3694), .ZN(n2058) );
  INV_X1 U2756 ( .A(n2564), .ZN(n2685) );
  INV_X1 U2757 ( .A(n2151), .ZN(n2152) );
  INV_X1 U2758 ( .A(n3667), .ZN(n2124) );
  INV_X1 U2759 ( .A(IR_REG_15__SCAN_IN), .ZN(n2247) );
  NAND2_X1 U2760 ( .A1(n2159), .A2(n2161), .ZN(n4027) );
  AND2_X1 U2761 ( .A1(n3293), .A2(n3357), .ZN(n2059) );
  AND2_X1 U2762 ( .A1(n4337), .A2(n3945), .ZN(n2060) );
  INV_X1 U2763 ( .A(n2077), .ZN(n4345) );
  NOR3_X1 U2764 ( .A1(n4029), .A2(n3993), .A3(n2080), .ZN(n2077) );
  AND2_X1 U2765 ( .A1(n2180), .A2(n2178), .ZN(n2061) );
  NAND2_X1 U2766 ( .A1(n2474), .A2(n2225), .ZN(n2062) );
  AND2_X1 U2767 ( .A1(n2633), .A2(n2632), .ZN(n2063) );
  INV_X1 U2768 ( .A(n3652), .ZN(n2141) );
  INV_X1 U2769 ( .A(IR_REG_0__SCAN_IN), .ZN(n2291) );
  INV_X1 U2770 ( .A(n4009), .ZN(n4016) );
  NAND2_X1 U2771 ( .A1(n3255), .A2(n3254), .ZN(n2064) );
  INV_X1 U2772 ( .A(n4704), .ZN(n3328) );
  NOR2_X1 U2773 ( .A1(n2590), .A2(n2589), .ZN(n2065) );
  NOR3_X1 U2774 ( .A1(n4275), .A2(n2074), .A3(n4522), .ZN(n2073) );
  OR2_X1 U2775 ( .A1(n3602), .A2(n2155), .ZN(n2153) );
  INV_X1 U2776 ( .A(n2153), .ZN(n2149) );
  NOR2_X1 U2777 ( .A1(n4275), .A2(n3676), .ZN(n2075) );
  INV_X1 U2778 ( .A(n3993), .ZN(n3998) );
  INV_X1 U2779 ( .A(n2178), .ZN(n2177) );
  AND2_X1 U2780 ( .A1(n2179), .A2(n2182), .ZN(n2178) );
  AND2_X1 U2781 ( .A1(n3684), .A2(n2145), .ZN(n2066) );
  AND2_X1 U2782 ( .A1(n2980), .A2(n2978), .ZN(n4591) );
  INV_X1 U2783 ( .A(n3869), .ZN(n3863) );
  INV_X1 U2784 ( .A(n2898), .ZN(n3833) );
  OR2_X1 U2785 ( .A1(n3817), .A2(n2898), .ZN(n2067) );
  INV_X1 U2786 ( .A(n4568), .ZN(n2083) );
  INV_X1 U2787 ( .A(n4589), .ZN(n2084) );
  INV_X1 U2788 ( .A(IR_REG_30__SCAN_IN), .ZN(n2258) );
  OR2_X1 U2789 ( .A1(n4698), .A2(n3787), .ZN(n2068) );
  INV_X1 U2790 ( .A(n4381), .ZN(n4098) );
  NAND2_X1 U2791 ( .A1(n2527), .A2(REG3_REG_15__SCAN_IN), .ZN(n2544) );
  NOR2_X2 U2792 ( .A1(n3942), .A2(n2060), .ZN(n3909) );
  NAND3_X1 U2793 ( .A1(n2033), .A2(n2163), .A3(n2826), .ZN(n2072) );
  NOR2_X2 U2794 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2319)
         );
  INV_X1 U2795 ( .A(n2073), .ZN(n4052) );
  INV_X1 U2796 ( .A(n2075), .ZN(n4120) );
  NAND3_X1 U2797 ( .A1(n2095), .A2(n2985), .A3(n2094), .ZN(n2987) );
  NAND3_X1 U2798 ( .A1(n3754), .A2(n3753), .A3(n3032), .ZN(n2094) );
  NAND3_X1 U2799 ( .A1(n2099), .A2(n2321), .A3(n2982), .ZN(n2098) );
  NAND2_X1 U2800 ( .A1(n3333), .A2(n3332), .ZN(n3782) );
  INV_X1 U2801 ( .A(n4625), .ZN(n2100) );
  NAND2_X1 U2802 ( .A1(n2103), .A2(n2101), .ZN(n4636) );
  NAND2_X1 U2803 ( .A1(n4636), .A2(n2068), .ZN(n3788) );
  INV_X1 U2804 ( .A(n2106), .ZN(n3211) );
  OAI21_X1 U2805 ( .B1(n2106), .B2(REG1_REG_7__SCAN_IN), .A(n4515), .ZN(n3209)
         );
  NAND2_X1 U2806 ( .A1(n3005), .A2(n4516), .ZN(n2107) );
  NAND2_X1 U2807 ( .A1(n2319), .A2(n2092), .ZN(n2320) );
  NAND2_X1 U2808 ( .A1(n3843), .A2(n2109), .ZN(n2108) );
  OAI211_X1 U2809 ( .C1(n3843), .C2(n2058), .A(n2110), .B(n2108), .ZN(n2907)
         );
  NOR2_X1 U2810 ( .A1(n3843), .A2(n3842), .ZN(n3841) );
  NAND2_X1 U2811 ( .A1(n2859), .A2(n2040), .ZN(n2117) );
  NAND2_X1 U2812 ( .A1(n2117), .A2(n2118), .ZN(n4056) );
  OAI21_X1 U2813 ( .B1(n3894), .B2(n2122), .A(n2056), .ZN(n2878) );
  NAND2_X1 U2814 ( .A1(n2865), .A2(n2131), .ZN(n3967) );
  NAND2_X1 U2815 ( .A1(n3967), .A2(n3704), .ZN(n2870) );
  OAI21_X1 U2816 ( .B1(n3312), .B2(n3610), .A(n3606), .ZN(n3373) );
  AOI21_X1 U2817 ( .B1(n3610), .B2(n3606), .A(n2137), .ZN(n2136) );
  NAND3_X1 U2818 ( .A1(n2035), .A2(n2138), .A3(n2226), .ZN(n2140) );
  AND2_X2 U2819 ( .A1(n2472), .A2(n2244), .ZN(n2474) );
  NAND2_X1 U2820 ( .A1(n3147), .A2(n3148), .ZN(n3146) );
  NAND2_X1 U2821 ( .A1(n2870), .A2(n3635), .ZN(n3910) );
  NAND2_X1 U2822 ( .A1(n2878), .A2(n2877), .ZN(n3843) );
  NAND2_X1 U2823 ( .A1(n2850), .A2(n3616), .ZN(n3312) );
  INV_X1 U2824 ( .A(n4025), .ZN(n2865) );
  NAND2_X4 U2825 ( .A1(n2262), .A2(n2261), .ZN(n3652) );
  XNOR2_X2 U2826 ( .A(n2142), .B(n2258), .ZN(n2261) );
  OAI21_X1 U2827 ( .B1(n2151), .B2(n3272), .A(n2150), .ZN(n2814) );
  OAI22_X1 U2828 ( .A1(n3602), .A2(n2147), .B1(n2050), .B2(n2032), .ZN(n2150)
         );
  OR2_X1 U2829 ( .A1(n2155), .A2(n2050), .ZN(n2147) );
  CLKBUF_X1 U2830 ( .A(n2163), .Z(n2158) );
  NAND2_X1 U2831 ( .A1(n3857), .A2(n3679), .ZN(n2171) );
  NAND4_X1 U2832 ( .A1(n2035), .A2(n2474), .A3(n2228), .A4(n2031), .ZN(n2273)
         );
  OAI21_X1 U2833 ( .B1(n3437), .B2(n3584), .A(n2185), .ZN(U3211) );
  NAND2_X1 U2834 ( .A1(n2186), .A2(n2187), .ZN(n3349) );
  NAND2_X1 U2835 ( .A1(n3440), .A2(n2054), .ZN(n2186) );
  NAND2_X1 U2836 ( .A1(n3470), .A2(n2194), .ZN(n2192) );
  NAND2_X1 U2837 ( .A1(n2192), .A2(n2193), .ZN(n3165) );
  NAND2_X1 U2838 ( .A1(n3386), .A2(n2041), .ZN(n2197) );
  NAND2_X1 U2839 ( .A1(n2197), .A2(n2198), .ZN(n3414) );
  NAND2_X1 U2840 ( .A1(n3554), .A2(n2206), .ZN(n2204) );
  NAND2_X1 U2841 ( .A1(n2560), .A2(n2559), .ZN(n3510) );
  INV_X1 U2842 ( .A(n2559), .ZN(n2217) );
  OAI21_X1 U2843 ( .B1(n3529), .B2(n2220), .A(n2218), .ZN(n3556) );
  AND2_X1 U2844 ( .A1(n2279), .A2(n2229), .ZN(n2269) );
  NAND2_X1 U2845 ( .A1(n2801), .A2(n2844), .ZN(n3105) );
  NAND2_X1 U2846 ( .A1(n3589), .A2(n3586), .ZN(n2842) );
  MUX2_X1 U2847 ( .A(n2777), .B(n2776), .S(IR_REG_28__SCAN_IN), .Z(n4521) );
  AOI22_X2 U2848 ( .A1(n3876), .A2(n2835), .B1(n3879), .B2(n3900), .ZN(n3857)
         );
  INV_X1 U2849 ( .A(n2540), .ZN(n2543) );
  NAND2_X2 U2850 ( .A1(n2817), .A2(n2816), .ZN(n3372) );
  XNOR2_X1 U2851 ( .A(n2310), .B(n2729), .ZN(n2312) );
  AND2_X1 U2852 ( .A1(n3651), .A2(DATAI_30_), .ZN(n4296) );
  AND2_X1 U2853 ( .A1(n3651), .A2(DATAI_28_), .ZN(n2898) );
  AND2_X1 U2854 ( .A1(n3651), .A2(DATAI_21_), .ZN(n4336) );
  AND2_X1 U2855 ( .A1(n3651), .A2(DATAI_20_), .ZN(n3977) );
  AND2_X1 U2856 ( .A1(n3651), .A2(DATAI_27_), .ZN(n4302) );
  NAND2_X1 U2857 ( .A1(n3651), .A2(DATAI_23_), .ZN(n3917) );
  NAND2_X1 U2858 ( .A1(n3651), .A2(DATAI_0_), .ZN(n2292) );
  OR2_X1 U2859 ( .A1(n3651), .A2(n2291), .ZN(n2293) );
  NAND2_X1 U2860 ( .A1(n3651), .A2(DATAI_24_), .ZN(n3904) );
  NAND2_X1 U2861 ( .A1(n4524), .A2(n4034), .ZN(n2230) );
  AND2_X1 U2862 ( .A1(n4239), .A2(n2237), .ZN(n2231) );
  OR2_X1 U2863 ( .A1(n4395), .A2(n3676), .ZN(n2232) );
  AND2_X1 U2864 ( .A1(n2391), .A2(n2390), .ZN(n2233) );
  AND2_X1 U2865 ( .A1(n3988), .A2(n2866), .ZN(n2234) );
  INV_X1 U2866 ( .A(IR_REG_28__SCAN_IN), .ZN(n2287) );
  NOR2_X1 U2867 ( .A1(n2670), .A2(n3516), .ZN(n2235) );
  NOR2_X1 U2868 ( .A1(n2668), .A2(n2669), .ZN(n2236) );
  NAND2_X1 U2869 ( .A1(n2799), .A2(n3083), .ZN(n3586) );
  INV_X1 U2870 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2507) );
  OAI22_X1 U2871 ( .A1(n2797), .A2(n2678), .B1(n3083), .B2(n2026), .ZN(n2310)
         );
  INV_X1 U2872 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2466) );
  INV_X1 U2873 ( .A(IR_REG_13__SCAN_IN), .ZN(n2244) );
  INV_X1 U2874 ( .A(IR_REG_18__SCAN_IN), .ZN(n2249) );
  INV_X1 U2875 ( .A(n2452), .ZN(n2453) );
  OR2_X1 U2876 ( .A1(n2622), .A2(n3492), .ZN(n2634) );
  OR2_X1 U2877 ( .A1(n2360), .A2(n4734), .ZN(n2345) );
  AND2_X1 U2878 ( .A1(n2578), .A2(REG3_REG_18__SCAN_IN), .ZN(n2607) );
  NAND2_X1 U2879 ( .A1(n2697), .A2(n2696), .ZN(n2702) );
  INV_X1 U2880 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3492) );
  AND2_X1 U2881 ( .A1(n2296), .A2(n2295), .ZN(n2303) );
  INV_X1 U2882 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3558) );
  OR2_X1 U2883 ( .A1(n2683), .A2(n3571), .ZN(n2703) );
  AND2_X1 U2884 ( .A1(n2644), .A2(REG3_REG_23__SCAN_IN), .ZN(n2654) );
  NOR2_X1 U2885 ( .A1(n2634), .A2(n3558), .ZN(n2644) );
  NAND2_X1 U2886 ( .A1(n2304), .A2(REG1_REG_2__SCAN_IN), .ZN(n2315) );
  INV_X1 U2887 ( .A(n4521), .ZN(n3020) );
  INV_X1 U2888 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2979) );
  INV_X1 U2889 ( .A(REG3_REG_8__SCAN_IN), .ZN(n3306) );
  INV_X1 U2890 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4528) );
  AND2_X1 U2891 ( .A1(n3651), .A2(n2943), .ZN(n2957) );
  INV_X1 U2892 ( .A(n3841), .ZN(n3845) );
  AND2_X1 U2893 ( .A1(n3665), .A2(n3858), .ZN(n3877) );
  OR2_X1 U2894 ( .A1(n3911), .A2(n3670), .ZN(n3957) );
  NAND2_X1 U2895 ( .A1(n4005), .A2(n4008), .ZN(n4004) );
  INV_X1 U2896 ( .A(n4279), .ZN(n4097) );
  AND2_X1 U2897 ( .A1(n2848), .A2(n3612), .ZN(n3602) );
  INV_X1 U2898 ( .A(n2885), .ZN(n2779) );
  INV_X1 U2899 ( .A(n4429), .ZN(n4414) );
  AND2_X1 U2900 ( .A1(n2734), .A2(n2952), .ZN(n2737) );
  INV_X1 U2901 ( .A(n2948), .ZN(n2749) );
  INV_X1 U2902 ( .A(n4522), .ZN(n4050) );
  INV_X1 U2903 ( .A(n4394), .ZN(n4273) );
  NAND2_X1 U2904 ( .A1(n4521), .A2(n2942), .ZN(n4429) );
  XNOR2_X1 U2905 ( .A(n2276), .B(n2275), .ZN(n2734) );
  NAND2_X1 U2906 ( .A1(n2521), .A2(n2519), .ZN(n3455) );
  AND2_X1 U2907 ( .A1(n3651), .A2(DATAI_25_), .ZN(n3879) );
  INV_X1 U2908 ( .A(n4034), .ZN(n4359) );
  AND2_X1 U2909 ( .A1(n3651), .A2(DATAI_22_), .ZN(n3945) );
  OAI21_X1 U2910 ( .B1(n3054), .B2(n3053), .A(n2313), .ZN(n3100) );
  AND2_X1 U2911 ( .A1(n2703), .A2(n2684), .ZN(n3871) );
  OR2_X1 U2912 ( .A1(n2318), .A2(n2772), .ZN(n3734) );
  AND2_X1 U2913 ( .A1(n2958), .A2(n2957), .ZN(n2980) );
  INV_X1 U2914 ( .A(n4643), .ZN(n4657) );
  INV_X1 U2915 ( .A(n4064), .ZN(n4290) );
  AND2_X1 U2916 ( .A1(n4022), .A2(n4414), .ZN(n4280) );
  AOI21_X1 U2917 ( .B1(n2749), .B2(n2738), .A(n2737), .ZN(n2892) );
  INV_X1 U2918 ( .A(n4302), .ZN(n3852) );
  INV_X1 U2919 ( .A(n4724), .ZN(n4350) );
  INV_X1 U2920 ( .A(n4372), .ZN(n4078) );
  AND3_X1 U2921 ( .A1(n2887), .A2(n2886), .A3(n3060), .ZN(n2893) );
  NAND2_X1 U2922 ( .A1(n2736), .A2(n2931), .ZN(n2948) );
  INV_X1 U2923 ( .A(n3223), .ZN(n3325) );
  AND2_X1 U2924 ( .A1(n2945), .A2(n2958), .ZN(n4635) );
  NAND2_X1 U2925 ( .A1(n2769), .A2(STATE_REG_SCAN_IN), .ZN(n4543) );
  INV_X1 U2926 ( .A(n4538), .ZN(n3584) );
  INV_X1 U2927 ( .A(n3997), .ZN(n4360) );
  INV_X1 U2928 ( .A(n4591), .ZN(n4630) );
  NAND2_X1 U2929 ( .A1(n2980), .A2(n4521), .ZN(n4641) );
  OR2_X1 U2930 ( .A1(n4018), .A2(n4719), .ZN(n4643) );
  AND2_X2 U2931 ( .A1(n3064), .A2(n4647), .ZN(n4663) );
  INV_X1 U2932 ( .A(n4739), .ZN(n4737) );
  INV_X1 U2933 ( .A(n4733), .ZN(n4732) );
  AND2_X2 U2934 ( .A1(n2948), .A2(n2947), .ZN(n4694) );
  AND2_X1 U2935 ( .A1(n2944), .A2(STATE_REG_SCAN_IN), .ZN(n4695) );
  OR2_X1 U2936 ( .A1(n2517), .A2(n2516), .ZN(n4704) );
  INV_X2 U2937 ( .A(n3747), .ZN(U4043) );
  INV_X1 U2938 ( .A(n2320), .ZN(n2238) );
  NAND2_X1 U2939 ( .A1(n2238), .A2(n2231), .ZN(n2366) );
  NOR2_X1 U2940 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2242)
         );
  NOR2_X1 U2941 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2241)
         );
  NOR2_X1 U2942 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2240)
         );
  NOR2_X1 U2943 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2239)
         );
  NAND4_X1 U2944 ( .A1(n2242), .A2(n2241), .A3(n2240), .A4(n2239), .ZN(n2243)
         );
  NOR2_X2 U2945 ( .A1(n2366), .A2(n2243), .ZN(n2472) );
  NAND2_X1 U2946 ( .A1(n2777), .A2(n2254), .ZN(n2256) );
  XNOR2_X2 U2947 ( .A(n2256), .B(n2255), .ZN(n2260) );
  NOR2_X1 U2948 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2257)
         );
  NAND2_X1 U2949 ( .A1(n2775), .A2(n2257), .ZN(n2928) );
  NAND2_X1 U2951 ( .A1(n4742), .A2(REG2_REG_0__SCAN_IN), .ZN(n2268) );
  INV_X1 U2952 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2959) );
  OR2_X1 U2953 ( .A1(n2360), .A2(n2959), .ZN(n2267) );
  INV_X1 U2954 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2263) );
  OR2_X1 U2955 ( .A1(n3652), .A2(n2263), .ZN(n2266) );
  NAND2_X2 U2956 ( .A1(n2260), .A2(n2939), .ZN(n2564) );
  INV_X1 U2957 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2264) );
  OR2_X1 U2958 ( .A1(n2564), .A2(n2264), .ZN(n2265) );
  NAND2_X1 U2959 ( .A1(n2270), .A2(IR_REG_31__SCAN_IN), .ZN(n2271) );
  NAND2_X1 U2960 ( .A1(n2751), .A2(n2271), .ZN(n2272) );
  NAND2_X1 U2961 ( .A1(n2273), .A2(IR_REG_31__SCAN_IN), .ZN(n2274) );
  INV_X1 U2962 ( .A(n2279), .ZN(n2280) );
  NAND2_X1 U2963 ( .A1(n2280), .A2(IR_REG_31__SCAN_IN), .ZN(n2281) );
  MUX2_X1 U2964 ( .A(IR_REG_31__SCAN_IN), .B(n2281), .S(IR_REG_21__SCAN_IN), 
        .Z(n2282) );
  NAND2_X1 U2965 ( .A1(n2283), .A2(IR_REG_31__SCAN_IN), .ZN(n2302) );
  NAND2_X1 U2966 ( .A1(n2302), .A2(n4241), .ZN(n2284) );
  INV_X1 U2967 ( .A(n2837), .ZN(n3066) );
  NAND2_X1 U2968 ( .A1(n3748), .A2(n2710), .ZN(n2296) );
  NAND2_X1 U2969 ( .A1(n2287), .A2(IR_REG_27__SCAN_IN), .ZN(n2288) );
  NAND2_X1 U2970 ( .A1(n3093), .A2(n2711), .ZN(n2295) );
  OR2_X1 U2971 ( .A1(n2294), .A2(n2959), .ZN(n2297) );
  NAND2_X1 U2972 ( .A1(n2303), .A2(n2297), .ZN(n3019) );
  NAND2_X1 U2973 ( .A1(n2036), .A2(IR_REG_31__SCAN_IN), .ZN(n2298) );
  NAND2_X1 U2974 ( .A1(n3748), .A2(n2718), .ZN(n2301) );
  NOR2_X1 U2975 ( .A1(n2294), .A2(n2291), .ZN(n2299) );
  AOI21_X1 U2976 ( .B1(n3093), .B2(n2716), .A(n2299), .ZN(n2300) );
  NAND2_X1 U2977 ( .A1(n2301), .A2(n2300), .ZN(n3018) );
  NAND2_X1 U2978 ( .A1(n3736), .A2(n3802), .ZN(n2770) );
  AOI22_X1 U2979 ( .A1(n3019), .A2(n3018), .B1(n2303), .B2(n2714), .ZN(n3054)
         );
  NAND2_X1 U2980 ( .A1(n2304), .A2(REG1_REG_1__SCAN_IN), .ZN(n2309) );
  INV_X1 U2981 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2305) );
  INV_X1 U2982 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3124) );
  NAND2_X1 U2983 ( .A1(n4742), .A2(REG2_REG_1__SCAN_IN), .ZN(n2306) );
  MUX2_X1 U2984 ( .A(n4519), .B(DATAI_1_), .S(n3651), .Z(n3126) );
  OAI22_X1 U2985 ( .A1(n2797), .A2(n2731), .B1(n3083), .B2(n2678), .ZN(n2311)
         );
  XNOR2_X1 U2986 ( .A(n2312), .B(n2311), .ZN(n3053) );
  NAND2_X1 U2987 ( .A1(n2312), .A2(n2311), .ZN(n2313) );
  INV_X1 U2988 ( .A(n3100), .ZN(n2329) );
  NAND2_X1 U2989 ( .A1(n4742), .A2(REG2_REG_2__SCAN_IN), .ZN(n2317) );
  INV_X1 U2990 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3136) );
  OR2_X1 U2991 ( .A1(n2564), .A2(n3136), .ZN(n2316) );
  INV_X1 U2992 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3115) );
  OR2_X1 U2993 ( .A1(n3652), .A2(n3115), .ZN(n2314) );
  INV_X1 U2994 ( .A(n2321), .ZN(n2322) );
  MUX2_X1 U2995 ( .A(n4518), .B(DATAI_2_), .S(n3651), .Z(n3152) );
  OAI22_X1 U2996 ( .A1(n3084), .A2(n2678), .B1(n3137), .B2(n2026), .ZN(n2324)
         );
  XNOR2_X1 U2997 ( .A(n2324), .B(n2729), .ZN(n2326) );
  OAI22_X1 U2998 ( .A1(n3084), .A2(n2731), .B1(n3137), .B2(n2678), .ZN(n2325)
         );
  OR2_X1 U2999 ( .A1(n2326), .A2(n2325), .ZN(n2330) );
  NAND2_X1 U3000 ( .A1(n2326), .A2(n2325), .ZN(n2327) );
  NAND2_X1 U3001 ( .A1(n2330), .A2(n2327), .ZN(n3099) );
  NAND2_X1 U3002 ( .A1(n2329), .A2(n2328), .ZN(n3097) );
  NAND2_X1 U3003 ( .A1(n3097), .A2(n2330), .ZN(n3471) );
  NAND2_X1 U3004 ( .A1(n4742), .A2(REG2_REG_3__SCAN_IN), .ZN(n2335) );
  OR2_X1 U3005 ( .A1(n2564), .A2(REG3_REG_3__SCAN_IN), .ZN(n2334) );
  INV_X1 U3006 ( .A(REG1_REG_3__SCAN_IN), .ZN(n3156) );
  OR2_X1 U3007 ( .A1(n2360), .A2(n3156), .ZN(n2333) );
  INV_X1 U3008 ( .A(REG0_REG_3__SCAN_IN), .ZN(n3159) );
  OR2_X1 U3009 ( .A1(n3652), .A2(n3159), .ZN(n2332) );
  NAND2_X1 U3010 ( .A1(n3745), .A2(n2710), .ZN(n2337) );
  NAND2_X1 U3011 ( .A1(n2321), .A2(IR_REG_31__SCAN_IN), .ZN(n2347) );
  XNOR2_X1 U3012 ( .A(n2347), .B(IR_REG_3__SCAN_IN), .ZN(n3759) );
  MUX2_X1 U3013 ( .A(n3759), .B(DATAI_3_), .S(n3651), .Z(n3475) );
  NAND2_X1 U3014 ( .A1(n3475), .A2(n2711), .ZN(n2336) );
  NAND2_X1 U3015 ( .A1(n2337), .A2(n2336), .ZN(n2338) );
  XNOR2_X1 U3016 ( .A(n2338), .B(n2729), .ZN(n2351) );
  AOI22_X1 U3017 ( .A1(n3745), .A2(n2718), .B1(n3475), .B2(n2710), .ZN(n2352)
         );
  XNOR2_X1 U3018 ( .A(n2351), .B(n2352), .ZN(n3472) );
  NAND2_X1 U3019 ( .A1(n4742), .A2(REG2_REG_4__SCAN_IN), .ZN(n2346) );
  INV_X1 U3020 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2339) );
  INV_X1 U3021 ( .A(n2361), .ZN(n2342) );
  INV_X1 U3022 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3474) );
  INV_X1 U3023 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2340) );
  NAND2_X1 U3024 ( .A1(n3474), .A2(n2340), .ZN(n2341) );
  NAND2_X1 U3025 ( .A1(n2342), .A2(n2341), .ZN(n3267) );
  OR2_X1 U3026 ( .A1(n2564), .A2(n3267), .ZN(n2343) );
  NAND2_X1 U3027 ( .A1(n2347), .A2(n4239), .ZN(n2348) );
  NAND2_X1 U3028 ( .A1(n2348), .A2(IR_REG_31__SCAN_IN), .ZN(n2349) );
  XNOR2_X1 U3029 ( .A(n2349), .B(IR_REG_4__SCAN_IN), .ZN(n4517) );
  MUX2_X1 U3030 ( .A(n4517), .B(DATAI_4_), .S(n3651), .Z(n3258) );
  OAI22_X1 U3031 ( .A1(n2802), .A2(n2678), .B1(n3265), .B2(n2026), .ZN(n2350)
         );
  XNOR2_X1 U3032 ( .A(n2350), .B(n2714), .ZN(n2355) );
  OAI22_X1 U3033 ( .A1(n2802), .A2(n2731), .B1(n3265), .B2(n2678), .ZN(n2356)
         );
  XNOR2_X1 U3034 ( .A(n2355), .B(n2356), .ZN(n3189) );
  INV_X1 U3035 ( .A(n2351), .ZN(n2353) );
  NAND2_X1 U3036 ( .A1(n2353), .A2(n2352), .ZN(n3190) );
  AND2_X1 U3037 ( .A1(n3189), .A2(n3190), .ZN(n2354) );
  INV_X1 U3038 ( .A(n2355), .ZN(n2357) );
  NAND2_X1 U3039 ( .A1(n2357), .A2(n2356), .ZN(n2358) );
  NAND2_X1 U3040 ( .A1(n2781), .A2(REG2_REG_5__SCAN_IN), .ZN(n2365) );
  INV_X1 U3041 ( .A(REG0_REG_5__SCAN_IN), .ZN(n2359) );
  OR2_X1 U3042 ( .A1(n3652), .A2(n2359), .ZN(n2364) );
  INV_X1 U3043 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2991) );
  OR2_X1 U3044 ( .A1(n2360), .A2(n2991), .ZN(n2363) );
  NAND2_X1 U3045 ( .A1(n2361), .A2(REG3_REG_5__SCAN_IN), .ZN(n2376) );
  OAI21_X1 U3046 ( .B1(n2361), .B2(REG3_REG_5__SCAN_IN), .A(n2376), .ZN(n3178)
         );
  OR2_X1 U3047 ( .A1(n2709), .A2(n3178), .ZN(n2362) );
  NAND2_X1 U3048 ( .A1(n2366), .A2(IR_REG_31__SCAN_IN), .ZN(n2368) );
  INV_X1 U3049 ( .A(IR_REG_5__SCAN_IN), .ZN(n2367) );
  XNOR2_X1 U3050 ( .A(n2368), .B(n2367), .ZN(n3770) );
  INV_X1 U3051 ( .A(DATAI_5_), .ZN(n2369) );
  MUX2_X1 U3052 ( .A(n3770), .B(n2369), .S(n3651), .Z(n2846) );
  OAI22_X1 U3053 ( .A1(n3276), .A2(n2678), .B1(n2846), .B2(n2026), .ZN(n2370)
         );
  XNOR2_X1 U3054 ( .A(n2370), .B(n2714), .ZN(n2371) );
  OAI22_X1 U3055 ( .A1(n3276), .A2(n2731), .B1(n2846), .B2(n2678), .ZN(n2372)
         );
  XNOR2_X1 U3056 ( .A(n2371), .B(n2372), .ZN(n3118) );
  INV_X1 U3057 ( .A(n2371), .ZN(n2373) );
  INV_X1 U3058 ( .A(n3165), .ZN(n2393) );
  NAND2_X1 U3059 ( .A1(n2781), .A2(REG2_REG_6__SCAN_IN), .ZN(n2381) );
  INV_X1 U3060 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2374) );
  OR2_X1 U3061 ( .A1(n3652), .A2(n2374), .ZN(n2380) );
  INV_X1 U3062 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2375) );
  OR2_X1 U3063 ( .A1(n2360), .A2(n2375), .ZN(n2379) );
  AND2_X1 U3064 ( .A1(n2376), .A2(n2979), .ZN(n2377) );
  NOR2_X1 U3065 ( .A1(n2376), .A2(n2979), .ZN(n2395) );
  OR2_X1 U3066 ( .A1(n2377), .A2(n2395), .ZN(n3283) );
  OR2_X1 U3067 ( .A1(n2564), .A2(n3283), .ZN(n2378) );
  NAND4_X1 U3068 ( .A1(n2381), .A2(n2380), .A3(n2379), .A4(n2378), .ZN(n3743)
         );
  NAND2_X1 U3069 ( .A1(n3743), .A2(n2710), .ZN(n2384) );
  NOR2_X1 U3070 ( .A1(n2366), .A2(IR_REG_5__SCAN_IN), .ZN(n2402) );
  OR2_X1 U3071 ( .A1(n2402), .A2(n2774), .ZN(n2382) );
  XNOR2_X1 U3072 ( .A(n2382), .B(IR_REG_6__SCAN_IN), .ZN(n4516) );
  MUX2_X1 U3073 ( .A(n4516), .B(DATAI_6_), .S(n3651), .Z(n3274) );
  NAND2_X1 U3074 ( .A1(n3274), .A2(n2711), .ZN(n2383) );
  NAND2_X1 U3075 ( .A1(n2384), .A2(n2383), .ZN(n2385) );
  XNOR2_X1 U3076 ( .A(n2385), .B(n2729), .ZN(n2388) );
  NAND2_X1 U3077 ( .A1(n3743), .A2(n2718), .ZN(n2387) );
  NAND2_X1 U3078 ( .A1(n3274), .A2(n2710), .ZN(n2386) );
  NAND2_X1 U3079 ( .A1(n2387), .A2(n2386), .ZN(n2389) );
  AND2_X1 U3080 ( .A1(n2388), .A2(n2389), .ZN(n3163) );
  INV_X1 U3081 ( .A(n3163), .ZN(n2392) );
  INV_X1 U3082 ( .A(n2388), .ZN(n2391) );
  INV_X1 U3083 ( .A(n2389), .ZN(n2390) );
  NAND2_X1 U3084 ( .A1(n2781), .A2(REG2_REG_7__SCAN_IN), .ZN(n2400) );
  INV_X1 U3085 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2394) );
  OR2_X1 U3086 ( .A1(n3652), .A2(n2394), .ZN(n2399) );
  INV_X1 U3087 ( .A(REG1_REG_7__SCAN_IN), .ZN(n3210) );
  OR2_X1 U3088 ( .A1(n2360), .A2(n3210), .ZN(n2398) );
  OR2_X1 U3089 ( .A1(n2395), .A2(REG3_REG_7__SCAN_IN), .ZN(n2396) );
  NAND2_X1 U3090 ( .A1(n2408), .A2(n2396), .ZN(n3443) );
  OR2_X1 U3091 ( .A1(n2709), .A2(n3443), .ZN(n2397) );
  NAND2_X1 U3092 ( .A1(n2402), .A2(n2401), .ZN(n2430) );
  NAND2_X1 U3093 ( .A1(n2430), .A2(IR_REG_31__SCAN_IN), .ZN(n2417) );
  XNOR2_X1 U3094 ( .A(n2417), .B(IR_REG_7__SCAN_IN), .ZN(n4515) );
  MUX2_X1 U3095 ( .A(n4515), .B(DATAI_7_), .S(n3651), .Z(n3442) );
  OAI22_X1 U3096 ( .A1(n2812), .A2(n2678), .B1(n2026), .B2(n3293), .ZN(n2403)
         );
  XNOR2_X1 U3097 ( .A(n2403), .B(n2714), .ZN(n2404) );
  OAI22_X1 U3098 ( .A1(n2812), .A2(n2731), .B1(n2678), .B2(n3293), .ZN(n2405)
         );
  XNOR2_X1 U3099 ( .A(n2404), .B(n2405), .ZN(n3439) );
  INV_X1 U3100 ( .A(n2404), .ZN(n2406) );
  NAND2_X1 U3101 ( .A1(n2406), .A2(n2405), .ZN(n2407) );
  NAND2_X1 U3102 ( .A1(n2781), .A2(REG2_REG_8__SCAN_IN), .ZN(n2415) );
  NAND2_X1 U3103 ( .A1(n2408), .A2(n3306), .ZN(n2409) );
  AND2_X1 U3104 ( .A1(n2424), .A2(n2409), .ZN(n4654) );
  INV_X1 U3105 ( .A(n4654), .ZN(n3307) );
  OR2_X1 U3106 ( .A1(n2709), .A2(n3307), .ZN(n2414) );
  INV_X1 U3107 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2410) );
  OR2_X1 U3108 ( .A1(n2360), .A2(n2410), .ZN(n2413) );
  INV_X1 U3109 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2411) );
  OR2_X1 U3110 ( .A1(n3652), .A2(n2411), .ZN(n2412) );
  OR2_X1 U3111 ( .A1(n3398), .A2(n2731), .ZN(n2421) );
  INV_X1 U3112 ( .A(IR_REG_7__SCAN_IN), .ZN(n2416) );
  NAND2_X1 U3113 ( .A1(n2417), .A2(n2416), .ZN(n2418) );
  NAND2_X1 U3114 ( .A1(n2418), .A2(IR_REG_31__SCAN_IN), .ZN(n2419) );
  XNOR2_X1 U3115 ( .A(n2419), .B(IR_REG_8__SCAN_IN), .ZN(n3229) );
  INV_X1 U3116 ( .A(n3229), .ZN(n4712) );
  INV_X1 U3117 ( .A(DATAI_8_), .ZN(n4711) );
  MUX2_X1 U3118 ( .A(n4712), .B(n4711), .S(n3651), .Z(n3357) );
  INV_X1 U3119 ( .A(n3357), .ZN(n3361) );
  NAND2_X1 U3120 ( .A1(n3361), .A2(n2716), .ZN(n2420) );
  NAND2_X1 U3121 ( .A1(n2421), .A2(n2420), .ZN(n3303) );
  OAI22_X1 U3122 ( .A1(n3398), .A2(n2678), .B1(n3357), .B2(n2026), .ZN(n2422)
         );
  XNOR2_X1 U3123 ( .A(n2422), .B(n2729), .ZN(n3302) );
  NAND2_X1 U3124 ( .A1(n2781), .A2(REG2_REG_9__SCAN_IN), .ZN(n2429) );
  AND2_X1 U3125 ( .A1(n2424), .A2(n2423), .ZN(n2425) );
  OR2_X1 U3126 ( .A1(n2425), .A2(n2437), .ZN(n3351) );
  OR2_X1 U3127 ( .A1(n2709), .A2(n3351), .ZN(n2428) );
  OR2_X1 U3128 ( .A1(n2360), .A2(n4186), .ZN(n2427) );
  INV_X1 U3129 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3401) );
  OR2_X1 U3130 ( .A1(n3652), .A2(n3401), .ZN(n2426) );
  NAND4_X1 U3131 ( .A1(n2429), .A2(n2428), .A3(n2427), .A4(n2426), .ZN(n4433)
         );
  NAND2_X1 U3132 ( .A1(n4433), .A2(n2716), .ZN(n2433) );
  NAND2_X1 U3133 ( .A1(n2443), .A2(IR_REG_31__SCAN_IN), .ZN(n2431) );
  XNOR2_X1 U3134 ( .A(n2431), .B(IR_REG_9__SCAN_IN), .ZN(n3226) );
  MUX2_X1 U3135 ( .A(n3226), .B(DATAI_9_), .S(n3651), .Z(n3395) );
  NAND2_X1 U3136 ( .A1(n3395), .A2(n2711), .ZN(n2432) );
  NAND2_X1 U3137 ( .A1(n2433), .A2(n2432), .ZN(n2434) );
  XNOR2_X1 U3138 ( .A(n2434), .B(n2714), .ZN(n2449) );
  AOI22_X1 U3139 ( .A1(n4433), .A2(n2718), .B1(n3395), .B2(n2710), .ZN(n2448)
         );
  XNOR2_X1 U3140 ( .A(n2449), .B(n2448), .ZN(n3350) );
  NAND2_X1 U3141 ( .A1(n2781), .A2(REG2_REG_10__SCAN_IN), .ZN(n2442) );
  INV_X1 U3142 ( .A(REG0_REG_10__SCAN_IN), .ZN(n2435) );
  OR2_X1 U3143 ( .A1(n3652), .A2(n2435), .ZN(n2441) );
  INV_X1 U3144 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2436) );
  OR2_X1 U3145 ( .A1(n2360), .A2(n2436), .ZN(n2440) );
  NOR2_X1 U3146 ( .A1(n2437), .A2(REG3_REG_10__SCAN_IN), .ZN(n2438) );
  OR2_X1 U3147 ( .A1(n2455), .A2(n2438), .ZN(n3389) );
  OR2_X1 U31480 ( .A1(n2709), .A2(n3389), .ZN(n2439) );
  NAND4_X1 U31490 ( .A1(n2442), .A2(n2441), .A3(n2440), .A4(n2439), .ZN(n4416)
         );
  NAND2_X1 U3150 ( .A1(n4416), .A2(n2710), .ZN(n2446) );
  NOR2_X1 U3151 ( .A1(n2443), .A2(IR_REG_9__SCAN_IN), .ZN(n2461) );
  OR2_X1 U3152 ( .A1(n2461), .A2(n2774), .ZN(n2444) );
  XNOR2_X1 U3153 ( .A(n2444), .B(IR_REG_10__SCAN_IN), .ZN(n4568) );
  MUX2_X1 U3154 ( .A(n4568), .B(DATAI_10_), .S(n3651), .Z(n3387) );
  NAND2_X1 U3155 ( .A1(n3387), .A2(n2711), .ZN(n2445) );
  NAND2_X1 U3156 ( .A1(n2446), .A2(n2445), .ZN(n2447) );
  XNOR2_X1 U3157 ( .A(n2447), .B(n2729), .ZN(n2451) );
  AOI22_X1 U3158 ( .A1(n4416), .A2(n2718), .B1(n2716), .B2(n3387), .ZN(n2452)
         );
  XNOR2_X1 U3159 ( .A(n2451), .B(n2452), .ZN(n3384) );
  NAND2_X1 U3160 ( .A1(n2449), .A2(n2448), .ZN(n3385) );
  AND2_X1 U3161 ( .A1(n3384), .A2(n3385), .ZN(n2450) );
  NAND2_X1 U3162 ( .A1(n2781), .A2(REG2_REG_11__SCAN_IN), .ZN(n2460) );
  NAND2_X1 U3163 ( .A1(n2455), .A2(REG3_REG_11__SCAN_IN), .ZN(n2484) );
  OR2_X1 U3164 ( .A1(n2455), .A2(REG3_REG_11__SCAN_IN), .ZN(n2456) );
  NAND2_X1 U3165 ( .A1(n2484), .A2(n2456), .ZN(n4648) );
  OR2_X1 U3166 ( .A1(n2709), .A2(n4648), .ZN(n2459) );
  INV_X1 U3167 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4425) );
  OR2_X1 U3168 ( .A1(n2360), .A2(n4425), .ZN(n2458) );
  INV_X1 U3169 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4507) );
  OR2_X1 U3170 ( .A1(n3652), .A2(n4507), .ZN(n2457) );
  NAND2_X1 U3171 ( .A1(n2461), .A2(n4240), .ZN(n2462) );
  NAND2_X1 U3172 ( .A1(n2462), .A2(IR_REG_31__SCAN_IN), .ZN(n2492) );
  XNOR2_X1 U3173 ( .A(n2492), .B(IR_REG_11__SCAN_IN), .ZN(n3225) );
  MUX2_X1 U3174 ( .A(n3225), .B(DATAI_11_), .S(n3651), .Z(n4413) );
  OAI22_X1 U3175 ( .A1(n4430), .A2(n2678), .B1(n4407), .B2(n2026), .ZN(n2463)
         );
  XNOR2_X1 U3176 ( .A(n2463), .B(n2729), .ZN(n2465) );
  OAI22_X1 U3177 ( .A1(n4430), .A2(n2731), .B1(n4407), .B2(n2678), .ZN(n2464)
         );
  OR2_X1 U3178 ( .A1(n2465), .A2(n2464), .ZN(n3407) );
  NAND2_X1 U3179 ( .A1(n2465), .A2(n2464), .ZN(n3406) );
  NAND2_X1 U3180 ( .A1(n2781), .A2(REG2_REG_13__SCAN_IN), .ZN(n2471) );
  INV_X1 U3181 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4500) );
  OR2_X1 U3182 ( .A1(n3652), .A2(n4500), .ZN(n2470) );
  INV_X1 U3183 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4391) );
  OR2_X1 U3184 ( .A1(n2360), .A2(n4391), .ZN(n2469) );
  NAND2_X1 U3185 ( .A1(n2486), .A2(n2466), .ZN(n2467) );
  NAND2_X1 U3186 ( .A1(n2508), .A2(n2467), .ZN(n4104) );
  OR2_X1 U3187 ( .A1(n2709), .A2(n4104), .ZN(n2468) );
  NAND4_X1 U3188 ( .A1(n2471), .A2(n2470), .A3(n2469), .A4(n2468), .ZN(n4395)
         );
  NAND2_X1 U3189 ( .A1(n4395), .A2(n2716), .ZN(n2477) );
  NOR2_X1 U3190 ( .A1(n2472), .A2(n2774), .ZN(n2473) );
  MUX2_X1 U3191 ( .A(n2774), .B(n2473), .S(IR_REG_13__SCAN_IN), .Z(n2475) );
  OR2_X1 U3192 ( .A1(n2475), .A2(n2474), .ZN(n3223) );
  MUX2_X1 U3193 ( .A(n3325), .B(DATAI_13_), .S(n3651), .Z(n3676) );
  NAND2_X1 U3194 ( .A1(n3676), .A2(n2711), .ZN(n2476) );
  NAND2_X1 U3195 ( .A1(n2477), .A2(n2476), .ZN(n2478) );
  XNOR2_X1 U3196 ( .A(n2478), .B(n2729), .ZN(n2502) );
  NAND2_X1 U3197 ( .A1(n4395), .A2(n2718), .ZN(n2480) );
  NAND2_X1 U3198 ( .A1(n3676), .A2(n2716), .ZN(n2479) );
  NAND2_X1 U3199 ( .A1(n2480), .A2(n2479), .ZN(n2503) );
  AND2_X1 U3200 ( .A1(n2502), .A2(n2503), .ZN(n2501) );
  NAND2_X1 U3201 ( .A1(n2781), .A2(REG2_REG_12__SCAN_IN), .ZN(n2490) );
  INV_X1 U3202 ( .A(REG0_REG_12__SCAN_IN), .ZN(n2481) );
  OR2_X1 U3203 ( .A1(n3652), .A2(n2481), .ZN(n2489) );
  INV_X1 U3204 ( .A(REG1_REG_12__SCAN_IN), .ZN(n2482) );
  OR2_X1 U3205 ( .A1(n2360), .A2(n2482), .ZN(n2488) );
  NAND2_X1 U3206 ( .A1(n2484), .A2(n2483), .ZN(n2485) );
  NAND2_X1 U3207 ( .A1(n2486), .A2(n2485), .ZN(n4276) );
  OR2_X1 U3208 ( .A1(n2564), .A2(n4276), .ZN(n2487) );
  NAND4_X1 U3209 ( .A1(n2490), .A2(n2489), .A3(n2488), .A4(n2487), .ZN(n4415)
         );
  NAND2_X1 U32100 ( .A1(n4415), .A2(n2716), .ZN(n2496) );
  INV_X1 U32110 ( .A(IR_REG_11__SCAN_IN), .ZN(n2491) );
  NAND2_X1 U32120 ( .A1(n2492), .A2(n2491), .ZN(n2493) );
  NAND2_X1 U32130 ( .A1(n2493), .A2(IR_REG_31__SCAN_IN), .ZN(n2494) );
  XNOR2_X1 U32140 ( .A(n2494), .B(IR_REG_12__SCAN_IN), .ZN(n4589) );
  MUX2_X1 U32150 ( .A(n4589), .B(DATAI_12_), .S(n3651), .Z(n4394) );
  NAND2_X1 U32160 ( .A1(n4394), .A2(n2711), .ZN(n2495) );
  NAND2_X1 U32170 ( .A1(n2496), .A2(n2495), .ZN(n2497) );
  XNOR2_X1 U32180 ( .A(n2497), .B(n2729), .ZN(n3543) );
  NAND2_X1 U32190 ( .A1(n4415), .A2(n2718), .ZN(n2499) );
  NAND2_X1 U32200 ( .A1(n4394), .A2(n2716), .ZN(n2498) );
  NAND2_X1 U32210 ( .A1(n2499), .A2(n2498), .ZN(n3542) );
  AND2_X1 U32220 ( .A1(n3543), .A2(n3542), .ZN(n2500) );
  INV_X1 U32230 ( .A(n2501), .ZN(n3541) );
  INV_X1 U32240 ( .A(n3542), .ZN(n3415) );
  INV_X1 U32250 ( .A(n3543), .ZN(n3545) );
  NAND3_X1 U32260 ( .A1(n3541), .A2(n3415), .A3(n3545), .ZN(n2506) );
  INV_X1 U32270 ( .A(n2502), .ZN(n2505) );
  INV_X1 U32280 ( .A(n2503), .ZN(n2504) );
  NAND2_X1 U32290 ( .A1(n2505), .A2(n2504), .ZN(n3540) );
  AND2_X1 U32300 ( .A1(n2506), .A2(n3540), .ZN(n2519) );
  NAND2_X1 U32310 ( .A1(n2781), .A2(REG2_REG_14__SCAN_IN), .ZN(n2513) );
  INV_X1 U32320 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4496) );
  OR2_X1 U32330 ( .A1(n3652), .A2(n4496), .ZN(n2512) );
  INV_X1 U32340 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4387) );
  OR2_X1 U32350 ( .A1(n2360), .A2(n4387), .ZN(n2511) );
  AND2_X1 U32360 ( .A1(n2508), .A2(n2507), .ZN(n2509) );
  OR2_X1 U32370 ( .A1(n2509), .A2(n2527), .ZN(n4093) );
  OR2_X1 U32380 ( .A1(n2564), .A2(n4093), .ZN(n2510) );
  NOR2_X1 U32390 ( .A1(n2474), .A2(n2774), .ZN(n2514) );
  MUX2_X1 U32400 ( .A(n2774), .B(n2514), .S(IR_REG_14__SCAN_IN), .Z(n2517) );
  INV_X1 U32410 ( .A(n2515), .ZN(n2516) );
  OAI22_X1 U32420 ( .A1(n4376), .A2(n2678), .B1(n2026), .B2(n4098), .ZN(n2518)
         );
  XNOR2_X1 U32430 ( .A(n2518), .B(n2714), .ZN(n3451) );
  OAI22_X1 U32440 ( .A1(n4376), .A2(n2731), .B1(n2678), .B2(n4098), .ZN(n3452)
         );
  AND2_X1 U32450 ( .A1(n2519), .A2(n3452), .ZN(n2520) );
  NAND2_X1 U32460 ( .A1(n2521), .A2(n2520), .ZN(n2524) );
  INV_X1 U32470 ( .A(n3452), .ZN(n2522) );
  OR2_X1 U32480 ( .A1(n2522), .A2(n3451), .ZN(n2523) );
  AND2_X1 U32490 ( .A1(n2524), .A2(n2523), .ZN(n2525) );
  NAND2_X1 U32500 ( .A1(n2781), .A2(REG2_REG_15__SCAN_IN), .ZN(n2532) );
  INV_X1 U32510 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4491) );
  OR2_X1 U32520 ( .A1(n3652), .A2(n4491), .ZN(n2531) );
  INV_X1 U32530 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4379) );
  OR2_X1 U32540 ( .A1(n2360), .A2(n4379), .ZN(n2530) );
  OR2_X1 U32550 ( .A1(n2527), .A2(REG3_REG_15__SCAN_IN), .ZN(n2528) );
  NAND2_X1 U32560 ( .A1(n2544), .A2(n2528), .ZN(n4074) );
  OR2_X1 U32570 ( .A1(n2564), .A2(n4074), .ZN(n2529) );
  NAND4_X1 U32580 ( .A1(n2532), .A2(n2531), .A3(n2530), .A4(n2529), .ZN(n4526)
         );
  NAND2_X1 U32590 ( .A1(n4526), .A2(n2716), .ZN(n2536) );
  NAND2_X1 U32600 ( .A1(n2515), .A2(IR_REG_31__SCAN_IN), .ZN(n2533) );
  NAND2_X1 U32610 ( .A1(n2533), .A2(n2247), .ZN(n2552) );
  OR2_X1 U32620 ( .A1(n2533), .A2(n2247), .ZN(n2534) );
  MUX2_X1 U32630 ( .A(n3339), .B(DATAI_15_), .S(n3651), .Z(n4372) );
  NAND2_X1 U32640 ( .A1(n4372), .A2(n2711), .ZN(n2535) );
  NAND2_X1 U32650 ( .A1(n2536), .A2(n2535), .ZN(n2537) );
  XNOR2_X1 U32660 ( .A(n2537), .B(n2714), .ZN(n2541) );
  NAND2_X1 U32670 ( .A1(n2540), .A2(n2541), .ZN(n3578) );
  NAND2_X1 U32680 ( .A1(n4526), .A2(n2718), .ZN(n2539) );
  NAND2_X1 U32690 ( .A1(n4372), .A2(n2710), .ZN(n2538) );
  NAND2_X1 U32700 ( .A1(n2539), .A2(n2538), .ZN(n4534) );
  NAND2_X1 U32710 ( .A1(n3578), .A2(n4534), .ZN(n2555) );
  INV_X1 U32720 ( .A(n2541), .ZN(n2542) );
  NAND2_X1 U32730 ( .A1(n2781), .A2(REG2_REG_16__SCAN_IN), .ZN(n2551) );
  NAND2_X1 U32740 ( .A1(n2544), .A2(n4528), .ZN(n2545) );
  INV_X1 U32750 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2546) );
  OR2_X1 U32760 ( .A1(n2360), .A2(n2546), .ZN(n2549) );
  INV_X1 U32770 ( .A(REG0_REG_16__SCAN_IN), .ZN(n2547) );
  OR2_X1 U32780 ( .A1(n3652), .A2(n2547), .ZN(n2548) );
  NAND2_X1 U32790 ( .A1(n2552), .A2(IR_REG_31__SCAN_IN), .ZN(n2553) );
  XNOR2_X1 U32800 ( .A(n2553), .B(IR_REG_16__SCAN_IN), .ZN(n3794) );
  MUX2_X1 U32810 ( .A(n3794), .B(DATAI_16_), .S(n3651), .Z(n4522) );
  OAI22_X1 U32820 ( .A1(n4363), .A2(n2678), .B1(n4050), .B2(n2026), .ZN(n2554)
         );
  XNOR2_X1 U32830 ( .A(n2554), .B(n2714), .ZN(n2556) );
  OAI22_X1 U32840 ( .A1(n4363), .A2(n2731), .B1(n4050), .B2(n2678), .ZN(n2557)
         );
  XNOR2_X1 U32850 ( .A(n2556), .B(n2557), .ZN(n4536) );
  NAND3_X1 U32860 ( .A1(n2555), .A2(n4533), .A3(n4536), .ZN(n2560) );
  INV_X1 U32870 ( .A(n2556), .ZN(n2558) );
  OR2_X1 U32880 ( .A1(n2558), .A2(n2557), .ZN(n2559) );
  NAND2_X1 U32890 ( .A1(n2781), .A2(REG2_REG_17__SCAN_IN), .ZN(n2568) );
  AND2_X1 U32900 ( .A1(n2562), .A2(n2561), .ZN(n2563) );
  OR2_X1 U32910 ( .A1(n2563), .A2(n2578), .ZN(n4030) );
  OR2_X1 U32920 ( .A1(n2564), .A2(n4030), .ZN(n2567) );
  INV_X1 U32930 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4366) );
  OR2_X1 U32940 ( .A1(n2360), .A2(n4366), .ZN(n2566) );
  INV_X1 U32950 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4483) );
  OR2_X1 U32960 ( .A1(n3652), .A2(n4483), .ZN(n2565) );
  NAND2_X1 U32970 ( .A1(n2062), .A2(IR_REG_31__SCAN_IN), .ZN(n2569) );
  XNOR2_X1 U32980 ( .A(n2569), .B(IR_REG_17__SCAN_IN), .ZN(n4699) );
  INV_X1 U32990 ( .A(n4699), .ZN(n4629) );
  INV_X1 U33000 ( .A(DATAI_17_), .ZN(n2570) );
  MUX2_X1 U33010 ( .A(n4629), .B(n2570), .S(n3651), .Z(n4034) );
  OAI22_X1 U33020 ( .A1(n4059), .A2(n2678), .B1(n4034), .B2(n2026), .ZN(n2571)
         );
  XNOR2_X1 U33030 ( .A(n2571), .B(n2714), .ZN(n3508) );
  OR2_X1 U33040 ( .A1(n4059), .A2(n2731), .ZN(n2573) );
  NAND2_X1 U33050 ( .A1(n4359), .A2(n2716), .ZN(n2572) );
  NAND2_X1 U33060 ( .A1(n2573), .A2(n2572), .ZN(n2575) );
  INV_X1 U33070 ( .A(n2575), .ZN(n3507) );
  AND2_X1 U33080 ( .A1(n3508), .A2(n3507), .ZN(n2574) );
  INV_X1 U33090 ( .A(n3508), .ZN(n2576) );
  NAND2_X1 U33100 ( .A1(n2576), .A2(n2575), .ZN(n2577) );
  NAND2_X1 U33110 ( .A1(n2781), .A2(REG2_REG_18__SCAN_IN), .ZN(n2583) );
  INV_X1 U33120 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4159) );
  OR2_X1 U33130 ( .A1(n3652), .A2(n4159), .ZN(n2582) );
  INV_X1 U33140 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3787) );
  OR2_X1 U33150 ( .A1(n2360), .A2(n3787), .ZN(n2581) );
  NOR2_X1 U33160 ( .A1(n2578), .A2(REG3_REG_18__SCAN_IN), .ZN(n2579) );
  OR2_X1 U33170 ( .A1(n2607), .A2(n2579), .ZN(n4019) );
  OR2_X1 U33180 ( .A1(n2709), .A2(n4019), .ZN(n2580) );
  NOR2_X1 U33190 ( .A1(n2584), .A2(n2774), .ZN(n2585) );
  MUX2_X1 U33200 ( .A(n2774), .B(n2585), .S(IR_REG_18__SCAN_IN), .Z(n2586) );
  INV_X1 U33210 ( .A(n2586), .ZN(n2587) );
  AND2_X1 U33220 ( .A1(n2587), .A2(n2283), .ZN(n3797) );
  MUX2_X1 U33230 ( .A(n3797), .B(DATAI_18_), .S(n3651), .Z(n4009) );
  OAI22_X1 U33240 ( .A1(n3997), .A2(n2678), .B1(n4016), .B2(n2026), .ZN(n2588)
         );
  XNOR2_X1 U33250 ( .A(n2588), .B(n2729), .ZN(n2590) );
  OAI22_X1 U33260 ( .A1(n3997), .A2(n2731), .B1(n4016), .B2(n2678), .ZN(n2589)
         );
  AND2_X1 U33270 ( .A1(n2590), .A2(n2589), .ZN(n3422) );
  NAND2_X1 U33280 ( .A1(n2781), .A2(REG2_REG_19__SCAN_IN), .ZN(n2594) );
  INV_X1 U33290 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4479) );
  OR2_X1 U33300 ( .A1(n3652), .A2(n4479), .ZN(n2593) );
  INV_X1 U33310 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4354) );
  OR2_X1 U33320 ( .A1(n2360), .A2(n4354), .ZN(n2592) );
  XNOR2_X1 U33330 ( .A(n2607), .B(REG3_REG_19__SCAN_IN), .ZN(n3999) );
  OR2_X1 U33340 ( .A1(n2709), .A2(n3999), .ZN(n2591) );
  NAND4_X1 U33350 ( .A1(n2594), .A2(n2593), .A3(n2592), .A4(n2591), .ZN(n4010)
         );
  NAND2_X1 U33360 ( .A1(n4010), .A2(n2716), .ZN(n2596) );
  MUX2_X1 U33370 ( .A(n3732), .B(DATAI_19_), .S(n3651), .Z(n3993) );
  NAND2_X1 U33380 ( .A1(n3993), .A2(n2711), .ZN(n2595) );
  NAND2_X1 U33390 ( .A1(n2596), .A2(n2595), .ZN(n2597) );
  XNOR2_X1 U33400 ( .A(n2597), .B(n2729), .ZN(n2598) );
  AOI22_X1 U33410 ( .A1(n4010), .A2(n2718), .B1(n2716), .B2(n3993), .ZN(n2599)
         );
  XNOR2_X1 U33420 ( .A(n2598), .B(n2599), .ZN(n3481) );
  NAND2_X1 U33430 ( .A1(n3480), .A2(n3481), .ZN(n2602) );
  INV_X1 U33440 ( .A(n2598), .ZN(n2600) );
  NAND2_X1 U33450 ( .A1(n2600), .A2(n2599), .ZN(n2601) );
  NAND2_X1 U33460 ( .A1(n2602), .A2(n2601), .ZN(n3529) );
  NAND2_X1 U33470 ( .A1(n2781), .A2(REG2_REG_20__SCAN_IN), .ZN(n2612) );
  INV_X1 U33480 ( .A(REG0_REG_20__SCAN_IN), .ZN(n2603) );
  OR2_X1 U33490 ( .A1(n3652), .A2(n2603), .ZN(n2611) );
  INV_X1 U33500 ( .A(REG1_REG_20__SCAN_IN), .ZN(n2604) );
  OR2_X1 U33510 ( .A1(n2360), .A2(n2604), .ZN(n2610) );
  NAND2_X1 U33520 ( .A1(n2607), .A2(REG3_REG_19__SCAN_IN), .ZN(n2605) );
  INV_X1 U3353 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3534) );
  NAND2_X1 U33540 ( .A1(n2605), .A2(n3534), .ZN(n2608) );
  AND2_X1 U3355 ( .A1(REG3_REG_19__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2606) );
  NAND2_X1 U3356 ( .A1(n2607), .A2(n2606), .ZN(n2622) );
  NAND2_X1 U3357 ( .A1(n2608), .A2(n2622), .ZN(n3978) );
  OR2_X1 U3358 ( .A1(n2709), .A2(n3978), .ZN(n2609) );
  NAND4_X1 U3359 ( .A1(n2612), .A2(n2611), .A3(n2610), .A4(n2609), .ZN(n3994)
         );
  NAND2_X1 U3360 ( .A1(n3994), .A2(n2716), .ZN(n2614) );
  NAND2_X1 U3361 ( .A1(n2711), .A2(n3977), .ZN(n2613) );
  NAND2_X1 U3362 ( .A1(n2614), .A2(n2613), .ZN(n2615) );
  XNOR2_X1 U3363 ( .A(n2615), .B(n2729), .ZN(n2618) );
  NAND2_X1 U3364 ( .A1(n3994), .A2(n2718), .ZN(n2617) );
  NAND2_X1 U3365 ( .A1(n2716), .A2(n3977), .ZN(n2616) );
  NAND2_X1 U3366 ( .A1(n2617), .A2(n2616), .ZN(n2619) );
  NAND2_X1 U3367 ( .A1(n2618), .A2(n2619), .ZN(n3530) );
  INV_X1 U3368 ( .A(n2618), .ZN(n2621) );
  INV_X1 U3369 ( .A(n2619), .ZN(n2620) );
  NAND2_X1 U3370 ( .A1(n2621), .A2(n2620), .ZN(n3532) );
  NAND2_X1 U3371 ( .A1(n2781), .A2(REG2_REG_21__SCAN_IN), .ZN(n2627) );
  INV_X1 U3372 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4474) );
  OR2_X1 U3373 ( .A1(n3652), .A2(n4474), .ZN(n2626) );
  INV_X1 U3374 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4343) );
  OR2_X1 U3375 ( .A1(n2360), .A2(n4343), .ZN(n2625) );
  NAND2_X1 U3376 ( .A1(n2622), .A2(n3492), .ZN(n2623) );
  NAND2_X1 U3377 ( .A1(n2634), .A2(n2623), .ZN(n3491) );
  OR2_X1 U3378 ( .A1(n2564), .A2(n3491), .ZN(n2624) );
  INV_X1 U3379 ( .A(n4336), .ZN(n3961) );
  OAI22_X1 U3380 ( .A1(n3935), .A2(n2318), .B1(n3961), .B2(n2026), .ZN(n2628)
         );
  XNOR2_X1 U3381 ( .A(n2628), .B(n2714), .ZN(n3488) );
  OR2_X1 U3382 ( .A1(n3935), .A2(n2731), .ZN(n2630) );
  NAND2_X1 U3383 ( .A1(n2710), .A2(n4336), .ZN(n2629) );
  NAND2_X1 U3384 ( .A1(n2630), .A2(n2629), .ZN(n2632) );
  INV_X1 U3385 ( .A(n2632), .ZN(n3487) );
  AND2_X1 U3386 ( .A1(n3488), .A2(n3487), .ZN(n2631) );
  INV_X1 U3387 ( .A(n3488), .ZN(n2633) );
  AND2_X1 U3388 ( .A1(n2634), .A2(n3558), .ZN(n2635) );
  OR2_X1 U3389 ( .A1(n2635), .A2(n2644), .ZN(n3948) );
  INV_X1 U3390 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4470) );
  OR2_X1 U3391 ( .A1(n3652), .A2(n4470), .ZN(n2637) );
  INV_X1 U3392 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4334) );
  OR2_X1 U3393 ( .A1(n2360), .A2(n4334), .ZN(n2636) );
  AND2_X1 U3394 ( .A1(n2637), .A2(n2636), .ZN(n2639) );
  NAND2_X1 U3395 ( .A1(n2781), .A2(REG2_REG_22__SCAN_IN), .ZN(n2638) );
  NAND2_X1 U3396 ( .A1(n4337), .A2(n2716), .ZN(n2641) );
  NAND2_X1 U3397 ( .A1(n2711), .A2(n3945), .ZN(n2640) );
  NAND2_X1 U3398 ( .A1(n2641), .A2(n2640), .ZN(n2642) );
  XNOR2_X1 U3399 ( .A(n2642), .B(n2714), .ZN(n2653) );
  AND2_X1 U3400 ( .A1(n3945), .A2(n2716), .ZN(n2643) );
  AOI21_X1 U3401 ( .B1(n4337), .B2(n2718), .A(n2643), .ZN(n2652) );
  XNOR2_X1 U3402 ( .A(n2653), .B(n2652), .ZN(n3557) );
  OR2_X2 U3403 ( .A1(n3556), .A2(n3557), .ZN(n3554) );
  NOR2_X1 U3404 ( .A1(n2644), .A2(REG3_REG_23__SCAN_IN), .ZN(n2645) );
  OR2_X1 U3405 ( .A1(n2654), .A2(n2645), .ZN(n3925) );
  AOI22_X1 U3406 ( .A1(n2141), .A2(REG0_REG_23__SCAN_IN), .B1(n2304), .B2(
        REG1_REG_23__SCAN_IN), .ZN(n2647) );
  NAND2_X1 U3407 ( .A1(n2781), .A2(REG2_REG_23__SCAN_IN), .ZN(n2646) );
  OAI211_X1 U3408 ( .C1(n3925), .C2(n2709), .A(n2647), .B(n2646), .ZN(n4320)
         );
  NAND2_X1 U3409 ( .A1(n4320), .A2(n2716), .ZN(n2649) );
  NAND2_X1 U3410 ( .A1(n3922), .A2(n2711), .ZN(n2648) );
  NAND2_X1 U3411 ( .A1(n2649), .A2(n2648), .ZN(n2650) );
  XNOR2_X1 U3412 ( .A(n2650), .B(n2729), .ZN(n2663) );
  NOR2_X1 U3413 ( .A1(n3917), .A2(n2678), .ZN(n2651) );
  AOI21_X1 U3414 ( .B1(n4320), .B2(n2718), .A(n2651), .ZN(n2661) );
  XNOR2_X1 U3415 ( .A(n2663), .B(n2661), .ZN(n3462) );
  NAND2_X1 U3416 ( .A1(n2653), .A2(n2652), .ZN(n3463) );
  NAND2_X1 U3417 ( .A1(n2654), .A2(REG3_REG_24__SCAN_IN), .ZN(n2672) );
  OR2_X1 U3418 ( .A1(n2654), .A2(REG3_REG_24__SCAN_IN), .ZN(n2655) );
  NAND2_X1 U3419 ( .A1(n2672), .A2(n2655), .ZN(n3521) );
  INV_X1 U3420 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4462) );
  INV_X1 U3421 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4326) );
  OAI22_X1 U3422 ( .A1(n3652), .A2(n4462), .B1(n2360), .B2(n4326), .ZN(n2656)
         );
  INV_X1 U3423 ( .A(n2656), .ZN(n2658) );
  NAND2_X1 U3424 ( .A1(n2781), .A2(REG2_REG_24__SCAN_IN), .ZN(n2657) );
  NOR2_X1 U3425 ( .A1(n3904), .A2(n2678), .ZN(n2659) );
  AOI21_X1 U3426 ( .B1(n3880), .B2(n2718), .A(n2659), .ZN(n2668) );
  INV_X1 U3427 ( .A(n2668), .ZN(n2660) );
  AND2_X1 U3428 ( .A1(n3461), .A2(n2660), .ZN(n2664) );
  INV_X1 U3429 ( .A(n2661), .ZN(n2662) );
  NAND2_X1 U3430 ( .A1(n2663), .A2(n2662), .ZN(n2669) );
  NAND2_X1 U3431 ( .A1(n3880), .A2(n2710), .ZN(n2666) );
  INV_X1 U3432 ( .A(n3904), .ZN(n4319) );
  NAND2_X1 U3433 ( .A1(n4319), .A2(n2711), .ZN(n2665) );
  NAND2_X1 U3434 ( .A1(n2666), .A2(n2665), .ZN(n2667) );
  XNOR2_X1 U3435 ( .A(n2667), .B(n2729), .ZN(n3520) );
  AND2_X1 U3436 ( .A1(n3461), .A2(n3520), .ZN(n2671) );
  INV_X1 U3437 ( .A(n3520), .ZN(n2670) );
  AND2_X1 U3438 ( .A1(n2669), .A2(n2668), .ZN(n3516) );
  INV_X1 U3439 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3501) );
  NAND2_X1 U3440 ( .A1(n2672), .A2(n3501), .ZN(n2673) );
  NAND2_X1 U3441 ( .A1(n2683), .A2(n2673), .ZN(n3887) );
  OR2_X1 U3442 ( .A1(n3887), .A2(n2564), .ZN(n2676) );
  AOI22_X1 U3443 ( .A1(n2304), .A2(REG1_REG_25__SCAN_IN), .B1(n2781), .B2(
        REG2_REG_25__SCAN_IN), .ZN(n2675) );
  INV_X1 U3444 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4458) );
  OR2_X1 U3445 ( .A1(n3652), .A2(n4458), .ZN(n2674) );
  OAI22_X1 U3446 ( .A1(n4323), .A2(n2318), .B1(n3885), .B2(n2026), .ZN(n2677)
         );
  XNOR2_X1 U3447 ( .A(n2677), .B(n2714), .ZN(n2680) );
  OAI22_X1 U3448 ( .A1(n4323), .A2(n2731), .B1(n3885), .B2(n2678), .ZN(n2681)
         );
  INV_X1 U3449 ( .A(n2681), .ZN(n2679) );
  NAND2_X1 U3450 ( .A1(n2680), .A2(n2679), .ZN(n3497) );
  INV_X1 U3451 ( .A(n2680), .ZN(n2682) );
  NAND2_X1 U3452 ( .A1(n2682), .A2(n2681), .ZN(n3498) );
  INV_X1 U3453 ( .A(n3568), .ZN(n2697) );
  INV_X1 U3454 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3571) );
  NAND2_X1 U3455 ( .A1(n2683), .A2(n3571), .ZN(n2684) );
  NAND2_X1 U3456 ( .A1(n3871), .A2(n2685), .ZN(n2690) );
  INV_X1 U3457 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4454) );
  NAND2_X1 U34580 ( .A1(n4742), .A2(REG2_REG_26__SCAN_IN), .ZN(n2687) );
  INV_X1 U34590 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4313) );
  OR2_X1 U3460 ( .A1(n2360), .A2(n4313), .ZN(n2686) );
  OAI211_X1 U3461 ( .C1(n3652), .C2(n4454), .A(n2687), .B(n2686), .ZN(n2688)
         );
  INV_X1 U3462 ( .A(n2688), .ZN(n2689) );
  NAND2_X1 U3463 ( .A1(n4303), .A2(n2710), .ZN(n2692) );
  NAND2_X1 U3464 ( .A1(n3651), .A2(DATAI_26_), .ZN(n3869) );
  NAND2_X1 U3465 ( .A1(n3863), .A2(n2711), .ZN(n2691) );
  NAND2_X1 U3466 ( .A1(n2692), .A2(n2691), .ZN(n2693) );
  XNOR2_X1 U34670 ( .A(n2693), .B(n2729), .ZN(n2698) );
  NAND2_X1 U3468 ( .A1(n4303), .A2(n2718), .ZN(n2695) );
  NAND2_X1 U34690 ( .A1(n3863), .A2(n2710), .ZN(n2694) );
  NAND2_X1 U3470 ( .A1(n2695), .A2(n2694), .ZN(n2699) );
  AND2_X1 U34710 ( .A1(n2698), .A2(n2699), .ZN(n3565) );
  INV_X1 U3472 ( .A(n3565), .ZN(n2696) );
  INV_X1 U34730 ( .A(n2698), .ZN(n2701) );
  INV_X1 U3474 ( .A(n2699), .ZN(n2700) );
  NAND2_X1 U34750 ( .A1(n2701), .A2(n2700), .ZN(n3564) );
  INV_X1 U3476 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3432) );
  AND2_X1 U34770 ( .A1(n2703), .A2(n3432), .ZN(n2704) );
  INV_X1 U3478 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4450) );
  NAND2_X1 U34790 ( .A1(n2781), .A2(REG2_REG_27__SCAN_IN), .ZN(n2706) );
  INV_X1 U3480 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4309) );
  OR2_X1 U34810 ( .A1(n2360), .A2(n4309), .ZN(n2705) );
  OAI211_X1 U3482 ( .C1(n3652), .C2(n4450), .A(n2706), .B(n2705), .ZN(n2707)
         );
  INV_X1 U34830 ( .A(n2707), .ZN(n2708) );
  OAI21_X1 U3484 ( .B1(n3431), .B2(n2709), .A(n2708), .ZN(n3828) );
  NAND2_X1 U34850 ( .A1(n3828), .A2(n2710), .ZN(n2713) );
  NAND2_X1 U3486 ( .A1(n2711), .A2(n4302), .ZN(n2712) );
  NAND2_X1 U34870 ( .A1(n2713), .A2(n2712), .ZN(n2715) );
  XNOR2_X1 U3488 ( .A(n2715), .B(n2714), .ZN(n2755) );
  AND2_X1 U34890 ( .A1(n4302), .A2(n2716), .ZN(n2717) );
  AOI21_X1 U3490 ( .B1(n3828), .B2(n2718), .A(n2717), .ZN(n2756) );
  XNOR2_X1 U34910 ( .A(n2755), .B(n2756), .ZN(n3429) );
  NAND2_X1 U3492 ( .A1(n2719), .A2(REG3_REG_28__SCAN_IN), .ZN(n3819) );
  INV_X1 U34930 ( .A(n2719), .ZN(n2721) );
  INV_X1 U3494 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2720) );
  NAND2_X1 U34950 ( .A1(n2721), .A2(n2720), .ZN(n2722) );
  NAND2_X1 U3496 ( .A1(n3819), .A2(n2722), .ZN(n3829) );
  INV_X1 U34970 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4208) );
  NAND2_X1 U3498 ( .A1(n4742), .A2(REG2_REG_28__SCAN_IN), .ZN(n2724) );
  INV_X1 U34990 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4222) );
  OR2_X1 U3500 ( .A1(n2360), .A2(n4222), .ZN(n2723) );
  OAI211_X1 U35010 ( .C1(n3652), .C2(n4208), .A(n2724), .B(n2723), .ZN(n2725)
         );
  INV_X1 U3502 ( .A(n2725), .ZN(n2726) );
  OAI22_X1 U35030 ( .A1(n4305), .A2(n2318), .B1(n3833), .B2(n2026), .ZN(n2730)
         );
  XNOR2_X1 U3504 ( .A(n2730), .B(n2729), .ZN(n2733) );
  OAI22_X1 U35050 ( .A1(n4305), .A2(n2731), .B1(n3833), .B2(n2318), .ZN(n2732)
         );
  XNOR2_X1 U35060 ( .A(n2733), .B(n2732), .ZN(n2792) );
  INV_X1 U35070 ( .A(n2792), .ZN(n2759) );
  NAND2_X1 U35080 ( .A1(n2734), .A2(n2949), .ZN(n2735) );
  MUX2_X1 U35090 ( .A(n2734), .B(n2735), .S(B_REG_SCAN_IN), .Z(n2736) );
  OAI22_X1 U35100 ( .A1(n2948), .A2(D_REG_1__SCAN_IN), .B1(n2931), .B2(n2934), 
        .ZN(n2887) );
  INV_X1 U35110 ( .A(n2887), .ZN(n3062) );
  INV_X1 U35120 ( .A(D_REG_0__SCAN_IN), .ZN(n2738) );
  INV_X1 U35130 ( .A(n2931), .ZN(n2952) );
  NOR4_X1 U35140 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2747) );
  NOR4_X1 U35150 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2746) );
  INV_X1 U35160 ( .A(D_REG_25__SCAN_IN), .ZN(n4670) );
  INV_X1 U35170 ( .A(D_REG_11__SCAN_IN), .ZN(n4684) );
  INV_X1 U35180 ( .A(D_REG_15__SCAN_IN), .ZN(n4680) );
  INV_X1 U35190 ( .A(D_REG_3__SCAN_IN), .ZN(n4692) );
  NAND4_X1 U35200 ( .A1(n4670), .A2(n4684), .A3(n4680), .A4(n4692), .ZN(n2744)
         );
  NOR4_X1 U35210 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2742) );
  NOR4_X1 U35220 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2741) );
  NOR4_X1 U35230 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2740) );
  NOR4_X1 U35240 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2739) );
  NAND4_X1 U35250 ( .A1(n2742), .A2(n2741), .A3(n2740), .A4(n2739), .ZN(n2743)
         );
  NOR4_X1 U35260 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(n2744), 
        .A4(n2743), .ZN(n2745) );
  NAND3_X1 U35270 ( .A1(n2747), .A2(n2746), .A3(n2745), .ZN(n2748) );
  NAND2_X1 U35280 ( .A1(n2749), .A2(n2748), .ZN(n3060) );
  NAND3_X1 U35290 ( .A1(n3062), .A2(n2892), .A3(n3060), .ZN(n2773) );
  AND2_X1 U35300 ( .A1(n2778), .A2(n3802), .ZN(n2765) );
  INV_X1 U35310 ( .A(n2765), .ZN(n2752) );
  NAND2_X1 U35320 ( .A1(n3065), .A2(n2752), .ZN(n2753) );
  NAND2_X1 U35330 ( .A1(n3736), .A2(n3727), .ZN(n2839) );
  NAND2_X1 U35340 ( .A1(n2753), .A2(n2839), .ZN(n2754) );
  INV_X1 U35350 ( .A(n2755), .ZN(n2758) );
  INV_X1 U35360 ( .A(n2756), .ZN(n2757) );
  NAND2_X1 U35370 ( .A1(n2758), .A2(n2757), .ZN(n2761) );
  NAND3_X1 U35380 ( .A1(n2759), .A2(n4538), .A3(n2761), .ZN(n2795) );
  AND2_X1 U35390 ( .A1(n2792), .A2(n4538), .ZN(n2760) );
  NAND2_X1 U35400 ( .A1(n2796), .A2(n2760), .ZN(n2794) );
  NOR2_X1 U35410 ( .A1(n2761), .A2(n3584), .ZN(n2791) );
  AND2_X1 U35420 ( .A1(n2778), .A2(n3732), .ZN(n2762) );
  NAND2_X1 U35430 ( .A1(n2773), .A2(n2779), .ZN(n3056) );
  NOR2_X1 U35440 ( .A1(n2839), .A2(n2765), .ZN(n2884) );
  INV_X1 U35450 ( .A(n2944), .ZN(n2766) );
  NOR2_X1 U35460 ( .A1(n2884), .A2(n2766), .ZN(n2767) );
  AND2_X1 U35470 ( .A1(n2294), .A2(n2767), .ZN(n2768) );
  NAND2_X1 U35480 ( .A1(n3056), .A2(n2768), .ZN(n2769) );
  INV_X1 U35490 ( .A(n2770), .ZN(n2771) );
  NAND2_X1 U35500 ( .A1(n4695), .A2(n2771), .ZN(n2772) );
  NOR2_X1 U35510 ( .A1(n2775), .A2(n2774), .ZN(n2776) );
  INV_X1 U35520 ( .A(n2778), .ZN(n4514) );
  AOI22_X1 U35530 ( .A1(n3828), .A2(n4527), .B1(n2898), .B2(n3569), .ZN(n2789)
         );
  OR2_X1 U35540 ( .A1(n3819), .A2(n2564), .ZN(n2786) );
  INV_X1 U35550 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2909) );
  NAND2_X1 U35560 ( .A1(n2141), .A2(REG0_REG_29__SCAN_IN), .ZN(n2783) );
  NAND2_X1 U35570 ( .A1(n2781), .A2(REG2_REG_29__SCAN_IN), .ZN(n2782) );
  OAI211_X1 U35580 ( .C1(n2909), .C2(n2360), .A(n2783), .B(n2782), .ZN(n2784)
         );
  INV_X1 U35590 ( .A(n2784), .ZN(n2785) );
  NAND2_X1 U35600 ( .A1(n2786), .A2(n2785), .ZN(n3827) );
  AOI22_X1 U35610 ( .A1(n3827), .A2(n3570), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n2788) );
  OAI211_X1 U35620 ( .C1(n3829), .C2(n4543), .A(n2789), .B(n2788), .ZN(n2790)
         );
  AOI21_X1 U35630 ( .B1(n2792), .B2(n2791), .A(n2790), .ZN(n2793) );
  OAI211_X1 U35640 ( .C1(n2796), .C2(n2795), .A(n2794), .B(n2793), .ZN(U3217)
         );
  INV_X1 U35650 ( .A(n3880), .ZN(n3918) );
  NAND2_X1 U35660 ( .A1(n2797), .A2(n3126), .ZN(n3589) );
  AND2_X1 U35670 ( .A1(n3748), .A2(n3093), .ZN(n3075) );
  NAND2_X1 U35680 ( .A1(n2842), .A2(n3075), .ZN(n3077) );
  NAND2_X1 U35690 ( .A1(n2799), .A2(n3126), .ZN(n2800) );
  NAND2_X1 U35700 ( .A1(n3077), .A2(n2800), .ZN(n3107) );
  INV_X1 U35710 ( .A(n3107), .ZN(n2801) );
  NAND2_X1 U35720 ( .A1(n3746), .A2(n3137), .ZN(n3593) );
  NAND2_X1 U35730 ( .A1(n3084), .A2(n3152), .ZN(n3590) );
  NAND2_X1 U35740 ( .A1(n2802), .A2(n3258), .ZN(n3596) );
  NAND2_X1 U35750 ( .A1(n3084), .A2(n3137), .ZN(n3144) );
  AND2_X1 U35760 ( .A1(n3144), .A2(n2803), .ZN(n3251) );
  NAND2_X1 U35770 ( .A1(n3105), .A2(n2805), .ZN(n3255) );
  NAND2_X1 U35780 ( .A1(n2806), .A2(n3258), .ZN(n2807) );
  NAND2_X1 U35790 ( .A1(n3745), .A2(n3475), .ZN(n3252) );
  NAND2_X1 U35800 ( .A1(n3255), .A2(n2808), .ZN(n3174) );
  NAND2_X1 U35810 ( .A1(n3276), .A2(n2846), .ZN(n2809) );
  NAND2_X1 U3582 ( .A1(n3174), .A2(n2809), .ZN(n2811) );
  NAND2_X1 U3583 ( .A1(n3744), .A2(n3242), .ZN(n2810) );
  NAND2_X1 U3584 ( .A1(n2811), .A2(n2810), .ZN(n3272) );
  NAND2_X1 U3585 ( .A1(n2812), .A2(n3442), .ZN(n2848) );
  INV_X2 U3586 ( .A(n2812), .ZN(n3742) );
  NAND2_X1 U3587 ( .A1(n3742), .A2(n3293), .ZN(n3612) );
  NAND2_X1 U3588 ( .A1(n3441), .A2(n3361), .ZN(n2813) );
  NAND2_X1 U3589 ( .A1(n2814), .A2(n2813), .ZN(n3314) );
  AND2_X1 U3590 ( .A1(n4433), .A2(n3395), .ZN(n2815) );
  INV_X1 U3591 ( .A(n4433), .ZN(n3363) );
  INV_X1 U3592 ( .A(n3395), .ZN(n2851) );
  NAND2_X1 U3593 ( .A1(n3363), .A2(n2851), .ZN(n2816) );
  INV_X1 U3594 ( .A(n4416), .ZN(n3318) );
  INV_X1 U3595 ( .A(n3387), .ZN(n4427) );
  NAND2_X1 U3596 ( .A1(n4430), .A2(n4413), .ZN(n4105) );
  NAND2_X1 U3597 ( .A1(n4281), .A2(n4407), .ZN(n4107) );
  INV_X1 U3598 ( .A(n4415), .ZN(n2854) );
  NAND2_X1 U3599 ( .A1(n2854), .A2(n4273), .ZN(n2818) );
  NAND2_X1 U3600 ( .A1(n2819), .A2(n2818), .ZN(n4118) );
  NAND2_X1 U3601 ( .A1(n4376), .A2(n4381), .ZN(n4065) );
  NAND2_X1 U3602 ( .A1(n4073), .A2(n4098), .ZN(n3608) );
  NAND2_X1 U3603 ( .A1(n4065), .A2(n3608), .ZN(n4088) );
  NAND2_X1 U3604 ( .A1(n4373), .A2(n4522), .ZN(n2821) );
  NAND2_X1 U3605 ( .A1(n4363), .A2(n4522), .ZN(n3699) );
  NAND2_X1 U3606 ( .A1(n4373), .A2(n4050), .ZN(n3701) );
  INV_X1 U3607 ( .A(n4526), .ZN(n2861) );
  NAND2_X1 U3608 ( .A1(n2861), .A2(n4078), .ZN(n4044) );
  NAND2_X1 U3609 ( .A1(n4526), .A2(n4372), .ZN(n4043) );
  OR2_X1 U3610 ( .A1(n2820), .A2(n4043), .ZN(n4040) );
  AND2_X1 U3611 ( .A1(n2821), .A2(n4040), .ZN(n2822) );
  AND2_X1 U3612 ( .A1(n4088), .A2(n2822), .ZN(n2825) );
  INV_X1 U3613 ( .A(n2822), .ZN(n2824) );
  NAND2_X1 U3614 ( .A1(n4376), .A2(n4098), .ZN(n4042) );
  AND2_X1 U3615 ( .A1(n4042), .A2(n2823), .ZN(n4039) );
  NAND2_X1 U3616 ( .A1(n4059), .A2(n4034), .ZN(n2826) );
  NAND2_X1 U3617 ( .A1(n3997), .A2(n4009), .ZN(n3987) );
  NAND2_X1 U3618 ( .A1(n4360), .A2(n4016), .ZN(n3988) );
  NAND2_X1 U3619 ( .A1(n3987), .A2(n3988), .ZN(n4008) );
  NAND2_X1 U3620 ( .A1(n3997), .A2(n4016), .ZN(n2827) );
  NAND2_X1 U3621 ( .A1(n4004), .A2(n2827), .ZN(n3984) );
  NAND2_X1 U3622 ( .A1(n4010), .A2(n3993), .ZN(n2829) );
  NOR2_X1 U3623 ( .A1(n4010), .A2(n3993), .ZN(n2828) );
  AND2_X1 U3624 ( .A1(n3994), .A2(n3977), .ZN(n3668) );
  INV_X1 U3625 ( .A(n3935), .ZN(n3969) );
  AND2_X1 U3626 ( .A1(n3969), .A2(n4336), .ZN(n3940) );
  INV_X1 U3627 ( .A(n3940), .ZN(n2833) );
  INV_X1 U3628 ( .A(n3994), .ZN(n4340) );
  NAND2_X1 U3629 ( .A1(n4340), .A2(n2889), .ZN(n3936) );
  INV_X1 U3630 ( .A(n4337), .ZN(n2830) );
  NAND2_X1 U3631 ( .A1(n2830), .A2(n3945), .ZN(n3914) );
  INV_X1 U3632 ( .A(n3945), .ZN(n2831) );
  NAND2_X1 U3633 ( .A1(n4337), .A2(n2831), .ZN(n2872) );
  NAND2_X1 U3634 ( .A1(n3914), .A2(n2872), .ZN(n3941) );
  NAND2_X1 U3635 ( .A1(n3935), .A2(n3961), .ZN(n3939) );
  OAI211_X1 U3636 ( .C1(n3940), .C2(n3936), .A(n3941), .B(n3939), .ZN(n2832)
         );
  NOR2_X1 U3637 ( .A1(n4320), .A2(n3922), .ZN(n2834) );
  INV_X1 U3638 ( .A(n4320), .ZN(n3523) );
  NAND2_X1 U3639 ( .A1(n4323), .A2(n3885), .ZN(n2835) );
  NAND2_X1 U3640 ( .A1(n4303), .A2(n3863), .ZN(n3679) );
  INV_X1 U3641 ( .A(n4303), .ZN(n3433) );
  NAND2_X1 U3642 ( .A1(n3433), .A2(n3869), .ZN(n3680) );
  NOR2_X1 U3643 ( .A1(n3828), .A2(n4302), .ZN(n2836) );
  INV_X1 U3644 ( .A(n3828), .ZN(n3866) );
  NAND2_X1 U3645 ( .A1(n3848), .A2(n3833), .ZN(n3642) );
  NAND2_X1 U3646 ( .A1(n4305), .A2(n2898), .ZN(n3650) );
  NAND2_X1 U3647 ( .A1(n3642), .A2(n3650), .ZN(n3693) );
  XNOR2_X1 U3648 ( .A(n2837), .B(n3736), .ZN(n2838) );
  INV_X1 U3649 ( .A(n4726), .ZN(n4437) );
  NOR2_X2 U3650 ( .A1(n4521), .A2(n2839), .ZN(n4434) );
  INV_X1 U3651 ( .A(n3827), .ZN(n2840) );
  INV_X1 U3652 ( .A(n2839), .ZN(n2942) );
  OAI22_X1 U3653 ( .A1(n2840), .A2(n4429), .B1(n4428), .B2(n3833), .ZN(n2841)
         );
  AOI21_X1 U3654 ( .B1(n4434), .B2(n3828), .A(n2841), .ZN(n2883) );
  INV_X1 U3655 ( .A(n3748), .ZN(n2843) );
  NAND2_X1 U3656 ( .A1(n2843), .A2(n3093), .ZN(n3078) );
  NAND2_X1 U3657 ( .A1(n3079), .A2(n3589), .ZN(n3110) );
  NAND2_X1 U3658 ( .A1(n3110), .A2(n3684), .ZN(n3109) );
  NAND2_X1 U3659 ( .A1(n3109), .A2(n3590), .ZN(n3147) );
  NAND2_X1 U3660 ( .A1(n3193), .A2(n3475), .ZN(n3595) );
  NAND2_X1 U3661 ( .A1(n3745), .A2(n3200), .ZN(n3592) );
  AND2_X1 U3662 ( .A1(n3595), .A2(n3592), .ZN(n3148) );
  INV_X1 U3663 ( .A(n3596), .ZN(n2845) );
  AND2_X1 U3664 ( .A1(n3744), .A2(n2846), .ZN(n3171) );
  NAND2_X1 U3665 ( .A1(n3276), .A2(n3242), .ZN(n3613) );
  INV_X1 U3666 ( .A(n3274), .ZN(n3281) );
  NAND2_X1 U3667 ( .A1(n3743), .A2(n3281), .ZN(n3615) );
  NAND2_X1 U3668 ( .A1(n3273), .A2(n3615), .ZN(n2847) );
  INV_X1 U3669 ( .A(n3743), .ZN(n3445) );
  NAND2_X1 U3670 ( .A1(n3445), .A2(n3274), .ZN(n3601) );
  INV_X1 U3671 ( .A(n2848), .ZN(n2849) );
  NAND2_X1 U3672 ( .A1(n3398), .A2(n3361), .ZN(n3605) );
  NAND2_X1 U3673 ( .A1(n3441), .A2(n3357), .ZN(n3616) );
  AND2_X1 U3674 ( .A1(n4433), .A2(n2851), .ZN(n3610) );
  NAND2_X1 U3675 ( .A1(n3363), .A2(n3395), .ZN(n3606) );
  NAND2_X1 U3676 ( .A1(n4416), .A2(n4427), .ZN(n3623) );
  NAND2_X1 U3677 ( .A1(n3318), .A2(n3387), .ZN(n3621) );
  NAND2_X1 U3678 ( .A1(n4415), .A2(n4273), .ZN(n4109) );
  INV_X1 U3679 ( .A(n3676), .ZN(n4121) );
  NAND2_X1 U3680 ( .A1(n4395), .A2(n4121), .ZN(n2852) );
  NAND2_X1 U3681 ( .A1(n4109), .A2(n2852), .ZN(n2855) );
  INV_X1 U3682 ( .A(n4107), .ZN(n2853) );
  NOR2_X1 U3683 ( .A1(n2855), .A2(n2853), .ZN(n3624) );
  NAND2_X1 U3684 ( .A1(n2854), .A2(n4394), .ZN(n4111) );
  NAND2_X1 U3685 ( .A1(n4105), .A2(n4111), .ZN(n2858) );
  INV_X1 U3686 ( .A(n2855), .ZN(n2857) );
  NOR2_X1 U3687 ( .A1(n4395), .A2(n4121), .ZN(n2856) );
  AOI21_X1 U3688 ( .B1(n2858), .B2(n2857), .A(n2856), .ZN(n3627) );
  INV_X1 U3689 ( .A(n4088), .ZN(n2860) );
  NAND2_X1 U3690 ( .A1(n2861), .A2(n4372), .ZN(n3628) );
  NAND2_X1 U3691 ( .A1(n4526), .A2(n4078), .ZN(n3609) );
  NAND2_X1 U3692 ( .A1(n3628), .A2(n3609), .ZN(n4069) );
  INV_X1 U3693 ( .A(n4065), .ZN(n2862) );
  NOR2_X1 U3694 ( .A1(n4069), .A2(n2862), .ZN(n2863) );
  NAND2_X1 U3695 ( .A1(n4056), .A2(n4046), .ZN(n2864) );
  NAND2_X1 U3696 ( .A1(n2864), .A2(n3701), .ZN(n4025) );
  NAND2_X1 U3697 ( .A1(n4010), .A2(n3998), .ZN(n2866) );
  NAND2_X1 U3698 ( .A1(n4059), .A2(n4359), .ZN(n3985) );
  NAND2_X1 U3699 ( .A1(n3987), .A2(n3985), .ZN(n2868) );
  NOR2_X1 U3700 ( .A1(n4010), .A2(n3998), .ZN(n2867) );
  AOI21_X1 U3701 ( .B1(n2868), .B2(n2234), .A(n2867), .ZN(n3966) );
  NAND2_X1 U3702 ( .A1(n4340), .A2(n3977), .ZN(n2869) );
  AND2_X1 U3703 ( .A1(n3966), .A2(n2869), .ZN(n3704) );
  NAND2_X1 U3704 ( .A1(n3994), .A2(n2889), .ZN(n3635) );
  NAND2_X1 U3705 ( .A1(n3935), .A2(n4336), .ZN(n3912) );
  NAND2_X1 U3706 ( .A1(n3914), .A2(n3912), .ZN(n3708) );
  INV_X1 U3707 ( .A(n3708), .ZN(n2871) );
  NAND2_X1 U3708 ( .A1(n3910), .A2(n2871), .ZN(n2875) );
  NOR2_X1 U3709 ( .A1(n3935), .A2(n4336), .ZN(n3911) );
  AND2_X1 U3710 ( .A1(n3911), .A2(n3914), .ZN(n2874) );
  NAND2_X1 U3711 ( .A1(n4320), .A2(n3917), .ZN(n2873) );
  NAND2_X1 U3712 ( .A1(n2873), .A2(n2872), .ZN(n3638) );
  NOR2_X1 U3713 ( .A1(n2874), .A2(n3638), .ZN(n3706) );
  NAND2_X1 U3714 ( .A1(n2875), .A2(n3706), .ZN(n3894) );
  OR2_X1 U3715 ( .A1(n3880), .A2(n3904), .ZN(n3666) );
  OR2_X1 U3716 ( .A1(n4320), .A2(n3917), .ZN(n3893) );
  AND2_X1 U3717 ( .A1(n3666), .A2(n3893), .ZN(n3709) );
  NAND2_X1 U3718 ( .A1(n3880), .A2(n3904), .ZN(n3667) );
  AND2_X1 U3719 ( .A1(n3900), .A2(n3885), .ZN(n3664) );
  NAND2_X1 U3720 ( .A1(n3433), .A2(n3863), .ZN(n2876) );
  NAND2_X1 U3721 ( .A1(n4323), .A2(n3879), .ZN(n3858) );
  AND2_X1 U3722 ( .A1(n2876), .A2(n3858), .ZN(n3719) );
  AND2_X1 U3723 ( .A1(n4303), .A2(n3869), .ZN(n3643) );
  INV_X1 U3724 ( .A(n3643), .ZN(n2877) );
  XNOR2_X1 U3725 ( .A(n3828), .B(n4302), .ZN(n3716) );
  OR2_X1 U3726 ( .A1(n3828), .A2(n3852), .ZN(n3649) );
  XNOR2_X1 U3727 ( .A(n2053), .B(n3693), .ZN(n2882) );
  NAND2_X1 U3728 ( .A1(n3736), .A2(n3732), .ZN(n2881) );
  NAND2_X1 U3729 ( .A1(n3727), .A2(n4514), .ZN(n2880) );
  NAND2_X1 U3730 ( .A1(n2882), .A2(n4421), .ZN(n3834) );
  OAI211_X1 U3731 ( .C1(n3839), .C2(n4437), .A(n2883), .B(n3834), .ZN(n2894)
         );
  NOR2_X1 U3732 ( .A1(n3055), .A2(n2885), .ZN(n2886) );
  MUX2_X1 U3733 ( .A(REG1_REG_28__SCAN_IN), .B(n2894), .S(n4739), .Z(n2888) );
  INV_X1 U3734 ( .A(n2888), .ZN(n2891) );
  NAND2_X1 U3735 ( .A1(n3083), .A2(n3073), .ZN(n3153) );
  NAND2_X1 U3736 ( .A1(n4405), .A2(n4273), .ZN(n4275) );
  NAND2_X1 U3737 ( .A1(n3923), .A2(n3904), .ZN(n3899) );
  OAI21_X1 U3738 ( .B1(n3846), .B2(n3833), .A(n2910), .ZN(n3826) );
  NAND2_X1 U3739 ( .A1(n2891), .A2(n2890), .ZN(U3546) );
  INV_X1 U3740 ( .A(n2892), .ZN(n3063) );
  MUX2_X1 U3741 ( .A(REG0_REG_28__SCAN_IN), .B(n2894), .S(n4733), .Z(n2895) );
  INV_X1 U3742 ( .A(n2895), .ZN(n2897) );
  NAND2_X1 U3743 ( .A1(n2897), .A2(n2896), .ZN(U3514) );
  NAND2_X1 U3744 ( .A1(n3651), .A2(DATAI_29_), .ZN(n3657) );
  XNOR2_X1 U3745 ( .A(n3827), .B(n3657), .ZN(n3694) );
  XNOR2_X1 U3746 ( .A(n2900), .B(n3694), .ZN(n3813) );
  INV_X1 U3747 ( .A(n3642), .ZN(n2901) );
  INV_X1 U3748 ( .A(n3694), .ZN(n2902) );
  AOI21_X1 U3749 ( .B1(n4513), .B2(B_REG_SCAN_IN), .A(n4429), .ZN(n3808) );
  INV_X1 U3750 ( .A(REG0_REG_30__SCAN_IN), .ZN(n2906) );
  NAND2_X1 U3751 ( .A1(n4742), .A2(REG2_REG_30__SCAN_IN), .ZN(n2905) );
  INV_X1 U3752 ( .A(REG1_REG_30__SCAN_IN), .ZN(n2903) );
  OR2_X1 U3753 ( .A1(n2360), .A2(n2903), .ZN(n2904) );
  OAI211_X1 U3754 ( .C1(n3652), .C2(n2906), .A(n2905), .B(n2904), .ZN(n3741)
         );
  NAND2_X1 U3755 ( .A1(n3848), .A2(n4434), .ZN(n2908) );
  INV_X1 U3756 ( .A(n2910), .ZN(n2911) );
  INV_X1 U3757 ( .A(n3657), .ZN(n3817) );
  OAI21_X1 U3758 ( .B1(n2911), .B2(n3657), .A(n2029), .ZN(n3820) );
  INV_X1 U3759 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2914) );
  MUX2_X1 U3760 ( .A(n2914), .B(n2913), .S(n4733), .Z(n2916) );
  NAND2_X1 U3761 ( .A1(n2916), .A2(n2915), .ZN(U3515) );
  INV_X1 U3762 ( .A(n4695), .ZN(n2917) );
  INV_X1 U3763 ( .A(DATAI_3_), .ZN(n2918) );
  INV_X1 U3764 ( .A(n3759), .ZN(n2986) );
  MUX2_X1 U3765 ( .A(n2918), .B(n2986), .S(STATE_REG_SCAN_IN), .Z(n2919) );
  INV_X1 U3766 ( .A(n2919), .ZN(U3349) );
  MUX2_X1 U3767 ( .A(n3770), .B(n2369), .S(U3149), .Z(n2920) );
  INV_X1 U3768 ( .A(n2920), .ZN(U3347) );
  INV_X1 U3769 ( .A(DATAI_15_), .ZN(n4174) );
  NAND2_X1 U3770 ( .A1(n3339), .A2(STATE_REG_SCAN_IN), .ZN(n2921) );
  OAI21_X1 U3771 ( .B1(STATE_REG_SCAN_IN), .B2(n4174), .A(n2921), .ZN(U3337)
         );
  INV_X1 U3772 ( .A(DATAI_13_), .ZN(n2923) );
  NAND2_X1 U3773 ( .A1(n3325), .A2(STATE_REG_SCAN_IN), .ZN(n2922) );
  OAI21_X1 U3774 ( .B1(STATE_REG_SCAN_IN), .B2(n2923), .A(n2922), .ZN(U3339)
         );
  INV_X1 U3775 ( .A(DATAI_19_), .ZN(n4220) );
  MUX2_X1 U3776 ( .A(n4220), .B(n3802), .S(STATE_REG_SCAN_IN), .Z(n2924) );
  INV_X1 U3777 ( .A(n2924), .ZN(U3333) );
  INV_X1 U3778 ( .A(DATAI_21_), .ZN(n2926) );
  NAND2_X1 U3779 ( .A1(n3727), .A2(STATE_REG_SCAN_IN), .ZN(n2925) );
  OAI21_X1 U3780 ( .B1(STATE_REG_SCAN_IN), .B2(n2926), .A(n2925), .ZN(U3331)
         );
  NAND3_X1 U3781 ( .A1(IR_REG_31__SCAN_IN), .A2(STATE_REG_SCAN_IN), .A3(n2258), 
        .ZN(n2927) );
  INV_X1 U3782 ( .A(DATAI_31_), .ZN(n4192) );
  OAI22_X1 U3783 ( .A1(n2928), .A2(n2927), .B1(STATE_REG_SCAN_IN), .B2(n4192), 
        .ZN(U3321) );
  INV_X1 U3784 ( .A(DATAI_22_), .ZN(n2930) );
  NAND2_X1 U3785 ( .A1(n3736), .A2(STATE_REG_SCAN_IN), .ZN(n2929) );
  OAI21_X1 U3786 ( .B1(STATE_REG_SCAN_IN), .B2(n2930), .A(n2929), .ZN(U3330)
         );
  INV_X1 U3787 ( .A(DATAI_26_), .ZN(n2933) );
  NAND2_X1 U3788 ( .A1(n2931), .A2(STATE_REG_SCAN_IN), .ZN(n2932) );
  OAI21_X1 U3789 ( .B1(STATE_REG_SCAN_IN), .B2(n2933), .A(n2932), .ZN(U3326)
         );
  INV_X1 U3790 ( .A(DATAI_25_), .ZN(n2936) );
  NAND2_X1 U3791 ( .A1(n2934), .A2(STATE_REG_SCAN_IN), .ZN(n2935) );
  OAI21_X1 U3792 ( .B1(STATE_REG_SCAN_IN), .B2(n2936), .A(n2935), .ZN(U3327)
         );
  INV_X1 U3793 ( .A(DATAI_24_), .ZN(n2937) );
  MUX2_X1 U3794 ( .A(n2734), .B(n2937), .S(U3149), .Z(n2938) );
  INV_X1 U3795 ( .A(n2938), .ZN(U3328) );
  INV_X1 U3796 ( .A(DATAI_30_), .ZN(n2941) );
  NAND2_X1 U3797 ( .A1(n2939), .A2(STATE_REG_SCAN_IN), .ZN(n2940) );
  OAI21_X1 U3798 ( .B1(STATE_REG_SCAN_IN), .B2(n2941), .A(n2940), .ZN(U3322)
         );
  NAND2_X1 U3799 ( .A1(n2944), .A2(n2942), .ZN(n2943) );
  INV_X1 U3800 ( .A(n2957), .ZN(n2945) );
  OR2_X1 U3801 ( .A1(n2944), .A2(U3149), .ZN(n3739) );
  NAND2_X1 U3802 ( .A1(n2946), .A2(n3739), .ZN(n2958) );
  NOR2_X1 U3803 ( .A1(n4635), .A2(U4043), .ZN(U3148) );
  INV_X1 U3804 ( .A(n2946), .ZN(n2947) );
  NAND3_X1 U3805 ( .A1(n4695), .A2(n2952), .A3(n2949), .ZN(n2950) );
  OAI21_X1 U3806 ( .B1(n4694), .B2(D_REG_1__SCAN_IN), .A(n2950), .ZN(n2951) );
  INV_X1 U3807 ( .A(n2951), .ZN(U3459) );
  NAND3_X1 U3808 ( .A1(n4695), .A2(n2734), .A3(n2952), .ZN(n2953) );
  OAI21_X1 U3809 ( .B1(n4694), .B2(D_REG_0__SCAN_IN), .A(n2953), .ZN(n2954) );
  INV_X1 U3810 ( .A(n2954), .ZN(U3458) );
  INV_X1 U3811 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3070) );
  AND2_X1 U3812 ( .A1(n4513), .A2(n3070), .ZN(n2955) );
  NOR2_X1 U3813 ( .A1(n4521), .A2(n2955), .ZN(n3025) );
  OAI21_X1 U3814 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4513), .A(n3025), .ZN(n2956)
         );
  MUX2_X1 U3815 ( .A(n2956), .B(n3025), .S(IR_REG_0__SCAN_IN), .Z(n2963) );
  INV_X1 U3816 ( .A(n2980), .ZN(n2962) );
  INV_X1 U3817 ( .A(n4513), .ZN(n3021) );
  NAND3_X1 U3818 ( .A1(n4637), .A2(IR_REG_0__SCAN_IN), .A3(n2959), .ZN(n2961)
         );
  AOI22_X1 U3819 ( .A1(n4635), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n2960) );
  OAI211_X1 U3820 ( .C1(n2963), .C2(n2962), .A(n2961), .B(n2960), .ZN(U3240)
         );
  INV_X1 U3821 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n2965) );
  NAND2_X1 U3822 ( .A1(n4416), .A2(U4043), .ZN(n2964) );
  OAI21_X1 U3823 ( .B1(U4043), .B2(n2965), .A(n2964), .ZN(U3560) );
  INV_X1 U3824 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2966) );
  MUX2_X1 U3825 ( .A(REG2_REG_2__SCAN_IN), .B(n2966), .S(n4518), .Z(n3029) );
  INV_X1 U3826 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3131) );
  MUX2_X1 U3827 ( .A(REG2_REG_1__SCAN_IN), .B(n3131), .S(n4519), .Z(n3751) );
  AND2_X1 U3828 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2967)
         );
  NAND2_X1 U3829 ( .A1(n3751), .A2(n2967), .ZN(n3750) );
  NAND2_X1 U3830 ( .A1(n4519), .A2(REG2_REG_1__SCAN_IN), .ZN(n2968) );
  NAND2_X1 U3831 ( .A1(n3750), .A2(n2968), .ZN(n3028) );
  NAND2_X1 U3832 ( .A1(n3029), .A2(n3028), .ZN(n3027) );
  NAND2_X1 U3833 ( .A1(n4518), .A2(REG2_REG_2__SCAN_IN), .ZN(n2969) );
  NAND2_X1 U3834 ( .A1(n3027), .A2(n2969), .ZN(n2970) );
  XNOR2_X1 U3835 ( .A(n2970), .B(n2986), .ZN(n3764) );
  NAND2_X1 U3836 ( .A1(n3764), .A2(REG2_REG_3__SCAN_IN), .ZN(n2972) );
  NAND2_X1 U3837 ( .A1(n2970), .A2(n3759), .ZN(n2971) );
  NAND2_X1 U3838 ( .A1(n2972), .A2(n2971), .ZN(n2973) );
  INV_X1 U3839 ( .A(n4517), .ZN(n3044) );
  XNOR2_X1 U3840 ( .A(n2973), .B(n3044), .ZN(n3038) );
  NAND2_X1 U3841 ( .A1(n3038), .A2(REG2_REG_4__SCAN_IN), .ZN(n2975) );
  NAND2_X1 U3842 ( .A1(n2973), .A2(n4517), .ZN(n2974) );
  NAND2_X1 U3843 ( .A1(n2975), .A2(n2974), .ZN(n3777) );
  INV_X1 U3844 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2976) );
  MUX2_X1 U3845 ( .A(n2976), .B(REG2_REG_5__SCAN_IN), .S(n3770), .Z(n3778) );
  NAND2_X1 U3846 ( .A1(n3777), .A2(n3778), .ZN(n3776) );
  OR2_X1 U3847 ( .A1(n3770), .A2(n2976), .ZN(n2977) );
  NAND2_X1 U3848 ( .A1(n3776), .A2(n2977), .ZN(n3008) );
  INV_X1 U3849 ( .A(n4516), .ZN(n2992) );
  XNOR2_X1 U3850 ( .A(n3008), .B(n2992), .ZN(n3010) );
  XNOR2_X1 U3851 ( .A(n3010), .B(REG2_REG_6__SCAN_IN), .ZN(n2996) );
  NAND2_X1 U3852 ( .A1(n3020), .A2(n4513), .ZN(n3735) );
  INV_X1 U3853 ( .A(n3735), .ZN(n2978) );
  NOR2_X1 U3854 ( .A1(STATE_REG_SCAN_IN), .A2(n2979), .ZN(n3167) );
  NOR2_X1 U3855 ( .A1(n4641), .A2(n2992), .ZN(n2981) );
  AOI211_X1 U3856 ( .C1(n4635), .C2(ADDR_REG_6__SCAN_IN), .A(n3167), .B(n2981), 
        .ZN(n2995) );
  INV_X1 U3857 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2982) );
  INV_X1 U3858 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2983) );
  XNOR2_X1 U3859 ( .A(n4519), .B(n2983), .ZN(n3754) );
  AND2_X1 U3860 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3753)
         );
  NAND2_X1 U3861 ( .A1(n4519), .A2(REG1_REG_1__SCAN_IN), .ZN(n2984) );
  NAND2_X1 U3862 ( .A1(n4518), .A2(REG1_REG_2__SCAN_IN), .ZN(n2985) );
  NAND2_X1 U3863 ( .A1(n3762), .A2(REG1_REG_3__SCAN_IN), .ZN(n3761) );
  NAND2_X1 U3864 ( .A1(n2987), .A2(n3759), .ZN(n2988) );
  NAND2_X1 U3865 ( .A1(n3761), .A2(n2988), .ZN(n2989) );
  INV_X1 U3866 ( .A(n2989), .ZN(n2990) );
  XNOR2_X1 U3867 ( .A(n2989), .B(n3044), .ZN(n3040) );
  NAND2_X1 U3868 ( .A1(n3040), .A2(REG1_REG_4__SCAN_IN), .ZN(n3039) );
  OAI21_X1 U3869 ( .B1(n2990), .B2(n3044), .A(n3039), .ZN(n3774) );
  XNOR2_X1 U3870 ( .A(n3770), .B(REG1_REG_5__SCAN_IN), .ZN(n3775) );
  NAND2_X1 U3871 ( .A1(n3774), .A2(n3775), .ZN(n3773) );
  XNOR2_X1 U3872 ( .A(n3005), .B(n2992), .ZN(n2993) );
  NAND2_X1 U3873 ( .A1(n2993), .A2(REG1_REG_6__SCAN_IN), .ZN(n3004) );
  OAI211_X1 U3874 ( .C1(REG1_REG_6__SCAN_IN), .C2(n2993), .A(n4637), .B(n3004), 
        .ZN(n2994) );
  OAI211_X1 U3875 ( .C1(n2996), .C2(n4630), .A(n2995), .B(n2994), .ZN(U3246)
         );
  INV_X1 U3876 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n2998) );
  NAND2_X1 U3877 ( .A1(n4526), .A2(U4043), .ZN(n2997) );
  OAI21_X1 U3878 ( .B1(U4043), .B2(n2998), .A(n2997), .ZN(U3565) );
  INV_X1 U3879 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n4261) );
  NAND2_X1 U3880 ( .A1(n3441), .A2(U4043), .ZN(n2999) );
  OAI21_X1 U3881 ( .B1(U4043), .B2(n4261), .A(n2999), .ZN(U3558) );
  INV_X1 U3882 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n3001) );
  NAND2_X1 U3883 ( .A1(n4373), .A2(U4043), .ZN(n3000) );
  OAI21_X1 U3884 ( .B1(U4043), .B2(n3001), .A(n3000), .ZN(U3566) );
  INV_X1 U3885 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n3003) );
  NAND2_X1 U3886 ( .A1(n3880), .A2(U4043), .ZN(n3002) );
  OAI21_X1 U3887 ( .B1(U4043), .B2(n3003), .A(n3002), .ZN(U3574) );
  XNOR2_X1 U3888 ( .A(n4515), .B(REG1_REG_7__SCAN_IN), .ZN(n3007) );
  OAI21_X1 U3889 ( .B1(n3211), .B2(n3007), .A(n4637), .ZN(n3006) );
  AOI21_X1 U3890 ( .B1(n3211), .B2(n3007), .A(n3006), .ZN(n3017) );
  AND2_X1 U3891 ( .A1(n3008), .A2(n4516), .ZN(n3009) );
  AOI21_X1 U3892 ( .B1(n3010), .B2(REG2_REG_6__SCAN_IN), .A(n3009), .ZN(n3012)
         );
  INV_X1 U3893 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3295) );
  MUX2_X1 U3894 ( .A(n3295), .B(REG2_REG_7__SCAN_IN), .S(n4515), .Z(n3011) );
  NOR2_X1 U3895 ( .A1(n3012), .A2(n3011), .ZN(n3227) );
  AOI211_X1 U3896 ( .C1(n3012), .C2(n3011), .A(n3227), .B(n4630), .ZN(n3016)
         );
  INV_X1 U3897 ( .A(n4515), .ZN(n3228) );
  NAND2_X1 U3898 ( .A1(REG3_REG_7__SCAN_IN), .A2(U3149), .ZN(n3444) );
  INV_X1 U3899 ( .A(n3444), .ZN(n3013) );
  AOI21_X1 U3900 ( .B1(n4635), .B2(ADDR_REG_7__SCAN_IN), .A(n3013), .ZN(n3014)
         );
  OAI21_X1 U3901 ( .B1(n4641), .B2(n3228), .A(n3014), .ZN(n3015) );
  OR3_X1 U3902 ( .A1(n3017), .A2(n3016), .A3(n3015), .ZN(U3247) );
  XNOR2_X1 U3903 ( .A(n3019), .B(n3018), .ZN(n3096) );
  NAND3_X1 U3904 ( .A1(n3096), .A2(n3021), .A3(n3020), .ZN(n3024) );
  NAND2_X1 U3905 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3749) );
  OAI21_X1 U3906 ( .B1(n3735), .B2(n3749), .A(U4043), .ZN(n3022) );
  INV_X1 U3907 ( .A(n3022), .ZN(n3023) );
  OAI211_X1 U3908 ( .C1(IR_REG_0__SCAN_IN), .C2(n3025), .A(n3024), .B(n3023), 
        .ZN(n3047) );
  INV_X1 U3909 ( .A(n4641), .ZN(n3760) );
  NAND2_X1 U3910 ( .A1(n4635), .A2(ADDR_REG_2__SCAN_IN), .ZN(n3026) );
  OAI21_X1 U3911 ( .B1(STATE_REG_SCAN_IN), .B2(n3136), .A(n3026), .ZN(n3036)
         );
  OAI211_X1 U3912 ( .C1(n3029), .C2(n3028), .A(n4591), .B(n3027), .ZN(n3034)
         );
  OAI211_X1 U3913 ( .C1(n3032), .C2(n3031), .A(n4637), .B(n3030), .ZN(n3033)
         );
  NAND2_X1 U3914 ( .A1(n3034), .A2(n3033), .ZN(n3035) );
  AOI211_X1 U3915 ( .C1(n4518), .C2(n3760), .A(n3036), .B(n3035), .ZN(n3037)
         );
  NAND2_X1 U3916 ( .A1(n3047), .A2(n3037), .ZN(U3242) );
  INV_X1 U3917 ( .A(REG2_REG_4__SCAN_IN), .ZN(n4206) );
  MUX2_X1 U3918 ( .A(n4206), .B(REG2_REG_4__SCAN_IN), .S(n3038), .Z(n3048) );
  OAI211_X1 U3919 ( .C1(REG1_REG_4__SCAN_IN), .C2(n3040), .A(n4637), .B(n3039), 
        .ZN(n3043) );
  NAND2_X1 U3920 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3191) );
  INV_X1 U3921 ( .A(n3191), .ZN(n3041) );
  AOI21_X1 U3922 ( .B1(n4635), .B2(ADDR_REG_4__SCAN_IN), .A(n3041), .ZN(n3042)
         );
  OAI211_X1 U3923 ( .C1(n4641), .C2(n3044), .A(n3043), .B(n3042), .ZN(n3045)
         );
  INV_X1 U3924 ( .A(n3045), .ZN(n3046) );
  OAI211_X1 U3925 ( .C1(n3048), .C2(n4630), .A(n3047), .B(n3046), .ZN(U3244)
         );
  NAND2_X1 U3926 ( .A1(n3748), .A2(n3073), .ZN(n3587) );
  NAND2_X1 U3927 ( .A1(n3078), .A2(n3587), .ZN(n3672) );
  INV_X1 U3928 ( .A(n3065), .ZN(n3049) );
  NOR2_X1 U3929 ( .A1(n3073), .A2(n3049), .ZN(n3051) );
  INV_X1 U3930 ( .A(n4419), .ZN(n3261) );
  OAI21_X1 U3931 ( .B1(n3261), .B2(n4421), .A(n3672), .ZN(n3050) );
  OAI21_X1 U3932 ( .B1(n2797), .B2(n4429), .A(n3050), .ZN(n3068) );
  AOI211_X1 U3933 ( .C1(n4724), .C2(n3672), .A(n3051), .B(n3068), .ZN(n4714)
         );
  NAND2_X1 U3934 ( .A1(n4737), .A2(REG1_REG_0__SCAN_IN), .ZN(n3052) );
  OAI21_X1 U3935 ( .B1(n4714), .B2(n4737), .A(n3052), .ZN(U3518) );
  XNOR2_X1 U3936 ( .A(n3053), .B(n3054), .ZN(n3059) );
  INV_X1 U3937 ( .A(n3055), .ZN(n3061) );
  NAND2_X1 U3938 ( .A1(n3056), .A2(n3061), .ZN(n3101) );
  AOI22_X1 U3939 ( .A1(n3570), .A2(n3746), .B1(REG3_REG_1__SCAN_IN), .B2(n3101), .ZN(n3058) );
  AOI22_X1 U3940 ( .A1(n3126), .A2(n4523), .B1(n4527), .B2(n3748), .ZN(n3057)
         );
  OAI211_X1 U3941 ( .C1(n3059), .C2(n3584), .A(n3058), .B(n3057), .ZN(U3219)
         );
  NAND4_X1 U3942 ( .A1(n3063), .A2(n3062), .A3(n3061), .A4(n3060), .ZN(n3064)
         );
  INV_X2 U3943 ( .A(n4663), .ZN(n4022) );
  NAND2_X1 U3944 ( .A1(n4022), .A2(n3802), .ZN(n4018) );
  INV_X1 U3945 ( .A(n4018), .ZN(n3297) );
  AOI21_X1 U3946 ( .B1(n3297), .B2(n3065), .A(n4279), .ZN(n3074) );
  NAND2_X1 U3947 ( .A1(n3066), .A2(n3732), .ZN(n3175) );
  INV_X1 U3948 ( .A(n3175), .ZN(n3067) );
  AND2_X1 U3949 ( .A1(n4022), .A2(n3067), .ZN(n4658) );
  AOI22_X1 U3950 ( .A1(n3068), .A2(n4022), .B1(REG3_REG_0__SCAN_IN), .B2(n4653), .ZN(n3069) );
  OAI21_X1 U3951 ( .B1(n3070), .B2(n4022), .A(n3069), .ZN(n3071) );
  AOI21_X1 U3952 ( .B1(n4658), .B2(n3672), .A(n3071), .ZN(n3072) );
  OAI21_X1 U3953 ( .B1(n3074), .B2(n3073), .A(n3072), .ZN(U3290) );
  OR2_X1 U3954 ( .A1(n3075), .A2(n2842), .ZN(n3076) );
  NAND2_X1 U3955 ( .A1(n3077), .A2(n3076), .ZN(n3125) );
  INV_X1 U3956 ( .A(n3125), .ZN(n3082) );
  INV_X1 U3957 ( .A(n2842), .ZN(n3080) );
  INV_X1 U3958 ( .A(n3078), .ZN(n3588) );
  OAI21_X1 U3959 ( .B1(n3080), .B2(n3588), .A(n3079), .ZN(n3081) );
  AOI22_X1 U3960 ( .A1(n3261), .A2(n3082), .B1(n3081), .B2(n4421), .ZN(n3132)
         );
  OAI22_X1 U3961 ( .A1(n3084), .A2(n4429), .B1(n4428), .B2(n3083), .ZN(n3085)
         );
  AOI21_X1 U3962 ( .B1(n4434), .B2(n3748), .A(n3085), .ZN(n3086) );
  OAI211_X1 U3963 ( .C1(n4350), .C2(n3125), .A(n3132), .B(n3086), .ZN(n3091)
         );
  NAND2_X1 U3964 ( .A1(n3126), .A2(n3093), .ZN(n3087) );
  NAND2_X1 U3965 ( .A1(n3153), .A2(n3087), .ZN(n3128) );
  OAI22_X1 U3966 ( .A1(n4440), .A2(n3128), .B1(n4739), .B2(n2983), .ZN(n3088)
         );
  AOI21_X1 U3967 ( .B1(n3091), .B2(n4739), .A(n3088), .ZN(n3089) );
  INV_X1 U3968 ( .A(n3089), .ZN(U3519) );
  OAI22_X1 U3969 ( .A1(n4511), .A2(n3128), .B1(n4733), .B2(n2305), .ZN(n3090)
         );
  AOI21_X1 U3970 ( .B1(n3091), .B2(n4733), .A(n3090), .ZN(n3092) );
  INV_X1 U3971 ( .A(n3092), .ZN(U3469) );
  AOI22_X1 U3972 ( .A1(n3570), .A2(n2799), .B1(REG3_REG_0__SCAN_IN), .B2(n3101), .ZN(n3095) );
  NAND2_X1 U3973 ( .A1(n3569), .A2(n3093), .ZN(n3094) );
  OAI211_X1 U3974 ( .C1(n3584), .C2(n3096), .A(n3095), .B(n3094), .ZN(U3229)
         );
  INV_X1 U3975 ( .A(n3097), .ZN(n3098) );
  AOI21_X1 U3976 ( .B1(n3100), .B2(n3099), .A(n3098), .ZN(n3104) );
  AOI22_X1 U3977 ( .A1(n3570), .A2(n3745), .B1(REG3_REG_2__SCAN_IN), .B2(n3101), .ZN(n3103) );
  AOI22_X1 U3978 ( .A1(n3152), .A2(n3569), .B1(n4527), .B2(n2799), .ZN(n3102)
         );
  OAI211_X1 U3979 ( .C1(n3104), .C2(n3584), .A(n3103), .B(n3102), .ZN(U3234)
         );
  INV_X1 U3980 ( .A(n3105), .ZN(n3106) );
  AOI21_X1 U3981 ( .B1(n3684), .B2(n3107), .A(n3106), .ZN(n3113) );
  INV_X1 U3982 ( .A(n3113), .ZN(n3139) );
  AOI22_X1 U3983 ( .A1(n3745), .A2(n4414), .B1(n3152), .B2(n4412), .ZN(n3108)
         );
  OAI21_X1 U3984 ( .B1(n2797), .B2(n4397), .A(n3108), .ZN(n3114) );
  OAI21_X1 U3985 ( .B1(n3684), .B2(n3110), .A(n3109), .ZN(n3111) );
  NAND2_X1 U3986 ( .A1(n3111), .A2(n4421), .ZN(n3112) );
  OAI21_X1 U3987 ( .B1(n3113), .B2(n4419), .A(n3112), .ZN(n3135) );
  AOI211_X1 U3988 ( .C1(n4724), .C2(n3139), .A(n3114), .B(n3135), .ZN(n3185)
         );
  XNOR2_X1 U3989 ( .A(n3153), .B(n3152), .ZN(n3187) );
  OAI22_X1 U3990 ( .A1(n4511), .A2(n3187), .B1(n4733), .B2(n3115), .ZN(n3116)
         );
  INV_X1 U3991 ( .A(n3116), .ZN(n3117) );
  OAI21_X1 U3992 ( .B1(n3185), .B2(n4732), .A(n3117), .ZN(U3471) );
  XNOR2_X1 U3993 ( .A(n3119), .B(n3118), .ZN(n3123) );
  AOI22_X1 U3994 ( .A1(n3242), .A2(n4523), .B1(n4527), .B2(n2806), .ZN(n3122)
         );
  AND2_X1 U3995 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3772) );
  NOR2_X1 U3996 ( .A1(n4543), .A2(n3178), .ZN(n3120) );
  AOI211_X1 U3997 ( .C1(n3570), .C2(n3743), .A(n3772), .B(n3120), .ZN(n3121)
         );
  OAI211_X1 U3998 ( .C1(n3123), .C2(n3584), .A(n3122), .B(n3121), .ZN(U3224)
         );
  INV_X1 U3999 ( .A(n4658), .ZN(n4644) );
  OAI22_X1 U4000 ( .A1(n4644), .A2(n3125), .B1(n3124), .B2(n4647), .ZN(n3130)
         );
  INV_X1 U4001 ( .A(n4346), .ZN(n4719) );
  NAND2_X1 U4002 ( .A1(n4022), .A2(n4434), .ZN(n3815) );
  AOI22_X1 U4003 ( .A1(n4282), .A2(n3748), .B1(n4279), .B2(n3126), .ZN(n3127)
         );
  OAI21_X1 U4004 ( .B1(n4643), .B2(n3128), .A(n3127), .ZN(n3129) );
  AOI211_X1 U4005 ( .C1(n4280), .C2(n3746), .A(n3130), .B(n3129), .ZN(n3134)
         );
  MUX2_X1 U4006 ( .A(n3132), .B(n3131), .S(n4663), .Z(n3133) );
  NAND2_X1 U4007 ( .A1(n3134), .A2(n3133), .ZN(U3289) );
  MUX2_X1 U4008 ( .A(REG2_REG_2__SCAN_IN), .B(n3135), .S(n4022), .Z(n3143) );
  OAI22_X1 U4009 ( .A1(n4097), .A2(n3137), .B1(n3136), .B2(n4647), .ZN(n3138)
         );
  AOI21_X1 U4010 ( .B1(n3139), .B2(n4658), .A(n3138), .ZN(n3141) );
  AOI22_X1 U4011 ( .A1(n4282), .A2(n2799), .B1(n4280), .B2(n3745), .ZN(n3140)
         );
  OAI211_X1 U4012 ( .C1(n3187), .C2(n4643), .A(n3141), .B(n3140), .ZN(n3142)
         );
  OR2_X1 U4013 ( .A1(n3143), .A2(n3142), .ZN(U3288) );
  NAND2_X1 U4014 ( .A1(n3105), .A2(n3144), .ZN(n3145) );
  INV_X1 U4015 ( .A(n3148), .ZN(n3687) );
  XNOR2_X1 U4016 ( .A(n3145), .B(n3687), .ZN(n3199) );
  OAI22_X1 U4017 ( .A1(n2802), .A2(n4429), .B1(n4428), .B2(n3200), .ZN(n3151)
         );
  OAI21_X1 U4018 ( .B1(n3148), .B2(n3147), .A(n3146), .ZN(n3149) );
  AOI22_X1 U4019 ( .A1(n3149), .A2(n4421), .B1(n4434), .B2(n3746), .ZN(n3150)
         );
  INV_X1 U4020 ( .A(n3150), .ZN(n3206) );
  AOI211_X1 U4021 ( .C1(n4726), .C2(n3199), .A(n3151), .B(n3206), .ZN(n3162)
         );
  OAI21_X1 U4022 ( .B1(n3153), .B2(n3152), .A(n3475), .ZN(n3154) );
  INV_X1 U4023 ( .A(n3154), .ZN(n3155) );
  OR2_X1 U4024 ( .A1(n3155), .A2(n3266), .ZN(n3204) );
  OAI22_X1 U4025 ( .A1(n4440), .A2(n3204), .B1(n4739), .B2(n3156), .ZN(n3157)
         );
  INV_X1 U4026 ( .A(n3157), .ZN(n3158) );
  OAI21_X1 U4027 ( .B1(n3162), .B2(n4737), .A(n3158), .ZN(U3521) );
  OAI22_X1 U4028 ( .A1(n4511), .A2(n3204), .B1(n4733), .B2(n3159), .ZN(n3160)
         );
  INV_X1 U4029 ( .A(n3160), .ZN(n3161) );
  OAI21_X1 U4030 ( .B1(n3162), .B2(n4732), .A(n3161), .ZN(U3473) );
  NOR2_X1 U4031 ( .A1(n2233), .A2(n3163), .ZN(n3164) );
  XNOR2_X1 U4032 ( .A(n3165), .B(n3164), .ZN(n3170) );
  AOI22_X1 U4033 ( .A1(n3274), .A2(n3569), .B1(n4527), .B2(n3744), .ZN(n3169)
         );
  NOR2_X1 U4034 ( .A1(n4543), .A2(n3283), .ZN(n3166) );
  AOI211_X1 U4035 ( .C1(n3570), .C2(n3742), .A(n3167), .B(n3166), .ZN(n3168)
         );
  OAI211_X1 U4036 ( .C1(n3170), .C2(n3584), .A(n3169), .B(n3168), .ZN(U3236)
         );
  INV_X1 U4037 ( .A(n3171), .ZN(n3598) );
  AND2_X1 U4038 ( .A1(n3598), .A2(n3613), .ZN(n3685) );
  XOR2_X1 U4039 ( .A(n3685), .B(n3172), .Z(n3173) );
  NAND2_X1 U4040 ( .A1(n3173), .A2(n4421), .ZN(n3244) );
  XNOR2_X1 U4041 ( .A(n3174), .B(n3685), .ZN(n3246) );
  NAND2_X1 U4042 ( .A1(n4419), .A2(n3175), .ZN(n3176) );
  AOI21_X1 U40430 ( .B1(n3242), .B2(n3264), .A(n3282), .ZN(n3248) );
  INV_X1 U4044 ( .A(n3248), .ZN(n3182) );
  OAI22_X1 U4045 ( .A1(n4022), .A2(n2976), .B1(n3178), .B2(n4647), .ZN(n3180)
         );
  INV_X1 U4046 ( .A(n4280), .ZN(n3317) );
  OAI22_X1 U4047 ( .A1(n3317), .A2(n3445), .B1(n2802), .B2(n3815), .ZN(n3179)
         );
  AOI211_X1 U4048 ( .C1(n3242), .C2(n4279), .A(n3180), .B(n3179), .ZN(n3181)
         );
  OAI21_X1 U4049 ( .B1(n4643), .B2(n3182), .A(n3181), .ZN(n3183) );
  AOI21_X1 U4050 ( .B1(n3246), .B2(n4290), .A(n3183), .ZN(n3184) );
  OAI21_X1 U4051 ( .B1(n3244), .B2(n4663), .A(n3184), .ZN(U3285) );
  MUX2_X1 U4052 ( .A(n2982), .B(n3185), .S(n4739), .Z(n3186) );
  OAI21_X1 U4053 ( .B1(n3187), .B2(n4440), .A(n3186), .ZN(U3520) );
  NAND2_X1 U4054 ( .A1(n3188), .A2(n4538), .ZN(n3198) );
  AOI21_X1 U4055 ( .B1(n3470), .B2(n3190), .A(n3189), .ZN(n3197) );
  NAND2_X1 U4056 ( .A1(n4525), .A2(n3744), .ZN(n3192) );
  OAI211_X1 U4057 ( .C1(n4543), .C2(n3267), .A(n3192), .B(n3191), .ZN(n3195)
         );
  NOR2_X1 U4058 ( .A1(n3572), .A2(n3193), .ZN(n3194) );
  AOI211_X1 U4059 ( .C1(n3258), .C2(n3569), .A(n3195), .B(n3194), .ZN(n3196)
         );
  OAI21_X1 U4060 ( .B1(n3198), .B2(n3197), .A(n3196), .ZN(U3227) );
  INV_X1 U4061 ( .A(n3199), .ZN(n3208) );
  INV_X1 U4062 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3763) );
  OAI22_X1 U4063 ( .A1(n4022), .A2(n3763), .B1(REG3_REG_3__SCAN_IN), .B2(n4647), .ZN(n3202) );
  NOR2_X1 U4064 ( .A1(n4097), .A2(n3200), .ZN(n3201) );
  AOI211_X1 U4065 ( .C1(n4280), .C2(n2806), .A(n3202), .B(n3201), .ZN(n3203)
         );
  OAI21_X1 U4066 ( .B1(n4643), .B2(n3204), .A(n3203), .ZN(n3205) );
  AOI21_X1 U4067 ( .B1(n4022), .B2(n3206), .A(n3205), .ZN(n3207) );
  OAI21_X1 U4068 ( .B1(n4064), .B2(n3208), .A(n3207), .ZN(U3287) );
  NAND2_X1 U4069 ( .A1(n3225), .A2(REG1_REG_11__SCAN_IN), .ZN(n3216) );
  INV_X1 U4070 ( .A(n3225), .ZN(n4707) );
  AOI22_X1 U4071 ( .A1(n3225), .A2(REG1_REG_11__SCAN_IN), .B1(n4425), .B2(
        n4707), .ZN(n4580) );
  INV_X1 U4072 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4186) );
  INV_X1 U4073 ( .A(n3226), .ZN(n4710) );
  AOI22_X1 U4074 ( .A1(n3226), .A2(REG1_REG_9__SCAN_IN), .B1(n4186), .B2(n4710), .ZN(n4559) );
  OAI21_X1 U4075 ( .B1(n3211), .B2(n3210), .A(n3209), .ZN(n3212) );
  NAND2_X1 U4076 ( .A1(n3229), .A2(n3212), .ZN(n3213) );
  NAND2_X1 U4077 ( .A1(n4568), .A2(n3214), .ZN(n3215) );
  NAND2_X1 U4078 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4570), .ZN(n4569) );
  NAND2_X1 U4079 ( .A1(n3215), .A2(n4569), .ZN(n4579) );
  NAND2_X1 U4080 ( .A1(n4580), .A2(n4579), .ZN(n4578) );
  NAND2_X1 U4081 ( .A1(n3216), .A2(n4578), .ZN(n3217) );
  NAND2_X1 U4082 ( .A1(n4589), .A2(n3217), .ZN(n3218) );
  XOR2_X1 U4083 ( .A(n3217), .B(n4589), .Z(n4597) );
  NAND2_X1 U4084 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4597), .ZN(n4596) );
  XNOR2_X1 U4085 ( .A(n3223), .B(REG1_REG_13__SCAN_IN), .ZN(n3219) );
  OAI211_X1 U4086 ( .C1(n3220), .C2(n3219), .A(n4637), .B(n3326), .ZN(n3222)
         );
  AND2_X1 U4087 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n3550) );
  AOI21_X1 U4088 ( .B1(n4635), .B2(ADDR_REG_13__SCAN_IN), .A(n3550), .ZN(n3221) );
  OAI211_X1 U4089 ( .C1(n4641), .C2(n3223), .A(n3222), .B(n3221), .ZN(n3241)
         );
  AND2_X1 U4090 ( .A1(n3325), .A2(REG2_REG_13__SCAN_IN), .ZN(n3335) );
  INV_X1 U4091 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4123) );
  NAND2_X1 U4092 ( .A1(n3223), .A2(n4123), .ZN(n3334) );
  INV_X1 U4093 ( .A(n3334), .ZN(n3224) );
  NOR2_X1 U4094 ( .A1(n3335), .A2(n3224), .ZN(n3239) );
  NAND2_X1 U4095 ( .A1(n3225), .A2(REG2_REG_11__SCAN_IN), .ZN(n3235) );
  INV_X1 U4096 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4646) );
  AOI22_X1 U4097 ( .A1(n3225), .A2(REG2_REG_11__SCAN_IN), .B1(n4646), .B2(
        n4707), .ZN(n4583) );
  NAND2_X1 U4098 ( .A1(n3226), .A2(REG2_REG_9__SCAN_IN), .ZN(n3232) );
  INV_X1 U4099 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3319) );
  AOI22_X1 U4100 ( .A1(n3226), .A2(REG2_REG_9__SCAN_IN), .B1(n3319), .B2(n4710), .ZN(n4562) );
  NAND2_X1 U4101 ( .A1(n3229), .A2(n3230), .ZN(n3231) );
  NAND2_X1 U4102 ( .A1(n3231), .A2(n4550), .ZN(n4561) );
  NAND2_X1 U4103 ( .A1(n4562), .A2(n4561), .ZN(n4560) );
  NAND2_X1 U4104 ( .A1(n4568), .A2(n3233), .ZN(n3234) );
  NAND2_X1 U4105 ( .A1(n4583), .A2(n4582), .ZN(n4581) );
  NAND2_X1 U4106 ( .A1(n4589), .A2(n3236), .ZN(n3237) );
  OAI21_X1 U4107 ( .B1(n3239), .B2(n3336), .A(n4591), .ZN(n3238) );
  AOI21_X1 U4108 ( .B1(n3239), .B2(n3336), .A(n3238), .ZN(n3240) );
  OR2_X1 U4109 ( .A1(n3241), .A2(n3240), .ZN(U3253) );
  AOI22_X1 U4110 ( .A1(n3743), .A2(n4414), .B1(n3242), .B2(n4412), .ZN(n3243)
         );
  OAI211_X1 U4111 ( .C1(n2802), .C2(n4397), .A(n3244), .B(n3243), .ZN(n3245)
         );
  AOI21_X1 U4112 ( .B1(n3246), .B2(n4726), .A(n3245), .ZN(n3250) );
  INV_X1 U4113 ( .A(n4440), .ZN(n4297) );
  AOI22_X1 U4114 ( .A1(n3248), .A2(n4297), .B1(REG1_REG_5__SCAN_IN), .B2(n4737), .ZN(n3247) );
  OAI21_X1 U4115 ( .B1(n3250), .B2(n4737), .A(n3247), .ZN(U3523) );
  INV_X1 U4116 ( .A(n4511), .ZN(n4446) );
  AOI22_X1 U4117 ( .A1(n3248), .A2(n4446), .B1(REG0_REG_5__SCAN_IN), .B2(n4732), .ZN(n3249) );
  OAI21_X1 U4118 ( .B1(n3250), .B2(n4732), .A(n3249), .ZN(U3477) );
  NAND2_X1 U4119 ( .A1(n3105), .A2(n3251), .ZN(n3253) );
  AND2_X1 U4120 ( .A1(n3253), .A2(n3252), .ZN(n3256) );
  INV_X1 U4121 ( .A(n4718), .ZN(n3271) );
  AOI22_X1 U4122 ( .A1(n3745), .A2(n4434), .B1(n3258), .B2(n4412), .ZN(n3259)
         );
  OAI21_X1 U4123 ( .B1(n3276), .B2(n4429), .A(n3259), .ZN(n3260) );
  AOI21_X1 U4124 ( .B1(n4718), .B2(n3261), .A(n3260), .ZN(n3262) );
  OAI21_X1 U4125 ( .B1(n4115), .B2(n3263), .A(n3262), .ZN(n4716) );
  OAI211_X1 U4126 ( .C1(n3266), .C2(n3265), .A(n3264), .B(n4346), .ZN(n4715)
         );
  OAI22_X1 U4127 ( .A1(n4715), .A2(n3732), .B1(n4647), .B2(n3267), .ZN(n3268)
         );
  NOR2_X1 U4128 ( .A1(n4716), .A2(n3268), .ZN(n3269) );
  MUX2_X1 U4129 ( .A(n4206), .B(n3269), .S(n4022), .Z(n3270) );
  OAI21_X1 U4130 ( .B1(n3271), .B2(n4644), .A(n3270), .ZN(U3286) );
  NAND2_X1 U4131 ( .A1(n3601), .A2(n3615), .ZN(n3674) );
  XNOR2_X1 U4132 ( .A(n3272), .B(n3674), .ZN(n3280) );
  XOR2_X1 U4133 ( .A(n3674), .B(n3273), .Z(n3278) );
  AOI22_X1 U4134 ( .A1(n3742), .A2(n4414), .B1(n4412), .B2(n3274), .ZN(n3275)
         );
  OAI21_X1 U4135 ( .B1(n3276), .B2(n4397), .A(n3275), .ZN(n3277) );
  AOI21_X1 U4136 ( .B1(n3278), .B2(n4421), .A(n3277), .ZN(n3279) );
  OAI21_X1 U4137 ( .B1(n4419), .B2(n3280), .A(n3279), .ZN(n4722) );
  INV_X1 U4138 ( .A(n4722), .ZN(n3288) );
  INV_X1 U4139 ( .A(n3280), .ZN(n4725) );
  NOR2_X1 U4140 ( .A1(n3282), .A2(n3281), .ZN(n4721) );
  NOR3_X1 U4141 ( .A1(n4721), .A2(n4720), .A3(n4643), .ZN(n3286) );
  INV_X1 U4142 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3284) );
  OAI22_X1 U4143 ( .A1(n4022), .A2(n3284), .B1(n3283), .B2(n4647), .ZN(n3285)
         );
  AOI211_X1 U4144 ( .C1(n4725), .C2(n4658), .A(n3286), .B(n3285), .ZN(n3287)
         );
  OAI21_X1 U4145 ( .B1(n3288), .B2(n4663), .A(n3287), .ZN(U3284) );
  OAI22_X1 U4146 ( .A1(n3398), .A2(n4429), .B1(n3293), .B2(n4428), .ZN(n3292)
         );
  INV_X1 U4147 ( .A(n3602), .ZN(n3673) );
  XNOR2_X1 U4148 ( .A(n3289), .B(n3673), .ZN(n3290) );
  NOR2_X1 U4149 ( .A1(n3290), .A2(n4115), .ZN(n3291) );
  AOI211_X1 U4150 ( .C1(n4434), .C2(n3743), .A(n3292), .B(n3291), .ZN(n4731)
         );
  OAI21_X1 U4151 ( .B1(n4720), .B2(n3293), .A(n4346), .ZN(n3294) );
  OR2_X1 U4152 ( .A1(n3294), .A2(n3358), .ZN(n4730) );
  INV_X1 U4153 ( .A(n4730), .ZN(n3298) );
  OAI22_X1 U4154 ( .A1(n4022), .A2(n3295), .B1(n3443), .B2(n4647), .ZN(n3296)
         );
  AOI21_X1 U4155 ( .B1(n3298), .B2(n3297), .A(n3296), .ZN(n3301) );
  NAND2_X1 U4156 ( .A1(n3299), .A2(n3602), .ZN(n4727) );
  NAND3_X1 U4157 ( .A1(n4728), .A2(n4727), .A3(n4290), .ZN(n3300) );
  OAI211_X1 U4158 ( .C1(n4731), .C2(n4663), .A(n3301), .B(n3300), .ZN(U3283)
         );
  XOR2_X1 U4159 ( .A(n3303), .B(n3302), .Z(n3304) );
  XNOR2_X1 U4160 ( .A(n3305), .B(n3304), .ZN(n3311) );
  AOI22_X1 U4161 ( .A1(n3361), .A2(n4523), .B1(n4527), .B2(n3742), .ZN(n3310)
         );
  NOR2_X1 U4162 ( .A1(STATE_REG_SCAN_IN), .A2(n3306), .ZN(n4555) );
  NOR2_X1 U4163 ( .A1(n4543), .A2(n3307), .ZN(n3308) );
  AOI211_X1 U4164 ( .C1(n3570), .C2(n4433), .A(n4555), .B(n3308), .ZN(n3309)
         );
  OAI211_X1 U4165 ( .C1(n3311), .C2(n3584), .A(n3310), .B(n3309), .ZN(U3218)
         );
  INV_X1 U4166 ( .A(n3610), .ZN(n3617) );
  NAND2_X1 U4167 ( .A1(n3617), .A2(n3606), .ZN(n3686) );
  XNOR2_X1 U4168 ( .A(n3312), .B(n3686), .ZN(n3313) );
  NAND2_X1 U4169 ( .A1(n3313), .A2(n4421), .ZN(n3397) );
  XOR2_X1 U4170 ( .A(n3314), .B(n3686), .Z(n3400) );
  NAND2_X1 U4171 ( .A1(n3400), .A2(n4290), .ZN(n3324) );
  NAND2_X1 U4172 ( .A1(n3356), .A2(n3395), .ZN(n3315) );
  NAND2_X1 U4173 ( .A1(n3375), .A2(n3315), .ZN(n3405) );
  INV_X1 U4174 ( .A(n3405), .ZN(n3322) );
  AOI22_X1 U4175 ( .A1(n4282), .A2(n3441), .B1(n4279), .B2(n3395), .ZN(n3316)
         );
  OAI21_X1 U4176 ( .B1(n3318), .B2(n3317), .A(n3316), .ZN(n3321) );
  OAI22_X1 U4177 ( .A1(n3351), .A2(n4647), .B1(n3319), .B2(n4022), .ZN(n3320)
         );
  AOI211_X1 U4178 ( .C1(n3322), .C2(n4657), .A(n3321), .B(n3320), .ZN(n3323)
         );
  OAI211_X1 U4179 ( .C1(n4663), .C2(n3397), .A(n3324), .B(n3323), .ZN(U3281)
         );
  INV_X1 U4180 ( .A(n3339), .ZN(n3347) );
  NAND2_X1 U4181 ( .A1(n3325), .A2(REG1_REG_13__SCAN_IN), .ZN(n3327) );
  NAND2_X1 U4182 ( .A1(n3328), .A2(n3329), .ZN(n3330) );
  NAND2_X1 U4183 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4607), .ZN(n4606) );
  NAND2_X1 U4184 ( .A1(n3330), .A2(n4606), .ZN(n3333) );
  NAND2_X1 U4185 ( .A1(n3339), .A2(REG1_REG_15__SCAN_IN), .ZN(n3783) );
  INV_X1 U4186 ( .A(n3783), .ZN(n3331) );
  AOI21_X1 U4187 ( .B1(n4379), .B2(n3347), .A(n3331), .ZN(n3332) );
  OAI211_X1 U4188 ( .C1(n3333), .C2(n3332), .A(n4637), .B(n3782), .ZN(n3346)
         );
  AND2_X1 U4189 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n3581) );
  OAI21_X1 U4190 ( .B1(n3336), .B2(n3335), .A(n3334), .ZN(n3337) );
  NOR2_X1 U4191 ( .A1(n4704), .A2(n3337), .ZN(n3338) );
  INV_X1 U4192 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4603) );
  XNOR2_X1 U4193 ( .A(n4704), .B(n3337), .ZN(n4602) );
  NOR2_X1 U4194 ( .A1(n4603), .A2(n4602), .ZN(n4601) );
  NOR2_X1 U4195 ( .A1(n3338), .A2(n4601), .ZN(n3343) );
  NAND2_X1 U4196 ( .A1(n3339), .A2(REG2_REG_15__SCAN_IN), .ZN(n3792) );
  OR2_X1 U4197 ( .A1(n3339), .A2(REG2_REG_15__SCAN_IN), .ZN(n3340) );
  NAND2_X1 U4198 ( .A1(n3792), .A2(n3340), .ZN(n3342) );
  INV_X1 U4199 ( .A(n3793), .ZN(n3341) );
  AOI211_X1 U4200 ( .C1(n3343), .C2(n3342), .A(n3341), .B(n4630), .ZN(n3344)
         );
  AOI211_X1 U4201 ( .C1(n4635), .C2(ADDR_REG_15__SCAN_IN), .A(n3581), .B(n3344), .ZN(n3345) );
  OAI211_X1 U4202 ( .C1(n4641), .C2(n3347), .A(n3346), .B(n3345), .ZN(U3255)
         );
  INV_X1 U4203 ( .A(n3386), .ZN(n3348) );
  AOI21_X1 U4204 ( .B1(n3350), .B2(n3349), .A(n3348), .ZN(n3355) );
  AOI22_X1 U4205 ( .A1(n3395), .A2(n3569), .B1(n4527), .B2(n3441), .ZN(n3354)
         );
  AND2_X1 U4206 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4566) );
  NOR2_X1 U4207 ( .A1(n4543), .A2(n3351), .ZN(n3352) );
  AOI211_X1 U4208 ( .C1(n3570), .C2(n4416), .A(n4566), .B(n3352), .ZN(n3353)
         );
  OAI211_X1 U4209 ( .C1(n3355), .C2(n3584), .A(n3354), .B(n3353), .ZN(U3228)
         );
  OAI21_X1 U4210 ( .B1(n3358), .B2(n3357), .A(n3356), .ZN(n4655) );
  NAND2_X1 U4211 ( .A1(n3605), .A2(n3616), .ZN(n3675) );
  XNOR2_X1 U4212 ( .A(n3359), .B(n3675), .ZN(n3364) );
  INV_X1 U4213 ( .A(n3364), .ZN(n4659) );
  XNOR2_X1 U4214 ( .A(n3360), .B(n3675), .ZN(n3367) );
  AOI22_X1 U4215 ( .A1(n3742), .A2(n4434), .B1(n4412), .B2(n3361), .ZN(n3362)
         );
  OAI21_X1 U4216 ( .B1(n3363), .B2(n4429), .A(n3362), .ZN(n3366) );
  NOR2_X1 U4217 ( .A1(n3364), .A2(n4419), .ZN(n3365) );
  AOI211_X1 U4218 ( .C1(n4421), .C2(n3367), .A(n3366), .B(n3365), .ZN(n4662)
         );
  INV_X1 U4219 ( .A(n4662), .ZN(n3368) );
  AOI21_X1 U4220 ( .B1(n4724), .B2(n4659), .A(n3368), .ZN(n3370) );
  MUX2_X1 U4221 ( .A(n2411), .B(n3370), .S(n4733), .Z(n3369) );
  OAI21_X1 U4222 ( .B1(n4655), .B2(n4511), .A(n3369), .ZN(U3483) );
  MUX2_X1 U4223 ( .A(n2410), .B(n3370), .S(n4739), .Z(n3371) );
  OAI21_X1 U4224 ( .B1(n4655), .B2(n4440), .A(n3371), .ZN(U3526) );
  NAND2_X1 U4225 ( .A1(n3621), .A2(n3623), .ZN(n3683) );
  XOR2_X1 U4226 ( .A(n3683), .B(n3372), .Z(n4436) );
  XNOR2_X1 U4227 ( .A(n3373), .B(n3683), .ZN(n3374) );
  NOR2_X1 U4228 ( .A1(n3374), .A2(n4115), .ZN(n4431) );
  NAND2_X1 U4229 ( .A1(n3375), .A2(n3387), .ZN(n3376) );
  NAND2_X1 U4230 ( .A1(n4404), .A2(n3376), .ZN(n4512) );
  INV_X1 U4231 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3377) );
  OAI22_X1 U4232 ( .A1(n4022), .A2(n3377), .B1(n3389), .B2(n4647), .ZN(n3378)
         );
  AOI21_X1 U4233 ( .B1(n4280), .B2(n4281), .A(n3378), .ZN(n3380) );
  AOI22_X1 U4234 ( .A1(n4282), .A2(n4433), .B1(n4279), .B2(n3387), .ZN(n3379)
         );
  OAI211_X1 U4235 ( .C1(n4512), .C2(n4643), .A(n3380), .B(n3379), .ZN(n3381)
         );
  AOI21_X1 U4236 ( .B1(n4431), .B2(n4022), .A(n3381), .ZN(n3382) );
  OAI21_X1 U4237 ( .B1(n4436), .B2(n4064), .A(n3382), .ZN(U3280) );
  NAND2_X1 U4238 ( .A1(n3383), .A2(n4538), .ZN(n3394) );
  AOI21_X1 U4239 ( .B1(n3386), .B2(n3385), .A(n3384), .ZN(n3393) );
  AOI22_X1 U4240 ( .A1(n3387), .A2(n4523), .B1(n4525), .B2(n4281), .ZN(n3392)
         );
  INV_X1 U4241 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3388) );
  NOR2_X1 U4242 ( .A1(STATE_REG_SCAN_IN), .A2(n3388), .ZN(n4576) );
  NOR2_X1 U4243 ( .A1(n4543), .A2(n3389), .ZN(n3390) );
  AOI211_X1 U4244 ( .C1(n4527), .C2(n4433), .A(n4576), .B(n3390), .ZN(n3391)
         );
  OAI211_X1 U4245 ( .C1(n3394), .C2(n3393), .A(n3392), .B(n3391), .ZN(U3214)
         );
  AOI22_X1 U4246 ( .A1(n4416), .A2(n4414), .B1(n4412), .B2(n3395), .ZN(n3396)
         );
  OAI211_X1 U4247 ( .C1(n3398), .C2(n4397), .A(n3397), .B(n3396), .ZN(n3399)
         );
  AOI21_X1 U4248 ( .B1(n3400), .B2(n4726), .A(n3399), .ZN(n3403) );
  MUX2_X1 U4249 ( .A(n3401), .B(n3403), .S(n4733), .Z(n3402) );
  OAI21_X1 U4250 ( .B1(n3405), .B2(n4511), .A(n3402), .ZN(U3485) );
  MUX2_X1 U4251 ( .A(n4186), .B(n3403), .S(n4739), .Z(n3404) );
  OAI21_X1 U4252 ( .B1(n4440), .B2(n3405), .A(n3404), .ZN(U3527) );
  NAND2_X1 U4253 ( .A1(n3407), .A2(n3406), .ZN(n3409) );
  XOR2_X1 U4254 ( .A(n3409), .B(n3408), .Z(n3413) );
  AOI22_X1 U4255 ( .A1(n4413), .A2(n3569), .B1(n4525), .B2(n4415), .ZN(n3412)
         );
  INV_X1 U4256 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4191) );
  NOR2_X1 U4257 ( .A1(STATE_REG_SCAN_IN), .A2(n4191), .ZN(n4587) );
  NOR2_X1 U4258 ( .A1(n4543), .A2(n4648), .ZN(n3410) );
  AOI211_X1 U4259 ( .C1(n4527), .C2(n4416), .A(n4587), .B(n3410), .ZN(n3411)
         );
  OAI211_X1 U4260 ( .C1(n3413), .C2(n3584), .A(n3412), .B(n3411), .ZN(U3233)
         );
  XNOR2_X1 U4261 ( .A(n3543), .B(n3415), .ZN(n3416) );
  XNOR2_X1 U4262 ( .A(n3414), .B(n3416), .ZN(n3421) );
  AOI22_X1 U4263 ( .A1(n4394), .A2(n3569), .B1(n4525), .B2(n4395), .ZN(n3420)
         );
  INV_X1 U4264 ( .A(n4276), .ZN(n3418) );
  NAND2_X1 U4265 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4594) );
  OAI21_X1 U4266 ( .B1(n3572), .B2(n4430), .A(n4594), .ZN(n3417) );
  AOI21_X1 U4267 ( .B1(n3418), .B2(n3574), .A(n3417), .ZN(n3419) );
  OAI211_X1 U4268 ( .C1(n3421), .C2(n3584), .A(n3420), .B(n3419), .ZN(U3221)
         );
  NOR2_X1 U4269 ( .A1(n2065), .A2(n3422), .ZN(n3423) );
  XNOR2_X1 U4270 ( .A(n3424), .B(n3423), .ZN(n3428) );
  AOI22_X1 U4271 ( .A1(n4009), .A2(n3569), .B1(n4525), .B2(n4010), .ZN(n3427)
         );
  INV_X1 U4272 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4161) );
  NOR2_X1 U4273 ( .A1(STATE_REG_SCAN_IN), .A2(n4161), .ZN(n4634) );
  NOR2_X1 U4274 ( .A1(n4543), .A2(n4019), .ZN(n3425) );
  AOI211_X1 U4275 ( .C1(n4527), .C2(n4524), .A(n4634), .B(n3425), .ZN(n3426)
         );
  OAI211_X1 U4276 ( .C1(n3428), .C2(n3584), .A(n3427), .B(n3426), .ZN(U3235)
         );
  XNOR2_X1 U4277 ( .A(n3430), .B(n3429), .ZN(n3437) );
  AOI22_X1 U4278 ( .A1(n3848), .A2(n3570), .B1(n4302), .B2(n3569), .ZN(n3436)
         );
  INV_X1 U4279 ( .A(n3431), .ZN(n3849) );
  OAI22_X1 U4280 ( .A1(n3572), .A2(n3433), .B1(STATE_REG_SCAN_IN), .B2(n3432), 
        .ZN(n3434) );
  AOI21_X1 U4281 ( .B1(n3849), .B2(n3574), .A(n3434), .ZN(n3435) );
  OAI211_X1 U4282 ( .C1(n3440), .C2(n3439), .A(n3438), .B(n4538), .ZN(n3450)
         );
  AOI22_X1 U4283 ( .A1(n3442), .A2(n3569), .B1(n4525), .B2(n3441), .ZN(n3449)
         );
  INV_X1 U4284 ( .A(n3443), .ZN(n3447) );
  OAI21_X1 U4285 ( .B1(n3572), .B2(n3445), .A(n3444), .ZN(n3446) );
  AOI21_X1 U4286 ( .B1(n3447), .B2(n3574), .A(n3446), .ZN(n3448) );
  NAND3_X1 U4287 ( .A1(n3450), .A2(n3449), .A3(n3448), .ZN(U3210) );
  INV_X1 U4288 ( .A(n3451), .ZN(n3453) );
  XNOR2_X1 U4289 ( .A(n3453), .B(n3452), .ZN(n3454) );
  XNOR2_X1 U4290 ( .A(n3455), .B(n3454), .ZN(n3460) );
  NAND2_X1 U4291 ( .A1(n4525), .A2(n4526), .ZN(n3456) );
  NAND2_X1 U4292 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4600) );
  OAI211_X1 U4293 ( .C1(n4543), .C2(n4093), .A(n3456), .B(n4600), .ZN(n3458)
         );
  INV_X1 U4294 ( .A(n4395), .ZN(n4383) );
  NOR2_X1 U4295 ( .A1(n3572), .A2(n4383), .ZN(n3457) );
  AOI211_X1 U4296 ( .C1(n4381), .C2(n4523), .A(n3458), .B(n3457), .ZN(n3459)
         );
  OAI21_X1 U4297 ( .B1(n3460), .B2(n3584), .A(n3459), .ZN(U3212) );
  NAND2_X1 U4298 ( .A1(n3554), .A2(n3461), .ZN(n3517) );
  INV_X1 U4299 ( .A(n3517), .ZN(n3465) );
  AOI21_X1 U4300 ( .B1(n3554), .B2(n3463), .A(n3462), .ZN(n3464) );
  NOR3_X1 U4301 ( .A1(n3465), .A2(n3464), .A3(n3584), .ZN(n3469) );
  AOI22_X1 U4302 ( .A1(n3922), .A2(n3569), .B1(n4525), .B2(n3880), .ZN(n3467)
         );
  AOI22_X1 U4303 ( .A1(n4527), .A2(n4337), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3466) );
  OAI211_X1 U4304 ( .C1(n3925), .C2(n4543), .A(n3467), .B(n3466), .ZN(n3468)
         );
  OR2_X1 U4305 ( .A1(n3469), .A2(n3468), .ZN(U3213) );
  OAI21_X1 U4306 ( .B1(n3472), .B2(n3471), .A(n3470), .ZN(n3473) );
  NAND2_X1 U4307 ( .A1(n3473), .A2(n4538), .ZN(n3479) );
  AOI22_X1 U4308 ( .A1(n4527), .A2(n3746), .B1(n4525), .B2(n2806), .ZN(n3478)
         );
  MUX2_X1 U4309 ( .A(STATE_REG_SCAN_IN), .B(n4543), .S(n3474), .Z(n3477) );
  NAND2_X1 U4310 ( .A1(n3569), .A2(n3475), .ZN(n3476) );
  NAND4_X1 U4311 ( .A1(n3479), .A2(n3478), .A3(n3477), .A4(n3476), .ZN(U3215)
         );
  XOR2_X1 U4312 ( .A(n3481), .B(n3480), .Z(n3486) );
  AOI22_X1 U4313 ( .A1(n3993), .A2(n4523), .B1(n4525), .B2(n3994), .ZN(n3485)
         );
  INV_X1 U4314 ( .A(n3999), .ZN(n3483) );
  NAND2_X1 U4315 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3801) );
  OAI21_X1 U4316 ( .B1(n3572), .B2(n3997), .A(n3801), .ZN(n3482) );
  AOI21_X1 U4317 ( .B1(n3483), .B2(n3574), .A(n3482), .ZN(n3484) );
  OAI211_X1 U4318 ( .C1(n3486), .C2(n3584), .A(n3485), .B(n3484), .ZN(U3216)
         );
  XNOR2_X1 U4319 ( .A(n3488), .B(n3487), .ZN(n3489) );
  XNOR2_X1 U4320 ( .A(n3490), .B(n3489), .ZN(n3496) );
  AOI22_X1 U4321 ( .A1(n4336), .A2(n3569), .B1(n4525), .B2(n4337), .ZN(n3495)
         );
  INV_X1 U4322 ( .A(n3491), .ZN(n3958) );
  OAI22_X1 U4323 ( .A1(n3572), .A2(n4340), .B1(STATE_REG_SCAN_IN), .B2(n3492), 
        .ZN(n3493) );
  AOI21_X1 U4324 ( .B1(n3958), .B2(n3574), .A(n3493), .ZN(n3494) );
  OAI211_X1 U4325 ( .C1(n3496), .C2(n3584), .A(n3495), .B(n3494), .ZN(U3220)
         );
  NAND2_X1 U4326 ( .A1(n3498), .A2(n3497), .ZN(n3500) );
  XOR2_X1 U4327 ( .A(n3500), .B(n3499), .Z(n3506) );
  AOI22_X1 U4328 ( .A1(n3879), .A2(n4523), .B1(n4525), .B2(n4303), .ZN(n3505)
         );
  INV_X1 U4329 ( .A(n3887), .ZN(n3503) );
  OAI22_X1 U4330 ( .A1(n3572), .A2(n3918), .B1(STATE_REG_SCAN_IN), .B2(n3501), 
        .ZN(n3502) );
  AOI21_X1 U4331 ( .B1(n3503), .B2(n3574), .A(n3502), .ZN(n3504) );
  OAI211_X1 U4332 ( .C1(n3506), .C2(n3584), .A(n3505), .B(n3504), .ZN(U3222)
         );
  XNOR2_X1 U4333 ( .A(n3508), .B(n3507), .ZN(n3509) );
  XNOR2_X1 U4334 ( .A(n3510), .B(n3509), .ZN(n3514) );
  AOI22_X1 U4335 ( .A1(n4359), .A2(n3569), .B1(n4525), .B2(n4360), .ZN(n3513)
         );
  AND2_X1 U4336 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4623) );
  NOR2_X1 U4337 ( .A1(n4543), .A2(n4030), .ZN(n3511) );
  AOI211_X1 U4338 ( .C1(n4527), .C2(n4373), .A(n4623), .B(n3511), .ZN(n3512)
         );
  OAI211_X1 U4339 ( .C1(n3514), .C2(n3584), .A(n3513), .B(n3512), .ZN(U3225)
         );
  NAND2_X1 U4340 ( .A1(n3517), .A2(n3516), .ZN(n3518) );
  NAND2_X1 U4341 ( .A1(n3515), .A2(n3518), .ZN(n3519) );
  XOR2_X1 U4342 ( .A(n3520), .B(n3519), .Z(n3527) );
  AOI22_X1 U4343 ( .A1(n3570), .A2(n3900), .B1(n4523), .B2(n4319), .ZN(n3526)
         );
  INV_X1 U4344 ( .A(n3521), .ZN(n3901) );
  INV_X1 U4345 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3522) );
  OAI22_X1 U4346 ( .A1(n3572), .A2(n3523), .B1(STATE_REG_SCAN_IN), .B2(n3522), 
        .ZN(n3524) );
  AOI21_X1 U4347 ( .B1(n3901), .B2(n3574), .A(n3524), .ZN(n3525) );
  OAI211_X1 U4348 ( .C1(n3527), .C2(n3584), .A(n3526), .B(n3525), .ZN(U3226)
         );
  INV_X1 U4349 ( .A(n3528), .ZN(n3533) );
  AOI21_X1 U4350 ( .B1(n3532), .B2(n3530), .A(n3529), .ZN(n3531) );
  AOI21_X1 U4351 ( .B1(n3533), .B2(n3532), .A(n3531), .ZN(n3539) );
  AOI22_X1 U4352 ( .A1(n3977), .A2(n3569), .B1(n4525), .B2(n3969), .ZN(n3538)
         );
  INV_X1 U4353 ( .A(n3978), .ZN(n3536) );
  INV_X1 U4354 ( .A(n4010), .ZN(n3971) );
  OAI22_X1 U4355 ( .A1(n3572), .A2(n3971), .B1(STATE_REG_SCAN_IN), .B2(n3534), 
        .ZN(n3535) );
  AOI21_X1 U4356 ( .B1(n3536), .B2(n3574), .A(n3535), .ZN(n3537) );
  OAI211_X1 U4357 ( .C1(n3539), .C2(n3584), .A(n3538), .B(n3537), .ZN(U3230)
         );
  NAND2_X1 U4358 ( .A1(n3541), .A2(n3540), .ZN(n3548) );
  INV_X1 U4359 ( .A(n3414), .ZN(n3546) );
  OAI21_X1 U4360 ( .B1(n3414), .B2(n3543), .A(n3542), .ZN(n3544) );
  OAI21_X1 U4361 ( .B1(n3546), .B2(n3545), .A(n3544), .ZN(n3547) );
  XOR2_X1 U4362 ( .A(n3548), .B(n3547), .Z(n3553) );
  AOI22_X1 U4363 ( .A1(n3676), .A2(n3569), .B1(n4525), .B2(n4073), .ZN(n3552)
         );
  NOR2_X1 U4364 ( .A1(n4543), .A2(n4104), .ZN(n3549) );
  AOI211_X1 U4365 ( .C1(n4527), .C2(n4415), .A(n3550), .B(n3549), .ZN(n3551)
         );
  OAI211_X1 U4366 ( .C1(n3553), .C2(n3584), .A(n3552), .B(n3551), .ZN(U3231)
         );
  INV_X1 U4367 ( .A(n3554), .ZN(n3555) );
  AOI21_X1 U4368 ( .B1(n3557), .B2(n3556), .A(n3555), .ZN(n3563) );
  AOI22_X1 U4369 ( .A1(n3945), .A2(n3569), .B1(n4525), .B2(n4320), .ZN(n3562)
         );
  INV_X1 U4370 ( .A(n3948), .ZN(n3560) );
  OAI22_X1 U4371 ( .A1(n3572), .A2(n3935), .B1(STATE_REG_SCAN_IN), .B2(n3558), 
        .ZN(n3559) );
  AOI21_X1 U4372 ( .B1(n3560), .B2(n3574), .A(n3559), .ZN(n3561) );
  OAI211_X1 U4373 ( .C1(n3563), .C2(n3584), .A(n3562), .B(n3561), .ZN(U3232)
         );
  INV_X1 U4374 ( .A(n3564), .ZN(n3566) );
  NOR2_X1 U4375 ( .A1(n3566), .A2(n3565), .ZN(n3567) );
  XNOR2_X1 U4376 ( .A(n3568), .B(n3567), .ZN(n3577) );
  AOI22_X1 U4377 ( .A1(n3828), .A2(n3570), .B1(n3863), .B2(n3569), .ZN(n3576)
         );
  OAI22_X1 U4378 ( .A1(n3572), .A2(n4323), .B1(STATE_REG_SCAN_IN), .B2(n3571), 
        .ZN(n3573) );
  AOI21_X1 U4379 ( .B1(n3871), .B2(n3574), .A(n3573), .ZN(n3575) );
  OAI211_X1 U4380 ( .C1(n3577), .C2(n3584), .A(n3576), .B(n3575), .ZN(U3237)
         );
  NAND2_X1 U4381 ( .A1(n3578), .A2(n4533), .ZN(n3579) );
  XOR2_X1 U4382 ( .A(n4534), .B(n3579), .Z(n3585) );
  AOI22_X1 U4383 ( .A1(n4372), .A2(n4523), .B1(n4527), .B2(n4073), .ZN(n3583)
         );
  NOR2_X1 U4384 ( .A1(n4543), .A2(n4074), .ZN(n3580) );
  AOI211_X1 U4385 ( .C1(n4525), .C2(n4373), .A(n3581), .B(n3580), .ZN(n3582)
         );
  OAI211_X1 U4386 ( .C1(n3585), .C2(n3584), .A(n3583), .B(n3582), .ZN(U3238)
         );
  NOR2_X1 U4387 ( .A1(n3664), .A2(n2124), .ZN(n3714) );
  OAI211_X1 U4388 ( .C1(n3588), .C2(n3727), .A(n3587), .B(n3586), .ZN(n3591)
         );
  NAND3_X1 U4389 ( .A1(n3591), .A2(n3590), .A3(n3589), .ZN(n3594) );
  NAND3_X1 U4390 ( .A1(n3594), .A2(n3593), .A3(n3592), .ZN(n3597) );
  NAND3_X1 U4391 ( .A1(n3597), .A2(n3596), .A3(n3595), .ZN(n3599) );
  NAND4_X1 U4392 ( .A1(n3600), .A2(n3599), .A3(n3615), .A4(n3598), .ZN(n3603)
         );
  NAND3_X1 U4393 ( .A1(n3603), .A2(n3602), .A3(n3601), .ZN(n3604) );
  NAND3_X1 U4394 ( .A1(n3604), .A2(n3612), .A3(n3616), .ZN(n3607) );
  AND3_X1 U4395 ( .A1(n3607), .A2(n3606), .A3(n3605), .ZN(n3611) );
  NAND2_X1 U4396 ( .A1(n3609), .A2(n3608), .ZN(n3619) );
  NOR3_X1 U4397 ( .A1(n3611), .A2(n3610), .A3(n3619), .ZN(n3626) );
  INV_X1 U4398 ( .A(n3612), .ZN(n3614) );
  NOR2_X1 U4399 ( .A1(n3614), .A2(n3613), .ZN(n3618) );
  NAND4_X1 U4400 ( .A1(n3618), .A2(n3617), .A3(n3616), .A4(n3615), .ZN(n3622)
         );
  NAND2_X1 U4401 ( .A1(n3619), .A2(n3628), .ZN(n3697) );
  INV_X1 U4402 ( .A(n3697), .ZN(n3620) );
  AOI21_X1 U4403 ( .B1(n3622), .B2(n3621), .A(n3620), .ZN(n3625) );
  OAI211_X1 U4404 ( .C1(n3626), .C2(n3625), .A(n3624), .B(n3623), .ZN(n3632)
         );
  INV_X1 U4405 ( .A(n3627), .ZN(n3629) );
  NAND2_X1 U4406 ( .A1(n4065), .A2(n3628), .ZN(n3698) );
  OAI21_X1 U4407 ( .B1(n3629), .B2(n3698), .A(n3697), .ZN(n3631) );
  INV_X1 U4408 ( .A(n3701), .ZN(n3630) );
  AOI21_X1 U4409 ( .B1(n3632), .B2(n3631), .A(n3630), .ZN(n3634) );
  INV_X1 U4410 ( .A(n3699), .ZN(n3633) );
  OAI211_X1 U4411 ( .C1(n3634), .C2(n3633), .A(n2234), .B(n2230), .ZN(n3636)
         );
  INV_X1 U4412 ( .A(n3635), .ZN(n3703) );
  AOI211_X1 U4413 ( .C1(n3636), .C2(n3704), .A(n3703), .B(n3911), .ZN(n3637)
         );
  NOR2_X1 U4414 ( .A1(n3637), .A2(n3708), .ZN(n3639) );
  OAI21_X1 U4415 ( .B1(n3639), .B2(n3638), .A(n3709), .ZN(n3640) );
  NAND2_X1 U4416 ( .A1(n3714), .A2(n3640), .ZN(n3647) );
  NOR2_X1 U4417 ( .A1(n3866), .A2(n4302), .ZN(n3646) );
  NAND2_X1 U4418 ( .A1(n3827), .A2(n3657), .ZN(n3641) );
  AND2_X1 U4419 ( .A1(n3642), .A2(n3641), .ZN(n3658) );
  INV_X1 U4420 ( .A(n3658), .ZN(n3644) );
  NOR2_X1 U4421 ( .A1(n3644), .A2(n3643), .ZN(n3715) );
  INV_X1 U4422 ( .A(n3715), .ZN(n3645) );
  AOI211_X1 U4423 ( .C1(n3719), .C2(n3647), .A(n3646), .B(n3645), .ZN(n3648)
         );
  INV_X1 U4424 ( .A(n3648), .ZN(n3663) );
  NAND2_X1 U4425 ( .A1(n3650), .A2(n3649), .ZN(n3712) );
  INV_X1 U4426 ( .A(n4296), .ZN(n4299) );
  NAND2_X1 U4427 ( .A1(n4742), .A2(REG2_REG_31__SCAN_IN), .ZN(n3655) );
  INV_X1 U4428 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4292) );
  OR2_X1 U4429 ( .A1(n2360), .A2(n4292), .ZN(n3654) );
  INV_X1 U4430 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4441) );
  OR2_X1 U4431 ( .A1(n3652), .A2(n4441), .ZN(n3653) );
  NAND2_X1 U4432 ( .A1(n3651), .A2(DATAI_31_), .ZN(n3810) );
  NAND2_X1 U4433 ( .A1(n3809), .A2(n3810), .ZN(n3662) );
  OAI21_X1 U4434 ( .B1(n3741), .B2(n4299), .A(n3662), .ZN(n3682) );
  INV_X1 U4435 ( .A(n3682), .ZN(n3656) );
  OAI21_X1 U4436 ( .B1(n3827), .B2(n3657), .A(n3656), .ZN(n3711) );
  AOI21_X1 U4437 ( .B1(n3712), .B2(n3658), .A(n3711), .ZN(n3718) );
  NOR2_X1 U4438 ( .A1(n3809), .A2(n3810), .ZN(n3724) );
  INV_X1 U4439 ( .A(n3724), .ZN(n3661) );
  INV_X1 U4440 ( .A(n3741), .ZN(n3659) );
  NOR2_X1 U4441 ( .A1(n3659), .A2(n4296), .ZN(n3725) );
  INV_X1 U4442 ( .A(n3725), .ZN(n3660) );
  NAND2_X1 U4443 ( .A1(n3661), .A2(n3660), .ZN(n3681) );
  AOI22_X1 U4444 ( .A1(n3663), .A2(n3718), .B1(n3662), .B2(n3681), .ZN(n3731)
         );
  INV_X1 U4445 ( .A(n3664), .ZN(n3665) );
  INV_X1 U4446 ( .A(n3668), .ZN(n3669) );
  INV_X1 U4447 ( .A(n3912), .ZN(n3670) );
  XNOR2_X1 U4448 ( .A(n4010), .B(n3998), .ZN(n3990) );
  NOR4_X1 U4449 ( .A1(n3972), .A2(n3957), .A3(n4008), .A4(n3990), .ZN(n3671)
         );
  NAND3_X1 U4450 ( .A1(n3877), .A2(n3897), .A3(n3671), .ZN(n3696) );
  NOR4_X1 U4451 ( .A1(n3673), .A2(n3941), .A3(n3672), .A4(n4069), .ZN(n3678)
         );
  NOR4_X1 U4452 ( .A1(n4055), .A2(n4088), .A3(n3675), .A4(n3674), .ZN(n3677)
         );
  XNOR2_X1 U4453 ( .A(n4320), .B(n3922), .ZN(n3915) );
  XNOR2_X1 U4454 ( .A(n4395), .B(n3676), .ZN(n4119) );
  NAND4_X1 U4455 ( .A1(n3678), .A2(n3677), .A3(n3915), .A4(n4119), .ZN(n3692)
         );
  NAND2_X1 U4456 ( .A1(n3680), .A2(n3679), .ZN(n3860) );
  NAND2_X1 U4457 ( .A1(n4111), .A2(n4109), .ZN(n4285) );
  NOR4_X1 U4458 ( .A1(n4285), .A2(n3683), .A3(n3682), .A4(n3681), .ZN(n3690)
         );
  NAND2_X1 U4459 ( .A1(n2230), .A2(n3985), .ZN(n4028) );
  NOR4_X1 U4460 ( .A1(n3687), .A2(n4028), .A3(n3686), .A4(n2842), .ZN(n3688)
         );
  NAND4_X1 U4461 ( .A1(n3860), .A2(n3690), .A3(n3689), .A4(n3688), .ZN(n3691)
         );
  OR3_X1 U4462 ( .A1(n3693), .A2(n3692), .A3(n3691), .ZN(n3695) );
  NOR4_X1 U4463 ( .A1(n3696), .A2(n3695), .A3(n3842), .A4(n3694), .ZN(n3729)
         );
  INV_X1 U4464 ( .A(n3810), .ZN(n3726) );
  OAI21_X1 U4465 ( .B1(n4085), .B2(n3698), .A(n3697), .ZN(n3700) );
  NAND2_X1 U4466 ( .A1(n3700), .A2(n3699), .ZN(n3702) );
  NAND4_X1 U4467 ( .A1(n3702), .A2(n2234), .A3(n3701), .A4(n2230), .ZN(n3705)
         );
  AOI21_X1 U4468 ( .B1(n3705), .B2(n3704), .A(n3703), .ZN(n3707) );
  OAI21_X1 U4469 ( .B1(n3708), .B2(n3707), .A(n3706), .ZN(n3710) );
  NAND2_X1 U4470 ( .A1(n3710), .A2(n3709), .ZN(n3713) );
  NAND2_X1 U4471 ( .A1(n3716), .A2(n3715), .ZN(n3717) );
  AOI22_X1 U4472 ( .A1(n3720), .A2(n3719), .B1(n3718), .B2(n3717), .ZN(n3721)
         );
  AOI21_X1 U4473 ( .B1(n4296), .B2(n3722), .A(n3721), .ZN(n3723) );
  AOI211_X1 U4474 ( .C1(n3726), .C2(n3725), .A(n3724), .B(n3723), .ZN(n3728)
         );
  MUX2_X1 U4475 ( .A(n3729), .B(n3728), .S(n3727), .Z(n3730) );
  MUX2_X1 U4476 ( .A(n3731), .B(n3730), .S(n4514), .Z(n3733) );
  XNOR2_X1 U4477 ( .A(n3733), .B(n3732), .ZN(n3740) );
  NOR2_X1 U4478 ( .A1(n3735), .A2(n3734), .ZN(n3738) );
  OAI21_X1 U4479 ( .B1(n3739), .B2(n3736), .A(B_REG_SCAN_IN), .ZN(n3737) );
  OAI22_X1 U4480 ( .A1(n3740), .A2(n3739), .B1(n3738), .B2(n3737), .ZN(U3239)
         );
  MUX2_X1 U4481 ( .A(DATAO_REG_31__SCAN_IN), .B(n3809), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4482 ( .A(n3741), .B(DATAO_REG_30__SCAN_IN), .S(n3747), .Z(U3580)
         );
  MUX2_X1 U4483 ( .A(n3827), .B(DATAO_REG_29__SCAN_IN), .S(n3747), .Z(U3579)
         );
  MUX2_X1 U4484 ( .A(DATAO_REG_28__SCAN_IN), .B(n3848), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4485 ( .A(n3828), .B(DATAO_REG_27__SCAN_IN), .S(n3747), .Z(U3577)
         );
  MUX2_X1 U4486 ( .A(n4303), .B(DATAO_REG_26__SCAN_IN), .S(n3747), .Z(U3576)
         );
  MUX2_X1 U4487 ( .A(n3900), .B(DATAO_REG_25__SCAN_IN), .S(n3747), .Z(U3575)
         );
  MUX2_X1 U4488 ( .A(n4320), .B(DATAO_REG_23__SCAN_IN), .S(n3747), .Z(U3573)
         );
  MUX2_X1 U4489 ( .A(n4337), .B(DATAO_REG_22__SCAN_IN), .S(n3747), .Z(U3572)
         );
  MUX2_X1 U4490 ( .A(DATAO_REG_21__SCAN_IN), .B(n3969), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4491 ( .A(n3994), .B(DATAO_REG_20__SCAN_IN), .S(n3747), .Z(U3570)
         );
  MUX2_X1 U4492 ( .A(n4010), .B(DATAO_REG_19__SCAN_IN), .S(n3747), .Z(U3569)
         );
  MUX2_X1 U4493 ( .A(DATAO_REG_18__SCAN_IN), .B(n4360), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4494 ( .A(DATAO_REG_17__SCAN_IN), .B(n4524), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4495 ( .A(DATAO_REG_14__SCAN_IN), .B(n4073), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4496 ( .A(n4395), .B(DATAO_REG_13__SCAN_IN), .S(n3747), .Z(U3563)
         );
  MUX2_X1 U4497 ( .A(n4415), .B(DATAO_REG_12__SCAN_IN), .S(n3747), .Z(U3562)
         );
  MUX2_X1 U4498 ( .A(DATAO_REG_11__SCAN_IN), .B(n4281), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4499 ( .A(n4433), .B(DATAO_REG_9__SCAN_IN), .S(n3747), .Z(U3559) );
  MUX2_X1 U4500 ( .A(DATAO_REG_7__SCAN_IN), .B(n3742), .S(U4043), .Z(U3557) );
  MUX2_X1 U4501 ( .A(n3743), .B(DATAO_REG_6__SCAN_IN), .S(n3747), .Z(U3556) );
  MUX2_X1 U4502 ( .A(DATAO_REG_5__SCAN_IN), .B(n3744), .S(U4043), .Z(U3555) );
  MUX2_X1 U4503 ( .A(DATAO_REG_4__SCAN_IN), .B(n2806), .S(U4043), .Z(U3554) );
  MUX2_X1 U4504 ( .A(n3745), .B(DATAO_REG_3__SCAN_IN), .S(n3747), .Z(U3553) );
  MUX2_X1 U4505 ( .A(DATAO_REG_2__SCAN_IN), .B(n3746), .S(U4043), .Z(U3552) );
  MUX2_X1 U4506 ( .A(DATAO_REG_1__SCAN_IN), .B(n2799), .S(U4043), .Z(U3551) );
  MUX2_X1 U4507 ( .A(n3748), .B(DATAO_REG_0__SCAN_IN), .S(n3747), .Z(U3550) );
  NAND2_X1 U4508 ( .A1(n3760), .A2(n4519), .ZN(n3758) );
  OAI211_X1 U4509 ( .C1(n2967), .C2(n3751), .A(n4591), .B(n3750), .ZN(n3757)
         );
  OAI211_X1 U4510 ( .C1(n3754), .C2(n3753), .A(n4637), .B(n3752), .ZN(n3756)
         );
  AOI22_X1 U4511 ( .A1(n4635), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3755) );
  NAND4_X1 U4512 ( .A1(n3758), .A2(n3757), .A3(n3756), .A4(n3755), .ZN(U3241)
         );
  NAND2_X1 U4513 ( .A1(n3760), .A2(n3759), .ZN(n3769) );
  OAI211_X1 U4514 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3762), .A(n4637), .B(n3761), 
        .ZN(n3768) );
  AOI22_X1 U4515 ( .A1(n4635), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3767) );
  XNOR2_X1 U4516 ( .A(n3764), .B(n3763), .ZN(n3765) );
  NAND2_X1 U4517 ( .A1(n4591), .A2(n3765), .ZN(n3766) );
  NAND4_X1 U4518 ( .A1(n3769), .A2(n3768), .A3(n3767), .A4(n3766), .ZN(U3243)
         );
  NOR2_X1 U4519 ( .A1(n4641), .A2(n3770), .ZN(n3771) );
  AOI211_X1 U4520 ( .C1(n4635), .C2(ADDR_REG_5__SCAN_IN), .A(n3772), .B(n3771), 
        .ZN(n3781) );
  OAI211_X1 U4521 ( .C1(n3775), .C2(n3774), .A(n4637), .B(n3773), .ZN(n3780)
         );
  OAI211_X1 U4522 ( .C1(n3778), .C2(n3777), .A(n4591), .B(n3776), .ZN(n3779)
         );
  NAND3_X1 U4523 ( .A1(n3781), .A2(n3780), .A3(n3779), .ZN(U3245) );
  INV_X1 U4524 ( .A(n4637), .ZN(n3807) );
  MUX2_X1 U4525 ( .A(REG1_REG_19__SCAN_IN), .B(n4354), .S(n3802), .Z(n3789) );
  INV_X1 U4526 ( .A(n3797), .ZN(n4698) );
  AOI22_X1 U4527 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3797), .B1(n4698), .B2(
        n3787), .ZN(n4639) );
  NOR2_X1 U4528 ( .A1(n4699), .A2(REG1_REG_17__SCAN_IN), .ZN(n3786) );
  NOR2_X1 U4529 ( .A1(n3794), .A2(n3784), .ZN(n3785) );
  NOR2_X1 U4530 ( .A1(n3785), .A2(n4616), .ZN(n4625) );
  AOI22_X1 U4531 ( .A1(n4699), .A2(n4366), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4629), .ZN(n4624) );
  XOR2_X1 U4532 ( .A(n3789), .B(n3788), .Z(n3806) );
  INV_X1 U4533 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4534 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4698), .B1(n3797), .B2(
        n3790), .ZN(n4633) );
  NOR2_X1 U4535 ( .A1(n4699), .A2(REG2_REG_17__SCAN_IN), .ZN(n3791) );
  AOI21_X1 U4536 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4699), .A(n3791), .ZN(n4621) );
  INV_X1 U4537 ( .A(n3794), .ZN(n4702) );
  NAND2_X1 U4538 ( .A1(n3795), .A2(n4702), .ZN(n3796) );
  INV_X1 U4539 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4610) );
  OAI21_X1 U4540 ( .B1(n4699), .B2(REG2_REG_17__SCAN_IN), .A(n4620), .ZN(n4632) );
  AOI21_X1 U4541 ( .B1(REG2_REG_18__SCAN_IN), .B2(n3797), .A(n4631), .ZN(n3799) );
  INV_X1 U4542 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4170) );
  MUX2_X1 U4543 ( .A(n4170), .B(REG2_REG_19__SCAN_IN), .S(n3802), .Z(n3798) );
  XNOR2_X1 U4544 ( .A(n3799), .B(n3798), .ZN(n3804) );
  NAND2_X1 U4545 ( .A1(n4635), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3800) );
  OAI211_X1 U4546 ( .C1(n4641), .C2(n3802), .A(n3801), .B(n3800), .ZN(n3803)
         );
  AOI21_X1 U4547 ( .B1(n3804), .B2(n4591), .A(n3803), .ZN(n3805) );
  OAI21_X1 U4548 ( .B1(n3807), .B2(n3806), .A(n3805), .ZN(U3259) );
  XNOR2_X1 U4549 ( .A(n4295), .B(n3810), .ZN(n4445) );
  NAND2_X1 U4550 ( .A1(n3809), .A2(n3808), .ZN(n4298) );
  OAI21_X1 U4551 ( .B1(n3810), .B2(n4428), .A(n4298), .ZN(n4443) );
  NAND2_X1 U4552 ( .A1(n4443), .A2(n4022), .ZN(n3812) );
  NAND2_X1 U4553 ( .A1(n4663), .A2(REG2_REG_31__SCAN_IN), .ZN(n3811) );
  OAI211_X1 U4554 ( .C1(n4445), .C2(n4643), .A(n3812), .B(n3811), .ZN(U3260)
         );
  INV_X1 U4555 ( .A(n3813), .ZN(n3825) );
  INV_X1 U4556 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3814) );
  OAI22_X1 U4557 ( .A1(n4305), .A2(n3815), .B1(n3814), .B2(n4022), .ZN(n3816)
         );
  AOI21_X1 U4558 ( .B1(n3817), .B2(n4279), .A(n3816), .ZN(n3824) );
  INV_X1 U4559 ( .A(n3818), .ZN(n3822) );
  OAI22_X1 U4560 ( .A1(n3820), .A2(n4643), .B1(n3819), .B2(n4647), .ZN(n3821)
         );
  OAI21_X1 U4561 ( .B1(n3822), .B2(n3821), .A(n4022), .ZN(n3823) );
  OAI211_X1 U4562 ( .C1(n3825), .C2(n4064), .A(n3824), .B(n3823), .ZN(U3354)
         );
  INV_X1 U4563 ( .A(n3826), .ZN(n3837) );
  AOI22_X1 U4564 ( .A1(n3828), .A2(n4282), .B1(n3827), .B2(n4280), .ZN(n3832)
         );
  INV_X1 U4565 ( .A(n3829), .ZN(n3830) );
  AOI22_X1 U4566 ( .A1(n3830), .A2(n4653), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4663), .ZN(n3831) );
  OAI211_X1 U4567 ( .C1(n3833), .C2(n4097), .A(n3832), .B(n3831), .ZN(n3836)
         );
  NOR2_X1 U4568 ( .A1(n3834), .A2(n4663), .ZN(n3835) );
  AOI211_X1 U4569 ( .C1(n4657), .C2(n3837), .A(n3836), .B(n3835), .ZN(n3838)
         );
  OAI21_X1 U4570 ( .B1(n3839), .B2(n4064), .A(n3838), .ZN(U3262) );
  XNOR2_X1 U4571 ( .A(n3840), .B(n3842), .ZN(n4308) );
  INV_X1 U4572 ( .A(n4308), .ZN(n3856) );
  NAND2_X1 U4573 ( .A1(n3843), .A2(n3842), .ZN(n3844) );
  AOI21_X1 U4574 ( .B1(n3845), .B2(n3844), .A(n4115), .ZN(n4307) );
  INV_X1 U4575 ( .A(n3846), .ZN(n3847) );
  OAI21_X1 U4576 ( .B1(n3867), .B2(n3852), .A(n3847), .ZN(n4452) );
  NOR2_X1 U4577 ( .A1(n4452), .A2(n4643), .ZN(n3854) );
  AOI22_X1 U4578 ( .A1(n3848), .A2(n4280), .B1(n4282), .B2(n4303), .ZN(n3851)
         );
  AOI22_X1 U4579 ( .A1(n3849), .A2(n4653), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4663), .ZN(n3850) );
  OAI211_X1 U4580 ( .C1(n3852), .C2(n4097), .A(n3851), .B(n3850), .ZN(n3853)
         );
  AOI211_X1 U4581 ( .C1(n4307), .C2(n4022), .A(n3854), .B(n3853), .ZN(n3855)
         );
  OAI21_X1 U4582 ( .B1(n3856), .B2(n4064), .A(n3855), .ZN(U3263) );
  XOR2_X1 U4583 ( .A(n3860), .B(n3857), .Z(n4312) );
  INV_X1 U4584 ( .A(n4312), .ZN(n3875) );
  NAND2_X1 U4585 ( .A1(n3859), .A2(n3858), .ZN(n3861) );
  XNOR2_X1 U4586 ( .A(n3861), .B(n3860), .ZN(n3862) );
  NAND2_X1 U4587 ( .A1(n3862), .A2(n4421), .ZN(n3865) );
  AOI22_X1 U4588 ( .A1(n3900), .A2(n4434), .B1(n3863), .B2(n4412), .ZN(n3864)
         );
  OAI211_X1 U4589 ( .C1(n3866), .C2(n4429), .A(n3865), .B(n3864), .ZN(n4311)
         );
  INV_X1 U4590 ( .A(n3884), .ZN(n3870) );
  INV_X1 U4591 ( .A(n3867), .ZN(n3868) );
  OAI21_X1 U4592 ( .B1(n3870), .B2(n3869), .A(n3868), .ZN(n4456) );
  AOI22_X1 U4593 ( .A1(n4663), .A2(REG2_REG_26__SCAN_IN), .B1(n3871), .B2(
        n4653), .ZN(n3872) );
  OAI21_X1 U4594 ( .B1(n4456), .B2(n4643), .A(n3872), .ZN(n3873) );
  AOI21_X1 U4595 ( .B1(n4311), .B2(n4022), .A(n3873), .ZN(n3874) );
  OAI21_X1 U4596 ( .B1(n3875), .B2(n4064), .A(n3874), .ZN(U3264) );
  XNOR2_X1 U4597 ( .A(n3876), .B(n3877), .ZN(n4316) );
  INV_X1 U4598 ( .A(n4316), .ZN(n3892) );
  XNOR2_X1 U4599 ( .A(n3878), .B(n3877), .ZN(n3883) );
  AOI22_X1 U4600 ( .A1(n3880), .A2(n4434), .B1(n3879), .B2(n4412), .ZN(n3882)
         );
  NAND2_X1 U4601 ( .A1(n4303), .A2(n4414), .ZN(n3881) );
  OAI211_X1 U4602 ( .C1(n3883), .C2(n4115), .A(n3882), .B(n3881), .ZN(n4315)
         );
  INV_X1 U4603 ( .A(n3899), .ZN(n3886) );
  OAI21_X1 U4604 ( .B1(n3886), .B2(n3885), .A(n3884), .ZN(n4460) );
  NOR2_X1 U4605 ( .A1(n4460), .A2(n4643), .ZN(n3890) );
  INV_X1 U4606 ( .A(REG2_REG_25__SCAN_IN), .ZN(n3888) );
  OAI22_X1 U4607 ( .A1(n4022), .A2(n3888), .B1(n3887), .B2(n4647), .ZN(n3889)
         );
  AOI211_X1 U4608 ( .C1(n4315), .C2(n4022), .A(n3890), .B(n3889), .ZN(n3891)
         );
  OAI21_X1 U4609 ( .B1(n3892), .B2(n4064), .A(n3891), .ZN(U3265) );
  NAND2_X1 U4610 ( .A1(n3894), .A2(n3893), .ZN(n3895) );
  XNOR2_X1 U4611 ( .A(n3895), .B(n3897), .ZN(n3896) );
  NAND2_X1 U4612 ( .A1(n3896), .A2(n4421), .ZN(n4322) );
  XNOR2_X1 U4613 ( .A(n3898), .B(n3897), .ZN(n4325) );
  NAND2_X1 U4614 ( .A1(n4325), .A2(n4290), .ZN(n3908) );
  OAI21_X1 U4615 ( .B1(n3923), .B2(n3904), .A(n3899), .ZN(n4464) );
  INV_X1 U4616 ( .A(n4464), .ZN(n3906) );
  AOI22_X1 U4617 ( .A1(n4280), .A2(n3900), .B1(n4282), .B2(n4320), .ZN(n3903)
         );
  AOI22_X1 U4618 ( .A1(n4663), .A2(REG2_REG_24__SCAN_IN), .B1(n3901), .B2(
        n4653), .ZN(n3902) );
  OAI211_X1 U4619 ( .C1(n3904), .C2(n4097), .A(n3903), .B(n3902), .ZN(n3905)
         );
  AOI21_X1 U4620 ( .B1(n3906), .B2(n4657), .A(n3905), .ZN(n3907) );
  OAI211_X1 U4621 ( .C1(n4663), .C2(n4322), .A(n3908), .B(n3907), .ZN(U3266)
         );
  XOR2_X1 U4622 ( .A(n3915), .B(n3909), .Z(n4329) );
  INV_X1 U4623 ( .A(n4329), .ZN(n3930) );
  OR2_X1 U4624 ( .A1(n3910), .A2(n3911), .ZN(n3913) );
  OAI21_X1 U4625 ( .B1(n3931), .B2(n3941), .A(n3914), .ZN(n3916) );
  XOR2_X1 U4626 ( .A(n3916), .B(n3915), .Z(n3921) );
  OAI22_X1 U4627 ( .A1(n3918), .A2(n4429), .B1(n4428), .B2(n3917), .ZN(n3919)
         );
  AOI21_X1 U4628 ( .B1(n4434), .B2(n4337), .A(n3919), .ZN(n3920) );
  OAI21_X1 U4629 ( .B1(n3921), .B2(n4115), .A(n3920), .ZN(n4328) );
  AND2_X1 U4630 ( .A1(n3947), .A2(n3922), .ZN(n3924) );
  OR2_X1 U4631 ( .A1(n3924), .A2(n3923), .ZN(n4468) );
  INV_X1 U4632 ( .A(n3925), .ZN(n3926) );
  AOI22_X1 U4633 ( .A1(n4663), .A2(REG2_REG_23__SCAN_IN), .B1(n3926), .B2(
        n4653), .ZN(n3927) );
  OAI21_X1 U4634 ( .B1(n4468), .B2(n4643), .A(n3927), .ZN(n3928) );
  AOI21_X1 U4635 ( .B1(n4328), .B2(n4022), .A(n3928), .ZN(n3929) );
  OAI21_X1 U4636 ( .B1(n3930), .B2(n4064), .A(n3929), .ZN(U3267) );
  XNOR2_X1 U4637 ( .A(n3931), .B(n3941), .ZN(n3932) );
  NAND2_X1 U4638 ( .A1(n3932), .A2(n4421), .ZN(n3934) );
  AOI22_X1 U4639 ( .A1(n4320), .A2(n4414), .B1(n3945), .B2(n4412), .ZN(n3933)
         );
  OAI211_X1 U4640 ( .C1(n3935), .C2(n4397), .A(n3934), .B(n3933), .ZN(n4332)
         );
  INV_X1 U4641 ( .A(n4332), .ZN(n3954) );
  INV_X1 U4642 ( .A(n3936), .ZN(n3937) );
  NOR2_X1 U4643 ( .A1(n3938), .A2(n3937), .ZN(n3956) );
  OAI21_X1 U4644 ( .B1(n3956), .B2(n3940), .A(n3939), .ZN(n3944) );
  INV_X1 U4645 ( .A(n3941), .ZN(n3943) );
  AOI21_X1 U4646 ( .B1(n3944), .B2(n3943), .A(n3942), .ZN(n4333) );
  NAND2_X1 U4647 ( .A1(n4333), .A2(n4290), .ZN(n3953) );
  NAND2_X1 U4648 ( .A1(n2027), .A2(n3945), .ZN(n3946) );
  NAND2_X1 U4649 ( .A1(n3947), .A2(n3946), .ZN(n4472) );
  INV_X1 U4650 ( .A(n4472), .ZN(n3951) );
  INV_X1 U4651 ( .A(REG2_REG_22__SCAN_IN), .ZN(n3949) );
  OAI22_X1 U4652 ( .A1(n4022), .A2(n3949), .B1(n3948), .B2(n4647), .ZN(n3950)
         );
  AOI21_X1 U4653 ( .B1(n3951), .B2(n4657), .A(n3950), .ZN(n3952) );
  OAI211_X1 U4654 ( .C1(n4663), .C2(n3954), .A(n3953), .B(n3952), .ZN(U3268)
         );
  XNOR2_X1 U4655 ( .A(n3910), .B(n3957), .ZN(n3955) );
  NAND2_X1 U4656 ( .A1(n3955), .A2(n4421), .ZN(n4339) );
  XOR2_X1 U4657 ( .A(n3957), .B(n3956), .Z(n4342) );
  NAND2_X1 U4658 ( .A1(n4342), .A2(n4290), .ZN(n3965) );
  OAI21_X1 U4659 ( .B1(n2077), .B2(n3961), .A(n2027), .ZN(n4476) );
  INV_X1 U4660 ( .A(n4476), .ZN(n3963) );
  AOI22_X1 U4661 ( .A1(n4282), .A2(n3994), .B1(n4280), .B2(n4337), .ZN(n3960)
         );
  AOI22_X1 U4662 ( .A1(n4663), .A2(REG2_REG_21__SCAN_IN), .B1(n3958), .B2(
        n4653), .ZN(n3959) );
  OAI211_X1 U4663 ( .C1(n3961), .C2(n4097), .A(n3960), .B(n3959), .ZN(n3962)
         );
  AOI21_X1 U4664 ( .B1(n3963), .B2(n4657), .A(n3962), .ZN(n3964) );
  OAI211_X1 U4665 ( .C1(n4663), .C2(n4339), .A(n3965), .B(n3964), .ZN(U3269)
         );
  NAND2_X1 U4666 ( .A1(n3967), .A2(n3966), .ZN(n3968) );
  XOR2_X1 U4667 ( .A(n3968), .B(n3972), .Z(n3976) );
  AOI22_X1 U4668 ( .A1(n3969), .A2(n4414), .B1(n4412), .B2(n3977), .ZN(n3970)
         );
  OAI21_X1 U4669 ( .B1(n3971), .B2(n4397), .A(n3970), .ZN(n3975) );
  XNOR2_X1 U4670 ( .A(n3973), .B(n3972), .ZN(n4351) );
  NOR2_X1 U4671 ( .A1(n4351), .A2(n4419), .ZN(n3974) );
  AOI211_X1 U4672 ( .C1(n4421), .C2(n3976), .A(n3975), .B(n3974), .ZN(n4349)
         );
  INV_X1 U4673 ( .A(n4351), .ZN(n3982) );
  NAND2_X1 U4674 ( .A1(n2034), .A2(n3977), .ZN(n4347) );
  AND3_X1 U4675 ( .A1(n4347), .A2(n4657), .A3(n4345), .ZN(n3981) );
  INV_X1 U4676 ( .A(REG2_REG_20__SCAN_IN), .ZN(n3979) );
  OAI22_X1 U4677 ( .A1(n4022), .A2(n3979), .B1(n3978), .B2(n4647), .ZN(n3980)
         );
  AOI211_X1 U4678 ( .C1(n3982), .C2(n4658), .A(n3981), .B(n3980), .ZN(n3983)
         );
  OAI21_X1 U4679 ( .B1(n4349), .B2(n4663), .A(n3983), .ZN(U3270) );
  XNOR2_X1 U4680 ( .A(n3984), .B(n3990), .ZN(n4353) );
  INV_X1 U4681 ( .A(n4353), .ZN(n4003) );
  NAND2_X1 U4682 ( .A1(n3986), .A2(n3985), .ZN(n4007) );
  INV_X1 U4683 ( .A(n3987), .ZN(n3989) );
  OAI21_X1 U4684 ( .B1(n4007), .B2(n3989), .A(n3988), .ZN(n3991) );
  XNOR2_X1 U4685 ( .A(n3991), .B(n3990), .ZN(n3992) );
  NAND2_X1 U4686 ( .A1(n3992), .A2(n4421), .ZN(n3996) );
  AOI22_X1 U4687 ( .A1(n3994), .A2(n4414), .B1(n4412), .B2(n3993), .ZN(n3995)
         );
  OAI211_X1 U4688 ( .C1(n3997), .C2(n4397), .A(n3996), .B(n3995), .ZN(n4352)
         );
  OAI21_X1 U4689 ( .B1(n4014), .B2(n3998), .A(n2034), .ZN(n4481) );
  NOR2_X1 U4690 ( .A1(n4481), .A2(n4643), .ZN(n4001) );
  OAI22_X1 U4691 ( .A1(n4022), .A2(n4170), .B1(n3999), .B2(n4647), .ZN(n4000)
         );
  AOI211_X1 U4692 ( .C1(n4352), .C2(n4022), .A(n4001), .B(n4000), .ZN(n4002)
         );
  OAI21_X1 U4693 ( .B1(n4003), .B2(n4064), .A(n4002), .ZN(U3271) );
  OAI21_X1 U4694 ( .B1(n4005), .B2(n4008), .A(n4004), .ZN(n4006) );
  INV_X1 U4695 ( .A(n4006), .ZN(n4358) );
  XOR2_X1 U4696 ( .A(n4008), .B(n4007), .Z(n4013) );
  AOI22_X1 U4697 ( .A1(n4010), .A2(n4414), .B1(n4009), .B2(n4412), .ZN(n4011)
         );
  OAI21_X1 U4698 ( .B1(n4059), .B2(n4397), .A(n4011), .ZN(n4012) );
  AOI21_X1 U4699 ( .B1(n4013), .B2(n4421), .A(n4012), .ZN(n4357) );
  INV_X1 U4700 ( .A(n4357), .ZN(n4023) );
  INV_X1 U4701 ( .A(n4029), .ZN(n4017) );
  INV_X1 U4702 ( .A(n4014), .ZN(n4015) );
  OAI211_X1 U4703 ( .C1(n4017), .C2(n4016), .A(n4015), .B(n4346), .ZN(n4356)
         );
  NOR2_X1 U4704 ( .A1(n4356), .A2(n4018), .ZN(n4021) );
  OAI22_X1 U4705 ( .A1(n4022), .A2(n3790), .B1(n4019), .B2(n4647), .ZN(n4020)
         );
  AOI211_X1 U4706 ( .C1(n4023), .C2(n4022), .A(n4021), .B(n4020), .ZN(n4024)
         );
  OAI21_X1 U4707 ( .B1(n4358), .B2(n4064), .A(n4024), .ZN(U3272) );
  XNOR2_X1 U4708 ( .A(n4025), .B(n4028), .ZN(n4026) );
  NAND2_X1 U4709 ( .A1(n4026), .A2(n4421), .ZN(n4362) );
  XOR2_X1 U4710 ( .A(n4028), .B(n4027), .Z(n4365) );
  NAND2_X1 U4711 ( .A1(n4365), .A2(n4290), .ZN(n4038) );
  OAI21_X1 U4712 ( .B1(n2073), .B2(n4034), .A(n4029), .ZN(n4486) );
  INV_X1 U4713 ( .A(n4486), .ZN(n4036) );
  AOI22_X1 U4714 ( .A1(n4282), .A2(n4373), .B1(n4280), .B2(n4360), .ZN(n4033)
         );
  INV_X1 U4715 ( .A(n4030), .ZN(n4031) );
  AOI22_X1 U4716 ( .A1(n4663), .A2(REG2_REG_17__SCAN_IN), .B1(n4031), .B2(
        n4653), .ZN(n4032) );
  OAI211_X1 U4717 ( .C1(n4034), .C2(n4097), .A(n4033), .B(n4032), .ZN(n4035)
         );
  AOI21_X1 U4718 ( .B1(n4036), .B2(n4657), .A(n4035), .ZN(n4037) );
  OAI211_X1 U4719 ( .C1(n4663), .C2(n4362), .A(n4038), .B(n4037), .ZN(U3273)
         );
  NAND2_X1 U4720 ( .A1(n4084), .A2(n4088), .ZN(n4083) );
  NAND2_X1 U4721 ( .A1(n4083), .A2(n4039), .ZN(n4041) );
  AND2_X1 U4722 ( .A1(n4041), .A2(n4040), .ZN(n4049) );
  NAND2_X1 U4723 ( .A1(n4083), .A2(n4042), .ZN(n4070) );
  NAND2_X1 U4724 ( .A1(n4070), .A2(n4043), .ZN(n4045) );
  NAND2_X1 U4725 ( .A1(n4045), .A2(n4044), .ZN(n4047) );
  NAND2_X1 U4726 ( .A1(n4047), .A2(n4046), .ZN(n4048) );
  NAND2_X1 U4727 ( .A1(n4049), .A2(n4048), .ZN(n4369) );
  OR2_X1 U4728 ( .A1(n4071), .A2(n4050), .ZN(n4051) );
  NAND2_X1 U4729 ( .A1(n4052), .A2(n4051), .ZN(n4490) );
  INV_X1 U4730 ( .A(n4490), .ZN(n4054) );
  OAI22_X1 U4731 ( .A1(n4022), .A2(n4610), .B1(n4542), .B2(n4647), .ZN(n4053)
         );
  AOI21_X1 U4732 ( .B1(n4054), .B2(n4657), .A(n4053), .ZN(n4063) );
  XNOR2_X1 U4733 ( .A(n4056), .B(n4055), .ZN(n4061) );
  NAND2_X1 U4734 ( .A1(n4522), .A2(n4412), .ZN(n4058) );
  NAND2_X1 U4735 ( .A1(n4526), .A2(n4434), .ZN(n4057) );
  OAI211_X1 U4736 ( .C1(n4059), .C2(n4429), .A(n4058), .B(n4057), .ZN(n4060)
         );
  AOI21_X1 U4737 ( .B1(n4061), .B2(n4421), .A(n4060), .ZN(n4368) );
  OR2_X1 U4738 ( .A1(n4368), .A2(n4663), .ZN(n4062) );
  OAI211_X1 U4739 ( .C1(n4369), .C2(n4064), .A(n4063), .B(n4062), .ZN(U3274)
         );
  NAND2_X1 U4740 ( .A1(n4086), .A2(n4065), .ZN(n4067) );
  INV_X1 U4741 ( .A(n4069), .ZN(n4066) );
  XNOR2_X1 U4742 ( .A(n4067), .B(n4066), .ZN(n4068) );
  NAND2_X1 U4743 ( .A1(n4068), .A2(n4421), .ZN(n4375) );
  XNOR2_X1 U4744 ( .A(n4070), .B(n4069), .ZN(n4378) );
  NAND2_X1 U4745 ( .A1(n4378), .A2(n4290), .ZN(n4082) );
  INV_X1 U4746 ( .A(n4071), .ZN(n4072) );
  OAI21_X1 U4747 ( .B1(n4091), .B2(n4078), .A(n4072), .ZN(n4494) );
  INV_X1 U4748 ( .A(n4494), .ZN(n4080) );
  AOI22_X1 U4749 ( .A1(n4282), .A2(n4073), .B1(n4280), .B2(n4373), .ZN(n4077)
         );
  INV_X1 U4750 ( .A(n4074), .ZN(n4075) );
  AOI22_X1 U4751 ( .A1(n4663), .A2(REG2_REG_15__SCAN_IN), .B1(n4075), .B2(
        n4653), .ZN(n4076) );
  OAI211_X1 U4752 ( .C1(n4078), .C2(n4097), .A(n4077), .B(n4076), .ZN(n4079)
         );
  AOI21_X1 U4753 ( .B1(n4080), .B2(n4657), .A(n4079), .ZN(n4081) );
  OAI211_X1 U4754 ( .C1(n4663), .C2(n4375), .A(n4082), .B(n4081), .ZN(U3275)
         );
  OAI21_X1 U4755 ( .B1(n4084), .B2(n4088), .A(n4083), .ZN(n4386) );
  INV_X1 U4756 ( .A(n4386), .ZN(n4103) );
  INV_X1 U4757 ( .A(n4085), .ZN(n4089) );
  INV_X1 U4758 ( .A(n4086), .ZN(n4087) );
  AOI21_X1 U4759 ( .B1(n4089), .B2(n4088), .A(n4087), .ZN(n4090) );
  OAI22_X1 U4760 ( .A1(n4103), .A2(n4419), .B1(n4115), .B2(n4090), .ZN(n4384)
         );
  NAND2_X1 U4761 ( .A1(n4384), .A2(n4022), .ZN(n4102) );
  INV_X1 U4762 ( .A(n4091), .ZN(n4092) );
  OAI21_X1 U4763 ( .B1(n2075), .B2(n4098), .A(n4092), .ZN(n4498) );
  INV_X1 U4764 ( .A(n4498), .ZN(n4100) );
  AOI22_X1 U4765 ( .A1(n4282), .A2(n4395), .B1(n4280), .B2(n4526), .ZN(n4096)
         );
  INV_X1 U4766 ( .A(n4093), .ZN(n4094) );
  AOI22_X1 U4767 ( .A1(n4663), .A2(REG2_REG_14__SCAN_IN), .B1(n4094), .B2(
        n4653), .ZN(n4095) );
  OAI211_X1 U4768 ( .C1(n4098), .C2(n4097), .A(n4096), .B(n4095), .ZN(n4099)
         );
  AOI21_X1 U4769 ( .B1(n4100), .B2(n4657), .A(n4099), .ZN(n4101) );
  OAI211_X1 U4770 ( .C1(n4103), .C2(n4644), .A(n4102), .B(n4101), .ZN(U3276)
         );
  INV_X1 U4771 ( .A(n4104), .ZN(n4117) );
  INV_X1 U4772 ( .A(n4105), .ZN(n4106) );
  OR2_X1 U4773 ( .A1(n4411), .A2(n4106), .ZN(n4108) );
  NAND2_X1 U4774 ( .A1(n4108), .A2(n4107), .ZN(n4286) );
  INV_X1 U4775 ( .A(n4109), .ZN(n4110) );
  AOI21_X1 U4776 ( .B1(n4286), .B2(n4111), .A(n4110), .ZN(n4112) );
  XOR2_X1 U4777 ( .A(n4119), .B(n4112), .Z(n4116) );
  OAI22_X1 U4778 ( .A1(n4376), .A2(n4429), .B1(n4428), .B2(n4121), .ZN(n4113)
         );
  AOI21_X1 U4779 ( .B1(n4434), .B2(n4415), .A(n4113), .ZN(n4114) );
  OAI21_X1 U4780 ( .B1(n4116), .B2(n4115), .A(n4114), .ZN(n4389) );
  AOI21_X1 U4781 ( .B1(n4117), .B2(n4653), .A(n4389), .ZN(n4126) );
  XOR2_X1 U4782 ( .A(n4119), .B(n4118), .Z(n4390) );
  INV_X1 U4783 ( .A(n4275), .ZN(n4122) );
  OAI21_X1 U4784 ( .B1(n4122), .B2(n4121), .A(n4120), .ZN(n4502) );
  OAI22_X1 U4785 ( .A1(n4502), .A2(n4643), .B1(n4123), .B2(n4022), .ZN(n4124)
         );
  AOI21_X1 U4786 ( .B1(n4390), .B2(n4290), .A(n4124), .ZN(n4125) );
  OAI21_X1 U4787 ( .B1(n4126), .B2(n4663), .A(n4125), .ZN(n4271) );
  INV_X1 U4788 ( .A(keyinput3), .ZN(n4169) );
  NOR3_X1 U4789 ( .A1(keyinput51), .A2(keyinput49), .A3(keyinput1), .ZN(n4130)
         );
  NAND3_X1 U4790 ( .A1(keyinput48), .A2(keyinput33), .A3(keyinput41), .ZN(
        n4128) );
  NAND3_X1 U4791 ( .A1(keyinput23), .A2(keyinput30), .A3(keyinput14), .ZN(
        n4127) );
  NOR4_X1 U4792 ( .A1(keyinput44), .A2(keyinput52), .A3(n4128), .A4(n4127), 
        .ZN(n4129) );
  NAND3_X1 U4793 ( .A1(keyinput17), .A2(n4130), .A3(n4129), .ZN(n4131) );
  NOR4_X1 U4794 ( .A1(keyinput58), .A2(keyinput13), .A3(n4169), .A4(n4131), 
        .ZN(n4154) );
  NAND3_X1 U4795 ( .A1(keyinput57), .A2(keyinput54), .A3(keyinput38), .ZN(
        n4152) );
  NOR2_X1 U4796 ( .A1(keyinput18), .A2(keyinput6), .ZN(n4135) );
  NAND4_X1 U4797 ( .A1(keyinput20), .A2(keyinput7), .A3(keyinput39), .A4(
        keyinput29), .ZN(n4133) );
  NAND2_X1 U4798 ( .A1(keyinput26), .A2(keyinput25), .ZN(n4132) );
  NOR4_X1 U4799 ( .A1(keyinput62), .A2(keyinput61), .A3(n4133), .A4(n4132), 
        .ZN(n4134) );
  NAND4_X1 U4800 ( .A1(keyinput46), .A2(keyinput42), .A3(n4135), .A4(n4134), 
        .ZN(n4151) );
  NAND2_X1 U4801 ( .A1(keyinput10), .A2(keyinput8), .ZN(n4141) );
  NOR2_X1 U4802 ( .A1(keyinput56), .A2(keyinput40), .ZN(n4139) );
  NAND3_X1 U4803 ( .A1(keyinput60), .A2(keyinput11), .A3(keyinput63), .ZN(
        n4137) );
  NAND3_X1 U4804 ( .A1(keyinput0), .A2(keyinput16), .A3(keyinput31), .ZN(n4136) );
  NOR4_X1 U4805 ( .A1(keyinput2), .A2(keyinput21), .A3(n4137), .A4(n4136), 
        .ZN(n4138) );
  NAND4_X1 U4806 ( .A1(keyinput15), .A2(keyinput36), .A3(n4139), .A4(n4138), 
        .ZN(n4140) );
  NOR4_X1 U4807 ( .A1(keyinput47), .A2(keyinput19), .A3(n4141), .A4(n4140), 
        .ZN(n4149) );
  NOR3_X1 U4808 ( .A1(keyinput55), .A2(keyinput50), .A3(keyinput59), .ZN(n4148) );
  NOR2_X1 U4809 ( .A1(keyinput34), .A2(keyinput35), .ZN(n4142) );
  NAND3_X1 U4810 ( .A1(keyinput43), .A2(keyinput32), .A3(n4142), .ZN(n4146) );
  NAND3_X1 U4811 ( .A1(keyinput28), .A2(keyinput4), .A3(keyinput53), .ZN(n4145) );
  INV_X1 U4812 ( .A(keyinput37), .ZN(n4143) );
  NAND4_X1 U4813 ( .A1(keyinput45), .A2(keyinput5), .A3(keyinput9), .A4(n4143), 
        .ZN(n4144) );
  NOR4_X1 U4814 ( .A1(keyinput12), .A2(n4146), .A3(n4145), .A4(n4144), .ZN(
        n4147) );
  NAND4_X1 U4815 ( .A1(n4149), .A2(keyinput22), .A3(n4148), .A4(n4147), .ZN(
        n4150) );
  NOR4_X1 U4816 ( .A1(keyinput27), .A2(n4152), .A3(n4151), .A4(n4150), .ZN(
        n4153) );
  AOI21_X1 U4817 ( .B1(n4154), .B2(n4153), .A(keyinput24), .ZN(n4269) );
  INV_X1 U4818 ( .A(DATAI_23_), .ZN(n4696) );
  INV_X1 U4819 ( .A(keyinput25), .ZN(n4156) );
  OAI22_X1 U4820 ( .A1(n4696), .A2(keyinput61), .B1(n4156), .B2(
        ADDR_REG_18__SCAN_IN), .ZN(n4155) );
  AOI221_X1 U4821 ( .B1(n4696), .B2(keyinput61), .C1(ADDR_REG_18__SCAN_IN), 
        .C2(n4156), .A(n4155), .ZN(n4167) );
  INV_X1 U4822 ( .A(keyinput62), .ZN(n4158) );
  OAI22_X1 U4823 ( .A1(n4159), .A2(keyinput57), .B1(n4158), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4157) );
  AOI221_X1 U4824 ( .B1(n4159), .B2(keyinput57), .C1(DATAO_REG_16__SCAN_IN), 
        .C2(n4158), .A(n4157), .ZN(n4166) );
  OAI22_X1 U4825 ( .A1(n4161), .A2(keyinput54), .B1(n4470), .B2(keyinput38), 
        .ZN(n4160) );
  AOI221_X1 U4826 ( .B1(n4161), .B2(keyinput54), .C1(keyinput38), .C2(n4470), 
        .A(n4160), .ZN(n4165) );
  INV_X1 U4827 ( .A(keyinput27), .ZN(n4163) );
  OAI22_X1 U4828 ( .A1(n4326), .A2(keyinput60), .B1(n4163), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4162) );
  AOI221_X1 U4829 ( .B1(n4326), .B2(keyinput60), .C1(DATAO_REG_24__SCAN_IN), 
        .C2(n4163), .A(n4162), .ZN(n4164) );
  NAND4_X1 U4830 ( .A1(n4167), .A2(n4166), .A3(n4165), .A4(n4164), .ZN(n4182)
         );
  AOI22_X1 U4831 ( .A1(n4170), .A2(keyinput48), .B1(ADDR_REG_19__SCAN_IN), 
        .B2(n4169), .ZN(n4168) );
  OAI221_X1 U4832 ( .B1(n4170), .B2(keyinput48), .C1(n4169), .C2(
        ADDR_REG_19__SCAN_IN), .A(n4168), .ZN(n4181) );
  AOI22_X1 U4833 ( .A1(n3284), .A2(keyinput1), .B1(n2375), .B2(keyinput46), 
        .ZN(n4171) );
  OAI221_X1 U4834 ( .B1(n3284), .B2(keyinput1), .C1(n2375), .C2(keyinput46), 
        .A(n4171), .ZN(n4180) );
  AOI22_X1 U4835 ( .A1(n4670), .A2(keyinput31), .B1(keyinput56), .B2(n4684), 
        .ZN(n4172) );
  OAI221_X1 U4836 ( .B1(n4670), .B2(keyinput31), .C1(n4684), .C2(keyinput56), 
        .A(n4172), .ZN(n4178) );
  AOI22_X1 U4837 ( .A1(n4174), .A2(keyinput4), .B1(n4711), .B2(keyinput12), 
        .ZN(n4173) );
  OAI221_X1 U4838 ( .B1(n4174), .B2(keyinput4), .C1(n4711), .C2(keyinput12), 
        .A(n4173), .ZN(n4177) );
  INV_X1 U4839 ( .A(keyinput51), .ZN(n4175) );
  XNOR2_X1 U4840 ( .A(n4175), .B(ADDR_REG_1__SCAN_IN), .ZN(n4176) );
  OR3_X1 U4841 ( .A1(n4178), .A2(n4177), .A3(n4176), .ZN(n4179) );
  NOR4_X1 U4842 ( .A1(n4182), .A2(n4181), .A3(n4180), .A4(n4179), .ZN(n4217)
         );
  INV_X1 U4843 ( .A(DATAI_9_), .ZN(n4709) );
  AOI22_X1 U4844 ( .A1(n4709), .A2(keyinput16), .B1(n2436), .B2(keyinput21), 
        .ZN(n4183) );
  OAI221_X1 U4845 ( .B1(n4709), .B2(keyinput16), .C1(n2436), .C2(keyinput21), 
        .A(n4183), .ZN(n4196) );
  INV_X1 U4846 ( .A(keyinput29), .ZN(n4185) );
  AOI22_X1 U4847 ( .A1(n4186), .A2(keyinput26), .B1(ADDR_REG_17__SCAN_IN), 
        .B2(n4185), .ZN(n4184) );
  OAI221_X1 U4848 ( .B1(n4186), .B2(keyinput26), .C1(n4185), .C2(
        ADDR_REG_17__SCAN_IN), .A(n4184), .ZN(n4195) );
  INV_X1 U4849 ( .A(keyinput7), .ZN(n4189) );
  INV_X1 U4850 ( .A(keyinput39), .ZN(n4188) );
  AOI22_X1 U4851 ( .A1(n4189), .A2(ADDR_REG_15__SCAN_IN), .B1(
        ADDR_REG_16__SCAN_IN), .B2(n4188), .ZN(n4187) );
  OAI221_X1 U4852 ( .B1(n4189), .B2(ADDR_REG_15__SCAN_IN), .C1(n4188), .C2(
        ADDR_REG_16__SCAN_IN), .A(n4187), .ZN(n4194) );
  AOI22_X1 U4853 ( .A1(n4192), .A2(keyinput30), .B1(n4191), .B2(keyinput14), 
        .ZN(n4190) );
  OAI221_X1 U4854 ( .B1(n4192), .B2(keyinput30), .C1(n4191), .C2(keyinput14), 
        .A(n4190), .ZN(n4193) );
  NOR4_X1 U4855 ( .A1(n4196), .A2(n4195), .A3(n4194), .A4(n4193), .ZN(n4216)
         );
  INV_X1 U4856 ( .A(keyinput6), .ZN(n4199) );
  INV_X1 U4857 ( .A(keyinput20), .ZN(n4198) );
  AOI22_X1 U4858 ( .A1(n4199), .A2(ADDR_REG_13__SCAN_IN), .B1(
        ADDR_REG_14__SCAN_IN), .B2(n4198), .ZN(n4197) );
  OAI221_X1 U4859 ( .B1(n4199), .B2(ADDR_REG_13__SCAN_IN), .C1(n4198), .C2(
        ADDR_REG_14__SCAN_IN), .A(n4197), .ZN(n4203) );
  INV_X1 U4860 ( .A(keyinput42), .ZN(n4201) );
  AOI22_X1 U4861 ( .A1(n3377), .A2(keyinput18), .B1(ADDR_REG_12__SCAN_IN), 
        .B2(n4201), .ZN(n4200) );
  OAI221_X1 U4862 ( .B1(n3377), .B2(keyinput18), .C1(n4201), .C2(
        ADDR_REG_12__SCAN_IN), .A(n4200), .ZN(n4202) );
  NOR2_X1 U4863 ( .A1(n4203), .A2(n4202), .ZN(n4215) );
  INV_X1 U4864 ( .A(keyinput17), .ZN(n4205) );
  AOI22_X1 U4865 ( .A1(n4206), .A2(keyinput49), .B1(ADDR_REG_2__SCAN_IN), .B2(
        n4205), .ZN(n4204) );
  OAI221_X1 U4866 ( .B1(n4206), .B2(keyinput49), .C1(n4205), .C2(
        ADDR_REG_2__SCAN_IN), .A(n4204), .ZN(n4213) );
  AOI22_X1 U4867 ( .A1(n4454), .A2(keyinput11), .B1(n4208), .B2(keyinput2), 
        .ZN(n4207) );
  OAI221_X1 U4868 ( .B1(n4454), .B2(keyinput11), .C1(n4208), .C2(keyinput2), 
        .A(n4207), .ZN(n4212) );
  INV_X1 U4869 ( .A(DATAI_7_), .ZN(n4209) );
  XNOR2_X1 U4870 ( .A(keyinput35), .B(n4209), .ZN(n4211) );
  XNOR2_X1 U4871 ( .A(keyinput47), .B(n4441), .ZN(n4210) );
  NOR4_X1 U4872 ( .A1(n4213), .A2(n4212), .A3(n4211), .A4(n4210), .ZN(n4214)
         );
  NAND4_X1 U4873 ( .A1(n4217), .A2(n4216), .A3(n4215), .A4(n4214), .ZN(n4267)
         );
  INV_X1 U4874 ( .A(IR_REG_25__SCAN_IN), .ZN(n4219) );
  AOI22_X1 U4875 ( .A1(n4220), .A2(keyinput13), .B1(n4219), .B2(keyinput9), 
        .ZN(n4218) );
  OAI221_X1 U4876 ( .B1(n4220), .B2(keyinput13), .C1(n4219), .C2(keyinput9), 
        .A(n4218), .ZN(n4230) );
  AOI22_X1 U4877 ( .A1(n4222), .A2(keyinput63), .B1(n2909), .B2(keyinput10), 
        .ZN(n4221) );
  OAI221_X1 U4878 ( .B1(n4222), .B2(keyinput63), .C1(n2909), .C2(keyinput10), 
        .A(n4221), .ZN(n4229) );
  INV_X1 U4879 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4224) );
  AOI22_X1 U4880 ( .A1(n2359), .A2(keyinput19), .B1(n4224), .B2(keyinput0), 
        .ZN(n4223) );
  OAI221_X1 U4881 ( .B1(n2359), .B2(keyinput19), .C1(n4224), .C2(keyinput0), 
        .A(n4223), .ZN(n4228) );
  INV_X1 U4882 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4547) );
  INV_X1 U4883 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4226) );
  AOI22_X1 U4884 ( .A1(n4547), .A2(keyinput41), .B1(n4226), .B2(keyinput23), 
        .ZN(n4225) );
  OAI221_X1 U4885 ( .B1(n4547), .B2(keyinput41), .C1(n4226), .C2(keyinput23), 
        .A(n4225), .ZN(n4227) );
  NOR4_X1 U4886 ( .A1(n4230), .A2(n4229), .A3(n4228), .A4(n4227), .ZN(n4255)
         );
  XOR2_X1 U4887 ( .A(DATAI_2_), .B(keyinput37), .Z(n4238) );
  XNOR2_X1 U4888 ( .A(DATAI_14_), .B(keyinput22), .ZN(n4234) );
  XNOR2_X1 U4889 ( .A(REG3_REG_21__SCAN_IN), .B(keyinput5), .ZN(n4233) );
  XNOR2_X1 U4890 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput45), .ZN(n4232) );
  XNOR2_X1 U4891 ( .A(IR_REG_4__SCAN_IN), .B(keyinput43), .ZN(n4231) );
  NAND4_X1 U4892 ( .A1(n4234), .A2(n4233), .A3(n4232), .A4(n4231), .ZN(n4237)
         );
  INV_X1 U4893 ( .A(DATAI_18_), .ZN(n4697) );
  XNOR2_X1 U4894 ( .A(n4697), .B(keyinput59), .ZN(n4236) );
  XNOR2_X1 U4895 ( .A(keyinput32), .B(n2258), .ZN(n4235) );
  NOR4_X1 U4896 ( .A1(n4238), .A2(n4237), .A3(n4236), .A4(n4235), .ZN(n4254)
         );
  XNOR2_X1 U4897 ( .A(n4239), .B(keyinput8), .ZN(n4245) );
  XOR2_X1 U4898 ( .A(IR_REG_16__SCAN_IN), .B(keyinput34), .Z(n4244) );
  XNOR2_X1 U4899 ( .A(n4240), .B(keyinput53), .ZN(n4243) );
  XNOR2_X1 U4900 ( .A(n4241), .B(keyinput40), .ZN(n4242) );
  NOR4_X1 U4901 ( .A1(n4245), .A2(n4244), .A3(n4243), .A4(n4242), .ZN(n4253)
         );
  XOR2_X1 U4902 ( .A(IR_REG_26__SCAN_IN), .B(keyinput28), .Z(n4251) );
  XOR2_X1 U4903 ( .A(REG3_REG_2__SCAN_IN), .B(keyinput52), .Z(n4250) );
  XNOR2_X1 U4904 ( .A(n4246), .B(keyinput50), .ZN(n4249) );
  XNOR2_X1 U4905 ( .A(n4247), .B(keyinput55), .ZN(n4248) );
  NOR4_X1 U4906 ( .A1(n4251), .A2(n4250), .A3(n4249), .A4(n4248), .ZN(n4252)
         );
  NAND4_X1 U4907 ( .A1(n4255), .A2(n4254), .A3(n4253), .A4(n4252), .ZN(n4266)
         );
  INV_X1 U4908 ( .A(keyinput33), .ZN(n4258) );
  INV_X1 U4909 ( .A(keyinput44), .ZN(n4257) );
  OAI22_X1 U4910 ( .A1(n4258), .A2(DATAO_REG_10__SCAN_IN), .B1(n4257), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n4256) );
  AOI221_X1 U4911 ( .B1(n4258), .B2(DATAO_REG_10__SCAN_IN), .C1(
        DATAO_REG_15__SCAN_IN), .C2(n4257), .A(n4256), .ZN(n4260) );
  XNOR2_X1 U4912 ( .A(REG2_REG_17__SCAN_IN), .B(keyinput58), .ZN(n4259) );
  OAI211_X1 U4913 ( .C1(keyinput24), .C2(n4261), .A(n4260), .B(n4259), .ZN(
        n4265) );
  OAI22_X1 U4914 ( .A1(n4680), .A2(keyinput15), .B1(n4692), .B2(keyinput36), 
        .ZN(n4262) );
  AOI221_X1 U4915 ( .B1(n4680), .B2(keyinput15), .C1(keyinput36), .C2(n4692), 
        .A(n4262), .ZN(n4263) );
  INV_X1 U4916 ( .A(n4263), .ZN(n4264) );
  NOR4_X1 U4917 ( .A1(n4267), .A2(n4266), .A3(n4265), .A4(n4264), .ZN(n4268)
         );
  OAI21_X1 U4918 ( .B1(n4269), .B2(DATAO_REG_8__SCAN_IN), .A(n4268), .ZN(n4270) );
  XNOR2_X1 U4919 ( .A(n4271), .B(n4270), .ZN(U3277) );
  XNOR2_X1 U4920 ( .A(n4272), .B(n4285), .ZN(n4393) );
  OR2_X1 U4921 ( .A1(n4405), .A2(n4273), .ZN(n4274) );
  NAND2_X1 U4922 ( .A1(n4275), .A2(n4274), .ZN(n4505) );
  INV_X1 U4923 ( .A(REG2_REG_12__SCAN_IN), .ZN(n4277) );
  OAI22_X1 U4924 ( .A1(n4022), .A2(n4277), .B1(n4276), .B2(n4647), .ZN(n4278)
         );
  AOI21_X1 U4925 ( .B1(n4394), .B2(n4279), .A(n4278), .ZN(n4284) );
  AOI22_X1 U4926 ( .A1(n4282), .A2(n4281), .B1(n4280), .B2(n4395), .ZN(n4283)
         );
  OAI211_X1 U4927 ( .C1(n4505), .C2(n4643), .A(n4284), .B(n4283), .ZN(n4289)
         );
  XNOR2_X1 U4928 ( .A(n4286), .B(n4285), .ZN(n4287) );
  NAND2_X1 U4929 ( .A1(n4287), .A2(n4421), .ZN(n4400) );
  NOR2_X1 U4930 ( .A1(n4400), .A2(n4663), .ZN(n4288) );
  AOI211_X1 U4931 ( .C1(n4290), .C2(n4393), .A(n4289), .B(n4288), .ZN(n4291)
         );
  INV_X1 U4932 ( .A(n4291), .ZN(U3278) );
  NOR2_X1 U4933 ( .A1(n4739), .A2(n4292), .ZN(n4293) );
  AOI21_X1 U4934 ( .B1(n4739), .B2(n4443), .A(n4293), .ZN(n4294) );
  OAI21_X1 U4935 ( .B1(n4445), .B2(n4440), .A(n4294), .ZN(U3549) );
  AOI21_X1 U4936 ( .B1(n4296), .B2(n2029), .A(n4295), .ZN(n4545) );
  NAND2_X1 U4937 ( .A1(n4545), .A2(n4297), .ZN(n4301) );
  OAI21_X1 U4938 ( .B1(n4299), .B2(n4428), .A(n4298), .ZN(n4544) );
  NAND2_X1 U4939 ( .A1(n4544), .A2(n4739), .ZN(n4300) );
  OAI211_X1 U4940 ( .C1(n4739), .C2(n2903), .A(n4301), .B(n4300), .ZN(U3548)
         );
  AOI22_X1 U4941 ( .A1(n4303), .A2(n4434), .B1(n4302), .B2(n4412), .ZN(n4304)
         );
  OAI21_X1 U4942 ( .B1(n4305), .B2(n4429), .A(n4304), .ZN(n4306) );
  AOI211_X1 U4943 ( .C1(n4308), .C2(n4726), .A(n4307), .B(n4306), .ZN(n4449)
         );
  MUX2_X1 U4944 ( .A(n4309), .B(n4449), .S(n4739), .Z(n4310) );
  OAI21_X1 U4945 ( .B1(n4440), .B2(n4452), .A(n4310), .ZN(U3545) );
  AOI21_X1 U4946 ( .B1(n4312), .B2(n4726), .A(n4311), .ZN(n4453) );
  MUX2_X1 U4947 ( .A(n4313), .B(n4453), .S(n4739), .Z(n4314) );
  OAI21_X1 U4948 ( .B1(n4440), .B2(n4456), .A(n4314), .ZN(U3544) );
  INV_X1 U4949 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4317) );
  AOI21_X1 U4950 ( .B1(n4316), .B2(n4726), .A(n4315), .ZN(n4457) );
  MUX2_X1 U4951 ( .A(n4317), .B(n4457), .S(n4739), .Z(n4318) );
  OAI21_X1 U4952 ( .B1(n4440), .B2(n4460), .A(n4318), .ZN(U3543) );
  AOI22_X1 U4953 ( .A1(n4320), .A2(n4434), .B1(n4319), .B2(n4412), .ZN(n4321)
         );
  OAI211_X1 U4954 ( .C1(n4323), .C2(n4429), .A(n4322), .B(n4321), .ZN(n4324)
         );
  AOI21_X1 U4955 ( .B1(n4325), .B2(n4726), .A(n4324), .ZN(n4461) );
  MUX2_X1 U4956 ( .A(n4326), .B(n4461), .S(n4739), .Z(n4327) );
  OAI21_X1 U4957 ( .B1(n4440), .B2(n4464), .A(n4327), .ZN(U3542) );
  INV_X1 U4958 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4330) );
  AOI21_X1 U4959 ( .B1(n4329), .B2(n4726), .A(n4328), .ZN(n4465) );
  MUX2_X1 U4960 ( .A(n4330), .B(n4465), .S(n4739), .Z(n4331) );
  OAI21_X1 U4961 ( .B1(n4440), .B2(n4468), .A(n4331), .ZN(U3541) );
  AOI21_X1 U4962 ( .B1(n4333), .B2(n4726), .A(n4332), .ZN(n4469) );
  MUX2_X1 U4963 ( .A(n4334), .B(n4469), .S(n4739), .Z(n4335) );
  OAI21_X1 U4964 ( .B1(n4440), .B2(n4472), .A(n4335), .ZN(U3540) );
  AOI22_X1 U4965 ( .A1(n4337), .A2(n4414), .B1(n4336), .B2(n4412), .ZN(n4338)
         );
  OAI211_X1 U4966 ( .C1(n4340), .C2(n4397), .A(n4339), .B(n4338), .ZN(n4341)
         );
  AOI21_X1 U4967 ( .B1(n4342), .B2(n4726), .A(n4341), .ZN(n4473) );
  MUX2_X1 U4968 ( .A(n4343), .B(n4473), .S(n4739), .Z(n4344) );
  OAI21_X1 U4969 ( .B1(n4440), .B2(n4476), .A(n4344), .ZN(U3539) );
  NAND3_X1 U4970 ( .A1(n4347), .A2(n4346), .A3(n4345), .ZN(n4348) );
  OAI211_X1 U4971 ( .C1(n4351), .C2(n4350), .A(n4349), .B(n4348), .ZN(n4477)
         );
  MUX2_X1 U4972 ( .A(REG1_REG_20__SCAN_IN), .B(n4477), .S(n4739), .Z(U3538) );
  AOI21_X1 U4973 ( .B1(n4353), .B2(n4726), .A(n4352), .ZN(n4478) );
  MUX2_X1 U4974 ( .A(n4354), .B(n4478), .S(n4739), .Z(n4355) );
  OAI21_X1 U4975 ( .B1(n4440), .B2(n4481), .A(n4355), .ZN(U3537) );
  OAI211_X1 U4976 ( .C1(n4358), .C2(n4437), .A(n4357), .B(n4356), .ZN(n4482)
         );
  MUX2_X1 U4977 ( .A(REG1_REG_18__SCAN_IN), .B(n4482), .S(n4739), .Z(U3536) );
  AOI22_X1 U4978 ( .A1(n4360), .A2(n4414), .B1(n4412), .B2(n4359), .ZN(n4361)
         );
  OAI211_X1 U4979 ( .C1(n4363), .C2(n4397), .A(n4362), .B(n4361), .ZN(n4364)
         );
  AOI21_X1 U4980 ( .B1(n4365), .B2(n4726), .A(n4364), .ZN(n4484) );
  MUX2_X1 U4981 ( .A(n4484), .B(n4366), .S(n4737), .Z(n4367) );
  OAI21_X1 U4982 ( .B1(n4440), .B2(n4486), .A(n4367), .ZN(U3535) );
  OAI21_X1 U4983 ( .B1(n4369), .B2(n4437), .A(n4368), .ZN(n4487) );
  MUX2_X1 U4984 ( .A(REG1_REG_16__SCAN_IN), .B(n4487), .S(n4739), .Z(n4370) );
  INV_X1 U4985 ( .A(n4370), .ZN(n4371) );
  OAI21_X1 U4986 ( .B1(n4440), .B2(n4490), .A(n4371), .ZN(U3534) );
  AOI22_X1 U4987 ( .A1(n4373), .A2(n4414), .B1(n4412), .B2(n4372), .ZN(n4374)
         );
  OAI211_X1 U4988 ( .C1(n4376), .C2(n4397), .A(n4375), .B(n4374), .ZN(n4377)
         );
  AOI21_X1 U4989 ( .B1(n4378), .B2(n4726), .A(n4377), .ZN(n4492) );
  MUX2_X1 U4990 ( .A(n4492), .B(n4379), .S(n4737), .Z(n4380) );
  OAI21_X1 U4991 ( .B1(n4440), .B2(n4494), .A(n4380), .ZN(U3533) );
  AOI22_X1 U4992 ( .A1(n4526), .A2(n4414), .B1(n4381), .B2(n4412), .ZN(n4382)
         );
  OAI21_X1 U4993 ( .B1(n4383), .B2(n4397), .A(n4382), .ZN(n4385) );
  AOI211_X1 U4994 ( .C1(n4724), .C2(n4386), .A(n4385), .B(n4384), .ZN(n4495)
         );
  MUX2_X1 U4995 ( .A(n4387), .B(n4495), .S(n4739), .Z(n4388) );
  OAI21_X1 U4996 ( .B1(n4440), .B2(n4498), .A(n4388), .ZN(U3532) );
  AOI21_X1 U4997 ( .B1(n4726), .B2(n4390), .A(n4389), .ZN(n4499) );
  MUX2_X1 U4998 ( .A(n4391), .B(n4499), .S(n4739), .Z(n4392) );
  OAI21_X1 U4999 ( .B1(n4440), .B2(n4502), .A(n4392), .ZN(U3531) );
  NAND2_X1 U5000 ( .A1(n4393), .A2(n4726), .ZN(n4402) );
  AOI22_X1 U5001 ( .A1(n4395), .A2(n4414), .B1(n4412), .B2(n4394), .ZN(n4396)
         );
  OAI21_X1 U5002 ( .B1(n4430), .B2(n4397), .A(n4396), .ZN(n4398) );
  INV_X1 U5003 ( .A(n4398), .ZN(n4399) );
  AND2_X1 U5004 ( .A1(n4400), .A2(n4399), .ZN(n4401) );
  AND2_X1 U5005 ( .A1(n4402), .A2(n4401), .ZN(n4503) );
  MUX2_X1 U5006 ( .A(n2482), .B(n4503), .S(n4739), .Z(n4403) );
  OAI21_X1 U5007 ( .B1(n4505), .B2(n4440), .A(n4403), .ZN(U3530) );
  INV_X1 U5008 ( .A(n4404), .ZN(n4408) );
  INV_X1 U5009 ( .A(n4405), .ZN(n4406) );
  OAI21_X1 U5010 ( .B1(n4408), .B2(n4407), .A(n4406), .ZN(n4642) );
  AOI21_X1 U5011 ( .B1(n4410), .B2(n4409), .A(n2061), .ZN(n4645) );
  INV_X1 U5012 ( .A(n4645), .ZN(n4424) );
  XNOR2_X1 U5013 ( .A(n4411), .B(n4410), .ZN(n4422) );
  AOI22_X1 U5014 ( .A1(n4415), .A2(n4414), .B1(n4413), .B2(n4412), .ZN(n4418)
         );
  NAND2_X1 U5015 ( .A1(n4416), .A2(n4434), .ZN(n4417) );
  OAI211_X1 U5016 ( .C1(n4645), .C2(n4419), .A(n4418), .B(n4417), .ZN(n4420)
         );
  AOI21_X1 U5017 ( .B1(n4422), .B2(n4421), .A(n4420), .ZN(n4652) );
  INV_X1 U5018 ( .A(n4652), .ZN(n4423) );
  AOI21_X1 U5019 ( .B1(n4724), .B2(n4424), .A(n4423), .ZN(n4506) );
  MUX2_X1 U5020 ( .A(n4425), .B(n4506), .S(n4739), .Z(n4426) );
  OAI21_X1 U5021 ( .B1(n4440), .B2(n4642), .A(n4426), .ZN(U3529) );
  OAI22_X1 U5022 ( .A1(n4430), .A2(n4429), .B1(n4428), .B2(n4427), .ZN(n4432)
         );
  AOI211_X1 U5023 ( .C1(n4434), .C2(n4433), .A(n4432), .B(n4431), .ZN(n4435)
         );
  OAI21_X1 U5024 ( .B1(n4437), .B2(n4436), .A(n4435), .ZN(n4438) );
  INV_X1 U5025 ( .A(n4438), .ZN(n4509) );
  MUX2_X1 U5026 ( .A(n2436), .B(n4509), .S(n4739), .Z(n4439) );
  OAI21_X1 U5027 ( .B1(n4512), .B2(n4440), .A(n4439), .ZN(U3528) );
  NOR2_X1 U5028 ( .A1(n4733), .A2(n4441), .ZN(n4442) );
  AOI21_X1 U5029 ( .B1(n4733), .B2(n4443), .A(n4442), .ZN(n4444) );
  OAI21_X1 U5030 ( .B1(n4445), .B2(n4511), .A(n4444), .ZN(U3517) );
  NAND2_X1 U5031 ( .A1(n4545), .A2(n4446), .ZN(n4448) );
  NAND2_X1 U5032 ( .A1(n4544), .A2(n4733), .ZN(n4447) );
  OAI211_X1 U5033 ( .C1(n4733), .C2(n2906), .A(n4448), .B(n4447), .ZN(U3516)
         );
  MUX2_X1 U5034 ( .A(n4450), .B(n4449), .S(n4733), .Z(n4451) );
  OAI21_X1 U5035 ( .B1(n4452), .B2(n4511), .A(n4451), .ZN(U3513) );
  MUX2_X1 U5036 ( .A(n4454), .B(n4453), .S(n4733), .Z(n4455) );
  OAI21_X1 U5037 ( .B1(n4456), .B2(n4511), .A(n4455), .ZN(U3512) );
  MUX2_X1 U5038 ( .A(n4458), .B(n4457), .S(n4733), .Z(n4459) );
  OAI21_X1 U5039 ( .B1(n4460), .B2(n4511), .A(n4459), .ZN(U3511) );
  MUX2_X1 U5040 ( .A(n4462), .B(n4461), .S(n4733), .Z(n4463) );
  OAI21_X1 U5041 ( .B1(n4464), .B2(n4511), .A(n4463), .ZN(U3510) );
  INV_X1 U5042 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4466) );
  MUX2_X1 U5043 ( .A(n4466), .B(n4465), .S(n4733), .Z(n4467) );
  OAI21_X1 U5044 ( .B1(n4468), .B2(n4511), .A(n4467), .ZN(U3509) );
  MUX2_X1 U5045 ( .A(n4470), .B(n4469), .S(n4733), .Z(n4471) );
  OAI21_X1 U5046 ( .B1(n4472), .B2(n4511), .A(n4471), .ZN(U3508) );
  MUX2_X1 U5047 ( .A(n4474), .B(n4473), .S(n4733), .Z(n4475) );
  OAI21_X1 U5048 ( .B1(n4476), .B2(n4511), .A(n4475), .ZN(U3507) );
  MUX2_X1 U5049 ( .A(REG0_REG_20__SCAN_IN), .B(n4477), .S(n4733), .Z(U3506) );
  MUX2_X1 U5050 ( .A(n4479), .B(n4478), .S(n4733), .Z(n4480) );
  OAI21_X1 U5051 ( .B1(n4481), .B2(n4511), .A(n4480), .ZN(U3505) );
  MUX2_X1 U5052 ( .A(REG0_REG_18__SCAN_IN), .B(n4482), .S(n4733), .Z(U3503) );
  MUX2_X1 U5053 ( .A(n4484), .B(n4483), .S(n4732), .Z(n4485) );
  OAI21_X1 U5054 ( .B1(n4486), .B2(n4511), .A(n4485), .ZN(U3501) );
  MUX2_X1 U5055 ( .A(REG0_REG_16__SCAN_IN), .B(n4487), .S(n4733), .Z(n4488) );
  INV_X1 U5056 ( .A(n4488), .ZN(n4489) );
  OAI21_X1 U5057 ( .B1(n4490), .B2(n4511), .A(n4489), .ZN(U3499) );
  MUX2_X1 U5058 ( .A(n4492), .B(n4491), .S(n4732), .Z(n4493) );
  OAI21_X1 U5059 ( .B1(n4494), .B2(n4511), .A(n4493), .ZN(U3497) );
  MUX2_X1 U5060 ( .A(n4496), .B(n4495), .S(n4733), .Z(n4497) );
  OAI21_X1 U5061 ( .B1(n4498), .B2(n4511), .A(n4497), .ZN(U3495) );
  MUX2_X1 U5062 ( .A(n4500), .B(n4499), .S(n4733), .Z(n4501) );
  OAI21_X1 U5063 ( .B1(n4502), .B2(n4511), .A(n4501), .ZN(U3493) );
  MUX2_X1 U5064 ( .A(n4503), .B(n2481), .S(n4732), .Z(n4504) );
  OAI21_X1 U5065 ( .B1(n4505), .B2(n4511), .A(n4504), .ZN(U3491) );
  MUX2_X1 U5066 ( .A(n4507), .B(n4506), .S(n4733), .Z(n4508) );
  OAI21_X1 U5067 ( .B1(n4642), .B2(n4511), .A(n4508), .ZN(U3489) );
  MUX2_X1 U5068 ( .A(n2435), .B(n4509), .S(n4733), .Z(n4510) );
  OAI21_X1 U5069 ( .B1(n4512), .B2(n4511), .A(n4510), .ZN(U3487) );
  MUX2_X1 U5070 ( .A(n2260), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5071 ( .A(n4513), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U5072 ( .A(DATAI_20_), .B(n4514), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5073 ( .A(DATAI_7_), .B(n4515), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U5074 ( .A(n4516), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5075 ( .A(DATAI_4_), .B(n4517), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5076 ( .A(DATAI_2_), .B(n4518), .S(STATE_REG_SCAN_IN), .Z(U3350) );
  MUX2_X1 U5077 ( .A(n4519), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U5078 ( .A(DATAI_28_), .ZN(n4520) );
  AOI22_X1 U5079 ( .A1(STATE_REG_SCAN_IN), .A2(n4521), .B1(n4520), .B2(U3149), 
        .ZN(U3324) );
  NAND2_X1 U5080 ( .A1(n4523), .A2(n4522), .ZN(n4532) );
  NAND2_X1 U5081 ( .A1(n4525), .A2(n4524), .ZN(n4531) );
  NAND2_X1 U5082 ( .A1(n4527), .A2(n4526), .ZN(n4530) );
  NOR2_X1 U5083 ( .A1(STATE_REG_SCAN_IN), .A2(n4528), .ZN(n4614) );
  INV_X1 U5084 ( .A(n4614), .ZN(n4529) );
  AND4_X1 U5085 ( .A1(n4532), .A2(n4531), .A3(n4530), .A4(n4529), .ZN(n4541)
         );
  INV_X1 U5086 ( .A(n4533), .ZN(n4535) );
  OAI21_X1 U5087 ( .B1(n4535), .B2(n4534), .A(n3578), .ZN(n4537) );
  XNOR2_X1 U5088 ( .A(n4537), .B(n4536), .ZN(n4539) );
  NAND2_X1 U5089 ( .A1(n4539), .A2(n4538), .ZN(n4540) );
  OAI211_X1 U5090 ( .C1(n4543), .C2(n4542), .A(n4541), .B(n4540), .ZN(U3223)
         );
  AOI22_X1 U5091 ( .A1(n4545), .A2(n4657), .B1(n4022), .B2(n4544), .ZN(n4546)
         );
  OAI21_X1 U5092 ( .B1(n4547), .B2(n4022), .A(n4546), .ZN(U3261) );
  OAI211_X1 U5093 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4549), .A(n4637), .B(n4548), 
        .ZN(n4553) );
  OAI211_X1 U5094 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4551), .A(n4591), .B(n4550), 
        .ZN(n4552) );
  OAI211_X1 U5095 ( .C1(n4641), .C2(n4712), .A(n4553), .B(n4552), .ZN(n4554)
         );
  AOI211_X1 U5096 ( .C1(n4635), .C2(ADDR_REG_8__SCAN_IN), .A(n4555), .B(n4554), 
        .ZN(n4556) );
  INV_X1 U5097 ( .A(n4556), .ZN(U3248) );
  OAI211_X1 U5098 ( .C1(n4559), .C2(n4558), .A(n4637), .B(n4557), .ZN(n4564)
         );
  OAI211_X1 U5099 ( .C1(n4562), .C2(n4561), .A(n4591), .B(n4560), .ZN(n4563)
         );
  OAI211_X1 U5100 ( .C1(n4641), .C2(n4710), .A(n4564), .B(n4563), .ZN(n4565)
         );
  AOI211_X1 U5101 ( .C1(n4635), .C2(ADDR_REG_9__SCAN_IN), .A(n4566), .B(n4565), 
        .ZN(n4567) );
  INV_X1 U5102 ( .A(n4567), .ZN(U3249) );
  OAI211_X1 U5103 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4570), .A(n4637), .B(n4569), .ZN(n4574) );
  OAI211_X1 U5104 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4572), .A(n4591), .B(n4571), .ZN(n4573) );
  OAI211_X1 U5105 ( .C1(n4641), .C2(n2083), .A(n4574), .B(n4573), .ZN(n4575)
         );
  AOI211_X1 U5106 ( .C1(n4635), .C2(ADDR_REG_10__SCAN_IN), .A(n4576), .B(n4575), .ZN(n4577) );
  INV_X1 U5107 ( .A(n4577), .ZN(U3250) );
  OAI211_X1 U5108 ( .C1(n4580), .C2(n4579), .A(n4637), .B(n4578), .ZN(n4585)
         );
  OAI211_X1 U5109 ( .C1(n4583), .C2(n4582), .A(n4591), .B(n4581), .ZN(n4584)
         );
  OAI211_X1 U5110 ( .C1(n4641), .C2(n4707), .A(n4585), .B(n4584), .ZN(n4586)
         );
  AOI211_X1 U5111 ( .C1(n4635), .C2(ADDR_REG_11__SCAN_IN), .A(n4587), .B(n4586), .ZN(n4588) );
  INV_X1 U5112 ( .A(n4588), .ZN(U3251) );
  OAI211_X1 U5113 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4592), .A(n4591), .B(n4590), .ZN(n4593) );
  NAND2_X1 U5114 ( .A1(n4594), .A2(n4593), .ZN(n4595) );
  AOI21_X1 U5115 ( .B1(n4635), .B2(ADDR_REG_12__SCAN_IN), .A(n4595), .ZN(n4599) );
  OAI211_X1 U5116 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4597), .A(n4637), .B(n4596), .ZN(n4598) );
  OAI211_X1 U5117 ( .C1(n4641), .C2(n2084), .A(n4599), .B(n4598), .ZN(U3252)
         );
  INV_X1 U5118 ( .A(n4600), .ZN(n4605) );
  AOI211_X1 U5119 ( .C1(n4603), .C2(n4602), .A(n4601), .B(n4630), .ZN(n4604)
         );
  AOI211_X1 U5120 ( .C1(ADDR_REG_14__SCAN_IN), .C2(n4635), .A(n4605), .B(n4604), .ZN(n4609) );
  OAI211_X1 U5121 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4607), .A(n4637), .B(n4606), .ZN(n4608) );
  OAI211_X1 U5122 ( .C1(n4641), .C2(n4704), .A(n4609), .B(n4608), .ZN(U3254)
         );
  AOI221_X1 U5123 ( .B1(n4612), .B2(n4611), .C1(n4610), .C2(n4611), .A(n4630), 
        .ZN(n4613) );
  AOI211_X1 U5124 ( .C1(ADDR_REG_16__SCAN_IN), .C2(n4635), .A(n4614), .B(n4613), .ZN(n4618) );
  OAI221_X1 U5125 ( .B1(n4616), .B2(REG1_REG_16__SCAN_IN), .C1(n4616), .C2(
        n4615), .A(n4637), .ZN(n4617) );
  OAI211_X1 U5126 ( .C1(n4641), .C2(n4702), .A(n4618), .B(n4617), .ZN(U3256)
         );
  AOI221_X1 U5127 ( .B1(n4621), .B2(n4620), .C1(n4619), .C2(n4620), .A(n4630), 
        .ZN(n4622) );
  AOI211_X1 U5128 ( .C1(ADDR_REG_17__SCAN_IN), .C2(n4635), .A(n4623), .B(n4622), .ZN(n4628) );
  OAI221_X1 U5129 ( .B1(n4626), .B2(n4625), .C1(n4626), .C2(n4624), .A(n4637), 
        .ZN(n4627) );
  OAI211_X1 U5130 ( .C1(n4641), .C2(n4629), .A(n4628), .B(n4627), .ZN(U3257)
         );
  OAI211_X1 U5131 ( .C1(n4639), .C2(n4638), .A(n4637), .B(n4636), .ZN(n4640)
         );
  OAI22_X1 U5132 ( .A1(n4645), .A2(n4644), .B1(n4643), .B2(n4642), .ZN(n4650)
         );
  OAI22_X1 U5133 ( .A1(n4648), .A2(n4647), .B1(n4646), .B2(n4022), .ZN(n4649)
         );
  NOR2_X1 U5134 ( .A1(n4650), .A2(n4649), .ZN(n4651) );
  OAI21_X1 U5135 ( .B1(n4652), .B2(n4663), .A(n4651), .ZN(U3279) );
  AOI22_X1 U5136 ( .A1(n4654), .A2(n4653), .B1(REG2_REG_8__SCAN_IN), .B2(n4663), .ZN(n4661) );
  INV_X1 U5137 ( .A(n4655), .ZN(n4656) );
  AOI22_X1 U5138 ( .A1(n4659), .A2(n4658), .B1(n4657), .B2(n4656), .ZN(n4660)
         );
  OAI211_X1 U5139 ( .C1(n4663), .C2(n4662), .A(n4661), .B(n4660), .ZN(U3282)
         );
  INV_X1 U5140 ( .A(D_REG_31__SCAN_IN), .ZN(n4664) );
  NOR2_X1 U5141 ( .A1(n4694), .A2(n4664), .ZN(U3291) );
  INV_X1 U5142 ( .A(D_REG_30__SCAN_IN), .ZN(n4665) );
  NOR2_X1 U5143 ( .A1(n4694), .A2(n4665), .ZN(U3292) );
  INV_X1 U5144 ( .A(D_REG_29__SCAN_IN), .ZN(n4666) );
  NOR2_X1 U5145 ( .A1(n4694), .A2(n4666), .ZN(U3293) );
  INV_X1 U5146 ( .A(D_REG_28__SCAN_IN), .ZN(n4667) );
  NOR2_X1 U5147 ( .A1(n4694), .A2(n4667), .ZN(U3294) );
  INV_X1 U5148 ( .A(D_REG_27__SCAN_IN), .ZN(n4668) );
  NOR2_X1 U5149 ( .A1(n4694), .A2(n4668), .ZN(U3295) );
  INV_X1 U5150 ( .A(D_REG_26__SCAN_IN), .ZN(n4669) );
  NOR2_X1 U5151 ( .A1(n4694), .A2(n4669), .ZN(U3296) );
  NOR2_X1 U5152 ( .A1(n4694), .A2(n4670), .ZN(U3297) );
  INV_X1 U5153 ( .A(D_REG_24__SCAN_IN), .ZN(n4671) );
  NOR2_X1 U5154 ( .A1(n4694), .A2(n4671), .ZN(U3298) );
  INV_X1 U5155 ( .A(D_REG_23__SCAN_IN), .ZN(n4672) );
  NOR2_X1 U5156 ( .A1(n4694), .A2(n4672), .ZN(U3299) );
  INV_X1 U5157 ( .A(D_REG_22__SCAN_IN), .ZN(n4673) );
  NOR2_X1 U5158 ( .A1(n4694), .A2(n4673), .ZN(U3300) );
  INV_X1 U5159 ( .A(D_REG_21__SCAN_IN), .ZN(n4674) );
  NOR2_X1 U5160 ( .A1(n4694), .A2(n4674), .ZN(U3301) );
  INV_X1 U5161 ( .A(D_REG_20__SCAN_IN), .ZN(n4675) );
  NOR2_X1 U5162 ( .A1(n4694), .A2(n4675), .ZN(U3302) );
  INV_X1 U5163 ( .A(D_REG_19__SCAN_IN), .ZN(n4676) );
  NOR2_X1 U5164 ( .A1(n4694), .A2(n4676), .ZN(U3303) );
  INV_X1 U5165 ( .A(D_REG_18__SCAN_IN), .ZN(n4677) );
  NOR2_X1 U5166 ( .A1(n4694), .A2(n4677), .ZN(U3304) );
  INV_X1 U5167 ( .A(D_REG_17__SCAN_IN), .ZN(n4678) );
  NOR2_X1 U5168 ( .A1(n4694), .A2(n4678), .ZN(U3305) );
  INV_X1 U5169 ( .A(D_REG_16__SCAN_IN), .ZN(n4679) );
  NOR2_X1 U5170 ( .A1(n4694), .A2(n4679), .ZN(U3306) );
  NOR2_X1 U5171 ( .A1(n4694), .A2(n4680), .ZN(U3307) );
  INV_X1 U5172 ( .A(D_REG_14__SCAN_IN), .ZN(n4681) );
  NOR2_X1 U5173 ( .A1(n4694), .A2(n4681), .ZN(U3308) );
  INV_X1 U5174 ( .A(D_REG_13__SCAN_IN), .ZN(n4682) );
  NOR2_X1 U5175 ( .A1(n4694), .A2(n4682), .ZN(U3309) );
  INV_X1 U5176 ( .A(D_REG_12__SCAN_IN), .ZN(n4683) );
  NOR2_X1 U5177 ( .A1(n4694), .A2(n4683), .ZN(U3310) );
  NOR2_X1 U5178 ( .A1(n4694), .A2(n4684), .ZN(U3311) );
  INV_X1 U5179 ( .A(D_REG_10__SCAN_IN), .ZN(n4685) );
  NOR2_X1 U5180 ( .A1(n4694), .A2(n4685), .ZN(U3312) );
  INV_X1 U5181 ( .A(D_REG_9__SCAN_IN), .ZN(n4686) );
  NOR2_X1 U5182 ( .A1(n4694), .A2(n4686), .ZN(U3313) );
  INV_X1 U5183 ( .A(D_REG_8__SCAN_IN), .ZN(n4687) );
  NOR2_X1 U5184 ( .A1(n4694), .A2(n4687), .ZN(U3314) );
  INV_X1 U5185 ( .A(D_REG_7__SCAN_IN), .ZN(n4688) );
  NOR2_X1 U5186 ( .A1(n4694), .A2(n4688), .ZN(U3315) );
  INV_X1 U5187 ( .A(D_REG_6__SCAN_IN), .ZN(n4689) );
  NOR2_X1 U5188 ( .A1(n4694), .A2(n4689), .ZN(U3316) );
  INV_X1 U5189 ( .A(D_REG_5__SCAN_IN), .ZN(n4690) );
  NOR2_X1 U5190 ( .A1(n4694), .A2(n4690), .ZN(U3317) );
  INV_X1 U5191 ( .A(D_REG_4__SCAN_IN), .ZN(n4691) );
  NOR2_X1 U5192 ( .A1(n4694), .A2(n4691), .ZN(U3318) );
  NOR2_X1 U5193 ( .A1(n4694), .A2(n4692), .ZN(U3319) );
  INV_X1 U5194 ( .A(D_REG_2__SCAN_IN), .ZN(n4693) );
  NOR2_X1 U5195 ( .A1(n4694), .A2(n4693), .ZN(U3320) );
  AOI21_X1 U5196 ( .B1(U3149), .B2(n4696), .A(n4695), .ZN(U3329) );
  AOI22_X1 U5197 ( .A1(STATE_REG_SCAN_IN), .A2(n4698), .B1(n4697), .B2(U3149), 
        .ZN(U3334) );
  OAI22_X1 U5198 ( .A1(U3149), .A2(n4699), .B1(DATAI_17_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4700) );
  INV_X1 U5199 ( .A(n4700), .ZN(U3335) );
  INV_X1 U5200 ( .A(DATAI_16_), .ZN(n4701) );
  AOI22_X1 U5201 ( .A1(STATE_REG_SCAN_IN), .A2(n4702), .B1(n4701), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5202 ( .A(DATAI_14_), .ZN(n4703) );
  AOI22_X1 U5203 ( .A1(STATE_REG_SCAN_IN), .A2(n4704), .B1(n4703), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5204 ( .A(DATAI_12_), .ZN(n4705) );
  AOI22_X1 U5205 ( .A1(STATE_REG_SCAN_IN), .A2(n2084), .B1(n4705), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5206 ( .A(DATAI_11_), .ZN(n4706) );
  AOI22_X1 U5207 ( .A1(STATE_REG_SCAN_IN), .A2(n4707), .B1(n4706), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5208 ( .A(DATAI_10_), .ZN(n4708) );
  AOI22_X1 U5209 ( .A1(STATE_REG_SCAN_IN), .A2(n2083), .B1(n4708), .B2(U3149), 
        .ZN(U3342) );
  AOI22_X1 U5210 ( .A1(STATE_REG_SCAN_IN), .A2(n4710), .B1(n4709), .B2(U3149), 
        .ZN(U3343) );
  AOI22_X1 U5211 ( .A1(STATE_REG_SCAN_IN), .A2(n4712), .B1(n4711), .B2(U3149), 
        .ZN(U3344) );
  INV_X1 U5212 ( .A(DATAI_0_), .ZN(n4713) );
  AOI22_X1 U5213 ( .A1(STATE_REG_SCAN_IN), .A2(n2291), .B1(n4713), .B2(U3149), 
        .ZN(U3352) );
  AOI22_X1 U5214 ( .A1(n4733), .A2(n4714), .B1(n2263), .B2(n4732), .ZN(U3467)
         );
  INV_X1 U5215 ( .A(n4715), .ZN(n4717) );
  AOI211_X1 U5216 ( .C1(n4718), .C2(n4724), .A(n4717), .B(n4716), .ZN(n4735)
         );
  AOI22_X1 U5217 ( .A1(n4733), .A2(n4735), .B1(n2339), .B2(n4732), .ZN(U3475)
         );
  NOR3_X1 U5218 ( .A1(n4721), .A2(n4720), .A3(n4719), .ZN(n4723) );
  AOI211_X1 U5219 ( .C1(n4725), .C2(n4724), .A(n4723), .B(n4722), .ZN(n4736)
         );
  AOI22_X1 U5220 ( .A1(n4733), .A2(n4736), .B1(n2374), .B2(n4732), .ZN(U3479)
         );
  NAND3_X1 U5221 ( .A1(n4728), .A2(n4727), .A3(n4726), .ZN(n4729) );
  AND3_X1 U5222 ( .A1(n4731), .A2(n4730), .A3(n4729), .ZN(n4738) );
  AOI22_X1 U5223 ( .A1(n4733), .A2(n4738), .B1(n2394), .B2(n4732), .ZN(U3481)
         );
  INV_X1 U5224 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4734) );
  AOI22_X1 U5225 ( .A1(n4739), .A2(n4735), .B1(n4734), .B2(n4737), .ZN(U3522)
         );
  AOI22_X1 U5226 ( .A1(n4739), .A2(n4736), .B1(n2375), .B2(n4737), .ZN(U3524)
         );
  AOI22_X1 U5227 ( .A1(n4739), .A2(n4738), .B1(n3210), .B2(n4737), .ZN(U3525)
         );
  CLKBUF_X3 U2272 ( .A(n2318), .Z(n2678) );
  INV_X1 U2281 ( .A(n3177), .ZN(n3282) );
  AND2_X2 U2710 ( .A1(n2262), .A2(n2939), .ZN(n4742) );
endmodule

