

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, 
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, 
        keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, 
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, 
        keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, 
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, 
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2133, n2134, n2135, n2136, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081;

  INV_X1 U2375 ( .A(n3405), .ZN(n3553) );
  NAND2_X1 U2376 ( .A1(n2819), .A2(n2723), .ZN(n4190) );
  NAND2_X1 U2377 ( .A1(n2575), .A2(n2464), .ZN(n4207) );
  NAND2_X1 U2378 ( .A1(n2861), .A2(n4948), .ZN(n2947) );
  INV_X1 U2379 ( .A(n2534), .ZN(n2748) );
  OAI21_X2 U2380 ( .B1(n4056), .B2(n2560), .A(n2559), .ZN(n2583) );
  CLKBUF_X2 U2381 ( .A(n4208), .Z(n2135) );
  INV_X1 U2382 ( .A(n3012), .ZN(n2979) );
  XNOR2_X1 U2383 ( .A(n3235), .B(n3513), .ZN(n3510) );
  NAND2_X1 U2384 ( .A1(n4116), .A2(n4119), .ZN(n4099) );
  OAI21_X1 U2385 ( .B1(n4056), .B2(n2178), .A(n2177), .ZN(n3577) );
  OR2_X1 U2386 ( .A1(n2686), .A2(n4761), .ZN(n2695) );
  INV_X2 U2387 ( .A(n3035), .ZN(n3088) );
  AND2_X1 U2388 ( .A1(n2272), .A2(n2266), .ZN(n4983) );
  AND2_X1 U2389 ( .A1(n4397), .A2(n4382), .ZN(n4377) );
  INV_X1 U2390 ( .A(n3812), .ZN(n4200) );
  NAND2_X2 U2391 ( .A1(n4512), .A2(n2760), .ZN(n4315) );
  NAND2_X2 U2392 ( .A1(n4341), .A2(n4340), .ZN(n4512) );
  NOR2_X2 U2393 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2227)
         );
  NAND2_X1 U2394 ( .A1(n2415), .A2(n2496), .ZN(n2133) );
  INV_X1 U2395 ( .A(n2133), .ZN(n2134) );
  NOR2_X2 U2396 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2718)
         );
  NAND4_X1 U2397 ( .A1(n2541), .A2(n2540), .A3(n2539), .A4(n2538), .ZN(n4208)
         );
  NAND3_X2 U2398 ( .A1(n2292), .A2(n4608), .A3(n2291), .ZN(n4210) );
  NAND2_X2 U2399 ( .A1(n2532), .A2(n2294), .ZN(n4608) );
  XNOR2_X2 U2400 ( .A(n3244), .B(n3800), .ZN(n3797) );
  NAND2_X2 U2401 ( .A1(n4226), .A2(n3243), .ZN(n3244) );
  NAND2_X2 U2402 ( .A1(n2579), .A2(n2348), .ZN(n3345) );
  NOR2_X2 U2403 ( .A1(n3209), .A2(n5010), .ZN(n5020) );
  OAI21_X2 U2404 ( .B1(n4995), .B2(n2343), .A(n2342), .ZN(n5010) );
  OAI211_X1 U2405 ( .C1(n3837), .C2(n5069), .A(n2864), .B(n3846), .ZN(n3265)
         );
  INV_X1 U2406 ( .A(n4483), .ZN(n4497) );
  OAI21_X1 U2407 ( .B1(n2323), .B2(REG1_REG_7__SCAN_IN), .A(n2178), .ZN(n3193)
         );
  NOR2_X1 U2408 ( .A1(n3446), .A2(n3449), .ZN(n2581) );
  NAND2_X1 U2409 ( .A1(n3302), .A2(n3229), .ZN(n3231) );
  NAND2_X2 U2410 ( .A1(n4136), .A2(n2845), .ZN(n4131) );
  INV_X2 U2411 ( .A(n2979), .ZN(n3029) );
  AND2_X1 U2412 ( .A1(n4551), .A2(n3112), .ZN(n2972) );
  INV_X4 U2413 ( .A(n3112), .ZN(n2955) );
  INV_X2 U2414 ( .A(n3531), .ZN(n2567) );
  INV_X2 U2415 ( .A(n2941), .ZN(n4551) );
  CLKBUF_X2 U2416 ( .A(n2550), .Z(n3330) );
  INV_X1 U2417 ( .A(IR_REG_20__SCAN_IN), .ZN(n2820) );
  CLKBUF_X1 U2418 ( .A(IR_REG_0__SCAN_IN), .Z(n5060) );
  AND2_X1 U2419 ( .A1(n3845), .A2(n2308), .ZN(n2307) );
  OAI21_X1 U2420 ( .B1(n3265), .B2(n5075), .A(n3267), .ZN(n3268) );
  NAND2_X1 U2421 ( .A1(n2191), .A2(n2193), .ZN(n4276) );
  AND2_X1 U2422 ( .A1(n2858), .A2(n2385), .ZN(n2384) );
  AND2_X1 U2423 ( .A1(n2818), .A2(n2817), .ZN(n4486) );
  NAND2_X1 U2424 ( .A1(n2799), .A2(n2798), .ZN(n4483) );
  NAND2_X1 U2425 ( .A1(n2779), .A2(n2778), .ZN(n4494) );
  AND2_X1 U2426 ( .A1(n4377), .A2(n2143), .ZN(n4301) );
  NAND2_X1 U2427 ( .A1(n2447), .A2(n2446), .ZN(n3793) );
  INV_X1 U2428 ( .A(n4417), .ZN(n4527) );
  AND2_X1 U2429 ( .A1(n2716), .A2(n2715), .ZN(n4417) );
  OR2_X1 U2430 ( .A1(n3477), .A2(n3478), .ZN(n2366) );
  AOI21_X1 U2431 ( .B1(n3232), .B2(n3563), .A(n2285), .ZN(n2282) );
  OR2_X1 U2432 ( .A1(n3406), .A2(n2301), .ZN(n3575) );
  NAND2_X1 U2433 ( .A1(n3231), .A2(n3230), .ZN(n3232) );
  XNOR2_X1 U2434 ( .A(n3231), .B(n3392), .ZN(n3390) );
  OAI21_X2 U2435 ( .B1(n3155), .B2(n3154), .A(n4451), .ZN(n3156) );
  AND2_X1 U2436 ( .A1(n4131), .A2(n2467), .ZN(n2605) );
  CLKBUF_X3 U2437 ( .A(n2972), .Z(n3116) );
  BUF_X1 U2438 ( .A(U4043), .Z(n4202) );
  NAND2_X1 U2439 ( .A1(n2225), .A2(n2175), .ZN(n3832) );
  AND2_X1 U2440 ( .A1(n3188), .A2(n2560), .ZN(n2465) );
  OR2_X1 U2441 ( .A1(n4465), .A2(n3318), .ZN(n4119) );
  NAND4_X2 U2442 ( .A1(n2555), .A2(n2554), .A3(n2553), .A4(n2552), .ZN(n4470)
         );
  NOR2_X4 U2443 ( .A1(n4949), .A2(n3310), .ZN(n2941) );
  XNOR2_X1 U2444 ( .A(n3222), .B(n3184), .ZN(n3292) );
  NAND4_X2 U2445 ( .A1(n2522), .A2(n2523), .A3(n2521), .A4(n2520), .ZN(n4465)
         );
  INV_X1 U2446 ( .A(n2861), .ZN(n4949) );
  OR2_X1 U2447 ( .A1(n2946), .A2(n4948), .ZN(n3310) );
  OR2_X1 U2448 ( .A1(n2923), .A2(n2493), .ZN(n2495) );
  NAND2_X1 U2449 ( .A1(n2819), .A2(IR_REG_31__SCAN_IN), .ZN(n2821) );
  NAND2_X1 U2450 ( .A1(n3346), .A2(n3182), .ZN(n3183) );
  XNOR2_X1 U2451 ( .A(n2827), .B(IR_REG_22__SCAN_IN), .ZN(n2946) );
  INV_X1 U2452 ( .A(n3419), .ZN(n2285) );
  NAND2_X1 U2454 ( .A1(n3348), .A2(n3347), .ZN(n3346) );
  AND2_X1 U2455 ( .A1(n2556), .A2(n2549), .ZN(n4957) );
  NAND2_X1 U2456 ( .A1(n2881), .A2(IR_REG_31__SCAN_IN), .ZN(n2827) );
  NAND2_X1 U2457 ( .A1(n3220), .A2(n3219), .ZN(n3351) );
  XNOR2_X1 U2458 ( .A(n2824), .B(IR_REG_21__SCAN_IN), .ZN(n4948) );
  OR2_X1 U2459 ( .A1(n2826), .A2(n2293), .ZN(n2824) );
  NAND2_X1 U2460 ( .A1(n2826), .A2(n2825), .ZN(n2881) );
  INV_X1 U2461 ( .A(n2596), .ZN(n2136) );
  INV_X1 U2462 ( .A(IR_REG_22__SCAN_IN), .ZN(n2486) );
  NOR2_X1 U2463 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2488)
         );
  INV_X1 U2464 ( .A(IR_REG_21__SCAN_IN), .ZN(n2825) );
  NOR2_X1 U2465 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2489)
         );
  NOR2_X1 U2466 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_2__SCAN_IN), .ZN(n2478)
         );
  NOR2_X1 U2467 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2354)
         );
  INV_X1 U2468 ( .A(IR_REG_3__SCAN_IN), .ZN(n2576) );
  INV_X1 U2469 ( .A(IR_REG_27__SCAN_IN), .ZN(n2506) );
  NOR2_X1 U2470 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2228)
         );
  NOR2_X2 U2471 ( .A1(n3300), .A2(n3189), .ZN(n3190) );
  OAI21_X2 U2472 ( .B1(n4234), .B2(n4760), .A(n2332), .ZN(n4987) );
  BUF_X4 U2473 ( .A(n2536), .Z(n2812) );
  NAND2_X2 U2474 ( .A1(n3282), .A2(n3280), .ZN(n2536) );
  AND2_X1 U2475 ( .A1(n2247), .A2(n2166), .ZN(n2246) );
  NAND2_X1 U2476 ( .A1(n2249), .A2(n2161), .ZN(n2247) );
  AOI21_X1 U2477 ( .B1(n2391), .B2(n2389), .A(n2388), .ZN(n2387) );
  INV_X1 U2478 ( .A(n4172), .ZN(n2388) );
  XNOR2_X1 U2479 ( .A(n2484), .B(IR_REG_17__SCAN_IN), .ZN(n3254) );
  INV_X1 U2480 ( .A(n3039), .ZN(n3040) );
  INV_X1 U2481 ( .A(n2742), .ZN(n2458) );
  NAND2_X1 U2482 ( .A1(n2249), .A2(n3054), .ZN(n2245) );
  INV_X1 U2483 ( .A(n2242), .ZN(n2241) );
  OAI21_X1 U2484 ( .B1(n2246), .B2(n2244), .A(n2243), .ZN(n2242) );
  NAND2_X1 U2485 ( .A1(n3418), .A2(n3234), .ZN(n3235) );
  INV_X1 U2486 ( .A(n3599), .ZN(n2288) );
  AOI21_X1 U2487 ( .B1(n2933), .B2(n2441), .A(n2932), .ZN(n2440) );
  NAND2_X1 U2488 ( .A1(n2444), .A2(n2806), .ZN(n2441) );
  NAND2_X1 U2489 ( .A1(n2192), .A2(n4173), .ZN(n2191) );
  OR2_X1 U2490 ( .A1(n2910), .A2(n2896), .ZN(n2909) );
  INV_X1 U2491 ( .A(IR_REG_8__SCAN_IN), .ZN(n2477) );
  NOR2_X1 U2492 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2229)
         );
  INV_X1 U2493 ( .A(IR_REG_23__SCAN_IN), .ZN(n2883) );
  INV_X1 U2494 ( .A(n3865), .ZN(n2262) );
  OAI21_X1 U2495 ( .B1(n3990), .B2(n3991), .A(n3992), .ZN(n3025) );
  NAND2_X1 U2496 ( .A1(n3990), .A2(n3991), .ZN(n3024) );
  NAND2_X1 U2497 ( .A1(n2197), .A2(n4160), .ZN(n3735) );
  NAND2_X1 U2498 ( .A1(n3769), .A2(n4156), .ZN(n2197) );
  AOI21_X1 U2499 ( .B1(n2431), .B2(n2429), .A(n2163), .ZN(n2428) );
  INV_X1 U2500 ( .A(n2537), .ZN(n2813) );
  AND2_X1 U2501 ( .A1(n4091), .A2(n2533), .ZN(n2426) );
  NAND2_X1 U2502 ( .A1(n2943), .A2(n5049), .ZN(n3211) );
  AND2_X1 U2503 ( .A1(n2900), .A2(n2899), .ZN(n3132) );
  OR2_X1 U2504 ( .A1(n2910), .A2(D_REG_0__SCAN_IN), .ZN(n2900) );
  NAND2_X1 U2505 ( .A1(n3862), .A2(IR_REG_31__SCAN_IN), .ZN(n2509) );
  NAND2_X1 U2506 ( .A1(n2543), .A2(n2542), .ZN(n2579) );
  NAND2_X1 U2507 ( .A1(n2344), .A2(n4794), .ZN(n2343) );
  NAND2_X1 U2508 ( .A1(n3208), .A2(n2344), .ZN(n2342) );
  INV_X1 U2509 ( .A(n5011), .ZN(n2344) );
  NAND2_X1 U2510 ( .A1(n3992), .A2(n3991), .ZN(n2250) );
  AND2_X1 U2511 ( .A1(n3040), .A2(n2383), .ZN(n2379) );
  INV_X1 U2512 ( .A(n2496), .ZN(n2414) );
  NOR2_X1 U2513 ( .A1(n2762), .A2(n2761), .ZN(n2187) );
  OR2_X1 U2514 ( .A1(n3068), .A2(n3067), .ZN(n3069) );
  INV_X1 U2515 ( .A(n4193), .ZN(n3150) );
  OAI21_X1 U2516 ( .B1(n3236), .B2(n2288), .A(n3238), .ZN(n2287) );
  NAND2_X1 U2517 ( .A1(n2404), .A2(n2403), .ZN(n2402) );
  NAND2_X1 U2518 ( .A1(n2387), .A2(n2390), .ZN(n2385) );
  INV_X1 U2519 ( .A(n2391), .ZN(n2390) );
  AOI21_X1 U2520 ( .B1(n4049), .B2(n4165), .A(n2392), .ZN(n2391) );
  INV_X1 U2521 ( .A(n4169), .ZN(n2392) );
  AND2_X1 U2522 ( .A1(n2459), .A2(n2455), .ZN(n2454) );
  NAND2_X1 U2523 ( .A1(n2458), .A2(n2456), .ZN(n2455) );
  INV_X1 U2524 ( .A(n2460), .ZN(n2456) );
  NAND2_X1 U2525 ( .A1(n2458), .A2(n2707), .ZN(n2457) );
  NAND2_X1 U2526 ( .A1(n4555), .A2(n4541), .ZN(n2460) );
  NAND2_X1 U2527 ( .A1(n4443), .A2(n4162), .ZN(n4368) );
  INV_X1 U2528 ( .A(n4149), .ZN(n2213) );
  INV_X1 U2529 ( .A(n2468), .ZN(n2430) );
  NAND2_X1 U2530 ( .A1(n3546), .A2(n2618), .ZN(n2418) );
  NOR2_X1 U2531 ( .A1(n4207), .A2(n3534), .ZN(n3449) );
  NOR2_X1 U2532 ( .A1(n2206), .A2(n2203), .ZN(n2201) );
  NAND2_X1 U2533 ( .A1(n3488), .A2(n2585), .ZN(n3447) );
  NAND2_X1 U2534 ( .A1(n2840), .A2(n2426), .ZN(n2425) );
  AND2_X1 U2535 ( .A1(n2547), .A2(n2423), .ZN(n2422) );
  NOR2_X1 U2536 ( .A1(n2318), .A2(n4317), .ZN(n2317) );
  INV_X1 U2537 ( .A(n2319), .ZN(n2318) );
  AND2_X1 U2538 ( .A1(n3644), .A2(n3689), .ZN(n2316) );
  AND2_X1 U2539 ( .A1(n2946), .A2(n4948), .ZN(n3213) );
  NOR2_X1 U2540 ( .A1(IR_REG_25__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .ZN(n2421)
         );
  OR3_X1 U2541 ( .A1(n2691), .A2(IR_REG_15__SCAN_IN), .A3(n2483), .ZN(n2733)
         );
  NAND4_X1 U2542 ( .A1(n2478), .A2(n2532), .A3(n2576), .A4(n2354), .ZN(n2596)
         );
  INV_X1 U2543 ( .A(n2237), .ZN(n2236) );
  NOR2_X1 U2544 ( .A1(n2236), .A2(n2232), .ZN(n2231) );
  INV_X1 U2545 ( .A(n2357), .ZN(n2232) );
  NAND2_X1 U2546 ( .A1(n2238), .A2(n2151), .ZN(n2237) );
  INV_X1 U2547 ( .A(n3698), .ZN(n2238) );
  NAND2_X1 U2548 ( .A1(n2188), .A2(REG3_REG_21__SCAN_IN), .ZN(n2753) );
  INV_X1 U2549 ( .A(n3069), .ZN(n2376) );
  NOR2_X1 U2550 ( .A1(n2373), .A2(n2377), .ZN(n2372) );
  INV_X1 U2551 ( .A(n3964), .ZN(n2377) );
  INV_X1 U2552 ( .A(n3893), .ZN(n2373) );
  NAND2_X1 U2553 ( .A1(n2783), .A2(REG3_REG_25__SCAN_IN), .ZN(n2793) );
  INV_X1 U2554 ( .A(n2785), .ZN(n2783) );
  NAND2_X1 U2555 ( .A1(n2986), .A2(n2987), .ZN(n2368) );
  INV_X1 U2556 ( .A(n2369), .ZN(n2365) );
  INV_X1 U2557 ( .A(n3529), .ZN(n2367) );
  NAND2_X1 U2558 ( .A1(n2502), .A2(REG3_REG_16__SCAN_IN), .ZN(n2697) );
  INV_X1 U2559 ( .A(n2695), .ZN(n2502) );
  NAND2_X1 U2560 ( .A1(n2187), .A2(REG3_REG_24__SCAN_IN), .ZN(n2785) );
  INV_X1 U2561 ( .A(n2187), .ZN(n2772) );
  AND2_X1 U2562 ( .A1(n2359), .A2(n3632), .ZN(n2356) );
  NAND2_X1 U2563 ( .A1(n2360), .A2(n3633), .ZN(n2359) );
  INV_X1 U2564 ( .A(n2361), .ZN(n2360) );
  INV_X1 U2565 ( .A(n2188), .ZN(n2744) );
  INV_X1 U2566 ( .A(n3919), .ZN(n2383) );
  OR2_X1 U2567 ( .A1(n3910), .A2(n3085), .ZN(n2258) );
  OR2_X1 U2568 ( .A1(n3021), .A2(n3020), .ZN(n3022) );
  NAND2_X1 U2569 ( .A1(n2148), .A2(n3085), .ZN(n2256) );
  INV_X1 U2570 ( .A(n3155), .ZN(n3144) );
  NAND2_X1 U2572 ( .A1(n2546), .A2(REG1_REG_2__SCAN_IN), .ZN(n3182) );
  INV_X1 U2573 ( .A(n4957), .ZN(n3184) );
  INV_X1 U2574 ( .A(n4959), .ZN(n3341) );
  AND2_X1 U2575 ( .A1(n4956), .A2(REG1_REG_5__SCAN_IN), .ZN(n3189) );
  NAND2_X1 U2576 ( .A1(n3510), .A2(REG2_REG_8__SCAN_IN), .ZN(n3237) );
  INV_X1 U2577 ( .A(n2321), .ZN(n2320) );
  OAI21_X1 U2578 ( .B1(n3200), .B2(n2322), .A(n3202), .ZN(n2321) );
  NOR2_X1 U2579 ( .A1(n4240), .A2(n2271), .ZN(n2269) );
  OR2_X1 U2580 ( .A1(n4972), .A2(n2264), .ZN(n2267) );
  NAND2_X1 U2581 ( .A1(n4240), .A2(n2265), .ZN(n2264) );
  INV_X1 U2582 ( .A(n4970), .ZN(n2265) );
  AND2_X1 U2583 ( .A1(n3250), .A2(REG2_REG_15__SCAN_IN), .ZN(n2290) );
  INV_X1 U2584 ( .A(n3210), .ZN(n2341) );
  INV_X1 U2585 ( .A(n2440), .ZN(n2439) );
  INV_X1 U2586 ( .A(n2812), .ZN(n2830) );
  NOR2_X1 U2587 ( .A1(n4348), .A2(n4310), .ZN(n4328) );
  NAND2_X1 U2588 ( .A1(n2503), .A2(REG3_REG_17__SCAN_IN), .ZN(n2725) );
  INV_X1 U2589 ( .A(n2697), .ZN(n2503) );
  NAND2_X1 U2590 ( .A1(n4564), .A2(n4455), .ZN(n2706) );
  OR2_X1 U2591 ( .A1(n4574), .A2(n4560), .ZN(n2693) );
  NAND2_X1 U2592 ( .A1(n3735), .A2(n3736), .ZN(n2851) );
  NAND2_X1 U2593 ( .A1(n2851), .A2(n2393), .ZN(n3784) );
  NOR2_X1 U2594 ( .A1(n4080), .A2(n2394), .ZN(n2393) );
  INV_X1 U2595 ( .A(n4043), .ZN(n2394) );
  NAND2_X1 U2596 ( .A1(n2849), .A2(n4154), .ZN(n3769) );
  OR2_X1 U2597 ( .A1(n3703), .A2(n3708), .ZN(n2176) );
  AOI21_X1 U2598 ( .B1(n2408), .B2(n2407), .A(n2406), .ZN(n2405) );
  INV_X1 U2599 ( .A(n4136), .ZN(n2407) );
  INV_X1 U2600 ( .A(n4135), .ZN(n2406) );
  NAND2_X2 U2601 ( .A1(n4206), .A2(n3577), .ZN(n4136) );
  AOI21_X1 U2602 ( .B1(n2207), .B2(n2843), .A(n2205), .ZN(n2204) );
  INV_X1 U2603 ( .A(n4143), .ZN(n2205) );
  NAND2_X1 U2604 ( .A1(n3401), .A2(n4125), .ZN(n3433) );
  INV_X1 U2605 ( .A(n3433), .ZN(n2211) );
  NAND2_X1 U2606 ( .A1(n2720), .A2(IR_REG_31__SCAN_IN), .ZN(n2722) );
  INV_X1 U2607 ( .A(IR_REG_19__SCAN_IN), .ZN(n2721) );
  NAND2_X1 U2608 ( .A1(n3402), .A2(n4094), .ZN(n3401) );
  NAND2_X1 U2609 ( .A1(n2226), .A2(n3832), .ZN(n3314) );
  INV_X1 U2610 ( .A(n2963), .ZN(n2226) );
  AND2_X1 U2611 ( .A1(n2909), .A2(n3290), .ZN(n3133) );
  INV_X1 U2612 ( .A(n3832), .ZN(n3311) );
  INV_X1 U2613 ( .A(n2437), .ZN(n2436) );
  INV_X1 U2614 ( .A(n3125), .ZN(n4482) );
  OR2_X1 U2615 ( .A1(n3815), .A2(n4019), .ZN(n4263) );
  NAND2_X1 U2616 ( .A1(n4301), .A2(n4285), .ZN(n3815) );
  INV_X1 U2617 ( .A(n4378), .ZN(n4530) );
  AND2_X1 U2618 ( .A1(n3786), .A2(n2169), .ZN(n4397) );
  AND3_X1 U2619 ( .A1(n2684), .A2(n2683), .A3(n2682), .ZN(n4562) );
  OR2_X1 U2620 ( .A1(n3778), .A2(n4571), .ZN(n3787) );
  INV_X1 U2621 ( .A(n4589), .ZN(n4573) );
  OR2_X1 U2622 ( .A1(n5026), .A2(n2946), .ZN(n3740) );
  INV_X1 U2623 ( .A(n3211), .ZN(n3827) );
  NAND2_X1 U2624 ( .A1(n2877), .A2(n4947), .ZN(n2910) );
  INV_X1 U2625 ( .A(IR_REG_29__SCAN_IN), .ZN(n2507) );
  INV_X1 U2626 ( .A(IR_REG_24__SCAN_IN), .ZN(n2485) );
  XNOR2_X1 U2627 ( .A(n2884), .B(n2883), .ZN(n3212) );
  NAND2_X1 U2628 ( .A1(n2882), .A2(IR_REG_31__SCAN_IN), .ZN(n2884) );
  NAND2_X1 U2629 ( .A1(n2692), .A2(IR_REG_31__SCAN_IN), .ZN(n2702) );
  OR2_X1 U2630 ( .A1(n2691), .A2(IR_REG_14__SCAN_IN), .ZN(n2692) );
  OR2_X1 U2631 ( .A1(n2643), .A2(IR_REG_10__SCAN_IN), .ZN(n2652) );
  INV_X1 U2632 ( .A(IR_REG_4__SCAN_IN), .ZN(n2577) );
  INV_X1 U2633 ( .A(IR_REG_1__SCAN_IN), .ZN(n2294) );
  NOR2_X1 U2634 ( .A1(n2141), .A2(n2261), .ZN(n2259) );
  INV_X1 U2635 ( .A(n3156), .ZN(n3985) );
  INV_X1 U2636 ( .A(n4033), .ZN(n3934) );
  OR2_X1 U2637 ( .A1(n3152), .A2(n3341), .ZN(n4033) );
  OAI21_X1 U2638 ( .B1(n3366), .B2(n2346), .A(n2345), .ZN(n3300) );
  NAND2_X1 U2639 ( .A1(n2347), .A2(REG1_REG_4__SCAN_IN), .ZN(n2346) );
  NAND2_X1 U2640 ( .A1(n2465), .A2(n2347), .ZN(n2345) );
  INV_X1 U2641 ( .A(n3301), .ZN(n2347) );
  NAND2_X1 U2642 ( .A1(n5018), .A2(ADDR_REG_17__SCAN_IN), .ZN(n2182) );
  NAND2_X1 U2643 ( .A1(n5007), .A2(n2184), .ZN(n2183) );
  OR2_X1 U2644 ( .A1(n5006), .A2(n5008), .ZN(n2184) );
  NAND2_X1 U2645 ( .A1(n2298), .A2(n5001), .ZN(n2297) );
  NAND2_X1 U2646 ( .A1(n5007), .A2(n2300), .ZN(n2299) );
  AND2_X1 U2647 ( .A1(n5007), .A2(n2279), .ZN(n5015) );
  AOI21_X1 U2648 ( .B1(n5018), .B2(ADDR_REG_18__SCAN_IN), .A(n5017), .ZN(n2296) );
  NAND2_X1 U2649 ( .A1(n5020), .A2(n5021), .ZN(n5019) );
  NAND2_X1 U2650 ( .A1(n5019), .A2(n2335), .ZN(n2333) );
  NOR2_X1 U2651 ( .A1(n2340), .A2(n2337), .ZN(n2335) );
  NOR2_X1 U2652 ( .A1(n2338), .A2(n3210), .ZN(n2337) );
  INV_X1 U2653 ( .A(n2466), .ZN(n2338) );
  AND2_X1 U2654 ( .A1(n2276), .A2(n2277), .ZN(n3257) );
  AOI21_X1 U2655 ( .B1(n2279), .B2(n2278), .A(n2281), .ZN(n2277) );
  INV_X1 U2656 ( .A(n3846), .ZN(n2312) );
  NAND2_X1 U2657 ( .A1(n2311), .A2(n2310), .ZN(n2309) );
  INV_X1 U2658 ( .A(n3844), .ZN(n2311) );
  NAND2_X1 U2659 ( .A1(n4200), .A2(n4466), .ZN(n2310) );
  NAND2_X1 U2660 ( .A1(n2196), .A2(n2397), .ZN(n4259) );
  OR2_X1 U2661 ( .A1(n2536), .A2(n2518), .ZN(n2523) );
  OR2_X1 U2662 ( .A1(n2537), .A2(n3216), .ZN(n2522) );
  NAND2_X1 U2663 ( .A1(n5032), .A2(n2915), .ZN(n4458) );
  NAND2_X1 U2664 ( .A1(n2906), .A2(n2313), .ZN(n3843) );
  OR2_X1 U2665 ( .A1(n4264), .A2(n3128), .ZN(n2313) );
  INV_X1 U2666 ( .A(n3255), .ZN(n5052) );
  INV_X1 U2667 ( .A(n3991), .ZN(n2251) );
  INV_X1 U2668 ( .A(n3992), .ZN(n2252) );
  NAND2_X1 U2669 ( .A1(n3040), .A2(n2382), .ZN(n2381) );
  INV_X1 U2670 ( .A(n3054), .ZN(n2244) );
  INV_X1 U2671 ( .A(n3053), .ZN(n2243) );
  AND2_X1 U2672 ( .A1(n3633), .A2(n2149), .ZN(n2357) );
  NOR2_X1 U2673 ( .A1(n2735), .A2(n4812), .ZN(n2188) );
  OAI21_X1 U2674 ( .B1(n3990), .B2(n2248), .A(n2246), .ZN(n3928) );
  NOR2_X1 U2675 ( .A1(n2668), .A2(n2501), .ZN(n2189) );
  INV_X1 U2676 ( .A(n4223), .ZN(n2322) );
  INV_X1 U2677 ( .A(n3248), .ZN(n2271) );
  NOR2_X1 U2678 ( .A1(n2932), .A2(n2443), .ZN(n2442) );
  NAND2_X1 U2679 ( .A1(n2806), .A2(n3805), .ZN(n2443) );
  NOR2_X1 U2680 ( .A1(n4175), .A2(n4063), .ZN(n2399) );
  NOR2_X1 U2681 ( .A1(n2725), .A2(n4658), .ZN(n2709) );
  AND2_X1 U2682 ( .A1(n3767), .A2(n3765), .ZN(n4156) );
  INV_X1 U2683 ( .A(n2469), .ZN(n2429) );
  INV_X1 U2684 ( .A(n3314), .ZN(n4118) );
  NAND2_X1 U2685 ( .A1(n2445), .A2(n2805), .ZN(n2444) );
  OAI21_X1 U2686 ( .B1(n2444), .B2(n3805), .A(n2806), .ZN(n2437) );
  NAND2_X1 U2687 ( .A1(n4258), .A2(n2399), .ZN(n2398) );
  INV_X1 U2688 ( .A(n2402), .ZN(n2401) );
  NOR2_X1 U2689 ( .A1(n4516), .A2(n4334), .ZN(n2319) );
  AND2_X1 U2690 ( .A1(n2142), .A2(n4411), .ZN(n2306) );
  INV_X1 U2691 ( .A(IR_REG_6__SCAN_IN), .ZN(n2595) );
  INV_X1 U2692 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2761) );
  INV_X1 U2693 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2635) );
  NAND2_X1 U2694 ( .A1(n2362), .A2(n2149), .ZN(n2361) );
  INV_X1 U2695 ( .A(n3654), .ZN(n2362) );
  NAND2_X1 U2696 ( .A1(n2414), .A2(n4621), .ZN(n2413) );
  NAND2_X1 U2697 ( .A1(n2415), .A2(n2412), .ZN(n2411) );
  NOR2_X1 U2698 ( .A1(n4958), .A2(n2414), .ZN(n2412) );
  NAND2_X1 U2699 ( .A1(n2352), .A2(n3105), .ZN(n2351) );
  NAND2_X1 U2700 ( .A1(n2498), .A2(REG3_REG_5__SCAN_IN), .ZN(n4618) );
  NAND2_X1 U2701 ( .A1(n2366), .A2(n2363), .ZN(n2364) );
  NAND2_X1 U2702 ( .A1(n2370), .A2(n2983), .ZN(n2369) );
  INV_X1 U2703 ( .A(n2984), .ZN(n2370) );
  NAND2_X1 U2704 ( .A1(n2499), .A2(REG3_REG_8__SCAN_IN), .ZN(n2622) );
  INV_X1 U2705 ( .A(n2608), .ZN(n2499) );
  NAND2_X1 U2706 ( .A1(n2500), .A2(REG3_REG_9__SCAN_IN), .ZN(n2636) );
  INV_X1 U2707 ( .A(n2622), .ZN(n2500) );
  NAND2_X1 U2708 ( .A1(n2378), .A2(n3069), .ZN(n3963) );
  NAND2_X1 U2709 ( .A1(n3892), .A2(n3893), .ZN(n2378) );
  NAND2_X1 U2710 ( .A1(n2709), .A2(REG3_REG_19__SCAN_IN), .ZN(n2735) );
  AND2_X1 U2711 ( .A1(n3037), .A2(n3036), .ZN(n3971) );
  INV_X1 U2712 ( .A(n2189), .ZN(n2680) );
  NAND2_X1 U2713 ( .A1(n2957), .A2(n2956), .ZN(n2958) );
  OR2_X1 U2714 ( .A1(n3382), .A2(n2955), .ZN(n2956) );
  INV_X1 U2715 ( .A(n2240), .ZN(n3058) );
  OR2_X1 U2716 ( .A1(n3106), .A2(n3853), .ZN(n3109) );
  INV_X1 U2717 ( .A(n3116), .ZN(n3126) );
  NAND2_X1 U2718 ( .A1(n2189), .A2(REG3_REG_14__SCAN_IN), .ZN(n2686) );
  OR2_X1 U2719 ( .A1(n2812), .A2(REG3_REG_3__SCAN_IN), .ZN(n2553) );
  NOR2_X1 U2720 ( .A1(n3185), .A2(n3184), .ZN(n3186) );
  INV_X1 U2721 ( .A(n3183), .ZN(n3185) );
  NAND2_X1 U2722 ( .A1(n3303), .A2(n3304), .ZN(n3302) );
  AND2_X1 U2723 ( .A1(n3191), .A2(n3230), .ZN(n2324) );
  NAND2_X1 U2724 ( .A1(n2275), .A2(n2286), .ZN(n3240) );
  NOR2_X1 U2725 ( .A1(n2288), .A2(n4850), .ZN(n2274) );
  XNOR2_X1 U2726 ( .A(n3240), .B(n3675), .ZN(n3672) );
  NAND2_X1 U2727 ( .A1(n4240), .A2(n2271), .ZN(n2270) );
  OR2_X1 U2728 ( .A1(n4978), .A2(n2173), .ZN(n2326) );
  OAI211_X1 U2729 ( .C1(n4977), .C2(n2172), .A(n2329), .B(n2328), .ZN(n4234)
         );
  AOI21_X1 U2730 ( .B1(n2330), .B2(n2173), .A(n2144), .ZN(n2329) );
  AND2_X1 U2731 ( .A1(n2331), .A2(n3273), .ZN(n2330) );
  INV_X1 U2732 ( .A(REG3_REG_15__SCAN_IN), .ZN(n4761) );
  INV_X1 U2733 ( .A(n2289), .ZN(n3251) );
  INV_X1 U2734 ( .A(n5008), .ZN(n2278) );
  OR2_X1 U2735 ( .A1(n5006), .A2(n2280), .ZN(n2276) );
  INV_X1 U2736 ( .A(n2399), .ZN(n2397) );
  NOR2_X1 U2737 ( .A1(n2194), .A2(n2402), .ZN(n2190) );
  NAND2_X1 U2738 ( .A1(n2386), .A2(n2384), .ZN(n4292) );
  NAND2_X1 U2739 ( .A1(n4325), .A2(n4312), .ZN(n2219) );
  NAND2_X1 U2740 ( .A1(n2215), .A2(n2391), .ZN(n4348) );
  AOI21_X1 U2741 ( .B1(n2454), .B2(n2457), .A(n2451), .ZN(n2450) );
  INV_X1 U2742 ( .A(n4085), .ZN(n2451) );
  OR2_X1 U2743 ( .A1(n4427), .A2(n2708), .ZN(n2453) );
  AND2_X1 U2744 ( .A1(n2517), .A2(n2516), .ZN(n4010) );
  NAND2_X1 U2745 ( .A1(n3784), .A2(n4045), .ZN(n4444) );
  AOI21_X1 U2746 ( .B1(n2138), .B2(n2676), .A(n2162), .ZN(n2446) );
  INV_X1 U2747 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2645) );
  AOI21_X1 U2748 ( .B1(n4144), .B2(n4138), .A(n2213), .ZN(n2212) );
  NAND2_X1 U2749 ( .A1(n2433), .A2(n2431), .ZN(n3680) );
  NAND2_X1 U2750 ( .A1(n2434), .A2(n2469), .ZN(n2433) );
  INV_X1 U2751 ( .A(n3703), .ZN(n3612) );
  NAND2_X1 U2752 ( .A1(n2418), .A2(n2619), .ZN(n2417) );
  NAND2_X1 U2753 ( .A1(n2588), .A2(REG3_REG_7__SCAN_IN), .ZN(n2608) );
  NAND2_X1 U2754 ( .A1(n4056), .A2(n3276), .ZN(n2177) );
  NAND2_X1 U2755 ( .A1(n2200), .A2(n2198), .ZN(n3576) );
  INV_X1 U2756 ( .A(n2199), .ZN(n2198) );
  OAI21_X1 U2757 ( .B1(n2204), .B2(n2203), .A(n4130), .ZN(n2199) );
  NAND2_X1 U2758 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2570) );
  CLKBUF_X1 U2759 ( .A(n3399), .Z(n3400) );
  OR2_X1 U2760 ( .A1(n2550), .A2(n2519), .ZN(n2521) );
  INV_X1 U2761 ( .A(n3839), .ZN(n3128) );
  NOR2_X2 U2762 ( .A1(n4263), .A2(n4482), .ZN(n4264) );
  INV_X1 U2763 ( .A(n4493), .ZN(n4285) );
  NAND2_X1 U2764 ( .A1(n4377), .A2(n2317), .ZN(n4319) );
  NAND2_X1 U2765 ( .A1(n4377), .A2(n2319), .ZN(n4336) );
  NAND2_X1 U2766 ( .A1(n4377), .A2(n4350), .ZN(n4352) );
  NAND2_X1 U2767 ( .A1(n3786), .A2(n2306), .ZN(n4410) );
  NAND2_X1 U2768 ( .A1(n3786), .A2(n2142), .ZN(n4429) );
  AND2_X1 U2769 ( .A1(n3786), .A2(n4550), .ZN(n4450) );
  INV_X1 U2770 ( .A(n4455), .ZN(n4550) );
  NOR2_X1 U2771 ( .A1(n2139), .A2(n3976), .ZN(n2315) );
  NOR2_X1 U2772 ( .A1(n3609), .A2(n2139), .ZN(n3776) );
  NAND2_X1 U2773 ( .A1(n2314), .A2(n2316), .ZN(n3753) );
  NAND2_X1 U2774 ( .A1(n2314), .A2(n3644), .ZN(n3688) );
  AND4_X1 U2775 ( .A1(n2651), .A2(n2650), .A3(n2649), .A4(n2648), .ZN(n3722)
         );
  NOR2_X2 U2776 ( .A1(n3575), .A2(n3659), .ZN(n3574) );
  NAND2_X1 U2777 ( .A1(n2305), .A2(n3497), .ZN(n2302) );
  NOR2_X1 U2778 ( .A1(n3406), .A2(n2304), .ZN(n3491) );
  INV_X1 U2779 ( .A(n4561), .ZN(n4590) );
  INV_X1 U2780 ( .A(n4598), .ZN(n5069) );
  INV_X1 U2781 ( .A(n4570), .ZN(n4593) );
  AND3_X1 U2782 ( .A1(n2898), .A2(n2897), .A3(n2909), .ZN(n3174) );
  NAND2_X1 U2783 ( .A1(n2876), .A2(n2875), .ZN(n2878) );
  MUX2_X1 U2784 ( .A(n2873), .B(IR_REG_31__SCAN_IN), .S(n2872), .Z(n2876) );
  CLKBUF_X1 U2785 ( .A(n2874), .Z(n2875) );
  XNOR2_X1 U2786 ( .A(n2702), .B(IR_REG_15__SCAN_IN), .ZN(n3250) );
  INV_X1 U2787 ( .A(IR_REG_13__SCAN_IN), .ZN(n2480) );
  OR2_X1 U2788 ( .A1(n2632), .A2(IR_REG_9__SCAN_IN), .ZN(n2643) );
  INV_X1 U2789 ( .A(IR_REG_7__SCAN_IN), .ZN(n2614) );
  NAND2_X1 U2790 ( .A1(n2524), .A2(n2293), .ZN(n2292) );
  INV_X1 U2791 ( .A(n3090), .ZN(n4317) );
  NAND2_X1 U2792 ( .A1(n2230), .A2(n2234), .ZN(n3717) );
  AND2_X1 U2793 ( .A1(n2235), .A2(n3718), .ZN(n2234) );
  OR2_X1 U2794 ( .A1(n2154), .A2(n2236), .ZN(n2235) );
  NAND2_X1 U2795 ( .A1(n2233), .A2(n2237), .ZN(n3719) );
  NAND2_X1 U2796 ( .A1(n2239), .A2(n2154), .ZN(n2233) );
  OR2_X1 U2797 ( .A1(n3337), .A2(n3007), .ZN(n2967) );
  AND2_X1 U2798 ( .A1(n2375), .A2(n3966), .ZN(n2374) );
  NAND2_X1 U2799 ( .A1(n2376), .A2(n3964), .ZN(n2375) );
  NAND2_X1 U2800 ( .A1(n3025), .A2(n3024), .ZN(n3921) );
  NAND2_X1 U2801 ( .A1(n2253), .A2(n2254), .ZN(n3528) );
  NAND2_X1 U2802 ( .A1(n2367), .A2(n2255), .ZN(n2254) );
  INV_X1 U2803 ( .A(n2368), .ZN(n2255) );
  AND2_X1 U2804 ( .A1(n2732), .A2(n2731), .ZN(n4543) );
  AND3_X1 U2805 ( .A1(n2700), .A2(n2699), .A3(n2698), .ZN(n4435) );
  AND2_X1 U2806 ( .A1(n2769), .A2(n2768), .ZN(n4333) );
  AND2_X1 U2807 ( .A1(n2785), .A2(n2773), .ZN(n4305) );
  INV_X1 U2808 ( .A(n2364), .ZN(n3470) );
  NAND2_X1 U2809 ( .A1(n2366), .A2(n2369), .ZN(n3471) );
  NAND2_X1 U2810 ( .A1(n4056), .A2(DATAI_0_), .ZN(n2225) );
  NAND2_X1 U2811 ( .A1(n2134), .A2(n5060), .ZN(n2175) );
  INV_X1 U2812 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4812) );
  NAND2_X1 U2813 ( .A1(n2380), .A2(n3918), .ZN(n3974) );
  INV_X1 U2814 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4810) );
  NAND2_X1 U2815 ( .A1(n2258), .A2(n3084), .ZN(n3981) );
  AND2_X1 U2816 ( .A1(n3153), .A2(n3341), .ZN(n4025) );
  INV_X1 U2817 ( .A(n4560), .ZN(n4036) );
  NAND2_X1 U2818 ( .A1(n3151), .A2(n3826), .ZN(n4038) );
  NAND2_X1 U2819 ( .A1(n2837), .A2(n2836), .ZN(n4199) );
  INV_X1 U2820 ( .A(n4486), .ZN(n4271) );
  NAND2_X1 U2821 ( .A1(n2791), .A2(n2790), .ZN(n4298) );
  INV_X1 U2822 ( .A(n4333), .ZN(n4201) );
  OR2_X1 U2823 ( .A1(n4354), .A2(n2812), .ZN(n2751) );
  NAND2_X1 U2824 ( .A1(n2741), .A2(n2740), .ZN(n4517) );
  INV_X1 U2825 ( .A(n4543), .ZN(n4438) );
  INV_X1 U2826 ( .A(n4435), .ZN(n4564) );
  INV_X1 U2827 ( .A(n4574), .ZN(n4454) );
  INV_X1 U2828 ( .A(n3722), .ZN(n4591) );
  AND2_X1 U2829 ( .A1(n2574), .A2(n2475), .ZN(n2464) );
  OR2_X1 U2830 ( .A1(n2550), .A2(n2525), .ZN(n2531) );
  OR2_X1 U2831 ( .A1(n3287), .A2(n2943), .ZN(n4209) );
  NAND2_X1 U2832 ( .A1(n4218), .A2(n3217), .ZN(n4217) );
  NOR2_X1 U2833 ( .A1(n3366), .A2(n5077), .ZN(n3365) );
  INV_X1 U2834 ( .A(n2323), .ZN(n3417) );
  NAND2_X1 U2835 ( .A1(n3232), .A2(n2284), .ZN(n3420) );
  NAND2_X1 U2836 ( .A1(n3390), .A2(REG2_REG_6__SCAN_IN), .ZN(n2284) );
  NAND2_X1 U2837 ( .A1(n3237), .A2(n3236), .ZN(n3598) );
  NAND2_X1 U2838 ( .A1(n3196), .A2(n3195), .ZN(n3597) );
  NAND2_X1 U2839 ( .A1(n4224), .A2(n4223), .ZN(n4222) );
  NAND2_X1 U2840 ( .A1(n3201), .A2(n3200), .ZN(n4224) );
  NAND2_X1 U2841 ( .A1(n4977), .A2(n4978), .ZN(n4976) );
  NAND2_X1 U2842 ( .A1(n2327), .A2(n2325), .ZN(n2332) );
  AND2_X1 U2843 ( .A1(n2326), .A2(n3273), .ZN(n2325) );
  OR2_X1 U2844 ( .A1(n4977), .A2(n2173), .ZN(n2327) );
  NAND2_X1 U2845 ( .A1(n4987), .A2(n4988), .ZN(n4986) );
  NAND2_X1 U2846 ( .A1(n2273), .A2(n2185), .ZN(n2266) );
  AND2_X1 U2847 ( .A1(n3248), .A2(n3273), .ZN(n2185) );
  XNOR2_X1 U2848 ( .A(n2289), .B(n4996), .ZN(n4993) );
  NAND2_X1 U2849 ( .A1(n4993), .A2(n4992), .ZN(n4991) );
  INV_X1 U2850 ( .A(n5009), .ZN(n2181) );
  NAND2_X1 U2851 ( .A1(n2339), .A2(n2341), .ZN(n2336) );
  CLKBUF_X1 U2852 ( .A(n4278), .Z(n4279) );
  OAI21_X1 U2853 ( .B1(n2218), .B2(n4425), .A(n2216), .ZN(n4506) );
  INV_X1 U2854 ( .A(n2217), .ZN(n2216) );
  XNOR2_X1 U2855 ( .A(n2219), .B(n4316), .ZN(n2218) );
  OAI21_X1 U2856 ( .B1(n4314), .B2(n4573), .A(n4313), .ZN(n2217) );
  INV_X1 U2857 ( .A(n4526), .ZN(n4382) );
  INV_X1 U2858 ( .A(n4010), .ZN(n4555) );
  NAND2_X1 U2859 ( .A1(n2851), .A2(n4043), .ZN(n3783) );
  NAND2_X1 U2860 ( .A1(n2448), .A2(n2138), .ZN(n3729) );
  OR2_X1 U2861 ( .A1(n3774), .A2(n2676), .ZN(n2448) );
  AND2_X1 U2862 ( .A1(n5032), .A2(n4589), .ZN(n4471) );
  NAND2_X1 U2863 ( .A1(n2202), .A2(n2204), .ZN(n3445) );
  NAND2_X1 U2864 ( .A1(n3433), .A2(n2207), .ZN(n2202) );
  INV_X1 U2865 ( .A(n4467), .ZN(n4433) );
  NAND2_X1 U2866 ( .A1(n2209), .A2(n2844), .ZN(n3486) );
  NAND2_X1 U2867 ( .A1(n2211), .A2(n2210), .ZN(n2209) );
  OR2_X1 U2868 ( .A1(n2722), .A2(n2721), .ZN(n2723) );
  INV_X1 U2869 ( .A(n4458), .ZN(n4473) );
  INV_X1 U2870 ( .A(n4460), .ZN(n4423) );
  INV_X1 U2871 ( .A(n3382), .ZN(n4468) );
  AND2_X1 U2872 ( .A1(n5032), .A2(n4590), .ZN(n4466) );
  AND2_X1 U2873 ( .A1(n5032), .A2(n4570), .ZN(n4467) );
  AND2_X1 U2874 ( .A1(n3321), .A2(n2533), .ZN(n3377) );
  NAND2_X1 U2875 ( .A1(n4485), .A2(n2223), .ZN(n2179) );
  INV_X1 U2876 ( .A(n2224), .ZN(n2223) );
  OAI21_X1 U2877 ( .B1(n4486), .B2(n4573), .A(n4484), .ZN(n2224) );
  INV_X1 U2878 ( .A(n4945), .ZN(n4935) );
  AND2_X1 U2879 ( .A1(n2507), .A2(n2493), .ZN(n2508) );
  INV_X1 U2880 ( .A(IR_REG_30__SCAN_IN), .ZN(n3863) );
  INV_X1 U2881 ( .A(n2878), .ZN(n4947) );
  OAI21_X1 U2882 ( .B1(n2881), .B2(n2869), .A(IR_REG_31__SCAN_IN), .ZN(n2870)
         );
  OR2_X1 U2883 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2869)
         );
  AND2_X1 U2884 ( .A1(n3212), .A2(STATE_REG_SCAN_IN), .ZN(n5049) );
  INV_X1 U2885 ( .A(n4190), .ZN(n4950) );
  INV_X1 U2886 ( .A(DATAI_18_), .ZN(n5051) );
  INV_X1 U2887 ( .A(n3250), .ZN(n5057) );
  AND2_X1 U2888 ( .A1(n2656), .A2(n2662), .ZN(n4953) );
  XNOR2_X1 U2889 ( .A(n2580), .B(IR_REG_5__SCAN_IN), .ZN(n4956) );
  AOI21_X1 U2890 ( .B1(n4608), .B2(n2158), .A(n2349), .ZN(n2348) );
  NOR2_X1 U2891 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_2__SCAN_IN), .ZN(n2349)
         );
  NAND2_X1 U2892 ( .A1(n3123), .A2(n2259), .ZN(n3165) );
  AOI21_X1 U2893 ( .B1(n2183), .B2(n5001), .A(n2180), .ZN(n5013) );
  NAND2_X1 U2894 ( .A1(n2182), .A2(n2181), .ZN(n2180) );
  OAI21_X1 U2895 ( .B1(n5015), .B2(n2297), .A(n2296), .ZN(n2295) );
  NOR2_X1 U2896 ( .A1(n5032), .A2(n2937), .ZN(n2938) );
  OAI21_X1 U2897 ( .B1(n3843), .B2(n4458), .A(n2307), .ZN(U3262) );
  AOI21_X1 U2898 ( .B1(n2312), .B2(n5032), .A(n2309), .ZN(n2308) );
  AND2_X1 U2899 ( .A1(n2152), .A2(n2903), .ZN(n2904) );
  OAI21_X1 U2900 ( .B1(n4887), .B2(n5079), .A(n2220), .ZN(U3545) );
  AOI21_X1 U2901 ( .B1(n2222), .B2(n4582), .A(n2221), .ZN(n2220) );
  NOR2_X1 U2902 ( .A1(n5081), .A2(n4488), .ZN(n2221) );
  INV_X1 U2903 ( .A(n4890), .ZN(n2222) );
  INV_X2 U2904 ( .A(n2979), .ZN(n3035) );
  OAI211_X1 U2905 ( .C1(n2415), .C2(DATAI_1_), .A(n2413), .B(n2411), .ZN(n3318) );
  AND2_X1 U2906 ( .A1(n2147), .A2(n4100), .ZN(n2138) );
  NAND2_X1 U2907 ( .A1(n2492), .A2(n2491), .ZN(n2867) );
  NAND2_X1 U2908 ( .A1(n2316), .A2(n4594), .ZN(n2139) );
  INV_X1 U2909 ( .A(n3567), .ZN(n2303) );
  OR2_X1 U2910 ( .A1(n4298), .A2(n4493), .ZN(n2140) );
  INV_X1 U2911 ( .A(n2452), .ZN(n4362) );
  INV_X1 U2912 ( .A(n4173), .ZN(n2195) );
  INV_X1 U2913 ( .A(n4075), .ZN(n2403) );
  NAND2_X1 U2914 ( .A1(n3137), .A2(n3994), .ZN(n2141) );
  AND2_X1 U2915 ( .A1(n4166), .A2(n4162), .ZN(n4448) );
  NAND2_X2 U2916 ( .A1(n2914), .A2(n4451), .ZN(n5032) );
  INV_X1 U2917 ( .A(n3423), .ZN(n2178) );
  AND2_X1 U2918 ( .A1(n4550), .A2(n4432), .ZN(n2142) );
  AND2_X1 U2919 ( .A1(n2317), .A2(n4303), .ZN(n2143) );
  NOR2_X1 U2920 ( .A1(n2172), .A2(n4978), .ZN(n2144) );
  NOR2_X1 U2921 ( .A1(n3406), .A2(n3405), .ZN(n2145) );
  AND2_X1 U2922 ( .A1(n2270), .A2(REG2_REG_14__SCAN_IN), .ZN(n2146) );
  NAND2_X4 U2923 ( .A1(n2947), .A2(n3143), .ZN(n3007) );
  NAND2_X1 U2924 ( .A1(n4588), .A2(n3976), .ZN(n2147) );
  AND2_X1 U2925 ( .A1(n3087), .A2(n3084), .ZN(n2148) );
  NAND2_X1 U2926 ( .A1(n3004), .A2(n3003), .ZN(n2149) );
  AND2_X1 U2927 ( .A1(n2258), .A2(n2148), .ZN(n2150) );
  NAND2_X1 U2928 ( .A1(n3018), .A2(n3017), .ZN(n2151) );
  NAND4_X1 U2929 ( .A1(n2531), .A2(n2530), .A3(n2529), .A4(n2528), .ZN(n2963)
         );
  AND2_X1 U2930 ( .A1(n2479), .A2(n2136), .ZN(n2823) );
  OR2_X1 U2931 ( .A1(n3843), .A2(n4873), .ZN(n2152) );
  OR2_X1 U2932 ( .A1(n3843), .A2(n4945), .ZN(n2153) );
  AND2_X1 U2933 ( .A1(n2356), .A2(n2151), .ZN(n2154) );
  NOR2_X1 U2934 ( .A1(n3058), .A2(n3057), .ZN(n4004) );
  INV_X1 U2935 ( .A(n4049), .ZN(n2389) );
  INV_X1 U2936 ( .A(n3105), .ZN(n3954) );
  NAND2_X1 U2937 ( .A1(n2453), .A2(n2460), .ZN(n2452) );
  AND2_X1 U2938 ( .A1(n3093), .A2(n2256), .ZN(n2155) );
  AND2_X1 U2939 ( .A1(n3963), .A2(n3964), .ZN(n2156) );
  XNOR2_X1 U2940 ( .A(n2958), .B(n3007), .ZN(n2960) );
  AND2_X1 U2941 ( .A1(n3852), .A2(n3104), .ZN(n2157) );
  INV_X1 U2942 ( .A(n2843), .ZN(n2210) );
  AND2_X1 U2943 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_2__SCAN_IN), .ZN(n2158)
         );
  NOR2_X1 U2944 ( .A1(n4994), .A2(n3208), .ZN(n2159) );
  AND2_X1 U2945 ( .A1(n4298), .A2(n4493), .ZN(n2160) );
  INV_X1 U2946 ( .A(n2194), .ZN(n2193) );
  OAI21_X1 U2947 ( .B1(n2384), .B2(n2195), .A(n4077), .ZN(n2194) );
  AND2_X1 U2948 ( .A1(n2252), .A2(n2251), .ZN(n2161) );
  AND2_X1 U2949 ( .A1(n4562), .A2(n3880), .ZN(n2162) );
  AND2_X1 U2950 ( .A1(n3722), .A2(n3689), .ZN(n2163) );
  INV_X1 U2951 ( .A(n2707), .ZN(n2708) );
  AND2_X1 U2952 ( .A1(n4078), .A2(n4291), .ZN(n4173) );
  INV_X1 U2953 ( .A(n3999), .ZN(n3689) );
  INV_X1 U2954 ( .A(n4063), .ZN(n2404) );
  INV_X1 U2955 ( .A(n2261), .ZN(n2260) );
  NAND2_X1 U2956 ( .A1(n2262), .A2(n4017), .ZN(n2261) );
  INV_X1 U2957 ( .A(IR_REG_26__SCAN_IN), .ZN(n2872) );
  INV_X1 U2958 ( .A(n2249), .ZN(n2248) );
  AND2_X1 U2959 ( .A1(n2379), .A2(n2250), .ZN(n2249) );
  INV_X1 U2960 ( .A(IR_REG_31__SCAN_IN), .ZN(n2293) );
  AND3_X1 U2961 ( .A1(n2491), .A2(n2506), .A3(n2872), .ZN(n2164) );
  INV_X1 U2962 ( .A(n3806), .ZN(n2445) );
  NOR2_X1 U2963 ( .A1(n2432), .A2(n2468), .ZN(n2431) );
  XNOR2_X1 U2964 ( .A(n2971), .B(n3007), .ZN(n2973) );
  OR2_X1 U2965 ( .A1(n4454), .A2(n4036), .ZN(n2165) );
  AND2_X1 U2966 ( .A1(n2381), .A2(n2471), .ZN(n2166) );
  AND2_X1 U2967 ( .A1(n2398), .A2(n2917), .ZN(n2167) );
  INV_X1 U2968 ( .A(n2409), .ZN(n2408) );
  NAND2_X1 U2969 ( .A1(n4137), .A2(n2410), .ZN(n2409) );
  INV_X1 U2970 ( .A(IR_REG_28__SCAN_IN), .ZN(n2493) );
  INV_X1 U2971 ( .A(n4128), .ZN(n2203) );
  NOR2_X1 U2972 ( .A1(n3787), .A2(n4036), .ZN(n3786) );
  AND2_X1 U2973 ( .A1(n3574), .A2(n3637), .ZN(n3540) );
  NAND2_X1 U2974 ( .A1(n2995), .A2(n2461), .ZN(n3653) );
  INV_X1 U2975 ( .A(n2844), .ZN(n2208) );
  NAND2_X1 U2976 ( .A1(n3717), .A2(n3022), .ZN(n3990) );
  NAND2_X1 U2977 ( .A1(n2239), .A2(n2356), .ZN(n3697) );
  NAND2_X1 U2978 ( .A1(n2358), .A2(n2361), .ZN(n3631) );
  INV_X1 U2979 ( .A(n4516), .ZN(n4350) );
  INV_X1 U2980 ( .A(n4399), .ZN(n2902) );
  AND2_X1 U2981 ( .A1(n2416), .A2(n2420), .ZN(n3545) );
  INV_X1 U2982 ( .A(n3976), .ZN(n3775) );
  INV_X1 U2983 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2186) );
  AND2_X1 U2984 ( .A1(n2364), .A2(n2368), .ZN(n2168) );
  INV_X1 U2985 ( .A(n4411), .ZN(n4415) );
  AND2_X1 U2986 ( .A1(n2306), .A2(n4399), .ZN(n2169) );
  AND2_X1 U2987 ( .A1(n2448), .A2(n2147), .ZN(n2170) );
  AND2_X1 U2988 ( .A1(n2433), .A2(n2430), .ZN(n2171) );
  NOR2_X1 U2989 ( .A1(n2949), .A2(n3405), .ZN(n2305) );
  AND2_X2 U2990 ( .A1(n3174), .A2(n3173), .ZN(n5076) );
  OR2_X1 U2991 ( .A1(n3406), .A2(n2302), .ZN(n3454) );
  AND2_X2 U2992 ( .A1(n3174), .A2(n3132), .ZN(n5081) );
  OR2_X1 U2993 ( .A1(n2173), .A2(n3273), .ZN(n2172) );
  INV_X1 U2994 ( .A(n3918), .ZN(n2382) );
  AND2_X1 U2995 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3247), .ZN(n2173) );
  NAND2_X1 U2996 ( .A1(n4099), .A2(n3322), .ZN(n3321) );
  NAND2_X1 U2997 ( .A1(n3321), .A2(n2426), .ZN(n3376) );
  INV_X1 U2998 ( .A(n2207), .ZN(n2206) );
  NOR2_X1 U2999 ( .A1(n4129), .A2(n2208), .ZN(n2207) );
  INV_X1 U3000 ( .A(n2340), .ZN(n2339) );
  NOR2_X1 U3001 ( .A1(n2466), .A2(n2341), .ZN(n2340) );
  OR2_X1 U3002 ( .A1(n3254), .A2(REG2_REG_17__SCAN_IN), .ZN(n2300) );
  INV_X1 U3003 ( .A(n2280), .ZN(n2279) );
  OR2_X1 U3004 ( .A1(n5016), .A2(n3253), .ZN(n2280) );
  NOR2_X1 U3005 ( .A1(n3365), .A2(n2465), .ZN(n2174) );
  NAND2_X1 U3006 ( .A1(n2863), .A2(n4577), .ZN(n3846) );
  INV_X1 U3007 ( .A(n4577), .ZN(n4425) );
  INV_X1 U3008 ( .A(n2295), .ZN(n5023) );
  NAND2_X1 U3009 ( .A1(n4991), .A2(n3252), .ZN(n5006) );
  NOR2_X1 U3010 ( .A1(n4983), .A2(n4982), .ZN(n4981) );
  NAND2_X1 U3011 ( .A1(n3227), .A2(n3226), .ZN(n3303) );
  NAND2_X1 U3012 ( .A1(n2299), .A2(n5016), .ZN(n2298) );
  NAND2_X1 U3013 ( .A1(n4217), .A2(n3218), .ZN(n3350) );
  MUX2_X2 U3014 ( .A(n4888), .B(n4887), .S(n5076), .Z(n4889) );
  INV_X1 U3015 ( .A(n3322), .ZN(n2424) );
  NAND2_X1 U3016 ( .A1(n2425), .A2(n2422), .ZN(n3399) );
  AOI21_X2 U3017 ( .B1(n2792), .B2(n2140), .A(n2160), .ZN(n3808) );
  OAI21_X2 U3018 ( .B1(n3608), .B2(n2634), .A(n2176), .ZN(n3643) );
  AOI22_X1 U3019 ( .A1(n4346), .A2(n2752), .B1(n4530), .B2(n4350), .ZN(n4341)
         );
  AOI21_X1 U3020 ( .B1(n4487), .B2(n4598), .A(n2179), .ZN(n4887) );
  NAND2_X1 U3021 ( .A1(n3350), .A2(n3351), .ZN(n3349) );
  INV_X1 U3022 ( .A(n2287), .ZN(n2286) );
  XNOR2_X2 U3023 ( .A(n3194), .B(n4955), .ZN(n3509) );
  XNOR2_X2 U3024 ( .A(n3199), .B(n3675), .ZN(n3671) );
  NOR2_X1 U3025 ( .A1(n4995), .A2(REG1_REG_16__SCAN_IN), .ZN(n4994) );
  NAND2_X1 U3026 ( .A1(n3167), .A2(n3168), .ZN(n3175) );
  AOI21_X2 U3027 ( .B1(n2929), .B2(n4577), .A(n2928), .ZN(n3167) );
  NOR2_X2 U3028 ( .A1(n4618), .A2(n2186), .ZN(n2588) );
  NAND2_X1 U3029 ( .A1(n4258), .A2(n2401), .ZN(n2400) );
  NAND2_X1 U3030 ( .A1(n2438), .A2(n2436), .ZN(n2934) );
  NAND2_X1 U3031 ( .A1(n2191), .A2(n2190), .ZN(n2196) );
  INV_X1 U3032 ( .A(n2386), .ZN(n2192) );
  NAND2_X1 U3033 ( .A1(n3433), .A2(n2201), .ZN(n2200) );
  OAI21_X1 U3034 ( .B1(n3606), .B2(n4144), .A(n4138), .ZN(n3642) );
  NAND2_X1 U3035 ( .A1(n2214), .A2(n2212), .ZN(n2848) );
  NAND2_X1 U3036 ( .A1(n3606), .A2(n4138), .ZN(n2214) );
  NAND2_X1 U3037 ( .A1(n4368), .A2(n4049), .ZN(n2215) );
  NAND4_X1 U3038 ( .A1(n2229), .A2(n2228), .A3(n2227), .A4(n2477), .ZN(n2487)
         );
  NAND3_X1 U3039 ( .A1(n2995), .A2(n2461), .A3(n2357), .ZN(n2239) );
  NAND3_X1 U3040 ( .A1(n2995), .A2(n2461), .A3(n2231), .ZN(n2230) );
  OAI21_X1 U3041 ( .B1(n3990), .B2(n2245), .A(n2241), .ZN(n2240) );
  NAND3_X1 U3042 ( .A1(n2366), .A2(n2363), .A3(n2367), .ZN(n2253) );
  NAND2_X1 U3043 ( .A1(n3910), .A2(n2148), .ZN(n2257) );
  NAND2_X2 U3044 ( .A1(n2257), .A2(n2155), .ZN(n3851) );
  NAND2_X1 U3045 ( .A1(n3123), .A2(n2260), .ZN(n3142) );
  NAND2_X1 U3046 ( .A1(n3123), .A2(n4017), .ZN(n3866) );
  NAND4_X1 U3047 ( .A1(n2490), .A2(n2263), .A3(n2136), .A4(n2508), .ZN(n3862)
         );
  NAND3_X1 U3048 ( .A1(n2263), .A2(n2490), .A3(n2136), .ZN(n2395) );
  AND2_X2 U3049 ( .A1(n2822), .A2(n2164), .ZN(n2263) );
  MUX2_X1 U3050 ( .A(n3216), .B(REG2_REG_1__SCAN_IN), .S(n4210), .Z(n4218) );
  OR2_X2 U3051 ( .A1(n4972), .A2(n4970), .ZN(n2273) );
  NAND3_X1 U3052 ( .A1(n2267), .A2(n2146), .A3(n2268), .ZN(n2272) );
  NAND2_X1 U3053 ( .A1(n2273), .A2(n2269), .ZN(n2268) );
  NAND3_X1 U3054 ( .A1(n2268), .A2(n2267), .A3(n2270), .ZN(n4236) );
  INV_X1 U3055 ( .A(n2272), .ZN(n4235) );
  NAND2_X1 U3056 ( .A1(n3510), .A2(n2274), .ZN(n2275) );
  NAND2_X1 U3057 ( .A1(n5006), .A2(n5008), .ZN(n5007) );
  AND2_X1 U3058 ( .A1(n3255), .A2(REG2_REG_18__SCAN_IN), .ZN(n2281) );
  INV_X1 U3059 ( .A(n3232), .ZN(n2283) );
  OAI21_X1 U3060 ( .B1(n3390), .B2(n2283), .A(n2282), .ZN(n3418) );
  OR2_X2 U3061 ( .A1(n4981), .A2(n2290), .ZN(n2289) );
  NAND3_X1 U3062 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .A3(
        IR_REG_0__SCAN_IN), .ZN(n2291) );
  NAND2_X2 U3063 ( .A1(n3246), .A2(n3245), .ZN(n4972) );
  NAND3_X1 U3064 ( .A1(n2305), .A2(n2303), .A3(n3497), .ZN(n2301) );
  INV_X1 U3065 ( .A(n2305), .ZN(n2304) );
  INV_X1 U3066 ( .A(n3609), .ZN(n2314) );
  NAND2_X1 U3067 ( .A1(n2314), .A2(n2315), .ZN(n3778) );
  NOR2_X2 U3068 ( .A1(n3295), .A2(n3413), .ZN(n3294) );
  XNOR2_X2 U3069 ( .A(n3183), .B(n4957), .ZN(n3295) );
  XNOR2_X1 U3070 ( .A(n3203), .B(n3800), .ZN(n3796) );
  OAI21_X2 U3071 ( .B1(n3201), .B2(n2322), .A(n2320), .ZN(n3203) );
  OR2_X2 U3072 ( .A1(n3393), .A2(n2324), .ZN(n2323) );
  NOR2_X1 U3073 ( .A1(n3394), .A2(n3457), .ZN(n3393) );
  NAND2_X1 U3074 ( .A1(n4977), .A2(n2330), .ZN(n2328) );
  OR2_X1 U3075 ( .A1(n4978), .A2(n2173), .ZN(n2331) );
  OAI211_X1 U3076 ( .C1(n5019), .C2(n2336), .A(n3215), .B(n2333), .ZN(n2334)
         );
  NAND2_X1 U3077 ( .A1(n3264), .A2(n2334), .ZN(U3259) );
  XNOR2_X2 U3078 ( .A(n3207), .B(n5054), .ZN(n4995) );
  XNOR2_X2 U3079 ( .A(n3187), .B(n3369), .ZN(n3366) );
  XNOR2_X1 U3080 ( .A(n2350), .B(n3855), .ZN(n3856) );
  NAND2_X1 U3081 ( .A1(n2353), .A2(n2351), .ZN(n2350) );
  INV_X1 U3082 ( .A(n3952), .ZN(n2352) );
  AND2_X2 U3083 ( .A1(n3851), .A2(n3848), .ZN(n3952) );
  INV_X1 U3084 ( .A(n3953), .ZN(n2353) );
  AOI21_X1 U3085 ( .B1(n3851), .B2(n3850), .A(n3849), .ZN(n3953) );
  NOR2_X2 U3086 ( .A1(n2487), .A2(n2355), .ZN(n2490) );
  NAND4_X1 U3087 ( .A1(n2485), .A2(n2486), .A3(n2825), .A4(n2883), .ZN(n2355)
         );
  NAND3_X1 U3088 ( .A1(n2995), .A2(n2461), .A3(n2149), .ZN(n2358) );
  NOR2_X1 U3089 ( .A1(n3472), .A2(n2365), .ZN(n2363) );
  NAND2_X1 U3090 ( .A1(n3892), .A2(n2372), .ZN(n2371) );
  NAND2_X1 U3091 ( .A1(n2371), .A2(n2374), .ZN(n3910) );
  NAND3_X1 U3092 ( .A1(n3025), .A2(n3024), .A3(n2383), .ZN(n2380) );
  NAND2_X1 U3093 ( .A1(n4368), .A2(n2387), .ZN(n2386) );
  NAND3_X1 U3094 ( .A1(n2490), .A2(n2136), .A3(n2822), .ZN(n2865) );
  OAI21_X2 U3095 ( .B1(n2395), .B2(IR_REG_28__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2510) );
  NAND2_X1 U3096 ( .A1(n2396), .A2(n2398), .ZN(n4261) );
  OR2_X2 U3097 ( .A1(n4276), .A2(n2400), .ZN(n2396) );
  NAND2_X1 U3098 ( .A1(n2396), .A2(n2167), .ZN(n2860) );
  OR2_X1 U3099 ( .A1(n4276), .A2(n4075), .ZN(n3809) );
  OAI21_X1 U3100 ( .B1(n3576), .B2(n2409), .A(n2405), .ZN(n3606) );
  OAI21_X1 U3101 ( .B1(n3576), .B2(n2846), .A(n4136), .ZN(n3539) );
  NAND2_X1 U3102 ( .A1(n2846), .A2(n4136), .ZN(n2410) );
  NAND2_X1 U3103 ( .A1(n4465), .A2(n3318), .ZN(n4116) );
  NAND2_X4 U3104 ( .A1(n2415), .A2(n2496), .ZN(n4056) );
  NAND2_X2 U3105 ( .A1(n2495), .A2(n2494), .ZN(n2415) );
  NAND4_X1 U3106 ( .A1(n2582), .A2(n2581), .A3(n2605), .A4(n2619), .ZN(n2419)
         );
  NAND3_X1 U3107 ( .A1(n2582), .A2(n2581), .A3(n2605), .ZN(n2416) );
  OAI211_X1 U3108 ( .C1(n2420), .C2(n2620), .A(n2419), .B(n2417), .ZN(n3608)
         );
  NAND3_X1 U3109 ( .A1(n2605), .A2(n3447), .A3(n2586), .ZN(n2420) );
  NAND2_X2 U3110 ( .A1(n2874), .A2(IR_REG_31__SCAN_IN), .ZN(n2923) );
  NAND2_X1 U3111 ( .A1(n2492), .A2(n2421), .ZN(n2874) );
  NAND3_X1 U3112 ( .A1(n2424), .A2(n4091), .A3(n2533), .ZN(n2423) );
  INV_X1 U3113 ( .A(n3643), .ZN(n2434) );
  NAND2_X1 U3114 ( .A1(n2427), .A2(n2428), .ZN(n3752) );
  NAND2_X1 U3115 ( .A1(n3643), .A2(n2431), .ZN(n2427) );
  INV_X1 U3116 ( .A(n2470), .ZN(n2432) );
  OR2_X1 U3117 ( .A1(n3808), .A2(n2444), .ZN(n2438) );
  NAND2_X1 U3118 ( .A1(n2435), .A2(n2439), .ZN(n2935) );
  NAND2_X1 U3119 ( .A1(n3808), .A2(n2442), .ZN(n2435) );
  AOI21_X1 U3120 ( .B1(n3808), .B2(n3805), .A(n3806), .ZN(n4257) );
  NAND2_X1 U3121 ( .A1(n3774), .A2(n2138), .ZN(n2447) );
  NAND2_X1 U3122 ( .A1(n4427), .A2(n2454), .ZN(n2449) );
  NAND2_X1 U3123 ( .A1(n2449), .A2(n2450), .ZN(n4346) );
  INV_X1 U3124 ( .A(n2743), .ZN(n2459) );
  OAI21_X1 U3125 ( .B1(n2931), .B2(n2930), .A(n5032), .ZN(n2940) );
  NOR2_X1 U3126 ( .A1(n2472), .A2(n2938), .ZN(n2939) );
  INV_X1 U3127 ( .A(n2906), .ZN(n2907) );
  OR2_X1 U3128 ( .A1(n2907), .A2(n2925), .ZN(n2908) );
  NAND2_X1 U3129 ( .A1(n2907), .A2(n2925), .ZN(n4251) );
  NAND2_X1 U3130 ( .A1(n2901), .A2(n3382), .ZN(n3406) );
  INV_X1 U3131 ( .A(n3386), .ZN(n2901) );
  AND2_X1 U3132 ( .A1(n4056), .A2(DATAI_26_), .ZN(n4019) );
  AND2_X1 U3133 ( .A1(n4056), .A2(DATAI_25_), .ZN(n4493) );
  AND2_X1 U3134 ( .A1(n2133), .A2(DATAI_24_), .ZN(n3957) );
  AND2_X1 U3135 ( .A1(n4056), .A2(DATAI_21_), .ZN(n4516) );
  AND2_X1 U3136 ( .A1(n4056), .A2(DATAI_20_), .ZN(n4526) );
  NAND2_X1 U3137 ( .A1(n2133), .A2(n2544), .ZN(n2545) );
  OR2_X1 U3138 ( .A1(n3521), .A2(n2993), .ZN(n2461) );
  AND2_X1 U3139 ( .A1(n3160), .A2(n3141), .ZN(n2462) );
  AND3_X1 U3140 ( .A1(n2719), .A2(n2718), .A3(n2717), .ZN(n2463) );
  INV_X1 U3141 ( .A(n3007), .ZN(n2998) );
  INV_X1 U3142 ( .A(n4997), .ZN(n3215) );
  INV_X1 U3143 ( .A(n4041), .ZN(n3994) );
  NAND2_X1 U3144 ( .A1(n3144), .A2(n3136), .ZN(n4041) );
  OR2_X1 U3145 ( .A1(n5052), .A2(n4827), .ZN(n2466) );
  INV_X1 U3146 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3266) );
  OR2_X1 U3147 ( .A1(n3567), .A2(n3582), .ZN(n2467) );
  AND2_X1 U31480 ( .A1(n3693), .A2(n3725), .ZN(n2468) );
  OR2_X1 U31490 ( .A1(n3693), .A2(n3725), .ZN(n2469) );
  NAND2_X1 U3150 ( .A1(n4154), .A2(n4150), .ZN(n2470) );
  AND2_X1 U3151 ( .A1(n2759), .A2(n2758), .ZN(n4520) );
  INV_X1 U3152 ( .A(n4520), .ZN(n4356) );
  INV_X1 U3153 ( .A(n3369), .ZN(n2560) );
  INV_X1 U3154 ( .A(n3345), .ZN(n2546) );
  AND2_X1 U3155 ( .A1(n3043), .A2(n3875), .ZN(n2471) );
  AND2_X1 U3156 ( .A1(n4056), .A2(DATAI_22_), .ZN(n4334) );
  INV_X1 U3157 ( .A(IR_REG_25__SCAN_IN), .ZN(n2491) );
  AND2_X1 U3158 ( .A1(n3166), .A2(n4460), .ZN(n2472) );
  OR2_X1 U3159 ( .A1(n3178), .A2(n4945), .ZN(n2473) );
  OR2_X1 U3160 ( .A1(n3178), .A2(n4873), .ZN(n2474) );
  AND2_X1 U3161 ( .A1(n2573), .A2(n2572), .ZN(n2475) );
  AND2_X1 U3162 ( .A1(n2949), .A2(n3531), .ZN(n2476) );
  OAI21_X1 U3163 ( .B1(n3972), .B2(n3971), .A(n3876), .ZN(n3039) );
  INV_X1 U3164 ( .A(n3318), .ZN(n2968) );
  NAND2_X1 U3165 ( .A1(n4010), .A2(n4432), .ZN(n2707) );
  AND2_X1 U3166 ( .A1(n2859), .A2(n4076), .ZN(n4175) );
  INV_X1 U3167 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4829) );
  INV_X1 U3168 ( .A(n3159), .ZN(n3140) );
  NAND2_X1 U3169 ( .A1(n4056), .A2(n2558), .ZN(n2559) );
  INV_X1 U3170 ( .A(n3982), .ZN(n3087) );
  AND2_X1 U3171 ( .A1(n3109), .A2(n3108), .ZN(n3110) );
  INV_X1 U3172 ( .A(n2619), .ZN(n2620) );
  NAND2_X1 U3173 ( .A1(n3345), .A2(REG2_REG_2__SCAN_IN), .ZN(n3219) );
  NAND2_X1 U3174 ( .A1(n2323), .A2(REG1_REG_7__SCAN_IN), .ZN(n3192) );
  AND2_X1 U3175 ( .A1(n2810), .A2(n2794), .ZN(n4020) );
  NAND2_X1 U3176 ( .A1(n4356), .A2(n4334), .ZN(n2760) );
  NAND2_X1 U3177 ( .A1(n2506), .A2(IR_REG_28__SCAN_IN), .ZN(n2496) );
  OR2_X1 U3178 ( .A1(n2910), .A2(D_REG_1__SCAN_IN), .ZN(n3131) );
  OR2_X1 U3179 ( .A1(n2881), .A2(IR_REG_22__SCAN_IN), .ZN(n2882) );
  INV_X1 U3180 ( .A(n3675), .ZN(n3239) );
  OR2_X1 U3181 ( .A1(n4282), .A2(n2812), .ZN(n2791) );
  AND3_X1 U3182 ( .A1(n2690), .A2(n2689), .A3(n2688), .ZN(n4574) );
  AND2_X1 U3183 ( .A1(n2917), .A2(n4179), .ZN(n4258) );
  INV_X1 U3184 ( .A(n3009), .ZN(n3637) );
  INV_X1 U3185 ( .A(n3534), .ZN(n3497) );
  AND2_X1 U3186 ( .A1(n4125), .A2(n4122), .ZN(n4094) );
  OR2_X1 U3187 ( .A1(n3740), .A2(n4948), .ZN(n2913) );
  OR2_X1 U3188 ( .A1(n4947), .A2(n2879), .ZN(n2899) );
  NAND2_X1 U3189 ( .A1(n4251), .A2(n2908), .ZN(n3178) );
  AND2_X1 U3190 ( .A1(n3213), .A2(n3341), .ZN(n4589) );
  INV_X1 U3191 ( .A(n3577), .ZN(n3659) );
  AOI21_X1 U3192 ( .B1(n2990), .B2(n2989), .A(n3528), .ZN(n3521) );
  OR3_X1 U3193 ( .A1(n3088), .A2(n3287), .A3(n3143), .ZN(n4193) );
  INV_X1 U3194 ( .A(n5014), .ZN(n5001) );
  OR2_X1 U3195 ( .A1(n3807), .A2(n3806), .ZN(n4108) );
  AND2_X1 U3196 ( .A1(n2727), .A2(n2726), .ZN(n4409) );
  AND2_X1 U3197 ( .A1(n5032), .A2(n2936), .ZN(n4460) );
  OR2_X1 U3198 ( .A1(n2913), .A2(n3211), .ZN(n4451) );
  INV_X1 U3199 ( .A(n4873), .ZN(n4582) );
  INV_X1 U3200 ( .A(n3957), .ZN(n4303) );
  INV_X1 U3201 ( .A(n3756), .ZN(n4594) );
  NAND2_X1 U3202 ( .A1(n4188), .A2(n2862), .ZN(n4577) );
  NAND2_X1 U3203 ( .A1(n3323), .A2(n3740), .ZN(n4598) );
  INV_X1 U3204 ( .A(n3132), .ZN(n3173) );
  INV_X1 U3205 ( .A(n5049), .ZN(n3287) );
  XNOR2_X1 U3206 ( .A(n2870), .B(IR_REG_24__SCAN_IN), .ZN(n2879) );
  AND2_X1 U3207 ( .A1(n3260), .A2(n3259), .ZN(n5018) );
  INV_X1 U3208 ( .A(n4025), .ZN(n4034) );
  INV_X1 U3209 ( .A(n4038), .ZN(n4003) );
  NAND2_X1 U32100 ( .A1(n2751), .A2(n2750), .ZN(n4378) );
  OR2_X1 U32110 ( .A1(n4969), .A2(n4192), .ZN(n5014) );
  OR2_X1 U32120 ( .A1(n4969), .A2(n4966), .ZN(n4997) );
  OR2_X1 U32130 ( .A1(n4969), .A2(n4959), .ZN(n5024) );
  INV_X1 U32140 ( .A(n5032), .ZN(n4462) );
  INV_X1 U32150 ( .A(n5032), .ZN(n4337) );
  NAND2_X1 U32160 ( .A1(n3265), .A2(n5081), .ZN(n2905) );
  NAND2_X1 U32170 ( .A1(n5081), .A2(n2941), .ZN(n4873) );
  INV_X1 U32180 ( .A(n5081), .ZN(n5079) );
  NAND2_X1 U32190 ( .A1(n5076), .A2(n2941), .ZN(n4945) );
  INV_X1 U32200 ( .A(n5076), .ZN(n5075) );
  INV_X1 U32210 ( .A(n5048), .ZN(n5047) );
  NAND2_X1 U32220 ( .A1(n2910), .A2(n3827), .ZN(n5048) );
  INV_X1 U32230 ( .A(n3254), .ZN(n5053) );
  AND2_X1 U32240 ( .A1(n2633), .A2(n2643), .ZN(n4954) );
  INV_X1 U32250 ( .A(n4209), .ZN(U4043) );
  NAND2_X1 U32260 ( .A1(n2940), .A2(n2939), .ZN(U3354) );
  NAND2_X1 U32270 ( .A1(n2905), .A2(n2904), .ZN(U3546) );
  INV_X1 U32280 ( .A(n2487), .ZN(n2479) );
  NAND2_X1 U32290 ( .A1(n2823), .A2(n2480), .ZN(n2691) );
  INV_X1 U32300 ( .A(IR_REG_14__SCAN_IN), .ZN(n2482) );
  INV_X1 U32310 ( .A(IR_REG_16__SCAN_IN), .ZN(n2481) );
  NAND2_X1 U32320 ( .A1(n2482), .A2(n2481), .ZN(n2483) );
  NAND2_X1 U32330 ( .A1(n2733), .A2(IR_REG_31__SCAN_IN), .ZN(n2484) );
  INV_X1 U32340 ( .A(DATAI_17_), .ZN(n2497) );
  NOR2_X2 U32350 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2717) );
  AND4_X2 U32360 ( .A1(n2718), .A2(n2717), .A3(n2489), .A4(n2488), .ZN(n2822)
         );
  INV_X1 U32370 ( .A(n2865), .ZN(n2492) );
  NAND2_X1 U32380 ( .A1(n2923), .A2(n2506), .ZN(n2494) );
  MUX2_X1 U32390 ( .A(n5053), .B(n2497), .S(n4056), .Z(n4432) );
  INV_X1 U32400 ( .A(n4432), .ZN(n4541) );
  INV_X1 U32410 ( .A(n2570), .ZN(n2498) );
  OR2_X2 U32420 ( .A1(n2636), .A2(n2635), .ZN(n2646) );
  OR2_X2 U32430 ( .A1(n2646), .A2(n2645), .ZN(n2668) );
  NAND2_X1 U32440 ( .A1(REG3_REG_13__SCAN_IN), .A2(REG3_REG_12__SCAN_IN), .ZN(
        n2501) );
  INV_X1 U32450 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2504) );
  NAND2_X1 U32460 ( .A1(n2697), .A2(n2504), .ZN(n2505) );
  NAND2_X1 U32470 ( .A1(n2725), .A2(n2505), .ZN(n4430) );
  XNOR2_X2 U32480 ( .A(n2509), .B(n3863), .ZN(n2512) );
  INV_X1 U32490 ( .A(n2512), .ZN(n3282) );
  XNOR2_X2 U32500 ( .A(n2510), .B(IR_REG_29__SCAN_IN), .ZN(n3280) );
  OR2_X1 U32510 ( .A1(n4430), .A2(n2812), .ZN(n2517) );
  OR2_X2 U32520 ( .A1(n2512), .A2(n3280), .ZN(n2537) );
  INV_X1 U32530 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4431) );
  INV_X1 U32540 ( .A(n3280), .ZN(n2511) );
  NAND2_X2 U32550 ( .A1(n2511), .A2(n2512), .ZN(n2550) );
  INV_X1 U32560 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4925) );
  OR2_X1 U32570 ( .A1(n3330), .A2(n4925), .ZN(n2514) );
  NAND2_X1 U32580 ( .A1(n3280), .A2(n2512), .ZN(n2551) );
  INV_X1 U32590 ( .A(n2551), .ZN(n2534) );
  INV_X1 U32600 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4547) );
  OR2_X1 U32610 ( .A1(n2748), .A2(n4547), .ZN(n2513) );
  OAI211_X1 U32620 ( .C1(n3334), .C2(n4431), .A(n2514), .B(n2513), .ZN(n2515)
         );
  INV_X1 U32630 ( .A(n2515), .ZN(n2516) );
  INV_X1 U32640 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2518) );
  INV_X1 U32650 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3216) );
  INV_X1 U32660 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U32670 ( .A1(n2534), .A2(REG1_REG_1__SCAN_IN), .ZN(n2520) );
  INV_X2 U32680 ( .A(IR_REG_0__SCAN_IN), .ZN(n2532) );
  INV_X1 U32690 ( .A(IR_REG_1__SCAN_IN), .ZN(n2524) );
  INV_X1 U32700 ( .A(DATAI_1_), .ZN(n4621) );
  INV_X1 U32710 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2525) );
  INV_X1 U32720 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2526) );
  OR2_X1 U32730 ( .A1(n2551), .A2(n2526), .ZN(n2530) );
  INV_X1 U32740 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2527) );
  OR2_X1 U32750 ( .A1(n2536), .A2(n2527), .ZN(n2529) );
  INV_X1 U32760 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4623) );
  OR2_X1 U32770 ( .A1(n2537), .A2(n4623), .ZN(n2528) );
  AND2_X1 U32780 ( .A1(n2963), .A2(n3832), .ZN(n3322) );
  NAND2_X1 U32790 ( .A1(n4465), .A2(n2968), .ZN(n2533) );
  NAND2_X1 U32800 ( .A1(n2534), .A2(REG1_REG_2__SCAN_IN), .ZN(n2541) );
  INV_X1 U32810 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4705) );
  OR2_X1 U32820 ( .A1(n2550), .A2(n4705), .ZN(n2540) );
  INV_X1 U32830 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2535) );
  OR2_X1 U32840 ( .A1(n2536), .A2(n2535), .ZN(n2539) );
  INV_X1 U32850 ( .A(REG2_REG_2__SCAN_IN), .ZN(n4464) );
  OR2_X1 U32860 ( .A1(n2537), .A2(n4464), .ZN(n2538) );
  INV_X1 U32870 ( .A(n4608), .ZN(n2543) );
  INV_X1 U32880 ( .A(IR_REG_2__SCAN_IN), .ZN(n2542) );
  INV_X1 U32890 ( .A(DATAI_2_), .ZN(n2544) );
  OAI21_X2 U32900 ( .B1(n4056), .B2(n2546), .A(n2545), .ZN(n3382) );
  OR2_X2 U32910 ( .A1(n2135), .A2(n3382), .ZN(n4120) );
  NAND2_X1 U32920 ( .A1(n2135), .A2(n3382), .ZN(n4123) );
  NAND2_X2 U32930 ( .A1(n4120), .A2(n4123), .ZN(n4091) );
  OR2_X1 U32940 ( .A1(n2135), .A2(n4468), .ZN(n2547) );
  INV_X1 U32950 ( .A(n3399), .ZN(n2582) );
  NAND2_X1 U32960 ( .A1(n2579), .A2(IR_REG_31__SCAN_IN), .ZN(n2548) );
  NAND2_X1 U32970 ( .A1(n2548), .A2(n2576), .ZN(n2556) );
  OR2_X1 U32980 ( .A1(n2548), .A2(n2576), .ZN(n2549) );
  MUX2_X1 U32990 ( .A(n4957), .B(DATAI_3_), .S(n4056), .Z(n3405) );
  INV_X1 U33000 ( .A(n2550), .ZN(n2920) );
  NAND2_X1 U33010 ( .A1(n2920), .A2(REG0_REG_3__SCAN_IN), .ZN(n2555) );
  INV_X1 U33020 ( .A(REG1_REG_3__SCAN_IN), .ZN(n3413) );
  OR2_X1 U33030 ( .A1(n2551), .A2(n3413), .ZN(n2554) );
  INV_X1 U33040 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3552) );
  OR2_X1 U33050 ( .A1(n2537), .A2(n3552), .ZN(n2552) );
  NAND2_X1 U33060 ( .A1(n2556), .A2(IR_REG_31__SCAN_IN), .ZN(n2557) );
  XNOR2_X1 U33070 ( .A(n2557), .B(n2577), .ZN(n3369) );
  INV_X1 U33080 ( .A(DATAI_4_), .ZN(n2558) );
  OAI21_X1 U33090 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2570), .ZN(n3467) );
  OR2_X1 U33100 ( .A1(n2812), .A2(n3467), .ZN(n2566) );
  INV_X1 U33110 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2561) );
  OR2_X1 U33120 ( .A1(n2550), .A2(n2561), .ZN(n2565) );
  NAND2_X1 U33130 ( .A1(n2534), .A2(REG1_REG_4__SCAN_IN), .ZN(n2564) );
  INV_X1 U33140 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2562) );
  OR2_X1 U33150 ( .A1(n2537), .A2(n2562), .ZN(n2563) );
  NAND4_X2 U33160 ( .A1(n2566), .A2(n2565), .A3(n2564), .A4(n2563), .ZN(n3531)
         );
  NAND2_X2 U33170 ( .A1(n2949), .A2(n2567), .ZN(n4126) );
  NAND2_X1 U33180 ( .A1(n3531), .A2(n2583), .ZN(n2844) );
  NAND2_X2 U33190 ( .A1(n4126), .A2(n2844), .ZN(n4096) );
  OAI21_X1 U33200 ( .B1(n3405), .B2(n4470), .A(n4096), .ZN(n3446) );
  INV_X1 U33210 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2568) );
  OR2_X1 U33220 ( .A1(n2748), .A2(n2568), .ZN(n2575) );
  INV_X1 U33230 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3228) );
  OR2_X1 U33240 ( .A1(n3334), .A2(n3228), .ZN(n2574) );
  NAND2_X1 U33250 ( .A1(n2920), .A2(REG0_REG_5__SCAN_IN), .ZN(n2573) );
  INV_X1 U33260 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2569) );
  NAND2_X1 U33270 ( .A1(n2570), .A2(n2569), .ZN(n2571) );
  NAND2_X1 U33280 ( .A1(n4618), .A2(n2571), .ZN(n3537) );
  OR2_X1 U33290 ( .A1(n2812), .A2(n3537), .ZN(n2572) );
  NAND2_X1 U33300 ( .A1(n2577), .A2(n2576), .ZN(n2578) );
  OAI21_X1 U33310 ( .B1(n2579), .B2(n2578), .A(IR_REG_31__SCAN_IN), .ZN(n2580)
         );
  MUX2_X1 U33320 ( .A(n4956), .B(DATAI_5_), .S(n4056), .Z(n3534) );
  AND2_X1 U33330 ( .A1(n4470), .A2(n3405), .ZN(n2584) );
  INV_X1 U33340 ( .A(n2583), .ZN(n2949) );
  AOI21_X1 U33350 ( .B1(n4096), .B2(n2584), .A(n2476), .ZN(n3488) );
  NAND2_X1 U33360 ( .A1(n4207), .A2(n3534), .ZN(n2585) );
  INV_X1 U33370 ( .A(n3449), .ZN(n2586) );
  NAND2_X1 U33380 ( .A1(n2534), .A2(REG1_REG_7__SCAN_IN), .ZN(n2594) );
  INV_X1 U33390 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2587) );
  OR2_X1 U33400 ( .A1(n2550), .A2(n2587), .ZN(n2593) );
  INV_X1 U33410 ( .A(n2588), .ZN(n2600) );
  INV_X1 U33420 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2589) );
  NAND2_X1 U33430 ( .A1(n2600), .A2(n2589), .ZN(n2590) );
  NAND2_X1 U33440 ( .A1(n2608), .A2(n2590), .ZN(n3662) );
  OR2_X1 U33450 ( .A1(n2812), .A2(n3662), .ZN(n2592) );
  INV_X1 U33460 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3233) );
  OR2_X1 U33470 ( .A1(n2537), .A2(n3233), .ZN(n2591) );
  NAND4_X4 U33480 ( .A1(n2594), .A2(n2593), .A3(n2592), .A4(n2591), .ZN(n4206)
         );
  NAND2_X1 U33490 ( .A1(n2136), .A2(n2595), .ZN(n2628) );
  NAND2_X1 U33500 ( .A1(n2628), .A2(IR_REG_31__SCAN_IN), .ZN(n2615) );
  XNOR2_X1 U33510 ( .A(n2615), .B(n2614), .ZN(n3423) );
  INV_X1 U33520 ( .A(DATAI_7_), .ZN(n3276) );
  OR2_X1 U3353 ( .A1(n4206), .A2(n3577), .ZN(n2845) );
  NAND2_X1 U33540 ( .A1(n2596), .A2(IR_REG_31__SCAN_IN), .ZN(n2597) );
  XNOR2_X1 U3355 ( .A(n2597), .B(IR_REG_6__SCAN_IN), .ZN(n3230) );
  MUX2_X1 U3356 ( .A(n3230), .B(DATAI_6_), .S(n4056), .Z(n3567) );
  NAND2_X1 U3357 ( .A1(n3329), .A2(REG1_REG_6__SCAN_IN), .ZN(n2604) );
  INV_X1 U3358 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2598) );
  OR2_X1 U3359 ( .A1(n3330), .A2(n2598), .ZN(n2603) );
  NAND2_X1 U3360 ( .A1(n4618), .A2(n2186), .ZN(n2599) );
  NAND2_X1 U3361 ( .A1(n2600), .A2(n2599), .ZN(n3562) );
  OR2_X1 U3362 ( .A1(n2812), .A2(n3562), .ZN(n2602) );
  INV_X1 U3363 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3563) );
  OR2_X1 U3364 ( .A1(n3334), .A2(n3563), .ZN(n2601) );
  NAND4_X2 U3365 ( .A1(n2604), .A2(n2603), .A3(n2602), .A4(n2601), .ZN(n3582)
         );
  AND2_X1 U3366 ( .A1(n3582), .A2(n3567), .ZN(n2606) );
  AOI22_X1 U3367 ( .A1(n4131), .A2(n2606), .B1(n3659), .B2(n4206), .ZN(n3546)
         );
  NAND2_X1 U3368 ( .A1(n2813), .A2(REG2_REG_8__SCAN_IN), .ZN(n2613) );
  INV_X1 U3369 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4797) );
  OR2_X1 U3370 ( .A1(n3330), .A2(n4797), .ZN(n2612) );
  INV_X1 U3371 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4796) );
  OR2_X1 U3372 ( .A1(n2748), .A2(n4796), .ZN(n2611) );
  INV_X1 U3373 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2607) );
  NAND2_X1 U3374 ( .A1(n2608), .A2(n2607), .ZN(n2609) );
  NAND2_X1 U3375 ( .A1(n2622), .A2(n2609), .ZN(n3542) );
  OR2_X1 U3376 ( .A1(n2812), .A2(n3542), .ZN(n2610) );
  NAND4_X1 U3377 ( .A1(n2613), .A2(n2612), .A3(n2611), .A4(n2610), .ZN(n4205)
         );
  NAND2_X1 U3378 ( .A1(n2615), .A2(n2614), .ZN(n2616) );
  NAND2_X1 U3379 ( .A1(n2616), .A2(IR_REG_31__SCAN_IN), .ZN(n2617) );
  XNOR2_X1 U3380 ( .A(n2617), .B(IR_REG_8__SCAN_IN), .ZN(n4955) );
  MUX2_X1 U3381 ( .A(n4955), .B(DATAI_8_), .S(n4056), .Z(n3009) );
  NAND2_X1 U3382 ( .A1(n4205), .A2(n3009), .ZN(n2618) );
  OR2_X1 U3383 ( .A1(n4205), .A2(n3009), .ZN(n2619) );
  NAND2_X1 U3384 ( .A1(n2920), .A2(REG0_REG_9__SCAN_IN), .ZN(n2627) );
  INV_X1 U3385 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3197) );
  OR2_X1 U3386 ( .A1(n2748), .A2(n3197), .ZN(n2626) );
  INV_X1 U3387 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2621) );
  NAND2_X1 U3388 ( .A1(n2622), .A2(n2621), .ZN(n2623) );
  NAND2_X1 U3389 ( .A1(n2636), .A2(n2623), .ZN(n3706) );
  OR2_X1 U3390 ( .A1(n2812), .A2(n3706), .ZN(n2625) );
  INV_X1 U3391 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3611) );
  OR2_X1 U3392 ( .A1(n2537), .A2(n3611), .ZN(n2624) );
  NAND4_X1 U3393 ( .A1(n2627), .A2(n2626), .A3(n2625), .A4(n2624), .ZN(n3708)
         );
  INV_X1 U3394 ( .A(n2628), .ZN(n2630) );
  NOR2_X1 U3395 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2629)
         );
  NAND2_X1 U3396 ( .A1(n2630), .A2(n2629), .ZN(n2632) );
  NAND2_X1 U3397 ( .A1(n2632), .A2(IR_REG_31__SCAN_IN), .ZN(n2631) );
  MUX2_X1 U3398 ( .A(IR_REG_31__SCAN_IN), .B(n2631), .S(IR_REG_9__SCAN_IN), 
        .Z(n2633) );
  MUX2_X1 U3399 ( .A(n4954), .B(DATAI_9_), .S(n4056), .Z(n3703) );
  AND2_X1 U3400 ( .A1(n3708), .A2(n3703), .ZN(n2634) );
  NAND2_X1 U3401 ( .A1(n2813), .A2(REG2_REG_10__SCAN_IN), .ZN(n2641) );
  INV_X1 U3402 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4765) );
  OR2_X1 U3403 ( .A1(n3330), .A2(n4765), .ZN(n2640) );
  INV_X1 U3404 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4763) );
  OR2_X1 U3405 ( .A1(n2748), .A2(n4763), .ZN(n2639) );
  NAND2_X1 U3406 ( .A1(n2636), .A2(n2635), .ZN(n2637) );
  NAND2_X1 U3407 ( .A1(n2646), .A2(n2637), .ZN(n3728) );
  OR2_X1 U3408 ( .A1(n2812), .A2(n3728), .ZN(n2638) );
  NAND4_X1 U3409 ( .A1(n2641), .A2(n2640), .A3(n2639), .A4(n2638), .ZN(n3693)
         );
  NAND2_X1 U3410 ( .A1(n2643), .A2(IR_REG_31__SCAN_IN), .ZN(n2642) );
  MUX2_X1 U3411 ( .A(IR_REG_31__SCAN_IN), .B(n2642), .S(IR_REG_10__SCAN_IN), 
        .Z(n2644) );
  NAND2_X1 U3412 ( .A1(n2644), .A2(n2652), .ZN(n3675) );
  MUX2_X1 U3413 ( .A(n3239), .B(DATAI_10_), .S(n4056), .Z(n3725) );
  NAND2_X1 U3414 ( .A1(n2920), .A2(REG0_REG_11__SCAN_IN), .ZN(n2651) );
  INV_X1 U3415 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3747) );
  OR2_X1 U3416 ( .A1(n2748), .A2(n3747), .ZN(n2650) );
  NAND2_X1 U3417 ( .A1(n2646), .A2(n2645), .ZN(n2647) );
  NAND2_X1 U3418 ( .A1(n2668), .A2(n2647), .ZN(n4002) );
  OR2_X1 U3419 ( .A1(n2812), .A2(n4002), .ZN(n2649) );
  INV_X1 U3420 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3687) );
  OR2_X1 U3421 ( .A1(n2537), .A2(n3687), .ZN(n2648) );
  NAND2_X1 U3422 ( .A1(n2652), .A2(IR_REG_31__SCAN_IN), .ZN(n2655) );
  INV_X1 U3423 ( .A(n2655), .ZN(n2653) );
  NAND2_X1 U3424 ( .A1(n2653), .A2(IR_REG_11__SCAN_IN), .ZN(n2656) );
  INV_X1 U3425 ( .A(IR_REG_11__SCAN_IN), .ZN(n2654) );
  NAND2_X1 U3426 ( .A1(n2655), .A2(n2654), .ZN(n2662) );
  MUX2_X1 U3427 ( .A(n4953), .B(DATAI_11_), .S(n4056), .Z(n3999) );
  NAND2_X1 U3428 ( .A1(n3722), .A2(n3999), .ZN(n4154) );
  NAND2_X1 U3429 ( .A1(n4591), .A2(n3689), .ZN(n4150) );
  XNOR2_X1 U3430 ( .A(n2668), .B(REG3_REG_12__SCAN_IN), .ZN(n3925) );
  NAND2_X1 U3431 ( .A1(n2830), .A2(n3925), .ZN(n2661) );
  INV_X1 U3432 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4599) );
  OR2_X1 U3433 ( .A1(n2748), .A2(n4599), .ZN(n2660) );
  INV_X1 U3434 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4943) );
  OR2_X1 U3435 ( .A1(n3330), .A2(n4943), .ZN(n2659) );
  INV_X1 U3436 ( .A(REG2_REG_12__SCAN_IN), .ZN(n2657) );
  OR2_X1 U3437 ( .A1(n3334), .A2(n2657), .ZN(n2658) );
  NAND4_X1 U3438 ( .A1(n2661), .A2(n2660), .A3(n2659), .A4(n2658), .ZN(n4204)
         );
  NAND2_X1 U3439 ( .A1(n2662), .A2(IR_REG_31__SCAN_IN), .ZN(n2663) );
  XNOR2_X1 U3440 ( .A(n2663), .B(IR_REG_12__SCAN_IN), .ZN(n4951) );
  MUX2_X1 U3441 ( .A(n4951), .B(DATAI_12_), .S(n4056), .Z(n3756) );
  NAND2_X1 U3442 ( .A1(n4204), .A2(n3756), .ZN(n2664) );
  NAND2_X1 U3443 ( .A1(n3752), .A2(n2664), .ZN(n2666) );
  INV_X1 U3444 ( .A(n4204), .ZN(n3997) );
  NAND2_X1 U3445 ( .A1(n3997), .A2(n4594), .ZN(n2665) );
  NAND2_X1 U3446 ( .A1(n2666), .A2(n2665), .ZN(n3774) );
  INV_X1 U3447 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2667) );
  INV_X1 U3448 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4758) );
  OAI21_X1 U3449 ( .B1(n2668), .B2(n2667), .A(n4758), .ZN(n2669) );
  AND2_X1 U3450 ( .A1(n2680), .A2(n2669), .ZN(n3977) );
  NAND2_X1 U3451 ( .A1(n2830), .A2(n3977), .ZN(n2674) );
  INV_X1 U3452 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4939) );
  OR2_X1 U3453 ( .A1(n3330), .A2(n4939), .ZN(n2673) );
  INV_X1 U3454 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4586) );
  OR2_X1 U3455 ( .A1(n2748), .A2(n4586), .ZN(n2672) );
  INV_X1 U3456 ( .A(REG2_REG_13__SCAN_IN), .ZN(n2670) );
  OR2_X1 U3457 ( .A1(n3334), .A2(n2670), .ZN(n2671) );
  NAND4_X1 U34580 ( .A1(n2674), .A2(n2673), .A3(n2672), .A4(n2671), .ZN(n4588)
         );
  OR2_X1 U34590 ( .A1(n2823), .A2(n2293), .ZN(n2675) );
  XNOR2_X1 U3460 ( .A(n2675), .B(IR_REG_13__SCAN_IN), .ZN(n3247) );
  MUX2_X1 U3461 ( .A(n3247), .B(DATAI_13_), .S(n4056), .Z(n3976) );
  NOR2_X1 U3462 ( .A1(n4588), .A2(n3976), .ZN(n2676) );
  INV_X1 U3463 ( .A(REG0_REG_14__SCAN_IN), .ZN(n2677) );
  OR2_X1 U3464 ( .A1(n3330), .A2(n2677), .ZN(n2679) );
  INV_X1 U3465 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4760) );
  OR2_X1 U3466 ( .A1(n2748), .A2(n4760), .ZN(n2678) );
  AND2_X1 U34670 ( .A1(n2679), .A2(n2678), .ZN(n2684) );
  INV_X1 U3468 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4837) );
  NAND2_X1 U34690 ( .A1(n2680), .A2(n4837), .ZN(n2681) );
  NAND2_X1 U3470 ( .A1(n2686), .A2(n2681), .ZN(n3731) );
  OR2_X1 U34710 ( .A1(n3731), .A2(n2812), .ZN(n2683) );
  NAND2_X1 U3472 ( .A1(n2813), .A2(REG2_REG_14__SCAN_IN), .ZN(n2682) );
  NAND2_X1 U34730 ( .A1(n2691), .A2(IR_REG_31__SCAN_IN), .ZN(n2685) );
  XNOR2_X1 U3474 ( .A(n2685), .B(IR_REG_14__SCAN_IN), .ZN(n3273) );
  MUX2_X1 U34750 ( .A(n3273), .B(DATAI_14_), .S(n4056), .Z(n4571) );
  NAND2_X1 U3476 ( .A1(n4562), .A2(n4571), .ZN(n4043) );
  INV_X1 U34770 ( .A(n4562), .ZN(n4203) );
  INV_X1 U3478 ( .A(n4571), .ZN(n3880) );
  NAND2_X1 U34790 ( .A1(n4203), .A2(n3880), .ZN(n4044) );
  NAND2_X1 U3480 ( .A1(n4043), .A2(n4044), .ZN(n4100) );
  NAND2_X1 U34810 ( .A1(n2686), .A2(n4761), .ZN(n2687) );
  AND2_X1 U3482 ( .A1(n2695), .A2(n2687), .ZN(n4037) );
  NAND2_X1 U34830 ( .A1(n4037), .A2(n2830), .ZN(n2690) );
  AOI22_X1 U3484 ( .A1(n3329), .A2(REG1_REG_15__SCAN_IN), .B1(n2920), .B2(
        REG0_REG_15__SCAN_IN), .ZN(n2689) );
  INV_X1 U34850 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3790) );
  OR2_X1 U3486 ( .A1(n3334), .A2(n3790), .ZN(n2688) );
  INV_X1 U34870 ( .A(DATAI_15_), .ZN(n5056) );
  MUX2_X1 U3488 ( .A(n5057), .B(n5056), .S(n4056), .Z(n4560) );
  NAND2_X1 U34890 ( .A1(n3793), .A2(n2693), .ZN(n2694) );
  NAND2_X1 U3490 ( .A1(n2694), .A2(n2165), .ZN(n4447) );
  INV_X1 U34910 ( .A(n4447), .ZN(n2705) );
  INV_X1 U3492 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4691) );
  NAND2_X1 U34930 ( .A1(n2695), .A2(n4691), .ZN(n2696) );
  NAND2_X1 U3494 ( .A1(n2697), .A2(n2696), .ZN(n4452) );
  OR2_X1 U34950 ( .A1(n4452), .A2(n2812), .ZN(n2700) );
  AOI22_X1 U3496 ( .A1(n3329), .A2(REG1_REG_16__SCAN_IN), .B1(n2920), .B2(
        REG0_REG_16__SCAN_IN), .ZN(n2699) );
  NAND2_X1 U34970 ( .A1(n2813), .A2(REG2_REG_16__SCAN_IN), .ZN(n2698) );
  INV_X1 U3498 ( .A(IR_REG_15__SCAN_IN), .ZN(n2701) );
  NAND2_X1 U34990 ( .A1(n2702), .A2(n2701), .ZN(n2703) );
  NAND2_X1 U3500 ( .A1(n2703), .A2(IR_REG_31__SCAN_IN), .ZN(n2704) );
  XNOR2_X1 U35010 ( .A(n2704), .B(IR_REG_16__SCAN_IN), .ZN(n5054) );
  MUX2_X1 U3502 ( .A(n5054), .B(DATAI_16_), .S(n4056), .Z(n4455) );
  NAND2_X1 U35030 ( .A1(n4435), .A2(n4455), .ZN(n4166) );
  NAND2_X1 U3504 ( .A1(n4564), .A2(n4550), .ZN(n4162) );
  NAND2_X1 U35050 ( .A1(n2705), .A2(n4081), .ZN(n4445) );
  AND2_X2 U35060 ( .A1(n4445), .A2(n2706), .ZN(n4427) );
  INV_X1 U35070 ( .A(n2709), .ZN(n2727) );
  INV_X1 U35080 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4784) );
  NAND2_X1 U35090 ( .A1(n2727), .A2(n4784), .ZN(n2710) );
  NAND2_X1 U35100 ( .A1(n2735), .A2(n2710), .ZN(n3894) );
  OR2_X1 U35110 ( .A1(n3894), .A2(n2812), .ZN(n2716) );
  INV_X1 U35120 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2713) );
  NAND2_X1 U35130 ( .A1(n2920), .A2(REG0_REG_19__SCAN_IN), .ZN(n2712) );
  INV_X1 U35140 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4536) );
  OR2_X1 U35150 ( .A1(n2748), .A2(n4536), .ZN(n2711) );
  OAI211_X1 U35160 ( .C1(n2713), .C2(n3334), .A(n2712), .B(n2711), .ZN(n2714)
         );
  INV_X1 U35170 ( .A(n2714), .ZN(n2715) );
  NOR2_X1 U35180 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2719) );
  NAND2_X1 U35190 ( .A1(n2823), .A2(n2463), .ZN(n2720) );
  NAND2_X1 U35200 ( .A1(n2722), .A2(n2721), .ZN(n2819) );
  INV_X1 U35210 ( .A(DATAI_19_), .ZN(n2724) );
  MUX2_X1 U35220 ( .A(n4190), .B(n2724), .S(n4056), .Z(n4399) );
  NAND2_X1 U35230 ( .A1(n4417), .A2(n4399), .ZN(n4364) );
  INV_X1 U35240 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4658) );
  NAND2_X1 U35250 ( .A1(n2725), .A2(n4658), .ZN(n2726) );
  NAND2_X1 U35260 ( .A1(n4409), .A2(n2830), .ZN(n2732) );
  INV_X1 U35270 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4827) );
  NAND2_X1 U35280 ( .A1(n2920), .A2(REG0_REG_18__SCAN_IN), .ZN(n2729) );
  NAND2_X1 U35290 ( .A1(n2813), .A2(REG2_REG_18__SCAN_IN), .ZN(n2728) );
  OAI211_X1 U35300 ( .C1(n2748), .C2(n4827), .A(n2729), .B(n2728), .ZN(n2730)
         );
  INV_X1 U35310 ( .A(n2730), .ZN(n2731) );
  OAI21_X1 U35320 ( .B1(n2733), .B2(IR_REG_17__SCAN_IN), .A(IR_REG_31__SCAN_IN), .ZN(n2734) );
  XNOR2_X1 U35330 ( .A(n2734), .B(IR_REG_18__SCAN_IN), .ZN(n3255) );
  MUX2_X1 U35340 ( .A(n5052), .B(n5051), .S(n4056), .Z(n4411) );
  NAND2_X1 U35350 ( .A1(n4543), .A2(n4411), .ZN(n4363) );
  NAND2_X1 U35360 ( .A1(n4364), .A2(n4363), .ZN(n2742) );
  OR2_X1 U35370 ( .A1(n4438), .A2(n4411), .ZN(n4390) );
  NAND2_X1 U35380 ( .A1(n4438), .A2(n4411), .ZN(n4388) );
  NAND2_X1 U35390 ( .A1(n4390), .A2(n4388), .ZN(n4413) );
  NAND2_X1 U35400 ( .A1(n4527), .A2(n2902), .ZN(n4366) );
  NAND2_X1 U35410 ( .A1(n2735), .A2(n4812), .ZN(n2736) );
  AND2_X1 U35420 ( .A1(n2744), .A2(n2736), .ZN(n4379) );
  NAND2_X1 U35430 ( .A1(n4379), .A2(n2830), .ZN(n2741) );
  INV_X1 U35440 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4783) );
  NAND2_X1 U35450 ( .A1(n2813), .A2(REG2_REG_20__SCAN_IN), .ZN(n2738) );
  NAND2_X1 U35460 ( .A1(n2920), .A2(REG0_REG_20__SCAN_IN), .ZN(n2737) );
  OAI211_X1 U35470 ( .C1(n2748), .C2(n4783), .A(n2738), .B(n2737), .ZN(n2739)
         );
  INV_X1 U35480 ( .A(n2739), .ZN(n2740) );
  NAND2_X1 U35490 ( .A1(n4517), .A2(n4526), .ZN(n4084) );
  OAI211_X1 U35500 ( .C1(n2742), .C2(n4413), .A(n4366), .B(n4084), .ZN(n2743)
         );
  INV_X1 U35510 ( .A(n4517), .ZN(n3912) );
  NAND2_X1 U35520 ( .A1(n3912), .A2(n4382), .ZN(n4085) );
  INV_X1 U35530 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3911) );
  NAND2_X1 U35540 ( .A1(n2744), .A2(n3911), .ZN(n2745) );
  NAND2_X1 U35550 ( .A1(n2753), .A2(n2745), .ZN(n4354) );
  INV_X1 U35560 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4523) );
  NAND2_X1 U35570 ( .A1(n2813), .A2(REG2_REG_21__SCAN_IN), .ZN(n2747) );
  OR2_X1 U35580 ( .A1(n3330), .A2(n4781), .ZN(n2746) );
  OAI211_X1 U35590 ( .C1(n2748), .C2(n4523), .A(n2747), .B(n2746), .ZN(n2749)
         );
  INV_X1 U35600 ( .A(n2749), .ZN(n2750) );
  NAND2_X1 U35610 ( .A1(n4378), .A2(n4516), .ZN(n2752) );
  OR2_X2 U35620 ( .A1(n2753), .A2(n4810), .ZN(n2762) );
  NAND2_X1 U35630 ( .A1(n2753), .A2(n4810), .ZN(n2754) );
  NAND2_X1 U35640 ( .A1(n2762), .A2(n2754), .ZN(n3983) );
  OR2_X1 U35650 ( .A1(n3983), .A2(n2812), .ZN(n2759) );
  INV_X1 U35660 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4909) );
  NAND2_X1 U35670 ( .A1(n2813), .A2(REG2_REG_22__SCAN_IN), .ZN(n2756) );
  NAND2_X1 U35680 ( .A1(n3329), .A2(REG1_REG_22__SCAN_IN), .ZN(n2755) );
  OAI211_X1 U35690 ( .C1(n3330), .C2(n4909), .A(n2756), .B(n2755), .ZN(n2757)
         );
  INV_X1 U35700 ( .A(n2757), .ZN(n2758) );
  NAND2_X1 U35710 ( .A1(n4520), .A2(n4334), .ZN(n4312) );
  INV_X1 U35720 ( .A(n4334), .ZN(n3984) );
  NAND2_X1 U35730 ( .A1(n4356), .A2(n3984), .ZN(n2857) );
  NAND2_X1 U35740 ( .A1(n4312), .A2(n2857), .ZN(n4340) );
  NAND2_X1 U35750 ( .A1(n2762), .A2(n2761), .ZN(n2763) );
  AND2_X1 U35760 ( .A1(n2772), .A2(n2763), .ZN(n4320) );
  NAND2_X1 U35770 ( .A1(n4320), .A2(n2830), .ZN(n2769) );
  INV_X1 U35780 ( .A(REG2_REG_23__SCAN_IN), .ZN(n2766) );
  NAND2_X1 U35790 ( .A1(n2920), .A2(REG0_REG_23__SCAN_IN), .ZN(n2765) );
  NAND2_X1 U35800 ( .A1(n3329), .A2(REG1_REG_23__SCAN_IN), .ZN(n2764) );
  OAI211_X1 U35810 ( .C1(n2766), .C2(n3334), .A(n2765), .B(n2764), .ZN(n2767)
         );
  INV_X1 U3582 ( .A(n2767), .ZN(n2768) );
  NAND2_X1 U3583 ( .A1(n2133), .A2(DATAI_23_), .ZN(n3090) );
  NAND2_X1 U3584 ( .A1(n4333), .A2(n3090), .ZN(n2771) );
  NOR2_X1 U3585 ( .A1(n4333), .A2(n3090), .ZN(n2770) );
  AOI21_X2 U3586 ( .B1(n4315), .B2(n2771), .A(n2770), .ZN(n4290) );
  INV_X1 U3587 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4813) );
  NAND2_X1 U3588 ( .A1(n2772), .A2(n4813), .ZN(n2773) );
  NAND2_X1 U3589 ( .A1(n4305), .A2(n2830), .ZN(n2779) );
  INV_X1 U3590 ( .A(REG2_REG_24__SCAN_IN), .ZN(n2776) );
  NAND2_X1 U3591 ( .A1(n3329), .A2(REG1_REG_24__SCAN_IN), .ZN(n2775) );
  NAND2_X1 U3592 ( .A1(n2920), .A2(REG0_REG_24__SCAN_IN), .ZN(n2774) );
  OAI211_X1 U3593 ( .C1(n2776), .C2(n3334), .A(n2775), .B(n2774), .ZN(n2777)
         );
  INV_X1 U3594 ( .A(n2777), .ZN(n2778) );
  NAND2_X1 U3595 ( .A1(n4494), .A2(n3957), .ZN(n2780) );
  NAND2_X1 U3596 ( .A1(n4290), .A2(n2780), .ZN(n2782) );
  INV_X1 U3597 ( .A(n4494), .ZN(n4314) );
  NAND2_X1 U3598 ( .A1(n4314), .A2(n4303), .ZN(n2781) );
  NAND2_X1 U3599 ( .A1(n2782), .A2(n2781), .ZN(n4278) );
  INV_X1 U3600 ( .A(n4278), .ZN(n2792) );
  INV_X1 U3601 ( .A(REG3_REG_25__SCAN_IN), .ZN(n2784) );
  NAND2_X1 U3602 ( .A1(n2785), .A2(n2784), .ZN(n2786) );
  NAND2_X1 U3603 ( .A1(n2793), .A2(n2786), .ZN(n4282) );
  INV_X1 U3604 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4281) );
  NAND2_X1 U3605 ( .A1(n2920), .A2(REG0_REG_25__SCAN_IN), .ZN(n2788) );
  NAND2_X1 U3606 ( .A1(n3329), .A2(REG1_REG_25__SCAN_IN), .ZN(n2787) );
  OAI211_X1 U3607 ( .C1(n4281), .C2(n3334), .A(n2788), .B(n2787), .ZN(n2789)
         );
  INV_X1 U3608 ( .A(n2789), .ZN(n2790) );
  OR2_X2 U3609 ( .A1(n2793), .A2(n4829), .ZN(n2810) );
  NAND2_X1 U3610 ( .A1(n2793), .A2(n4829), .ZN(n2794) );
  NAND2_X1 U3611 ( .A1(n4020), .A2(n2830), .ZN(n2799) );
  INV_X1 U3612 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4893) );
  NAND2_X1 U3613 ( .A1(n2813), .A2(REG2_REG_26__SCAN_IN), .ZN(n2796) );
  NAND2_X1 U3614 ( .A1(n3329), .A2(REG1_REG_26__SCAN_IN), .ZN(n2795) );
  OAI211_X1 U3615 ( .C1(n3330), .C2(n4893), .A(n2796), .B(n2795), .ZN(n2797)
         );
  INV_X1 U3616 ( .A(n2797), .ZN(n2798) );
  NAND2_X1 U3617 ( .A1(n4483), .A2(n4019), .ZN(n3805) );
  NOR2_X1 U3618 ( .A1(n4483), .A2(n4019), .ZN(n3806) );
  XNOR2_X1 U3619 ( .A(n2810), .B(REG3_REG_27__SCAN_IN), .ZN(n4266) );
  NAND2_X1 U3620 ( .A1(n4266), .A2(n2830), .ZN(n2804) );
  INV_X1 U3621 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4888) );
  NAND2_X1 U3622 ( .A1(n2813), .A2(REG2_REG_27__SCAN_IN), .ZN(n2801) );
  NAND2_X1 U3623 ( .A1(n3329), .A2(REG1_REG_27__SCAN_IN), .ZN(n2800) );
  OAI211_X1 U3624 ( .C1(n3330), .C2(n4888), .A(n2801), .B(n2800), .ZN(n2802)
         );
  INV_X1 U3625 ( .A(n2802), .ZN(n2803) );
  AND2_X2 U3626 ( .A1(n2804), .A2(n2803), .ZN(n3812) );
  NAND2_X1 U3627 ( .A1(n2133), .A2(DATAI_27_), .ZN(n3125) );
  NAND2_X1 U3628 ( .A1(n3812), .A2(n3125), .ZN(n2805) );
  NAND2_X1 U3629 ( .A1(n4200), .A2(n4482), .ZN(n2806) );
  INV_X1 U3630 ( .A(n2810), .ZN(n2808) );
  AND2_X1 U3631 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_28__SCAN_IN), .ZN(
        n2807) );
  NAND2_X1 U3632 ( .A1(n2808), .A2(n2807), .ZN(n2916) );
  INV_X1 U3633 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4652) );
  INV_X1 U3634 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2809) );
  OAI21_X1 U3635 ( .B1(n2810), .B2(n4652), .A(n2809), .ZN(n2811) );
  NAND2_X1 U3636 ( .A1(n2916), .A2(n2811), .ZN(n3842) );
  OR2_X1 U3637 ( .A1(n3842), .A2(n2812), .ZN(n2818) );
  INV_X1 U3638 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4654) );
  NAND2_X1 U3639 ( .A1(n2813), .A2(REG2_REG_28__SCAN_IN), .ZN(n2815) );
  OR2_X1 U3640 ( .A1(n3330), .A2(n3266), .ZN(n2814) );
  OAI211_X1 U3641 ( .C1(n2748), .C2(n4654), .A(n2815), .B(n2814), .ZN(n2816)
         );
  INV_X1 U3642 ( .A(n2816), .ZN(n2817) );
  AND2_X1 U3643 ( .A1(n2133), .A2(DATAI_28_), .ZN(n3839) );
  NAND2_X1 U3644 ( .A1(n4486), .A2(n3839), .ZN(n2918) );
  NAND2_X1 U3645 ( .A1(n4271), .A2(n3128), .ZN(n4062) );
  NAND2_X1 U3646 ( .A1(n2918), .A2(n4062), .ZN(n2933) );
  XNOR2_X1 U3647 ( .A(n2934), .B(n2933), .ZN(n3837) );
  XNOR2_X2 U3648 ( .A(n2821), .B(n2820), .ZN(n2861) );
  AND2_X2 U3649 ( .A1(n2823), .A2(n2822), .ZN(n2826) );
  XNOR2_X1 U3650 ( .A(n2947), .B(n2946), .ZN(n2828) );
  NAND2_X1 U3651 ( .A1(n2828), .A2(n4190), .ZN(n3323) );
  NAND2_X1 U3652 ( .A1(n2861), .A2(n4950), .ZN(n5026) );
  NAND2_X1 U3653 ( .A1(n2395), .A2(IR_REG_31__SCAN_IN), .ZN(n2829) );
  XNOR2_X1 U3654 ( .A(n2829), .B(IR_REG_28__SCAN_IN), .ZN(n4959) );
  NAND2_X1 U3655 ( .A1(n3213), .A2(n4959), .ZN(n4561) );
  INV_X1 U3656 ( .A(n2916), .ZN(n2831) );
  NAND2_X1 U3657 ( .A1(n2831), .A2(n2830), .ZN(n2837) );
  INV_X1 U3658 ( .A(REG2_REG_29__SCAN_IN), .ZN(n2937) );
  NAND2_X1 U3659 ( .A1(n3329), .A2(REG1_REG_29__SCAN_IN), .ZN(n2834) );
  INV_X1 U3660 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2832) );
  OR2_X1 U3661 ( .A1(n3330), .A2(n2832), .ZN(n2833) );
  OAI211_X1 U3662 ( .C1(n2937), .C2(n3334), .A(n2834), .B(n2833), .ZN(n2835)
         );
  INV_X1 U3663 ( .A(n2835), .ZN(n2836) );
  INV_X1 U3664 ( .A(n4199), .ZN(n2838) );
  NOR2_X2 U3665 ( .A1(n3310), .A2(n2861), .ZN(n4570) );
  OAI22_X1 U3666 ( .A1(n2838), .A2(n4573), .B1(n4593), .B2(n3128), .ZN(n2839)
         );
  AOI21_X1 U3667 ( .B1(n4590), .B2(n4200), .A(n2839), .ZN(n2864) );
  INV_X1 U3668 ( .A(n4099), .ZN(n2840) );
  NAND2_X1 U3669 ( .A1(n4118), .A2(n2840), .ZN(n3378) );
  NAND2_X1 U3670 ( .A1(n3378), .A2(n4119), .ZN(n2842) );
  INV_X1 U3671 ( .A(n4091), .ZN(n2841) );
  NAND2_X1 U3672 ( .A1(n2842), .A2(n2841), .ZN(n3380) );
  NAND2_X1 U3673 ( .A1(n3380), .A2(n4120), .ZN(n3402) );
  OR2_X1 U3674 ( .A1(n4470), .A2(n3553), .ZN(n4125) );
  NAND2_X1 U3675 ( .A1(n4470), .A2(n3553), .ZN(n4122) );
  INV_X1 U3676 ( .A(n4126), .ZN(n2843) );
  AND2_X1 U3677 ( .A1(n4207), .A2(n3497), .ZN(n4129) );
  OR2_X1 U3678 ( .A1(n4207), .A2(n3497), .ZN(n4143) );
  NAND2_X1 U3679 ( .A1(n3582), .A2(n2303), .ZN(n4128) );
  OR2_X1 U3680 ( .A1(n3582), .A2(n2303), .ZN(n4130) );
  INV_X1 U3681 ( .A(n2845), .ZN(n2846) );
  OR2_X1 U3682 ( .A1(n4205), .A2(n3637), .ZN(n4137) );
  NAND2_X1 U3683 ( .A1(n4205), .A2(n3637), .ZN(n4135) );
  AND2_X1 U3684 ( .A1(n3708), .A2(n3612), .ZN(n4144) );
  INV_X1 U3685 ( .A(n4144), .ZN(n2847) );
  OR2_X1 U3686 ( .A1(n3708), .A2(n3612), .ZN(n4138) );
  INV_X1 U3687 ( .A(n3725), .ZN(n3644) );
  NAND2_X1 U3688 ( .A1(n3693), .A2(n3644), .ZN(n4149) );
  OR2_X1 U3689 ( .A1(n3693), .A2(n3644), .ZN(n4146) );
  NAND2_X1 U3690 ( .A1(n2848), .A2(n4146), .ZN(n3681) );
  NAND2_X1 U3691 ( .A1(n3681), .A2(n4150), .ZN(n2849) );
  NAND2_X1 U3692 ( .A1(n4204), .A2(n4594), .ZN(n3767) );
  NAND2_X1 U3693 ( .A1(n4588), .A2(n3775), .ZN(n3765) );
  NOR2_X1 U3694 ( .A1(n4204), .A2(n4594), .ZN(n3768) );
  OR2_X1 U3695 ( .A1(n4588), .A2(n3775), .ZN(n3766) );
  INV_X1 U3696 ( .A(n3766), .ZN(n2850) );
  AOI21_X1 U3697 ( .B1(n4156), .B2(n3768), .A(n2850), .ZN(n4160) );
  INV_X1 U3698 ( .A(n4100), .ZN(n3736) );
  OR2_X1 U3699 ( .A1(n4454), .A2(n4560), .ZN(n4046) );
  NAND2_X1 U3700 ( .A1(n4454), .A2(n4560), .ZN(n4045) );
  NAND2_X1 U3701 ( .A1(n4046), .A2(n4045), .ZN(n4080) );
  NAND2_X1 U3702 ( .A1(n4444), .A2(n4448), .ZN(n4443) );
  NAND2_X1 U3703 ( .A1(n4527), .A2(n4399), .ZN(n2852) );
  AND2_X1 U3704 ( .A1(n2852), .A2(n4388), .ZN(n2855) );
  INV_X1 U3705 ( .A(n2855), .ZN(n4373) );
  AND2_X1 U3706 ( .A1(n4555), .A2(n4432), .ZN(n4369) );
  OR2_X1 U3707 ( .A1(n4373), .A2(n4369), .ZN(n4165) );
  NOR2_X1 U3708 ( .A1(n4555), .A2(n4432), .ZN(n4370) );
  AOI22_X1 U3709 ( .A1(n2855), .A2(n4370), .B1(n3912), .B2(n4526), .ZN(n2856)
         );
  INV_X1 U3710 ( .A(n4390), .ZN(n2854) );
  NOR2_X1 U3711 ( .A1(n4527), .A2(n4399), .ZN(n2853) );
  AOI21_X1 U3712 ( .B1(n2855), .B2(n2854), .A(n2853), .ZN(n4372) );
  AND2_X1 U3713 ( .A1(n2856), .A2(n4372), .ZN(n4049) );
  NAND2_X1 U3714 ( .A1(n4517), .A2(n4382), .ZN(n4169) );
  NAND2_X1 U3715 ( .A1(n4530), .A2(n4516), .ZN(n4311) );
  AND2_X1 U3716 ( .A1(n4312), .A2(n4311), .ZN(n4172) );
  NAND2_X1 U3717 ( .A1(n4201), .A2(n3090), .ZN(n4079) );
  NAND2_X1 U3718 ( .A1(n4079), .A2(n2857), .ZN(n4054) );
  AND2_X1 U3719 ( .A1(n4378), .A2(n4350), .ZN(n4310) );
  AND2_X1 U3720 ( .A1(n4312), .A2(n4310), .ZN(n4051) );
  NOR2_X1 U3721 ( .A1(n4054), .A2(n4051), .ZN(n2858) );
  OR2_X1 U3722 ( .A1(n4494), .A2(n4303), .ZN(n4078) );
  OR2_X1 U3723 ( .A1(n4201), .A2(n3090), .ZN(n4291) );
  NAND2_X1 U3724 ( .A1(n4494), .A2(n4303), .ZN(n4077) );
  AND2_X1 U3725 ( .A1(n4298), .A2(n4285), .ZN(n4075) );
  NAND2_X1 U3726 ( .A1(n4497), .A2(n4019), .ZN(n2859) );
  INV_X1 U3727 ( .A(n4298), .ZN(n4023) );
  NAND2_X1 U3728 ( .A1(n4023), .A2(n4493), .ZN(n4076) );
  INV_X1 U3729 ( .A(n4019), .ZN(n3816) );
  AND2_X1 U3730 ( .A1(n4483), .A2(n3816), .ZN(n4063) );
  NAND2_X1 U3731 ( .A1(n3812), .A2(n4482), .ZN(n2917) );
  NAND2_X1 U3732 ( .A1(n4200), .A2(n3125), .ZN(n4179) );
  INV_X1 U3733 ( .A(n2933), .ZN(n4111) );
  XNOR2_X1 U3734 ( .A(n2860), .B(n4111), .ZN(n2863) );
  NAND2_X1 U3735 ( .A1(n4949), .A2(n4948), .ZN(n4188) );
  NAND2_X1 U3736 ( .A1(n2946), .A2(n4950), .ZN(n2862) );
  NAND2_X1 U3737 ( .A1(n2865), .A2(IR_REG_31__SCAN_IN), .ZN(n2866) );
  MUX2_X1 U3738 ( .A(IR_REG_31__SCAN_IN), .B(n2866), .S(IR_REG_25__SCAN_IN), 
        .Z(n2868) );
  NAND2_X1 U3739 ( .A1(n2868), .A2(n2867), .ZN(n3279) );
  NAND2_X1 U3740 ( .A1(n3279), .A2(B_REG_SCAN_IN), .ZN(n2871) );
  MUX2_X1 U3741 ( .A(n2871), .B(B_REG_SCAN_IN), .S(n2879), .Z(n2877) );
  NAND2_X1 U3742 ( .A1(n2867), .A2(IR_REG_31__SCAN_IN), .ZN(n2873) );
  NAND2_X1 U3743 ( .A1(n2878), .A2(n3279), .ZN(n3290) );
  NAND2_X1 U3744 ( .A1(n3131), .A2(n3290), .ZN(n2898) );
  NOR2_X1 U3745 ( .A1(n2878), .A2(n3279), .ZN(n2880) );
  NAND2_X1 U3746 ( .A1(n2880), .A2(n2879), .ZN(n2943) );
  NAND2_X1 U3747 ( .A1(n2861), .A2(n4190), .ZN(n2885) );
  NAND2_X1 U3748 ( .A1(n3213), .A2(n2885), .ZN(n3147) );
  NAND2_X1 U3749 ( .A1(n2913), .A2(n3147), .ZN(n2886) );
  NOR2_X1 U3750 ( .A1(n3211), .A2(n2886), .ZN(n2897) );
  INV_X1 U3751 ( .A(D_REG_31__SCAN_IN), .ZN(n5034) );
  INV_X1 U3752 ( .A(D_REG_29__SCAN_IN), .ZN(n5036) );
  INV_X1 U3753 ( .A(D_REG_9__SCAN_IN), .ZN(n5046) );
  INV_X1 U3754 ( .A(D_REG_11__SCAN_IN), .ZN(n5045) );
  NAND4_X1 U3755 ( .A1(n5034), .A2(n5036), .A3(n5046), .A4(n5045), .ZN(n2887)
         );
  NOR4_X1 U3756 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(n2887), .ZN(n4650) );
  NOR4_X1 U3757 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2889) );
  NOR3_X1 U3758 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .ZN(n2888) );
  NAND3_X1 U3759 ( .A1(n4650), .A2(n2889), .A3(n2888), .ZN(n2895) );
  NOR4_X1 U3760 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2893) );
  NOR4_X1 U3761 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_7__SCAN_IN), .ZN(n2892) );
  NOR4_X1 U3762 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n2891) );
  NOR4_X1 U3763 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2890) );
  NAND4_X1 U3764 ( .A1(n2893), .A2(n2892), .A3(n2891), .A4(n2890), .ZN(n2894)
         );
  NOR2_X1 U3765 ( .A1(n2895), .A2(n2894), .ZN(n2896) );
  NAND2_X1 U3766 ( .A1(n3318), .A2(n3311), .ZN(n3386) );
  NAND2_X1 U3767 ( .A1(n3540), .A2(n3612), .ZN(n3609) );
  NAND2_X1 U3768 ( .A1(n4264), .A2(n3128), .ZN(n2906) );
  NAND2_X1 U3769 ( .A1(n5079), .A2(REG1_REG_28__SCAN_IN), .ZN(n2903) );
  NAND2_X1 U3770 ( .A1(n2133), .A2(DATAI_29_), .ZN(n2925) );
  INV_X1 U3771 ( .A(D_REG_1__SCAN_IN), .ZN(n2911) );
  OAI21_X1 U3772 ( .B1(n3211), .B2(n2911), .A(n5048), .ZN(n2912) );
  NAND4_X1 U3773 ( .A1(n3173), .A2(n3133), .A3(n3147), .A4(n2912), .ZN(n2914)
         );
  AND2_X1 U3774 ( .A1(n2941), .A2(n4190), .ZN(n2915) );
  OAI22_X1 U3775 ( .A1(n3178), .A2(n4458), .B1(n2916), .B2(n4451), .ZN(n2931)
         );
  NAND2_X1 U3776 ( .A1(n2918), .A2(n2917), .ZN(n4066) );
  OAI21_X1 U3777 ( .B1(n4261), .B2(n4066), .A(n4062), .ZN(n2919) );
  OR2_X1 U3778 ( .A1(n4199), .A2(n2925), .ZN(n4058) );
  NAND2_X1 U3779 ( .A1(n4199), .A2(n2925), .ZN(n4061) );
  NAND2_X1 U3780 ( .A1(n4058), .A2(n4061), .ZN(n4074) );
  XNOR2_X1 U3781 ( .A(n2919), .B(n4074), .ZN(n2929) );
  INV_X1 U3782 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4819) );
  INV_X1 U3783 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4656) );
  OR2_X1 U3784 ( .A1(n2748), .A2(n4656), .ZN(n2922) );
  NAND2_X1 U3785 ( .A1(n2920), .A2(REG0_REG_30__SCAN_IN), .ZN(n2921) );
  OAI211_X1 U3786 ( .C1(n3334), .C2(n4819), .A(n2922), .B(n2921), .ZN(n4198)
         );
  XNOR2_X1 U3787 ( .A(n2923), .B(IR_REG_27__SCAN_IN), .ZN(n4966) );
  NAND2_X1 U3788 ( .A1(n4966), .A2(B_REG_SCAN_IN), .ZN(n2924) );
  AND2_X1 U3789 ( .A1(n4589), .A2(n2924), .ZN(n4245) );
  INV_X1 U3790 ( .A(n2925), .ZN(n2926) );
  AOI22_X1 U3791 ( .A1(n4198), .A2(n4245), .B1(n2926), .B2(n4570), .ZN(n2927)
         );
  OAI21_X1 U3792 ( .B1(n4486), .B2(n4561), .A(n2927), .ZN(n2928) );
  INV_X1 U3793 ( .A(n3167), .ZN(n2930) );
  NOR2_X1 U3794 ( .A1(n4486), .A2(n3128), .ZN(n2932) );
  XNOR2_X1 U3795 ( .A(n2935), .B(n4074), .ZN(n3166) );
  OR2_X1 U3796 ( .A1(n2947), .A2(n4190), .ZN(n3441) );
  NAND2_X1 U3797 ( .A1(n3323), .A2(n3441), .ZN(n2936) );
  INV_X2 U3798 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  AND2_X4 U3799 ( .A1(n2943), .A2(n2947), .ZN(n3112) );
  INV_X1 U3800 ( .A(n2947), .ZN(n2942) );
  AND2_X2 U3801 ( .A1(n2943), .A2(n2942), .ZN(n3012) );
  AOI22_X1 U3802 ( .A1(n3116), .A2(n4207), .B1(n3534), .B2(n3035), .ZN(n2988)
         );
  INV_X1 U3803 ( .A(n2988), .ZN(n2990) );
  NAND2_X1 U3804 ( .A1(n4207), .A2(n3029), .ZN(n2945) );
  NAND2_X1 U3805 ( .A1(n3534), .A2(n3112), .ZN(n2944) );
  NAND2_X1 U3806 ( .A1(n2945), .A2(n2944), .ZN(n2948) );
  NAND2_X1 U3807 ( .A1(n2946), .A2(n4190), .ZN(n3143) );
  XNOR2_X1 U3808 ( .A(n2948), .B(n3007), .ZN(n2989) );
  AOI22_X1 U3809 ( .A1(n3035), .A2(n2949), .B1(n3116), .B2(n3531), .ZN(n2985)
         );
  INV_X1 U3810 ( .A(n2985), .ZN(n2987) );
  NAND2_X1 U3811 ( .A1(n3531), .A2(n3029), .ZN(n2951) );
  OR2_X1 U3812 ( .A1(n2583), .A2(n2955), .ZN(n2950) );
  NAND2_X1 U3813 ( .A1(n2951), .A2(n2950), .ZN(n2952) );
  XNOR2_X1 U3814 ( .A(n2952), .B(n3007), .ZN(n2986) );
  NAND2_X1 U3815 ( .A1(n3116), .A2(n2135), .ZN(n2954) );
  OR2_X1 U3816 ( .A1(n3382), .A2(n2979), .ZN(n2953) );
  NAND2_X1 U3817 ( .A1(n2954), .A2(n2953), .ZN(n2959) );
  INV_X1 U3818 ( .A(n2959), .ZN(n2978) );
  NAND2_X1 U3819 ( .A1(n2135), .A2(n3029), .ZN(n2957) );
  INV_X1 U3820 ( .A(n2960), .ZN(n2977) );
  XNOR2_X1 U3821 ( .A(n2960), .B(n2959), .ZN(n3824) );
  NAND2_X1 U3822 ( .A1(n2972), .A2(n2963), .ZN(n2962) );
  NAND2_X1 U3823 ( .A1(n3832), .A2(n3012), .ZN(n2961) );
  NAND2_X1 U3824 ( .A1(n2962), .A2(n2961), .ZN(n3338) );
  NAND2_X1 U3825 ( .A1(n2963), .A2(n3012), .ZN(n2965) );
  NAND2_X1 U3826 ( .A1(n3832), .A2(n3112), .ZN(n2964) );
  NAND2_X1 U3827 ( .A1(n2965), .A2(n2964), .ZN(n3337) );
  NAND2_X1 U3828 ( .A1(n5060), .A2(REG1_REG_0__SCAN_IN), .ZN(n3180) );
  NOR2_X1 U3829 ( .A1(n2943), .A2(n3180), .ZN(n2966) );
  AOI21_X1 U3830 ( .B1(n3338), .B2(n3337), .A(n2966), .ZN(n3340) );
  NAND2_X1 U3831 ( .A1(n3340), .A2(n2967), .ZN(n3902) );
  NAND2_X1 U3832 ( .A1(n2968), .A2(n3112), .ZN(n2970) );
  NAND2_X1 U3833 ( .A1(n4465), .A2(n3012), .ZN(n2969) );
  NAND2_X1 U3834 ( .A1(n2970), .A2(n2969), .ZN(n2971) );
  AOI22_X1 U3835 ( .A1(n2968), .A2(n3012), .B1(n2972), .B2(n4465), .ZN(n2974)
         );
  XNOR2_X1 U3836 ( .A(n2973), .B(n2974), .ZN(n3901) );
  NAND2_X1 U3837 ( .A1(n3902), .A2(n3901), .ZN(n3903) );
  INV_X1 U3838 ( .A(n2974), .ZN(n2975) );
  NAND2_X1 U3839 ( .A1(n2973), .A2(n2975), .ZN(n2976) );
  NAND2_X1 U3840 ( .A1(n3903), .A2(n2976), .ZN(n3823) );
  NOR2_X2 U3841 ( .A1(n3824), .A2(n3823), .ZN(n3822) );
  AOI21_X1 U3842 ( .B1(n2978), .B2(n2977), .A(n3822), .ZN(n3477) );
  AOI22_X1 U3843 ( .A1(n3116), .A2(n4470), .B1(n3405), .B2(n3035), .ZN(n2983)
         );
  NAND2_X1 U3844 ( .A1(n4470), .A2(n3029), .ZN(n2981) );
  NAND2_X1 U3845 ( .A1(n3405), .A2(n3112), .ZN(n2980) );
  NAND2_X1 U3846 ( .A1(n2981), .A2(n2980), .ZN(n2982) );
  XNOR2_X1 U3847 ( .A(n2982), .B(n3007), .ZN(n2984) );
  XOR2_X1 U3848 ( .A(n2983), .B(n2984), .Z(n3478) );
  XOR2_X1 U3849 ( .A(n2986), .B(n2985), .Z(n3472) );
  XOR2_X1 U3850 ( .A(n2988), .B(n2989), .Z(n3529) );
  INV_X1 U3851 ( .A(n3582), .ZN(n3656) );
  OAI22_X1 U3852 ( .A1(n3656), .A2(n3126), .B1(n2303), .B2(n3088), .ZN(n3518)
         );
  INV_X1 U3853 ( .A(n3518), .ZN(n2993) );
  AOI22_X1 U3854 ( .A1(n3029), .A2(n3582), .B1(n3567), .B2(n3112), .ZN(n2991)
         );
  XOR2_X1 U3855 ( .A(n3007), .B(n2991), .Z(n3519) );
  INV_X1 U3856 ( .A(n3519), .ZN(n2992) );
  AOI21_X1 U3857 ( .B1(n3521), .B2(n2993), .A(n2992), .ZN(n2994) );
  INV_X1 U3858 ( .A(n2994), .ZN(n2995) );
  NAND2_X1 U3859 ( .A1(n4206), .A2(n3035), .ZN(n2997) );
  OR2_X1 U3860 ( .A1(n3577), .A2(n2955), .ZN(n2996) );
  NAND2_X1 U3861 ( .A1(n2997), .A2(n2996), .ZN(n2999) );
  XNOR2_X1 U3862 ( .A(n2999), .B(n2998), .ZN(n3002) );
  NAND2_X1 U3863 ( .A1(n3116), .A2(n4206), .ZN(n3001) );
  OR2_X1 U3864 ( .A1(n3577), .A2(n3088), .ZN(n3000) );
  NAND2_X1 U3865 ( .A1(n3001), .A2(n3000), .ZN(n3003) );
  XNOR2_X1 U3866 ( .A(n3002), .B(n3003), .ZN(n3654) );
  INV_X1 U3867 ( .A(n3002), .ZN(n3004) );
  NAND2_X1 U3868 ( .A1(n4205), .A2(n3035), .ZN(n3006) );
  NAND2_X1 U3869 ( .A1(n3009), .A2(n3112), .ZN(n3005) );
  NAND2_X1 U3870 ( .A1(n3006), .A2(n3005), .ZN(n3008) );
  XNOR2_X1 U3871 ( .A(n3008), .B(n2998), .ZN(n3011) );
  AOI22_X1 U3872 ( .A1(n3116), .A2(n4205), .B1(n3009), .B2(n3029), .ZN(n3010)
         );
  OR2_X1 U3873 ( .A1(n3011), .A2(n3010), .ZN(n3633) );
  NAND2_X1 U3874 ( .A1(n3011), .A2(n3010), .ZN(n3632) );
  NAND2_X1 U3875 ( .A1(n3708), .A2(n3012), .ZN(n3014) );
  NAND2_X1 U3876 ( .A1(n3703), .A2(n3112), .ZN(n3013) );
  NAND2_X1 U3877 ( .A1(n3014), .A2(n3013), .ZN(n3015) );
  XNOR2_X1 U3878 ( .A(n3015), .B(n3007), .ZN(n3016) );
  AOI22_X1 U3879 ( .A1(n3116), .A2(n3708), .B1(n3703), .B2(n3035), .ZN(n3017)
         );
  XNOR2_X1 U3880 ( .A(n3016), .B(n3017), .ZN(n3698) );
  INV_X1 U3881 ( .A(n3016), .ZN(n3018) );
  AOI22_X1 U3882 ( .A1(n3116), .A2(n3693), .B1(n3725), .B2(n3035), .ZN(n3020)
         );
  AOI22_X1 U3883 ( .A1(n3035), .A2(n3693), .B1(n3725), .B2(n3112), .ZN(n3019)
         );
  XNOR2_X1 U3884 ( .A(n3019), .B(n3007), .ZN(n3021) );
  XOR2_X1 U3885 ( .A(n3020), .B(n3021), .Z(n3718) );
  OAI22_X1 U3886 ( .A1(n3722), .A2(n3126), .B1(n3689), .B2(n3088), .ZN(n3991)
         );
  OAI22_X1 U3887 ( .A1(n3722), .A2(n3088), .B1(n3689), .B2(n2955), .ZN(n3023)
         );
  XNOR2_X1 U3888 ( .A(n3023), .B(n3007), .ZN(n3992) );
  NAND2_X1 U3889 ( .A1(n4204), .A2(n3035), .ZN(n3027) );
  NAND2_X1 U3890 ( .A1(n3756), .A2(n3112), .ZN(n3026) );
  NAND2_X1 U3891 ( .A1(n3027), .A2(n3026), .ZN(n3028) );
  XNOR2_X1 U3892 ( .A(n3028), .B(n2998), .ZN(n3031) );
  AOI22_X1 U3893 ( .A1(n3116), .A2(n4204), .B1(n3756), .B2(n3029), .ZN(n3030)
         );
  NOR2_X1 U3894 ( .A1(n3031), .A2(n3030), .ZN(n3919) );
  NAND2_X1 U3895 ( .A1(n3031), .A2(n3030), .ZN(n3918) );
  NAND2_X1 U3896 ( .A1(n4588), .A2(n3029), .ZN(n3033) );
  NAND2_X1 U3897 ( .A1(n3976), .A2(n3112), .ZN(n3032) );
  NAND2_X1 U3898 ( .A1(n3033), .A2(n3032), .ZN(n3034) );
  XNOR2_X1 U3899 ( .A(n3034), .B(n2998), .ZN(n3972) );
  NAND2_X1 U3900 ( .A1(n3116), .A2(n4588), .ZN(n3037) );
  NAND2_X1 U3901 ( .A1(n3976), .A2(n3035), .ZN(n3036) );
  OAI22_X1 U3902 ( .A1(n4562), .A2(n3088), .B1(n3880), .B2(n2955), .ZN(n3038)
         );
  XNOR2_X1 U3903 ( .A(n3038), .B(n3007), .ZN(n3042) );
  OAI22_X1 U3904 ( .A1(n4562), .A2(n3126), .B1(n3880), .B2(n3088), .ZN(n3041)
         );
  NAND2_X1 U3905 ( .A1(n3042), .A2(n3041), .ZN(n3876) );
  NAND3_X1 U3906 ( .A1(n3876), .A2(n3971), .A3(n3972), .ZN(n3043) );
  OR2_X1 U3907 ( .A1(n3042), .A2(n3041), .ZN(n3875) );
  OAI22_X1 U3908 ( .A1(n4574), .A2(n3126), .B1(n3088), .B2(n4560), .ZN(n4031)
         );
  OAI22_X1 U3909 ( .A1(n4574), .A2(n3088), .B1(n2955), .B2(n4560), .ZN(n3044)
         );
  XNOR2_X1 U3910 ( .A(n3044), .B(n3007), .ZN(n3929) );
  OAI22_X1 U3911 ( .A1(n4435), .A2(n3088), .B1(n2955), .B2(n4550), .ZN(n3045)
         );
  XNOR2_X1 U3912 ( .A(n3045), .B(n3007), .ZN(n3932) );
  OAI22_X1 U3913 ( .A1(n4435), .A2(n3126), .B1(n3088), .B2(n4550), .ZN(n3050)
         );
  AND2_X1 U3914 ( .A1(n3932), .A2(n3050), .ZN(n3047) );
  AOI21_X1 U3915 ( .B1(n4031), .B2(n3929), .A(n3047), .ZN(n3054) );
  OAI22_X1 U3916 ( .A1(n4010), .A2(n3088), .B1(n4432), .B2(n2955), .ZN(n3046)
         );
  XNOR2_X1 U3917 ( .A(n3046), .B(n3007), .ZN(n3945) );
  OAI22_X1 U3918 ( .A1(n4010), .A2(n3126), .B1(n4432), .B2(n3088), .ZN(n3055)
         );
  INV_X1 U3919 ( .A(n3047), .ZN(n3049) );
  INV_X1 U3920 ( .A(n3929), .ZN(n3048) );
  INV_X1 U3921 ( .A(n4031), .ZN(n3941) );
  NAND3_X1 U3922 ( .A1(n3049), .A2(n3048), .A3(n3941), .ZN(n3052) );
  INV_X1 U3923 ( .A(n3932), .ZN(n3051) );
  INV_X1 U3924 ( .A(n3050), .ZN(n3931) );
  NAND2_X1 U3925 ( .A1(n3051), .A2(n3931), .ZN(n3942) );
  OAI211_X1 U3926 ( .C1(n3945), .C2(n3055), .A(n3052), .B(n3942), .ZN(n3053)
         );
  INV_X1 U3927 ( .A(n3945), .ZN(n3056) );
  INV_X1 U3928 ( .A(n3055), .ZN(n3944) );
  NOR2_X1 U3929 ( .A1(n3056), .A2(n3944), .ZN(n3057) );
  OAI22_X1 U3930 ( .A1(n4543), .A2(n3088), .B1(n2955), .B2(n4411), .ZN(n3059)
         );
  XNOR2_X1 U3931 ( .A(n3059), .B(n3007), .ZN(n3061) );
  OAI22_X1 U3932 ( .A1(n4543), .A2(n3126), .B1(n3088), .B2(n4411), .ZN(n3062)
         );
  AND2_X1 U3933 ( .A1(n3061), .A2(n3062), .ZN(n4006) );
  INV_X1 U3934 ( .A(n4006), .ZN(n3060) );
  NAND2_X1 U3935 ( .A1(n4004), .A2(n3060), .ZN(n3065) );
  INV_X1 U3936 ( .A(n3061), .ZN(n3064) );
  INV_X1 U3937 ( .A(n3062), .ZN(n3063) );
  NAND2_X1 U3938 ( .A1(n3064), .A2(n3063), .ZN(n4005) );
  NAND2_X1 U3939 ( .A1(n3065), .A2(n4005), .ZN(n3892) );
  OAI22_X1 U3940 ( .A1(n4417), .A2(n3088), .B1(n2955), .B2(n4399), .ZN(n3066)
         );
  XNOR2_X1 U3941 ( .A(n3066), .B(n3007), .ZN(n3068) );
  OAI22_X1 U3942 ( .A1(n4417), .A2(n3126), .B1(n3088), .B2(n4399), .ZN(n3067)
         );
  XOR2_X1 U3943 ( .A(n3068), .B(n3067), .Z(n3893) );
  NAND2_X1 U3944 ( .A1(n4517), .A2(n3035), .ZN(n3071) );
  NAND2_X1 U3945 ( .A1(n3112), .A2(n4526), .ZN(n3070) );
  NAND2_X1 U3946 ( .A1(n3071), .A2(n3070), .ZN(n3072) );
  XNOR2_X1 U3947 ( .A(n3072), .B(n3007), .ZN(n3075) );
  NAND2_X1 U3948 ( .A1(n4517), .A2(n3116), .ZN(n3074) );
  NAND2_X1 U3949 ( .A1(n3029), .A2(n4526), .ZN(n3073) );
  NAND2_X1 U3950 ( .A1(n3074), .A2(n3073), .ZN(n3076) );
  NAND2_X1 U3951 ( .A1(n3075), .A2(n3076), .ZN(n3964) );
  INV_X1 U3952 ( .A(n3075), .ZN(n3078) );
  INV_X1 U3953 ( .A(n3076), .ZN(n3077) );
  NAND2_X1 U3954 ( .A1(n3078), .A2(n3077), .ZN(n3966) );
  NAND2_X1 U3955 ( .A1(n4378), .A2(n3035), .ZN(n3080) );
  NAND2_X1 U3956 ( .A1(n3112), .A2(n4516), .ZN(n3079) );
  NAND2_X1 U3957 ( .A1(n3080), .A2(n3079), .ZN(n3081) );
  XNOR2_X1 U3958 ( .A(n3081), .B(n3007), .ZN(n3908) );
  NAND2_X1 U3959 ( .A1(n4378), .A2(n3116), .ZN(n3083) );
  NAND2_X1 U3960 ( .A1(n3035), .A2(n4516), .ZN(n3082) );
  NAND2_X1 U3961 ( .A1(n3083), .A2(n3082), .ZN(n3907) );
  NOR2_X1 U3962 ( .A1(n3908), .A2(n3907), .ZN(n3085) );
  NAND2_X1 U3963 ( .A1(n3908), .A2(n3907), .ZN(n3084) );
  OAI22_X1 U3964 ( .A1(n4520), .A2(n3088), .B1(n3984), .B2(n2955), .ZN(n3086)
         );
  XNOR2_X1 U3965 ( .A(n3086), .B(n3007), .ZN(n3092) );
  OAI22_X1 U3966 ( .A1(n4520), .A2(n3126), .B1(n3984), .B2(n3088), .ZN(n3091)
         );
  XNOR2_X1 U3967 ( .A(n3092), .B(n3091), .ZN(n3982) );
  OAI22_X1 U3968 ( .A1(n4333), .A2(n3088), .B1(n3090), .B2(n2955), .ZN(n3089)
         );
  XNOR2_X1 U3969 ( .A(n3089), .B(n3007), .ZN(n3098) );
  OAI22_X1 U3970 ( .A1(n4333), .A2(n3126), .B1(n3090), .B2(n3088), .ZN(n3097)
         );
  XNOR2_X1 U3971 ( .A(n3098), .B(n3097), .ZN(n3885) );
  NOR2_X1 U3972 ( .A1(n3092), .A2(n3091), .ZN(n3886) );
  NOR2_X1 U3973 ( .A1(n3885), .A2(n3886), .ZN(n3093) );
  NAND2_X1 U3974 ( .A1(n4298), .A2(n3035), .ZN(n3095) );
  NAND2_X1 U3975 ( .A1(n3112), .A2(n4493), .ZN(n3094) );
  NAND2_X1 U3976 ( .A1(n3095), .A2(n3094), .ZN(n3096) );
  XNOR2_X1 U3977 ( .A(n3096), .B(n3007), .ZN(n3853) );
  OAI22_X1 U3978 ( .A1(n4023), .A2(n3126), .B1(n3088), .B2(n4285), .ZN(n3854)
         );
  NAND2_X1 U3979 ( .A1(n3853), .A2(n3854), .ZN(n3852) );
  NAND2_X1 U3980 ( .A1(n3098), .A2(n3097), .ZN(n3850) );
  INV_X1 U3981 ( .A(n3850), .ZN(n3103) );
  NAND2_X1 U3982 ( .A1(n4494), .A2(n3035), .ZN(n3100) );
  NAND2_X1 U3983 ( .A1(n3112), .A2(n3957), .ZN(n3099) );
  NAND2_X1 U3984 ( .A1(n3100), .A2(n3099), .ZN(n3101) );
  XNOR2_X1 U3985 ( .A(n3101), .B(n3007), .ZN(n3105) );
  NOR2_X1 U3986 ( .A1(n4303), .A2(n3088), .ZN(n3102) );
  AOI21_X1 U3987 ( .B1(n4494), .B2(n3116), .A(n3102), .ZN(n3849) );
  NAND2_X1 U3988 ( .A1(n3850), .A2(n3849), .ZN(n3847) );
  OAI21_X1 U3989 ( .B1(n3103), .B2(n3105), .A(n3847), .ZN(n3104) );
  NAND2_X1 U3990 ( .A1(n3851), .A2(n2157), .ZN(n3111) );
  INV_X1 U3991 ( .A(n3854), .ZN(n3107) );
  AOI21_X1 U3992 ( .B1(n3954), .B2(n3849), .A(n3107), .ZN(n3106) );
  NAND3_X1 U3993 ( .A1(n3954), .A2(n3107), .A3(n3849), .ZN(n3108) );
  NAND2_X1 U3994 ( .A1(n3111), .A2(n3110), .ZN(n4015) );
  NAND2_X1 U3995 ( .A1(n4483), .A2(n3035), .ZN(n3114) );
  NAND2_X1 U3996 ( .A1(n3112), .A2(n4019), .ZN(n3113) );
  NAND2_X1 U3997 ( .A1(n3114), .A2(n3113), .ZN(n3115) );
  XNOR2_X1 U3998 ( .A(n3115), .B(n3007), .ZN(n3119) );
  NAND2_X1 U3999 ( .A1(n4483), .A2(n3116), .ZN(n3118) );
  NAND2_X1 U4000 ( .A1(n3035), .A2(n4019), .ZN(n3117) );
  NAND2_X1 U4001 ( .A1(n3118), .A2(n3117), .ZN(n3120) );
  NAND2_X1 U4002 ( .A1(n3119), .A2(n3120), .ZN(n4016) );
  NAND2_X1 U4003 ( .A1(n4015), .A2(n4016), .ZN(n3123) );
  INV_X1 U4004 ( .A(n3119), .ZN(n3122) );
  INV_X1 U4005 ( .A(n3120), .ZN(n3121) );
  NAND2_X1 U4006 ( .A1(n3122), .A2(n3121), .ZN(n4017) );
  OAI22_X1 U4007 ( .A1(n3812), .A2(n3088), .B1(n2955), .B2(n3125), .ZN(n3124)
         );
  XNOR2_X1 U4008 ( .A(n3124), .B(n3007), .ZN(n3139) );
  OAI22_X1 U4009 ( .A1(n3812), .A2(n3126), .B1(n3088), .B2(n3125), .ZN(n3138)
         );
  XNOR2_X1 U4010 ( .A(n3139), .B(n3138), .ZN(n3865) );
  OAI22_X1 U4011 ( .A1(n4486), .A2(n3126), .B1(n3128), .B2(n3088), .ZN(n3127)
         );
  XNOR2_X1 U4012 ( .A(n3127), .B(n3007), .ZN(n3130) );
  OAI22_X1 U4013 ( .A1(n4486), .A2(n3088), .B1(n3128), .B2(n2955), .ZN(n3129)
         );
  XNOR2_X1 U4014 ( .A(n3130), .B(n3129), .ZN(n3137) );
  NAND3_X1 U4015 ( .A1(n3133), .A2(n3132), .A3(n3131), .ZN(n3155) );
  INV_X1 U4016 ( .A(n3213), .ZN(n3134) );
  OAI21_X1 U4017 ( .B1(n4190), .B2(n3310), .A(n3134), .ZN(n3135) );
  OR2_X1 U4018 ( .A1(n3135), .A2(n4570), .ZN(n3145) );
  NOR2_X1 U4019 ( .A1(n3211), .A2(n3145), .ZN(n3136) );
  INV_X1 U4020 ( .A(n3137), .ZN(n3160) );
  NAND2_X1 U4021 ( .A1(n3139), .A2(n3138), .ZN(n3159) );
  NOR2_X1 U4022 ( .A1(n3140), .A2(n4041), .ZN(n3141) );
  NAND2_X1 U4023 ( .A1(n3142), .A2(n2462), .ZN(n3164) );
  NAND2_X1 U4024 ( .A1(n3144), .A2(n3150), .ZN(n3152) );
  NAND2_X1 U4025 ( .A1(n3145), .A2(n4593), .ZN(n3146) );
  NAND2_X1 U4026 ( .A1(n3155), .A2(n3146), .ZN(n3148) );
  NAND2_X1 U4027 ( .A1(n3148), .A2(n3147), .ZN(n3825) );
  NAND2_X1 U4028 ( .A1(n2943), .A2(n3212), .ZN(n3149) );
  OAI21_X1 U4029 ( .B1(n3825), .B2(n3149), .A(STATE_REG_SCAN_IN), .ZN(n3151)
         );
  NAND2_X1 U4030 ( .A1(n3155), .A2(n3150), .ZN(n3826) );
  INV_X1 U4031 ( .A(n3152), .ZN(n3153) );
  NAND2_X1 U4032 ( .A1(n4199), .A2(n4025), .ZN(n3158) );
  NAND2_X1 U4033 ( .A1(n3827), .A2(n4570), .ZN(n3154) );
  AOI22_X1 U4034 ( .A1(n3156), .A2(n3839), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3157) );
  OAI211_X1 U4035 ( .C1(n4003), .C2(n3842), .A(n3158), .B(n3157), .ZN(n3162)
         );
  NOR3_X1 U4036 ( .A1(n3160), .A2(n4041), .A3(n3159), .ZN(n3161) );
  AOI211_X1 U4037 ( .C1(n3934), .C2(n4200), .A(n3162), .B(n3161), .ZN(n3163)
         );
  NAND3_X1 U4038 ( .A1(n3165), .A2(n3164), .A3(n3163), .ZN(U3217) );
  NAND2_X1 U4039 ( .A1(n3166), .A2(n4598), .ZN(n3168) );
  OR2_X1 U4040 ( .A1(n3175), .A2(n5079), .ZN(n3171) );
  INV_X1 U4041 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3169) );
  NAND2_X1 U4042 ( .A1(n5079), .A2(n3169), .ZN(n3170) );
  NAND2_X1 U40430 ( .A1(n3171), .A2(n3170), .ZN(n3172) );
  NAND2_X1 U4044 ( .A1(n3172), .A2(n2474), .ZN(U3547) );
  OR2_X1 U4045 ( .A1(n3175), .A2(n5075), .ZN(n3177) );
  NAND2_X1 U4046 ( .A1(n5075), .A2(n2832), .ZN(n3176) );
  NAND2_X1 U4047 ( .A1(n3177), .A2(n3176), .ZN(n3179) );
  NAND2_X1 U4048 ( .A1(n3179), .A2(n2473), .ZN(U3515) );
  NOR2_X1 U4049 ( .A1(n3254), .A2(REG1_REG_17__SCAN_IN), .ZN(n3209) );
  NAND2_X1 U4050 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3250), .ZN(n3206) );
  INV_X1 U4051 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4871) );
  MUX2_X1 U4052 ( .A(n4871), .B(REG1_REG_2__SCAN_IN), .S(n3345), .Z(n3348) );
  XNOR2_X1 U4053 ( .A(n4210), .B(REG1_REG_1__SCAN_IN), .ZN(n4215) );
  INV_X1 U4054 ( .A(n3180), .ZN(n4214) );
  NAND2_X1 U4055 ( .A1(n4215), .A2(n4214), .ZN(n4213) );
  INV_X1 U4056 ( .A(n4210), .ZN(n4958) );
  NAND2_X1 U4057 ( .A1(n4958), .A2(REG1_REG_1__SCAN_IN), .ZN(n3181) );
  NAND2_X1 U4058 ( .A1(n4213), .A2(n3181), .ZN(n3347) );
  NOR2_X2 U4059 ( .A1(n3294), .A2(n3186), .ZN(n3187) );
  INV_X1 U4060 ( .A(REG1_REG_4__SCAN_IN), .ZN(n5077) );
  INV_X1 U4061 ( .A(n3187), .ZN(n3188) );
  XNOR2_X1 U4062 ( .A(n4956), .B(REG1_REG_5__SCAN_IN), .ZN(n3301) );
  INV_X1 U4063 ( .A(n3190), .ZN(n3191) );
  INV_X1 U4064 ( .A(n3230), .ZN(n3392) );
  XNOR2_X1 U4065 ( .A(n3190), .B(n3392), .ZN(n3394) );
  INV_X1 U4066 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3457) );
  INV_X1 U4067 ( .A(REG1_REG_7__SCAN_IN), .ZN(n3414) );
  AND2_X2 U4068 ( .A1(n3193), .A2(n3192), .ZN(n3194) );
  NAND2_X1 U4069 ( .A1(n3509), .A2(REG1_REG_8__SCAN_IN), .ZN(n3196) );
  INV_X1 U4070 ( .A(n4955), .ZN(n3513) );
  OR2_X1 U4071 ( .A1(n3194), .A2(n3513), .ZN(n3195) );
  MUX2_X1 U4072 ( .A(REG1_REG_9__SCAN_IN), .B(n3197), .S(n4954), .Z(n3596) );
  NAND2_X1 U4073 ( .A1(n3597), .A2(n3596), .ZN(n3595) );
  NAND2_X1 U4074 ( .A1(n4954), .A2(REG1_REG_9__SCAN_IN), .ZN(n3198) );
  NAND2_X2 U4075 ( .A1(n3595), .A2(n3198), .ZN(n3199) );
  NAND2_X1 U4076 ( .A1(n3671), .A2(REG1_REG_10__SCAN_IN), .ZN(n3201) );
  NAND2_X1 U4077 ( .A1(n3199), .A2(n3239), .ZN(n3200) );
  MUX2_X1 U4078 ( .A(REG1_REG_11__SCAN_IN), .B(n3747), .S(n4953), .Z(n4223) );
  NAND2_X1 U4079 ( .A1(n4953), .A2(REG1_REG_11__SCAN_IN), .ZN(n3202) );
  INV_X1 U4080 ( .A(n4951), .ZN(n3800) );
  NAND2_X1 U4081 ( .A1(n3796), .A2(REG1_REG_12__SCAN_IN), .ZN(n3205) );
  NAND2_X1 U4082 ( .A1(n3203), .A2(n4951), .ZN(n3204) );
  NAND2_X2 U4083 ( .A1(n3205), .A2(n3204), .ZN(n4977) );
  INV_X1 U4084 ( .A(n3247), .ZN(n5059) );
  AOI22_X1 U4085 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3247), .B1(n5059), .B2(
        n4586), .ZN(n4978) );
  INV_X1 U4086 ( .A(n3273), .ZN(n4240) );
  INV_X1 U4087 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4842) );
  AOI22_X1 U4088 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3250), .B1(n5057), .B2(
        n4842), .ZN(n4988) );
  NAND2_X1 U4089 ( .A1(n3206), .A2(n4986), .ZN(n3207) );
  NOR2_X1 U4090 ( .A1(n5054), .A2(n3207), .ZN(n3208) );
  AOI22_X1 U4091 ( .A1(n3254), .A2(n4547), .B1(REG1_REG_17__SCAN_IN), .B2(
        n5053), .ZN(n5011) );
  AOI22_X1 U4092 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3255), .B1(n5052), .B2(
        n4827), .ZN(n5021) );
  MUX2_X1 U4093 ( .A(REG1_REG_19__SCAN_IN), .B(n4536), .S(n4190), .Z(n3210) );
  OR2_X1 U4094 ( .A1(n3212), .A2(U3149), .ZN(n4196) );
  NAND2_X1 U4095 ( .A1(n3211), .A2(n4196), .ZN(n3260) );
  NAND2_X1 U4096 ( .A1(n3213), .A2(n3212), .ZN(n3214) );
  AND2_X1 U4097 ( .A1(n4056), .A2(n3214), .ZN(n3258) );
  NAND2_X1 U4098 ( .A1(n3260), .A2(n3258), .ZN(n4969) );
  INV_X1 U4099 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4831) );
  AOI22_X1 U4100 ( .A1(REG2_REG_18__SCAN_IN), .A2(n5052), .B1(n3255), .B2(
        n4831), .ZN(n5016) );
  AND2_X1 U4101 ( .A1(n5060), .A2(REG2_REG_0__SCAN_IN), .ZN(n3217) );
  NAND2_X1 U4102 ( .A1(n4958), .A2(REG2_REG_1__SCAN_IN), .ZN(n3218) );
  OR2_X1 U4103 ( .A1(n3345), .A2(REG2_REG_2__SCAN_IN), .ZN(n3220) );
  NAND2_X1 U4104 ( .A1(n2546), .A2(REG2_REG_2__SCAN_IN), .ZN(n3221) );
  NAND2_X1 U4105 ( .A1(n3349), .A2(n3221), .ZN(n3222) );
  NAND2_X1 U4106 ( .A1(n3292), .A2(REG2_REG_3__SCAN_IN), .ZN(n3224) );
  NAND2_X1 U4107 ( .A1(n3222), .A2(n4957), .ZN(n3223) );
  NAND2_X1 U4108 ( .A1(n3224), .A2(n3223), .ZN(n3225) );
  XNOR2_X1 U4109 ( .A(n3225), .B(n3369), .ZN(n3364) );
  NAND2_X1 U4110 ( .A1(n3364), .A2(REG2_REG_4__SCAN_IN), .ZN(n3227) );
  NAND2_X1 U4111 ( .A1(n3225), .A2(n2560), .ZN(n3226) );
  MUX2_X1 U4112 ( .A(REG2_REG_5__SCAN_IN), .B(n3228), .S(n4956), .Z(n3304) );
  NAND2_X1 U4113 ( .A1(n4956), .A2(REG2_REG_5__SCAN_IN), .ZN(n3229) );
  MUX2_X1 U4114 ( .A(n3233), .B(REG2_REG_7__SCAN_IN), .S(n3423), .Z(n3419) );
  OR2_X1 U4115 ( .A1(n3423), .A2(n3233), .ZN(n3234) );
  NAND2_X1 U4116 ( .A1(n3235), .A2(n4955), .ZN(n3236) );
  XNOR2_X1 U4117 ( .A(n4954), .B(n3611), .ZN(n3599) );
  NAND2_X1 U4118 ( .A1(n4954), .A2(REG2_REG_9__SCAN_IN), .ZN(n3238) );
  NAND2_X1 U4119 ( .A1(n3672), .A2(REG2_REG_10__SCAN_IN), .ZN(n3242) );
  NAND2_X1 U4120 ( .A1(n3240), .A2(n3239), .ZN(n3241) );
  NAND2_X1 U4121 ( .A1(n3242), .A2(n3241), .ZN(n4228) );
  MUX2_X1 U4122 ( .A(REG2_REG_11__SCAN_IN), .B(n3687), .S(n4953), .Z(n4227) );
  NAND2_X1 U4123 ( .A1(n4228), .A2(n4227), .ZN(n4226) );
  NAND2_X1 U4124 ( .A1(n4953), .A2(REG2_REG_11__SCAN_IN), .ZN(n3243) );
  NAND2_X1 U4125 ( .A1(n3797), .A2(REG2_REG_12__SCAN_IN), .ZN(n3246) );
  NAND2_X1 U4126 ( .A1(n3244), .A2(n4951), .ZN(n3245) );
  NOR2_X1 U4127 ( .A1(n2670), .A2(n5059), .ZN(n4970) );
  OR2_X1 U4128 ( .A1(n3247), .A2(REG2_REG_13__SCAN_IN), .ZN(n3248) );
  INV_X1 U4129 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4237) );
  NAND2_X1 U4130 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3250), .ZN(n3249) );
  OAI21_X1 U4131 ( .B1(REG2_REG_15__SCAN_IN), .B2(n3250), .A(n3249), .ZN(n4982) );
  INV_X1 U4132 ( .A(n5054), .ZN(n4996) );
  INV_X1 U4133 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4992) );
  NAND2_X1 U4134 ( .A1(n3251), .A2(n4996), .ZN(n3252) );
  NOR2_X1 U4135 ( .A1(n3254), .A2(REG2_REG_17__SCAN_IN), .ZN(n3253) );
  AOI21_X1 U4136 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3254), .A(n3253), .ZN(n5008) );
  MUX2_X1 U4137 ( .A(n2713), .B(REG2_REG_19__SCAN_IN), .S(n4190), .Z(n3256) );
  XNOR2_X1 U4138 ( .A(n3257), .B(n3256), .ZN(n3263) );
  NAND2_X1 U4139 ( .A1(n4966), .A2(n4959), .ZN(n4192) );
  NAND2_X1 U4140 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3895) );
  INV_X1 U4141 ( .A(n3258), .ZN(n3259) );
  NAND2_X1 U4142 ( .A1(n5018), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3261) );
  OAI211_X1 U4143 ( .C1(n5024), .C2(n4190), .A(n3895), .B(n3261), .ZN(n3262)
         );
  AOI21_X1 U4144 ( .B1(n3263), .B2(n5001), .A(n3262), .ZN(n3264) );
  NAND2_X1 U4145 ( .A1(n5075), .A2(n3266), .ZN(n3267) );
  NAND2_X1 U4146 ( .A1(n3268), .A2(n2153), .ZN(U3514) );
  MUX2_X1 U4147 ( .A(n3345), .B(n2544), .S(U3149), .Z(n3269) );
  INV_X1 U4148 ( .A(n3269), .ZN(U3350) );
  INV_X1 U4149 ( .A(DATAI_6_), .ZN(n3270) );
  MUX2_X1 U4150 ( .A(n3392), .B(n3270), .S(U3149), .Z(n3271) );
  INV_X1 U4151 ( .A(n3271), .ZN(U3346) );
  MUX2_X1 U4152 ( .A(n2558), .B(n3369), .S(STATE_REG_SCAN_IN), .Z(n3272) );
  INV_X1 U4153 ( .A(n3272), .ZN(U3348) );
  INV_X1 U4154 ( .A(DATAI_14_), .ZN(n3275) );
  NAND2_X1 U4155 ( .A1(n3273), .A2(STATE_REG_SCAN_IN), .ZN(n3274) );
  OAI21_X1 U4156 ( .B1(STATE_REG_SCAN_IN), .B2(n3275), .A(n3274), .ZN(U3338)
         );
  MUX2_X1 U4157 ( .A(n3276), .B(n3423), .S(STATE_REG_SCAN_IN), .Z(n3277) );
  INV_X1 U4158 ( .A(n3277), .ZN(U3345) );
  NAND2_X1 U4159 ( .A1(U3149), .A2(DATAI_25_), .ZN(n3278) );
  OAI21_X1 U4160 ( .B1(n3279), .B2(U3149), .A(n3278), .ZN(U3327) );
  INV_X1 U4161 ( .A(DATAI_29_), .ZN(n4815) );
  NAND2_X1 U4162 ( .A1(n3280), .A2(STATE_REG_SCAN_IN), .ZN(n3281) );
  OAI21_X1 U4163 ( .B1(STATE_REG_SCAN_IN), .B2(n4815), .A(n3281), .ZN(U3323)
         );
  INV_X1 U4164 ( .A(DATAI_30_), .ZN(n3284) );
  NAND2_X1 U4165 ( .A1(n3282), .A2(STATE_REG_SCAN_IN), .ZN(n3283) );
  OAI21_X1 U4166 ( .B1(STATE_REG_SCAN_IN), .B2(n3284), .A(n3283), .ZN(U3322)
         );
  INV_X1 U4167 ( .A(DATAI_10_), .ZN(n3285) );
  MUX2_X1 U4168 ( .A(n3675), .B(n3285), .S(U3149), .Z(n3286) );
  INV_X1 U4169 ( .A(n3286), .ZN(U3342) );
  INV_X1 U4170 ( .A(D_REG_0__SCAN_IN), .ZN(n3289) );
  NOR3_X1 U4171 ( .A1(n3287), .A2(n4947), .A3(n2879), .ZN(n3288) );
  AOI21_X1 U4172 ( .B1(n5048), .B2(n3289), .A(n3288), .ZN(U3458) );
  INV_X1 U4173 ( .A(n3290), .ZN(n3291) );
  AOI22_X1 U4174 ( .A1(n5048), .A2(n2911), .B1(n3291), .B2(n5049), .ZN(U3459)
         );
  XNOR2_X1 U4175 ( .A(n3292), .B(n3552), .ZN(n3298) );
  AOI22_X1 U4176 ( .A1(n5018), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3293) );
  OAI21_X1 U4177 ( .B1(n3184), .B2(n5024), .A(n3293), .ZN(n3297) );
  AOI211_X1 U4178 ( .C1(n3413), .C2(n3295), .A(n3294), .B(n4997), .ZN(n3296)
         );
  AOI211_X1 U4179 ( .C1(n5001), .C2(n3298), .A(n3297), .B(n3296), .ZN(n3299)
         );
  INV_X1 U4180 ( .A(n3299), .ZN(U3243) );
  AOI211_X1 U4181 ( .C1(n2174), .C2(n3301), .A(n4997), .B(n3300), .ZN(n3309)
         );
  INV_X1 U4182 ( .A(n4956), .ZN(n3307) );
  OAI211_X1 U4183 ( .C1(n3304), .C2(n3303), .A(n5001), .B(n3302), .ZN(n3306)
         );
  NOR2_X1 U4184 ( .A1(STATE_REG_SCAN_IN), .A2(n2569), .ZN(n3533) );
  AOI21_X1 U4185 ( .B1(n5018), .B2(ADDR_REG_5__SCAN_IN), .A(n3533), .ZN(n3305)
         );
  OAI211_X1 U4186 ( .C1(n5024), .C2(n3307), .A(n3306), .B(n3305), .ZN(n3308)
         );
  OR2_X1 U4187 ( .A1(n3309), .A2(n3308), .ZN(U3245) );
  INV_X1 U4188 ( .A(n3740), .ZN(n5064) );
  NAND2_X1 U4189 ( .A1(n3311), .A2(n2963), .ZN(n4117) );
  NAND2_X1 U4190 ( .A1(n4117), .A2(n3314), .ZN(n5029) );
  NOR2_X1 U4191 ( .A1(n3311), .A2(n3310), .ZN(n5027) );
  INV_X1 U4192 ( .A(n4465), .ZN(n3836) );
  INV_X1 U4193 ( .A(n3323), .ZN(n3683) );
  OAI21_X1 U4194 ( .B1(n3683), .B2(n4577), .A(n5029), .ZN(n3312) );
  OAI21_X1 U4195 ( .B1(n3836), .B2(n4573), .A(n3312), .ZN(n5025) );
  AOI211_X1 U4196 ( .C1(n5064), .C2(n5029), .A(n5027), .B(n5025), .ZN(n5062)
         );
  NAND2_X1 U4197 ( .A1(n5079), .A2(REG1_REG_0__SCAN_IN), .ZN(n3313) );
  OAI21_X1 U4198 ( .B1(n5062), .B2(n5079), .A(n3313), .ZN(U3518) );
  NOR2_X1 U4199 ( .A1(n5018), .A2(n4202), .ZN(U3148) );
  NAND2_X1 U4200 ( .A1(n4099), .A2(n3314), .ZN(n3315) );
  NAND2_X1 U4201 ( .A1(n3378), .A2(n3315), .ZN(n3320) );
  NAND2_X1 U4202 ( .A1(n2963), .A2(n4590), .ZN(n3317) );
  NAND2_X1 U4203 ( .A1(n2135), .A2(n4589), .ZN(n3316) );
  OAI211_X1 U4204 ( .C1(n3318), .C2(n4593), .A(n3317), .B(n3316), .ZN(n3319)
         );
  AOI21_X1 U4205 ( .B1(n3320), .B2(n4577), .A(n3319), .ZN(n3325) );
  OAI21_X1 U4206 ( .B1(n4099), .B2(n3322), .A(n3321), .ZN(n3460) );
  OR2_X1 U4207 ( .A1(n3460), .A2(n3323), .ZN(n3324) );
  NAND2_X1 U4208 ( .A1(n3325), .A2(n3324), .ZN(n3462) );
  NAND2_X1 U4209 ( .A1(n2968), .A2(n3832), .ZN(n3326) );
  NAND2_X1 U4210 ( .A1(n3326), .A2(n3386), .ZN(n3461) );
  OAI22_X1 U4211 ( .A1(n3460), .A2(n3740), .B1(n4551), .B2(n3461), .ZN(n3327)
         );
  NOR2_X1 U4212 ( .A1(n3462), .A2(n3327), .ZN(n5063) );
  NAND2_X1 U4213 ( .A1(n5079), .A2(REG1_REG_1__SCAN_IN), .ZN(n3328) );
  OAI21_X1 U4214 ( .B1(n5063), .B2(n5079), .A(n3328), .ZN(U3519) );
  INV_X1 U4215 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4686) );
  INV_X1 U4216 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3333) );
  NAND2_X1 U4217 ( .A1(n3329), .A2(REG1_REG_31__SCAN_IN), .ZN(n3332) );
  INV_X1 U4218 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4729) );
  OR2_X1 U4219 ( .A1(n3330), .A2(n4729), .ZN(n3331) );
  OAI211_X1 U4220 ( .C1(n3334), .C2(n3333), .A(n3332), .B(n3331), .ZN(n4246)
         );
  NAND2_X1 U4221 ( .A1(n4202), .A2(n4246), .ZN(n3335) );
  OAI21_X1 U4222 ( .B1(U4043), .B2(n4686), .A(n3335), .ZN(U3581) );
  NOR2_X1 U4223 ( .A1(n5060), .A2(REG1_REG_0__SCAN_IN), .ZN(n4961) );
  NOR2_X1 U4224 ( .A1(n2943), .A2(n4961), .ZN(n3336) );
  OR3_X1 U4225 ( .A1(n3338), .A2(n3337), .A3(n3336), .ZN(n3339) );
  AND2_X1 U4226 ( .A1(n3340), .A2(n3339), .ZN(n3833) );
  NOR3_X1 U4227 ( .A1(n3833), .A2(n4966), .A3(n3341), .ZN(n3343) );
  AOI21_X1 U4228 ( .B1(n4966), .B2(n4623), .A(n3341), .ZN(n4963) );
  NAND2_X1 U4229 ( .A1(n5060), .A2(REG2_REG_0__SCAN_IN), .ZN(n4216) );
  OAI22_X1 U4230 ( .A1(n4963), .A2(n5060), .B1(n4216), .B2(n4192), .ZN(n3342)
         );
  NOR3_X1 U4231 ( .A1(n3343), .A2(n4209), .A3(n3342), .ZN(n3372) );
  AOI22_X1 U4232 ( .A1(n5018), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3344) );
  OAI21_X1 U4233 ( .B1(n3345), .B2(n5024), .A(n3344), .ZN(n3355) );
  OAI21_X1 U4234 ( .B1(n3348), .B2(n3347), .A(n3346), .ZN(n3353) );
  OAI21_X1 U4235 ( .B1(n3351), .B2(n3350), .A(n3349), .ZN(n3352) );
  OAI22_X1 U4236 ( .A1(n4997), .A2(n3353), .B1(n5014), .B2(n3352), .ZN(n3354)
         );
  OR3_X1 U4237 ( .A1(n3372), .A2(n3355), .A3(n3354), .ZN(U3242) );
  INV_X1 U4238 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n4743) );
  NAND2_X1 U4239 ( .A1(n3582), .A2(n4202), .ZN(n3356) );
  OAI21_X1 U4240 ( .B1(n4202), .B2(n4743), .A(n3356), .ZN(U3556) );
  INV_X1 U4241 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4726) );
  NAND2_X1 U4242 ( .A1(n4555), .A2(n4202), .ZN(n3357) );
  OAI21_X1 U4243 ( .B1(n4202), .B2(n4726), .A(n3357), .ZN(U3567) );
  INV_X1 U4244 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n4733) );
  NAND2_X1 U4245 ( .A1(n3708), .A2(n4202), .ZN(n3358) );
  OAI21_X1 U4246 ( .B1(n4202), .B2(n4733), .A(n3358), .ZN(U3559) );
  INV_X1 U4247 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n4732) );
  NAND2_X1 U4248 ( .A1(n4454), .A2(n4202), .ZN(n3359) );
  OAI21_X1 U4249 ( .B1(n4202), .B2(n4732), .A(n3359), .ZN(U3565) );
  INV_X1 U4250 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n4664) );
  NAND2_X1 U4251 ( .A1(n3693), .A2(n4202), .ZN(n3360) );
  OAI21_X1 U4252 ( .B1(n4202), .B2(n4664), .A(n3360), .ZN(U3560) );
  INV_X1 U4253 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n4745) );
  NAND2_X1 U4254 ( .A1(n4588), .A2(n4202), .ZN(n3361) );
  OAI21_X1 U4255 ( .B1(n4202), .B2(n4745), .A(n3361), .ZN(U3563) );
  INV_X1 U4256 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n4744) );
  NAND2_X1 U4257 ( .A1(n3531), .A2(n4202), .ZN(n3362) );
  OAI21_X1 U4258 ( .B1(U4043), .B2(n4744), .A(n3362), .ZN(U3554) );
  INV_X1 U4259 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4666) );
  NAND2_X1 U4260 ( .A1(n4470), .A2(n4202), .ZN(n3363) );
  OAI21_X1 U4261 ( .B1(U4043), .B2(n4666), .A(n3363), .ZN(U3553) );
  XNOR2_X1 U4262 ( .A(n3364), .B(REG2_REG_4__SCAN_IN), .ZN(n3374) );
  AOI211_X1 U4263 ( .C1(n5077), .C2(n3366), .A(n4997), .B(n3365), .ZN(n3371)
         );
  NAND2_X1 U4264 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3468) );
  INV_X1 U4265 ( .A(n3468), .ZN(n3367) );
  AOI21_X1 U4266 ( .B1(n5018), .B2(ADDR_REG_4__SCAN_IN), .A(n3367), .ZN(n3368)
         );
  OAI21_X1 U4267 ( .B1(n5024), .B2(n3369), .A(n3368), .ZN(n3370) );
  NOR3_X1 U4268 ( .A1(n3372), .A2(n3371), .A3(n3370), .ZN(n3373) );
  OAI21_X1 U4269 ( .B1(n3374), .B2(n5014), .A(n3373), .ZN(U3244) );
  INV_X1 U4270 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4730) );
  NAND2_X1 U4271 ( .A1(n4517), .A2(n4202), .ZN(n3375) );
  OAI21_X1 U4272 ( .B1(U4043), .B2(n4730), .A(n3375), .ZN(U3570) );
  OAI21_X1 U4273 ( .B1(n3377), .B2(n4091), .A(n3376), .ZN(n4469) );
  INV_X1 U4274 ( .A(n4469), .ZN(n3385) );
  NAND3_X1 U4275 ( .A1(n3378), .A2(n4091), .A3(n4119), .ZN(n3379) );
  NAND2_X1 U4276 ( .A1(n3380), .A2(n3379), .ZN(n3381) );
  AOI22_X1 U4277 ( .A1(n4469), .A2(n3683), .B1(n4577), .B2(n3381), .ZN(n4463)
         );
  OAI22_X1 U4278 ( .A1(n3836), .A2(n4561), .B1(n3382), .B2(n4593), .ZN(n3383)
         );
  AOI21_X1 U4279 ( .B1(n4589), .B2(n4470), .A(n3383), .ZN(n3384) );
  OAI211_X1 U4280 ( .C1(n3385), .C2(n3740), .A(n4463), .B(n3384), .ZN(n4875)
         );
  NAND2_X1 U4281 ( .A1(n3386), .A2(n4468), .ZN(n3387) );
  NAND2_X1 U4282 ( .A1(n3406), .A2(n3387), .ZN(n4872) );
  OAI22_X1 U4283 ( .A1(n4945), .A2(n4872), .B1(n5076), .B2(n4705), .ZN(n3388)
         );
  AOI21_X1 U4284 ( .B1(n4875), .B2(n5076), .A(n3388), .ZN(n3389) );
  INV_X1 U4285 ( .A(n3389), .ZN(U3471) );
  XOR2_X1 U4286 ( .A(n3390), .B(REG2_REG_6__SCAN_IN), .Z(n3397) );
  NAND2_X1 U4287 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3522) );
  NAND2_X1 U4288 ( .A1(n5018), .A2(ADDR_REG_6__SCAN_IN), .ZN(n3391) );
  OAI211_X1 U4289 ( .C1(n5024), .C2(n3392), .A(n3522), .B(n3391), .ZN(n3396)
         );
  AOI211_X1 U4290 ( .C1(n3394), .C2(n3457), .A(n4997), .B(n3393), .ZN(n3395)
         );
  AOI211_X1 U4291 ( .C1(n5001), .C2(n3397), .A(n3396), .B(n3395), .ZN(n3398)
         );
  INV_X1 U4292 ( .A(n3398), .ZN(U3246) );
  XNOR2_X1 U4293 ( .A(n3400), .B(n4094), .ZN(n3557) );
  OAI21_X1 U4294 ( .B1(n4094), .B2(n3402), .A(n3401), .ZN(n3403) );
  AOI22_X1 U4295 ( .A1(n3403), .A2(n4577), .B1(n4590), .B2(n2135), .ZN(n3560)
         );
  AOI22_X1 U4296 ( .A1(n4589), .A2(n3531), .B1(n3405), .B2(n4570), .ZN(n3404)
         );
  OAI211_X1 U4297 ( .C1(n5069), .C2(n3557), .A(n3560), .B(n3404), .ZN(n3410)
         );
  INV_X1 U4298 ( .A(n3410), .ZN(n3409) );
  AND2_X1 U4299 ( .A1(n3406), .A2(n3405), .ZN(n3407) );
  NOR2_X1 U4300 ( .A1(n2145), .A2(n3407), .ZN(n3556) );
  AOI22_X1 U4301 ( .A1(n4935), .A2(n3556), .B1(REG0_REG_3__SCAN_IN), .B2(n5075), .ZN(n3408) );
  OAI21_X1 U4302 ( .B1(n3409), .B2(n5075), .A(n3408), .ZN(U3473) );
  NAND2_X1 U4303 ( .A1(n3410), .A2(n5081), .ZN(n3412) );
  NAND2_X1 U4304 ( .A1(n4582), .A2(n3556), .ZN(n3411) );
  OAI211_X1 U4305 ( .C1(n5081), .C2(n3413), .A(n3412), .B(n3411), .ZN(U3521)
         );
  XNOR2_X1 U4306 ( .A(n3423), .B(n3414), .ZN(n3416) );
  OAI21_X1 U4307 ( .B1(n3417), .B2(n3416), .A(n3215), .ZN(n3415) );
  AOI21_X1 U4308 ( .B1(n3417), .B2(n3416), .A(n3415), .ZN(n3425) );
  OAI211_X1 U4309 ( .C1(n3420), .C2(n3419), .A(n3418), .B(n5001), .ZN(n3422)
         );
  AND2_X1 U4310 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3658) );
  AOI21_X1 U4311 ( .B1(n5018), .B2(ADDR_REG_7__SCAN_IN), .A(n3658), .ZN(n3421)
         );
  OAI211_X1 U4312 ( .C1(n5024), .C2(n3423), .A(n3422), .B(n3421), .ZN(n3424)
         );
  OR2_X1 U4313 ( .A1(n3425), .A2(n3424), .ZN(U3247) );
  INV_X1 U4314 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4741) );
  NAND2_X1 U4315 ( .A1(n4356), .A2(n4202), .ZN(n3426) );
  OAI21_X1 U4316 ( .B1(n4202), .B2(n4741), .A(n3426), .ZN(U3572) );
  OAI21_X1 U4317 ( .B1(n2145), .B2(n2583), .A(n2941), .ZN(n3427) );
  NOR2_X1 U4318 ( .A1(n3427), .A2(n3491), .ZN(n5066) );
  NOR2_X1 U4319 ( .A1(n4451), .A2(n3467), .ZN(n3440) );
  INV_X1 U4320 ( .A(n4470), .ZN(n3428) );
  OAI21_X1 U4321 ( .B1(n3400), .B2(n3428), .A(n3553), .ZN(n3430) );
  NAND2_X1 U4322 ( .A1(n3400), .A2(n3428), .ZN(n3429) );
  NAND2_X1 U4323 ( .A1(n3430), .A2(n3429), .ZN(n3431) );
  XNOR2_X1 U4324 ( .A(n3431), .B(n4096), .ZN(n5065) );
  NAND2_X1 U4325 ( .A1(n5065), .A2(n3683), .ZN(n3439) );
  INV_X1 U4326 ( .A(n4096), .ZN(n3432) );
  XNOR2_X1 U4327 ( .A(n3433), .B(n3432), .ZN(n3437) );
  NAND2_X1 U4328 ( .A1(n4207), .A2(n4589), .ZN(n3435) );
  NAND2_X1 U4329 ( .A1(n4470), .A2(n4590), .ZN(n3434) );
  OAI211_X1 U4330 ( .C1(n2583), .C2(n4593), .A(n3435), .B(n3434), .ZN(n3436)
         );
  AOI21_X1 U4331 ( .B1(n3437), .B2(n4577), .A(n3436), .ZN(n3438) );
  NAND2_X1 U4332 ( .A1(n3439), .A2(n3438), .ZN(n5068) );
  AOI211_X1 U4333 ( .C1(n5066), .C2(n4190), .A(n3440), .B(n5068), .ZN(n3444)
         );
  INV_X1 U4334 ( .A(n3441), .ZN(n3442) );
  NAND2_X1 U4335 ( .A1(n5032), .A2(n3442), .ZN(n3696) );
  INV_X1 U4336 ( .A(n3696), .ZN(n5030) );
  AOI22_X1 U4337 ( .A1(n5065), .A2(n5030), .B1(REG2_REG_4__SCAN_IN), .B2(n4337), .ZN(n3443) );
  OAI21_X1 U4338 ( .B1(n3444), .B2(n4337), .A(n3443), .ZN(U3286) );
  NAND2_X1 U4339 ( .A1(n4130), .A2(n4128), .ZN(n4098) );
  XOR2_X1 U4340 ( .A(n4098), .B(n3445), .Z(n3572) );
  OR2_X1 U4341 ( .A1(n3446), .A2(n3400), .ZN(n3489) );
  INV_X1 U4342 ( .A(n3447), .ZN(n3448) );
  NAND2_X1 U4343 ( .A1(n3489), .A2(n3448), .ZN(n3450) );
  AND2_X1 U4344 ( .A1(n3450), .A2(n2586), .ZN(n3583) );
  XNOR2_X1 U4345 ( .A(n3583), .B(n4098), .ZN(n3570) );
  AOI22_X1 U4346 ( .A1(n4590), .A2(n4207), .B1(n3567), .B2(n4570), .ZN(n3452)
         );
  NAND2_X1 U4347 ( .A1(n4206), .A2(n4589), .ZN(n3451) );
  OAI211_X1 U4348 ( .C1(n3570), .C2(n5069), .A(n3452), .B(n3451), .ZN(n3453)
         );
  AOI21_X1 U4349 ( .B1(n3572), .B2(n4577), .A(n3453), .ZN(n3459) );
  INV_X1 U4350 ( .A(n3575), .ZN(n3455) );
  AOI21_X1 U4351 ( .B1(n3567), .B2(n3454), .A(n3455), .ZN(n3566) );
  AOI22_X1 U4352 ( .A1(n3566), .A2(n4935), .B1(n5075), .B2(REG0_REG_6__SCAN_IN), .ZN(n3456) );
  OAI21_X1 U4353 ( .B1(n3459), .B2(n5075), .A(n3456), .ZN(U3479) );
  AOI22_X1 U4354 ( .A1(n3566), .A2(n4582), .B1(n5079), .B2(REG1_REG_6__SCAN_IN), .ZN(n3458) );
  OAI21_X1 U4355 ( .B1(n3459), .B2(n5079), .A(n3458), .ZN(U3524) );
  INV_X1 U4356 ( .A(n3460), .ZN(n3465) );
  OAI22_X1 U4357 ( .A1(n4458), .A2(n3461), .B1(n2518), .B2(n4451), .ZN(n3464)
         );
  MUX2_X1 U4358 ( .A(n3462), .B(REG2_REG_1__SCAN_IN), .S(n4337), .Z(n3463) );
  AOI211_X1 U4359 ( .C1(n3465), .C2(n5030), .A(n3464), .B(n3463), .ZN(n3466)
         );
  INV_X1 U4360 ( .A(n3466), .ZN(U3289) );
  INV_X1 U4361 ( .A(n3467), .ZN(n3475) );
  AOI22_X1 U4362 ( .A1(n3934), .A2(n4470), .B1(n4025), .B2(n4207), .ZN(n3469)
         );
  OAI211_X1 U4363 ( .C1(n3985), .C2(n2583), .A(n3469), .B(n3468), .ZN(n3474)
         );
  AOI211_X1 U4364 ( .C1(n3472), .C2(n3471), .A(n4041), .B(n3470), .ZN(n3473)
         );
  AOI211_X1 U4365 ( .C1(n3475), .C2(n4038), .A(n3474), .B(n3473), .ZN(n3476)
         );
  INV_X1 U4366 ( .A(n3476), .ZN(U3227) );
  XOR2_X1 U4367 ( .A(n3478), .B(n3477), .Z(n3484) );
  INV_X1 U4368 ( .A(n2135), .ZN(n3479) );
  OAI22_X1 U4369 ( .A1(n3985), .A2(n3553), .B1(n4033), .B2(n3479), .ZN(n3482)
         );
  INV_X1 U4370 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3480) );
  MUX2_X1 U4371 ( .A(U3149), .B(n4038), .S(n3480), .Z(n3481) );
  AOI211_X1 U4372 ( .C1(n4025), .C2(n3531), .A(n3482), .B(n3481), .ZN(n3483)
         );
  OAI21_X1 U4373 ( .B1(n3484), .B2(n4041), .A(n3483), .ZN(U3215) );
  INV_X1 U4374 ( .A(n4129), .ZN(n3485) );
  NAND2_X1 U4375 ( .A1(n3485), .A2(n4143), .ZN(n4089) );
  XOR2_X1 U4376 ( .A(n4089), .B(n3486), .Z(n3487) );
  NOR2_X1 U4377 ( .A1(n3487), .A2(n4425), .ZN(n3502) );
  INV_X1 U4378 ( .A(n3502), .ZN(n3500) );
  NAND2_X1 U4379 ( .A1(n3489), .A2(n3488), .ZN(n3490) );
  XOR2_X1 U4380 ( .A(n4089), .B(n3490), .Z(n3504) );
  INV_X1 U4381 ( .A(n3491), .ZN(n3493) );
  INV_X1 U4382 ( .A(n3454), .ZN(n3492) );
  AOI21_X1 U4383 ( .B1(n3534), .B2(n3493), .A(n3492), .ZN(n3506) );
  OAI22_X1 U4384 ( .A1(n5032), .A2(n3228), .B1(n3537), .B2(n4451), .ZN(n3494)
         );
  AOI21_X1 U4385 ( .B1(n3506), .B2(n4473), .A(n3494), .ZN(n3496) );
  AOI22_X1 U4386 ( .A1(n4471), .A2(n3582), .B1(n4466), .B2(n3531), .ZN(n3495)
         );
  OAI211_X1 U4387 ( .C1(n3497), .C2(n4433), .A(n3496), .B(n3495), .ZN(n3498)
         );
  AOI21_X1 U4388 ( .B1(n4460), .B2(n3504), .A(n3498), .ZN(n3499) );
  OAI21_X1 U4389 ( .B1(n3500), .B2(n4337), .A(n3499), .ZN(U3285) );
  AOI22_X1 U4390 ( .A1(n4590), .A2(n3531), .B1(n3534), .B2(n4570), .ZN(n3501)
         );
  OAI21_X1 U4391 ( .B1(n3656), .B2(n4573), .A(n3501), .ZN(n3503) );
  AOI211_X1 U4392 ( .C1(n3504), .C2(n4598), .A(n3503), .B(n3502), .ZN(n3508)
         );
  AOI22_X1 U4393 ( .A1(n3506), .A2(n4935), .B1(REG0_REG_5__SCAN_IN), .B2(n5075), .ZN(n3505) );
  OAI21_X1 U4394 ( .B1(n3508), .B2(n5075), .A(n3505), .ZN(U3477) );
  AOI22_X1 U4395 ( .A1(n3506), .A2(n4582), .B1(REG1_REG_5__SCAN_IN), .B2(n5079), .ZN(n3507) );
  OAI21_X1 U4396 ( .B1(n3508), .B2(n5079), .A(n3507), .ZN(U3523) );
  XNOR2_X1 U4397 ( .A(n3509), .B(REG1_REG_8__SCAN_IN), .ZN(n3517) );
  XOR2_X1 U4398 ( .A(n3510), .B(REG2_REG_8__SCAN_IN), .Z(n3511) );
  NAND2_X1 U4399 ( .A1(n5001), .A2(n3511), .ZN(n3512) );
  NAND2_X1 U4400 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3635) );
  NAND2_X1 U4401 ( .A1(n3512), .A2(n3635), .ZN(n3515) );
  NOR2_X1 U4402 ( .A1(n5024), .A2(n3513), .ZN(n3514) );
  AOI211_X1 U4403 ( .C1(n5018), .C2(ADDR_REG_8__SCAN_IN), .A(n3515), .B(n3514), 
        .ZN(n3516) );
  OAI21_X1 U4404 ( .B1(n3517), .B2(n4997), .A(n3516), .ZN(U3248) );
  XNOR2_X1 U4405 ( .A(n3519), .B(n3518), .ZN(n3520) );
  XNOR2_X1 U4406 ( .A(n3521), .B(n3520), .ZN(n3527) );
  INV_X1 U4407 ( .A(n3562), .ZN(n3525) );
  AOI22_X1 U4408 ( .A1(n3934), .A2(n4207), .B1(n4025), .B2(n4206), .ZN(n3523)
         );
  OAI211_X1 U4409 ( .C1(n3985), .C2(n2303), .A(n3523), .B(n3522), .ZN(n3524)
         );
  AOI21_X1 U4410 ( .B1(n3525), .B2(n4038), .A(n3524), .ZN(n3526) );
  OAI21_X1 U4411 ( .B1(n3527), .B2(n4041), .A(n3526), .ZN(U3236) );
  AOI211_X1 U4412 ( .C1(n2168), .C2(n3529), .A(n4041), .B(n3528), .ZN(n3530)
         );
  INV_X1 U4413 ( .A(n3530), .ZN(n3536) );
  OAI22_X1 U4414 ( .A1(n4034), .A2(n3656), .B1(n2567), .B2(n4033), .ZN(n3532)
         );
  AOI211_X1 U4415 ( .C1(n3534), .C2(n3156), .A(n3533), .B(n3532), .ZN(n3535)
         );
  OAI211_X1 U4416 ( .C1(n4003), .C2(n3537), .A(n3536), .B(n3535), .ZN(U3224)
         );
  INV_X1 U4417 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4727) );
  NAND2_X1 U4418 ( .A1(n4298), .A2(n4202), .ZN(n3538) );
  OAI21_X1 U4419 ( .B1(U4043), .B2(n4727), .A(n3538), .ZN(U3575) );
  NAND2_X1 U4420 ( .A1(n4137), .A2(n4135), .ZN(n4095) );
  XOR2_X1 U4421 ( .A(n3539), .B(n4095), .Z(n3624) );
  AND2_X1 U4422 ( .A1(n5032), .A2(n4577), .ZN(n4385) );
  INV_X1 U4423 ( .A(n4385), .ZN(n3651) );
  NOR2_X1 U4424 ( .A1(n3574), .A2(n3637), .ZN(n3541) );
  OR2_X1 U4425 ( .A1(n3540), .A2(n3541), .ZN(n3627) );
  INV_X1 U4426 ( .A(n3627), .ZN(n3550) );
  AOI22_X1 U4427 ( .A1(n4466), .A2(n4206), .B1(n4471), .B2(n3708), .ZN(n3544)
         );
  INV_X1 U4428 ( .A(n3542), .ZN(n3639) );
  INV_X1 U4429 ( .A(n4451), .ZN(n5028) );
  AOI22_X1 U4430 ( .A1(n4337), .A2(REG2_REG_8__SCAN_IN), .B1(n3639), .B2(n5028), .ZN(n3543) );
  OAI211_X1 U4431 ( .C1(n3637), .C2(n4433), .A(n3544), .B(n3543), .ZN(n3549)
         );
  NAND2_X1 U4432 ( .A1(n3545), .A2(n3546), .ZN(n3547) );
  XNOR2_X1 U4433 ( .A(n3547), .B(n4095), .ZN(n3620) );
  NOR2_X1 U4434 ( .A1(n3620), .A2(n4423), .ZN(n3548) );
  AOI211_X1 U4435 ( .C1(n3550), .C2(n4473), .A(n3549), .B(n3548), .ZN(n3551)
         );
  OAI21_X1 U4436 ( .B1(n3624), .B2(n3651), .A(n3551), .ZN(U3282) );
  OAI22_X1 U4437 ( .A1(n5032), .A2(n3552), .B1(REG3_REG_3__SCAN_IN), .B2(n4451), .ZN(n3555) );
  INV_X1 U4438 ( .A(n4471), .ZN(n3759) );
  OAI22_X1 U4439 ( .A1(n2567), .A2(n3759), .B1(n4433), .B2(n3553), .ZN(n3554)
         );
  AOI211_X1 U4440 ( .C1(n4473), .C2(n3556), .A(n3555), .B(n3554), .ZN(n3559)
         );
  OR2_X1 U4441 ( .A1(n3557), .A2(n4423), .ZN(n3558) );
  OAI211_X1 U4442 ( .C1(n4337), .C2(n3560), .A(n3559), .B(n3558), .ZN(U3287)
         );
  INV_X1 U4443 ( .A(n4466), .ZN(n4434) );
  INV_X1 U4444 ( .A(n4207), .ZN(n3561) );
  NOR2_X1 U4445 ( .A1(n4434), .A2(n3561), .ZN(n3565) );
  OAI22_X1 U4446 ( .A1(n5032), .A2(n3563), .B1(n3562), .B2(n4451), .ZN(n3564)
         );
  AOI211_X1 U4447 ( .C1(n3566), .C2(n4473), .A(n3565), .B(n3564), .ZN(n3569)
         );
  AOI22_X1 U4448 ( .A1(n4467), .A2(n3567), .B1(n4471), .B2(n4206), .ZN(n3568)
         );
  OAI211_X1 U4449 ( .C1(n4423), .C2(n3570), .A(n3569), .B(n3568), .ZN(n3571)
         );
  AOI21_X1 U4450 ( .B1(n3572), .B2(n4385), .A(n3571), .ZN(n3573) );
  INV_X1 U4451 ( .A(n3573), .ZN(U3284) );
  AOI211_X1 U4452 ( .C1(n3659), .C2(n3575), .A(n4551), .B(n3574), .ZN(n5072)
         );
  XNOR2_X1 U4453 ( .A(n3576), .B(n4131), .ZN(n3580) );
  OAI22_X1 U4454 ( .A1(n3656), .A2(n4561), .B1(n3577), .B2(n4593), .ZN(n3578)
         );
  AOI21_X1 U4455 ( .B1(n4589), .B2(n4205), .A(n3578), .ZN(n3579) );
  OAI21_X1 U4456 ( .B1(n3580), .B2(n4425), .A(n3579), .ZN(n5074) );
  AOI21_X1 U4457 ( .B1(n5072), .B2(n4190), .A(n5074), .ZN(n3593) );
  INV_X1 U4458 ( .A(n3583), .ZN(n3581) );
  NAND2_X1 U4459 ( .A1(n3581), .A2(n3656), .ZN(n3586) );
  NAND2_X1 U4460 ( .A1(n3583), .A2(n3582), .ZN(n3584) );
  NAND2_X1 U4461 ( .A1(n3584), .A2(n2303), .ZN(n3585) );
  AND2_X1 U4462 ( .A1(n3586), .A2(n3585), .ZN(n3587) );
  NOR2_X1 U4463 ( .A1(n3587), .A2(n4131), .ZN(n5071) );
  INV_X1 U4464 ( .A(n3587), .ZN(n3589) );
  INV_X1 U4465 ( .A(n4131), .ZN(n3588) );
  NOR2_X1 U4466 ( .A1(n3589), .A2(n3588), .ZN(n5070) );
  NOR3_X1 U4467 ( .A1(n5071), .A2(n5070), .A3(n4423), .ZN(n3591) );
  OAI22_X1 U4468 ( .A1(n5032), .A2(n3233), .B1(n3662), .B2(n4451), .ZN(n3590)
         );
  NOR2_X1 U4469 ( .A1(n3591), .A2(n3590), .ZN(n3592) );
  OAI21_X1 U4470 ( .B1(n3593), .B2(n4337), .A(n3592), .ZN(U3283) );
  INV_X1 U4471 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4704) );
  NAND2_X1 U4472 ( .A1(n4483), .A2(n4202), .ZN(n3594) );
  OAI21_X1 U4473 ( .B1(n4202), .B2(n4704), .A(n3594), .ZN(U3576) );
  INV_X1 U4474 ( .A(n4954), .ZN(n3605) );
  OAI211_X1 U4475 ( .C1(n3597), .C2(n3596), .A(n3595), .B(n3215), .ZN(n3604)
         );
  AND2_X1 U4476 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3702) );
  INV_X1 U4477 ( .A(n5018), .ZN(n5005) );
  INV_X1 U4478 ( .A(ADDR_REG_9__SCAN_IN), .ZN(n4852) );
  XOR2_X1 U4479 ( .A(n3599), .B(n3598), .Z(n3600) );
  NAND2_X1 U4480 ( .A1(n3600), .A2(n5001), .ZN(n3601) );
  OAI21_X1 U4481 ( .B1(n5005), .B2(n4852), .A(n3601), .ZN(n3602) );
  NOR2_X1 U4482 ( .A1(n3702), .A2(n3602), .ZN(n3603) );
  OAI211_X1 U4483 ( .C1(n5024), .C2(n3605), .A(n3604), .B(n3603), .ZN(U3249)
         );
  NAND2_X1 U4484 ( .A1(n2847), .A2(n4138), .ZN(n4101) );
  XOR2_X1 U4485 ( .A(n3606), .B(n4101), .Z(n3607) );
  NOR2_X1 U4486 ( .A1(n3607), .A2(n4425), .ZN(n3664) );
  INV_X1 U4487 ( .A(n3664), .ZN(n3619) );
  XOR2_X1 U4488 ( .A(n3608), .B(n4101), .Z(n3666) );
  INV_X1 U4489 ( .A(n3540), .ZN(n3610) );
  AOI21_X1 U4490 ( .B1(n3703), .B2(n3610), .A(n2314), .ZN(n3668) );
  INV_X1 U4491 ( .A(n3668), .ZN(n3616) );
  OAI22_X1 U4492 ( .A1(n5032), .A2(n3611), .B1(n3706), .B2(n4451), .ZN(n3614)
         );
  INV_X1 U4493 ( .A(n4205), .ZN(n3700) );
  OAI22_X1 U4494 ( .A1(n3700), .A2(n4434), .B1(n4433), .B2(n3612), .ZN(n3613)
         );
  AOI211_X1 U4495 ( .C1(n4471), .C2(n3693), .A(n3614), .B(n3613), .ZN(n3615)
         );
  OAI21_X1 U4496 ( .B1(n3616), .B2(n4458), .A(n3615), .ZN(n3617) );
  AOI21_X1 U4497 ( .B1(n4460), .B2(n3666), .A(n3617), .ZN(n3618) );
  OAI21_X1 U4498 ( .B1(n3619), .B2(n4337), .A(n3618), .ZN(U3281) );
  INV_X1 U4499 ( .A(n3708), .ZN(n3721) );
  OAI22_X1 U4500 ( .A1(n3721), .A2(n4573), .B1(n3637), .B2(n4593), .ZN(n3622)
         );
  NOR2_X1 U4501 ( .A1(n3620), .A2(n5069), .ZN(n3621) );
  AOI211_X1 U4502 ( .C1(n4590), .C2(n4206), .A(n3622), .B(n3621), .ZN(n3623)
         );
  OAI21_X1 U4503 ( .B1(n3624), .B2(n4425), .A(n3623), .ZN(n3629) );
  OAI22_X1 U4504 ( .A1(n3627), .A2(n4945), .B1(n5076), .B2(n4797), .ZN(n3625)
         );
  AOI21_X1 U4505 ( .B1(n3629), .B2(n5076), .A(n3625), .ZN(n3626) );
  INV_X1 U4506 ( .A(n3626), .ZN(U3483) );
  OAI22_X1 U4507 ( .A1(n3627), .A2(n4873), .B1(n5081), .B2(n4796), .ZN(n3628)
         );
  AOI21_X1 U4508 ( .B1(n3629), .B2(n5081), .A(n3628), .ZN(n3630) );
  INV_X1 U4509 ( .A(n3630), .ZN(U3526) );
  NAND2_X1 U4510 ( .A1(n3633), .A2(n3632), .ZN(n3634) );
  XNOR2_X1 U4511 ( .A(n3631), .B(n3634), .ZN(n3641) );
  AOI22_X1 U4512 ( .A1(n3934), .A2(n4206), .B1(n4025), .B2(n3708), .ZN(n3636)
         );
  OAI211_X1 U4513 ( .C1(n3985), .C2(n3637), .A(n3636), .B(n3635), .ZN(n3638)
         );
  AOI21_X1 U4514 ( .B1(n3639), .B2(n4038), .A(n3638), .ZN(n3640) );
  OAI21_X1 U4515 ( .B1(n3641), .B2(n4041), .A(n3640), .ZN(U3218) );
  NAND2_X1 U4516 ( .A1(n4146), .A2(n4149), .ZN(n4088) );
  XOR2_X1 U4517 ( .A(n4088), .B(n3642), .Z(n3712) );
  INV_X1 U4518 ( .A(n3712), .ZN(n3652) );
  XNOR2_X1 U4519 ( .A(n3643), .B(n4088), .ZN(n3707) );
  OAI21_X1 U4520 ( .B1(n2314), .B2(n3644), .A(n3688), .ZN(n3716) );
  INV_X1 U4521 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3645) );
  OAI22_X1 U4522 ( .A1(n5032), .A2(n3645), .B1(n3728), .B2(n4451), .ZN(n3647)
         );
  OAI22_X1 U4523 ( .A1(n3721), .A2(n4434), .B1(n3759), .B2(n3722), .ZN(n3646)
         );
  AOI211_X1 U4524 ( .C1(n3725), .C2(n4467), .A(n3647), .B(n3646), .ZN(n3648)
         );
  OAI21_X1 U4525 ( .B1(n3716), .B2(n4458), .A(n3648), .ZN(n3649) );
  AOI21_X1 U4526 ( .B1(n3707), .B2(n4460), .A(n3649), .ZN(n3650) );
  OAI21_X1 U4527 ( .B1(n3652), .B2(n3651), .A(n3650), .ZN(U3280) );
  XOR2_X1 U4528 ( .A(n3654), .B(n3653), .Z(n3655) );
  NAND2_X1 U4529 ( .A1(n3655), .A2(n3994), .ZN(n3661) );
  OAI22_X1 U4530 ( .A1(n4034), .A2(n3700), .B1(n3656), .B2(n4033), .ZN(n3657)
         );
  AOI211_X1 U4531 ( .C1(n3659), .C2(n3156), .A(n3658), .B(n3657), .ZN(n3660)
         );
  OAI211_X1 U4532 ( .C1(n4003), .C2(n3662), .A(n3661), .B(n3660), .ZN(U3210)
         );
  INV_X1 U4533 ( .A(n3693), .ZN(n3996) );
  AOI22_X1 U4534 ( .A1(n4590), .A2(n4205), .B1(n3703), .B2(n4570), .ZN(n3663)
         );
  OAI21_X1 U4535 ( .B1(n3996), .B2(n4573), .A(n3663), .ZN(n3665) );
  AOI211_X1 U4536 ( .C1(n3666), .C2(n4598), .A(n3665), .B(n3664), .ZN(n3670)
         );
  AOI22_X1 U4537 ( .A1(n3668), .A2(n4935), .B1(REG0_REG_9__SCAN_IN), .B2(n5075), .ZN(n3667) );
  OAI21_X1 U4538 ( .B1(n3670), .B2(n5075), .A(n3667), .ZN(U3485) );
  AOI22_X1 U4539 ( .A1(n3668), .A2(n4582), .B1(REG1_REG_9__SCAN_IN), .B2(n5079), .ZN(n3669) );
  OAI21_X1 U4540 ( .B1(n3670), .B2(n5079), .A(n3669), .ZN(U3527) );
  XNOR2_X1 U4541 ( .A(n3671), .B(REG1_REG_10__SCAN_IN), .ZN(n3679) );
  XOR2_X1 U4542 ( .A(n3672), .B(REG2_REG_10__SCAN_IN), .Z(n3673) );
  NAND2_X1 U4543 ( .A1(n5001), .A2(n3673), .ZN(n3674) );
  NAND2_X1 U4544 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n3720) );
  NAND2_X1 U4545 ( .A1(n3674), .A2(n3720), .ZN(n3677) );
  NOR2_X1 U4546 ( .A1(n5024), .A2(n3675), .ZN(n3676) );
  AOI211_X1 U4547 ( .C1(n5018), .C2(ADDR_REG_10__SCAN_IN), .A(n3677), .B(n3676), .ZN(n3678) );
  OAI21_X1 U4548 ( .B1(n3679), .B2(n4997), .A(n3678), .ZN(U3250) );
  OAI21_X1 U4549 ( .B1(n2171), .B2(n2470), .A(n3680), .ZN(n3684) );
  INV_X1 U4550 ( .A(n3684), .ZN(n3741) );
  XNOR2_X1 U4551 ( .A(n3681), .B(n2470), .ZN(n3686) );
  OAI22_X1 U4552 ( .A1(n3997), .A2(n4573), .B1(n3689), .B2(n4593), .ZN(n3682)
         );
  AOI21_X1 U4553 ( .B1(n3684), .B2(n3683), .A(n3682), .ZN(n3685) );
  OAI21_X1 U4554 ( .B1(n3686), .B2(n4425), .A(n3685), .ZN(n3743) );
  NAND2_X1 U4555 ( .A1(n3743), .A2(n5032), .ZN(n3695) );
  OAI22_X1 U4556 ( .A1(n5032), .A2(n3687), .B1(n4002), .B2(n4451), .ZN(n3692)
         );
  INV_X1 U4557 ( .A(n3688), .ZN(n3690) );
  OAI21_X1 U4558 ( .B1(n3690), .B2(n3689), .A(n3753), .ZN(n3749) );
  NOR2_X1 U4559 ( .A1(n3749), .A2(n4458), .ZN(n3691) );
  AOI211_X1 U4560 ( .C1(n4466), .C2(n3693), .A(n3692), .B(n3691), .ZN(n3694)
         );
  OAI211_X1 U4561 ( .C1(n3741), .C2(n3696), .A(n3695), .B(n3694), .ZN(U3279)
         );
  XNOR2_X1 U4562 ( .A(n3697), .B(n3698), .ZN(n3699) );
  NAND2_X1 U4563 ( .A1(n3699), .A2(n3994), .ZN(n3705) );
  OAI22_X1 U4564 ( .A1(n4034), .A2(n3996), .B1(n3700), .B2(n4033), .ZN(n3701)
         );
  AOI211_X1 U4565 ( .C1(n3703), .C2(n3156), .A(n3702), .B(n3701), .ZN(n3704)
         );
  OAI211_X1 U4566 ( .C1(n4003), .C2(n3706), .A(n3705), .B(n3704), .ZN(U3228)
         );
  NAND2_X1 U4567 ( .A1(n3707), .A2(n4598), .ZN(n3710) );
  AOI22_X1 U4568 ( .A1(n4590), .A2(n3708), .B1(n3725), .B2(n4570), .ZN(n3709)
         );
  OAI211_X1 U4569 ( .C1(n3722), .C2(n4573), .A(n3710), .B(n3709), .ZN(n3711)
         );
  AOI21_X1 U4570 ( .B1(n3712), .B2(n4577), .A(n3711), .ZN(n3714) );
  MUX2_X1 U4571 ( .A(n4765), .B(n3714), .S(n5076), .Z(n3713) );
  OAI21_X1 U4572 ( .B1(n3716), .B2(n4945), .A(n3713), .ZN(U3487) );
  MUX2_X1 U4573 ( .A(n4763), .B(n3714), .S(n5081), .Z(n3715) );
  OAI21_X1 U4574 ( .B1(n4873), .B2(n3716), .A(n3715), .ZN(U3528) );
  OAI211_X1 U4575 ( .C1(n3719), .C2(n3718), .A(n3717), .B(n3994), .ZN(n3727)
         );
  INV_X1 U4576 ( .A(n3720), .ZN(n3724) );
  OAI22_X1 U4577 ( .A1(n4034), .A2(n3722), .B1(n3721), .B2(n4033), .ZN(n3723)
         );
  AOI211_X1 U4578 ( .C1(n3725), .C2(n3156), .A(n3724), .B(n3723), .ZN(n3726)
         );
  OAI211_X1 U4579 ( .C1(n4003), .C2(n3728), .A(n3727), .B(n3726), .ZN(U3214)
         );
  OAI21_X1 U4580 ( .B1(n2170), .B2(n4100), .A(n3729), .ZN(n4576) );
  INV_X1 U4581 ( .A(n4576), .ZN(n3739) );
  INV_X1 U4582 ( .A(n3787), .ZN(n3730) );
  AOI21_X1 U4583 ( .B1(n4571), .B2(n3778), .A(n3730), .ZN(n4936) );
  AOI22_X1 U4584 ( .A1(n4471), .A2(n4454), .B1(n4466), .B2(n4588), .ZN(n3733)
         );
  INV_X1 U4585 ( .A(n3731), .ZN(n3882) );
  AOI22_X1 U4586 ( .A1(n4462), .A2(REG2_REG_14__SCAN_IN), .B1(n3882), .B2(
        n5028), .ZN(n3732) );
  OAI211_X1 U4587 ( .C1(n3880), .C2(n4433), .A(n3733), .B(n3732), .ZN(n3734)
         );
  AOI21_X1 U4588 ( .B1(n4936), .B2(n4473), .A(n3734), .ZN(n3738) );
  XNOR2_X1 U4589 ( .A(n3735), .B(n3736), .ZN(n4578) );
  NAND2_X1 U4590 ( .A1(n4578), .A2(n4385), .ZN(n3737) );
  OAI211_X1 U4591 ( .C1(n3739), .C2(n4423), .A(n3738), .B(n3737), .ZN(U3276)
         );
  INV_X1 U4592 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3744) );
  OAI22_X1 U4593 ( .A1(n3741), .A2(n3740), .B1(n3996), .B2(n4561), .ZN(n3742)
         );
  NOR2_X1 U4594 ( .A1(n3743), .A2(n3742), .ZN(n3746) );
  MUX2_X1 U4595 ( .A(n3744), .B(n3746), .S(n5076), .Z(n3745) );
  OAI21_X1 U4596 ( .B1(n3749), .B2(n4945), .A(n3745), .ZN(U3489) );
  MUX2_X1 U4597 ( .A(n3747), .B(n3746), .S(n5081), .Z(n3748) );
  OAI21_X1 U4598 ( .B1(n4873), .B2(n3749), .A(n3748), .ZN(U3529) );
  INV_X1 U4599 ( .A(n3767), .ZN(n3750) );
  NOR2_X1 U4600 ( .A1(n3768), .A2(n3750), .ZN(n4082) );
  XOR2_X1 U4601 ( .A(n4082), .B(n3769), .Z(n3751) );
  NOR2_X1 U4602 ( .A1(n3751), .A2(n4425), .ZN(n4595) );
  INV_X1 U4603 ( .A(n4595), .ZN(n3764) );
  XOR2_X1 U4604 ( .A(n4082), .B(n3752), .Z(n4597) );
  INV_X1 U4605 ( .A(n3753), .ZN(n3755) );
  INV_X1 U4606 ( .A(n3776), .ZN(n3754) );
  OAI21_X1 U4607 ( .B1(n3755), .B2(n4594), .A(n3754), .ZN(n4946) );
  NOR2_X1 U4608 ( .A1(n4946), .A2(n4458), .ZN(n3762) );
  INV_X1 U4609 ( .A(n4588), .ZN(n3760) );
  AOI22_X1 U4610 ( .A1(n4467), .A2(n3756), .B1(n4466), .B2(n4591), .ZN(n3758)
         );
  AOI22_X1 U4611 ( .A1(n4337), .A2(REG2_REG_12__SCAN_IN), .B1(n3925), .B2(
        n5028), .ZN(n3757) );
  OAI211_X1 U4612 ( .C1(n3760), .C2(n3759), .A(n3758), .B(n3757), .ZN(n3761)
         );
  AOI211_X1 U4613 ( .C1(n4597), .C2(n4460), .A(n3762), .B(n3761), .ZN(n3763)
         );
  OAI21_X1 U4614 ( .B1(n3764), .B2(n4462), .A(n3763), .ZN(U3278) );
  NAND2_X1 U4615 ( .A1(n3766), .A2(n3765), .ZN(n4090) );
  OAI21_X1 U4616 ( .B1(n3769), .B2(n3768), .A(n3767), .ZN(n3770) );
  XOR2_X1 U4617 ( .A(n4090), .B(n3770), .Z(n3773) );
  OAI22_X1 U4618 ( .A1(n3997), .A2(n4561), .B1(n3775), .B2(n4593), .ZN(n3771)
         );
  AOI21_X1 U4619 ( .B1(n4589), .B2(n4203), .A(n3771), .ZN(n3772) );
  OAI21_X1 U4620 ( .B1(n3773), .B2(n4425), .A(n3772), .ZN(n4584) );
  INV_X1 U4621 ( .A(n4584), .ZN(n3782) );
  XNOR2_X1 U4622 ( .A(n3774), .B(n4090), .ZN(n4585) );
  OR2_X1 U4623 ( .A1(n3776), .A2(n3775), .ZN(n3777) );
  NAND2_X1 U4624 ( .A1(n3778), .A2(n3777), .ZN(n4941) );
  AOI22_X1 U4625 ( .A1(n4337), .A2(REG2_REG_13__SCAN_IN), .B1(n3977), .B2(
        n5028), .ZN(n3779) );
  OAI21_X1 U4626 ( .B1(n4941), .B2(n4458), .A(n3779), .ZN(n3780) );
  AOI21_X1 U4627 ( .B1(n4585), .B2(n4460), .A(n3780), .ZN(n3781) );
  OAI21_X1 U4628 ( .B1(n3782), .B2(n4462), .A(n3781), .ZN(U3277) );
  AOI21_X1 U4629 ( .B1(n3783), .B2(n4080), .A(n4425), .ZN(n3785) );
  NAND2_X1 U4630 ( .A1(n3785), .A2(n3784), .ZN(n4565) );
  AOI21_X1 U4631 ( .B1(n4036), .B2(n3787), .A(n3786), .ZN(n4931) );
  NAND2_X1 U4632 ( .A1(n4471), .A2(n4564), .ZN(n3789) );
  NAND2_X1 U4633 ( .A1(n5028), .A2(n4037), .ZN(n3788) );
  OAI211_X1 U4634 ( .C1(n5032), .C2(n3790), .A(n3789), .B(n3788), .ZN(n3792)
         );
  OAI22_X1 U4635 ( .A1(n4562), .A2(n4434), .B1(n4433), .B2(n4560), .ZN(n3791)
         );
  AOI211_X1 U4636 ( .C1(n4931), .C2(n4473), .A(n3792), .B(n3791), .ZN(n3795)
         );
  XNOR2_X1 U4637 ( .A(n3793), .B(n4080), .ZN(n4559) );
  NAND2_X1 U4638 ( .A1(n4559), .A2(n4460), .ZN(n3794) );
  OAI211_X1 U4639 ( .C1(n4565), .C2(n4462), .A(n3795), .B(n3794), .ZN(U3275)
         );
  XNOR2_X1 U4640 ( .A(n3796), .B(REG1_REG_12__SCAN_IN), .ZN(n3804) );
  XOR2_X1 U4641 ( .A(REG2_REG_12__SCAN_IN), .B(n3797), .Z(n3798) );
  NAND2_X1 U4642 ( .A1(n5001), .A2(n3798), .ZN(n3799) );
  NAND2_X1 U4643 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n3922) );
  NAND2_X1 U4644 ( .A1(n3799), .A2(n3922), .ZN(n3802) );
  NOR2_X1 U4645 ( .A1(n5024), .A2(n3800), .ZN(n3801) );
  AOI211_X1 U4646 ( .C1(n5018), .C2(ADDR_REG_12__SCAN_IN), .A(n3802), .B(n3801), .ZN(n3803) );
  OAI21_X1 U4647 ( .B1(n3804), .B2(n4997), .A(n3803), .ZN(U3252) );
  INV_X1 U4648 ( .A(n3805), .ZN(n3807) );
  XNOR2_X1 U4649 ( .A(n3808), .B(n4108), .ZN(n4490) );
  NAND2_X1 U4650 ( .A1(n3809), .A2(n4076), .ZN(n3810) );
  XNOR2_X1 U4651 ( .A(n3810), .B(n4108), .ZN(n3814) );
  AOI22_X1 U4652 ( .A1(n4298), .A2(n4590), .B1(n4019), .B2(n4570), .ZN(n3811)
         );
  OAI21_X1 U4653 ( .B1(n3812), .B2(n4573), .A(n3811), .ZN(n3813) );
  AOI21_X1 U4654 ( .B1(n3814), .B2(n4577), .A(n3813), .ZN(n4489) );
  INV_X1 U4655 ( .A(n4489), .ZN(n3820) );
  INV_X1 U4656 ( .A(n3815), .ZN(n3817) );
  OAI21_X1 U4657 ( .B1(n3817), .B2(n3816), .A(n4263), .ZN(n4895) );
  AOI22_X1 U4658 ( .A1(n4020), .A2(n5028), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4337), .ZN(n3818) );
  OAI21_X1 U4659 ( .B1(n4895), .B2(n4458), .A(n3818), .ZN(n3819) );
  AOI21_X1 U4660 ( .B1(n3820), .B2(n5032), .A(n3819), .ZN(n3821) );
  OAI21_X1 U4661 ( .B1(n4490), .B2(n4423), .A(n3821), .ZN(U3264) );
  AOI21_X1 U4662 ( .B1(n3824), .B2(n3823), .A(n3822), .ZN(n3831) );
  AOI22_X1 U4663 ( .A1(n3934), .A2(n4465), .B1(n4468), .B2(n3156), .ZN(n3830)
         );
  INV_X1 U4664 ( .A(n3825), .ZN(n3828) );
  NAND3_X1 U4665 ( .A1(n3828), .A2(n3827), .A3(n3826), .ZN(n3900) );
  AOI22_X1 U4666 ( .A1(n3900), .A2(REG3_REG_2__SCAN_IN), .B1(n4025), .B2(n4470), .ZN(n3829) );
  OAI211_X1 U4667 ( .C1(n3831), .C2(n4041), .A(n3830), .B(n3829), .ZN(U3234)
         );
  AOI22_X1 U4668 ( .A1(n3994), .A2(n3833), .B1(n3156), .B2(n3832), .ZN(n3835)
         );
  NAND2_X1 U4669 ( .A1(n3900), .A2(REG3_REG_0__SCAN_IN), .ZN(n3834) );
  OAI211_X1 U4670 ( .C1(n4034), .C2(n3836), .A(n3835), .B(n3834), .ZN(U3229)
         );
  INV_X1 U4671 ( .A(n3837), .ZN(n3838) );
  NAND2_X1 U4672 ( .A1(n3838), .A2(n4460), .ZN(n3845) );
  NAND2_X1 U4673 ( .A1(n4199), .A2(n4471), .ZN(n3841) );
  AOI22_X1 U4674 ( .A1(n4467), .A2(n3839), .B1(n4462), .B2(
        REG2_REG_28__SCAN_IN), .ZN(n3840) );
  OAI211_X1 U4675 ( .C1(n4451), .C2(n3842), .A(n3841), .B(n3840), .ZN(n3844)
         );
  INV_X1 U4676 ( .A(n3847), .ZN(n3848) );
  OAI21_X1 U4677 ( .B1(n3854), .B2(n3853), .A(n3852), .ZN(n3855) );
  NAND2_X1 U4678 ( .A1(n3856), .A2(n3994), .ZN(n3861) );
  NOR2_X1 U4679 ( .A1(n4282), .A2(n4003), .ZN(n3859) );
  AOI22_X1 U4680 ( .A1(n3156), .A2(n4493), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3857) );
  OAI21_X1 U4681 ( .B1(n4314), .B2(n4033), .A(n3857), .ZN(n3858) );
  AOI211_X1 U4682 ( .C1(n4025), .C2(n4483), .A(n3859), .B(n3858), .ZN(n3860)
         );
  NAND2_X1 U4683 ( .A1(n3861), .A2(n3860), .ZN(U3222) );
  NAND3_X1 U4684 ( .A1(n3863), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3864) );
  INV_X1 U4685 ( .A(DATAI_31_), .ZN(n4687) );
  OAI22_X1 U4686 ( .A1(n3862), .A2(n3864), .B1(STATE_REG_SCAN_IN), .B2(n4687), 
        .ZN(U3321) );
  XNOR2_X1 U4687 ( .A(n3866), .B(n3865), .ZN(n3871) );
  AOI22_X1 U4688 ( .A1(n3156), .A2(n4482), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3868) );
  NAND2_X1 U4689 ( .A1(n4266), .A2(n4038), .ZN(n3867) );
  OAI211_X1 U4690 ( .C1(n4497), .C2(n4033), .A(n3868), .B(n3867), .ZN(n3869)
         );
  AOI21_X1 U4691 ( .B1(n4025), .B2(n4271), .A(n3869), .ZN(n3870) );
  OAI21_X1 U4692 ( .B1(n3871), .B2(n4041), .A(n3870), .ZN(U3211) );
  INV_X1 U4693 ( .A(n3974), .ZN(n3874) );
  INV_X1 U4694 ( .A(n3972), .ZN(n3873) );
  AOI21_X1 U4695 ( .B1(n3974), .B2(n3972), .A(n3971), .ZN(n3872) );
  AOI21_X1 U4696 ( .B1(n3874), .B2(n3873), .A(n3872), .ZN(n3878) );
  NAND2_X1 U4697 ( .A1(n3876), .A2(n3875), .ZN(n3877) );
  XNOR2_X1 U4698 ( .A(n3878), .B(n3877), .ZN(n3884) );
  AOI22_X1 U4699 ( .A1(n3934), .A2(n4588), .B1(n4025), .B2(n4454), .ZN(n3879)
         );
  NAND2_X1 U4700 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n4239) );
  OAI211_X1 U4701 ( .C1(n3985), .C2(n3880), .A(n3879), .B(n4239), .ZN(n3881)
         );
  AOI21_X1 U4702 ( .B1(n3882), .B2(n4038), .A(n3881), .ZN(n3883) );
  OAI21_X1 U4703 ( .B1(n3884), .B2(n4041), .A(n3883), .ZN(U3212) );
  OAI21_X1 U4704 ( .B1(n2150), .B2(n3886), .A(n3885), .ZN(n3887) );
  NAND3_X1 U4705 ( .A1(n3887), .A2(n3994), .A3(n3851), .ZN(n3891) );
  AOI22_X1 U4706 ( .A1(n3156), .A2(n4317), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3890) );
  AOI22_X1 U4707 ( .A1(n4494), .A2(n4025), .B1(n3934), .B2(n4356), .ZN(n3889)
         );
  NAND2_X1 U4708 ( .A1(n4320), .A2(n4038), .ZN(n3888) );
  NAND4_X1 U4709 ( .A1(n3891), .A2(n3890), .A3(n3889), .A4(n3888), .ZN(U3213)
         );
  XOR2_X1 U4710 ( .A(n3893), .B(n3892), .Z(n3899) );
  INV_X1 U4711 ( .A(n3894), .ZN(n4401) );
  AOI22_X1 U4712 ( .A1(n4517), .A2(n4025), .B1(n3934), .B2(n4438), .ZN(n3896)
         );
  OAI211_X1 U4713 ( .C1(n3985), .C2(n4399), .A(n3896), .B(n3895), .ZN(n3897)
         );
  AOI21_X1 U4714 ( .B1(n4401), .B2(n4038), .A(n3897), .ZN(n3898) );
  OAI21_X1 U4715 ( .B1(n3899), .B2(n4041), .A(n3898), .ZN(U3216) );
  AOI22_X1 U4716 ( .A1(n3900), .A2(REG3_REG_1__SCAN_IN), .B1(n4025), .B2(n2135), .ZN(n3906) );
  AOI22_X1 U4717 ( .A1(n3934), .A2(n2963), .B1(n2968), .B2(n3156), .ZN(n3905)
         );
  OAI211_X1 U4718 ( .C1(n3901), .C2(n3902), .A(n3903), .B(n3994), .ZN(n3904)
         );
  NAND3_X1 U4719 ( .A1(n3906), .A2(n3905), .A3(n3904), .ZN(U3219) );
  XNOR2_X1 U4720 ( .A(n3908), .B(n3907), .ZN(n3909) );
  XNOR2_X1 U4721 ( .A(n3910), .B(n3909), .ZN(n3917) );
  INV_X1 U4722 ( .A(n4354), .ZN(n3915) );
  OAI22_X1 U4723 ( .A1(n3985), .A2(n4350), .B1(STATE_REG_SCAN_IN), .B2(n3911), 
        .ZN(n3914) );
  OAI22_X1 U4724 ( .A1(n4520), .A2(n4034), .B1(n3912), .B2(n4033), .ZN(n3913)
         );
  AOI211_X1 U4725 ( .C1(n3915), .C2(n4038), .A(n3914), .B(n3913), .ZN(n3916)
         );
  OAI21_X1 U4726 ( .B1(n3917), .B2(n4041), .A(n3916), .ZN(U3220) );
  NOR2_X1 U4727 ( .A1(n3919), .A2(n2382), .ZN(n3920) );
  XNOR2_X1 U4728 ( .A(n3921), .B(n3920), .ZN(n3927) );
  AOI22_X1 U4729 ( .A1(n3934), .A2(n4591), .B1(n4025), .B2(n4588), .ZN(n3923)
         );
  OAI211_X1 U4730 ( .C1(n3985), .C2(n4594), .A(n3923), .B(n3922), .ZN(n3924)
         );
  AOI21_X1 U4731 ( .B1(n3925), .B2(n4038), .A(n3924), .ZN(n3926) );
  OAI21_X1 U4732 ( .B1(n3927), .B2(n4041), .A(n3926), .ZN(U3221) );
  INV_X1 U4733 ( .A(n3928), .ZN(n3930) );
  NAND2_X1 U4734 ( .A1(n3930), .A2(n3929), .ZN(n4028) );
  NOR2_X1 U4735 ( .A1(n3930), .A2(n3929), .ZN(n4030) );
  AOI21_X1 U4736 ( .B1(n3941), .B2(n4028), .A(n4030), .ZN(n3933) );
  XNOR2_X1 U4737 ( .A(n3932), .B(n3931), .ZN(n3940) );
  XNOR2_X1 U4738 ( .A(n3933), .B(n3940), .ZN(n3939) );
  INV_X1 U4739 ( .A(n4452), .ZN(n3937) );
  AOI22_X1 U4740 ( .A1(n3934), .A2(n4454), .B1(n4025), .B2(n4555), .ZN(n3935)
         );
  NAND2_X1 U4741 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n5002) );
  OAI211_X1 U4742 ( .C1(n3985), .C2(n4550), .A(n3935), .B(n5002), .ZN(n3936)
         );
  AOI21_X1 U4743 ( .B1(n3937), .B2(n4038), .A(n3936), .ZN(n3938) );
  OAI21_X1 U4744 ( .B1(n3939), .B2(n4041), .A(n3938), .ZN(U3223) );
  OAI211_X1 U4745 ( .C1(n4030), .C2(n3941), .A(n3940), .B(n4028), .ZN(n3943)
         );
  NAND2_X1 U4746 ( .A1(n3943), .A2(n3942), .ZN(n3947) );
  XNOR2_X1 U4747 ( .A(n3945), .B(n3944), .ZN(n3946) );
  XNOR2_X1 U4748 ( .A(n3947), .B(n3946), .ZN(n3948) );
  NAND2_X1 U4749 ( .A1(n3948), .A2(n3994), .ZN(n3951) );
  AND2_X1 U4750 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n5009) );
  OAI22_X1 U4751 ( .A1(n4034), .A2(n4543), .B1(n4435), .B2(n4033), .ZN(n3949)
         );
  AOI211_X1 U4752 ( .C1(n4541), .C2(n3156), .A(n5009), .B(n3949), .ZN(n3950)
         );
  OAI211_X1 U4753 ( .C1(n4003), .C2(n4430), .A(n3951), .B(n3950), .ZN(U3225)
         );
  NOR2_X1 U4754 ( .A1(n3953), .A2(n3952), .ZN(n3955) );
  XNOR2_X1 U4755 ( .A(n3955), .B(n3954), .ZN(n3956) );
  NAND2_X1 U4756 ( .A1(n3956), .A2(n3994), .ZN(n3962) );
  NAND2_X1 U4757 ( .A1(n4298), .A2(n4025), .ZN(n3959) );
  AOI22_X1 U4758 ( .A1(n3156), .A2(n3957), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3958) );
  OAI211_X1 U4759 ( .C1(n4333), .C2(n4033), .A(n3959), .B(n3958), .ZN(n3960)
         );
  AOI21_X1 U4760 ( .B1(n4305), .B2(n4038), .A(n3960), .ZN(n3961) );
  NAND2_X1 U4761 ( .A1(n3962), .A2(n3961), .ZN(U3226) );
  AOI21_X1 U4762 ( .B1(n3966), .B2(n3964), .A(n3963), .ZN(n3965) );
  AOI21_X1 U4763 ( .B1(n2156), .B2(n3966), .A(n3965), .ZN(n3970) );
  OAI22_X1 U4764 ( .A1(n3985), .A2(n4382), .B1(STATE_REG_SCAN_IN), .B2(n4812), 
        .ZN(n3968) );
  OAI22_X1 U4765 ( .A1(n4530), .A2(n4034), .B1(n4417), .B2(n4033), .ZN(n3967)
         );
  AOI211_X1 U4766 ( .C1(n4379), .C2(n4038), .A(n3968), .B(n3967), .ZN(n3969)
         );
  OAI21_X1 U4767 ( .B1(n3970), .B2(n4041), .A(n3969), .ZN(U3230) );
  XNOR2_X1 U4768 ( .A(n3972), .B(n3971), .ZN(n3973) );
  XNOR2_X1 U4769 ( .A(n3974), .B(n3973), .ZN(n3980) );
  NOR2_X1 U4770 ( .A1(n4758), .A2(STATE_REG_SCAN_IN), .ZN(n4975) );
  OAI22_X1 U4771 ( .A1(n4034), .A2(n4562), .B1(n3997), .B2(n4033), .ZN(n3975)
         );
  AOI211_X1 U4772 ( .C1(n3976), .C2(n3156), .A(n4975), .B(n3975), .ZN(n3979)
         );
  NAND2_X1 U4773 ( .A1(n4038), .A2(n3977), .ZN(n3978) );
  OAI211_X1 U4774 ( .C1(n3980), .C2(n4041), .A(n3979), .B(n3978), .ZN(U3231)
         );
  AOI21_X1 U4775 ( .B1(n3982), .B2(n3981), .A(n2150), .ZN(n3989) );
  INV_X1 U4776 ( .A(n3983), .ZN(n4338) );
  OAI22_X1 U4777 ( .A1(n3985), .A2(n3984), .B1(STATE_REG_SCAN_IN), .B2(n4810), 
        .ZN(n3987) );
  OAI22_X1 U4778 ( .A1(n4333), .A2(n4034), .B1(n4530), .B2(n4033), .ZN(n3986)
         );
  AOI211_X1 U4779 ( .C1(n4338), .C2(n4038), .A(n3987), .B(n3986), .ZN(n3988)
         );
  OAI21_X1 U4780 ( .B1(n3989), .B2(n4041), .A(n3988), .ZN(U3232) );
  XNOR2_X1 U4781 ( .A(n3992), .B(n3991), .ZN(n3993) );
  XNOR2_X1 U4782 ( .A(n3990), .B(n3993), .ZN(n3995) );
  NAND2_X1 U4783 ( .A1(n3995), .A2(n3994), .ZN(n4001) );
  AND2_X1 U4784 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4225) );
  OAI22_X1 U4785 ( .A1(n4034), .A2(n3997), .B1(n3996), .B2(n4033), .ZN(n3998)
         );
  AOI211_X1 U4786 ( .C1(n3999), .C2(n3156), .A(n4225), .B(n3998), .ZN(n4000)
         );
  OAI211_X1 U4787 ( .C1(n4003), .C2(n4002), .A(n4001), .B(n4000), .ZN(U3233)
         );
  INV_X1 U4788 ( .A(n4004), .ZN(n4009) );
  INV_X1 U4789 ( .A(n4005), .ZN(n4007) );
  NOR2_X1 U4790 ( .A1(n4007), .A2(n4006), .ZN(n4008) );
  XNOR2_X1 U4791 ( .A(n4009), .B(n4008), .ZN(n4014) );
  NOR2_X1 U4792 ( .A1(n4658), .A2(STATE_REG_SCAN_IN), .ZN(n5017) );
  OAI22_X1 U4793 ( .A1(n4034), .A2(n4417), .B1(n4010), .B2(n4033), .ZN(n4011)
         );
  AOI211_X1 U4794 ( .C1(n4415), .C2(n3156), .A(n5017), .B(n4011), .ZN(n4013)
         );
  NAND2_X1 U4795 ( .A1(n4038), .A2(n4409), .ZN(n4012) );
  OAI211_X1 U4796 ( .C1(n4014), .C2(n4041), .A(n4013), .B(n4012), .ZN(U3235)
         );
  NAND2_X1 U4797 ( .A1(n4017), .A2(n4016), .ZN(n4018) );
  XNOR2_X1 U4798 ( .A(n4015), .B(n4018), .ZN(n4027) );
  AOI22_X1 U4799 ( .A1(n3156), .A2(n4019), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n4022) );
  NAND2_X1 U4800 ( .A1(n4020), .A2(n4038), .ZN(n4021) );
  OAI211_X1 U4801 ( .C1(n4023), .C2(n4033), .A(n4022), .B(n4021), .ZN(n4024)
         );
  AOI21_X1 U4802 ( .B1(n4200), .B2(n4025), .A(n4024), .ZN(n4026) );
  OAI21_X1 U4803 ( .B1(n4027), .B2(n4041), .A(n4026), .ZN(U3237) );
  INV_X1 U4804 ( .A(n4028), .ZN(n4029) );
  NOR2_X1 U4805 ( .A1(n4030), .A2(n4029), .ZN(n4032) );
  XNOR2_X1 U4806 ( .A(n4032), .B(n4031), .ZN(n4042) );
  NOR2_X1 U4807 ( .A1(n4761), .A2(STATE_REG_SCAN_IN), .ZN(n4985) );
  OAI22_X1 U4808 ( .A1(n4034), .A2(n4435), .B1(n4562), .B2(n4033), .ZN(n4035)
         );
  AOI211_X1 U4809 ( .C1(n4036), .C2(n3156), .A(n4985), .B(n4035), .ZN(n4040)
         );
  NAND2_X1 U4810 ( .A1(n4038), .A2(n4037), .ZN(n4039) );
  OAI211_X1 U4811 ( .C1(n4042), .C2(n4041), .A(n4040), .B(n4039), .ZN(U3238)
         );
  NAND2_X1 U4812 ( .A1(n4046), .A2(n4043), .ZN(n4155) );
  NAND2_X1 U4813 ( .A1(n4045), .A2(n4044), .ZN(n4140) );
  NAND2_X1 U4814 ( .A1(n4140), .A2(n4046), .ZN(n4158) );
  OAI21_X1 U4815 ( .B1(n3735), .B2(n4155), .A(n4158), .ZN(n4048) );
  INV_X1 U4816 ( .A(n4162), .ZN(n4047) );
  AOI211_X1 U4817 ( .C1(n4048), .C2(n4166), .A(n4047), .B(n4165), .ZN(n4050)
         );
  OAI21_X1 U4818 ( .B1(n4050), .B2(n2389), .A(n4169), .ZN(n4052) );
  AOI21_X1 U4819 ( .B1(n4052), .B2(n4172), .A(n4051), .ZN(n4055) );
  INV_X1 U4820 ( .A(n4077), .ZN(n4053) );
  AOI211_X1 U4821 ( .C1(n4173), .C2(n4054), .A(n4053), .B(n4075), .ZN(n4174)
         );
  OAI21_X1 U4822 ( .B1(n4055), .B2(n2195), .A(n4174), .ZN(n4060) );
  INV_X1 U4823 ( .A(n4066), .ZN(n4059) );
  NAND2_X1 U4824 ( .A1(n4056), .A2(DATAI_31_), .ZN(n4247) );
  NAND2_X1 U4825 ( .A1(n4246), .A2(n4247), .ZN(n4182) );
  AND2_X1 U4826 ( .A1(n4056), .A2(DATAI_30_), .ZN(n4252) );
  INV_X1 U4827 ( .A(n4252), .ZN(n4071) );
  OR2_X1 U4828 ( .A1(n4198), .A2(n4071), .ZN(n4057) );
  AND2_X1 U4829 ( .A1(n4182), .A2(n4057), .ZN(n4086) );
  AND2_X1 U4830 ( .A1(n4058), .A2(n4086), .ZN(n4064) );
  NAND4_X1 U4831 ( .A1(n4060), .A2(n4059), .A3(n4175), .A4(n4064), .ZN(n4070)
         );
  INV_X1 U4832 ( .A(n4258), .ZN(n4113) );
  AND2_X1 U4833 ( .A1(n4062), .A2(n4061), .ZN(n4067) );
  NAND2_X1 U4834 ( .A1(n4067), .A2(n2404), .ZN(n4115) );
  INV_X1 U4835 ( .A(n4064), .ZN(n4065) );
  AOI21_X1 U4836 ( .B1(n4067), .B2(n4066), .A(n4065), .ZN(n4184) );
  OAI21_X1 U4837 ( .B1(n4113), .B2(n4115), .A(n4184), .ZN(n4069) );
  INV_X1 U4838 ( .A(n4246), .ZN(n4068) );
  AOI22_X1 U4839 ( .A1(n4070), .A2(n4069), .B1(n4068), .B2(n4252), .ZN(n4073)
         );
  NAND2_X1 U4840 ( .A1(n4198), .A2(n4071), .ZN(n4087) );
  AOI21_X1 U4841 ( .B1(n4087), .B2(n4246), .A(n4247), .ZN(n4072) );
  NOR2_X1 U4842 ( .A1(n4073), .A2(n4072), .ZN(n4189) );
  INV_X1 U4843 ( .A(n4074), .ZN(n4110) );
  NAND2_X1 U4844 ( .A1(n2403), .A2(n4076), .ZN(n4280) );
  NAND2_X1 U4845 ( .A1(n4078), .A2(n4077), .ZN(n4293) );
  NAND2_X1 U4846 ( .A1(n4291), .A2(n4079), .ZN(n4316) );
  INV_X1 U4847 ( .A(n4310), .ZN(n4168) );
  NAND2_X1 U4848 ( .A1(n4168), .A2(n4311), .ZN(n4347) );
  INV_X1 U4849 ( .A(n4448), .ZN(n4081) );
  NOR4_X1 U4850 ( .A1(n4081), .A2(n4131), .A3(n4080), .A4(n5029), .ZN(n4083)
         );
  NAND2_X1 U4851 ( .A1(n4364), .A2(n4366), .ZN(n4396) );
  INV_X1 U4852 ( .A(n4413), .ZN(n4408) );
  NAND4_X1 U4853 ( .A1(n4083), .A2(n4396), .A3(n4408), .A4(n4082), .ZN(n4106)
         );
  NAND2_X1 U4854 ( .A1(n4085), .A2(n4084), .ZN(n4374) );
  OR2_X1 U4855 ( .A1(n4369), .A2(n4370), .ZN(n4428) );
  INV_X1 U4856 ( .A(n4086), .ZN(n4093) );
  OAI21_X1 U4857 ( .B1(n4246), .B2(n4247), .A(n4087), .ZN(n4181) );
  OR4_X1 U4858 ( .A1(n4091), .A2(n4090), .A3(n4089), .A4(n4088), .ZN(n4092) );
  NOR4_X1 U4859 ( .A1(n4428), .A2(n4093), .A3(n4181), .A4(n4092), .ZN(n4104)
         );
  INV_X1 U4860 ( .A(n4094), .ZN(n4097) );
  NOR4_X1 U4861 ( .A1(n2470), .A2(n4097), .A3(n4096), .A4(n4095), .ZN(n4103)
         );
  NOR4_X1 U4862 ( .A1(n4101), .A2(n4100), .A3(n4099), .A4(n4098), .ZN(n4102)
         );
  NAND4_X1 U4863 ( .A1(n4374), .A2(n4104), .A3(n4103), .A4(n4102), .ZN(n4105)
         );
  OR4_X1 U4864 ( .A1(n4340), .A2(n4347), .A3(n4106), .A4(n4105), .ZN(n4107) );
  NOR4_X1 U4865 ( .A1(n4280), .A2(n4293), .A3(n4316), .A4(n4107), .ZN(n4109)
         );
  NAND4_X1 U4866 ( .A1(n4111), .A2(n4110), .A3(n4109), .A4(n4108), .ZN(n4114)
         );
  INV_X1 U4867 ( .A(n4948), .ZN(n4112) );
  OAI21_X1 U4868 ( .B1(n4114), .B2(n4113), .A(n4112), .ZN(n4186) );
  INV_X1 U4869 ( .A(n4115), .ZN(n4180) );
  OAI211_X1 U4870 ( .C1(n4118), .C2(n4948), .A(n4117), .B(n4116), .ZN(n4121)
         );
  NAND3_X1 U4871 ( .A1(n4121), .A2(n4120), .A3(n4119), .ZN(n4124) );
  NAND3_X1 U4872 ( .A1(n4124), .A2(n4123), .A3(n4122), .ZN(n4127) );
  NAND3_X1 U4873 ( .A1(n4127), .A2(n4126), .A3(n4125), .ZN(n4134) );
  NOR3_X1 U4874 ( .A1(n2203), .A2(n2208), .A3(n4129), .ZN(n4133) );
  INV_X1 U4875 ( .A(n4130), .ZN(n4132) );
  AOI211_X1 U4876 ( .C1(n4134), .C2(n4133), .A(n4132), .B(n4131), .ZN(n4139)
         );
  NAND2_X1 U4877 ( .A1(n4136), .A2(n4135), .ZN(n4145) );
  OAI211_X1 U4878 ( .C1(n4139), .C2(n4145), .A(n4138), .B(n4137), .ZN(n4142)
         );
  INV_X1 U4879 ( .A(n4140), .ZN(n4141) );
  NAND3_X1 U4880 ( .A1(n4142), .A2(n4141), .A3(n2847), .ZN(n4153) );
  NOR4_X1 U4881 ( .A1(n2203), .A2(n4145), .A3(n4144), .A4(n4143), .ZN(n4148)
         );
  INV_X1 U4882 ( .A(n4146), .ZN(n4147) );
  OAI21_X1 U4883 ( .B1(n4148), .B2(n4147), .A(n4158), .ZN(n4152) );
  NAND3_X1 U4884 ( .A1(n4156), .A2(n4150), .A3(n4149), .ZN(n4151) );
  AOI21_X1 U4885 ( .B1(n4153), .B2(n4152), .A(n4151), .ZN(n4164) );
  INV_X1 U4886 ( .A(n4154), .ZN(n4157) );
  AOI21_X1 U4887 ( .B1(n4157), .B2(n4156), .A(n4155), .ZN(n4161) );
  INV_X1 U4888 ( .A(n4158), .ZN(n4159) );
  AOI21_X1 U4889 ( .B1(n4161), .B2(n4160), .A(n4159), .ZN(n4163) );
  OAI21_X1 U4890 ( .B1(n4164), .B2(n4163), .A(n4162), .ZN(n4167) );
  AOI21_X1 U4891 ( .B1(n4167), .B2(n4166), .A(n4165), .ZN(n4170) );
  OAI211_X1 U4892 ( .C1(n4170), .C2(n2389), .A(n4169), .B(n4168), .ZN(n4171)
         );
  NAND4_X1 U4893 ( .A1(n4175), .A2(n4173), .A3(n4172), .A4(n4171), .ZN(n4178)
         );
  INV_X1 U4894 ( .A(n4174), .ZN(n4176) );
  NAND2_X1 U4895 ( .A1(n4176), .A2(n4175), .ZN(n4177) );
  NAND4_X1 U4896 ( .A1(n4180), .A2(n4179), .A3(n4178), .A4(n4177), .ZN(n4183)
         );
  AOI22_X1 U4897 ( .A1(n4184), .A2(n4183), .B1(n4182), .B2(n4181), .ZN(n4185)
         );
  MUX2_X1 U4898 ( .A(n4186), .B(n4185), .S(n2861), .Z(n4187) );
  OAI21_X1 U4899 ( .B1(n4189), .B2(n4188), .A(n4187), .ZN(n4191) );
  XNOR2_X1 U4900 ( .A(n4191), .B(n4190), .ZN(n4197) );
  NOR2_X1 U4901 ( .A1(n4193), .A2(n4192), .ZN(n4195) );
  OAI21_X1 U4902 ( .B1(n4196), .B2(n2946), .A(B_REG_SCAN_IN), .ZN(n4194) );
  OAI22_X1 U4903 ( .A1(n4197), .A2(n4196), .B1(n4195), .B2(n4194), .ZN(U3239)
         );
  MUX2_X1 U4904 ( .A(n4198), .B(DATAO_REG_30__SCAN_IN), .S(n4209), .Z(U3580)
         );
  MUX2_X1 U4905 ( .A(n4199), .B(DATAO_REG_29__SCAN_IN), .S(n4209), .Z(U3579)
         );
  MUX2_X1 U4906 ( .A(n4271), .B(DATAO_REG_28__SCAN_IN), .S(n4209), .Z(U3578)
         );
  MUX2_X1 U4907 ( .A(n4200), .B(DATAO_REG_27__SCAN_IN), .S(n4209), .Z(U3577)
         );
  MUX2_X1 U4908 ( .A(n4494), .B(DATAO_REG_24__SCAN_IN), .S(n4209), .Z(U3574)
         );
  MUX2_X1 U4909 ( .A(n4201), .B(DATAO_REG_23__SCAN_IN), .S(n4209), .Z(U3573)
         );
  MUX2_X1 U4910 ( .A(n4378), .B(DATAO_REG_21__SCAN_IN), .S(n4209), .Z(U3571)
         );
  MUX2_X1 U4911 ( .A(DATAO_REG_19__SCAN_IN), .B(n4527), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4912 ( .A(DATAO_REG_18__SCAN_IN), .B(n4438), .S(n4202), .Z(U3568)
         );
  MUX2_X1 U4913 ( .A(n4564), .B(DATAO_REG_16__SCAN_IN), .S(n4209), .Z(U3566)
         );
  MUX2_X1 U4914 ( .A(DATAO_REG_14__SCAN_IN), .B(n4203), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4915 ( .A(n4204), .B(DATAO_REG_12__SCAN_IN), .S(n4209), .Z(U3562)
         );
  MUX2_X1 U4916 ( .A(DATAO_REG_11__SCAN_IN), .B(n4591), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4917 ( .A(n4205), .B(DATAO_REG_8__SCAN_IN), .S(n4209), .Z(U3558) );
  MUX2_X1 U4918 ( .A(n4206), .B(DATAO_REG_7__SCAN_IN), .S(n4209), .Z(U3557) );
  MUX2_X1 U4919 ( .A(n4207), .B(DATAO_REG_5__SCAN_IN), .S(n4209), .Z(U3555) );
  MUX2_X1 U4920 ( .A(n2135), .B(DATAO_REG_2__SCAN_IN), .S(n4209), .Z(U3552) );
  MUX2_X1 U4921 ( .A(n4465), .B(DATAO_REG_1__SCAN_IN), .S(n4209), .Z(U3551) );
  MUX2_X1 U4922 ( .A(n2963), .B(DATAO_REG_0__SCAN_IN), .S(n4209), .Z(U3550) );
  INV_X1 U4923 ( .A(ADDR_REG_1__SCAN_IN), .ZN(n4856) );
  NOR2_X1 U4924 ( .A1(n5005), .A2(n4856), .ZN(n4212) );
  NOR2_X1 U4925 ( .A1(n5024), .A2(n4210), .ZN(n4211) );
  AOI211_X1 U4926 ( .C1(REG3_REG_1__SCAN_IN), .C2(U3149), .A(n4212), .B(n4211), 
        .ZN(n4221) );
  OAI211_X1 U4927 ( .C1(n4215), .C2(n4214), .A(n3215), .B(n4213), .ZN(n4220)
         );
  OAI211_X1 U4928 ( .C1(n3217), .C2(n4218), .A(n5001), .B(n4217), .ZN(n4219)
         );
  NAND3_X1 U4929 ( .A1(n4221), .A2(n4220), .A3(n4219), .ZN(U3241) );
  OAI211_X1 U4930 ( .C1(n4224), .C2(n4223), .A(n4222), .B(n3215), .ZN(n4233)
         );
  AOI21_X1 U4931 ( .B1(n5018), .B2(ADDR_REG_11__SCAN_IN), .A(n4225), .ZN(n4232) );
  OAI211_X1 U4932 ( .C1(n4228), .C2(n4227), .A(n4226), .B(n5001), .ZN(n4231)
         );
  INV_X1 U4933 ( .A(n4953), .ZN(n4229) );
  OR2_X1 U4934 ( .A1(n5024), .A2(n4229), .ZN(n4230) );
  NAND4_X1 U4935 ( .A1(n4233), .A2(n4232), .A3(n4231), .A4(n4230), .ZN(U3251)
         );
  XNOR2_X1 U4936 ( .A(n4234), .B(REG1_REG_14__SCAN_IN), .ZN(n4243) );
  AOI211_X1 U4937 ( .C1(n4237), .C2(n4236), .A(n5014), .B(n4235), .ZN(n4242)
         );
  NAND2_X1 U4938 ( .A1(n5018), .A2(ADDR_REG_14__SCAN_IN), .ZN(n4238) );
  OAI211_X1 U4939 ( .C1(n5024), .C2(n4240), .A(n4239), .B(n4238), .ZN(n4241)
         );
  AOI211_X1 U4940 ( .C1(n4243), .C2(n3215), .A(n4242), .B(n4241), .ZN(n4244)
         );
  INV_X1 U4941 ( .A(n4244), .ZN(U3254) );
  NOR2_X2 U4942 ( .A1(n4251), .A2(n4252), .ZN(n4250) );
  XNOR2_X1 U4943 ( .A(n4250), .B(n4247), .ZN(n4881) );
  NAND2_X1 U4944 ( .A1(n4246), .A2(n4245), .ZN(n4254) );
  OAI21_X1 U4945 ( .B1(n4247), .B2(n4593), .A(n4254), .ZN(n4878) );
  NAND2_X1 U4946 ( .A1(n5032), .A2(n4878), .ZN(n4249) );
  NAND2_X1 U4947 ( .A1(n4462), .A2(REG2_REG_31__SCAN_IN), .ZN(n4248) );
  OAI211_X1 U4948 ( .C1(n4881), .C2(n4458), .A(n4249), .B(n4248), .ZN(U3260)
         );
  AOI21_X1 U4949 ( .B1(n4252), .B2(n4251), .A(n4250), .ZN(n4882) );
  NAND2_X1 U4950 ( .A1(n4882), .A2(n4473), .ZN(n4256) );
  NAND2_X1 U4951 ( .A1(n4252), .A2(n4570), .ZN(n4253) );
  NAND2_X1 U4952 ( .A1(n4254), .A2(n4253), .ZN(n4883) );
  NAND2_X1 U4953 ( .A1(n5032), .A2(n4883), .ZN(n4255) );
  OAI211_X1 U4954 ( .C1(n5032), .C2(n4819), .A(n4256), .B(n4255), .ZN(U3261)
         );
  XNOR2_X1 U4955 ( .A(n4257), .B(n4258), .ZN(n4487) );
  NOR2_X1 U4956 ( .A1(n4259), .A2(n4258), .ZN(n4260) );
  OR2_X1 U4957 ( .A1(n4261), .A2(n4260), .ZN(n4262) );
  NAND2_X1 U4958 ( .A1(n4262), .A2(n4577), .ZN(n4485) );
  NOR2_X1 U4959 ( .A1(n4485), .A2(n4337), .ZN(n4274) );
  AND2_X1 U4960 ( .A1(n4263), .A2(n4482), .ZN(n4265) );
  OR2_X1 U4961 ( .A1(n4265), .A2(n4264), .ZN(n4890) );
  NAND2_X1 U4962 ( .A1(n4483), .A2(n4466), .ZN(n4269) );
  AOI22_X1 U4963 ( .A1(n4467), .A2(n4482), .B1(n4462), .B2(
        REG2_REG_27__SCAN_IN), .ZN(n4268) );
  NAND2_X1 U4964 ( .A1(n4266), .A2(n5028), .ZN(n4267) );
  NAND3_X1 U4965 ( .A1(n4269), .A2(n4268), .A3(n4267), .ZN(n4270) );
  AOI21_X1 U4966 ( .B1(n4271), .B2(n4471), .A(n4270), .ZN(n4272) );
  OAI21_X1 U4967 ( .B1(n4890), .B2(n4458), .A(n4272), .ZN(n4273) );
  AOI211_X1 U4968 ( .C1(n4487), .C2(n4460), .A(n4274), .B(n4273), .ZN(n4275)
         );
  INV_X1 U4969 ( .A(n4275), .ZN(U3263) );
  XNOR2_X1 U4970 ( .A(n4276), .B(n4280), .ZN(n4277) );
  NAND2_X1 U4971 ( .A1(n4277), .A2(n4577), .ZN(n4496) );
  XNOR2_X1 U4972 ( .A(n4279), .B(n4280), .ZN(n4499) );
  NAND2_X1 U4973 ( .A1(n4499), .A2(n4460), .ZN(n4289) );
  OAI22_X1 U4974 ( .A1(n4282), .A2(n4451), .B1(n4281), .B2(n5032), .ZN(n4283)
         );
  AOI21_X1 U4975 ( .B1(n4493), .B2(n4467), .A(n4283), .ZN(n4284) );
  OAI21_X1 U4976 ( .B1(n4314), .B2(n4434), .A(n4284), .ZN(n4287) );
  OAI21_X1 U4977 ( .B1(n4301), .B2(n4285), .A(n3815), .ZN(n4899) );
  NOR2_X1 U4978 ( .A1(n4899), .A2(n4458), .ZN(n4286) );
  AOI211_X1 U4979 ( .C1(n4471), .C2(n4483), .A(n4287), .B(n4286), .ZN(n4288)
         );
  OAI211_X1 U4980 ( .C1(n4462), .C2(n4496), .A(n4289), .B(n4288), .ZN(U3265)
         );
  XNOR2_X1 U4981 ( .A(n4290), .B(n4293), .ZN(n4503) );
  INV_X1 U4982 ( .A(n4503), .ZN(n4309) );
  NAND2_X1 U4983 ( .A1(n4292), .A2(n4291), .ZN(n4295) );
  INV_X1 U4984 ( .A(n4293), .ZN(n4294) );
  XNOR2_X1 U4985 ( .A(n4295), .B(n4294), .ZN(n4296) );
  NAND2_X1 U4986 ( .A1(n4296), .A2(n4577), .ZN(n4300) );
  OAI22_X1 U4987 ( .A1(n4333), .A2(n4561), .B1(n4303), .B2(n4593), .ZN(n4297)
         );
  AOI21_X1 U4988 ( .B1(n4589), .B2(n4298), .A(n4297), .ZN(n4299) );
  NAND2_X1 U4989 ( .A1(n4300), .A2(n4299), .ZN(n4502) );
  INV_X1 U4990 ( .A(n4319), .ZN(n4304) );
  INV_X1 U4991 ( .A(n4301), .ZN(n4302) );
  OAI21_X1 U4992 ( .B1(n4304), .B2(n4303), .A(n4302), .ZN(n4903) );
  AOI22_X1 U4993 ( .A1(n4305), .A2(n5028), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4337), .ZN(n4306) );
  OAI21_X1 U4994 ( .B1(n4903), .B2(n4458), .A(n4306), .ZN(n4307) );
  AOI21_X1 U4995 ( .B1(n4502), .B2(n5032), .A(n4307), .ZN(n4308) );
  OAI21_X1 U4996 ( .B1(n4309), .B2(n4423), .A(n4308), .ZN(U3266) );
  INV_X1 U4997 ( .A(n4311), .ZN(n4326) );
  INV_X1 U4998 ( .A(n4340), .ZN(n4327) );
  OAI21_X1 U4999 ( .B1(n4328), .B2(n4326), .A(n4327), .ZN(n4325) );
  AOI22_X1 U5000 ( .A1(n4356), .A2(n4590), .B1(n4570), .B2(n4317), .ZN(n4313)
         );
  INV_X1 U5001 ( .A(n4506), .ZN(n4324) );
  XOR2_X1 U5002 ( .A(n4316), .B(n4315), .Z(n4507) );
  NAND2_X1 U5003 ( .A1(n4336), .A2(n4317), .ZN(n4318) );
  NAND2_X1 U5004 ( .A1(n4319), .A2(n4318), .ZN(n4907) );
  AOI22_X1 U5005 ( .A1(n4320), .A2(n5028), .B1(REG2_REG_23__SCAN_IN), .B2(
        n4337), .ZN(n4321) );
  OAI21_X1 U5006 ( .B1(n4907), .B2(n4458), .A(n4321), .ZN(n4322) );
  AOI21_X1 U5007 ( .B1(n4507), .B2(n4460), .A(n4322), .ZN(n4323) );
  OAI21_X1 U5008 ( .B1(n4462), .B2(n4324), .A(n4323), .ZN(U3267) );
  INV_X1 U5009 ( .A(n4325), .ZN(n4330) );
  NOR3_X1 U5010 ( .A1(n4328), .A2(n4327), .A3(n4326), .ZN(n4329) );
  OAI21_X1 U5011 ( .B1(n4330), .B2(n4329), .A(n4577), .ZN(n4332) );
  AOI22_X1 U5012 ( .A1(n4378), .A2(n4590), .B1(n4334), .B2(n4570), .ZN(n4331)
         );
  OAI211_X1 U5013 ( .C1(n4333), .C2(n4573), .A(n4332), .B(n4331), .ZN(n4511)
         );
  NAND2_X1 U5014 ( .A1(n4352), .A2(n4334), .ZN(n4335) );
  NAND2_X1 U5015 ( .A1(n4336), .A2(n4335), .ZN(n4911) );
  AOI22_X1 U5016 ( .A1(n4338), .A2(n5028), .B1(REG2_REG_22__SCAN_IN), .B2(
        n4337), .ZN(n4339) );
  OAI21_X1 U5017 ( .B1(n4911), .B2(n4458), .A(n4339), .ZN(n4344) );
  NOR2_X1 U5018 ( .A1(n4341), .A2(n4340), .ZN(n4510) );
  INV_X1 U5019 ( .A(n4512), .ZN(n4342) );
  NOR3_X1 U5020 ( .A1(n4510), .A2(n4342), .A3(n4423), .ZN(n4343) );
  AOI211_X1 U5021 ( .C1(n5032), .C2(n4511), .A(n4344), .B(n4343), .ZN(n4345)
         );
  INV_X1 U5022 ( .A(n4345), .ZN(U3268) );
  XNOR2_X1 U5023 ( .A(n4346), .B(n4347), .ZN(n4522) );
  XNOR2_X1 U5024 ( .A(n4348), .B(n4347), .ZN(n4349) );
  NAND2_X1 U5025 ( .A1(n4349), .A2(n4577), .ZN(n4519) );
  NOR2_X1 U5026 ( .A1(n4519), .A2(n4337), .ZN(n4360) );
  OR2_X1 U5027 ( .A1(n4377), .A2(n4350), .ZN(n4351) );
  NAND2_X1 U5028 ( .A1(n4352), .A2(n4351), .ZN(n4914) );
  INV_X1 U5029 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4353) );
  OAI22_X1 U5030 ( .A1(n4354), .A2(n4451), .B1(n4353), .B2(n5032), .ZN(n4355)
         );
  AOI21_X1 U5031 ( .B1(n4356), .B2(n4471), .A(n4355), .ZN(n4358) );
  AOI22_X1 U5032 ( .A1(n4517), .A2(n4466), .B1(n4467), .B2(n4516), .ZN(n4357)
         );
  OAI211_X1 U5033 ( .C1(n4914), .C2(n4458), .A(n4358), .B(n4357), .ZN(n4359)
         );
  AOI211_X1 U5034 ( .C1(n4522), .C2(n4460), .A(n4360), .B(n4359), .ZN(n4361)
         );
  INV_X1 U5035 ( .A(n4361), .ZN(U3269) );
  NAND2_X1 U5036 ( .A1(n4362), .A2(n4413), .ZN(n4406) );
  NAND2_X1 U5037 ( .A1(n4406), .A2(n4363), .ZN(n4395) );
  INV_X1 U5038 ( .A(n4364), .ZN(n4365) );
  AOI21_X1 U5039 ( .B1(n4395), .B2(n4366), .A(n4365), .ZN(n4367) );
  XNOR2_X1 U5040 ( .A(n4367), .B(n4374), .ZN(n4532) );
  INV_X1 U5041 ( .A(n4532), .ZN(n4387) );
  INV_X1 U5042 ( .A(n4368), .ZN(n4424) );
  INV_X1 U5043 ( .A(n4369), .ZN(n4371) );
  AOI21_X1 U5044 ( .B1(n4424), .B2(n4371), .A(n4370), .ZN(n4414) );
  OAI21_X1 U5045 ( .B1(n4414), .B2(n4373), .A(n4372), .ZN(n4375) );
  XNOR2_X1 U5046 ( .A(n4375), .B(n4374), .ZN(n4525) );
  NOR2_X1 U5047 ( .A1(n4397), .A2(n4382), .ZN(n4376) );
  OR2_X1 U5048 ( .A1(n4377), .A2(n4376), .ZN(n4918) );
  NOR2_X1 U5049 ( .A1(n4918), .A2(n4458), .ZN(n4384) );
  AOI22_X1 U5050 ( .A1(n4378), .A2(n4471), .B1(n4466), .B2(n4527), .ZN(n4381)
         );
  AOI22_X1 U5051 ( .A1(n4379), .A2(n5028), .B1(n4462), .B2(
        REG2_REG_20__SCAN_IN), .ZN(n4380) );
  OAI211_X1 U5052 ( .C1(n4382), .C2(n4433), .A(n4381), .B(n4380), .ZN(n4383)
         );
  AOI211_X1 U5053 ( .C1(n4525), .C2(n4385), .A(n4384), .B(n4383), .ZN(n4386)
         );
  OAI21_X1 U5054 ( .B1(n4387), .B2(n4423), .A(n4386), .ZN(U3270) );
  INV_X1 U5055 ( .A(n4388), .ZN(n4389) );
  AOI21_X1 U5056 ( .B1(n4414), .B2(n4390), .A(n4389), .ZN(n4391) );
  XOR2_X1 U5057 ( .A(n4396), .B(n4391), .Z(n4394) );
  OAI22_X1 U5058 ( .A1(n4543), .A2(n4561), .B1(n4399), .B2(n4593), .ZN(n4392)
         );
  AOI21_X1 U5059 ( .B1(n4517), .B2(n4589), .A(n4392), .ZN(n4393) );
  OAI21_X1 U5060 ( .B1(n4394), .B2(n4425), .A(n4393), .ZN(n4534) );
  INV_X1 U5061 ( .A(n4534), .ZN(n4405) );
  XOR2_X1 U5062 ( .A(n4396), .B(n4395), .Z(n4535) );
  INV_X1 U5063 ( .A(n4410), .ZN(n4400) );
  INV_X1 U5064 ( .A(n4397), .ZN(n4398) );
  OAI21_X1 U5065 ( .B1(n4400), .B2(n4399), .A(n4398), .ZN(n4922) );
  AOI22_X1 U5066 ( .A1(n4337), .A2(REG2_REG_19__SCAN_IN), .B1(n4401), .B2(
        n5028), .ZN(n4402) );
  OAI21_X1 U5067 ( .B1(n4922), .B2(n4458), .A(n4402), .ZN(n4403) );
  AOI21_X1 U5068 ( .B1(n4535), .B2(n4460), .A(n4403), .ZN(n4404) );
  OAI21_X1 U5069 ( .B1(n4462), .B2(n4405), .A(n4404), .ZN(U3271) );
  INV_X1 U5070 ( .A(n4406), .ZN(n4407) );
  AOI21_X1 U5071 ( .B1(n4408), .B2(n2452), .A(n4407), .ZN(n4540) );
  AOI22_X1 U5072 ( .A1(n4462), .A2(REG2_REG_18__SCAN_IN), .B1(n4409), .B2(
        n5028), .ZN(n4422) );
  INV_X1 U5073 ( .A(n4429), .ZN(n4412) );
  OAI211_X1 U5074 ( .C1(n4412), .C2(n4411), .A(n4410), .B(n2941), .ZN(n4538)
         );
  XNOR2_X1 U5075 ( .A(n4414), .B(n4413), .ZN(n4419) );
  AOI22_X1 U5076 ( .A1(n4555), .A2(n4590), .B1(n4570), .B2(n4415), .ZN(n4416)
         );
  OAI21_X1 U5077 ( .B1(n4417), .B2(n4573), .A(n4416), .ZN(n4418) );
  AOI21_X1 U5078 ( .B1(n4419), .B2(n4577), .A(n4418), .ZN(n4539) );
  OAI21_X1 U5079 ( .B1(n4950), .B2(n4538), .A(n4539), .ZN(n4420) );
  NAND2_X1 U5080 ( .A1(n4420), .A2(n5032), .ZN(n4421) );
  OAI211_X1 U5081 ( .C1(n4540), .C2(n4423), .A(n4422), .B(n4421), .ZN(U3272)
         );
  XNOR2_X1 U5082 ( .A(n4424), .B(n4428), .ZN(n4426) );
  NOR2_X1 U5083 ( .A1(n4426), .A2(n4425), .ZN(n4544) );
  INV_X1 U5084 ( .A(n4544), .ZN(n4442) );
  XNOR2_X1 U5085 ( .A(n4427), .B(n4428), .ZN(n4546) );
  OAI21_X1 U5086 ( .B1(n4450), .B2(n4432), .A(n4429), .ZN(n4927) );
  OAI22_X1 U5087 ( .A1(n5032), .A2(n4431), .B1(n4430), .B2(n4451), .ZN(n4437)
         );
  OAI22_X1 U5088 ( .A1(n4435), .A2(n4434), .B1(n4433), .B2(n4432), .ZN(n4436)
         );
  AOI211_X1 U5089 ( .C1(n4471), .C2(n4438), .A(n4437), .B(n4436), .ZN(n4439)
         );
  OAI21_X1 U5090 ( .B1(n4927), .B2(n4458), .A(n4439), .ZN(n4440) );
  AOI21_X1 U5091 ( .B1(n4546), .B2(n4460), .A(n4440), .ZN(n4441) );
  OAI21_X1 U5092 ( .B1(n4462), .B2(n4442), .A(n4441), .ZN(U3273) );
  OAI211_X1 U5093 ( .C1(n4444), .C2(n4448), .A(n4443), .B(n4577), .ZN(n4556)
         );
  INV_X1 U5094 ( .A(n4445), .ZN(n4446) );
  AOI21_X1 U5095 ( .B1(n4448), .B2(n4447), .A(n4446), .ZN(n4549) );
  NOR2_X1 U5096 ( .A1(n3786), .A2(n4550), .ZN(n4449) );
  OR2_X1 U5097 ( .A1(n4450), .A2(n4449), .ZN(n4552) );
  OAI22_X1 U5098 ( .A1(n5032), .A2(n4992), .B1(n4452), .B2(n4451), .ZN(n4453)
         );
  AOI21_X1 U5099 ( .B1(n4471), .B2(n4555), .A(n4453), .ZN(n4457) );
  AOI22_X1 U5100 ( .A1(n4455), .A2(n4467), .B1(n4466), .B2(n4454), .ZN(n4456)
         );
  OAI211_X1 U5101 ( .C1(n4552), .C2(n4458), .A(n4457), .B(n4456), .ZN(n4459)
         );
  AOI21_X1 U5102 ( .B1(n4549), .B2(n4460), .A(n4459), .ZN(n4461) );
  OAI21_X1 U5103 ( .B1(n4462), .B2(n4556), .A(n4461), .ZN(U3274) );
  MUX2_X1 U5104 ( .A(n4464), .B(n4463), .S(n5032), .Z(n4477) );
  AOI22_X1 U5105 ( .A1(n4468), .A2(n4467), .B1(n4466), .B2(n4465), .ZN(n4476)
         );
  AOI22_X1 U5106 ( .A1(n5030), .A2(n4469), .B1(REG3_REG_2__SCAN_IN), .B2(n5028), .ZN(n4475) );
  INV_X1 U5107 ( .A(n4872), .ZN(n4472) );
  AOI22_X1 U5108 ( .A1(n4473), .A2(n4472), .B1(n4471), .B2(n4470), .ZN(n4474)
         );
  NAND4_X1 U5109 ( .A1(n4477), .A2(n4476), .A3(n4475), .A4(n4474), .ZN(U3288)
         );
  NAND2_X1 U5110 ( .A1(n5081), .A2(n4878), .ZN(n4479) );
  NAND2_X1 U5111 ( .A1(n5079), .A2(REG1_REG_31__SCAN_IN), .ZN(n4478) );
  OAI211_X1 U5112 ( .C1(n4881), .C2(n4873), .A(n4479), .B(n4478), .ZN(U3549)
         );
  NAND2_X1 U5113 ( .A1(n4882), .A2(n4582), .ZN(n4481) );
  NAND2_X1 U5114 ( .A1(n5081), .A2(n4883), .ZN(n4480) );
  OAI211_X1 U5115 ( .C1(n5081), .C2(n4656), .A(n4481), .B(n4480), .ZN(U3548)
         );
  INV_X1 U5116 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4488) );
  AOI22_X1 U5117 ( .A1(n4483), .A2(n4590), .B1(n4482), .B2(n4570), .ZN(n4484)
         );
  OAI21_X1 U5118 ( .B1(n4490), .B2(n5069), .A(n4489), .ZN(n4891) );
  MUX2_X1 U5119 ( .A(REG1_REG_26__SCAN_IN), .B(n4891), .S(n5081), .Z(n4491) );
  INV_X1 U5120 ( .A(n4491), .ZN(n4492) );
  OAI21_X1 U5121 ( .B1(n4873), .B2(n4895), .A(n4492), .ZN(U3544) );
  INV_X1 U5122 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4500) );
  AOI22_X1 U5123 ( .A1(n4494), .A2(n4590), .B1(n4493), .B2(n4570), .ZN(n4495)
         );
  OAI211_X1 U5124 ( .C1(n4497), .C2(n4573), .A(n4496), .B(n4495), .ZN(n4498)
         );
  AOI21_X1 U5125 ( .B1(n4499), .B2(n4598), .A(n4498), .ZN(n4896) );
  MUX2_X1 U5126 ( .A(n4500), .B(n4896), .S(n5081), .Z(n4501) );
  OAI21_X1 U5127 ( .B1(n4873), .B2(n4899), .A(n4501), .ZN(U3543) );
  INV_X1 U5128 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4504) );
  AOI21_X1 U5129 ( .B1(n4503), .B2(n4598), .A(n4502), .ZN(n4900) );
  MUX2_X1 U5130 ( .A(n4504), .B(n4900), .S(n5081), .Z(n4505) );
  OAI21_X1 U5131 ( .B1(n4873), .B2(n4903), .A(n4505), .ZN(U3542) );
  INV_X1 U5132 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4508) );
  AOI21_X1 U5133 ( .B1(n4507), .B2(n4598), .A(n4506), .ZN(n4904) );
  MUX2_X1 U5134 ( .A(n4508), .B(n4904), .S(n5081), .Z(n4509) );
  OAI21_X1 U5135 ( .B1(n4873), .B2(n4907), .A(n4509), .ZN(U3541) );
  INV_X1 U5136 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4514) );
  NOR2_X1 U5137 ( .A1(n4510), .A2(n5069), .ZN(n4513) );
  AOI21_X1 U5138 ( .B1(n4513), .B2(n4512), .A(n4511), .ZN(n4908) );
  MUX2_X1 U5139 ( .A(n4514), .B(n4908), .S(n5081), .Z(n4515) );
  OAI21_X1 U5140 ( .B1(n4873), .B2(n4911), .A(n4515), .ZN(U3540) );
  AOI22_X1 U5141 ( .A1(n4517), .A2(n4590), .B1(n4570), .B2(n4516), .ZN(n4518)
         );
  OAI211_X1 U5142 ( .C1(n4520), .C2(n4573), .A(n4519), .B(n4518), .ZN(n4521)
         );
  AOI21_X1 U5143 ( .B1(n4522), .B2(n4598), .A(n4521), .ZN(n4912) );
  MUX2_X1 U5144 ( .A(n4523), .B(n4912), .S(n5081), .Z(n4524) );
  OAI21_X1 U5145 ( .B1(n4873), .B2(n4914), .A(n4524), .ZN(U3539) );
  NAND2_X1 U5146 ( .A1(n4525), .A2(n4577), .ZN(n4529) );
  AOI22_X1 U5147 ( .A1(n4527), .A2(n4590), .B1(n4526), .B2(n4570), .ZN(n4528)
         );
  OAI211_X1 U5148 ( .C1(n4530), .C2(n4573), .A(n4529), .B(n4528), .ZN(n4531)
         );
  AOI21_X1 U5149 ( .B1(n4532), .B2(n4598), .A(n4531), .ZN(n4915) );
  MUX2_X1 U5150 ( .A(n4783), .B(n4915), .S(n5081), .Z(n4533) );
  OAI21_X1 U5151 ( .B1(n4873), .B2(n4918), .A(n4533), .ZN(U3538) );
  AOI21_X1 U5152 ( .B1(n4535), .B2(n4598), .A(n4534), .ZN(n4919) );
  MUX2_X1 U5153 ( .A(n4536), .B(n4919), .S(n5081), .Z(n4537) );
  OAI21_X1 U5154 ( .B1(n4873), .B2(n4922), .A(n4537), .ZN(U3537) );
  OAI211_X1 U5155 ( .C1(n4540), .C2(n5069), .A(n4539), .B(n4538), .ZN(n4923)
         );
  MUX2_X1 U5156 ( .A(REG1_REG_18__SCAN_IN), .B(n4923), .S(n5081), .Z(U3536) );
  AOI22_X1 U5157 ( .A1(n4564), .A2(n4590), .B1(n4570), .B2(n4541), .ZN(n4542)
         );
  OAI21_X1 U5158 ( .B1(n4543), .B2(n4573), .A(n4542), .ZN(n4545) );
  AOI211_X1 U5159 ( .C1(n4546), .C2(n4598), .A(n4545), .B(n4544), .ZN(n4924)
         );
  MUX2_X1 U5160 ( .A(n4547), .B(n4924), .S(n5081), .Z(n4548) );
  OAI21_X1 U5161 ( .B1(n4873), .B2(n4927), .A(n4548), .ZN(U3535) );
  INV_X1 U5162 ( .A(n4549), .ZN(n4558) );
  OAI22_X1 U5163 ( .A1(n4574), .A2(n4561), .B1(n4550), .B2(n4593), .ZN(n4554)
         );
  NOR2_X1 U5164 ( .A1(n4552), .A2(n4551), .ZN(n4553) );
  AOI211_X1 U5165 ( .C1(n4589), .C2(n4555), .A(n4554), .B(n4553), .ZN(n4557)
         );
  OAI211_X1 U5166 ( .C1(n4558), .C2(n5069), .A(n4557), .B(n4556), .ZN(n4928)
         );
  MUX2_X1 U5167 ( .A(REG1_REG_16__SCAN_IN), .B(n4928), .S(n5081), .Z(U3534) );
  NAND2_X1 U5168 ( .A1(n4559), .A2(n4598), .ZN(n4567) );
  OAI22_X1 U5169 ( .A1(n4562), .A2(n4561), .B1(n4593), .B2(n4560), .ZN(n4563)
         );
  AOI21_X1 U5170 ( .B1(n4564), .B2(n4589), .A(n4563), .ZN(n4566) );
  NAND3_X1 U5171 ( .A1(n4567), .A2(n4566), .A3(n4565), .ZN(n4929) );
  MUX2_X1 U5172 ( .A(REG1_REG_15__SCAN_IN), .B(n4929), .S(n5081), .Z(n4568) );
  AOI21_X1 U5173 ( .B1(n4582), .B2(n4931), .A(n4568), .ZN(n4569) );
  INV_X1 U5174 ( .A(n4569), .ZN(U3533) );
  AOI22_X1 U5175 ( .A1(n4590), .A2(n4588), .B1(n4571), .B2(n4570), .ZN(n4572)
         );
  OAI21_X1 U5176 ( .B1(n4574), .B2(n4573), .A(n4572), .ZN(n4575) );
  AOI21_X1 U5177 ( .B1(n4576), .B2(n4598), .A(n4575), .ZN(n4580) );
  NAND2_X1 U5178 ( .A1(n4578), .A2(n4577), .ZN(n4579) );
  NAND2_X1 U5179 ( .A1(n4580), .A2(n4579), .ZN(n4933) );
  MUX2_X1 U5180 ( .A(REG1_REG_14__SCAN_IN), .B(n4933), .S(n5081), .Z(n4581) );
  AOI21_X1 U5181 ( .B1(n4582), .B2(n4936), .A(n4581), .ZN(n4583) );
  INV_X1 U5182 ( .A(n4583), .ZN(U3532) );
  AOI21_X1 U5183 ( .B1(n4598), .B2(n4585), .A(n4584), .ZN(n4938) );
  MUX2_X1 U5184 ( .A(n4586), .B(n4938), .S(n5081), .Z(n4587) );
  OAI21_X1 U5185 ( .B1(n4873), .B2(n4941), .A(n4587), .ZN(U3531) );
  AOI22_X1 U5186 ( .A1(n4591), .A2(n4590), .B1(n4589), .B2(n4588), .ZN(n4592)
         );
  OAI21_X1 U5187 ( .B1(n4594), .B2(n4593), .A(n4592), .ZN(n4596) );
  AOI211_X1 U5188 ( .C1(n4598), .C2(n4597), .A(n4596), .B(n4595), .ZN(n4942)
         );
  MUX2_X1 U5189 ( .A(n4599), .B(n4942), .S(n5081), .Z(n4600) );
  OAI21_X1 U5190 ( .B1(n4873), .B2(n4946), .A(n4600), .ZN(U3530) );
  NAND4_X1 U5191 ( .A1(REG1_REG_17__SCAN_IN), .A2(REG1_REG_13__SCAN_IN), .A3(
        ADDR_REG_17__SCAN_IN), .A4(n4842), .ZN(n4607) );
  INV_X1 U5192 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n5004) );
  NAND4_X1 U5193 ( .A1(REG2_REG_12__SCAN_IN), .A2(REG3_REG_14__SCAN_IN), .A3(
        ADDR_REG_12__SCAN_IN), .A4(n5004), .ZN(n4606) );
  INV_X1 U5194 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4818) );
  NOR4_X1 U5195 ( .A1(REG3_REG_22__SCAN_IN), .A2(n4812), .A3(n4818), .A4(n4819), .ZN(n4604) );
  NOR4_X1 U5196 ( .A1(REG2_REG_29__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .A3(
        REG3_REG_24__SCAN_IN), .A4(n4831), .ZN(n4603) );
  INV_X1 U5197 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4850) );
  NOR4_X1 U5198 ( .A1(REG2_REG_10__SCAN_IN), .A2(ADDR_REG_9__SCAN_IN), .A3(
        ADDR_REG_11__SCAN_IN), .A4(n4850), .ZN(n4602) );
  NOR4_X1 U5199 ( .A1(DATAI_20_), .A2(REG2_REG_20__SCAN_IN), .A3(n4815), .A4(
        n4856), .ZN(n4601) );
  NAND4_X1 U5200 ( .A1(n4604), .A2(n4603), .A3(n4602), .A4(n4601), .ZN(n4605)
         );
  NOR3_X1 U5201 ( .A1(n4607), .A2(n4606), .A3(n4605), .ZN(n4648) );
  INV_X1 U5202 ( .A(IR_REG_18__SCAN_IN), .ZN(n4678) );
  NOR4_X1 U5203 ( .A1(IR_REG_21__SCAN_IN), .A2(DATAO_REG_6__SCAN_IN), .A3(
        n4678), .A4(n4608), .ZN(n4647) );
  INV_X1 U5204 ( .A(DATAI_11_), .ZN(n4711) );
  NAND4_X1 U5205 ( .A1(DATAO_REG_25__SCAN_IN), .A2(DATAO_REG_17__SCAN_IN), 
        .A3(DATAO_REG_20__SCAN_IN), .A4(n4711), .ZN(n4616) );
  NOR4_X1 U5206 ( .A1(REG2_REG_19__SCAN_IN), .A2(REG1_REG_18__SCAN_IN), .A3(
        n4536), .A4(n4431), .ZN(n4610) );
  NOR4_X1 U5207 ( .A1(REG2_REG_11__SCAN_IN), .A2(REG1_REG_7__SCAN_IN), .A3(
        REG1_REG_5__SCAN_IN), .A4(REG2_REG_5__SCAN_IN), .ZN(n4609) );
  AND3_X1 U5208 ( .A1(n2507), .A2(n4610), .A3(n4609), .ZN(n4611) );
  AND3_X1 U5209 ( .A1(IR_REG_26__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(n4611), 
        .ZN(n4613) );
  NOR2_X1 U5210 ( .A1(REG3_REG_6__SCAN_IN), .A2(DATAI_22_), .ZN(n4612) );
  NAND4_X1 U5211 ( .A1(n4613), .A2(IR_REG_22__SCAN_IN), .A3(IR_REG_27__SCAN_IN), .A4(n4612), .ZN(n4615) );
  INV_X1 U5212 ( .A(B_REG_SCAN_IN), .ZN(n4809) );
  NAND4_X1 U5213 ( .A1(D_REG_1__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(n4809), .ZN(n4614) );
  NOR3_X1 U5214 ( .A1(n4616), .A2(n4615), .A3(n4614), .ZN(n4633) );
  NAND4_X1 U5215 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .A3(
        IR_REG_4__SCAN_IN), .A4(n2614), .ZN(n4619) );
  NAND4_X1 U5216 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n4617) );
  NOR3_X1 U5217 ( .A1(n4619), .A2(n4618), .A3(n4617), .ZN(n4632) );
  INV_X1 U5218 ( .A(DATAI_8_), .ZN(n4620) );
  INV_X1 U5219 ( .A(DATAI_12_), .ZN(n4692) );
  NAND4_X1 U5220 ( .A1(n4705), .A2(n4621), .A3(n4620), .A4(n4692), .ZN(n4625)
         );
  INV_X1 U5221 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4622) );
  NAND4_X1 U5222 ( .A1(n4623), .A2(n4622), .A3(REG1_REG_0__SCAN_IN), .A4(
        DATAI_31_), .ZN(n4624) );
  NOR3_X1 U5223 ( .A1(n4744), .A2(n4625), .A3(n4624), .ZN(n4631) );
  INV_X1 U5224 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n4712) );
  NAND4_X1 U5225 ( .A1(ADDR_REG_0__SCAN_IN), .A2(REG3_REG_16__SCAN_IN), .A3(
        DATAO_REG_26__SCAN_IN), .A4(n4712), .ZN(n4629) );
  NAND4_X1 U5226 ( .A1(DATAI_23_), .A2(REG0_REG_31__SCAN_IN), .A3(
        DATAO_REG_9__SCAN_IN), .A4(DATAO_REG_15__SCAN_IN), .ZN(n4628) );
  INV_X1 U5227 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n4626) );
  NAND4_X1 U5228 ( .A1(n4626), .A2(n4745), .A3(DATAO_REG_31__SCAN_IN), .A4(
        DATAO_REG_22__SCAN_IN), .ZN(n4627) );
  NOR3_X1 U5229 ( .A1(n4629), .A2(n4628), .A3(n4627), .ZN(n4630) );
  AND4_X1 U5230 ( .A1(n4633), .A2(n4632), .A3(n4631), .A4(n4630), .ZN(n4637)
         );
  INV_X1 U5231 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4773) );
  NOR4_X1 U5232 ( .A1(REG1_REG_14__SCAN_IN), .A2(REG0_REG_13__SCAN_IN), .A3(
        n4773), .A4(n4761), .ZN(n4636) );
  INV_X1 U5233 ( .A(DATAI_24_), .ZN(n4668) );
  INV_X1 U5234 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n4677) );
  NOR4_X1 U5235 ( .A1(DATAI_17_), .A2(n5051), .A3(n4668), .A4(n4677), .ZN(
        n4635) );
  NOR4_X1 U5236 ( .A1(DATAO_REG_3__SCAN_IN), .A2(DATAO_REG_10__SCAN_IN), .A3(
        n2724), .A4(n4658), .ZN(n4634) );
  AND4_X1 U5237 ( .A1(n4637), .A2(n4636), .A3(n4635), .A4(n4634), .ZN(n4646)
         );
  NAND4_X1 U5238 ( .A1(DATAI_9_), .A2(REG0_REG_8__SCAN_IN), .A3(
        REG0_REG_6__SCAN_IN), .A4(n4796), .ZN(n4644) );
  NAND4_X1 U5239 ( .A1(DATAI_13_), .A2(REG3_REG_13__SCAN_IN), .A3(
        REG1_REG_10__SCAN_IN), .A4(n4765), .ZN(n4643) );
  NOR4_X1 U5240 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG1_REG_21__SCAN_IN), .A3(
        REG0_REG_21__SCAN_IN), .A4(n4353), .ZN(n4641) );
  INV_X1 U5241 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4794) );
  NOR4_X1 U5242 ( .A1(REG0_REG_17__SCAN_IN), .A2(n4783), .A3(n4784), .A4(n4794), .ZN(n4640) );
  NOR4_X1 U5243 ( .A1(REG0_REG_29__SCAN_IN), .A2(REG1_REG_28__SCAN_IN), .A3(
        n3266), .A4(n4656), .ZN(n4639) );
  NOR4_X1 U5244 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG0_REG_27__SCAN_IN), .A3(
        REG0_REG_26__SCAN_IN), .A4(REG0_REG_22__SCAN_IN), .ZN(n4638) );
  NAND4_X1 U5245 ( .A1(n4641), .A2(n4640), .A3(n4639), .A4(n4638), .ZN(n4642)
         );
  NOR3_X1 U5246 ( .A1(n4644), .A2(n4643), .A3(n4642), .ZN(n4645) );
  AND4_X1 U5247 ( .A1(n4648), .A2(n4647), .A3(n4646), .A4(n4645), .ZN(n4649)
         );
  AOI21_X1 U5248 ( .B1(n4650), .B2(n4649), .A(IR_REG_12__SCAN_IN), .ZN(n4870)
         );
  AOI22_X1 U5249 ( .A1(n4888), .A2(keyinput11), .B1(n4652), .B2(keyinput41), 
        .ZN(n4651) );
  OAI221_X1 U5250 ( .B1(n4888), .B2(keyinput11), .C1(n4652), .C2(keyinput41), 
        .A(n4651), .ZN(n4662) );
  AOI22_X1 U5251 ( .A1(n3266), .A2(keyinput27), .B1(n4654), .B2(keyinput110), 
        .ZN(n4653) );
  OAI221_X1 U5252 ( .B1(n3266), .B2(keyinput27), .C1(n4654), .C2(keyinput110), 
        .A(n4653), .ZN(n4661) );
  AOI22_X1 U5253 ( .A1(n2832), .A2(keyinput112), .B1(keyinput47), .B2(n4656), 
        .ZN(n4655) );
  OAI221_X1 U5254 ( .B1(n2832), .B2(keyinput112), .C1(n4656), .C2(keyinput47), 
        .A(n4655), .ZN(n4660) );
  AOI22_X1 U5255 ( .A1(n4658), .A2(keyinput126), .B1(n2701), .B2(keyinput122), 
        .ZN(n4657) );
  OAI221_X1 U5256 ( .B1(n4658), .B2(keyinput126), .C1(n2701), .C2(keyinput122), 
        .A(n4657), .ZN(n4659) );
  NOR4_X1 U5257 ( .A1(n4662), .A2(n4661), .A3(n4660), .A4(n4659), .ZN(n4702)
         );
  AOI22_X1 U5258 ( .A1(n5046), .A2(keyinput118), .B1(keyinput117), .B2(n4664), 
        .ZN(n4663) );
  OAI221_X1 U5259 ( .B1(n5046), .B2(keyinput118), .C1(n4664), .C2(keyinput117), 
        .A(n4663), .ZN(n4674) );
  AOI22_X1 U5260 ( .A1(n4666), .A2(keyinput120), .B1(n2724), .B2(keyinput116), 
        .ZN(n4665) );
  OAI221_X1 U5261 ( .B1(n4666), .B2(keyinput120), .C1(n2724), .C2(keyinput116), 
        .A(n4665), .ZN(n4673) );
  INV_X1 U5262 ( .A(D_REG_18__SCAN_IN), .ZN(n5041) );
  AOI22_X1 U5263 ( .A1(n4668), .A2(keyinput100), .B1(n5041), .B2(keyinput102), 
        .ZN(n4667) );
  OAI221_X1 U5264 ( .B1(n4668), .B2(keyinput100), .C1(n5041), .C2(keyinput102), 
        .A(n4667), .ZN(n4672) );
  XOR2_X1 U5265 ( .A(n2497), .B(keyinput104), .Z(n4670) );
  XNOR2_X1 U5266 ( .A(IR_REG_21__SCAN_IN), .B(keyinput109), .ZN(n4669) );
  NAND2_X1 U5267 ( .A1(n4670), .A2(n4669), .ZN(n4671) );
  NOR4_X1 U5268 ( .A1(n4674), .A2(n4673), .A3(n4672), .A4(n4671), .ZN(n4701)
         );
  INV_X1 U5269 ( .A(D_REG_17__SCAN_IN), .ZN(n5042) );
  INV_X1 U5270 ( .A(D_REG_25__SCAN_IN), .ZN(n5038) );
  AOI22_X1 U5271 ( .A1(n5042), .A2(keyinput97), .B1(keyinput93), .B2(n5038), 
        .ZN(n4675) );
  OAI221_X1 U5272 ( .B1(n5042), .B2(keyinput97), .C1(n5038), .C2(keyinput93), 
        .A(n4675), .ZN(n4684) );
  AOI22_X1 U5273 ( .A1(n4678), .A2(keyinput84), .B1(keyinput82), .B2(n4677), 
        .ZN(n4676) );
  OAI221_X1 U5274 ( .B1(n4678), .B2(keyinput84), .C1(n4677), .C2(keyinput82), 
        .A(n4676), .ZN(n4683) );
  AOI22_X1 U5275 ( .A1(n5036), .A2(keyinput81), .B1(n2524), .B2(keyinput78), 
        .ZN(n4679) );
  OAI221_X1 U5276 ( .B1(n5036), .B2(keyinput81), .C1(n2524), .C2(keyinput78), 
        .A(n4679), .ZN(n4682) );
  AOI22_X1 U5277 ( .A1(n5051), .A2(keyinput77), .B1(n2507), .B2(keyinput73), 
        .ZN(n4680) );
  OAI221_X1 U5278 ( .B1(n5051), .B2(keyinput77), .C1(n2507), .C2(keyinput73), 
        .A(n4680), .ZN(n4681) );
  NOR4_X1 U5279 ( .A1(n4684), .A2(n4683), .A3(n4682), .A4(n4681), .ZN(n4700)
         );
  AOI22_X1 U5280 ( .A1(n4687), .A2(keyinput72), .B1(keyinput68), .B2(n4686), 
        .ZN(n4685) );
  OAI221_X1 U5281 ( .B1(n4687), .B2(keyinput72), .C1(n4686), .C2(keyinput68), 
        .A(n4685), .ZN(n4698) );
  INV_X1 U5282 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n4689) );
  AOI22_X1 U5283 ( .A1(n5045), .A2(keyinput54), .B1(keyinput48), .B2(n4689), 
        .ZN(n4688) );
  OAI221_X1 U5284 ( .B1(n5045), .B2(keyinput54), .C1(n4689), .C2(keyinput48), 
        .A(n4688), .ZN(n4697) );
  AOI22_X1 U5285 ( .A1(n4692), .A2(keyinput62), .B1(n4691), .B2(keyinput52), 
        .ZN(n4690) );
  OAI221_X1 U5286 ( .B1(n4692), .B2(keyinput62), .C1(n4691), .C2(keyinput52), 
        .A(n4690), .ZN(n4696) );
  XNOR2_X1 U5287 ( .A(IR_REG_27__SCAN_IN), .B(keyinput70), .ZN(n4694) );
  XNOR2_X1 U5288 ( .A(DATAI_8_), .B(keyinput60), .ZN(n4693) );
  NAND2_X1 U5289 ( .A1(n4694), .A2(n4693), .ZN(n4695) );
  NOR4_X1 U5290 ( .A1(n4698), .A2(n4697), .A3(n4696), .A4(n4695), .ZN(n4699)
         );
  NAND4_X1 U5291 ( .A1(n4702), .A2(n4701), .A3(n4700), .A4(n4699), .ZN(n4868)
         );
  AOI22_X1 U5292 ( .A1(n4704), .A2(keyinput45), .B1(n4621), .B2(keyinput36), 
        .ZN(n4703) );
  OAI221_X1 U5293 ( .B1(n4704), .B2(keyinput45), .C1(n4621), .C2(keyinput36), 
        .A(n4703), .ZN(n4708) );
  XNOR2_X1 U5294 ( .A(n4705), .B(keyinput42), .ZN(n4707) );
  XNOR2_X1 U5295 ( .A(n5034), .B(keyinput46), .ZN(n4706) );
  OR3_X1 U5296 ( .A1(n4708), .A2(n4707), .A3(n4706), .ZN(n4715) );
  INV_X1 U5297 ( .A(D_REG_16__SCAN_IN), .ZN(n5043) );
  INV_X1 U5298 ( .A(D_REG_24__SCAN_IN), .ZN(n5039) );
  AOI22_X1 U5299 ( .A1(n5043), .A2(keyinput14), .B1(keyinput67), .B2(n5039), 
        .ZN(n4709) );
  OAI221_X1 U5300 ( .B1(n5043), .B2(keyinput14), .C1(n5039), .C2(keyinput67), 
        .A(n4709), .ZN(n4714) );
  AOI22_X1 U5301 ( .A1(n4712), .A2(keyinput33), .B1(n4711), .B2(keyinput25), 
        .ZN(n4710) );
  OAI221_X1 U5302 ( .B1(n4712), .B2(keyinput33), .C1(n4711), .C2(keyinput25), 
        .A(n4710), .ZN(n4713) );
  NOR3_X1 U5303 ( .A1(n4715), .A2(n4714), .A3(n4713), .ZN(n4756) );
  INV_X1 U5304 ( .A(D_REG_15__SCAN_IN), .ZN(n5044) );
  AOI22_X1 U5305 ( .A1(n5044), .A2(keyinput123), .B1(n2911), .B2(keyinput22), 
        .ZN(n4716) );
  OAI221_X1 U5306 ( .B1(n5044), .B2(keyinput123), .C1(n2911), .C2(keyinput22), 
        .A(n4716), .ZN(n4724) );
  INV_X1 U5307 ( .A(D_REG_28__SCAN_IN), .ZN(n5037) );
  INV_X1 U5308 ( .A(D_REG_30__SCAN_IN), .ZN(n5035) );
  AOI22_X1 U5309 ( .A1(n5037), .A2(keyinput3), .B1(n5035), .B2(keyinput16), 
        .ZN(n4717) );
  OAI221_X1 U5310 ( .B1(n5037), .B2(keyinput3), .C1(n5035), .C2(keyinput16), 
        .A(n4717), .ZN(n4723) );
  XOR2_X1 U5311 ( .A(n2486), .B(keyinput21), .Z(n4720) );
  XNOR2_X1 U5312 ( .A(IR_REG_17__SCAN_IN), .B(keyinput119), .ZN(n4719) );
  XNOR2_X1 U5313 ( .A(IR_REG_26__SCAN_IN), .B(keyinput71), .ZN(n4718) );
  NAND3_X1 U5314 ( .A1(n4720), .A2(n4719), .A3(n4718), .ZN(n4722) );
  INV_X1 U5315 ( .A(D_REG_21__SCAN_IN), .ZN(n5040) );
  XNOR2_X1 U5316 ( .A(n5040), .B(keyinput26), .ZN(n4721) );
  NOR4_X1 U5317 ( .A1(n4724), .A2(n4723), .A3(n4722), .A4(n4721), .ZN(n4755)
         );
  AOI22_X1 U5318 ( .A1(n4727), .A2(keyinput31), .B1(keyinput12), .B2(n4726), 
        .ZN(n4725) );
  OAI221_X1 U5319 ( .B1(n4727), .B2(keyinput31), .C1(n4726), .C2(keyinput12), 
        .A(n4725), .ZN(n4739) );
  AOI22_X1 U5320 ( .A1(n4730), .A2(keyinput2), .B1(n4729), .B2(keyinput0), 
        .ZN(n4728) );
  OAI221_X1 U5321 ( .B1(n4730), .B2(keyinput2), .C1(n4729), .C2(keyinput0), 
        .A(n4728), .ZN(n4738) );
  AOI22_X1 U5322 ( .A1(n4733), .A2(keyinput1), .B1(keyinput34), .B2(n4732), 
        .ZN(n4731) );
  OAI221_X1 U5323 ( .B1(n4733), .B2(keyinput1), .C1(n4732), .C2(keyinput34), 
        .A(n4731), .ZN(n4737) );
  INV_X1 U5324 ( .A(DATAI_23_), .ZN(n5050) );
  INV_X1 U5325 ( .A(DATAI_22_), .ZN(n4735) );
  AOI22_X1 U5326 ( .A1(n5050), .A2(keyinput75), .B1(keyinput29), .B2(n4735), 
        .ZN(n4734) );
  OAI221_X1 U5327 ( .B1(n5050), .B2(keyinput75), .C1(n4735), .C2(keyinput29), 
        .A(n4734), .ZN(n4736) );
  NOR4_X1 U5328 ( .A1(n4739), .A2(n4738), .A3(n4737), .A4(n4736), .ZN(n4754)
         );
  AOI22_X1 U5329 ( .A1(n2569), .A2(keyinput24), .B1(keyinput9), .B2(n4741), 
        .ZN(n4740) );
  OAI221_X1 U5330 ( .B1(n2569), .B2(keyinput24), .C1(n4741), .C2(keyinput9), 
        .A(n4740), .ZN(n4752) );
  AOI22_X1 U5331 ( .A1(n4744), .A2(keyinput111), .B1(keyinput55), .B2(n4743), 
        .ZN(n4742) );
  OAI221_X1 U5332 ( .B1(n4744), .B2(keyinput111), .C1(n4743), .C2(keyinput55), 
        .A(n4742), .ZN(n4751) );
  XOR2_X1 U5333 ( .A(n4745), .B(keyinput127), .Z(n4749) );
  XOR2_X1 U5334 ( .A(n4626), .B(keyinput23), .Z(n4748) );
  XNOR2_X1 U5335 ( .A(REG3_REG_6__SCAN_IN), .B(keyinput17), .ZN(n4747) );
  XNOR2_X1 U5336 ( .A(IR_REG_4__SCAN_IN), .B(keyinput43), .ZN(n4746) );
  NAND4_X1 U5337 ( .A1(n4749), .A2(n4748), .A3(n4747), .A4(n4746), .ZN(n4750)
         );
  NOR3_X1 U5338 ( .A1(n4752), .A2(n4751), .A3(n4750), .ZN(n4753) );
  NAND4_X1 U5339 ( .A1(n4756), .A2(n4755), .A3(n4754), .A4(n4753), .ZN(n4867)
         );
  AOI22_X1 U5340 ( .A1(n4939), .A2(keyinput99), .B1(n4758), .B2(keyinput87), 
        .ZN(n4757) );
  OAI221_X1 U5341 ( .B1(n4939), .B2(keyinput99), .C1(n4758), .C2(keyinput87), 
        .A(n4757), .ZN(n4769) );
  AOI22_X1 U5342 ( .A1(n4761), .A2(keyinput89), .B1(keyinput30), .B2(n4760), 
        .ZN(n4759) );
  OAI221_X1 U5343 ( .B1(n4761), .B2(keyinput89), .C1(n4760), .C2(keyinput30), 
        .A(n4759), .ZN(n4768) );
  AOI22_X1 U5344 ( .A1(n4763), .A2(keyinput66), .B1(keyinput56), .B2(n2598), 
        .ZN(n4762) );
  OAI221_X1 U5345 ( .B1(n4763), .B2(keyinput66), .C1(n2598), .C2(keyinput56), 
        .A(n4762), .ZN(n4767) );
  INV_X1 U5346 ( .A(DATAI_13_), .ZN(n5058) );
  AOI22_X1 U5347 ( .A1(n5058), .A2(keyinput113), .B1(keyinput90), .B2(n4765), 
        .ZN(n4764) );
  OAI221_X1 U5348 ( .B1(n5058), .B2(keyinput113), .C1(n4765), .C2(keyinput90), 
        .A(n4764), .ZN(n4766) );
  NOR4_X1 U5349 ( .A1(n4769), .A2(n4768), .A3(n4767), .A4(n4766), .ZN(n4807)
         );
  AOI22_X1 U5350 ( .A1(n4623), .A2(keyinput76), .B1(n3228), .B2(keyinput19), 
        .ZN(n4770) );
  OAI221_X1 U5351 ( .B1(n4623), .B2(keyinput76), .C1(n3228), .C2(keyinput19), 
        .A(n4770), .ZN(n4779) );
  AOI22_X1 U5352 ( .A1(n4586), .A2(keyinput88), .B1(keyinput96), .B2(n3414), 
        .ZN(n4771) );
  OAI221_X1 U5353 ( .B1(n4586), .B2(keyinput88), .C1(n3414), .C2(keyinput96), 
        .A(n4771), .ZN(n4778) );
  AOI22_X1 U5354 ( .A1(n3687), .A2(keyinput15), .B1(n4773), .B2(keyinput40), 
        .ZN(n4772) );
  OAI221_X1 U5355 ( .B1(n3687), .B2(keyinput15), .C1(n4773), .C2(keyinput40), 
        .A(n4772), .ZN(n4777) );
  XOR2_X1 U5356 ( .A(n2568), .B(keyinput74), .Z(n4775) );
  XNOR2_X1 U5357 ( .A(REG1_REG_1__SCAN_IN), .B(keyinput83), .ZN(n4774) );
  NAND2_X1 U5358 ( .A1(n4775), .A2(n4774), .ZN(n4776) );
  NOR4_X1 U5359 ( .A1(n4779), .A2(n4778), .A3(n4777), .A4(n4776), .ZN(n4806)
         );
  INV_X1 U5360 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4781) );
  AOI22_X1 U5361 ( .A1(n4353), .A2(keyinput51), .B1(n4781), .B2(keyinput86), 
        .ZN(n4780) );
  OAI221_X1 U5362 ( .B1(n4353), .B2(keyinput51), .C1(n4781), .C2(keyinput86), 
        .A(n4780), .ZN(n4790) );
  AOI22_X1 U5363 ( .A1(n4784), .A2(keyinput114), .B1(keyinput35), .B2(n4783), 
        .ZN(n4782) );
  OAI221_X1 U5364 ( .B1(n4784), .B2(keyinput114), .C1(n4783), .C2(keyinput35), 
        .A(n4782), .ZN(n4789) );
  AOI22_X1 U5365 ( .A1(n4909), .A2(keyinput39), .B1(n4893), .B2(keyinput49), 
        .ZN(n4785) );
  OAI221_X1 U5366 ( .B1(n4909), .B2(keyinput39), .C1(n4893), .C2(keyinput49), 
        .A(n4785), .ZN(n4788) );
  AOI22_X1 U5367 ( .A1(n4523), .A2(keyinput91), .B1(n3911), .B2(keyinput20), 
        .ZN(n4786) );
  OAI221_X1 U5368 ( .B1(n4523), .B2(keyinput91), .C1(n3911), .C2(keyinput20), 
        .A(n4786), .ZN(n4787) );
  NOR4_X1 U5369 ( .A1(n4790), .A2(n4789), .A3(n4788), .A4(n4787), .ZN(n4805)
         );
  INV_X1 U5370 ( .A(DATAI_9_), .ZN(n4792) );
  AOI22_X1 U5371 ( .A1(n2614), .A2(keyinput38), .B1(keyinput18), .B2(n4792), 
        .ZN(n4791) );
  OAI221_X1 U5372 ( .B1(n2614), .B2(keyinput38), .C1(n4792), .C2(keyinput18), 
        .A(n4791), .ZN(n4803) );
  AOI22_X1 U5373 ( .A1(n4794), .A2(keyinput69), .B1(n4925), .B2(keyinput124), 
        .ZN(n4793) );
  OAI221_X1 U5374 ( .B1(n4794), .B2(keyinput69), .C1(n4925), .C2(keyinput124), 
        .A(n4793), .ZN(n4802) );
  AOI22_X1 U5375 ( .A1(n4797), .A2(keyinput106), .B1(n4796), .B2(keyinput92), 
        .ZN(n4795) );
  OAI221_X1 U5376 ( .B1(n4797), .B2(keyinput106), .C1(n4796), .C2(keyinput92), 
        .A(n4795), .ZN(n4801) );
  XNOR2_X1 U5377 ( .A(IR_REG_6__SCAN_IN), .B(keyinput53), .ZN(n4799) );
  XNOR2_X1 U5378 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput121), .ZN(n4798) );
  NAND2_X1 U5379 ( .A1(n4799), .A2(n4798), .ZN(n4800) );
  NOR4_X1 U5380 ( .A1(n4803), .A2(n4802), .A3(n4801), .A4(n4800), .ZN(n4804)
         );
  NAND4_X1 U5381 ( .A1(n4807), .A2(n4806), .A3(n4805), .A4(n4804), .ZN(n4866)
         );
  AOI22_X1 U5382 ( .A1(n4810), .A2(keyinput108), .B1(n4809), .B2(keyinput85), 
        .ZN(n4808) );
  OAI221_X1 U5383 ( .B1(n4810), .B2(keyinput108), .C1(n4809), .C2(keyinput85), 
        .A(n4808), .ZN(n4823) );
  AOI22_X1 U5384 ( .A1(n4813), .A2(keyinput98), .B1(keyinput37), .B2(n4812), 
        .ZN(n4811) );
  OAI221_X1 U5385 ( .B1(n4813), .B2(keyinput98), .C1(n4812), .C2(keyinput37), 
        .A(n4811), .ZN(n4822) );
  INV_X1 U5386 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4816) );
  AOI22_X1 U5387 ( .A1(n4816), .A2(keyinput103), .B1(n4815), .B2(keyinput57), 
        .ZN(n4814) );
  OAI221_X1 U5388 ( .B1(n4816), .B2(keyinput103), .C1(n4815), .C2(keyinput57), 
        .A(n4814), .ZN(n4821) );
  AOI22_X1 U5389 ( .A1(n4819), .A2(keyinput8), .B1(n4818), .B2(keyinput125), 
        .ZN(n4817) );
  OAI221_X1 U5390 ( .B1(n4819), .B2(keyinput8), .C1(n4818), .C2(keyinput125), 
        .A(n4817), .ZN(n4820) );
  NOR4_X1 U5391 ( .A1(n4823), .A2(n4822), .A3(n4821), .A4(n4820), .ZN(n4864)
         );
  INV_X1 U5392 ( .A(keyinput95), .ZN(n4825) );
  XOR2_X1 U5393 ( .A(n4431), .B(keyinput115), .Z(n4824) );
  OAI21_X1 U5394 ( .B1(IR_REG_12__SCAN_IN), .B2(n4825), .A(n4824), .ZN(n4835)
         );
  AOI22_X1 U5395 ( .A1(n4827), .A2(keyinput63), .B1(n4536), .B2(keyinput44), 
        .ZN(n4826) );
  OAI221_X1 U5396 ( .B1(n4827), .B2(keyinput63), .C1(n4536), .C2(keyinput44), 
        .A(n4826), .ZN(n4834) );
  AOI22_X1 U5397 ( .A1(n2937), .A2(keyinput79), .B1(keyinput65), .B2(n4829), 
        .ZN(n4828) );
  OAI221_X1 U5398 ( .B1(n2937), .B2(keyinput79), .C1(n4829), .C2(keyinput65), 
        .A(n4828), .ZN(n4833) );
  AOI22_X1 U5399 ( .A1(n2713), .A2(keyinput32), .B1(keyinput10), .B2(n4831), 
        .ZN(n4830) );
  OAI221_X1 U5400 ( .B1(n2713), .B2(keyinput32), .C1(n4831), .C2(keyinput10), 
        .A(n4830), .ZN(n4832) );
  NOR4_X1 U5401 ( .A1(n4835), .A2(n4834), .A3(n4833), .A4(n4832), .ZN(n4863)
         );
  INV_X1 U5402 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n4838) );
  AOI22_X1 U5403 ( .A1(n4838), .A2(keyinput28), .B1(n4837), .B2(keyinput105), 
        .ZN(n4836) );
  OAI221_X1 U5404 ( .B1(n4838), .B2(keyinput28), .C1(n4837), .C2(keyinput105), 
        .A(n4836), .ZN(n4848) );
  INV_X1 U5405 ( .A(ADDR_REG_11__SCAN_IN), .ZN(n4840) );
  AOI22_X1 U5406 ( .A1(n4840), .A2(keyinput6), .B1(n2657), .B2(keyinput13), 
        .ZN(n4839) );
  OAI221_X1 U5407 ( .B1(n4840), .B2(keyinput6), .C1(n2657), .C2(keyinput13), 
        .A(n4839), .ZN(n4847) );
  AOI22_X1 U5408 ( .A1(n4547), .A2(keyinput7), .B1(keyinput107), .B2(n4842), 
        .ZN(n4841) );
  OAI221_X1 U5409 ( .B1(n4547), .B2(keyinput7), .C1(n4842), .C2(keyinput107), 
        .A(n4841), .ZN(n4846) );
  INV_X1 U5410 ( .A(ADDR_REG_17__SCAN_IN), .ZN(n4844) );
  AOI22_X1 U5411 ( .A1(n5004), .A2(keyinput64), .B1(n4844), .B2(keyinput59), 
        .ZN(n4843) );
  OAI221_X1 U5412 ( .B1(n5004), .B2(keyinput64), .C1(n4844), .C2(keyinput59), 
        .A(n4843), .ZN(n4845) );
  NOR4_X1 U5413 ( .A1(n4848), .A2(n4847), .A3(n4846), .A4(n4845), .ZN(n4862)
         );
  AOI22_X1 U5414 ( .A1(n2532), .A2(keyinput4), .B1(keyinput58), .B2(n4850), 
        .ZN(n4849) );
  OAI221_X1 U5415 ( .B1(n2532), .B2(keyinput4), .C1(n4850), .C2(keyinput58), 
        .A(n4849), .ZN(n4860) );
  AOI22_X1 U5416 ( .A1(n4852), .A2(keyinput50), .B1(n3645), .B2(keyinput101), 
        .ZN(n4851) );
  OAI221_X1 U5417 ( .B1(n4852), .B2(keyinput50), .C1(n3645), .C2(keyinput101), 
        .A(n4851), .ZN(n4859) );
  XNOR2_X1 U5418 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput61), .ZN(n4855) );
  XNOR2_X1 U5419 ( .A(REG1_REG_0__SCAN_IN), .B(keyinput80), .ZN(n4854) );
  XNOR2_X1 U5420 ( .A(DATAI_20_), .B(keyinput5), .ZN(n4853) );
  NAND3_X1 U5421 ( .A1(n4855), .A2(n4854), .A3(n4853), .ZN(n4858) );
  XNOR2_X1 U5422 ( .A(n4856), .B(keyinput94), .ZN(n4857) );
  NOR4_X1 U5423 ( .A1(n4860), .A2(n4859), .A3(n4858), .A4(n4857), .ZN(n4861)
         );
  NAND4_X1 U5424 ( .A1(n4864), .A2(n4863), .A3(n4862), .A4(n4861), .ZN(n4865)
         );
  NOR4_X1 U5425 ( .A1(n4868), .A2(n4867), .A3(n4866), .A4(n4865), .ZN(n4869)
         );
  OAI21_X1 U5426 ( .B1(n4870), .B2(keyinput95), .A(n4869), .ZN(n4877) );
  OAI22_X1 U5427 ( .A1(n4873), .A2(n4872), .B1(n5081), .B2(n4871), .ZN(n4874)
         );
  AOI21_X1 U5428 ( .B1(n4875), .B2(n5081), .A(n4874), .ZN(n4876) );
  XOR2_X1 U5429 ( .A(n4877), .B(n4876), .Z(U3520) );
  NAND2_X1 U5430 ( .A1(n5076), .A2(n4878), .ZN(n4880) );
  NAND2_X1 U5431 ( .A1(n5075), .A2(REG0_REG_31__SCAN_IN), .ZN(n4879) );
  OAI211_X1 U5432 ( .C1(n4881), .C2(n4945), .A(n4880), .B(n4879), .ZN(U3517)
         );
  INV_X1 U5433 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4886) );
  NAND2_X1 U5434 ( .A1(n4882), .A2(n4935), .ZN(n4885) );
  NAND2_X1 U5435 ( .A1(n5076), .A2(n4883), .ZN(n4884) );
  OAI211_X1 U5436 ( .C1(n5076), .C2(n4886), .A(n4885), .B(n4884), .ZN(U3516)
         );
  OAI21_X1 U5437 ( .B1(n4890), .B2(n4945), .A(n4889), .ZN(U3513) );
  INV_X1 U5438 ( .A(n4891), .ZN(n4892) );
  MUX2_X1 U5439 ( .A(n4893), .B(n4892), .S(n5076), .Z(n4894) );
  OAI21_X1 U5440 ( .B1(n4895), .B2(n4945), .A(n4894), .ZN(U3512) );
  INV_X1 U5441 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4897) );
  MUX2_X1 U5442 ( .A(n4897), .B(n4896), .S(n5076), .Z(n4898) );
  OAI21_X1 U5443 ( .B1(n4899), .B2(n4945), .A(n4898), .ZN(U3511) );
  INV_X1 U5444 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4901) );
  MUX2_X1 U5445 ( .A(n4901), .B(n4900), .S(n5076), .Z(n4902) );
  OAI21_X1 U5446 ( .B1(n4903), .B2(n4945), .A(n4902), .ZN(U3510) );
  INV_X1 U5447 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4905) );
  MUX2_X1 U5448 ( .A(n4905), .B(n4904), .S(n5076), .Z(n4906) );
  OAI21_X1 U5449 ( .B1(n4907), .B2(n4945), .A(n4906), .ZN(U3509) );
  MUX2_X1 U5450 ( .A(n4909), .B(n4908), .S(n5076), .Z(n4910) );
  OAI21_X1 U5451 ( .B1(n4911), .B2(n4945), .A(n4910), .ZN(U3508) );
  MUX2_X1 U5452 ( .A(n4781), .B(n4912), .S(n5076), .Z(n4913) );
  OAI21_X1 U5453 ( .B1(n4914), .B2(n4945), .A(n4913), .ZN(U3507) );
  INV_X1 U5454 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4916) );
  MUX2_X1 U5455 ( .A(n4916), .B(n4915), .S(n5076), .Z(n4917) );
  OAI21_X1 U5456 ( .B1(n4918), .B2(n4945), .A(n4917), .ZN(U3506) );
  INV_X1 U5457 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4920) );
  MUX2_X1 U5458 ( .A(n4920), .B(n4919), .S(n5076), .Z(n4921) );
  OAI21_X1 U5459 ( .B1(n4922), .B2(n4945), .A(n4921), .ZN(U3505) );
  MUX2_X1 U5460 ( .A(REG0_REG_18__SCAN_IN), .B(n4923), .S(n5076), .Z(U3503) );
  MUX2_X1 U5461 ( .A(n4925), .B(n4924), .S(n5076), .Z(n4926) );
  OAI21_X1 U5462 ( .B1(n4927), .B2(n4945), .A(n4926), .ZN(U3501) );
  MUX2_X1 U5463 ( .A(REG0_REG_16__SCAN_IN), .B(n4928), .S(n5076), .Z(U3499) );
  MUX2_X1 U5464 ( .A(REG0_REG_15__SCAN_IN), .B(n4929), .S(n5076), .Z(n4930) );
  AOI21_X1 U5465 ( .B1(n4931), .B2(n4935), .A(n4930), .ZN(n4932) );
  INV_X1 U5466 ( .A(n4932), .ZN(U3497) );
  MUX2_X1 U5467 ( .A(REG0_REG_14__SCAN_IN), .B(n4933), .S(n5076), .Z(n4934) );
  AOI21_X1 U5468 ( .B1(n4936), .B2(n4935), .A(n4934), .ZN(n4937) );
  INV_X1 U5469 ( .A(n4937), .ZN(U3495) );
  MUX2_X1 U5470 ( .A(n4939), .B(n4938), .S(n5076), .Z(n4940) );
  OAI21_X1 U5471 ( .B1(n4941), .B2(n4945), .A(n4940), .ZN(U3493) );
  MUX2_X1 U5472 ( .A(n4943), .B(n4942), .S(n5076), .Z(n4944) );
  OAI21_X1 U5473 ( .B1(n4946), .B2(n4945), .A(n4944), .ZN(U3491) );
  MUX2_X1 U5474 ( .A(n4966), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U5475 ( .A(n4947), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5476 ( .A(n2879), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5477 ( .A(DATAI_22_), .B(n2946), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U5478 ( .A(DATAI_21_), .B(n4948), .S(STATE_REG_SCAN_IN), .Z(U3331)
         );
  MUX2_X1 U5479 ( .A(DATAI_20_), .B(n4949), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5480 ( .A(DATAI_19_), .B(n4950), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U5481 ( .A(n4951), .B(DATAI_12_), .S(U3149), .Z(U3340) );
  MUX2_X1 U5482 ( .A(n4953), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5483 ( .A(n4954), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5484 ( .A(DATAI_8_), .B(n4955), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5485 ( .A(DATAI_5_), .B(n4956), .S(STATE_REG_SCAN_IN), .Z(U3347) );
  MUX2_X1 U5486 ( .A(n4957), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5487 ( .A(n4958), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  OAI22_X1 U5488 ( .A1(U3149), .A2(n4959), .B1(DATAI_28_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4960) );
  INV_X1 U5489 ( .A(n4960), .ZN(U3324) );
  INV_X1 U5490 ( .A(n4961), .ZN(n4965) );
  OAI21_X1 U5491 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4966), .A(n4963), .ZN(n4962)
         );
  MUX2_X1 U5492 ( .A(n4963), .B(n4962), .S(n5060), .Z(n4964) );
  OAI21_X1 U5493 ( .B1(n4966), .B2(n4965), .A(n4964), .ZN(n4968) );
  AOI22_X1 U5494 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n5018), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4967) );
  OAI21_X1 U5495 ( .B1(n4969), .B2(n4968), .A(n4967), .ZN(U3240) );
  AOI21_X1 U5496 ( .B1(n2670), .B2(n5059), .A(n4970), .ZN(n4973) );
  OAI21_X1 U5497 ( .B1(n4973), .B2(n4972), .A(n5001), .ZN(n4971) );
  AOI21_X1 U5498 ( .B1(n4973), .B2(n4972), .A(n4971), .ZN(n4974) );
  AOI211_X1 U5499 ( .C1(n5018), .C2(ADDR_REG_13__SCAN_IN), .A(n4975), .B(n4974), .ZN(n4980) );
  OAI211_X1 U5500 ( .C1(n4978), .C2(n4977), .A(n3215), .B(n4976), .ZN(n4979)
         );
  OAI211_X1 U5501 ( .C1(n5024), .C2(n5059), .A(n4980), .B(n4979), .ZN(U3253)
         );
  AOI211_X1 U5502 ( .C1(n4983), .C2(n4982), .A(n4981), .B(n5014), .ZN(n4984)
         );
  AOI211_X1 U5503 ( .C1(n5018), .C2(ADDR_REG_15__SCAN_IN), .A(n4985), .B(n4984), .ZN(n4990) );
  OAI211_X1 U5504 ( .C1(n4988), .C2(n4987), .A(n3215), .B(n4986), .ZN(n4989)
         );
  OAI211_X1 U5505 ( .C1(n5024), .C2(n5057), .A(n4990), .B(n4989), .ZN(U3255)
         );
  OAI21_X1 U5506 ( .B1(n4993), .B2(n4992), .A(n4991), .ZN(n5000) );
  AOI21_X1 U5507 ( .B1(REG1_REG_16__SCAN_IN), .B2(n4995), .A(n4994), .ZN(n4998) );
  OAI22_X1 U5508 ( .A1(n4998), .A2(n4997), .B1(n4996), .B2(n5024), .ZN(n4999)
         );
  AOI21_X1 U5509 ( .B1(n5001), .B2(n5000), .A(n4999), .ZN(n5003) );
  OAI211_X1 U5510 ( .C1(n5005), .C2(n5004), .A(n5003), .B(n5002), .ZN(U3256)
         );
  OAI221_X1 U5511 ( .B1(n5010), .B2(n2159), .C1(n5010), .C2(n5011), .A(n3215), 
        .ZN(n5012) );
  OAI211_X1 U5512 ( .C1(n5024), .C2(n5053), .A(n5013), .B(n5012), .ZN(U3257)
         );
  OAI211_X1 U5513 ( .C1(n5021), .C2(n5020), .A(n3215), .B(n5019), .ZN(n5022)
         );
  OAI211_X1 U5514 ( .C1(n5024), .C2(n5052), .A(n5023), .B(n5022), .ZN(U3258)
         );
  AOI21_X1 U5515 ( .B1(n5027), .B2(n5026), .A(n5025), .ZN(n5033) );
  AOI22_X1 U5516 ( .A1(n5030), .A2(n5029), .B1(REG3_REG_0__SCAN_IN), .B2(n5028), .ZN(n5031) );
  OAI221_X1 U5517 ( .B1(n4337), .B2(n5033), .C1(n5032), .C2(n4623), .A(n5031), 
        .ZN(U3290) );
  NOR2_X1 U5518 ( .A1(n5047), .A2(n5034), .ZN(U3291) );
  NOR2_X1 U5519 ( .A1(n5047), .A2(n5035), .ZN(U3292) );
  NOR2_X1 U5520 ( .A1(n5047), .A2(n5036), .ZN(U3293) );
  NOR2_X1 U5521 ( .A1(n5047), .A2(n5037), .ZN(U3294) );
  AND2_X1 U5522 ( .A1(D_REG_27__SCAN_IN), .A2(n5048), .ZN(U3295) );
  AND2_X1 U5523 ( .A1(D_REG_26__SCAN_IN), .A2(n5048), .ZN(U3296) );
  NOR2_X1 U5524 ( .A1(n5047), .A2(n5038), .ZN(U3297) );
  NOR2_X1 U5525 ( .A1(n5047), .A2(n5039), .ZN(U3298) );
  AND2_X1 U5526 ( .A1(D_REG_23__SCAN_IN), .A2(n5048), .ZN(U3299) );
  AND2_X1 U5527 ( .A1(D_REG_22__SCAN_IN), .A2(n5048), .ZN(U3300) );
  NOR2_X1 U5528 ( .A1(n5047), .A2(n5040), .ZN(U3301) );
  AND2_X1 U5529 ( .A1(D_REG_20__SCAN_IN), .A2(n5048), .ZN(U3302) );
  AND2_X1 U5530 ( .A1(D_REG_19__SCAN_IN), .A2(n5048), .ZN(U3303) );
  NOR2_X1 U5531 ( .A1(n5047), .A2(n5041), .ZN(U3304) );
  NOR2_X1 U5532 ( .A1(n5047), .A2(n5042), .ZN(U3305) );
  NOR2_X1 U5533 ( .A1(n5047), .A2(n5043), .ZN(U3306) );
  NOR2_X1 U5534 ( .A1(n5047), .A2(n5044), .ZN(U3307) );
  AND2_X1 U5535 ( .A1(D_REG_14__SCAN_IN), .A2(n5048), .ZN(U3308) );
  AND2_X1 U5536 ( .A1(D_REG_13__SCAN_IN), .A2(n5048), .ZN(U3309) );
  AND2_X1 U5537 ( .A1(D_REG_12__SCAN_IN), .A2(n5048), .ZN(U3310) );
  NOR2_X1 U5538 ( .A1(n5047), .A2(n5045), .ZN(U3311) );
  AND2_X1 U5539 ( .A1(D_REG_10__SCAN_IN), .A2(n5048), .ZN(U3312) );
  NOR2_X1 U5540 ( .A1(n5047), .A2(n5046), .ZN(U3313) );
  AND2_X1 U5541 ( .A1(D_REG_8__SCAN_IN), .A2(n5048), .ZN(U3314) );
  AND2_X1 U5542 ( .A1(D_REG_7__SCAN_IN), .A2(n5048), .ZN(U3315) );
  AND2_X1 U5543 ( .A1(D_REG_6__SCAN_IN), .A2(n5048), .ZN(U3316) );
  AND2_X1 U5544 ( .A1(D_REG_5__SCAN_IN), .A2(n5048), .ZN(U3317) );
  AND2_X1 U5545 ( .A1(D_REG_4__SCAN_IN), .A2(n5048), .ZN(U3318) );
  AND2_X1 U5546 ( .A1(D_REG_3__SCAN_IN), .A2(n5048), .ZN(U3319) );
  AND2_X1 U5547 ( .A1(D_REG_2__SCAN_IN), .A2(n5048), .ZN(U3320) );
  AOI21_X1 U5548 ( .B1(U3149), .B2(n5050), .A(n5049), .ZN(U3329) );
  AOI22_X1 U5549 ( .A1(STATE_REG_SCAN_IN), .A2(n5052), .B1(n5051), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5550 ( .A1(STATE_REG_SCAN_IN), .A2(n5053), .B1(n2497), .B2(U3149), 
        .ZN(U3335) );
  OAI22_X1 U5551 ( .A1(U3149), .A2(n5054), .B1(DATAI_16_), .B2(
        STATE_REG_SCAN_IN), .ZN(n5055) );
  INV_X1 U5552 ( .A(n5055), .ZN(U3336) );
  AOI22_X1 U5553 ( .A1(STATE_REG_SCAN_IN), .A2(n5057), .B1(n5056), .B2(U3149), 
        .ZN(U3337) );
  AOI22_X1 U5554 ( .A1(STATE_REG_SCAN_IN), .A2(n5059), .B1(n5058), .B2(U3149), 
        .ZN(U3339) );
  OAI22_X1 U5555 ( .A1(U3149), .A2(n5060), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n5061) );
  INV_X1 U5556 ( .A(n5061), .ZN(U3352) );
  AOI22_X1 U5557 ( .A1(n5076), .A2(n5062), .B1(n2525), .B2(n5075), .ZN(U3467)
         );
  AOI22_X1 U5558 ( .A1(n5076), .A2(n5063), .B1(n2519), .B2(n5075), .ZN(U3469)
         );
  AND2_X1 U5559 ( .A1(n5065), .A2(n5064), .ZN(n5067) );
  NOR3_X1 U5560 ( .A1(n5068), .A2(n5067), .A3(n5066), .ZN(n5078) );
  AOI22_X1 U5561 ( .A1(n5076), .A2(n5078), .B1(n2561), .B2(n5075), .ZN(U3475)
         );
  NOR3_X1 U5562 ( .A1(n5071), .A2(n5070), .A3(n5069), .ZN(n5073) );
  NOR3_X1 U5563 ( .A1(n5074), .A2(n5073), .A3(n5072), .ZN(n5080) );
  AOI22_X1 U5564 ( .A1(n5076), .A2(n5080), .B1(n2587), .B2(n5075), .ZN(U3481)
         );
  AOI22_X1 U5565 ( .A1(n5081), .A2(n5078), .B1(n5077), .B2(n5079), .ZN(U3522)
         );
  AOI22_X1 U5566 ( .A1(n5081), .A2(n5080), .B1(n3414), .B2(n5079), .ZN(U3525)
         );
  CLKBUF_X1 U2453 ( .A(n2534), .Z(n3329) );
  CLKBUF_X2 U2571 ( .A(n2537), .Z(n3334) );
endmodule

