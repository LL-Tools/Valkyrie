

module b17_C_gen_AntiSAT_k_128_9 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, 
        keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, 
        keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, 
        keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, 
        keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, 
        keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, 
        keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, 
        keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, 
        keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, 
        keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, 
        keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, 
        keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, 
        keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, 
        keyinput_g61, keyinput_g62, keyinput_g63, U355, U356, U357, U358, U359, 
        U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, 
        U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, 
        U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, 
        U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, 
        U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, 
        U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, 
        U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, 
        U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
         n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
         n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
         n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
         n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
         n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
         n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
         n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
         n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
         n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
         n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142,
         n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214,
         n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
         n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
         n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
         n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
         n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014,
         n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
         n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
         n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
         n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
         n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
         n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
         n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
         n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
         n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
         n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
         n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
         n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
         n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
         n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
         n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
         n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
         n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
         n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
         n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
         n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
         n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294,
         n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
         n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
         n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
         n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
         n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
         n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
         n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
         n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
         n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
         n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982,
         n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
         n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
         n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
         n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
         n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
         n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
         n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
         n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
         n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
         n21119, n21120, n21121;

  NAND2_X1 U11074 ( .A1(n14545), .A2(n9817), .ZN(n14154) );
  BUF_X1 U11075 ( .A(n10418), .Z(n9665) );
  AND2_X1 U11076 ( .A1(n12242), .A2(n9780), .ZN(n14874) );
  OR2_X1 U11077 ( .A1(n13469), .A2(n9921), .ZN(n13366) );
  NAND2_X1 U11078 ( .A1(n10529), .A2(n10556), .ZN(n12218) );
  CLKBUF_X1 U11079 ( .A(n11312), .Z(n11375) );
  AND2_X1 U11080 ( .A1(n11521), .A2(n15841), .ZN(n11556) );
  AND2_X1 U11081 ( .A1(n15841), .A2(n11519), .ZN(n19613) );
  AND2_X1 U11082 ( .A1(n13138), .A2(n11511), .ZN(n11567) );
  AND2_X1 U11083 ( .A1(n11473), .A2(n11485), .ZN(n15823) );
  NAND2_X1 U11084 ( .A1(n10316), .A2(n10315), .ZN(n10362) );
  BUF_X2 U11085 ( .A(n12291), .Z(n9632) );
  CLKBUF_X2 U11086 ( .A(n14245), .Z(n14307) );
  INV_X1 U11087 ( .A(n12378), .ZN(n14301) );
  CLKBUF_X2 U11088 ( .A(n10363), .Z(n10977) );
  CLKBUF_X1 U11089 ( .A(n10981), .Z(n10820) );
  INV_X1 U11090 ( .A(n14289), .ZN(n12459) );
  INV_X1 U11091 ( .A(n14305), .ZN(n12466) );
  INV_X1 U11092 ( .A(n12408), .ZN(n14300) );
  INV_X1 U11093 ( .A(n14290), .ZN(n12460) );
  CLKBUF_X2 U11094 ( .A(n12596), .Z(n17231) );
  CLKBUF_X1 U11095 ( .A(n10979), .Z(n10831) );
  BUF_X2 U11096 ( .A(n10963), .Z(n9674) );
  CLKBUF_X2 U11097 ( .A(n10370), .Z(n9676) );
  CLKBUF_X2 U11098 ( .A(n9670), .Z(n10987) );
  CLKBUF_X2 U11100 ( .A(n12089), .Z(n9631) );
  INV_X1 U11101 ( .A(n12597), .ZN(n17114) );
  INV_X1 U11102 ( .A(n13246), .ZN(n20910) );
  INV_X1 U11103 ( .A(n17208), .ZN(n17142) );
  INV_X1 U11104 ( .A(n11305), .ZN(n19989) );
  BUF_X1 U11105 ( .A(n11398), .Z(n19288) );
  NAND2_X2 U11106 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18728) );
  NAND2_X1 U11107 ( .A1(n11342), .A2(n11341), .ZN(n19265) );
  AND2_X1 U11108 ( .A1(n10192), .A2(n10193), .ZN(n10369) );
  AND2_X1 U11109 ( .A1(n13431), .A2(n15163), .ZN(n10349) );
  OAI21_X1 U11110 ( .B1(n11395), .B2(n11394), .A(n11393), .ZN(n12519) );
  XNOR2_X1 U11111 ( .A(n10543), .B(n10553), .ZN(n12196) );
  AND4_X1 U11112 ( .A1(n10205), .A2(n10204), .A3(n10203), .A4(n10202), .ZN(
        n10206) );
  AND2_X1 U11113 ( .A1(n11221), .A2(n13761), .ZN(n9653) );
  OR2_X1 U11114 ( .A1(n11330), .A2(n16338), .ZN(n14305) );
  NAND2_X1 U11115 ( .A1(n10460), .A2(n10459), .ZN(n11024) );
  XNOR2_X1 U11116 ( .A(n12218), .B(n10559), .ZN(n12205) );
  AND2_X1 U11117 ( .A1(n10181), .A2(n10255), .ZN(n13315) );
  INV_X1 U11118 ( .A(n14303), .ZN(n12465) );
  NAND2_X1 U11119 ( .A1(n12553), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11856) );
  INV_X2 U11120 ( .A(n11388), .ZN(n16366) );
  NOR2_X1 U11121 ( .A1(n15859), .A2(n15823), .ZN(n11501) );
  OR2_X1 U11122 ( .A1(n10245), .A2(n10244), .ZN(n20267) );
  AND2_X1 U11123 ( .A1(n9875), .A2(n9872), .ZN(n9871) );
  NAND2_X1 U11124 ( .A1(n9969), .A2(n9970), .ZN(n11305) );
  AOI211_X1 U11126 ( .C1(n17230), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n12109), .B(n12108), .ZN(n18291) );
  INV_X1 U11127 ( .A(n20258), .ZN(n13310) );
  NOR2_X1 U11128 ( .A1(n14154), .A2(n11088), .ZN(n11008) );
  INV_X1 U11131 ( .A(n12601), .ZN(n17035) );
  AND2_X1 U11132 ( .A1(n10023), .A2(n10021), .ZN(n12692) );
  INV_X1 U11133 ( .A(n17815), .ZN(n10022) );
  NAND2_X1 U11134 ( .A1(n13177), .A2(n20244), .ZN(n12980) );
  INV_X1 U11135 ( .A(n20078), .ZN(n20093) );
  AND2_X1 U11136 ( .A1(n9831), .A2(n9830), .ZN(n14150) );
  NOR2_X2 U11137 ( .A1(n14775), .A2(n14692), .ZN(n14691) );
  NAND2_X2 U11138 ( .A1(n11261), .A2(n11260), .ZN(n11388) );
  INV_X1 U11139 ( .A(n19113), .ZN(n15544) );
  NOR2_X1 U11140 ( .A1(n18294), .A2(n17332), .ZN(n17328) );
  INV_X1 U11141 ( .A(n17184), .ZN(n17161) );
  INV_X1 U11142 ( .A(n17722), .ZN(n17748) );
  NOR2_X1 U11143 ( .A1(n18123), .A2(n18049), .ZN(n17743) );
  INV_X1 U11144 ( .A(n17912), .ZN(n17818) );
  INV_X1 U11145 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12022) );
  XNOR2_X1 U11146 ( .A(n14154), .B(n11088), .ZN(n14863) );
  BUF_X1 U11147 ( .A(n13115), .Z(n15841) );
  INV_X1 U11148 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19645) );
  NAND4_X1 U11149 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_24__SCAN_IN), .A4(n17003), .ZN(n16985) );
  AOI211_X1 U11150 ( .C1(n17225), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n12583), .B(n12582), .ZN(n17422) );
  AND3_X1 U11151 ( .A1(n9721), .A2(n10159), .A3(n10009), .ZN(n17434) );
  INV_X1 U11152 ( .A(n17696), .ZN(n17897) );
  INV_X1 U11153 ( .A(n17902), .ZN(n17916) );
  NAND2_X1 U11154 ( .A1(n10141), .A2(n10140), .ZN(n11330) );
  AND2_X1 U11155 ( .A1(n10193), .A2(n10190), .ZN(n10978) );
  INV_X1 U11156 ( .A(n12224), .ZN(n14972) );
  BUF_X4 U11157 ( .A(n17237), .Z(n9630) );
  INV_X1 U11158 ( .A(n17167), .ZN(n17237) );
  AOI21_X4 U11159 ( .B1(n11479), .B2(n11478), .A(n11848), .ZN(n11493) );
  NAND2_X2 U11161 ( .A1(n16067), .A2(n12204), .ZN(n16064) );
  AND2_X2 U11162 ( .A1(n9709), .A2(n10206), .ZN(n10300) );
  AOI211_X2 U11163 ( .C1(n16578), .C2(n18784), .A(n16577), .B(n16576), .ZN(
        n16581) );
  XNOR2_X1 U11164 ( .A(n12163), .B(n12164), .ZN(n13286) );
  NOR2_X2 U11165 ( .A1(n16854), .A2(n17257), .ZN(n17250) );
  OAI222_X1 U11166 ( .A1(n17280), .A2(n17279), .B1(n17278), .B2(n17285), .C1(
        n17277), .C2(n17274), .ZN(P3_U2702) );
  OR2_X1 U11167 ( .A1(n11184), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n11098) );
  NAND2_X2 U11168 ( .A1(n9658), .A2(n14490), .ZN(n11184) );
  NOR2_X1 U11169 ( .A1(n12014), .A2(n12017), .ZN(n12089) );
  AND2_X2 U11170 ( .A1(n14595), .A2(n10121), .ZN(n14545) );
  AND2_X2 U11171 ( .A1(n14609), .A2(n14608), .ZN(n14595) );
  NOR2_X2 U11172 ( .A1(n18728), .A2(n12020), .ZN(n12596) );
  INV_X1 U11173 ( .A(n11417), .ZN(n12291) );
  NAND2_X2 U11174 ( .A1(n13061), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12163) );
  AOI21_X2 U11175 ( .B1(n10418), .B2(n20914), .A(n9723), .ZN(n12156) );
  BUF_X4 U11176 ( .A(n15863), .Z(n9633) );
  AND2_X4 U11177 ( .A1(n11221), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11312) );
  OAI22_X2 U11178 ( .A1(n18123), .A2(n17916), .B1(n17758), .B2(n17782), .ZN(
        n17774) );
  NOR2_X2 U11179 ( .A1(n17511), .A2(n17313), .ZN(n17305) );
  NAND2_X2 U11180 ( .A1(n10473), .A2(n10474), .ZN(n10507) );
  AOI21_X2 U11181 ( .B1(n11797), .B2(n15461), .A(n19114), .ZN(n11680) );
  XNOR2_X1 U11182 ( .A(n10359), .B(n10358), .ZN(n9779) );
  OAI22_X2 U11183 ( .A1(n13775), .A2(n13776), .B1(n11680), .B2(n13789), .ZN(
        n13927) );
  XNOR2_X1 U11184 ( .A(n14356), .B(n14358), .ZN(n15259) );
  CLKBUF_X1 U11185 ( .A(n15532), .Z(n15533) );
  NAND2_X1 U11186 ( .A1(n12692), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17574) );
  OR2_X1 U11187 ( .A1(n10022), .A2(n17610), .ZN(n17601) );
  NAND2_X1 U11188 ( .A1(n11810), .A2(n11811), .ZN(n13597) );
  AND2_X2 U11189 ( .A1(n12218), .A2(n12217), .ZN(n12224) );
  OR2_X1 U11190 ( .A1(n15653), .A2(n15473), .ZN(n15648) );
  BUF_X1 U11192 ( .A(n11563), .Z(n11564) );
  AND2_X1 U11193 ( .A1(n14039), .A2(n14038), .ZN(n16115) );
  INV_X1 U11194 ( .A(n19250), .ZN(n19245) );
  AND2_X1 U11195 ( .A1(n11521), .A2(n13680), .ZN(n11555) );
  AND2_X1 U11196 ( .A1(n11519), .A2(n13680), .ZN(n19771) );
  OR2_X2 U11197 ( .A1(n9779), .A2(n10424), .ZN(n10475) );
  AND2_X1 U11198 ( .A1(n13138), .A2(n11517), .ZN(n11565) );
  INV_X1 U11199 ( .A(n15874), .ZN(n15877) );
  NAND2_X1 U11200 ( .A1(n13696), .A2(n13695), .ZN(n13746) );
  INV_X1 U11201 ( .A(n11482), .ZN(n11849) );
  OR2_X1 U11202 ( .A1(n17876), .A2(n9698), .ZN(n10013) );
  NAND2_X1 U11203 ( .A1(n11424), .A2(n15828), .ZN(n12553) );
  CLKBUF_X2 U11204 ( .A(n11463), .Z(n11897) );
  XOR2_X1 U11205 ( .A(n18207), .B(n12665), .Z(n17876) );
  NOR2_X1 U11206 ( .A1(n17291), .A2(n18277), .ZN(n12711) );
  AOI211_X2 U11207 ( .C1(n17225), .C2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n12052), .B(n12051), .ZN(n17291) );
  INV_X1 U11208 ( .A(n12725), .ZN(n17445) );
  NAND4_X1 U11209 ( .A1(n12656), .A2(n12655), .A3(n12654), .A4(n12653), .ZN(
        n17911) );
  INV_X8 U11210 ( .A(n12291), .ZN(n19275) );
  AND2_X1 U11211 ( .A1(n11418), .A2(n11413), .ZN(n12525) );
  OAI21_X1 U11212 ( .B1(n13315), .B2(n12247), .A(n9772), .ZN(n10258) );
  INV_X1 U11213 ( .A(n11390), .ZN(n11387) );
  CLKBUF_X1 U11214 ( .A(n11305), .Z(n11412) );
  INV_X1 U11215 ( .A(n14160), .ZN(n10304) );
  INV_X1 U11216 ( .A(n12969), .ZN(n9634) );
  AND3_X2 U11217 ( .A1(n9970), .A2(n9969), .A3(n19645), .ZN(n14168) );
  NAND2_X1 U11218 ( .A1(n11259), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11260) );
  NAND2_X1 U11219 ( .A1(n11327), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11328) );
  AND4_X1 U11220 ( .A1(n11321), .A2(n11320), .A3(n11319), .A4(n11318), .ZN(
        n11322) );
  AND4_X1 U11221 ( .A1(n11326), .A2(n11325), .A3(n11324), .A4(n11323), .ZN(
        n11327) );
  INV_X4 U11222 ( .A(n12100), .ZN(n17185) );
  INV_X4 U11223 ( .A(n17035), .ZN(n17202) );
  CLKBUF_X2 U11224 ( .A(n12644), .Z(n9652) );
  BUF_X1 U11225 ( .A(n12086), .Z(n17241) );
  INV_X4 U11226 ( .A(n17205), .ZN(n12616) );
  CLKBUF_X2 U11227 ( .A(n9631), .Z(n17204) );
  BUF_X2 U11228 ( .A(n10343), .Z(n10962) );
  CLKBUF_X2 U11229 ( .A(n10364), .Z(n10938) );
  CLKBUF_X2 U11230 ( .A(n10369), .Z(n10955) );
  BUF_X2 U11231 ( .A(n10348), .Z(n10986) );
  CLKBUF_X2 U11232 ( .A(n12033), .Z(n17235) );
  CLKBUF_X2 U11233 ( .A(n10250), .Z(n10980) );
  NOR2_X1 U11234 ( .A1(n12020), .A2(n12019), .ZN(n12644) );
  CLKBUF_X2 U11235 ( .A(n10349), .Z(n10988) );
  OR3_X1 U11236 ( .A1(n12014), .A2(n18897), .A3(n16926), .ZN(n12086) );
  AND2_X2 U11237 ( .A1(n10190), .A2(n10191), .ZN(n10289) );
  CLKBUF_X2 U11238 ( .A(n14271), .Z(n9657) );
  CLKBUF_X2 U11239 ( .A(n14271), .Z(n9656) );
  CLKBUF_X2 U11240 ( .A(n14271), .Z(n9655) );
  BUF_X2 U11241 ( .A(n10978), .Z(n9668) );
  AND3_X2 U11243 ( .A1(n13763), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14271) );
  INV_X8 U11244 ( .A(n12608), .ZN(n9635) );
  AND2_X2 U11245 ( .A1(n11221), .A2(n13761), .ZN(n14436) );
  AND2_X2 U11246 ( .A1(n11221), .A2(n13761), .ZN(n9654) );
  INV_X1 U11248 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13761) );
  INV_X4 U11249 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12023) );
  NOR2_X4 U11250 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10193) );
  NAND2_X1 U11251 ( .A1(n9915), .A2(n9913), .ZN(n15519) );
  NAND2_X1 U11252 ( .A1(n9788), .A2(n9786), .ZN(n15396) );
  OAI21_X1 U11253 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15413), .A(
        n15401), .ZN(n15579) );
  AND2_X1 U11254 ( .A1(n9915), .A2(n9914), .ZN(n15494) );
  NAND2_X1 U11255 ( .A1(n9915), .A2(n9740), .ZN(n15479) );
  NAND2_X1 U11256 ( .A1(n14874), .A2(n15044), .ZN(n9830) );
  AOI21_X1 U11257 ( .B1(n14572), .B2(n14583), .A(n14571), .ZN(n14901) );
  AND2_X1 U11258 ( .A1(n9912), .A2(n9909), .ZN(n15763) );
  AND2_X1 U11259 ( .A1(n15746), .A2(n15745), .ZN(n16243) );
  AND2_X1 U11260 ( .A1(n14892), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12242) );
  AND2_X2 U11261 ( .A1(n12241), .A2(n14923), .ZN(n14914) );
  CLKBUF_X1 U11262 ( .A(n15440), .Z(n9640) );
  OR2_X1 U11263 ( .A1(n15765), .A2(n15753), .ZN(n15746) );
  OR2_X2 U11264 ( .A1(n15472), .A2(n15473), .ZN(n15448) );
  OAI21_X1 U11265 ( .B1(n15453), .B2(n15451), .A(n15449), .ZN(n15440) );
  NOR2_X1 U11266 ( .A1(n15533), .A2(n11704), .ZN(n16257) );
  NAND2_X1 U11267 ( .A1(n14359), .A2(n14358), .ZN(n14360) );
  NAND2_X1 U11268 ( .A1(n15259), .A2(n15258), .ZN(n15257) );
  CLKBUF_X2 U11269 ( .A(n14964), .Z(n9671) );
  NAND2_X1 U11270 ( .A1(n11831), .A2(n11830), .ZN(n15553) );
  NAND2_X1 U11271 ( .A1(n9916), .A2(n10090), .ZN(n9865) );
  INV_X1 U11272 ( .A(n17300), .ZN(n17296) );
  NAND2_X1 U11273 ( .A1(n9816), .A2(n10629), .ZN(n14004) );
  AOI21_X1 U11274 ( .B1(n12238), .B2(n12237), .A(n10042), .ZN(n10041) );
  AND2_X1 U11275 ( .A1(n12550), .A2(n14200), .ZN(n15567) );
  OAI21_X1 U11276 ( .B1(n9918), .B2(n10090), .A(n10088), .ZN(n9917) );
  AND2_X1 U11277 ( .A1(n14318), .A2(n14335), .ZN(n14319) );
  AND2_X1 U11278 ( .A1(n14032), .A2(n12236), .ZN(n12237) );
  NAND2_X1 U11279 ( .A1(n10098), .A2(n15417), .ZN(n10097) );
  AND2_X1 U11280 ( .A1(n15024), .A2(n15023), .ZN(n9832) );
  NAND2_X1 U11281 ( .A1(n9811), .A2(n10119), .ZN(n13690) );
  NOR2_X1 U11282 ( .A1(n12223), .A2(n9839), .ZN(n9838) );
  NAND2_X1 U11283 ( .A1(n9775), .A2(n9717), .ZN(n14031) );
  INV_X1 U11284 ( .A(n13530), .ZN(n9811) );
  NAND2_X1 U11285 ( .A1(n12690), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10020) );
  OR2_X1 U11286 ( .A1(n16038), .A2(n12235), .ZN(n14983) );
  AND2_X1 U11287 ( .A1(n9810), .A2(n9809), .ZN(n11681) );
  XNOR2_X1 U11288 ( .A(n11823), .B(n11790), .ZN(n16287) );
  OAI21_X1 U11289 ( .B1(n11823), .B2(n15461), .A(n16336), .ZN(n16285) );
  AND2_X1 U11290 ( .A1(n11814), .A2(n13598), .ZN(n13780) );
  OR3_X2 U11291 ( .A1(n17627), .A2(n17610), .A3(n17631), .ZN(n12690) );
  AND2_X1 U11292 ( .A1(n11621), .A2(n11822), .ZN(n11819) );
  NAND2_X1 U11293 ( .A1(n12229), .A2(n14995), .ZN(n9776) );
  NOR2_X2 U11294 ( .A1(n9695), .A2(n12872), .ZN(n15267) );
  NOR2_X2 U11295 ( .A1(n13618), .A2(n13617), .ZN(n13668) );
  NAND2_X1 U11296 ( .A1(n17626), .A2(n12688), .ZN(n17611) );
  NAND2_X1 U11297 ( .A1(n13513), .A2(n13512), .ZN(n13618) );
  XNOR2_X1 U11298 ( .A(n11191), .B(n14489), .ZN(n14517) );
  AND2_X1 U11299 ( .A1(n9782), .A2(n11587), .ZN(n11659) );
  OAI22_X1 U11300 ( .A1(n14488), .A2(n11155), .B1(n11188), .B2(n11187), .ZN(
        n11191) );
  NOR2_X1 U11301 ( .A1(n13849), .A2(n13848), .ZN(n13893) );
  INV_X1 U11302 ( .A(n10551), .ZN(n10529) );
  AND4_X1 U11303 ( .A1(n11525), .A2(n11524), .A3(n11523), .A4(n11522), .ZN(
        n11526) );
  NAND4_X1 U11304 ( .A1(n10075), .A2(n10072), .A3(n10071), .A4(n10070), .ZN(
        n10069) );
  NOR2_X1 U11305 ( .A1(n17761), .A2(n12680), .ZN(n12683) );
  OAI22_X1 U11306 ( .A1(n19245), .A2(n19259), .B1(n11495), .B2(n12360), .ZN(
        n11500) );
  NAND2_X1 U11307 ( .A1(n9955), .A2(n9954), .ZN(n11757) );
  AND3_X1 U11308 ( .A1(n11550), .A2(n10079), .A3(n10078), .ZN(n9685) );
  AND2_X1 U11309 ( .A1(n10074), .A2(n10073), .ZN(n10072) );
  NAND2_X1 U11310 ( .A1(n11562), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10071) );
  NAND2_X1 U11311 ( .A1(n11572), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10070) );
  AND4_X1 U11312 ( .A1(n11514), .A2(n11513), .A3(n11512), .A4(n19989), .ZN(
        n11525) );
  AND2_X1 U11313 ( .A1(n12678), .A2(n12677), .ZN(n17771) );
  OR2_X1 U11314 ( .A1(n10910), .A2(n14561), .ZN(n10931) );
  INV_X1 U11315 ( .A(n11743), .ZN(n9955) );
  NOR2_X2 U11316 ( .A1(n13897), .A2(n13898), .ZN(n15220) );
  NOR2_X1 U11317 ( .A1(n13787), .A2(n12531), .ZN(n16311) );
  INV_X1 U11318 ( .A(n10475), .ZN(n10473) );
  AND2_X1 U11319 ( .A1(n11501), .A2(n11508), .ZN(n19338) );
  CLKBUF_X1 U11320 ( .A(n13474), .Z(n9677) );
  NAND2_X1 U11321 ( .A1(n17794), .A2(n17708), .ZN(n17827) );
  NAND3_X1 U11322 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(n15877), .ZN(n17127) );
  NOR2_X1 U11323 ( .A1(n15992), .A2(n17438), .ZN(n17409) );
  NOR2_X2 U11324 ( .A1(n11082), .A2(n20238), .ZN(n11080) );
  NOR2_X1 U11325 ( .A1(n10017), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10016) );
  AOI21_X1 U11326 ( .B1(n13123), .B2(n13122), .A(n13121), .ZN(n13521) );
  INV_X1 U11327 ( .A(n11729), .ZN(n11713) );
  NOR2_X2 U11328 ( .A1(n15987), .A2(n18200), .ZN(n18750) );
  NAND2_X1 U11329 ( .A1(n10454), .A2(n10342), .ZN(n13415) );
  NAND2_X1 U11330 ( .A1(n10045), .A2(n9684), .ZN(n20326) );
  AND2_X1 U11331 ( .A1(n13323), .A2(n20000), .ZN(n13340) );
  OR2_X1 U11332 ( .A1(n10421), .A2(n10420), .ZN(n10422) );
  AND2_X1 U11333 ( .A1(n15823), .A2(n11515), .ZN(n11520) );
  NAND2_X1 U11334 ( .A1(n12972), .A2(n12971), .ZN(n15826) );
  NAND2_X1 U11335 ( .A1(n10398), .A2(n10397), .ZN(n10421) );
  INV_X1 U11336 ( .A(n15823), .ZN(n19138) );
  INV_X2 U11337 ( .A(n18738), .ZN(n18128) );
  INV_X2 U11338 ( .A(n17282), .ZN(n17274) );
  NOR2_X1 U11339 ( .A1(n15888), .A2(n15886), .ZN(n12126) );
  NAND2_X1 U11340 ( .A1(n10458), .A2(n10457), .ZN(n20401) );
  NAND2_X1 U11341 ( .A1(n10014), .A2(n10013), .ZN(n17875) );
  NOR2_X2 U11342 ( .A1(n18945), .A2(n16555), .ZN(n15888) );
  OR2_X2 U11343 ( .A1(n17483), .A2(n18775), .ZN(n17551) );
  AND2_X1 U11344 ( .A1(n15987), .A2(n17485), .ZN(n15886) );
  AND2_X1 U11345 ( .A1(n13304), .A2(n13303), .ZN(n13471) );
  NAND2_X1 U11346 ( .A1(n11452), .A2(n11408), .ZN(n11466) );
  NAND2_X2 U11347 ( .A1(n16437), .A2(n12674), .ZN(n17815) );
  AND2_X1 U11348 ( .A1(n9927), .A2(n9926), .ZN(n13304) );
  AOI211_X1 U11349 ( .C1(n15905), .C2(n15992), .A(n12720), .B(n12719), .ZN(
        n15891) );
  NOR4_X2 U11350 ( .A1(n14066), .A2(n12720), .A3(n12110), .A4(n12112), .ZN(
        n17485) );
  AOI21_X1 U11351 ( .B1(n10442), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10110), 
        .ZN(n10109) );
  NOR2_X1 U11352 ( .A1(n17429), .A2(n12660), .ZN(n12664) );
  OR2_X1 U11353 ( .A1(n17291), .A2(n18267), .ZN(n12120) );
  INV_X1 U11354 ( .A(n11406), .ZN(n12524) );
  INV_X1 U11355 ( .A(n18281), .ZN(n15905) );
  NOR2_X1 U11356 ( .A1(n11664), .A2(n11658), .ZN(n9942) );
  NAND2_X1 U11357 ( .A1(n11429), .A2(n16386), .ZN(n11858) );
  AND2_X1 U11358 ( .A1(n17562), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11996) );
  AND2_X1 U11359 ( .A1(n19971), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11429) );
  INV_X1 U11360 ( .A(n11673), .ZN(n9943) );
  NAND2_X1 U11361 ( .A1(n12516), .A2(n11405), .ZN(n12273) );
  AND2_X1 U11362 ( .A1(n11966), .A2(n12525), .ZN(n12514) );
  OR2_X1 U11363 ( .A1(n11042), .A2(n10392), .ZN(n10395) );
  NAND3_X1 U11364 ( .A1(n9854), .A2(n9853), .A3(n12978), .ZN(n11406) );
  NOR2_X2 U11365 ( .A1(n11999), .A2(n17606), .ZN(n17562) );
  INV_X1 U11366 ( .A(n11387), .ZN(n12516) );
  NAND2_X1 U11367 ( .A1(n11386), .A2(n11385), .ZN(n9854) );
  BUF_X2 U11368 ( .A(n12315), .Z(n12503) );
  AND2_X1 U11369 ( .A1(n13310), .A2(n13632), .ZN(n14484) );
  NOR2_X1 U11370 ( .A1(n20267), .A2(n20263), .ZN(n13165) );
  NAND2_X1 U11371 ( .A1(n9634), .A2(n11389), .ZN(n12266) );
  INV_X2 U11372 ( .A(n14492), .ZN(n9636) );
  OR2_X1 U11373 ( .A1(n11275), .A2(n11274), .ZN(n11547) );
  AND2_X1 U11374 ( .A1(n11545), .A2(n11544), .ZN(n12302) );
  NOR2_X2 U11375 ( .A1(n19989), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12974) );
  AND2_X1 U11376 ( .A1(n12595), .A2(n12594), .ZN(n17429) );
  OR2_X1 U11377 ( .A1(n11302), .A2(n11301), .ZN(n12319) );
  NAND2_X1 U11378 ( .A1(n13329), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10460) );
  NAND3_X1 U11379 ( .A1(n10177), .A2(n12620), .A3(n10156), .ZN(n12725) );
  INV_X1 U11380 ( .A(n11305), .ZN(n14355) );
  OR2_X1 U11381 ( .A1(n13632), .A2(n20258), .ZN(n13246) );
  INV_X1 U11382 ( .A(n13315), .ZN(n20263) );
  AND2_X1 U11383 ( .A1(n12606), .A2(n10010), .ZN(n10009) );
  OR2_X1 U11384 ( .A1(n10376), .A2(n10375), .ZN(n12219) );
  NAND2_X1 U11385 ( .A1(n12969), .A2(n11398), .ZN(n13264) );
  CLKBUF_X1 U11386 ( .A(n12969), .Z(n19279) );
  OR2_X1 U11387 ( .A1(n10388), .A2(n10387), .ZN(n12157) );
  OR2_X2 U11388 ( .A1(n16500), .A2(n16453), .ZN(n16503) );
  OR2_X1 U11389 ( .A1(n11616), .A2(n11615), .ZN(n12332) );
  AND4_X2 U11390 ( .A1(n10279), .A2(n10278), .A3(n10277), .A4(n10276), .ZN(
        n13632) );
  NAND2_X2 U11391 ( .A1(n11354), .A2(n11353), .ZN(n12969) );
  NAND2_X1 U11392 ( .A1(n11366), .A2(n11365), .ZN(n11398) );
  AND4_X1 U11393 ( .A1(n12648), .A2(n12647), .A3(n12646), .A4(n12645), .ZN(
        n12656) );
  BUF_X2 U11394 ( .A(n10300), .Z(n13329) );
  NAND2_X2 U11395 ( .A1(n10182), .A2(n10180), .ZN(n20289) );
  AND4_X1 U11396 ( .A1(n10254), .A2(n10253), .A3(n10252), .A4(n10251), .ZN(
        n10255) );
  AND4_X1 U11397 ( .A1(n10293), .A2(n10292), .A3(n10291), .A4(n10290), .ZN(
        n10294) );
  AND4_X1 U11398 ( .A1(n10284), .A2(n10283), .A3(n10282), .A4(n10281), .ZN(
        n10296) );
  AND4_X1 U11399 ( .A1(n10267), .A2(n10266), .A3(n10265), .A4(n10264), .ZN(
        n10278) );
  AND4_X1 U11400 ( .A1(n10263), .A2(n10262), .A3(n10261), .A4(n10260), .ZN(
        n10279) );
  NAND4_X2 U11401 ( .A1(n10234), .A2(n10233), .A3(n10232), .A4(n10231), .ZN(
        n14160) );
  INV_X2 U11402 ( .A(U214), .ZN(n16500) );
  NOR2_X2 U11403 ( .A1(n18345), .A2(n18508), .ZN(n18304) );
  NAND2_X1 U11404 ( .A1(n11322), .A2(n16338), .ZN(n11329) );
  AND4_X1 U11405 ( .A1(n10275), .A2(n10274), .A3(n10273), .A4(n10272), .ZN(
        n10276) );
  AND4_X1 U11406 ( .A1(n10271), .A2(n10270), .A3(n10269), .A4(n10268), .ZN(
        n10277) );
  AND4_X1 U11407 ( .A1(n10288), .A2(n10287), .A3(n10286), .A4(n10285), .ZN(
        n10295) );
  AND4_X1 U11408 ( .A1(n10230), .A2(n10229), .A3(n10228), .A4(n10227), .ZN(
        n10231) );
  AND4_X1 U11409 ( .A1(n10226), .A2(n10225), .A3(n10224), .A4(n10223), .ZN(
        n10232) );
  AND4_X1 U11411 ( .A1(n10222), .A2(n10221), .A3(n10220), .A4(n10219), .ZN(
        n10233) );
  AND4_X1 U11412 ( .A1(n10218), .A2(n10217), .A3(n10216), .A4(n10215), .ZN(
        n10234) );
  AND4_X1 U11413 ( .A1(n10214), .A2(n10213), .A3(n10212), .A4(n10211), .ZN(
        n9680) );
  AND4_X1 U11414 ( .A1(n10197), .A2(n10196), .A3(n10195), .A4(n10194), .ZN(
        n10180) );
  AND4_X1 U11415 ( .A1(n10201), .A2(n10200), .A3(n10199), .A4(n10198), .ZN(
        n9709) );
  INV_X1 U11416 ( .A(n12644), .ZN(n17184) );
  AND2_X1 U11417 ( .A1(n11310), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9857) );
  INV_X2 U11418 ( .A(n12033), .ZN(n17209) );
  AND2_X1 U11419 ( .A1(n11316), .A2(n16338), .ZN(n9859) );
  INV_X2 U11420 ( .A(n9631), .ZN(n17227) );
  INV_X2 U11421 ( .A(n11539), .ZN(n14294) );
  BUF_X1 U11422 ( .A(n10289), .Z(n9670) );
  AND2_X2 U11423 ( .A1(n14417), .A2(n16338), .ZN(n14308) );
  NAND2_X2 U11424 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19918), .ZN(n19916) );
  AOI22_X1 U11425 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10212) );
  INV_X2 U11426 ( .A(n12086), .ZN(n17101) );
  NOR2_X1 U11427 ( .A1(n12020), .A2(n16926), .ZN(n12643) );
  NAND2_X1 U11428 ( .A1(n12018), .A2(n12014), .ZN(n17205) );
  OR2_X2 U11429 ( .A1(n16926), .A2(n10024), .ZN(n12562) );
  NAND3_X1 U11430 ( .A1(n18912), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n18712), .ZN(n12033) );
  OR2_X2 U11431 ( .A1(n18728), .A2(n12021), .ZN(n17099) );
  NAND2_X2 U11432 ( .A1(n18870), .A2(n18809), .ZN(n18862) );
  AND2_X2 U11433 ( .A1(n9651), .A2(n16338), .ZN(n14293) );
  NAND2_X2 U11434 ( .A1(n18870), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18873) );
  INV_X2 U11435 ( .A(n16543), .ZN(n16545) );
  NOR2_X1 U11436 ( .A1(n15684), .A2(n15501), .ZN(n11835) );
  NAND2_X1 U11437 ( .A1(n12022), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12019) );
  NAND3_X1 U11438 ( .A1(n12023), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12017) );
  NAND4_X2 U11439 ( .A1(n12023), .A2(n18897), .A3(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A4(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n17167) );
  NAND2_X1 U11440 ( .A1(n12014), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12021) );
  AND2_X1 U11441 ( .A1(n10184), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13425) );
  BUF_X4 U11442 ( .A(n14271), .Z(n9637) );
  AND2_X2 U11443 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13429) );
  NOR2_X1 U11444 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10141) );
  AND2_X2 U11445 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15163) );
  AND2_X1 U11446 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13431) );
  NAND2_X1 U11447 ( .A1(n12684), .A2(n12683), .ZN(n17709) );
  NAND2_X1 U11448 ( .A1(n17728), .A2(n16442), .ZN(n12684) );
  NAND2_X1 U11449 ( .A1(n11792), .A2(n9707), .ZN(n11770) );
  OR2_X2 U11450 ( .A1(n11775), .A2(n11774), .ZN(n11786) );
  NOR2_X1 U11451 ( .A1(n15532), .A2(n9638), .ZN(n15488) );
  NAND2_X1 U11452 ( .A1(n11833), .A2(n11835), .ZN(n9638) );
  XNOR2_X1 U11453 ( .A(n11475), .B(n11476), .ZN(n9639) );
  XNOR2_X1 U11454 ( .A(n11475), .B(n11476), .ZN(n11474) );
  NOR3_X2 U11455 ( .A1(n18294), .A2(n15905), .A3(n14064), .ZN(n14065) );
  NAND3_X2 U11456 ( .A1(n10087), .A2(n11850), .A3(n10086), .ZN(n10029) );
  OAI21_X1 U11457 ( .B1(n9919), .B2(n10090), .A(n9916), .ZN(n9641) );
  CLKBUF_X1 U11458 ( .A(n13776), .Z(n9642) );
  OAI21_X1 U11459 ( .B1(n9919), .B2(n10090), .A(n9916), .ZN(n15794) );
  NAND2_X2 U11460 ( .A1(n13668), .A2(n13667), .ZN(n13708) );
  INV_X2 U11461 ( .A(n11853), .ZN(n10087) );
  INV_X1 U11462 ( .A(n14969), .ZN(n9643) );
  OAI22_X1 U11463 ( .A1(n15154), .A2(n12176), .B1(n13246), .B2(n12175), .ZN(
        n9644) );
  INV_X1 U11464 ( .A(n10415), .ZN(n9645) );
  NAND2_X1 U11465 ( .A1(n14056), .A2(n12226), .ZN(n14009) );
  OAI22_X1 U11466 ( .A1(n15154), .A2(n12176), .B1(n13246), .B2(n12175), .ZN(
        n12177) );
  NAND2_X1 U11467 ( .A1(n11062), .A2(n13310), .ZN(n13176) );
  NAND2_X1 U11468 ( .A1(n13176), .A2(n11065), .ZN(n13325) );
  NOR2_X1 U11469 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9824) );
  AND3_X4 U11471 ( .A1(n11223), .A2(n13763), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14440) );
  OAI21_X2 U11473 ( .B1(n13487), .B2(n10034), .A(n11808), .ZN(n11810) );
  NAND2_X2 U11474 ( .A1(n13927), .A2(n13928), .ZN(n9919) );
  AND2_X1 U11475 ( .A1(n11504), .A2(n11496), .ZN(n11563) );
  AND2_X2 U11476 ( .A1(n11497), .A2(n9895), .ZN(n11554) );
  AND2_X4 U11477 ( .A1(n12974), .A2(n12296), .ZN(n12314) );
  AND2_X2 U11478 ( .A1(n10189), .A2(n13425), .ZN(n10963) );
  INV_X1 U11479 ( .A(n11330), .ZN(n9647) );
  NAND2_X4 U11481 ( .A1(n9705), .A2(n9680), .ZN(n20280) );
  NOR2_X2 U11482 ( .A1(n12764), .A2(n15399), .ZN(n12765) );
  BUF_X2 U11483 ( .A(n18291), .Z(n9649) );
  OR2_X1 U11484 ( .A1(n12247), .A2(n11099), .ZN(n13336) );
  AND4_X2 U11485 ( .A1(n10210), .A2(n10209), .A3(n10208), .A4(n10207), .ZN(
        n9705) );
  AND2_X1 U11486 ( .A1(n10193), .A2(n15163), .ZN(n9650) );
  OAI21_X2 U11488 ( .B1(n12980), .B2(n13183), .A(n13324), .ZN(n10103) );
  AND3_X1 U11489 ( .A1(n14484), .A2(n10304), .A3(n13165), .ZN(n13330) );
  AOI211_X2 U11490 ( .C1(n16306), .C2(n15404), .A(n15403), .B(n15402), .ZN(
        n15405) );
  XNOR2_X1 U11491 ( .A(n11680), .B(n13789), .ZN(n13775) );
  AOI22_X2 U11492 ( .A1(n13595), .A2(n13596), .B1(n11679), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13776) );
  AND2_X2 U11493 ( .A1(n15829), .A2(n11223), .ZN(n9651) );
  NOR2_X2 U11494 ( .A1(n14883), .A2(n12242), .ZN(n14875) );
  NAND2_X1 U11495 ( .A1(n10306), .A2(n20267), .ZN(n10259) );
  BUF_X4 U11496 ( .A(n9636), .Z(n9658) );
  XNOR2_X1 U11497 ( .A(n10314), .B(n10328), .ZN(n20366) );
  AND2_X1 U11498 ( .A1(n10356), .A2(n20271), .ZN(n11046) );
  XOR2_X1 U11499 ( .A(n14151), .B(n14150), .Z(n15042) );
  INV_X1 U11500 ( .A(n14440), .ZN(n9660) );
  INV_X1 U11501 ( .A(n9660), .ZN(n9661) );
  NOR2_X1 U11505 ( .A1(n14858), .A2(n14857), .ZN(n9778) );
  NAND2_X1 U11506 ( .A1(n14875), .A2(n15045), .ZN(n14858) );
  NAND2_X1 U11507 ( .A1(n10040), .A2(n10041), .ZN(n16082) );
  INV_X1 U11508 ( .A(n13476), .ZN(n10418) );
  NAND2_X1 U11509 ( .A1(n14160), .A2(n10300), .ZN(n12247) );
  INV_X2 U11510 ( .A(n20280), .ZN(n10318) );
  NOR2_X2 U11511 ( .A1(n11507), .A2(n15859), .ZN(n11566) );
  AND2_X2 U11512 ( .A1(n10193), .A2(n15163), .ZN(n9666) );
  AND2_X1 U11513 ( .A1(n10189), .A2(n10191), .ZN(n9675) );
  XNOR2_X1 U11514 ( .A(n12171), .B(n20204), .ZN(n13293) );
  NAND2_X2 U11515 ( .A1(n10338), .A2(n10339), .ZN(n10454) );
  NAND2_X2 U11516 ( .A1(n16064), .A2(n12212), .ZN(n9840) );
  NAND2_X1 U11517 ( .A1(n20366), .A2(n10413), .ZN(n10416) );
  AND2_X2 U11518 ( .A1(n14660), .A2(n14662), .ZN(n14648) );
  NOR2_X2 U11519 ( .A1(n14673), .A2(n14674), .ZN(n14660) );
  OAI21_X2 U11520 ( .B1(n9840), .B2(n9700), .A(n9836), .ZN(n14056) );
  OAI21_X2 U11521 ( .B1(n18714), .B2(n18727), .A(n18713), .ZN(n18738) );
  NAND2_X1 U11522 ( .A1(n20221), .A2(n12165), .ZN(n12171) );
  NAND3_X2 U11523 ( .A1(n10259), .A2(n10258), .A3(n10297), .ZN(n10307) );
  OAI21_X2 U11524 ( .B1(n9671), .B2(n9768), .A(n12224), .ZN(n14923) );
  XNOR2_X1 U11525 ( .A(n9777), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15032) );
  NOR2_X4 U11526 ( .A1(n10303), .A2(n12245), .ZN(n13177) );
  NAND2_X2 U11527 ( .A1(n10302), .A2(n10305), .ZN(n12245) );
  NAND2_X2 U11528 ( .A1(n10235), .A2(n13163), .ZN(n10306) );
  NAND2_X2 U11529 ( .A1(n10328), .A2(n10100), .ZN(n10332) );
  AND2_X1 U11530 ( .A1(n10193), .A2(n10190), .ZN(n9667) );
  AND2_X1 U11531 ( .A1(n10189), .A2(n13431), .ZN(n9669) );
  NAND2_X2 U11532 ( .A1(n10507), .A2(n10476), .ZN(n15154) );
  NAND2_X1 U11533 ( .A1(n12218), .A2(n12217), .ZN(n9672) );
  NAND2_X1 U11534 ( .A1(n12218), .A2(n12217), .ZN(n9673) );
  AND2_X4 U11535 ( .A1(n10189), .A2(n10193), .ZN(n10979) );
  NOR2_X2 U11536 ( .A1(n10307), .A2(n10280), .ZN(n11062) );
  OR2_X1 U11537 ( .A1(n9671), .A2(n9766), .ZN(n14931) );
  AND2_X1 U11538 ( .A1(n10189), .A2(n10191), .ZN(n10370) );
  NOR2_X4 U11539 ( .A1(n13690), .A2(n13742), .ZN(n13743) );
  NAND2_X1 U11540 ( .A1(n9919), .A2(n9916), .ZN(n9866) );
  AOI21_X1 U11541 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19938), .A(
        n11202), .ZN(n11211) );
  NOR2_X1 U11542 ( .A1(n11207), .A2(n11201), .ZN(n11202) );
  NAND2_X1 U11543 ( .A1(n11064), .A2(n11063), .ZN(n13193) );
  NOR2_X1 U11544 ( .A1(n12805), .A2(n12804), .ZN(n14170) );
  INV_X1 U11545 ( .A(n13565), .ZN(n9960) );
  NAND2_X1 U11546 ( .A1(n11387), .A2(n12978), .ZN(n9853) );
  NAND2_X1 U11547 ( .A1(n9781), .A2(n10508), .ZN(n10551) );
  AND2_X1 U11548 ( .A1(n10412), .A2(n10411), .ZN(n10419) );
  OR2_X1 U11549 ( .A1(n11042), .A2(n10410), .ZN(n10411) );
  OAI21_X1 U11550 ( .B1(n10445), .B2(n10111), .A(n10109), .ZN(n10398) );
  AND2_X1 U11551 ( .A1(n11619), .A2(n11659), .ZN(n10095) );
  NAND2_X1 U11552 ( .A1(n19265), .A2(n12266), .ZN(n11420) );
  NOR2_X1 U11553 ( .A1(n17422), .A2(n12667), .ZN(n12672) );
  AND2_X1 U11554 ( .A1(n10179), .A2(n14596), .ZN(n10123) );
  INV_X1 U11555 ( .A(n14626), .ZN(n10120) );
  AND2_X1 U11556 ( .A1(n10566), .A2(n10580), .ZN(n10119) );
  INV_X1 U11557 ( .A(n13693), .ZN(n10580) );
  NOR2_X1 U11558 ( .A1(n9949), .A2(n9751), .ZN(n9948) );
  INV_X1 U11559 ( .A(n9697), .ZN(n9795) );
  NAND2_X1 U11560 ( .A1(n15431), .A2(n15619), .ZN(n9878) );
  OAI21_X1 U11561 ( .B1(n15431), .B2(n15619), .A(n11765), .ZN(n9879) );
  NAND2_X1 U11562 ( .A1(n10065), .A2(n15290), .ZN(n10064) );
  INV_X1 U11563 ( .A(n15306), .ZN(n10065) );
  AND2_X1 U11564 ( .A1(n9737), .A2(n12859), .ZN(n9964) );
  INV_X1 U11565 ( .A(n9917), .ZN(n9916) );
  AOI21_X1 U11566 ( .B1(n10092), .B2(n10089), .A(n9728), .ZN(n10088) );
  INV_X1 U11567 ( .A(n11693), .ZN(n10089) );
  NOR2_X1 U11568 ( .A1(n13585), .A2(n9968), .ZN(n9967) );
  INV_X1 U11569 ( .A(n13257), .ZN(n9968) );
  OR2_X1 U11570 ( .A1(n11287), .A2(n11286), .ZN(n12324) );
  INV_X2 U11571 ( .A(n11873), .ZN(n11957) );
  NAND2_X1 U11573 ( .A1(n11228), .A2(n11229), .ZN(n9970) );
  AND4_X1 U11574 ( .A1(n11227), .A2(n11226), .A3(n11225), .A4(n16338), .ZN(
        n11228) );
  NAND2_X1 U11575 ( .A1(n11234), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9969) );
  AND4_X1 U11576 ( .A1(n11233), .A2(n11232), .A3(n11231), .A4(n11230), .ZN(
        n11234) );
  NAND2_X1 U11577 ( .A1(n11347), .A2(n16338), .ZN(n11354) );
  OAI22_X1 U11578 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15903), .B1(
        n11212), .B2(n11211), .ZN(n11984) );
  NAND2_X1 U11579 ( .A1(n17594), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11999) );
  NOR2_X1 U11580 ( .A1(n15991), .A2(n12111), .ZN(n15893) );
  NOR2_X1 U11581 ( .A1(n9734), .A2(n9818), .ZN(n9817) );
  INV_X1 U11582 ( .A(n14546), .ZN(n9818) );
  AND2_X2 U11583 ( .A1(n11054), .A2(n11053), .ZN(n14483) );
  INV_X1 U11584 ( .A(n11858), .ZN(n11873) );
  INV_X1 U11585 ( .A(n11790), .ZN(n15461) );
  AND2_X1 U11586 ( .A1(n9973), .A2(n15336), .ZN(n9971) );
  NOR2_X1 U11587 ( .A1(n9974), .A2(n9764), .ZN(n9973) );
  NOR2_X1 U11588 ( .A1(n9902), .A2(n9899), .ZN(n9898) );
  OAI21_X1 U11589 ( .B1(n9901), .B2(n9899), .A(n9897), .ZN(n9896) );
  NAND2_X1 U11590 ( .A1(n9646), .A2(n9908), .ZN(n9904) );
  NAND2_X1 U11591 ( .A1(n9646), .A2(n15777), .ZN(n9912) );
  AND2_X1 U11592 ( .A1(n13784), .A2(n9960), .ZN(n9959) );
  NOR2_X1 U11593 ( .A1(n19934), .A2(n19961), .ZN(n19606) );
  INV_X1 U11594 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19987) );
  OR2_X1 U11595 ( .A1(n14457), .A2(n19137), .ZN(n12829) );
  NAND2_X1 U11596 ( .A1(n19250), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10082) );
  NAND2_X1 U11597 ( .A1(n11565), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10081) );
  NAND2_X1 U11598 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10080) );
  NAND2_X1 U11599 ( .A1(n11553), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10078) );
  AND2_X1 U11600 ( .A1(n19966), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11204) );
  NOR2_X1 U11601 ( .A1(n11015), .A2(n11016), .ZN(n11014) );
  NAND2_X1 U11602 ( .A1(n10498), .A2(n10497), .ZN(n10508) );
  OR2_X1 U11603 ( .A1(n11042), .A2(n10486), .ZN(n10498) );
  NAND2_X1 U11604 ( .A1(n13336), .A2(n10308), .ZN(n10102) );
  AOI21_X1 U11605 ( .B1(n20645), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11014), .ZN(n11013) );
  AND4_X1 U11606 ( .A1(n11638), .A2(n11637), .A3(n11636), .A4(n11635), .ZN(
        n11644) );
  INV_X1 U11607 ( .A(n12332), .ZN(n11647) );
  AND4_X1 U11608 ( .A1(n11592), .A2(n11591), .A3(n11590), .A4(n11589), .ZN(
        n11606) );
  NAND2_X1 U11609 ( .A1(n9681), .A2(n9713), .ZN(n9782) );
  INV_X1 U11610 ( .A(n15408), .ZN(n10098) );
  NAND2_X1 U11611 ( .A1(n9854), .A2(n9853), .ZN(n11395) );
  NAND2_X1 U11612 ( .A1(n11200), .A2(n11199), .ZN(n11207) );
  NAND2_X1 U11613 ( .A1(n10256), .A2(n13315), .ZN(n9772) );
  INV_X1 U11614 ( .A(n11001), .ZN(n10970) );
  OR2_X1 U11615 ( .A1(n10306), .A2(n20914), .ZN(n11001) );
  NAND2_X1 U11616 ( .A1(n10116), .A2(n10115), .ZN(n10114) );
  INV_X1 U11617 ( .A(n10117), .ZN(n10116) );
  INV_X1 U11618 ( .A(n14690), .ZN(n10115) );
  INV_X1 U11619 ( .A(n14491), .ZN(n11176) );
  NOR2_X1 U11620 ( .A1(n10555), .A2(n10554), .ZN(n10556) );
  INV_X1 U11621 ( .A(n10552), .ZN(n10555) );
  INV_X1 U11622 ( .A(n13746), .ZN(n9925) );
  NAND2_X1 U11623 ( .A1(n9658), .A2(n11155), .ZN(n11175) );
  NAND2_X1 U11624 ( .A1(n11113), .A2(n9922), .ZN(n9921) );
  INV_X1 U11625 ( .A(n13367), .ZN(n11113) );
  INV_X1 U11626 ( .A(n13380), .ZN(n9922) );
  NAND2_X1 U11627 ( .A1(n10337), .A2(n10336), .ZN(n10339) );
  OAI21_X1 U11628 ( .B1(n15967), .B2(n13447), .A(n15187), .ZN(n20243) );
  OR3_X1 U11629 ( .A1(n9945), .A2(n11653), .A3(n9940), .ZN(n11661) );
  NAND2_X1 U11630 ( .A1(n9943), .A2(n9944), .ZN(n9940) );
  NAND2_X1 U11631 ( .A1(n9655), .A2(n16338), .ZN(n12408) );
  INV_X1 U11632 ( .A(n14395), .ZN(n10132) );
  NAND2_X1 U11633 ( .A1(n10143), .A2(n13846), .ZN(n10142) );
  INV_X1 U11634 ( .A(n10145), .ZN(n10143) );
  AND2_X1 U11635 ( .A1(n19989), .A2(n13041), .ZN(n14393) );
  NOR2_X1 U11636 ( .A1(n12551), .A2(n14198), .ZN(n10057) );
  NOR2_X1 U11637 ( .A1(n10062), .A2(n10061), .ZN(n10060) );
  INV_X1 U11638 ( .A(n15211), .ZN(n10061) );
  INV_X1 U11639 ( .A(n15266), .ZN(n10062) );
  NAND2_X1 U11640 ( .A1(n9999), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9998) );
  INV_X1 U11641 ( .A(n10000), .ZN(n9999) );
  NOR2_X1 U11642 ( .A1(n10053), .A2(n13203), .ZN(n10052) );
  INV_X1 U11643 ( .A(n10054), .ZN(n10053) );
  INV_X1 U11644 ( .A(n9876), .ZN(n9875) );
  OAI21_X1 U11645 ( .B1(n11780), .B2(n9795), .A(n12260), .ZN(n9876) );
  NAND2_X1 U11646 ( .A1(n9975), .A2(n12882), .ZN(n9974) );
  INV_X1 U11647 ( .A(n15189), .ZN(n9975) );
  NOR2_X1 U11648 ( .A1(n9794), .A2(n9796), .ZN(n9793) );
  NOR2_X1 U11649 ( .A1(n9952), .A2(n9795), .ZN(n9794) );
  NOR2_X1 U11650 ( .A1(n11746), .A2(n15802), .ZN(n9864) );
  NAND2_X1 U11651 ( .A1(n9862), .A2(n15795), .ZN(n9861) );
  INV_X1 U11652 ( .A(n11746), .ZN(n9862) );
  NOR2_X1 U11653 ( .A1(n15466), .A2(n11752), .ZN(n9956) );
  NOR2_X1 U11654 ( .A1(n13684), .A2(n13712), .ZN(n10068) );
  INV_X1 U11655 ( .A(n15539), .ZN(n9899) );
  INV_X1 U11656 ( .A(n15747), .ZN(n9965) );
  NOR2_X1 U11657 ( .A1(n9911), .A2(n15779), .ZN(n9910) );
  INV_X1 U11658 ( .A(n15760), .ZN(n9911) );
  NAND2_X1 U11659 ( .A1(n11421), .A2(n11420), .ZN(n11422) );
  NAND2_X1 U11660 ( .A1(n11419), .A2(n11418), .ZN(n11421) );
  AND2_X1 U11661 ( .A1(n13115), .A2(n11496), .ZN(n11508) );
  NOR2_X1 U11662 ( .A1(n12295), .A2(n12969), .ZN(n11400) );
  OAI211_X1 U11663 ( .C1(n17241), .C2(n9849), .A(n9848), .B(n9847), .ZN(n9846)
         );
  INV_X1 U11664 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n9849) );
  NAND2_X1 U11665 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n9847) );
  NAND2_X1 U11666 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n9848) );
  INV_X1 U11667 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17207) );
  NOR3_X1 U11668 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n12022), .ZN(n12018) );
  NAND2_X1 U11669 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12617) );
  NAND2_X1 U11670 ( .A1(n12616), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12618) );
  OR2_X1 U11671 ( .A1(n18714), .A2(n12717), .ZN(n14064) );
  NOR3_X1 U11672 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n12019), .ZN(n12601) );
  INV_X1 U11673 ( .A(n18286), .ZN(n12110) );
  OAI21_X1 U11674 ( .B1(n12137), .B2(n12708), .A(n12709), .ZN(n16553) );
  INV_X1 U11675 ( .A(n17794), .ZN(n12678) );
  AND2_X1 U11676 ( .A1(n12672), .A2(n12671), .ZN(n12674) );
  NAND2_X1 U11677 ( .A1(n17846), .A2(n9696), .ZN(n10026) );
  NAND2_X1 U11678 ( .A1(n10027), .A2(n9696), .ZN(n10025) );
  AND2_X1 U11679 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12665), .ZN(
        n12666) );
  XNOR2_X1 U11680 ( .A(n17445), .B(n17434), .ZN(n12658) );
  NOR3_X1 U11681 ( .A1(n12720), .A2(n15911), .A3(n18715), .ZN(n15896) );
  OR2_X1 U11682 ( .A1(n20916), .A2(n13630), .ZN(n14727) );
  NAND2_X1 U11683 ( .A1(n10104), .A2(n10617), .ZN(n10108) );
  NAND2_X1 U11684 ( .A1(n13743), .A2(n13825), .ZN(n10104) );
  AND2_X1 U11685 ( .A1(n10106), .A2(n13967), .ZN(n10105) );
  OR2_X1 U11686 ( .A1(n13825), .A2(n10107), .ZN(n10106) );
  XNOR2_X1 U11687 ( .A(n12255), .B(n12254), .ZN(n13641) );
  INV_X1 U11688 ( .A(n10905), .ZN(n11006) );
  OR2_X1 U11689 ( .A1(n10976), .A2(n10975), .ZN(n12253) );
  NOR2_X1 U11690 ( .A1(n10122), .A2(n14557), .ZN(n10121) );
  INV_X1 U11691 ( .A(n10123), .ZN(n10122) );
  NAND2_X1 U11692 ( .A1(n10814), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10876) );
  NAND2_X1 U11693 ( .A1(n14009), .A2(n12237), .ZN(n10040) );
  INV_X1 U11694 ( .A(n14963), .ZN(n10042) );
  INV_X1 U11695 ( .A(n14547), .ZN(n9935) );
  INV_X1 U11696 ( .A(n12213), .ZN(n9839) );
  OAI21_X1 U11697 ( .B1(n20326), .B2(n12176), .A(n12155), .ZN(n13061) );
  AND2_X1 U11698 ( .A1(n10393), .A2(n12215), .ZN(n10394) );
  NAND2_X1 U11699 ( .A1(n10475), .A2(n10425), .ZN(n20240) );
  INV_X1 U11700 ( .A(n12156), .ZN(n10435) );
  OR3_X1 U11701 ( .A1(n13194), .A2(n13193), .A3(n13192), .ZN(n15939) );
  CLKBUF_X1 U11702 ( .A(n13476), .Z(n20651) );
  NOR2_X1 U11703 ( .A1(n15154), .A2(n15155), .ZN(n20622) );
  OR2_X1 U11704 ( .A1(n9677), .A2(n20326), .ZN(n20698) );
  AND2_X1 U11705 ( .A1(n9677), .A2(n20326), .ZN(n20719) );
  OR2_X1 U11706 ( .A1(n20240), .A2(n15156), .ZN(n20778) );
  OR2_X1 U11707 ( .A1(n14483), .A2(n14472), .ZN(n15951) );
  INV_X1 U11708 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20645) );
  OR2_X1 U11709 ( .A1(n15205), .A2(n15425), .ZN(n9985) );
  NAND2_X1 U11710 ( .A1(n11744), .A2(n11757), .ZN(n18976) );
  AND2_X1 U11711 ( .A1(n19027), .A2(n19029), .ZN(n12791) );
  INV_X1 U11712 ( .A(n11728), .ZN(n11712) );
  NOR2_X1 U11713 ( .A1(n11734), .A2(n9949), .ZN(n11732) );
  NAND2_X1 U11714 ( .A1(n9947), .A2(n10172), .ZN(n11733) );
  NAND2_X1 U11715 ( .A1(n10032), .A2(n11486), .ZN(n11850) );
  NAND2_X1 U11716 ( .A1(n9639), .A2(n11485), .ZN(n10032) );
  OR3_X1 U11717 ( .A1(n10064), .A2(n10066), .A3(n12898), .ZN(n10063) );
  AND2_X1 U11718 ( .A1(n11934), .A2(n11933), .ZN(n12872) );
  NAND2_X1 U11719 ( .A1(n10125), .A2(n10131), .ZN(n10128) );
  INV_X1 U11720 ( .A(n10139), .ZN(n15274) );
  NAND2_X1 U11721 ( .A1(n13571), .A2(n13278), .ZN(n15783) );
  AND3_X1 U11722 ( .A1(n12354), .A2(n12353), .A3(n12352), .ZN(n13585) );
  NAND2_X1 U11723 ( .A1(n13261), .A2(n13260), .ZN(n13755) );
  INV_X1 U11724 ( .A(n19845), .ZN(n13262) );
  AND2_X1 U11725 ( .A1(n11944), .A2(n11943), .ZN(n15251) );
  NAND2_X1 U11726 ( .A1(n10048), .A2(n13665), .ZN(n10047) );
  INV_X1 U11727 ( .A(n13622), .ZN(n10048) );
  NAND2_X1 U11728 ( .A1(n12780), .A2(n10006), .ZN(n12789) );
  NOR2_X1 U11729 ( .A1(n10008), .A2(n9725), .ZN(n10006) );
  AND2_X1 U11730 ( .A1(n12780), .A2(n11842), .ZN(n12788) );
  INV_X1 U11731 ( .A(n10008), .ZN(n10007) );
  INV_X1 U11732 ( .A(n13782), .ZN(n11818) );
  INV_X1 U11733 ( .A(n11819), .ZN(n11817) );
  AOI21_X1 U11734 ( .B1(n10161), .B2(n13782), .A(n9726), .ZN(n9851) );
  AND2_X1 U11735 ( .A1(n11384), .A2(n11383), .ZN(n12283) );
  INV_X1 U11736 ( .A(n9783), .ZN(n9800) );
  AOI21_X1 U11737 ( .B1(n15420), .B2(n9793), .A(n9784), .ZN(n9783) );
  NAND2_X1 U11738 ( .A1(n9801), .A2(n9785), .ZN(n9784) );
  NAND2_X1 U11739 ( .A1(n9803), .A2(n12555), .ZN(n9801) );
  OAI21_X1 U11740 ( .B1(n15420), .B2(n9795), .A(n9793), .ZN(n9804) );
  NAND2_X1 U11741 ( .A1(n15420), .A2(n9787), .ZN(n9786) );
  INV_X1 U11742 ( .A(n9789), .ZN(n9788) );
  NOR2_X1 U11743 ( .A1(n10097), .A2(n14195), .ZN(n9787) );
  AND2_X1 U11744 ( .A1(n11836), .A2(n10039), .ZN(n15413) );
  AOI21_X1 U11745 ( .B1(n15527), .B2(n15528), .A(n15465), .ZN(n15516) );
  INV_X1 U11746 ( .A(n15466), .ZN(n9913) );
  AND2_X1 U11747 ( .A1(n9860), .A2(n9868), .ZN(n15460) );
  AND2_X1 U11748 ( .A1(n13256), .A2(n9967), .ZN(n13583) );
  AND3_X1 U11749 ( .A1(n12327), .A2(n12326), .A3(n12325), .ZN(n13565) );
  NAND2_X2 U11750 ( .A1(n9657), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14303) );
  NAND2_X1 U11751 ( .A1(n12970), .A2(n19645), .ZN(n13126) );
  INV_X1 U11752 ( .A(n13114), .ZN(n13132) );
  XNOR2_X1 U11753 ( .A(n15826), .B(n13119), .ZN(n13123) );
  OR2_X1 U11754 ( .A1(n13134), .A2(n13133), .ZN(n13201) );
  INV_X1 U11755 ( .A(n10135), .ZN(n10134) );
  AND2_X2 U11756 ( .A1(n11504), .A2(n11502), .ZN(n11557) );
  INV_X1 U11757 ( .A(n19781), .ZN(n19466) );
  NOR2_X1 U11758 ( .A1(n19934), .A2(n19297), .ZN(n19714) );
  OR2_X1 U11759 ( .A1(n11213), .A2(n11984), .ZN(n16357) );
  AOI21_X1 U11760 ( .B1(n16693), .B2(n16863), .A(n16862), .ZN(n16684) );
  OAI21_X1 U11761 ( .B1(n16593), .B2(n9893), .A(n9894), .ZN(n9891) );
  OR2_X1 U11762 ( .A1(n12021), .A2(n12019), .ZN(n9699) );
  INV_X1 U11763 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15873) );
  AOI21_X1 U11764 ( .B1(n15896), .B2(n18752), .A(n14065), .ZN(n15988) );
  NOR2_X1 U11765 ( .A1(n17241), .A2(n18597), .ZN(n12652) );
  NOR2_X1 U11766 ( .A1(n17558), .A2(n17557), .ZN(n17556) );
  NAND2_X1 U11767 ( .A1(n17638), .A2(n10168), .ZN(n17623) );
  INV_X1 U11768 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n9884) );
  INV_X1 U11769 ( .A(n16801), .ZN(n9885) );
  NOR2_X1 U11770 ( .A1(n17766), .A2(n17755), .ZN(n17749) );
  INV_X1 U11771 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17766) );
  AOI21_X1 U11772 ( .B1(n12695), .B2(n9691), .A(n10022), .ZN(n12701) );
  NOR2_X1 U11773 ( .A1(n17600), .A2(n17924), .ZN(n17920) );
  NAND2_X1 U11774 ( .A1(n17709), .A2(n12685), .ZN(n12687) );
  NAND2_X1 U11775 ( .A1(n17656), .A2(n12689), .ZN(n17627) );
  INV_X1 U11776 ( .A(n12113), .ZN(n15906) );
  OAI211_X1 U11777 ( .C1(n17163), .C2(n17113), .A(n12573), .B(n12572), .ZN(
        n16437) );
  NAND2_X1 U11778 ( .A1(n15917), .A2(n15891), .ZN(n18757) );
  AOI22_X1 U11779 ( .A1(n12616), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12043) );
  NAND2_X1 U11780 ( .A1(n11094), .A2(n20000), .ZN(n14769) );
  NAND2_X1 U11781 ( .A1(n11093), .A2(n11092), .ZN(n11094) );
  INV_X1 U11782 ( .A(n14769), .ZN(n14778) );
  INV_X2 U11783 ( .A(n16049), .ZN(n20239) );
  XNOR2_X1 U11784 ( .A(n9833), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15025) );
  OR2_X1 U11785 ( .A1(n10160), .A2(n15195), .ZN(n10003) );
  XNOR2_X1 U11786 ( .A(n12809), .B(n11960), .ZN(n16186) );
  NAND2_X1 U11787 ( .A1(n12810), .A2(n12809), .ZN(n14457) );
  NAND2_X1 U11788 ( .A1(n12808), .A2(n12552), .ZN(n16199) );
  XNOR2_X1 U11789 ( .A(n14170), .B(n14169), .ZN(n19148) );
  NAND2_X1 U11790 ( .A1(n9870), .A2(n9869), .ZN(n11796) );
  OR2_X1 U11791 ( .A1(n12806), .A2(n14170), .ZN(n14451) );
  INV_X1 U11792 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19966) );
  NAND2_X1 U11793 ( .A1(n12976), .A2(n12975), .ZN(n19961) );
  INV_X1 U11794 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19956) );
  AND2_X1 U11795 ( .A1(n19942), .A2(n19949), .ZN(n19941) );
  INV_X1 U11796 ( .A(n19494), .ZN(n19931) );
  INV_X1 U11797 ( .A(n16937), .ZN(n16929) );
  NAND2_X1 U11798 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17376), .ZN(n17372) );
  NAND2_X1 U11799 ( .A1(n20572), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11010) );
  INV_X1 U11800 ( .A(n10442), .ZN(n10111) );
  AND2_X1 U11801 ( .A1(n13182), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10192) );
  OR2_X1 U11802 ( .A1(n11021), .A2(n11026), .ZN(n11023) );
  NAND2_X1 U11803 ( .A1(n11023), .A2(n11010), .ZN(n11020) );
  AOI22_X1 U11804 ( .A1(n11020), .A2(n11011), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20646), .ZN(n11015) );
  OR2_X1 U11805 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20646), .ZN(
        n11011) );
  INV_X1 U11806 ( .A(n10114), .ZN(n10113) );
  NOR2_X1 U11807 ( .A1(n10355), .A2(n10354), .ZN(n12173) );
  OR2_X1 U11808 ( .A1(n11042), .A2(n10509), .ZN(n10521) );
  OR2_X1 U11809 ( .A1(n10496), .A2(n10495), .ZN(n12188) );
  NAND2_X1 U11810 ( .A1(n10423), .A2(n10422), .ZN(n10424) );
  NAND2_X1 U11811 ( .A1(n13417), .A2(n9773), .ZN(n13167) );
  AND2_X1 U11812 ( .A1(n13166), .A2(n9774), .ZN(n9773) );
  NAND2_X1 U11813 ( .A1(n13632), .A2(n12247), .ZN(n9774) );
  INV_X1 U11814 ( .A(n10097), .ZN(n9952) );
  INV_X1 U11815 ( .A(n16268), .ZN(n11703) );
  OR2_X1 U11816 ( .A1(n11585), .A2(n11584), .ZN(n11656) );
  NAND2_X1 U11817 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10075) );
  NAND2_X1 U11818 ( .A1(n11557), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10077) );
  OR2_X1 U11819 ( .A1(n11463), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11464) );
  NOR2_X1 U11820 ( .A1(n11389), .A2(n12969), .ZN(n9805) );
  INV_X1 U11821 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10140) );
  XNOR2_X1 U11822 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11206) );
  AND2_X1 U11823 ( .A1(n11205), .A2(n11197), .ZN(n11208) );
  NOR2_X1 U11824 ( .A1(n15905), .A2(n17292), .ZN(n12116) );
  INV_X1 U11825 ( .A(n12670), .ZN(n10027) );
  INV_X1 U11826 ( .A(n12834), .ZN(n10124) );
  NAND2_X1 U11827 ( .A1(n14004), .A2(n9813), .ZN(n14673) );
  NOR2_X1 U11828 ( .A1(n10112), .A2(n9814), .ZN(n9813) );
  INV_X1 U11829 ( .A(n14003), .ZN(n9814) );
  NAND2_X1 U11830 ( .A1(n10113), .A2(n10709), .ZN(n10112) );
  NAND2_X1 U11831 ( .A1(n14771), .A2(n10118), .ZN(n10117) );
  NAND2_X1 U11832 ( .A1(n10581), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10607) );
  INV_X1 U11833 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10606) );
  NOR2_X1 U11834 ( .A1(n9937), .A2(n14560), .ZN(n9936) );
  INV_X1 U11835 ( .A(n9938), .ZN(n9937) );
  NOR2_X1 U11836 ( .A1(n14575), .A2(n9939), .ZN(n9938) );
  INV_X1 U11837 ( .A(n14587), .ZN(n9939) );
  NOR2_X1 U11838 ( .A1(n9931), .A2(n14629), .ZN(n9930) );
  INV_X1 U11839 ( .A(n9932), .ZN(n9931) );
  NOR2_X1 U11840 ( .A1(n9934), .A2(n9933), .ZN(n9932) );
  INV_X1 U11841 ( .A(n14650), .ZN(n9934) );
  INV_X1 U11842 ( .A(n14640), .ZN(n9933) );
  INV_X1 U11843 ( .A(n9776), .ZN(n9775) );
  NOR2_X1 U11844 ( .A1(n13632), .A2(n20267), .ZN(n11180) );
  NOR2_X1 U11845 ( .A1(n13747), .A2(n13826), .ZN(n9924) );
  INV_X1 U11846 ( .A(n11180), .ZN(n11162) );
  NAND2_X1 U11847 ( .A1(n13329), .A2(n12219), .ZN(n12215) );
  XNOR2_X1 U11848 ( .A(n10421), .B(n10419), .ZN(n10434) );
  NAND2_X1 U11849 ( .A1(n10101), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10100) );
  NAND2_X1 U11850 ( .A1(n13423), .A2(n20914), .ZN(n10472) );
  NAND2_X1 U11851 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n9822) );
  NAND2_X1 U11852 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n9823) );
  NAND2_X1 U11853 ( .A1(n10343), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n9826) );
  NAND2_X1 U11854 ( .A1(n10415), .A2(n10414), .ZN(n20297) );
  INV_X1 U11855 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20572) );
  AND2_X1 U11856 ( .A1(n11046), .A2(n12214), .ZN(n11045) );
  AOI221_X1 U11857 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n11013), 
        .C1(n16175), .C2(n11013), .A(n11012), .ZN(n11061) );
  INV_X1 U11858 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20646) );
  NAND2_X1 U11859 ( .A1(n11741), .A2(n11740), .ZN(n11743) );
  NAND2_X1 U11860 ( .A1(n9742), .A2(n10172), .ZN(n9949) );
  AND2_X1 U11861 ( .A1(n9951), .A2(n11705), .ZN(n9950) );
  AND2_X1 U11862 ( .A1(n13360), .A2(n13519), .ZN(n9951) );
  AND4_X1 U11863 ( .A1(n11634), .A2(n11633), .A3(n11632), .A4(n11631), .ZN(
        n11645) );
  AND4_X1 U11864 ( .A1(n11642), .A2(n11641), .A3(n11640), .A4(n11639), .ZN(
        n11643) );
  NOR4_X2 U11865 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n15832), .A4(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14245) );
  NAND2_X1 U11866 ( .A1(n10136), .A2(n10138), .ZN(n14356) );
  NAND2_X1 U11867 ( .A1(n9690), .A2(n15262), .ZN(n10138) );
  NAND2_X1 U11868 ( .A1(n13819), .A2(n9689), .ZN(n10145) );
  NAND2_X1 U11869 ( .A1(n10001), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10000) );
  INV_X1 U11870 ( .A(n11845), .ZN(n10001) );
  NAND2_X1 U11871 ( .A1(n11842), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10008) );
  NAND2_X1 U11872 ( .A1(n11618), .A2(n11617), .ZN(n11816) );
  INV_X1 U11873 ( .A(n11547), .ZN(n12311) );
  OR2_X1 U11874 ( .A1(n11249), .A2(n11248), .ZN(n12292) );
  OR2_X1 U11875 ( .A1(n19969), .A2(n12288), .ZN(n11306) );
  OR2_X1 U11876 ( .A1(n11786), .A2(n11785), .ZN(n11791) );
  INV_X1 U11877 ( .A(n14185), .ZN(n9872) );
  NOR2_X1 U11878 ( .A1(n10097), .A2(n9718), .ZN(n10096) );
  OAI21_X1 U11879 ( .B1(n15420), .B2(n9791), .A(n9790), .ZN(n9789) );
  INV_X1 U11880 ( .A(n9792), .ZN(n9791) );
  AOI22_X1 U11881 ( .A1(n10097), .A2(n9792), .B1(n9796), .B2(n9795), .ZN(n9790) );
  NOR2_X1 U11882 ( .A1(n9795), .A2(n9796), .ZN(n9792) );
  NOR2_X1 U11883 ( .A1(n15607), .A2(n15414), .ZN(n10039) );
  NAND2_X1 U11884 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10038) );
  AND2_X1 U11885 ( .A1(n11931), .A2(n11930), .ZN(n12898) );
  INV_X1 U11886 ( .A(n15299), .ZN(n10066) );
  AND2_X1 U11887 ( .A1(n9980), .A2(n9979), .ZN(n9978) );
  INV_X1 U11888 ( .A(n15664), .ZN(n9979) );
  AND2_X1 U11889 ( .A1(n15219), .A2(n13991), .ZN(n9980) );
  OR2_X1 U11890 ( .A1(n19006), .A2(n15461), .ZN(n11747) );
  NOR2_X1 U11891 ( .A1(n11748), .A2(n15508), .ZN(n15466) );
  INV_X1 U11892 ( .A(n15741), .ZN(n9903) );
  NAND2_X1 U11893 ( .A1(n9702), .A2(n15551), .ZN(n10093) );
  NAND2_X1 U11894 ( .A1(n10050), .A2(n13515), .ZN(n10049) );
  INV_X1 U11895 ( .A(n13356), .ZN(n10050) );
  INV_X1 U11896 ( .A(n11824), .ZN(n11825) );
  NAND2_X1 U11897 ( .A1(n11818), .A2(n9720), .ZN(n9850) );
  NAND2_X1 U11898 ( .A1(n11682), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9918) );
  AND2_X1 U11899 ( .A1(n13211), .A2(n11854), .ZN(n10054) );
  INV_X1 U11900 ( .A(n13488), .ZN(n10034) );
  NAND2_X1 U11901 ( .A1(n11666), .A2(n11665), .ZN(n11809) );
  AND2_X1 U11902 ( .A1(n13074), .A2(n13073), .ZN(n13076) );
  NAND2_X1 U11903 ( .A1(n11454), .A2(n10146), .ZN(n11460) );
  OR2_X1 U11904 ( .A1(n12513), .A2(n12512), .ZN(n15836) );
  OAI21_X1 U11905 ( .B1(n13115), .B2(n13114), .A(n13113), .ZN(n13117) );
  AND2_X1 U11906 ( .A1(n11502), .A2(n13115), .ZN(n11497) );
  NAND2_X1 U11907 ( .A1(n18273), .A2(n12116), .ZN(n12112) );
  INV_X1 U11908 ( .A(n12711), .ZN(n12720) );
  NOR2_X1 U11909 ( .A1(n17623), .A2(n17622), .ZN(n17594) );
  NAND2_X1 U11910 ( .A1(n15906), .A2(n9843), .ZN(n12122) );
  NOR2_X1 U11911 ( .A1(n12120), .A2(n9844), .ZN(n9843) );
  NAND2_X1 U11912 ( .A1(n18277), .A2(n18281), .ZN(n9844) );
  NAND2_X1 U11913 ( .A1(n17626), .A2(n17655), .ZN(n17656) );
  NAND2_X1 U11914 ( .A1(n12757), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17708) );
  NOR2_X1 U11915 ( .A1(n12747), .A2(n17850), .ZN(n12750) );
  NOR2_X1 U11916 ( .A1(n12743), .A2(n17857), .ZN(n12745) );
  AND2_X1 U11917 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12742), .ZN(
        n12743) );
  NAND2_X1 U11918 ( .A1(n18277), .A2(n18273), .ZN(n18714) );
  AOI21_X1 U11919 ( .B1(n12713), .B2(n15987), .A(n12712), .ZN(n18713) );
  AOI211_X1 U11920 ( .C1(n17228), .C2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n12028), .B(n12027), .ZN(n12029) );
  NOR2_X1 U11921 ( .A1(n18909), .A2(n18788), .ZN(n18265) );
  NAND2_X1 U11922 ( .A1(n15888), .A2(n15907), .ZN(n17446) );
  NAND2_X1 U11923 ( .A1(n9771), .A2(n13632), .ZN(n10280) );
  INV_X1 U11924 ( .A(n12247), .ZN(n9771) );
  INV_X1 U11925 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20037) );
  INV_X1 U11926 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20066) );
  AND2_X1 U11927 ( .A1(n14665), .A2(n14650), .ZN(n14652) );
  AND2_X1 U11928 ( .A1(n11106), .A2(n11105), .ZN(n13470) );
  NAND2_X1 U11929 ( .A1(n13082), .A2(n9658), .ZN(n9926) );
  AND2_X1 U11930 ( .A1(n10744), .A2(n10743), .ZN(n14662) );
  AOI21_X1 U11931 ( .B1(n12179), .B2(n10684), .A(n10506), .ZN(n13377) );
  INV_X1 U11932 ( .A(n20127), .ZN(n13229) );
  NAND2_X1 U11933 ( .A1(n10932), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10976) );
  OR2_X1 U11934 ( .A1(n10909), .A2(n10908), .ZN(n10910) );
  OR2_X1 U11935 ( .A1(n10913), .A2(n10912), .ZN(n14557) );
  INV_X1 U11936 ( .A(n10876), .ZN(n10877) );
  OR2_X1 U11937 ( .A1(n10890), .A2(n10889), .ZN(n14585) );
  AOI21_X1 U11938 ( .B1(n10848), .B2(n10847), .A(n10846), .ZN(n14596) );
  AND2_X1 U11939 ( .A1(n14597), .A2(n13628), .ZN(n10846) );
  AND2_X1 U11940 ( .A1(n10813), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10814) );
  INV_X1 U11941 ( .A(n10812), .ZN(n10813) );
  AND2_X1 U11942 ( .A1(n10819), .A2(n10818), .ZN(n14608) );
  OR2_X1 U11943 ( .A1(n14926), .A2(n11004), .ZN(n10818) );
  NAND2_X1 U11944 ( .A1(n10776), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10812) );
  AND2_X1 U11945 ( .A1(n10759), .A2(n10758), .ZN(n14649) );
  INV_X1 U11946 ( .A(n10720), .ZN(n10738) );
  AOI21_X1 U11947 ( .B1(n10970), .B2(n10723), .A(n10722), .ZN(n14674) );
  NOR2_X1 U11948 ( .A1(n10705), .A2(n14696), .ZN(n10706) );
  NAND2_X1 U11949 ( .A1(n10675), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10705) );
  NOR2_X1 U11950 ( .A1(n10660), .A2(n10659), .ZN(n10675) );
  NAND2_X1 U11951 ( .A1(n10645), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10660) );
  INV_X1 U11952 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10659) );
  AND2_X1 U11953 ( .A1(n10612), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10613) );
  AOI21_X1 U11954 ( .B1(n20028), .B2(n13628), .A(n10595), .ZN(n13742) );
  CLKBUF_X1 U11955 ( .A(n13690), .Z(n13691) );
  NOR2_X1 U11956 ( .A1(n10560), .A2(n20037), .ZN(n10581) );
  AOI21_X1 U11957 ( .B1(n12205), .B2(n10684), .A(n10565), .ZN(n13653) );
  NAND2_X1 U11958 ( .A1(n10549), .A2(n10548), .ZN(n13531) );
  NOR2_X1 U11959 ( .A1(n10522), .A2(n20066), .ZN(n10544) );
  NAND2_X1 U11960 ( .A1(n10502), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10522) );
  NAND2_X1 U11961 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10478) );
  NOR2_X1 U11962 ( .A1(n10478), .A2(n10477), .ZN(n10502) );
  INV_X1 U11963 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10477) );
  INV_X1 U11964 ( .A(n13296), .ZN(n10451) );
  NAND2_X1 U11965 ( .A1(n13254), .A2(n13253), .ZN(n13296) );
  INV_X1 U11966 ( .A(n9830), .ZN(n9829) );
  NAND2_X1 U11967 ( .A1(n14858), .A2(n12224), .ZN(n9831) );
  NAND2_X1 U11968 ( .A1(n14601), .A2(n9936), .ZN(n14558) );
  NAND2_X1 U11969 ( .A1(n14601), .A2(n14587), .ZN(n14586) );
  NAND2_X1 U11970 ( .A1(n14601), .A2(n9938), .ZN(n14573) );
  AND2_X1 U11971 ( .A1(n14614), .A2(n14599), .ZN(n14601) );
  AND2_X1 U11972 ( .A1(n14665), .A2(n9928), .ZN(n14614) );
  NOR2_X1 U11973 ( .A1(n9929), .A2(n14612), .ZN(n9928) );
  INV_X1 U11974 ( .A(n9930), .ZN(n9929) );
  NAND2_X1 U11975 ( .A1(n10043), .A2(n14972), .ZN(n14922) );
  NAND2_X1 U11976 ( .A1(n14665), .A2(n9930), .ZN(n14627) );
  NAND2_X1 U11977 ( .A1(n14665), .A2(n9932), .ZN(n14639) );
  NOR2_X1 U11978 ( .A1(n14678), .A2(n14663), .ZN(n14665) );
  OR2_X1 U11979 ( .A1(n14676), .A2(n14675), .ZN(n14678) );
  NAND2_X1 U11980 ( .A1(n14691), .A2(n14030), .ZN(n14676) );
  NAND2_X1 U11981 ( .A1(n14007), .A2(n14006), .ZN(n14708) );
  NOR2_X2 U11982 ( .A1(n13746), .A2(n9923), .ZN(n14007) );
  NAND2_X1 U11983 ( .A1(n9924), .A2(n14000), .ZN(n9923) );
  INV_X1 U11984 ( .A(n9837), .ZN(n9836) );
  OAI21_X1 U11985 ( .B1(n9838), .B2(n9700), .A(n12225), .ZN(n9837) );
  NAND2_X1 U11986 ( .A1(n9925), .A2(n11124), .ZN(n13827) );
  INV_X1 U11987 ( .A(n20212), .ZN(n16142) );
  OR2_X1 U11988 ( .A1(n13469), .A2(n13380), .ZN(n13382) );
  AND2_X1 U11989 ( .A1(n15100), .A2(n15098), .ZN(n20212) );
  INV_X1 U11990 ( .A(n20209), .ZN(n20210) );
  NAND2_X1 U11991 ( .A1(n11162), .A2(n11155), .ZN(n14491) );
  CLKBUF_X1 U11992 ( .A(n13415), .Z(n13416) );
  INV_X1 U11993 ( .A(n20431), .ZN(n20490) );
  INV_X1 U11994 ( .A(n20698), .ZN(n20551) );
  INV_X1 U11995 ( .A(n20275), .ZN(n20290) );
  INV_X1 U11996 ( .A(n20778), .ZN(n20720) );
  AOI21_X1 U11997 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20692), .A(n20299), 
        .ZN(n20779) );
  INV_X1 U11998 ( .A(n13440), .ZN(n15949) );
  NAND2_X1 U11999 ( .A1(n11770), .A2(n11771), .ZN(n11775) );
  INV_X1 U12000 ( .A(n9984), .ZN(n9983) );
  AOI21_X1 U12001 ( .B1(n12794), .B2(n15425), .A(n16210), .ZN(n9984) );
  AND2_X1 U12002 ( .A1(n11695), .A2(n13360), .ZN(n11697) );
  AND2_X1 U12003 ( .A1(n11695), .A2(n9951), .ZN(n11706) );
  CLKBUF_X1 U12004 ( .A(n11684), .Z(n11691) );
  OR2_X1 U12005 ( .A1(n9946), .A2(n9945), .ZN(n11663) );
  AND2_X1 U12006 ( .A1(n11920), .A2(n11919), .ZN(n15306) );
  NOR2_X1 U12007 ( .A1(n9694), .A2(n15306), .ZN(n15307) );
  NAND2_X1 U12008 ( .A1(n10132), .A2(n10131), .ZN(n10130) );
  NAND2_X1 U12009 ( .A1(n14379), .A2(n10132), .ZN(n10129) );
  AND2_X1 U12010 ( .A1(n12480), .A2(n12479), .ZN(n13898) );
  AND2_X1 U12011 ( .A1(n14393), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13209) );
  AND2_X1 U12012 ( .A1(n13025), .A2(n19988), .ZN(n19197) );
  INV_X1 U12013 ( .A(n13003), .ZN(n13853) );
  INV_X1 U12014 ( .A(n12807), .ZN(n10056) );
  NAND2_X1 U12015 ( .A1(n12884), .A2(n10057), .ZN(n12808) );
  NAND2_X1 U12016 ( .A1(n12884), .A2(n14197), .ZN(n12550) );
  AND2_X1 U12017 ( .A1(n11947), .A2(n11946), .ZN(n12885) );
  NOR2_X1 U12018 ( .A1(n10059), .A2(n15251), .ZN(n10058) );
  INV_X1 U12019 ( .A(n10060), .ZN(n10059) );
  NAND2_X1 U12020 ( .A1(n9997), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9996) );
  INV_X1 U12021 ( .A(n9998), .ZN(n9997) );
  AND2_X1 U12022 ( .A1(n11917), .A2(n11916), .ZN(n13923) );
  AND2_X1 U12023 ( .A1(n11908), .A2(n11907), .ZN(n12860) );
  AND2_X1 U12024 ( .A1(n11905), .A2(n11904), .ZN(n13712) );
  INV_X1 U12025 ( .A(n10068), .ZN(n13714) );
  AND2_X1 U12026 ( .A1(n11891), .A2(n11890), .ZN(n13622) );
  AND2_X1 U12027 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11840) );
  AND2_X1 U12028 ( .A1(n11867), .A2(n11866), .ZN(n13203) );
  NAND2_X1 U12029 ( .A1(n9873), .A2(n9875), .ZN(n14182) );
  INV_X1 U12030 ( .A(n9974), .ZN(n9972) );
  NAND2_X1 U12031 ( .A1(n15334), .A2(n12882), .ZN(n15190) );
  NOR2_X1 U12032 ( .A1(n15356), .A2(n15203), .ZN(n15337) );
  NOR2_X1 U12033 ( .A1(n10038), .A2(n15619), .ZN(n10036) );
  OR2_X1 U12034 ( .A1(n15354), .A2(n15353), .ZN(n15356) );
  OR2_X1 U12035 ( .A1(n12869), .A2(n15461), .ZN(n11762) );
  NAND2_X1 U12036 ( .A1(n15220), .A2(n9976), .ZN(n12896) );
  AND2_X1 U12037 ( .A1(n9978), .A2(n9977), .ZN(n9976) );
  INV_X1 U12038 ( .A(n15378), .ZN(n9977) );
  NOR2_X1 U12039 ( .A1(n12896), .A2(n12897), .ZN(n12895) );
  NAND2_X1 U12040 ( .A1(n9863), .A2(n9861), .ZN(n9867) );
  NAND2_X1 U12041 ( .A1(n15459), .A2(n11704), .ZN(n9807) );
  NOR3_X1 U12042 ( .A1(n9694), .A2(n10066), .A3(n15306), .ZN(n15301) );
  NAND2_X1 U12043 ( .A1(n15220), .A2(n9978), .ZN(n15667) );
  NAND2_X1 U12044 ( .A1(n15220), .A2(n9980), .ZN(n15665) );
  NOR2_X1 U12045 ( .A1(n15505), .A2(n15466), .ZN(n9914) );
  NAND2_X1 U12046 ( .A1(n15782), .A2(n9741), .ZN(n13897) );
  INV_X1 U12047 ( .A(n13861), .ZN(n9963) );
  NAND2_X1 U12048 ( .A1(n10068), .A2(n10067), .ZN(n13849) );
  INV_X1 U12049 ( .A(n12860), .ZN(n10067) );
  AND2_X1 U12050 ( .A1(n11911), .A2(n11910), .ZN(n13848) );
  OR3_X1 U12051 ( .A1(n11749), .A2(n15461), .A3(n15543), .ZN(n15539) );
  OR2_X1 U12052 ( .A1(n9905), .A2(n9903), .ZN(n9901) );
  AOI21_X1 U12053 ( .B1(n9906), .B2(n11739), .A(n15463), .ZN(n9905) );
  OR2_X1 U12054 ( .A1(n9907), .A2(n9903), .ZN(n9902) );
  AND3_X1 U12055 ( .A1(n12458), .A2(n12457), .A3(n12456), .ZN(n15747) );
  NOR2_X1 U12056 ( .A1(n15783), .A2(n15784), .ZN(n15782) );
  NAND2_X1 U12057 ( .A1(n15782), .A2(n13506), .ZN(n15748) );
  INV_X1 U12058 ( .A(n10093), .ZN(n10091) );
  NOR2_X1 U12059 ( .A1(n13573), .A2(n13572), .ZN(n13571) );
  NAND2_X1 U12060 ( .A1(n13256), .A2(n9966), .ZN(n13573) );
  AND2_X1 U12061 ( .A1(n9967), .A2(n13276), .ZN(n9966) );
  OR2_X1 U12062 ( .A1(n11700), .A2(n15810), .ZN(n16268) );
  NAND2_X1 U12063 ( .A1(n9710), .A2(n11693), .ZN(n10094) );
  AND2_X1 U12064 ( .A1(n13607), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16278) );
  OAI21_X1 U12065 ( .B1(n13484), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n13485), .ZN(n11676) );
  NAND2_X1 U12066 ( .A1(n10055), .A2(n10054), .ZN(n13212) );
  XNOR2_X1 U12067 ( .A(n13076), .B(n12306), .ZN(n13050) );
  AOI21_X1 U12068 ( .B1(n11496), .B2(n13132), .A(n13043), .ZN(n13122) );
  CLKBUF_X1 U12069 ( .A(n13762), .Z(n15848) );
  NOR2_X2 U12070 ( .A1(n12263), .A2(n11985), .ZN(n16363) );
  NAND2_X1 U12071 ( .A1(n11335), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11342) );
  NOR2_X2 U12072 ( .A1(n13854), .A2(n13736), .ZN(n19292) );
  INV_X1 U12073 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19769) );
  NOR2_X1 U12074 ( .A1(n18273), .A2(n12122), .ZN(n15889) );
  NAND2_X1 U12075 ( .A1(n9841), .A2(n9739), .ZN(n18764) );
  NAND2_X1 U12076 ( .A1(n18750), .A2(n18752), .ZN(n9841) );
  AND2_X1 U12077 ( .A1(n16597), .A2(n12005), .ZN(n16586) );
  AND2_X1 U12078 ( .A1(n16628), .A2(n12005), .ZN(n16619) );
  OR2_X1 U12079 ( .A1(n16630), .A2(n17597), .ZN(n16628) );
  AND2_X1 U12080 ( .A1(n16649), .A2(n12005), .ZN(n16641) );
  NOR2_X1 U12081 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16744), .ZN(n16733) );
  NAND2_X1 U12082 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17158), .ZN(n15874) );
  AND3_X1 U12083 ( .A1(n12045), .A2(n9729), .A3(n12046), .ZN(n12048) );
  INV_X1 U12084 ( .A(n17285), .ZN(n14067) );
  OR3_X2 U12085 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18728), .ZN(n12608) );
  NAND2_X1 U12086 ( .A1(n12616), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10010) );
  INV_X1 U12087 ( .A(n12615), .ZN(n12620) );
  NOR2_X1 U12088 ( .A1(n17483), .A2(n17446), .ZN(n17464) );
  NOR2_X1 U12089 ( .A1(n18781), .A2(n16553), .ZN(n17484) );
  NOR2_X1 U12090 ( .A1(n11995), .A2(n16593), .ZN(n12001) );
  NAND2_X1 U12091 ( .A1(n11996), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12011) );
  INV_X1 U12092 ( .A(n17594), .ZN(n17605) );
  INV_X1 U12093 ( .A(n11999), .ZN(n12009) );
  AND2_X1 U12094 ( .A1(n17711), .A2(n9886), .ZN(n17638) );
  AND2_X1 U12095 ( .A1(n9683), .A2(n9745), .ZN(n9886) );
  NAND2_X1 U12096 ( .A1(n17711), .A2(n10170), .ZN(n17698) );
  AOI21_X1 U12097 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17664), .A(
        n18304), .ZN(n17722) );
  NOR2_X1 U12098 ( .A1(n17819), .A2(n9701), .ZN(n9883) );
  NOR2_X1 U12099 ( .A1(n17819), .A2(n16801), .ZN(n17788) );
  NAND2_X1 U12100 ( .A1(n17415), .A2(n9659), .ZN(n17758) );
  NOR2_X1 U12101 ( .A1(n17873), .A2(n11994), .ZN(n17853) );
  NAND2_X1 U12102 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11994) );
  NOR2_X1 U12103 ( .A1(n12741), .A2(n17870), .ZN(n17859) );
  NOR2_X1 U12104 ( .A1(n17859), .A2(n17858), .ZN(n17857) );
  NOR2_X1 U12105 ( .A1(n12701), .A2(n12697), .ZN(n15974) );
  NAND2_X1 U12106 ( .A1(n15974), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15973) );
  AOI21_X1 U12107 ( .B1(n12690), .B2(n10022), .A(n12691), .ZN(n10021) );
  NOR2_X1 U12108 ( .A1(n17782), .A2(n18035), .ZN(n17974) );
  NOR2_X1 U12109 ( .A1(n17720), .A2(n17618), .ZN(n17955) );
  NOR2_X1 U12110 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n12686), .ZN(
        n17657) );
  NAND2_X1 U12111 ( .A1(n12683), .A2(n12681), .ZN(n12682) );
  NAND2_X1 U12112 ( .A1(n10022), .A2(n18053), .ZN(n12681) );
  NAND2_X1 U12113 ( .A1(n17704), .A2(n18029), .ZN(n17703) );
  INV_X1 U12114 ( .A(n18121), .ZN(n17782) );
  NOR2_X1 U12115 ( .A1(n10022), .A2(n17771), .ZN(n17761) );
  INV_X1 U12116 ( .A(n18750), .ZN(n18097) );
  NAND2_X1 U12117 ( .A1(n17840), .A2(n10016), .ZN(n17794) );
  INV_X1 U12118 ( .A(n10150), .ZN(n10017) );
  NOR2_X1 U12119 ( .A1(n17783), .A2(n10018), .ZN(n18121) );
  NOR2_X1 U12120 ( .A1(n12755), .A2(n17825), .ZN(n18123) );
  NOR2_X1 U12121 ( .A1(n17852), .A2(n17851), .ZN(n17850) );
  OR2_X1 U12122 ( .A1(n17885), .A2(n18216), .ZN(n10015) );
  INV_X1 U12123 ( .A(n12120), .ZN(n12124) );
  NOR2_X1 U12124 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18265), .ZN(n18568) );
  OAI211_X1 U12125 ( .C1(n14519), .C2(n11192), .A(n14518), .B(n9704), .ZN(
        n14520) );
  AND2_X1 U12126 ( .A1(n14620), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n14605) );
  OR2_X1 U12127 ( .A1(n14644), .A2(n14503), .ZN(n14604) );
  AND2_X1 U12128 ( .A1(n13641), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13631) );
  NAND2_X1 U12129 ( .A1(n13640), .A2(n13635), .ZN(n20044) );
  AND2_X1 U12130 ( .A1(n14727), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20091) );
  NAND2_X1 U12131 ( .A1(n14727), .A2(n13642), .ZN(n20078) );
  XNOR2_X1 U12132 ( .A(n9927), .B(n13082), .ZN(n13648) );
  OR2_X1 U12133 ( .A1(n14488), .A2(n14167), .ZN(n14527) );
  INV_X1 U12134 ( .A(n14820), .ZN(n14840) );
  INV_X1 U12135 ( .A(n14823), .ZN(n14842) );
  OR2_X1 U12136 ( .A1(n13193), .A2(n11068), .ZN(n11069) );
  INV_X1 U12137 ( .A(n10629), .ZN(n9815) );
  INV_X2 U12138 ( .A(n14849), .ZN(n14853) );
  CLKBUF_X1 U12139 ( .A(n20125), .Z(n20919) );
  INV_X2 U12140 ( .A(n13386), .ZN(n20164) );
  INV_X1 U12141 ( .A(n20007), .ZN(n20174) );
  NOR2_X1 U12142 ( .A1(n14856), .A2(n9778), .ZN(n9777) );
  INV_X1 U12143 ( .A(n9835), .ZN(n13868) );
  AOI21_X1 U12144 ( .B1(n9840), .B2(n9838), .A(n9700), .ZN(n9835) );
  NAND2_X1 U12145 ( .A1(n9840), .A2(n12213), .ZN(n13799) );
  INV_X1 U12147 ( .A(n20222), .ZN(n20206) );
  AND2_X1 U12148 ( .A1(n13340), .A2(n14474), .ZN(n20209) );
  NAND2_X1 U12149 ( .A1(n20212), .A2(n20210), .ZN(n20220) );
  INV_X1 U12150 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20692) );
  NAND2_X1 U12151 ( .A1(n10046), .A2(n10442), .ZN(n10045) );
  NAND2_X1 U12152 ( .A1(n10441), .A2(n10443), .ZN(n10046) );
  CLKBUF_X1 U12153 ( .A(n12248), .Z(n20783) );
  OAI21_X1 U12154 ( .B1(n13445), .B2(n16182), .A(n20299), .ZN(n20235) );
  NOR2_X1 U12155 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16172) );
  OAI211_X1 U12156 ( .C1(n20291), .C2(n20525), .A(n20577), .B(n20250), .ZN(
        n20294) );
  NAND2_X1 U12157 ( .A1(n20369), .A2(n20719), .ZN(n20394) );
  INV_X1 U12158 ( .A(n20448), .ZN(n20451) );
  OAI211_X1 U12159 ( .C1(n20541), .C2(n20525), .A(n20577), .B(n20524), .ZN(
        n20543) );
  OAI22_X1 U12160 ( .A1(n20581), .A2(n20580), .B1(n20579), .B2(n20724), .ZN(
        n20605) );
  INV_X1 U12161 ( .A(n20647), .ZN(n20774) );
  INV_X1 U12162 ( .A(n20660), .ZN(n20789) );
  INV_X1 U12163 ( .A(n20664), .ZN(n20795) );
  INV_X1 U12164 ( .A(n20668), .ZN(n20801) );
  INV_X1 U12165 ( .A(n20672), .ZN(n20807) );
  INV_X1 U12166 ( .A(n20680), .ZN(n20819) );
  NOR2_X2 U12167 ( .A1(n20778), .A2(n20242), .ZN(n20829) );
  INV_X1 U12168 ( .A(n20685), .ZN(n20827) );
  NOR2_X1 U12169 ( .A1(n20525), .A2(n14483), .ZN(n15968) );
  NAND2_X1 U12171 ( .A1(n16181), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20835) );
  NOR2_X1 U12172 ( .A1(n16357), .A2(n12823), .ZN(n12905) );
  CLKBUF_X1 U12173 ( .A(n12515), .Z(n12913) );
  INV_X1 U12174 ( .A(n10005), .ZN(n16194) );
  NAND2_X1 U12175 ( .A1(n10005), .A2(n10004), .ZN(n16193) );
  INV_X1 U12176 ( .A(n9985), .ZN(n15206) );
  OAI21_X1 U12177 ( .B1(n18980), .B2(n9992), .A(n9991), .ZN(n12890) );
  NAND2_X1 U12178 ( .A1(n15456), .A2(n9993), .ZN(n9992) );
  NAND2_X1 U12179 ( .A1(n19105), .A2(n15456), .ZN(n9991) );
  INV_X1 U12180 ( .A(n18982), .ZN(n9993) );
  NOR2_X1 U12181 ( .A1(n18992), .A2(n19105), .ZN(n18980) );
  INV_X1 U12182 ( .A(n19017), .ZN(n9995) );
  NOR2_X1 U12183 ( .A1(n19105), .A2(n12791), .ZN(n19018) );
  NOR2_X1 U12184 ( .A1(n19018), .A2(n19017), .ZN(n19016) );
  INV_X1 U12185 ( .A(n19101), .ZN(n19131) );
  AND2_X1 U12186 ( .A1(n11731), .A2(n11730), .ZN(n19021) );
  OR2_X1 U12187 ( .A1(n19980), .A2(n12820), .ZN(n19133) );
  AND2_X1 U12188 ( .A1(n19980), .A2(n12812), .ZN(n19122) );
  NAND2_X1 U12189 ( .A1(n10144), .A2(n9689), .ZN(n13817) );
  INV_X1 U12190 ( .A(n13708), .ZN(n10144) );
  OR2_X1 U12191 ( .A1(n12440), .A2(n12439), .ZN(n13709) );
  OR2_X1 U12192 ( .A1(n12423), .A2(n12422), .ZN(n13667) );
  OR2_X1 U12193 ( .A1(n12403), .A2(n12402), .ZN(n13620) );
  NOR2_X1 U12194 ( .A1(n13511), .A2(n13510), .ZN(n13512) );
  AND2_X1 U12195 ( .A1(n9692), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10133) );
  OR2_X1 U12196 ( .A1(n12351), .A2(n12350), .ZN(n13348) );
  CLKBUF_X1 U12197 ( .A(n13509), .Z(n13508) );
  INV_X1 U12198 ( .A(n15312), .ZN(n15298) );
  CLKBUF_X1 U12199 ( .A(n13218), .Z(n13217) );
  OR2_X1 U12200 ( .A1(n15269), .A2(n12978), .ZN(n15312) );
  INV_X1 U12201 ( .A(n10128), .ZN(n15252) );
  NOR2_X1 U12202 ( .A1(n15274), .A2(n14319), .ZN(n15263) );
  INV_X1 U12203 ( .A(n15381), .ZN(n16235) );
  NAND2_X1 U12204 ( .A1(n13256), .A2(n13257), .ZN(n13584) );
  AND2_X1 U12205 ( .A1(n15381), .A2(n13855), .ZN(n19196) );
  INV_X1 U12206 ( .A(n19961), .ZN(n19297) );
  INV_X1 U12207 ( .A(n16237), .ZN(n19189) );
  NOR2_X1 U12208 ( .A1(n19197), .A2(n19982), .ZN(n19211) );
  CLKBUF_X1 U12210 ( .A(n19211), .Z(n19228) );
  AND2_X1 U12211 ( .A1(n12905), .A2(n11551), .ZN(n12963) );
  NAND2_X1 U12212 ( .A1(n13022), .A2(n12920), .ZN(n12982) );
  NAND2_X1 U12213 ( .A1(n9990), .A2(n11847), .ZN(n9986) );
  INV_X1 U12214 ( .A(n15497), .ZN(n19004) );
  AND2_X1 U12215 ( .A1(n11834), .A2(n15534), .ZN(n15542) );
  NAND2_X1 U12216 ( .A1(n13938), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13937) );
  NAND2_X1 U12217 ( .A1(n11818), .A2(n11817), .ZN(n9852) );
  NAND2_X1 U12218 ( .A1(n12916), .A2(n11838), .ZN(n16310) );
  AND2_X1 U12219 ( .A1(n16310), .A2(n13109), .ZN(n16301) );
  AND2_X1 U12220 ( .A1(n12283), .A2(n19970), .ZN(n19236) );
  NAND2_X1 U12221 ( .A1(n15396), .A2(n9798), .ZN(n9797) );
  AOI21_X1 U12222 ( .B1(n15479), .B2(n15467), .A(n15480), .ZN(n15470) );
  INV_X1 U12223 ( .A(n9915), .ZN(n15517) );
  NAND2_X1 U12224 ( .A1(n9904), .A2(n9906), .ZN(n15744) );
  INV_X1 U12225 ( .A(n15779), .ZN(n9909) );
  NOR2_X1 U12226 ( .A1(n13145), .A2(n9958), .ZN(n13785) );
  NAND2_X1 U12227 ( .A1(n9961), .A2(n9960), .ZN(n9958) );
  NAND2_X1 U12228 ( .A1(n9957), .A2(n9961), .ZN(n13564) );
  INV_X1 U12229 ( .A(n19952), .ZN(n19949) );
  INV_X1 U12230 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19946) );
  INV_X1 U12231 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19938) );
  NOR2_X1 U12232 ( .A1(n13145), .A2(n12318), .ZN(n13493) );
  NAND2_X1 U12233 ( .A1(n15823), .A2(n13132), .ZN(n12972) );
  XNOR2_X1 U12234 ( .A(n13123), .B(n13122), .ZN(n19952) );
  NAND2_X1 U12235 ( .A1(n13202), .A2(n13137), .ZN(n19934) );
  CLKBUF_X1 U12236 ( .A(n12264), .Z(n12265) );
  OR2_X1 U12237 ( .A1(n19341), .A2(n19466), .ZN(n19360) );
  AND2_X1 U12238 ( .A1(n19409), .A2(n19408), .ZN(n19415) );
  INV_X1 U12239 ( .A(n19415), .ZN(n19432) );
  OR3_X1 U12240 ( .A1(n19467), .A2(n19466), .A3(n19465), .ZN(n19486) );
  AND2_X1 U12241 ( .A1(n19489), .A2(n10178), .ZN(n19485) );
  INV_X1 U12242 ( .A(n19513), .ZN(n19516) );
  AND2_X1 U12243 ( .A1(n19489), .A2(n19931), .ZN(n19544) );
  OAI21_X1 U12244 ( .B1(n19556), .B2(n19555), .A(n19554), .ZN(n19573) );
  INV_X1 U12245 ( .A(n19642), .ZN(n19626) );
  OR2_X1 U12246 ( .A1(n19651), .A2(n19650), .ZN(n19678) );
  INV_X1 U12247 ( .A(n19668), .ZN(n19677) );
  AND2_X1 U12248 ( .A1(n19606), .A2(n10178), .ZN(n19745) );
  OAI22_X1 U12249 ( .A1(n20279), .A2(n19283), .B1(n19282), .B2(n19281), .ZN(
        n19754) );
  OAI21_X1 U12250 ( .B1(n19726), .B2(n19725), .A(n19724), .ZN(n19762) );
  INV_X1 U12251 ( .A(n19623), .ZN(n19784) );
  INV_X1 U12252 ( .A(n19694), .ZN(n19805) );
  INV_X1 U12253 ( .A(n19699), .ZN(n19812) );
  AND2_X1 U12254 ( .A1(n19606), .A2(n19931), .ZN(n19820) );
  INV_X1 U12255 ( .A(n19672), .ZN(n19819) );
  INV_X1 U12256 ( .A(n19820), .ZN(n19842) );
  INV_X1 U12257 ( .A(n19768), .ZN(n19837) );
  AND2_X1 U12258 ( .A1(n19714), .A2(n19931), .ZN(n19838) );
  AND2_X1 U12259 ( .A1(n11220), .A2(n19957), .ZN(n19968) );
  INV_X1 U12260 ( .A(n17484), .ZN(n17483) );
  NAND2_X1 U12261 ( .A1(n18764), .A2(n18927), .ZN(n16556) );
  AND2_X1 U12262 ( .A1(n16671), .A2(n12005), .ZN(n16663) );
  NOR2_X1 U12263 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16719), .ZN(n16707) );
  AOI211_X1 U12264 ( .C1(n11995), .C2(n9894), .A(n9889), .B(n9890), .ZN(n9888)
         );
  INV_X1 U12265 ( .A(n9891), .ZN(n9890) );
  NOR2_X1 U12266 ( .A1(n11995), .A2(n9892), .ZN(n9889) );
  NOR2_X1 U12267 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16796), .ZN(n16778) );
  NOR2_X1 U12268 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16808), .ZN(n16807) );
  INV_X1 U12269 ( .A(n16922), .ZN(n16885) );
  NAND3_X1 U12270 ( .A1(n18946), .A2(n16913), .A3(n12139), .ZN(n16937) );
  INV_X1 U12271 ( .A(n16891), .ZN(n16934) );
  NAND2_X1 U12272 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17051), .ZN(n17004) );
  NOR2_X1 U12273 ( .A1(n18294), .A2(n17065), .ZN(n17051) );
  NAND2_X1 U12274 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17082), .ZN(n17065) );
  INV_X1 U12275 ( .A(n17094), .ZN(n17068) );
  INV_X1 U12276 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17256) );
  NOR2_X1 U12277 ( .A1(n14067), .A2(n17263), .ZN(n17258) );
  NAND2_X1 U12278 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17258), .ZN(n17257) );
  NOR2_X2 U12279 ( .A1(n14067), .A2(n17291), .ZN(n17282) );
  NAND2_X1 U12280 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17318), .ZN(n17313) );
  NOR2_X1 U12281 ( .A1(n17507), .A2(n17322), .ZN(n17318) );
  INV_X1 U12282 ( .A(n17327), .ZN(n17323) );
  NAND2_X1 U12283 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17323), .ZN(n17322) );
  INV_X1 U12284 ( .A(n17291), .ZN(n18294) );
  INV_X1 U12285 ( .A(n17365), .ZN(n17360) );
  NOR2_X1 U12286 ( .A1(n18294), .A2(n17372), .ZN(n17366) );
  INV_X1 U12287 ( .A(n17369), .ZN(n17370) );
  INV_X1 U12288 ( .A(n17363), .ZN(n17371) );
  NAND2_X1 U12289 ( .A1(n17290), .A2(n17289), .ZN(n17382) );
  NOR2_X1 U12290 ( .A1(n17380), .A2(n17288), .ZN(n17289) );
  NOR2_X1 U12291 ( .A1(n12593), .A2(n12592), .ZN(n12594) );
  NOR3_X1 U12292 ( .A1(n17521), .A2(n17440), .A3(n17414), .ZN(n17436) );
  NAND2_X1 U12293 ( .A1(n15991), .A2(n15994), .ZN(n17437) );
  NOR3_X1 U12294 ( .A1(n15988), .A2(n18267), .A3(n15987), .ZN(n15989) );
  AOI21_X1 U12295 ( .B1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B2(n9630), .A(
        n12652), .ZN(n12653) );
  INV_X1 U12296 ( .A(n17441), .ZN(n17414) );
  INV_X1 U12297 ( .A(n17437), .ZN(n17439) );
  NOR2_X1 U12298 ( .A1(n18932), .A2(n17548), .ZN(n17540) );
  OAI211_X1 U12299 ( .C1(n18932), .C2(n18933), .A(n17485), .B(n17484), .ZN(
        n17545) );
  BUF_X1 U12300 ( .A(n17545), .Z(n17548) );
  AND2_X1 U12302 ( .A1(n17718), .A2(n9842), .ZN(n17571) );
  INV_X1 U12303 ( .A(n17917), .ZN(n9842) );
  INV_X1 U12304 ( .A(n17718), .ZN(n17587) );
  INV_X1 U12305 ( .A(n17562), .ZN(n11997) );
  NAND2_X1 U12306 ( .A1(n16710), .A2(n10169), .ZN(n17663) );
  AND2_X1 U12307 ( .A1(n17774), .A2(n16442), .ZN(n17718) );
  NOR2_X1 U12308 ( .A1(n9701), .A2(n9881), .ZN(n9880) );
  INV_X1 U12309 ( .A(n17749), .ZN(n9881) );
  INV_X1 U12310 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17755) );
  NAND2_X1 U12311 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17909), .ZN(n17754) );
  NOR2_X2 U12312 ( .A1(n17915), .A2(n17415), .ZN(n17810) );
  INV_X1 U12313 ( .A(n17774), .ZN(n17813) );
  AND2_X1 U12314 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17816) );
  INV_X1 U12315 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17821) );
  INV_X1 U12316 ( .A(n17758), .ZN(n17828) );
  INV_X1 U12317 ( .A(n17810), .ZN(n17831) );
  INV_X1 U12318 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17834) );
  NAND2_X1 U12319 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17873) );
  INV_X1 U12320 ( .A(n18304), .ZN(n18592) );
  NOR2_X1 U12321 ( .A1(n18932), .A2(n16556), .ZN(n17905) );
  INV_X1 U12322 ( .A(n9659), .ZN(n17915) );
  OAI21_X1 U12323 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18926), .A(n16556), 
        .ZN(n17912) );
  AOI21_X1 U12324 ( .B1(n16436), .B2(n10151), .A(n16435), .ZN(n16441) );
  AOI21_X1 U12325 ( .B1(n17994), .B2(n17561), .A(n17553), .ZN(n16443) );
  AND2_X1 U12326 ( .A1(n12127), .A2(n9845), .ZN(n18740) );
  INV_X1 U12327 ( .A(n18720), .ZN(n9845) );
  INV_X1 U12328 ( .A(n12690), .ZN(n17602) );
  AND2_X1 U12329 ( .A1(n18740), .A2(n18721), .ZN(n18138) );
  OAI221_X1 U12330 ( .B1(n15918), .B2(n18756), .C1(n15918), .C2(n15917), .A(
        n18927), .ZN(n18161) );
  NOR2_X1 U12331 ( .A1(n17860), .A2(n12670), .ZN(n17847) );
  NAND2_X1 U12332 ( .A1(n18128), .A2(n18138), .ZN(n18200) );
  INV_X1 U12333 ( .A(n18248), .ZN(n18240) );
  INV_X1 U12334 ( .A(n18740), .ZN(n18717) );
  INV_X1 U12335 ( .A(n18161), .ZN(n18243) );
  NOR2_X1 U12336 ( .A1(n18757), .A2(n18161), .ZN(n18248) );
  INV_X1 U12337 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18743) );
  INV_X1 U12338 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18761) );
  INV_X1 U12339 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18763) );
  CLKBUF_X1 U12340 ( .A(n12022), .Z(n18912) );
  INV_X1 U12341 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18905) );
  INV_X1 U12342 ( .A(n18910), .ZN(n18913) );
  OAI211_X1 U12343 ( .C1(n18781), .C2(n18766), .A(n18266), .B(n15897), .ZN(
        n18910) );
  INV_X1 U12344 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18605) );
  CLKBUF_X1 U12345 ( .A(n16529), .Z(n16539) );
  AOI21_X1 U12346 ( .B1(n11195), .B2(n11194), .A(n11193), .ZN(n11196) );
  NOR2_X1 U12347 ( .A1(n14778), .A2(n11192), .ZN(n11193) );
  AOI21_X1 U12348 ( .B1(n10171), .B2(n11194), .A(n12837), .ZN(n12838) );
  OAI21_X1 U12349 ( .B1(n15025), .B2(n20007), .A(n9820), .ZN(P1_U2968) );
  AOI21_X1 U12350 ( .B1(n14487), .B2(n20239), .A(n9821), .ZN(n9820) );
  INV_X1 U12351 ( .A(n12258), .ZN(n9821) );
  OAI21_X1 U12352 ( .B1(n15025), .B2(n20222), .A(n9832), .ZN(P1_U3000) );
  NAND2_X1 U12353 ( .A1(n12829), .A2(n10148), .ZN(n12830) );
  AOI21_X1 U12354 ( .B1(n19148), .B2(n16324), .A(n9962), .ZN(n14179) );
  NAND2_X1 U12355 ( .A1(n10176), .A2(n14176), .ZN(n9962) );
  AOI21_X1 U12356 ( .B1(n12558), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12557), .ZN(n12559) );
  INV_X1 U12357 ( .A(n12596), .ZN(n17217) );
  OR2_X1 U12358 ( .A1(n14002), .A2(n10117), .ZN(n14688) );
  NOR2_X1 U12359 ( .A1(n15448), .A2(n10038), .ZN(n15434) );
  AND2_X1 U12360 ( .A1(n9985), .A2(n12794), .ZN(n9678) );
  INV_X2 U12361 ( .A(n12853), .ZN(n19105) );
  NAND2_X1 U12362 ( .A1(n14545), .A2(n14546), .ZN(n12833) );
  AND2_X1 U12363 ( .A1(n16221), .A2(n12796), .ZN(n9679) );
  NAND2_X1 U12364 ( .A1(n14595), .A2(n14596), .ZN(n14570) );
  NAND2_X1 U12365 ( .A1(n14648), .A2(n14649), .ZN(n14636) );
  NAND2_X1 U12366 ( .A1(n14595), .A2(n10123), .ZN(n14556) );
  INV_X1 U12367 ( .A(n10092), .ZN(n10090) );
  NOR2_X1 U12368 ( .A1(n10093), .A2(n16269), .ZN(n10092) );
  AND2_X1 U12369 ( .A1(n12328), .A2(n11657), .ZN(n11664) );
  AND4_X1 U12370 ( .A1(n11561), .A2(n11560), .A3(n11559), .A4(n11558), .ZN(
        n9681) );
  NAND2_X1 U12371 ( .A1(n10037), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15445) );
  NAND2_X1 U12372 ( .A1(n14648), .A2(n9735), .ZN(n14625) );
  NAND2_X1 U12373 ( .A1(n13743), .A2(n9752), .ZN(n10629) );
  AND2_X1 U12374 ( .A1(n10108), .A2(n10629), .ZN(n9682) );
  AND2_X1 U12375 ( .A1(n10170), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9683) );
  OR2_X1 U12376 ( .A1(n10442), .A2(n10110), .ZN(n9684) );
  AND2_X1 U12377 ( .A1(n9961), .A2(n9959), .ZN(n9686) );
  INV_X1 U12378 ( .A(n13736), .ZN(n16306) );
  NAND3_X1 U12379 ( .A1(n19939), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19781), 
        .ZN(n13736) );
  OR2_X1 U12380 ( .A1(n12774), .A2(n11845), .ZN(n9687) );
  AND2_X1 U12381 ( .A1(n15782), .A2(n9737), .ZN(n12857) );
  OR2_X1 U12382 ( .A1(n12774), .A2(n9998), .ZN(n9688) );
  AND2_X1 U12383 ( .A1(n15761), .A2(n15777), .ZN(n9908) );
  OR2_X1 U12384 ( .A1(n18976), .A2(n9755), .ZN(n9953) );
  AND2_X1 U12385 ( .A1(n13709), .A2(n13710), .ZN(n9689) );
  NOR2_X1 U12386 ( .A1(n12318), .A2(n9763), .ZN(n9961) );
  OR3_X1 U12387 ( .A1(n14338), .A2(n14337), .A3(n15265), .ZN(n9690) );
  AND2_X1 U12388 ( .A1(n17558), .A2(n16419), .ZN(n9691) );
  NOR2_X1 U12389 ( .A1(n9994), .A2(n15512), .ZN(n15228) );
  INV_X1 U12390 ( .A(n10051), .ZN(n13204) );
  AND2_X1 U12391 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9692) );
  AND2_X1 U12392 ( .A1(n10044), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9693) );
  OR2_X1 U12393 ( .A1(n13891), .A2(n13923), .ZN(n9694) );
  NOR3_X1 U12394 ( .A1(n18728), .A2(n12014), .A3(n18897), .ZN(n12088) );
  INV_X2 U12395 ( .A(n12088), .ZN(n17208) );
  AND2_X2 U12396 ( .A1(n9654), .A2(n16338), .ZN(n11288) );
  OR2_X1 U12397 ( .A1(n9694), .A2(n10063), .ZN(n9695) );
  NAND2_X1 U12398 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12673), .ZN(
        n9696) );
  AND2_X1 U12399 ( .A1(n11783), .A2(n15418), .ZN(n9697) );
  AND2_X1 U12400 ( .A1(n12974), .A2(n9632), .ZN(n12473) );
  OR2_X1 U12401 ( .A1(n12662), .A2(n12661), .ZN(n9698) );
  NAND2_X1 U12402 ( .A1(n15553), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15554) );
  NOR2_X1 U12403 ( .A1(n13797), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9700) );
  NAND2_X1 U12404 ( .A1(n11685), .A2(n11792), .ZN(n11695) );
  NOR2_X1 U12405 ( .A1(n14002), .A2(n10114), .ZN(n14689) );
  INV_X1 U12406 ( .A(n11099), .ZN(n14490) );
  NAND2_X1 U12407 ( .A1(n15488), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15472) );
  INV_X1 U12408 ( .A(n11836), .ZN(n15426) );
  AND3_X1 U12409 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12784) );
  INV_X1 U12410 ( .A(n11398), .ZN(n12978) );
  OR2_X1 U12411 ( .A1(n16800), .A2(n9884), .ZN(n9701) );
  NOR2_X1 U12412 ( .A1(n16281), .A2(n13944), .ZN(n9702) );
  AND4_X1 U12413 ( .A1(n9826), .A2(n9825), .A3(n9823), .A4(n9822), .ZN(n9703)
         );
  OR2_X1 U12414 ( .A1(n14517), .A2(n20086), .ZN(n9704) );
  OAI211_X1 U12415 ( .C1(n12562), .C2(n17234), .A(n12043), .B(n12042), .ZN(
        n18267) );
  AND2_X1 U12416 ( .A1(n10094), .A2(n9702), .ZN(n9706) );
  OR2_X1 U12417 ( .A1(n11768), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n9707) );
  NAND2_X1 U12418 ( .A1(n9874), .A2(n9697), .ZN(n12259) );
  AND2_X1 U12419 ( .A1(n15267), .A2(n15266), .ZN(n15210) );
  XOR2_X1 U12420 ( .A(n14196), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .Z(
        n9708) );
  NAND2_X1 U12421 ( .A1(n10134), .A2(n13201), .ZN(n13202) );
  NAND2_X1 U12422 ( .A1(n11836), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15412) );
  AND2_X1 U12423 ( .A1(n9919), .A2(n9918), .ZN(n9710) );
  AND2_X1 U12424 ( .A1(n20910), .A2(n20271), .ZN(n9711) );
  OR3_X1 U12425 ( .A1(n11756), .A2(n15480), .A3(n15505), .ZN(n9712) );
  AND3_X1 U12426 ( .A1(n11574), .A2(n11575), .A3(n11573), .ZN(n9713) );
  INV_X1 U12427 ( .A(n15448), .ZN(n10037) );
  NAND2_X1 U12428 ( .A1(n10094), .A2(n10091), .ZN(n16267) );
  INV_X1 U12429 ( .A(n18932), .ZN(n15987) );
  AND3_X1 U12430 ( .A1(n11369), .A2(n16338), .A3(n11368), .ZN(n9714) );
  INV_X1 U12431 ( .A(n14195), .ZN(n9796) );
  NOR2_X1 U12432 ( .A1(n12880), .A2(n15461), .ZN(n14195) );
  NOR2_X1 U12433 ( .A1(n15263), .A2(n15262), .ZN(n9715) );
  NAND2_X1 U12434 ( .A1(n15334), .A2(n9972), .ZN(n9716) );
  NAND2_X1 U12435 ( .A1(n14972), .A2(n16114), .ZN(n9717) );
  NOR2_X1 U12436 ( .A1(n14195), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9718) );
  AND4_X1 U12437 ( .A1(n10083), .A2(n10082), .A3(n10081), .A4(n10080), .ZN(
        n9719) );
  AND2_X1 U12438 ( .A1(n11817), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9720) );
  AND4_X1 U12439 ( .A1(n12605), .A2(n12604), .A3(n12603), .A4(n12602), .ZN(
        n9721) );
  NOR3_X1 U12440 ( .A1(n12869), .A2(n15461), .A3(n15633), .ZN(n9722) );
  NOR2_X1 U12441 ( .A1(n10460), .A2(n10417), .ZN(n9723) );
  AND2_X1 U12442 ( .A1(n12791), .A2(n9995), .ZN(n9724) );
  NAND2_X1 U12443 ( .A1(n11710), .A2(n11709), .ZN(n11734) );
  NAND2_X1 U12444 ( .A1(n10395), .A2(n10394), .ZN(n10443) );
  INV_X1 U12445 ( .A(n10443), .ZN(n10110) );
  OAI21_X1 U12446 ( .B1(n14153), .B2(n14152), .A(n14154), .ZN(n14159) );
  OR2_X1 U12447 ( .A1(n11843), .A2(n19074), .ZN(n9725) );
  AND2_X1 U12448 ( .A1(n13781), .A2(n11816), .ZN(n9726) );
  NAND2_X1 U12449 ( .A1(n11439), .A2(n11438), .ZN(n11482) );
  NAND2_X1 U12450 ( .A1(n14183), .A2(n14181), .ZN(n9727) );
  OR2_X1 U12451 ( .A1(n11703), .A2(n10174), .ZN(n9728) );
  NAND2_X1 U12452 ( .A1(n15267), .A2(n10060), .ZN(n15209) );
  AND2_X1 U12453 ( .A1(n13124), .A2(n13118), .ZN(n13520) );
  OAI21_X1 U12454 ( .B1(n15254), .B2(n10130), .A(n10129), .ZN(n14398) );
  INV_X1 U12455 ( .A(n14398), .ZN(n10126) );
  NAND2_X1 U12456 ( .A1(n12126), .A2(n12125), .ZN(n18727) );
  INV_X1 U12457 ( .A(n18727), .ZN(n12127) );
  NAND2_X1 U12458 ( .A1(n11854), .A2(n10033), .ZN(n11853) );
  NOR2_X1 U12459 ( .A1(n9846), .A2(n12047), .ZN(n9729) );
  NOR2_X1 U12460 ( .A1(n14379), .A2(n10132), .ZN(n9730) );
  INV_X2 U12461 ( .A(n19265), .ZN(n11418) );
  INV_X2 U12462 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18897) );
  OR2_X1 U12463 ( .A1(n12152), .A2(n12151), .ZN(P3_U2640) );
  INV_X2 U12464 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n11444) );
  INV_X1 U12465 ( .A(n11900), .ZN(n11463) );
  NOR2_X2 U12466 ( .A1(n19288), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12315) );
  XNOR2_X1 U12467 ( .A(n10436), .B(n10435), .ZN(n13474) );
  NOR2_X1 U12468 ( .A1(n12782), .A2(n16309), .ZN(n12781) );
  INV_X1 U12469 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10183) );
  NAND2_X1 U12470 ( .A1(n12524), .A2(n11427), .ZN(n9732) );
  OR2_X1 U12471 ( .A1(n11747), .A2(n15684), .ZN(n9733) );
  NAND2_X1 U12472 ( .A1(n20267), .A2(n13315), .ZN(n13169) );
  NOR2_X1 U12473 ( .A1(n13708), .A2(n10145), .ZN(n13845) );
  NAND2_X1 U12474 ( .A1(n15782), .A2(n9964), .ZN(n12858) );
  NAND2_X1 U12475 ( .A1(n14004), .A2(n14003), .ZN(n14002) );
  NOR2_X1 U12476 ( .A1(n12789), .A2(n16253), .ZN(n12778) );
  NOR2_X1 U12477 ( .A1(n12776), .A2(n15545), .ZN(n12777) );
  NAND2_X1 U12478 ( .A1(n13893), .A2(n13892), .ZN(n13891) );
  INV_X1 U12479 ( .A(n12314), .ZN(n12476) );
  INV_X1 U12480 ( .A(n11664), .ZN(n9944) );
  NAND2_X1 U12481 ( .A1(n10124), .A2(n14152), .ZN(n9734) );
  AND2_X1 U12482 ( .A1(n10781), .A2(n14649), .ZN(n9735) );
  AND3_X1 U12483 ( .A1(n13372), .A2(n13373), .A3(n9812), .ZN(n13363) );
  NAND2_X1 U12484 ( .A1(n9858), .A2(n9856), .ZN(n11390) );
  NOR3_X1 U12485 ( .A1(n13355), .A2(n10049), .A3(n10047), .ZN(n13664) );
  AND2_X1 U12486 ( .A1(n15220), .A2(n15219), .ZN(n13990) );
  INV_X1 U12487 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20914) );
  NAND2_X1 U12488 ( .A1(n12780), .A2(n10007), .ZN(n12779) );
  AND2_X1 U12489 ( .A1(n12781), .A2(n11840), .ZN(n12780) );
  OAI211_X1 U12490 ( .C1(n12516), .C2(n12290), .A(n19288), .B(n12273), .ZN(
        n12521) );
  OR3_X1 U12491 ( .A1(n9694), .A2(n10064), .A3(n10066), .ZN(n9736) );
  AOI21_X1 U12492 ( .B1(n15205), .B2(n12794), .A(n9983), .ZN(n16209) );
  AND2_X1 U12493 ( .A1(n9965), .A2(n13506), .ZN(n9737) );
  NOR2_X1 U12494 ( .A1(n18980), .A2(n18982), .ZN(n18981) );
  OR2_X1 U12495 ( .A1(n15466), .A2(n15518), .ZN(n9738) );
  XNOR2_X1 U12496 ( .A(n11389), .B(n12969), .ZN(n12271) );
  INV_X1 U12497 ( .A(n15795), .ZN(n9868) );
  OR2_X1 U12498 ( .A1(n18757), .A2(n15916), .ZN(n9739) );
  OR2_X1 U12500 ( .A1(n11653), .A2(n11673), .ZN(n9946) );
  AND2_X1 U12501 ( .A1(n9733), .A2(n9914), .ZN(n9740) );
  AND2_X1 U12502 ( .A1(n9964), .A2(n9963), .ZN(n9741) );
  INV_X1 U12503 ( .A(n13747), .ZN(n11124) );
  INV_X1 U12504 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17699) );
  INV_X1 U12505 ( .A(n13632), .ZN(n20244) );
  NAND2_X1 U12506 ( .A1(n19275), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n9742) );
  INV_X1 U12507 ( .A(n18721), .ZN(n18751) );
  NAND2_X1 U12508 ( .A1(n18945), .A2(n15896), .ZN(n18721) );
  OR2_X1 U12509 ( .A1(n9816), .A2(n9815), .ZN(n9743) );
  OR2_X1 U12510 ( .A1(n14857), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9744) );
  INV_X1 U12511 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9920) );
  AND2_X1 U12512 ( .A1(n10169), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9745) );
  NOR2_X1 U12513 ( .A1(n18981), .A2(n19105), .ZN(n9746) );
  NAND2_X1 U12514 ( .A1(n10472), .A2(n10471), .ZN(n10474) );
  INV_X1 U12515 ( .A(n9907), .ZN(n9906) );
  NOR2_X1 U12516 ( .A1(n9910), .A2(n15462), .ZN(n9907) );
  AND2_X1 U12517 ( .A1(n9735), .A2(n10120), .ZN(n9747) );
  AND2_X1 U12518 ( .A1(n13201), .A2(n13135), .ZN(n9748) );
  INV_X1 U12519 ( .A(n9888), .ZN(n16862) );
  INV_X1 U12520 ( .A(n10426), .ZN(n11004) );
  INV_X1 U12521 ( .A(n11004), .ZN(n13628) );
  INV_X1 U12522 ( .A(n15302), .ZN(n15309) );
  NAND2_X1 U12523 ( .A1(n11855), .A2(n10087), .ZN(n10055) );
  NAND2_X1 U12524 ( .A1(n13270), .A2(n10162), .ZN(n13256) );
  NAND2_X1 U12525 ( .A1(n13219), .A2(n9692), .ZN(n13347) );
  INV_X1 U12526 ( .A(n10617), .ZN(n10107) );
  NOR3_X1 U12527 ( .A1(n13355), .A2(n10049), .A3(n13622), .ZN(n13623) );
  AND2_X1 U12528 ( .A1(n9925), .A2(n9924), .ZN(n9749) );
  NOR2_X1 U12529 ( .A1(n12774), .A2(n9996), .ZN(n12771) );
  INV_X1 U12530 ( .A(n15538), .ZN(n9897) );
  OR2_X1 U12531 ( .A1(n17815), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9750) );
  NOR2_X1 U12532 ( .A1(n13355), .A2(n13356), .ZN(n13357) );
  NOR2_X1 U12533 ( .A1(n13222), .A2(n13272), .ZN(n13271) );
  NOR2_X1 U12534 ( .A1(n12772), .A2(n15441), .ZN(n12793) );
  AND2_X1 U12535 ( .A1(n19275), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n9751) );
  AND2_X1 U12536 ( .A1(n13825), .A2(n10107), .ZN(n9752) );
  AND2_X1 U12537 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9753) );
  NOR2_X1 U12538 ( .A1(n12774), .A2(n10000), .ZN(n12773) );
  NOR2_X1 U12539 ( .A1(n19105), .A2(n9724), .ZN(n9994) );
  NOR2_X1 U12540 ( .A1(n17847), .A2(n17846), .ZN(n9754) );
  NAND2_X1 U12541 ( .A1(n11434), .A2(n11435), .ZN(n11854) );
  INV_X1 U12542 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19074) );
  OR2_X1 U12543 ( .A1(n15461), .A2(n15473), .ZN(n9755) );
  INV_X1 U12544 ( .A(n9990), .ZN(n9989) );
  NAND2_X1 U12545 ( .A1(n9753), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9990) );
  OR2_X1 U12546 ( .A1(n13355), .A2(n10049), .ZN(n9756) );
  AND2_X1 U12547 ( .A1(n14375), .A2(n14380), .ZN(n9757) );
  NAND2_X1 U12548 ( .A1(n10318), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10610) );
  INV_X1 U12549 ( .A(n10610), .ZN(n10684) );
  NAND2_X1 U12550 ( .A1(n10052), .A2(n10055), .ZN(n10051) );
  AND2_X1 U12551 ( .A1(n9936), .A2(n9935), .ZN(n9758) );
  AND2_X1 U12552 ( .A1(n10057), .A2(n10056), .ZN(n9759) );
  AND2_X1 U12553 ( .A1(n13219), .A2(n10133), .ZN(n9760) );
  AND2_X1 U12554 ( .A1(n13348), .A2(n10133), .ZN(n9761) );
  AND2_X1 U12555 ( .A1(n10055), .A2(n11854), .ZN(n9762) );
  AND2_X1 U12556 ( .A1(n12765), .A2(n9753), .ZN(n12799) );
  INV_X1 U12557 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10184) );
  AND4_X1 U12558 ( .A1(n12323), .A2(n12322), .A3(n12321), .A4(n12320), .ZN(
        n9763) );
  AND2_X1 U12559 ( .A1(n9885), .A2(n9883), .ZN(n16695) );
  INV_X1 U12560 ( .A(n19098), .ZN(n9809) );
  INV_X1 U12561 ( .A(n15253), .ZN(n10131) );
  AND2_X1 U12562 ( .A1(n12765), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12797) );
  AND2_X1 U12563 ( .A1(n12505), .A2(n12504), .ZN(n9764) );
  AND2_X1 U12564 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15829) );
  INV_X1 U12565 ( .A(n10160), .ZN(n10004) );
  AND2_X1 U12566 ( .A1(n10015), .A2(n9698), .ZN(n9765) );
  OR2_X1 U12567 ( .A1(n12240), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9766) );
  NAND2_X1 U12568 ( .A1(n17711), .A2(n9683), .ZN(n9887) );
  AND2_X1 U12569 ( .A1(n10039), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9767) );
  OR2_X1 U12570 ( .A1(n9766), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9768) );
  NAND2_X1 U12571 ( .A1(n17853), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17819) );
  AND2_X1 U12572 ( .A1(n11832), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9769) );
  AND2_X1 U12573 ( .A1(n9767), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9770) );
  INV_X1 U12574 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n9893) );
  INV_X1 U12575 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n9894) );
  INV_X1 U12576 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10019) );
  INV_X1 U12577 ( .A(n15061), .ZN(n9780) );
  INV_X1 U12578 ( .A(n15105), .ZN(n10044) );
  NAND2_X2 U12579 ( .A1(n18944), .A2(n18783), .ZN(n18140) );
  AOI22_X2 U12580 ( .A1(DATAI_16_), .A2(n20285), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20284), .ZN(n20734) );
  AOI22_X2 U12581 ( .A1(DATAI_19_), .A2(n20285), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20284), .ZN(n20746) );
  AOI221_X2 U12582 ( .B1(n18510), .B2(n18509), .C1(n18508), .C2(n18509), .A(
        n18507), .ZN(n18533) );
  AOI22_X2 U12583 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19292), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19291), .ZN(n19843) );
  NOR2_X2 U12584 ( .A1(n13853), .A2(n13736), .ZN(n19291) );
  NOR2_X2 U12585 ( .A1(n18883), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18653) );
  INV_X1 U12586 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18883) );
  AOI22_X2 U12587 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20284), .B1(DATAI_30_), 
        .B2(n20285), .ZN(n20823) );
  AOI21_X1 U12588 ( .B1(n9643), .B2(n16039), .A(n9776), .ZN(n16040) );
  NOR2_X2 U12589 ( .A1(n12244), .A2(n12243), .ZN(n14856) );
  NAND2_X1 U12590 ( .A1(n10424), .A2(n9779), .ZN(n10425) );
  INV_X1 U12591 ( .A(n10507), .ZN(n9781) );
  NAND3_X1 U12592 ( .A1(n10040), .A2(n10041), .A3(n9693), .ZN(n10043) );
  NAND2_X1 U12593 ( .A1(n9793), .A2(n9795), .ZN(n9785) );
  OAI211_X1 U12594 ( .C1(n9802), .C2(n15396), .A(n9799), .B(n9797), .ZN(n15578) );
  AND2_X1 U12595 ( .A1(n9708), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9798) );
  OAI21_X1 U12596 ( .B1(n9804), .B2(n9708), .A(n9800), .ZN(n9799) );
  NAND2_X1 U12597 ( .A1(n9804), .A2(n9803), .ZN(n9802) );
  INV_X1 U12598 ( .A(n9708), .ZN(n9803) );
  NAND2_X1 U12599 ( .A1(n16366), .A2(n9805), .ZN(n11419) );
  NAND2_X1 U12600 ( .A1(n9806), .A2(n11407), .ZN(n11454) );
  NAND2_X1 U12601 ( .A1(n12521), .A2(n19265), .ZN(n9806) );
  AOI21_X2 U12602 ( .B1(n9807), .B2(n9867), .A(n9712), .ZN(n15453) );
  NOR2_X2 U12603 ( .A1(n15794), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15459) );
  NAND3_X1 U12604 ( .A1(n11665), .A2(n12324), .A3(n11666), .ZN(n11660) );
  NAND2_X2 U12605 ( .A1(n9808), .A2(n11552), .ZN(n11666) );
  OAI21_X2 U12606 ( .B1(n10076), .B2(n10069), .A(n14355), .ZN(n9808) );
  NAND3_X1 U12607 ( .A1(n11621), .A2(n11822), .A3(n15461), .ZN(n9810) );
  AND2_X2 U12608 ( .A1(n9895), .A2(n13680), .ZN(n11504) );
  AND2_X2 U12609 ( .A1(n15859), .A2(n19138), .ZN(n9895) );
  AOI21_X2 U12610 ( .B1(n15440), .B2(n15439), .A(n9722), .ZN(n15431) );
  NAND2_X1 U12611 ( .A1(n9811), .A2(n10566), .ZN(n13652) );
  NAND2_X1 U12612 ( .A1(n13372), .A2(n13373), .ZN(n13378) );
  INV_X1 U12613 ( .A(n13377), .ZN(n9812) );
  INV_X1 U12614 ( .A(n13364), .ZN(n10550) );
  NAND2_X1 U12615 ( .A1(n13363), .A2(n13365), .ZN(n13364) );
  OAI21_X1 U12616 ( .B1(n13743), .B2(n10107), .A(n10105), .ZN(n9816) );
  NAND2_X1 U12617 ( .A1(n9819), .A2(n10432), .ZN(n10433) );
  NAND3_X1 U12618 ( .A1(n10475), .A2(n10425), .A3(n10684), .ZN(n9819) );
  AND3_X4 U12619 ( .A1(n13429), .A2(n13182), .A3(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10957) );
  AND2_X2 U12620 ( .A1(n13429), .A2(n9824), .ZN(n10981) );
  NAND2_X1 U12621 ( .A1(n10979), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n9825) );
  AND2_X2 U12622 ( .A1(n10183), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10189) );
  AND2_X2 U12623 ( .A1(n13425), .A2(n10192), .ZN(n10343) );
  NAND2_X1 U12624 ( .A1(n9834), .A2(n9827), .ZN(n9833) );
  NAND2_X1 U12625 ( .A1(n9831), .A2(n9828), .ZN(n9827) );
  NOR2_X1 U12626 ( .A1(n9744), .A2(n9829), .ZN(n9828) );
  NAND2_X1 U12627 ( .A1(n14856), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9834) );
  NOR2_X2 U12628 ( .A1(n16556), .A2(n15987), .ZN(n17902) );
  NAND2_X1 U12629 ( .A1(n9851), .A2(n9852), .ZN(n13938) );
  OAI211_X1 U12630 ( .C1(n9851), .C2(n13932), .A(n9850), .B(n11821), .ZN(
        n13951) );
  NAND2_X1 U12631 ( .A1(n10155), .A2(n11406), .ZN(n11455) );
  AND2_X2 U12632 ( .A1(n9855), .A2(n11548), .ZN(n11665) );
  NAND3_X1 U12633 ( .A1(n11527), .A2(n11528), .A3(n11526), .ZN(n9855) );
  AND2_X2 U12634 ( .A1(n10035), .A2(n10036), .ZN(n11836) );
  NAND4_X1 U12635 ( .A1(n9857), .A2(n11311), .A3(n11308), .A4(n11309), .ZN(
        n9856) );
  NAND4_X1 U12636 ( .A1(n9859), .A2(n11315), .A3(n11314), .A4(n11313), .ZN(
        n9858) );
  XNOR2_X2 U12637 ( .A(n11659), .B(n11660), .ZN(n11797) );
  NAND3_X1 U12638 ( .A1(n9866), .A2(n9865), .A3(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n9860) );
  NAND3_X1 U12639 ( .A1(n9866), .A2(n9865), .A3(n9864), .ZN(n9863) );
  OR2_X1 U12640 ( .A1(n11781), .A2(n9795), .ZN(n9873) );
  NAND2_X1 U12641 ( .A1(n11781), .A2(n9871), .ZN(n9870) );
  NAND2_X1 U12642 ( .A1(n11781), .A2(n11780), .ZN(n9874) );
  AOI21_X2 U12643 ( .B1(n9871), .B2(n9795), .A(n9727), .ZN(n9869) );
  AND2_X1 U12644 ( .A1(n9879), .A2(n9878), .ZN(n15420) );
  NAND2_X1 U12645 ( .A1(n9879), .A2(n9877), .ZN(n10099) );
  AND2_X1 U12646 ( .A1(n9878), .A2(n10096), .ZN(n9877) );
  NOR2_X2 U12647 ( .A1(n12011), .A2(n17565), .ZN(n12722) );
  INV_X1 U12648 ( .A(n17819), .ZN(n9882) );
  NAND3_X1 U12649 ( .A1(n9885), .A2(n9882), .A3(n9880), .ZN(n17739) );
  NAND3_X1 U12650 ( .A1(n9882), .A2(n9885), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16789) );
  INV_X1 U12651 ( .A(n9887), .ZN(n16710) );
  NAND3_X1 U12652 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n9892) );
  AND2_X2 U12653 ( .A1(n11508), .A2(n9895), .ZN(n11553) );
  OAI21_X1 U12654 ( .B1(n9646), .B2(n9902), .A(n9901), .ZN(n15541) );
  AOI21_X2 U12655 ( .B1(n9900), .B2(n9898), .A(n9896), .ZN(n15527) );
  INV_X1 U12656 ( .A(n9646), .ZN(n9900) );
  OR2_X2 U12657 ( .A1(n15516), .A2(n9738), .ZN(n9915) );
  AND2_X2 U12658 ( .A1(n9920), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10191) );
  NAND2_X1 U12659 ( .A1(n11098), .A2(n11097), .ZN(n9927) );
  AND2_X2 U12660 ( .A1(n14601), .A2(n9758), .ZN(n14549) );
  NOR3_X2 U12661 ( .A1(n9945), .A2(n11653), .A3(n9941), .ZN(n11684) );
  NAND2_X1 U12662 ( .A1(n9943), .A2(n9942), .ZN(n9941) );
  INV_X1 U12663 ( .A(n9946), .ZN(n11678) );
  INV_X1 U12664 ( .A(n11677), .ZN(n9945) );
  INV_X1 U12665 ( .A(n11734), .ZN(n9947) );
  NAND2_X1 U12666 ( .A1(n9947), .A2(n9948), .ZN(n11726) );
  NAND2_X1 U12667 ( .A1(n11695), .A2(n9950), .ZN(n11736) );
  NAND3_X1 U12668 ( .A1(n9733), .A2(n9956), .A3(n9953), .ZN(n11756) );
  INV_X1 U12669 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n9954) );
  INV_X1 U12670 ( .A(n13145), .ZN(n9957) );
  NAND2_X1 U12671 ( .A1(n9957), .A2(n9686), .ZN(n13783) );
  AND2_X1 U12672 ( .A1(n15337), .A2(n15336), .ZN(n15334) );
  NAND2_X1 U12673 ( .A1(n15337), .A2(n9971), .ZN(n12805) );
  NAND2_X1 U12674 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12783) );
  INV_X1 U12675 ( .A(n12783), .ZN(n9982) );
  NAND2_X1 U12676 ( .A1(n9982), .A2(n9981), .ZN(n12782) );
  AND2_X1 U12677 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n9981) );
  NOR2_X2 U12678 ( .A1(n9679), .A2(n19105), .ZN(n15205) );
  OR2_X1 U12679 ( .A1(n12765), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9988) );
  NAND3_X1 U12680 ( .A1(n9988), .A2(n9987), .A3(n9986), .ZN(n12763) );
  NAND3_X1 U12681 ( .A1(n12765), .A2(n9989), .A3(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n9987) );
  OR2_X1 U12682 ( .A1(n15192), .A2(n15195), .ZN(n15193) );
  NAND2_X1 U12683 ( .A1(n10002), .A2(n12794), .ZN(n12801) );
  OR2_X1 U12684 ( .A1(n15192), .A2(n10003), .ZN(n10002) );
  NAND2_X1 U12685 ( .A1(n15193), .A2(n12794), .ZN(n10005) );
  NOR2_X2 U12686 ( .A1(n17611), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17610) );
  NAND2_X2 U12687 ( .A1(n17703), .A2(n17815), .ZN(n17626) );
  NAND2_X1 U12688 ( .A1(n10012), .A2(n10011), .ZN(n10014) );
  NOR2_X1 U12689 ( .A1(n17876), .A2(n18216), .ZN(n10011) );
  INV_X1 U12690 ( .A(n17885), .ZN(n10012) );
  NOR2_X2 U12691 ( .A1(n17875), .A2(n12666), .ZN(n12669) );
  INV_X1 U12692 ( .A(n10015), .ZN(n17884) );
  NAND2_X1 U12693 ( .A1(n17840), .A2(n10150), .ZN(n12757) );
  INV_X1 U12694 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10018) );
  NAND3_X1 U12695 ( .A1(n10020), .A2(n17601), .A3(n9750), .ZN(n17586) );
  NAND4_X1 U12696 ( .A1(n10020), .A2(n17601), .A3(n9750), .A4(n10019), .ZN(
        n10023) );
  INV_X1 U12697 ( .A(n10023), .ZN(n17585) );
  NAND2_X1 U12698 ( .A1(n12014), .A2(n18897), .ZN(n10024) );
  NAND2_X2 U12699 ( .A1(n12022), .A2(n12023), .ZN(n16926) );
  XNOR2_X1 U12700 ( .A(n12676), .B(n12675), .ZN(n17842) );
  OAI21_X2 U12701 ( .B1(n17860), .B2(n10025), .A(n10026), .ZN(n12676) );
  NAND2_X1 U12702 ( .A1(n12695), .A2(n17558), .ZN(n15933) );
  NAND3_X4 U12703 ( .A1(n10030), .A2(n10029), .A3(n10028), .ZN(n15859) );
  NAND4_X1 U12704 ( .A1(n10032), .A2(n11486), .A3(n10084), .A4(n11853), .ZN(
        n10028) );
  NAND2_X2 U12705 ( .A1(n10031), .A2(n10085), .ZN(n10030) );
  NAND2_X1 U12706 ( .A1(n10087), .A2(n10084), .ZN(n10031) );
  NAND2_X1 U12707 ( .A1(n11437), .A2(n11436), .ZN(n10033) );
  NAND2_X2 U12708 ( .A1(n13780), .A2(n13777), .ZN(n13782) );
  XNOR2_X2 U12709 ( .A(n11665), .B(n11666), .ZN(n13487) );
  NAND2_X1 U12710 ( .A1(n15553), .A2(n9769), .ZN(n15532) );
  INV_X1 U12711 ( .A(n15532), .ZN(n11834) );
  INV_X1 U12712 ( .A(n15448), .ZN(n10035) );
  AND2_X1 U12713 ( .A1(n11836), .A2(n9767), .ZN(n15400) );
  NAND2_X1 U12714 ( .A1(n11836), .A2(n9770), .ZN(n14203) );
  OAI21_X1 U12715 ( .B1(n14009), .B2(n12238), .A(n12237), .ZN(n14964) );
  NAND3_X1 U12716 ( .A1(n10052), .A2(n13221), .A3(n10055), .ZN(n13222) );
  NAND2_X1 U12717 ( .A1(n12884), .A2(n9759), .ZN(n12809) );
  NAND2_X1 U12718 ( .A1(n15267), .A2(n10058), .ZN(n12883) );
  NAND2_X2 U12719 ( .A1(n11471), .A2(n11472), .ZN(n11485) );
  NAND2_X1 U12720 ( .A1(n11556), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10073) );
  NAND2_X1 U12721 ( .A1(n19771), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10074) );
  NAND4_X1 U12722 ( .A1(n9719), .A2(n9685), .A3(n10077), .A4(n11549), .ZN(
        n10076) );
  NAND2_X1 U12723 ( .A1(n11555), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10079) );
  NAND2_X1 U12724 ( .A1(n19613), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10083) );
  NAND2_X1 U12725 ( .A1(n11848), .A2(n11849), .ZN(n10084) );
  NAND2_X1 U12726 ( .A1(n10086), .A2(n11853), .ZN(n10085) );
  NAND2_X1 U12727 ( .A1(n11482), .A2(n11483), .ZN(n10086) );
  NAND2_X1 U12728 ( .A1(n11588), .A2(n10095), .ZN(n11822) );
  NAND2_X1 U12729 ( .A1(n11588), .A2(n11659), .ZN(n11620) );
  NAND3_X1 U12730 ( .A1(n12524), .A2(n11427), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n11900) );
  NAND2_X1 U12731 ( .A1(n15420), .A2(n15417), .ZN(n15406) );
  NAND2_X1 U12732 ( .A1(n10099), .A2(n11778), .ZN(n11781) );
  NOR2_X4 U12733 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10190) );
  NAND3_X1 U12734 ( .A1(n10322), .A2(n10310), .A3(n10309), .ZN(n10101) );
  NOR2_X1 U12735 ( .A1(n9711), .A2(n10102), .ZN(n10322) );
  OAI21_X2 U12736 ( .B1(n13325), .B2(n10103), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10328) );
  NAND2_X1 U12737 ( .A1(n10445), .A2(n20914), .ZN(n10441) );
  XNOR2_X2 U12738 ( .A(n10362), .B(n10361), .ZN(n10445) );
  NOR2_X1 U12739 ( .A1(n14002), .A2(n14702), .ZN(n14701) );
  INV_X1 U12740 ( .A(n14702), .ZN(n10118) );
  AND2_X2 U12741 ( .A1(n14648), .A2(n9747), .ZN(n14609) );
  INV_X1 U12743 ( .A(n15254), .ZN(n10125) );
  NAND2_X1 U12744 ( .A1(n9730), .A2(n10128), .ZN(n10127) );
  AND2_X2 U12745 ( .A1(n10127), .A2(n10126), .ZN(n15247) );
  INV_X1 U12746 ( .A(n13509), .ZN(n13513) );
  NAND2_X1 U12747 ( .A1(n13219), .A2(n9761), .ZN(n13509) );
  NAND2_X1 U12748 ( .A1(n13136), .A2(n13135), .ZN(n10135) );
  NAND3_X1 U12749 ( .A1(n10135), .A2(n13201), .A3(n13200), .ZN(n13210) );
  NAND2_X1 U12750 ( .A1(n13210), .A2(n13209), .ZN(n13218) );
  NAND3_X1 U12751 ( .A1(n10137), .A2(n9690), .A3(n10139), .ZN(n10136) );
  NAND2_X1 U12752 ( .A1(n15273), .A2(n15272), .ZN(n10139) );
  INV_X1 U12753 ( .A(n14319), .ZN(n10137) );
  INV_X2 U12754 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13763) );
  NOR2_X2 U12755 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11222) );
  INV_X2 U12756 ( .A(n11330), .ZN(n14399) );
  NOR2_X2 U12757 ( .A1(n13708), .A2(n10142), .ZN(n14270) );
  AOI21_X1 U12758 ( .B1(n15859), .B2(n13132), .A(n13131), .ZN(n13134) );
  AOI21_X1 U12759 ( .B1(n12684), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n12682), .ZN(n17704) );
  NAND2_X1 U12760 ( .A1(n12777), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12774) );
  NAND2_X1 U12761 ( .A1(n12895), .A2(n12870), .ZN(n15354) );
  AOI21_X1 U12762 ( .B1(n16186), .B2(n16331), .A(n14175), .ZN(n14176) );
  OAI211_X1 U12763 ( .C1(n14451), .C2(n15816), .A(n10175), .B(n14213), .ZN(
        n14214) );
  NAND2_X1 U12764 ( .A1(n12778), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12776) );
  INV_X1 U12765 ( .A(n11483), .ZN(n11848) );
  OAI21_X1 U12766 ( .B1(n11850), .B2(n11849), .A(n11848), .ZN(n11852) );
  CLKBUF_X1 U12767 ( .A(n13951), .Z(n16288) );
  NAND2_X1 U12768 ( .A1(n11276), .A2(n11973), .ZN(n11650) );
  NOR2_X1 U12769 ( .A1(n16926), .A2(n12021), .ZN(n12597) );
  AOI21_X1 U12770 ( .B1(n14526), .B2(n20239), .A(n14157), .ZN(n14158) );
  AND2_X2 U12771 ( .A1(n11684), .A2(n11689), .ZN(n11687) );
  INV_X2 U12772 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13182) );
  NAND2_X1 U12773 ( .A1(n10416), .A2(n20297), .ZN(n13476) );
  CLKBUF_X1 U12774 ( .A(n15488), .Z(n15680) );
  AND2_X1 U12775 ( .A1(n10362), .A2(n10360), .ZN(n10413) );
  OAI22_X2 U12776 ( .A1(n13415), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n12173), 
        .B2(n10460), .ZN(n10359) );
  NAND2_X1 U12777 ( .A1(n20289), .A2(n20280), .ZN(n13311) );
  AND2_X1 U12778 ( .A1(n14160), .A2(n20258), .ZN(n12214) );
  NAND2_X1 U12779 ( .A1(n20267), .A2(n20258), .ZN(n11099) );
  NOR2_X1 U12780 ( .A1(n13644), .A2(n13632), .ZN(n13640) );
  NAND2_X1 U12781 ( .A1(n13632), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10459) );
  NOR2_X1 U12782 ( .A1(n13632), .A2(n20914), .ZN(n10356) );
  OR2_X2 U12783 ( .A1(n13310), .A2(n13632), .ZN(n14492) );
  CLKBUF_X1 U12784 ( .A(n14270), .Z(n15287) );
  INV_X1 U12785 ( .A(n12651), .ZN(n12654) );
  NAND2_X1 U12786 ( .A1(n11834), .A2(n11833), .ZN(n15500) );
  NAND2_X1 U12787 ( .A1(n12196), .A2(n10684), .ZN(n10549) );
  OR2_X1 U12788 ( .A1(n13136), .A2(n9748), .ZN(n13137) );
  BUF_X1 U12789 ( .A(n11449), .Z(n13762) );
  NAND2_X1 U12790 ( .A1(n12509), .A2(n11415), .ZN(n11449) );
  INV_X1 U12791 ( .A(n10257), .ZN(n10235) );
  XNOR2_X1 U12792 ( .A(n11008), .B(n11007), .ZN(n14487) );
  XNOR2_X1 U12793 ( .A(n14450), .B(n14449), .ZN(n14460) );
  NAND2_X1 U12794 ( .A1(n15237), .A2(n14430), .ZN(n14450) );
  INV_X1 U12795 ( .A(n10434), .ZN(n10436) );
  NAND2_X1 U12796 ( .A1(n14355), .A2(n11388), .ZN(n11426) );
  OAI21_X2 U12797 ( .B1(n13141), .B2(n11856), .A(n11442), .ZN(n11483) );
  NAND2_X1 U12798 ( .A1(n14487), .A2(n10158), .ZN(n11087) );
  AND2_X1 U12799 ( .A1(n15859), .A2(n11520), .ZN(n11521) );
  INV_X1 U12800 ( .A(n15859), .ZN(n13138) );
  AND2_X1 U12801 ( .A1(n15859), .A2(n11509), .ZN(n11519) );
  AND2_X1 U12802 ( .A1(n11455), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10146) );
  INV_X1 U12803 ( .A(n15811), .ZN(n16331) );
  INV_X1 U12804 ( .A(n16324), .ZN(n15816) );
  INV_X1 U12805 ( .A(n14779), .ZN(n13662) );
  INV_X1 U12806 ( .A(n14777), .ZN(n11194) );
  AND3_X1 U12807 ( .A1(n20645), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10147) );
  INV_X1 U12808 ( .A(n13452), .ZN(n20135) );
  NOR2_X1 U12809 ( .A1(n12828), .A2(n12827), .ZN(n10148) );
  AND2_X1 U12810 ( .A1(n13640), .A2(n13636), .ZN(n20088) );
  NOR2_X1 U12811 ( .A1(n9677), .A2(n20241), .ZN(n10149) );
  OR2_X1 U12812 ( .A1(n12676), .A2(n12675), .ZN(n10150) );
  NOR2_X1 U12813 ( .A1(n16433), .A2(n10154), .ZN(n10151) );
  OR2_X1 U12814 ( .A1(n15975), .A2(n16419), .ZN(n10152) );
  AND2_X1 U12815 ( .A1(n18050), .A2(n17918), .ZN(n10153) );
  OR2_X1 U12816 ( .A1(n18757), .A2(n17415), .ZN(n10154) );
  NAND2_X1 U12817 ( .A1(n20914), .A2(n20243), .ZN(n20299) );
  AND2_X1 U12818 ( .A1(n12266), .A2(n11412), .ZN(n10155) );
  AND3_X1 U12819 ( .A1(n12619), .A2(n12618), .A3(n12617), .ZN(n10156) );
  AND2_X1 U12820 ( .A1(n12260), .A2(n14181), .ZN(n10157) );
  AND2_X1 U12821 ( .A1(n14853), .A2(n14161), .ZN(n10158) );
  AND2_X1 U12822 ( .A1(n12607), .A2(n10167), .ZN(n10159) );
  NOR2_X1 U12823 ( .A1(n12799), .A2(n12800), .ZN(n10160) );
  INV_X1 U12824 ( .A(n18870), .ZN(n18941) );
  AND2_X1 U12825 ( .A1(n11819), .A2(n13778), .ZN(n10161) );
  NAND2_X2 U12826 ( .A1(n14853), .A2(n13281), .ZN(n14848) );
  OR2_X1 U12827 ( .A1(n15461), .A2(n12336), .ZN(n10162) );
  NOR2_X1 U12828 ( .A1(n13624), .A2(n13623), .ZN(n10163) );
  AND2_X1 U12829 ( .A1(n11373), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10164) );
  AND3_X1 U12830 ( .A1(n12074), .A2(n12073), .A3(n12072), .ZN(n10165) );
  OR2_X1 U12831 ( .A1(n17217), .A2(n14082), .ZN(n10166) );
  OR2_X1 U12832 ( .A1(n17241), .A2(n18605), .ZN(n10167) );
  AND2_X1 U12833 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10168) );
  INV_X1 U12834 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11841) );
  INV_X1 U12835 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11846) );
  INV_X1 U12836 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12642) );
  AND2_X1 U12837 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10169) );
  AND2_X1 U12838 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10170) );
  INV_X1 U12839 ( .A(n10428), .ZN(n10905) );
  NOR2_X1 U12840 ( .A1(n14166), .A2(n12836), .ZN(n10171) );
  NAND2_X1 U12841 ( .A1(n19275), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10172) );
  INV_X1 U12842 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15557) );
  OR3_X1 U12843 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17644), .ZN(n10173) );
  AND2_X1 U12844 ( .A1(n11702), .A2(n11701), .ZN(n10174) );
  OR3_X1 U12845 ( .A1(n15570), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14207), .ZN(n10175) );
  OR4_X1 U12846 ( .A1(n15570), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14208), .A4(n14207), .ZN(n10176) );
  AND4_X1 U12847 ( .A1(n12612), .A2(n12611), .A3(n12610), .A4(n12609), .ZN(
        n10177) );
  NOR2_X1 U12848 ( .A1(n19942), .A2(n19952), .ZN(n10178) );
  NOR2_X1 U12849 ( .A1(n14572), .A2(n14585), .ZN(n10179) );
  NOR2_X2 U12850 ( .A1(n14203), .A2(n12287), .ZN(n14188) );
  OAI22_X1 U12851 ( .A1(n12763), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19987), 
        .B2(n12762), .ZN(n12853) );
  NOR2_X1 U12852 ( .A1(n18791), .A2(n17818), .ZN(n17664) );
  INV_X1 U12853 ( .A(n12766), .ZN(n12770) );
  AND2_X2 U12854 ( .A1(n13425), .A2(n15163), .ZN(n10348) );
  AND2_X2 U12855 ( .A1(n10191), .A2(n15163), .ZN(n13424) );
  AND4_X1 U12856 ( .A1(n10249), .A2(n10248), .A3(n10247), .A4(n10246), .ZN(
        n10181) );
  AND2_X2 U12857 ( .A1(n10189), .A2(n13431), .ZN(n10363) );
  AND4_X1 U12858 ( .A1(n10188), .A2(n10187), .A3(n10186), .A4(n10185), .ZN(
        n10182) );
  AOI22_X1 U12859 ( .A1(n19338), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11554), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U12860 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n10304), .B1(n11024), 
        .B2(n20258), .ZN(n11036) );
  OR2_X1 U12861 ( .A1(n11042), .A2(n10530), .ZN(n10542) );
  NAND2_X1 U12862 ( .A1(n11453), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11433) );
  AOI22_X1 U12863 ( .A1(n19338), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11554), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11498) );
  INV_X1 U12864 ( .A(n11024), .ZN(n11040) );
  NAND2_X1 U12865 ( .A1(n10542), .A2(n10541), .ZN(n10553) );
  NAND2_X1 U12866 ( .A1(n20289), .A2(n20271), .ZN(n10257) );
  NAND2_X1 U12867 ( .A1(n10332), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10316) );
  AOI22_X1 U12868 ( .A1(n11562), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11563), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11505) );
  INV_X1 U12869 ( .A(n11413), .ZN(n11391) );
  NAND2_X1 U12870 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20692), .ZN(
        n11026) );
  OR2_X1 U12871 ( .A1(n10519), .A2(n10518), .ZN(n12198) );
  INV_X1 U12872 ( .A(n10553), .ZN(n10554) );
  OR2_X1 U12873 ( .A1(n10540), .A2(n10539), .ZN(n12207) );
  NAND2_X1 U12874 ( .A1(n13311), .A2(n10257), .ZN(n10297) );
  OAI21_X1 U12875 ( .B1(n16287), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n16285), .ZN(n11824) );
  NAND2_X1 U12876 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12070) );
  OR2_X1 U12877 ( .A1(n12710), .A2(n12706), .ZN(n12128) );
  INV_X1 U12878 ( .A(n10297), .ZN(n10298) );
  INV_X1 U12879 ( .A(n14637), .ZN(n10781) );
  INV_X1 U12880 ( .A(n10547), .ZN(n10548) );
  OR2_X1 U12881 ( .A1(n10408), .A2(n10407), .ZN(n12158) );
  INV_X1 U12882 ( .A(n11046), .ZN(n11042) );
  INV_X1 U12883 ( .A(n14357), .ZN(n14358) );
  NAND2_X1 U12884 ( .A1(n11792), .A2(n11736), .ZN(n11710) );
  OR2_X1 U12885 ( .A1(n11984), .A2(n11979), .ZN(n11980) );
  OAI21_X1 U12886 ( .B1(n17163), .B2(n17034), .A(n12070), .ZN(n12071) );
  OAI21_X1 U12887 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n12023), .A(
        n12128), .ZN(n12133) );
  NAND2_X1 U12888 ( .A1(n10521), .A2(n10520), .ZN(n10552) );
  OR2_X1 U12889 ( .A1(n14483), .A2(n14471), .ZN(n11064) );
  NOR2_X1 U12890 ( .A1(n10931), .A2(n10930), .ZN(n10932) );
  AND2_X1 U12891 ( .A1(n10877), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10886) );
  NOR2_X1 U12892 ( .A1(n10775), .A2(n10774), .ZN(n10776) );
  INV_X1 U12893 ( .A(n10630), .ZN(n10645) );
  OR2_X1 U12894 ( .A1(n10470), .A2(n10469), .ZN(n12180) );
  AND2_X1 U12895 ( .A1(n11117), .A2(n11116), .ZN(n13656) );
  INV_X1 U12896 ( .A(n13311), .ZN(n13328) );
  NOR2_X1 U12897 ( .A1(n11426), .A2(n11425), .ZN(n11427) );
  AND2_X1 U12898 ( .A1(n14378), .A2(n9757), .ZN(n14379) );
  AND2_X1 U12899 ( .A1(n11829), .A2(n16284), .ZN(n11830) );
  INV_X1 U12900 ( .A(n12473), .ZN(n12336) );
  INV_X1 U12901 ( .A(n17654), .ZN(n12003) );
  INV_X1 U12902 ( .A(n12071), .ZN(n12072) );
  AND2_X1 U12903 ( .A1(n17815), .A2(n12679), .ZN(n12680) );
  NOR2_X1 U12904 ( .A1(n14684), .A2(n14683), .ZN(n14653) );
  NOR2_X1 U12905 ( .A1(n12253), .A2(n14515), .ZN(n12255) );
  NAND2_X1 U12906 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10293) );
  AND2_X1 U12907 ( .A1(n20837), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11005) );
  AOI22_X1 U12908 ( .A1(n10974), .A2(n10973), .B1(n13628), .B2(n14528), .ZN(
        n14152) );
  NAND2_X1 U12909 ( .A1(n10886), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10909) );
  AND2_X1 U12910 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n10738), .ZN(
        n10739) );
  OR2_X1 U12911 ( .A1(n15116), .A2(n15006), .ZN(n15086) );
  INV_X1 U12912 ( .A(n14490), .ZN(n11155) );
  AND2_X1 U12913 ( .A1(n11128), .A2(n11127), .ZN(n13826) );
  NAND2_X1 U12914 ( .A1(n13177), .A2(n9636), .ZN(n11065) );
  NAND2_X1 U12915 ( .A1(n13330), .A2(n13328), .ZN(n13324) );
  INV_X1 U12916 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15521) );
  AND2_X1 U12917 ( .A1(n11882), .A2(n11881), .ZN(n13356) );
  AND2_X1 U12918 ( .A1(n12904), .A2(n19985), .ZN(n12917) );
  NOR2_X2 U12919 ( .A1(n12883), .A2(n12885), .ZN(n12884) );
  XNOR2_X1 U12920 ( .A(n11483), .B(n11482), .ZN(n11488) );
  NOR2_X1 U12921 ( .A1(n12803), .A2(n12802), .ZN(n12806) );
  OR2_X1 U12922 ( .A1(n15615), .A2(n12548), .ZN(n15583) );
  AND2_X1 U12923 ( .A1(n19934), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19932) );
  AND2_X1 U12924 ( .A1(n11984), .A2(n13026), .ZN(n11985) );
  NAND2_X1 U12925 ( .A1(n17657), .A2(n18000), .ZN(n17644) );
  NOR2_X1 U12926 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n10022), .ZN(
        n17690) );
  NOR2_X1 U12927 ( .A1(n10022), .A2(n12757), .ZN(n17783) );
  NOR2_X1 U12928 ( .A1(n17891), .A2(n12659), .ZN(n12662) );
  OR2_X1 U12929 ( .A1(n14656), .A2(n14951), .ZN(n14643) );
  NOR2_X1 U12930 ( .A1(n20044), .A2(n14497), .ZN(n15995) );
  INV_X1 U12931 ( .A(n13870), .ZN(n20028) );
  INV_X1 U12932 ( .A(n20091), .ZN(n20067) );
  INV_X1 U12933 ( .A(n20916), .ZN(n13644) );
  AND2_X1 U12934 ( .A1(n11130), .A2(n11129), .ZN(n14000) );
  INV_X1 U12935 ( .A(n20238), .ZN(n20237) );
  NAND2_X1 U12936 ( .A1(n10739), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10775) );
  INV_X1 U12937 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14696) );
  NOR2_X1 U12938 ( .A1(n10607), .A2(n10606), .ZN(n10612) );
  AND3_X1 U12939 ( .A1(n10579), .A2(n10578), .A3(n10577), .ZN(n13693) );
  NAND2_X1 U12940 ( .A1(n20007), .A2(n12249), .ZN(n13067) );
  AND2_X1 U12941 ( .A1(n15164), .A2(n11089), .ZN(n14474) );
  OR2_X1 U12942 ( .A1(n20240), .A2(n10474), .ZN(n20431) );
  NOR2_X1 U12943 ( .A1(n20400), .A2(n20299), .ZN(n20577) );
  INV_X1 U12944 ( .A(n20240), .ZN(n15155) );
  AND2_X1 U12945 ( .A1(n20579), .A2(n20406), .ZN(n20729) );
  NAND2_X1 U12946 ( .A1(n11416), .A2(n11426), .ZN(n12515) );
  NAND2_X1 U12947 ( .A1(n11766), .A2(n15270), .ZN(n15208) );
  NAND2_X2 U12948 ( .A1(n11687), .A2(n9632), .ZN(n11792) );
  INV_X1 U12949 ( .A(n13620), .ZN(n13617) );
  OR2_X1 U12950 ( .A1(n12368), .A2(n12367), .ZN(n13354) );
  OAI21_X1 U12951 ( .B1(n12851), .B2(n12850), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13003) );
  INV_X1 U12952 ( .A(n15429), .ZN(n11765) );
  AND2_X1 U12953 ( .A1(n11754), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15480) );
  NOR2_X1 U12954 ( .A1(n15227), .A2(n11755), .ZN(n15505) );
  OR3_X1 U12955 ( .A1(n11750), .A2(n15461), .A3(n15769), .ZN(n15760) );
  INV_X1 U12956 ( .A(n16311), .ZN(n15797) );
  AND2_X1 U12957 ( .A1(n13757), .A2(n13756), .ZN(n16374) );
  OR2_X1 U12958 ( .A1(n19302), .A2(n19300), .ZN(n19328) );
  OR2_X1 U12959 ( .A1(n19942), .A2(n19949), .ZN(n19494) );
  OAI21_X2 U12960 ( .B1(n16388), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11986), 
        .ZN(n19781) );
  NOR2_X1 U12961 ( .A1(n18754), .A2(n17483), .ZN(n18943) );
  AOI21_X1 U12962 ( .B1(n16579), .B2(n12148), .A(n12147), .ZN(n12149) );
  NOR2_X1 U12963 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16769), .ZN(n16754) );
  NAND2_X1 U12964 ( .A1(n18943), .A2(n18267), .ZN(n12145) );
  NOR2_X1 U12965 ( .A1(n16797), .A2(n17177), .ZN(n14068) );
  INV_X1 U12966 ( .A(n17410), .ZN(n17290) );
  AOI211_X1 U12967 ( .C1(n12616), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n12571), .B(n12570), .ZN(n12572) );
  INV_X1 U12968 ( .A(n17974), .ZN(n18062) );
  INV_X1 U12969 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17740) );
  NOR2_X1 U12970 ( .A1(n12696), .A2(n17815), .ZN(n12697) );
  NAND2_X1 U12971 ( .A1(n12687), .A2(n10173), .ZN(n12688) );
  AOI222_X1 U12972 ( .A1(n18030), .A2(n16442), .B1(n18024), .B2(n18218), .C1(
        n18751), .C2(n17975), .ZN(n17982) );
  INV_X1 U12973 ( .A(n16442), .ZN(n18035) );
  INV_X1 U12974 ( .A(n17795), .ZN(n17803) );
  NOR2_X1 U12975 ( .A1(n17826), .A2(n10018), .ZN(n17825) );
  NAND2_X1 U12976 ( .A1(n18720), .A2(n12127), .ZN(n15898) );
  AOI211_X1 U12977 ( .C1(n9630), .C2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n12041), .B(n12040), .ZN(n12042) );
  NOR2_X1 U12978 ( .A1(n20835), .A2(n20914), .ZN(n20000) );
  AND2_X1 U12979 ( .A1(n14605), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14565) );
  NOR2_X1 U12980 ( .A1(n14643), .A2(n14496), .ZN(n14620) );
  INV_X1 U12981 ( .A(n20029), .ZN(n20058) );
  AND2_X1 U12982 ( .A1(n13640), .A2(n13639), .ZN(n20089) );
  NOR2_X1 U12983 ( .A1(n14778), .A2(n14540), .ZN(n12837) );
  NAND2_X1 U12984 ( .A1(n11069), .A2(n20000), .ZN(n14849) );
  INV_X1 U12985 ( .A(n13387), .ZN(n20149) );
  OR2_X1 U12986 ( .A1(n13248), .A2(n13247), .ZN(n20159) );
  NAND2_X1 U12987 ( .A1(n10706), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10720) );
  NAND2_X1 U12988 ( .A1(n10613), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10630) );
  NAND2_X1 U12989 ( .A1(n10544), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10560) );
  OAI21_X1 U12990 ( .B1(n20210), .B2(n20208), .A(n16144), .ZN(n20193) );
  OR2_X1 U12991 ( .A1(n13339), .A2(n13338), .ZN(n20214) );
  INV_X1 U12992 ( .A(n15968), .ZN(n15187) );
  INV_X1 U12993 ( .A(n20325), .ZN(n20314) );
  AND2_X1 U12994 ( .A1(n15154), .A2(n20240), .ZN(n20369) );
  AND2_X1 U12995 ( .A1(n20369), .A2(n20621), .ZN(n20420) );
  INV_X1 U12996 ( .A(n20512), .ZN(n20515) );
  INV_X1 U12997 ( .A(n20519), .ZN(n20542) );
  INV_X1 U12998 ( .A(n20609), .ZN(n20597) );
  INV_X1 U12999 ( .A(n20691), .ZN(n20640) );
  AND2_X1 U13000 ( .A1(n9677), .A2(n20241), .ZN(n20621) );
  OAI211_X1 U13001 ( .C1(n20760), .C2(n20730), .A(n20729), .B(n20728), .ZN(
        n20763) );
  INV_X1 U13002 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n10427) );
  INV_X1 U13003 ( .A(n16193), .ZN(n16188) );
  AOI21_X1 U13004 ( .B1(n16194), .B2(n10160), .A(n19851), .ZN(n16201) );
  INV_X1 U13005 ( .A(n19122), .ZN(n19137) );
  INV_X1 U13006 ( .A(n19133), .ZN(n19076) );
  AND2_X1 U13007 ( .A1(n19980), .A2(n16385), .ZN(n19129) );
  INV_X1 U13008 ( .A(n13115), .ZN(n13680) );
  OR2_X1 U13009 ( .A1(n13921), .A2(n13984), .ZN(n13988) );
  OR2_X1 U13010 ( .A1(n12472), .A2(n12471), .ZN(n13819) );
  INV_X1 U13011 ( .A(n14451), .ZN(n14455) );
  NOR2_X1 U13012 ( .A1(n13855), .A2(n13854), .ZN(n19149) );
  INV_X1 U13013 ( .A(n19196), .ZN(n19167) );
  INV_X1 U13014 ( .A(n12982), .ZN(n13017) );
  INV_X1 U13015 ( .A(n18988), .ZN(n15670) );
  INV_X1 U13016 ( .A(n16310), .ZN(n19231) );
  NOR2_X1 U13017 ( .A1(n15494), .A2(n15506), .ZN(n15495) );
  AND2_X1 U13018 ( .A1(n16273), .A2(n16272), .ZN(n16317) );
  AND2_X1 U13019 ( .A1(n12554), .A2(n12511), .ZN(n16324) );
  INV_X1 U13020 ( .A(n15798), .ZN(n15710) );
  OR2_X1 U13021 ( .A1(n16363), .A2(n19645), .ZN(n16388) );
  OAI21_X1 U13022 ( .B1(n19253), .B2(n19252), .A(n19251), .ZN(n19293) );
  AND2_X1 U13023 ( .A1(n19941), .A2(n19462), .ZN(n19330) );
  AND2_X1 U13024 ( .A1(n19934), .A2(n19297), .ZN(n19489) );
  INV_X1 U13025 ( .A(n19400), .ZN(n19388) );
  AND2_X1 U13026 ( .A1(n19489), .A2(n19619), .ZN(n19431) );
  AND2_X1 U13027 ( .A1(n19462), .A2(n10178), .ZN(n19455) );
  AND2_X1 U13028 ( .A1(n19934), .A2(n19961), .ZN(n19462) );
  AOI22_X1 U13029 ( .A1(n19527), .A2(n19526), .B1(n19525), .B2(n19524), .ZN(
        n19545) );
  INV_X1 U13030 ( .A(n19577), .ZN(n19569) );
  AND2_X1 U13031 ( .A1(n19606), .A2(n19941), .ZN(n19602) );
  AND2_X1 U13032 ( .A1(n19942), .A2(n19952), .ZN(n19619) );
  INV_X1 U13033 ( .A(n19787), .ZN(n19682) );
  INV_X1 U13034 ( .A(n19735), .ZN(n19791) );
  XNOR2_X1 U13035 ( .A(n18932), .B(n14066), .ZN(n18945) );
  NOR3_X1 U13036 ( .A1(n15888), .A2(n15886), .A3(n18730), .ZN(n18754) );
  INV_X1 U13037 ( .A(n16884), .ZN(n16924) );
  INV_X1 U13038 ( .A(n16665), .ZN(n16661) );
  NOR2_X1 U13039 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16701), .ZN(n16686) );
  INV_X1 U13040 ( .A(n16901), .ZN(n16933) );
  NOR2_X2 U13041 ( .A1(n18776), .A2(n12145), .ZN(n16884) );
  NOR2_X2 U13042 ( .A1(n18883), .A2(n16929), .ZN(n16922) );
  INV_X1 U13043 ( .A(n17178), .ZN(n17158) );
  INV_X1 U13044 ( .A(n18267), .ZN(n14066) );
  AND2_X1 U13045 ( .A1(n17338), .A2(n17360), .ZN(n17354) );
  AND2_X1 U13046 ( .A1(n12075), .A2(n10165), .ZN(n18286) );
  INV_X1 U13047 ( .A(n17389), .ZN(n17432) );
  NOR2_X1 U13048 ( .A1(n18062), .A2(n17917), .ZN(n17919) );
  NAND2_X1 U13049 ( .A1(n17743), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17720) );
  INV_X1 U13050 ( .A(n17754), .ZN(n17770) );
  NOR2_X1 U13051 ( .A1(n18071), .A2(n17555), .ZN(n16445) );
  NOR2_X1 U13052 ( .A1(n17982), .A2(n18161), .ZN(n17994) );
  INV_X1 U13053 ( .A(n18108), .ZN(n18075) );
  NOR2_X2 U13054 ( .A1(n18240), .A2(n17415), .ZN(n18151) );
  INV_X1 U13055 ( .A(n18230), .ZN(n18246) );
  INV_X1 U13056 ( .A(n18568), .ZN(n18345) );
  AND2_X1 U13057 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18304), .ZN(n18655) );
  INV_X1 U13058 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18799) );
  INV_X1 U13059 ( .A(n13853), .ZN(n13854) );
  OR3_X1 U13060 ( .A1(n14483), .A2(n13227), .A3(n12980), .ZN(n13248) );
  NAND2_X1 U13061 ( .A1(n13248), .A2(n13038), .ZN(n20916) );
  OR2_X1 U13062 ( .A1(n14555), .A2(n14507), .ZN(n14535) );
  NAND2_X1 U13063 ( .A1(n14727), .A2(n13631), .ZN(n20029) );
  INV_X1 U13064 ( .A(n20089), .ZN(n20086) );
  OR2_X1 U13065 ( .A1(n14769), .A2(n20289), .ZN(n14777) );
  INV_X1 U13066 ( .A(n14901), .ZN(n14802) );
  INV_X1 U13067 ( .A(n14945), .ZN(n14826) );
  OR2_X1 U13068 ( .A1(n14849), .A2(n13281), .ZN(n14852) );
  NAND2_X1 U13069 ( .A1(n13229), .A2(n20244), .ZN(n13555) );
  OR3_X1 U13070 ( .A1(n13228), .A2(n14483), .A3(n13227), .ZN(n20127) );
  INV_X1 U13071 ( .A(n20159), .ZN(n13452) );
  OR2_X2 U13072 ( .A1(n15951), .A2(n13227), .ZN(n20007) );
  INV_X1 U13073 ( .A(n20228), .ZN(n20182) );
  NAND2_X1 U13074 ( .A1(n13340), .A2(n13327), .ZN(n20222) );
  INV_X1 U13075 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16175) );
  NAND2_X1 U13076 ( .A1(n20369), .A2(n10149), .ZN(n20325) );
  NAND2_X1 U13077 ( .A1(n20369), .A2(n20551), .ZN(n20364) );
  INV_X1 U13078 ( .A(n20420), .ZN(n20428) );
  NAND2_X1 U13079 ( .A1(n20490), .A2(n10149), .ZN(n20448) );
  NAND2_X1 U13080 ( .A1(n20490), .A2(n20551), .ZN(n20489) );
  NAND2_X1 U13081 ( .A1(n20490), .A2(n20719), .ZN(n20512) );
  NAND2_X1 U13082 ( .A1(n20622), .A2(n10149), .ZN(n20571) );
  NAND2_X1 U13083 ( .A1(n20622), .A2(n20551), .ZN(n20609) );
  NAND2_X1 U13084 ( .A1(n20622), .A2(n20719), .ZN(n20644) );
  NAND2_X1 U13085 ( .A1(n20622), .A2(n20621), .ZN(n20691) );
  NAND2_X1 U13086 ( .A1(n20720), .A2(n10149), .ZN(n20718) );
  NAND2_X1 U13087 ( .A1(n20720), .A2(n20719), .ZN(n20833) );
  INV_X1 U13088 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16181) );
  INV_X1 U13089 ( .A(n20904), .ZN(n20839) );
  INV_X1 U13090 ( .A(n20899), .ZN(n20923) );
  AND2_X1 U13091 ( .A1(n13259), .A2(n13262), .ZN(n19980) );
  AOI21_X1 U13092 ( .B1(n14455), .B2(n19129), .A(n12830), .ZN(n12831) );
  INV_X1 U13093 ( .A(n19129), .ZN(n19127) );
  NAND2_X1 U13094 ( .A1(n12977), .A2(n13262), .ZN(n15269) );
  INV_X1 U13095 ( .A(n15269), .ZN(n15302) );
  XNOR2_X1 U13096 ( .A(n13520), .B(n13521), .ZN(n19942) );
  INV_X1 U13097 ( .A(n19188), .ZN(n15380) );
  OR2_X1 U13098 ( .A1(n19188), .A2(n12266), .ZN(n19183) );
  INV_X1 U13099 ( .A(n19197), .ZN(n19230) );
  INV_X1 U13100 ( .A(n12963), .ZN(n13022) );
  INV_X1 U13101 ( .A(n19236), .ZN(n16303) );
  INV_X1 U13102 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16253) );
  INV_X1 U13103 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16309) );
  INV_X1 U13104 ( .A(n16301), .ZN(n19240) );
  XNOR2_X1 U13105 ( .A(n12259), .B(n10157), .ZN(n15395) );
  INV_X1 U13106 ( .A(n16328), .ZN(n15804) );
  INV_X1 U13107 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15903) );
  AOI21_X1 U13108 ( .B1(n19249), .B2(n19252), .A(n19247), .ZN(n19296) );
  NAND2_X1 U13109 ( .A1(n19941), .A2(n19489), .ZN(n19356) );
  NAND2_X1 U13110 ( .A1(n19462), .A2(n19619), .ZN(n19400) );
  INV_X1 U13111 ( .A(n19431), .ZN(n19428) );
  INV_X1 U13112 ( .A(n19455), .ZN(n19454) );
  INV_X1 U13113 ( .A(n19485), .ZN(n19482) );
  NAND2_X1 U13114 ( .A1(n19931), .A2(n19462), .ZN(n19513) );
  INV_X1 U13115 ( .A(n19544), .ZN(n19540) );
  NAND2_X1 U13116 ( .A1(n19714), .A2(n19941), .ZN(n19577) );
  INV_X1 U13117 ( .A(n19602), .ZN(n19597) );
  NAND2_X1 U13118 ( .A1(n19714), .A2(n19619), .ZN(n19642) );
  NAND2_X1 U13119 ( .A1(n19714), .A2(n10178), .ZN(n19703) );
  INV_X1 U13120 ( .A(n19745), .ZN(n19767) );
  INV_X1 U13121 ( .A(n19838), .ZN(n19823) );
  INV_X1 U13122 ( .A(n16395), .ZN(n19848) );
  INV_X1 U13123 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16800) );
  INV_X1 U13124 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17862) );
  INV_X1 U13125 ( .A(n16893), .ZN(n18948) );
  AND2_X1 U13126 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17068), .ZN(n17082) );
  AND2_X1 U13127 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17222), .ZN(n17249) );
  NOR2_X1 U13128 ( .A1(n17438), .A2(n17291), .ZN(n17389) );
  INV_X1 U13129 ( .A(n12663), .ZN(n17426) );
  INV_X1 U13130 ( .A(n17409), .ZN(n17444) );
  INV_X1 U13131 ( .A(n17464), .ZN(n17482) );
  AND2_X1 U13132 ( .A1(n12760), .A2(n12759), .ZN(n12761) );
  INV_X1 U13133 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18134) );
  INV_X1 U13134 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17880) );
  NOR2_X1 U13135 ( .A1(n17818), .A2(n17820), .ZN(n17909) );
  INV_X1 U13136 ( .A(n18151), .ZN(n18170) );
  INV_X1 U13137 ( .A(n18242), .ZN(n18233) );
  INV_X1 U13138 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18539) );
  INV_X1 U13139 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18516) );
  INV_X1 U13140 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18601) );
  CLKBUF_X1 U13141 ( .A(n18792), .Z(n18879) );
  OAI21_X1 U13142 ( .B1(n14863), .B2(n14779), .A(n11196), .ZN(P1_U2842) );
  OAI21_X1 U13143 ( .B1(n14789), .B2(n14779), .A(n12838), .ZN(P1_U2844) );
  AND2_X2 U13144 ( .A1(n13425), .A2(n10190), .ZN(n10364) );
  AOI22_X1 U13145 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10364), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10188) );
  AOI22_X1 U13146 ( .A1(n10343), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10363), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U13147 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10186) );
  AND2_X2 U13148 ( .A1(n10190), .A2(n13431), .ZN(n10250) );
  AOI22_X1 U13149 ( .A1(n10370), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10250), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U13150 ( .A1(n10979), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10978), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10197) );
  AOI22_X1 U13151 ( .A1(n13424), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U13152 ( .A1(n10369), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10836), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10195) );
  AOI22_X1 U13153 ( .A1(n10348), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10349), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10194) );
  AOI22_X1 U13154 ( .A1(n10363), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10978), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10201) );
  AOI22_X1 U13155 ( .A1(n10364), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13424), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10200) );
  AOI22_X1 U13156 ( .A1(n10369), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10250), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10199) );
  AOI22_X1 U13157 ( .A1(n10348), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10349), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10198) );
  AOI22_X1 U13158 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10205) );
  AOI22_X1 U13159 ( .A1(n10343), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10204) );
  AOI22_X1 U13160 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U13161 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10836), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10202) );
  INV_X2 U13162 ( .A(n10300), .ZN(n20271) );
  AOI22_X1 U13163 ( .A1(n10250), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9650), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10210) );
  AOI22_X1 U13164 ( .A1(n13424), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10369), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10209) );
  AOI22_X1 U13165 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10349), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10208) );
  AOI22_X1 U13166 ( .A1(n10348), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10207) );
  AOI22_X1 U13167 ( .A1(n10364), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9667), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10214) );
  AOI22_X1 U13168 ( .A1(n10343), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9669), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10213) );
  AOI22_X1 U13169 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10211) );
  NAND2_X1 U13170 ( .A1(n10364), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10218) );
  NAND2_X1 U13171 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10217) );
  NAND2_X1 U13172 ( .A1(n10289), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10216) );
  NAND2_X1 U13173 ( .A1(n10978), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10215) );
  NAND2_X1 U13174 ( .A1(n10348), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10222) );
  NAND2_X1 U13175 ( .A1(n10370), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10221) );
  NAND2_X1 U13176 ( .A1(n10979), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10220) );
  NAND2_X1 U13177 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10219) );
  NAND2_X1 U13178 ( .A1(n13424), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10226) );
  NAND2_X1 U13179 ( .A1(n10369), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10225) );
  NAND2_X1 U13180 ( .A1(n10250), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10224) );
  NAND2_X1 U13181 ( .A1(n10836), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10223) );
  NAND2_X1 U13182 ( .A1(n10343), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10230) );
  NAND2_X1 U13183 ( .A1(n10363), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10229) );
  NAND2_X1 U13184 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10228) );
  NAND2_X1 U13185 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10227) );
  AND2_X2 U13186 ( .A1(n10318), .A2(n14160), .ZN(n13163) );
  AOI22_X1 U13187 ( .A1(n13424), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10369), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10239) );
  AOI22_X1 U13188 ( .A1(n10348), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10238) );
  AOI22_X1 U13189 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10349), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10237) );
  AOI22_X1 U13190 ( .A1(n10250), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9650), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10236) );
  NAND4_X1 U13191 ( .A1(n10239), .A2(n10238), .A3(n10237), .A4(n10236), .ZN(
        n10245) );
  AOI22_X1 U13192 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10289), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10243) );
  AOI22_X1 U13193 ( .A1(n10343), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10363), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10242) );
  AOI22_X1 U13194 ( .A1(n10364), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9667), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10241) );
  AOI22_X1 U13195 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10240) );
  NAND4_X1 U13196 ( .A1(n10243), .A2(n10242), .A3(n10241), .A4(n10240), .ZN(
        n10244) );
  NAND2_X1 U13197 ( .A1(n14160), .A2(n20280), .ZN(n10256) );
  AOI22_X1 U13198 ( .A1(n10364), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10363), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10249) );
  AOI22_X1 U13199 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13424), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10248) );
  AOI22_X1 U13200 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10247) );
  AOI22_X1 U13201 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10246) );
  AOI22_X1 U13202 ( .A1(n10369), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10250), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10254) );
  AOI22_X1 U13203 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10348), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10253) );
  AOI22_X1 U13204 ( .A1(n10343), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10978), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10252) );
  AOI22_X1 U13205 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10349), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10251) );
  NAND2_X1 U13206 ( .A1(n10364), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10263) );
  NAND2_X1 U13207 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10262) );
  NAND2_X1 U13208 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10261) );
  NAND2_X1 U13209 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10260) );
  NAND2_X1 U13210 ( .A1(n10348), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10267) );
  NAND2_X1 U13211 ( .A1(n10370), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10266) );
  NAND2_X1 U13212 ( .A1(n10979), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10265) );
  NAND2_X1 U13213 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10264) );
  NAND2_X1 U13214 ( .A1(n13424), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10271) );
  NAND2_X1 U13215 ( .A1(n10369), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10270) );
  NAND2_X1 U13216 ( .A1(n10250), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10269) );
  NAND2_X1 U13217 ( .A1(n10836), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10268) );
  NAND2_X1 U13218 ( .A1(n10343), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10275) );
  NAND2_X1 U13219 ( .A1(n10363), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10274) );
  NAND2_X1 U13220 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10273) );
  NAND2_X1 U13221 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10272) );
  NAND2_X1 U13222 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10284) );
  NAND2_X1 U13223 ( .A1(n10348), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10283) );
  NAND2_X1 U13224 ( .A1(n13424), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10282) );
  NAND2_X1 U13225 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10281) );
  NAND2_X1 U13226 ( .A1(n10836), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10288) );
  NAND2_X1 U13227 ( .A1(n10364), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10287) );
  NAND2_X1 U13228 ( .A1(n10363), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10286) );
  NAND2_X1 U13229 ( .A1(n10369), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10285) );
  NAND2_X1 U13230 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10292) );
  NAND2_X1 U13231 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10291) );
  NAND2_X1 U13232 ( .A1(n10250), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10290) );
  NAND4_X4 U13233 ( .A1(n10296), .A2(n10295), .A3(n10294), .A4(n9703), .ZN(
        n20258) );
  INV_X1 U13234 ( .A(n13169), .ZN(n10299) );
  NAND2_X1 U13235 ( .A1(n10299), .A2(n10298), .ZN(n10303) );
  NAND2_X1 U13236 ( .A1(n13163), .A2(n13329), .ZN(n10302) );
  NAND2_X1 U13237 ( .A1(n10304), .A2(n20280), .ZN(n10301) );
  AND2_X2 U13238 ( .A1(n10301), .A2(n20289), .ZN(n10305) );
  XNOR2_X1 U13239 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n13183) );
  INV_X1 U13240 ( .A(n13163), .ZN(n13280) );
  INV_X1 U13241 ( .A(n10305), .ZN(n10317) );
  NAND3_X1 U13242 ( .A1(n13280), .A2(n13329), .A3(n10305), .ZN(n13164) );
  AOI21_X1 U13243 ( .B1(n13164), .B2(n10306), .A(n13165), .ZN(n10310) );
  NAND2_X1 U13244 ( .A1(n10307), .A2(n13632), .ZN(n10309) );
  MUX2_X1 U13245 ( .A(n13315), .B(n13310), .S(n13632), .Z(n10308) );
  NAND2_X1 U13246 ( .A1(n10332), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10313) );
  NAND2_X1 U13247 ( .A1(n16172), .A2(n20914), .ZN(n12250) );
  NAND2_X1 U13248 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10334) );
  OAI21_X1 U13249 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n10334), .ZN(n20575) );
  NAND2_X1 U13250 ( .A1(n20835), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10329) );
  OAI21_X1 U13251 ( .B1(n12250), .B2(n20575), .A(n10329), .ZN(n10311) );
  INV_X1 U13252 ( .A(n10311), .ZN(n10312) );
  NAND2_X1 U13253 ( .A1(n10313), .A2(n10312), .ZN(n10314) );
  INV_X1 U13254 ( .A(n20835), .ZN(n15965) );
  MUX2_X1 U13255 ( .A(n15965), .B(n12250), .S(n20692), .Z(n10315) );
  NAND3_X1 U13256 ( .A1(n13164), .A2(n10306), .A3(n20258), .ZN(n10321) );
  INV_X1 U13257 ( .A(n16172), .ZN(n15184) );
  NOR2_X1 U13258 ( .A1(n15184), .A2(n20914), .ZN(n10320) );
  NAND2_X1 U13259 ( .A1(n20910), .A2(n10317), .ZN(n10319) );
  NAND2_X1 U13260 ( .A1(n13165), .A2(n10318), .ZN(n13334) );
  NAND4_X1 U13261 ( .A1(n10321), .A2(n10320), .A3(n10319), .A4(n13334), .ZN(
        n10324) );
  INV_X1 U13262 ( .A(n10322), .ZN(n10323) );
  NOR2_X1 U13263 ( .A1(n10324), .A2(n10323), .ZN(n10327) );
  INV_X1 U13264 ( .A(n14484), .ZN(n14482) );
  NAND3_X1 U13265 ( .A1(n14482), .A2(n13280), .A3(n20267), .ZN(n10325) );
  NAND2_X1 U13266 ( .A1(n10307), .A2(n10325), .ZN(n10326) );
  NAND2_X1 U13267 ( .A1(n10327), .A2(n10326), .ZN(n10360) );
  INV_X1 U13268 ( .A(n10328), .ZN(n10331) );
  NAND2_X1 U13269 ( .A1(n10329), .A2(n10183), .ZN(n10330) );
  NAND2_X1 U13270 ( .A1(n10331), .A2(n10330), .ZN(n10340) );
  NAND2_X1 U13271 ( .A1(n10416), .A2(n10340), .ZN(n10338) );
  NAND2_X1 U13272 ( .A1(n10332), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10337) );
  INV_X1 U13273 ( .A(n10334), .ZN(n10333) );
  NAND2_X1 U13274 ( .A1(n10333), .A2(n20646), .ZN(n20610) );
  NAND2_X1 U13275 ( .A1(n10334), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10335) );
  NAND2_X1 U13276 ( .A1(n20610), .A2(n10335), .ZN(n20252) );
  INV_X1 U13277 ( .A(n12250), .ZN(n10456) );
  AOI22_X1 U13278 ( .A1(n20252), .A2(n10456), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n20835), .ZN(n10336) );
  INV_X1 U13279 ( .A(n10339), .ZN(n10341) );
  NAND3_X1 U13280 ( .A1(n10416), .A2(n10341), .A3(n10340), .ZN(n10342) );
  AOI22_X1 U13281 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10347) );
  AOI22_X1 U13282 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U13283 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10345) );
  AOI22_X1 U13284 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10344) );
  NAND4_X1 U13285 ( .A1(n10347), .A2(n10346), .A3(n10345), .A4(n10344), .ZN(
        n10355) );
  INV_X1 U13286 ( .A(n13424), .ZN(n10382) );
  INV_X2 U13287 ( .A(n10382), .ZN(n10956) );
  AOI22_X1 U13288 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10353) );
  AOI22_X1 U13289 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10352) );
  AOI22_X1 U13290 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10351) );
  AOI22_X1 U13291 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9650), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10350) );
  NAND4_X1 U13292 ( .A1(n10353), .A2(n10352), .A3(n10351), .A4(n10350), .ZN(
        n10354) );
  INV_X1 U13293 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10357) );
  OAI22_X1 U13294 ( .A1(n11042), .A2(n10357), .B1(n12173), .B2(n10459), .ZN(
        n10358) );
  INV_X1 U13295 ( .A(n10360), .ZN(n10361) );
  AOI22_X1 U13296 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n9674), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10368) );
  AOI22_X1 U13297 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10363), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10367) );
  AOI22_X1 U13298 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n10938), .B1(
        n10978), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U13299 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10365) );
  NAND4_X1 U13300 ( .A1(n10368), .A2(n10367), .A3(n10366), .A4(n10365), .ZN(
        n10376) );
  AOI22_X1 U13301 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n13424), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10374) );
  AOI22_X1 U13302 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10986), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10373) );
  AOI22_X1 U13303 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10372) );
  AOI22_X1 U13304 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10980), .B1(
        n10836), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10371) );
  NAND4_X1 U13305 ( .A1(n10374), .A2(n10373), .A3(n10372), .A4(n10371), .ZN(
        n10375) );
  INV_X1 U13306 ( .A(n12219), .ZN(n10377) );
  NAND2_X1 U13307 ( .A1(n10377), .A2(n13329), .ZN(n10389) );
  AOI22_X1 U13308 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U13309 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U13310 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U13311 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10378) );
  NAND4_X1 U13312 ( .A1(n10381), .A2(n10380), .A3(n10379), .A4(n10378), .ZN(
        n10388) );
  AOI22_X1 U13313 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9676), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U13314 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10385) );
  AOI22_X1 U13315 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10978), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10384) );
  AOI22_X1 U13316 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9650), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10383) );
  NAND4_X1 U13317 ( .A1(n10386), .A2(n10385), .A3(n10384), .A4(n10383), .ZN(
        n10387) );
  MUX2_X1 U13318 ( .A(n12215), .B(n10389), .S(n12157), .Z(n10390) );
  INV_X1 U13319 ( .A(n10390), .ZN(n10391) );
  NAND2_X1 U13320 ( .A1(n10391), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10442) );
  INV_X1 U13321 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10392) );
  AOI21_X1 U13322 ( .B1(n13632), .B2(n12157), .A(n20914), .ZN(n10393) );
  INV_X1 U13323 ( .A(n12215), .ZN(n10396) );
  NAND2_X1 U13324 ( .A1(n10396), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U13325 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10402) );
  AOI22_X1 U13326 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10401) );
  AOI22_X1 U13327 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10400) );
  AOI22_X1 U13328 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10250), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10399) );
  NAND4_X1 U13329 ( .A1(n10402), .A2(n10401), .A3(n10400), .A4(n10399), .ZN(
        n10408) );
  AOI22_X1 U13330 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10986), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10406) );
  AOI22_X1 U13331 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10405) );
  AOI22_X1 U13332 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10836), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10404) );
  AOI22_X1 U13333 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10403) );
  NAND4_X1 U13334 ( .A1(n10406), .A2(n10405), .A3(n10404), .A4(n10403), .ZN(
        n10407) );
  INV_X1 U13335 ( .A(n12158), .ZN(n10417) );
  OAI22_X1 U13336 ( .A1(n10460), .A2(n12219), .B1(n10459), .B2(n10417), .ZN(
        n10409) );
  INV_X1 U13337 ( .A(n10409), .ZN(n10412) );
  INV_X1 U13338 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10410) );
  INV_X1 U13339 ( .A(n20366), .ZN(n10415) );
  INV_X1 U13340 ( .A(n10413), .ZN(n10414) );
  NAND2_X1 U13341 ( .A1(n10434), .A2(n12156), .ZN(n10423) );
  INV_X1 U13342 ( .A(n10419), .ZN(n10420) );
  NAND2_X1 U13343 ( .A1(n13328), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10483) );
  NOR2_X1 U13344 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n10426) );
  XNOR2_X1 U13345 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14729) );
  AOI21_X1 U13346 ( .B1(n13628), .B2(n14729), .A(n11005), .ZN(n10430) );
  NOR2_X2 U13347 ( .A1(n20289), .A2(n10427), .ZN(n10428) );
  NAND2_X1 U13348 ( .A1(n11006), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n10429) );
  OAI211_X1 U13349 ( .C1(n10483), .C2(n10184), .A(n10430), .B(n10429), .ZN(
        n10431) );
  INV_X1 U13350 ( .A(n10431), .ZN(n10432) );
  NAND2_X1 U13351 ( .A1(n11005), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10453) );
  NAND2_X1 U13352 ( .A1(n10433), .A2(n10453), .ZN(n13297) );
  INV_X1 U13353 ( .A(n13297), .ZN(n10452) );
  NAND2_X1 U13354 ( .A1(n13474), .A2(n10684), .ZN(n10440) );
  AOI22_X1 U13355 ( .A1(n11006), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20837), .ZN(n10438) );
  INV_X1 U13356 ( .A(n10483), .ZN(n10499) );
  NAND2_X1 U13357 ( .A1(n10499), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10437) );
  AND2_X1 U13358 ( .A1(n10438), .A2(n10437), .ZN(n10439) );
  NAND2_X1 U13359 ( .A1(n10440), .A2(n10439), .ZN(n13254) );
  NAND2_X1 U13360 ( .A1(n20326), .A2(n10318), .ZN(n10444) );
  NAND2_X1 U13361 ( .A1(n10444), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13057) );
  NAND2_X1 U13362 ( .A1(n20837), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10447) );
  NAND2_X1 U13363 ( .A1(n11006), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n10446) );
  OAI211_X1 U13364 ( .C1(n10483), .C2(n13182), .A(n10447), .B(n10446), .ZN(
        n10448) );
  AOI21_X1 U13365 ( .B1(n10445), .B2(n10684), .A(n10448), .ZN(n10449) );
  OR2_X1 U13366 ( .A1(n13057), .A2(n10449), .ZN(n13058) );
  INV_X1 U13367 ( .A(n10449), .ZN(n13059) );
  OR2_X1 U13368 ( .A1(n13059), .A2(n11004), .ZN(n10450) );
  NAND2_X1 U13369 ( .A1(n13058), .A2(n10450), .ZN(n13253) );
  NAND2_X1 U13370 ( .A1(n10452), .A2(n10451), .ZN(n13294) );
  NAND2_X1 U13371 ( .A1(n13294), .A2(n10453), .ZN(n13372) );
  NAND2_X1 U13372 ( .A1(n10332), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10458) );
  NAND2_X1 U13373 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10147), .ZN(
        n20492) );
  NAND2_X1 U13374 ( .A1(n20645), .A2(n20492), .ZN(n10455) );
  NOR3_X1 U13375 ( .A1(n20645), .A2(n20646), .A3(n20572), .ZN(n20782) );
  NAND2_X1 U13376 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20782), .ZN(
        n20769) );
  AND2_X1 U13377 ( .A1(n10455), .A2(n20769), .ZN(n20520) );
  AOI22_X1 U13378 ( .A1(n10456), .A2(n20520), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20835), .ZN(n10457) );
  XNOR2_X2 U13379 ( .A(n10454), .B(n20401), .ZN(n13423) );
  AOI22_X1 U13380 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10464) );
  AOI22_X1 U13381 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9676), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10463) );
  AOI22_X1 U13382 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10462) );
  AOI22_X1 U13383 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10836), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10461) );
  NAND4_X1 U13384 ( .A1(n10464), .A2(n10463), .A3(n10462), .A4(n10461), .ZN(
        n10470) );
  AOI22_X1 U13385 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10468) );
  AOI22_X1 U13386 ( .A1(n10987), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10467) );
  AOI22_X1 U13387 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10466) );
  AOI22_X1 U13388 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10465) );
  NAND4_X1 U13389 ( .A1(n10468), .A2(n10467), .A3(n10466), .A4(n10465), .ZN(
        n10469) );
  AOI22_X1 U13390 ( .A1(n11046), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11024), .B2(n12180), .ZN(n10471) );
  INV_X1 U13391 ( .A(n10474), .ZN(n15156) );
  NAND2_X1 U13392 ( .A1(n10475), .A2(n15156), .ZN(n10476) );
  INV_X1 U13393 ( .A(n10478), .ZN(n10480) );
  INV_X1 U13394 ( .A(n10502), .ZN(n10479) );
  OAI21_X1 U13395 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n10480), .A(
        n10479), .ZN(n20090) );
  AOI22_X1 U13396 ( .A1(n13628), .A2(n20090), .B1(n11005), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10482) );
  NAND2_X1 U13397 ( .A1(n11006), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n10481) );
  OAI211_X1 U13398 ( .C1(n10483), .C2(n9920), .A(n10482), .B(n10481), .ZN(
        n10484) );
  INV_X1 U13399 ( .A(n10484), .ZN(n10485) );
  OAI21_X1 U13400 ( .B1(n15154), .B2(n10610), .A(n10485), .ZN(n13373) );
  INV_X1 U13401 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13402 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13403 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U13404 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13405 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10487) );
  NAND4_X1 U13406 ( .A1(n10490), .A2(n10489), .A3(n10488), .A4(n10487), .ZN(
        n10496) );
  AOI22_X1 U13407 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10494) );
  AOI22_X1 U13408 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10493) );
  AOI22_X1 U13409 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13410 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10836), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10491) );
  NAND4_X1 U13411 ( .A1(n10494), .A2(n10493), .A3(n10492), .A4(n10491), .ZN(
        n10495) );
  NAND2_X1 U13412 ( .A1(n11024), .A2(n12188), .ZN(n10497) );
  XNOR2_X1 U13413 ( .A(n10507), .B(n10508), .ZN(n12179) );
  NAND2_X1 U13414 ( .A1(n10499), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10505) );
  INV_X1 U13415 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10500) );
  AOI21_X1 U13416 ( .B1(n10500), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10501) );
  AOI21_X1 U13417 ( .B1(n11006), .B2(P1_EAX_REG_4__SCAN_IN), .A(n10501), .ZN(
        n10504) );
  OAI21_X1 U13418 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n10502), .A(
        n10522), .ZN(n20177) );
  NOR2_X1 U13419 ( .A1(n20177), .A2(n11004), .ZN(n10503) );
  AOI21_X1 U13420 ( .B1(n10505), .B2(n10504), .A(n10503), .ZN(n10506) );
  INV_X1 U13421 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U13422 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9674), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U13423 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9676), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10512) );
  AOI22_X1 U13424 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10511) );
  AOI22_X1 U13425 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10250), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10510) );
  NAND4_X1 U13426 ( .A1(n10513), .A2(n10512), .A3(n10511), .A4(n10510), .ZN(
        n10519) );
  AOI22_X1 U13427 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10517) );
  AOI22_X1 U13428 ( .A1(n10987), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10516) );
  AOI22_X1 U13429 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U13430 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10514) );
  NAND4_X1 U13431 ( .A1(n10517), .A2(n10516), .A3(n10515), .A4(n10514), .ZN(
        n10518) );
  NAND2_X1 U13432 ( .A1(n11024), .A2(n12198), .ZN(n10520) );
  XNOR2_X1 U13433 ( .A(n10551), .B(n10552), .ZN(n12187) );
  NAND2_X1 U13434 ( .A1(n12187), .A2(n10684), .ZN(n10528) );
  INV_X1 U13435 ( .A(n11005), .ZN(n10689) );
  INV_X1 U13436 ( .A(n10522), .ZN(n10524) );
  INV_X1 U13437 ( .A(n10544), .ZN(n10523) );
  OAI21_X1 U13438 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n10524), .A(
        n10523), .ZN(n20074) );
  NAND2_X1 U13439 ( .A1(n20074), .A2(n13628), .ZN(n10525) );
  OAI21_X1 U13440 ( .B1(n20066), .B2(n10689), .A(n10525), .ZN(n10526) );
  AOI21_X1 U13441 ( .B1(n10428), .B2(P1_EAX_REG_5__SCAN_IN), .A(n10526), .ZN(
        n10527) );
  NAND2_X1 U13442 ( .A1(n10528), .A2(n10527), .ZN(n13365) );
  NAND2_X1 U13443 ( .A1(n10529), .A2(n10552), .ZN(n10543) );
  INV_X1 U13444 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10530) );
  AOI22_X1 U13445 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10534) );
  AOI22_X1 U13446 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10533) );
  AOI22_X1 U13447 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U13448 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10531) );
  NAND4_X1 U13449 ( .A1(n10534), .A2(n10533), .A3(n10532), .A4(n10531), .ZN(
        n10540) );
  AOI22_X1 U13450 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10538) );
  AOI22_X1 U13451 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13452 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13453 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10535) );
  NAND4_X1 U13454 ( .A1(n10538), .A2(n10537), .A3(n10536), .A4(n10535), .ZN(
        n10539) );
  NAND2_X1 U13455 ( .A1(n11024), .A2(n12207), .ZN(n10541) );
  INV_X1 U13456 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n10546) );
  OAI21_X1 U13457 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n10544), .A(
        n10560), .ZN(n20062) );
  AOI22_X1 U13458 ( .A1(n13628), .A2(n20062), .B1(n11005), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10545) );
  OAI21_X1 U13459 ( .B1(n10905), .B2(n10546), .A(n10545), .ZN(n10547) );
  NAND2_X1 U13460 ( .A1(n10550), .A2(n13531), .ZN(n13530) );
  INV_X1 U13461 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10558) );
  NAND2_X1 U13462 ( .A1(n11024), .A2(n12219), .ZN(n10557) );
  OAI21_X1 U13463 ( .B1(n11042), .B2(n10558), .A(n10557), .ZN(n10559) );
  INV_X1 U13464 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n10564) );
  INV_X1 U13465 ( .A(n10560), .ZN(n10562) );
  INV_X1 U13466 ( .A(n10581), .ZN(n10561) );
  OAI21_X1 U13467 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n10562), .A(
        n10561), .ZN(n20049) );
  AOI22_X1 U13468 ( .A1(n13628), .A2(n20049), .B1(n11005), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10563) );
  OAI21_X1 U13469 ( .B1(n10905), .B2(n10564), .A(n10563), .ZN(n10565) );
  INV_X1 U13470 ( .A(n13653), .ZN(n10566) );
  AOI22_X1 U13471 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10570) );
  AOI22_X1 U13472 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U13473 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U13474 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10250), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10567) );
  NAND4_X1 U13475 ( .A1(n10570), .A2(n10569), .A3(n10568), .A4(n10567), .ZN(
        n10576) );
  AOI22_X1 U13476 ( .A1(n10987), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10574) );
  AOI22_X1 U13477 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10573) );
  AOI22_X1 U13478 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13479 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10571) );
  NAND4_X1 U13480 ( .A1(n10574), .A2(n10573), .A3(n10572), .A4(n10571), .ZN(
        n10575) );
  OAI21_X1 U13481 ( .B1(n10576), .B2(n10575), .A(n10684), .ZN(n10579) );
  NAND2_X1 U13482 ( .A1(n11006), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n10578) );
  XNOR2_X1 U13483 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n10581), .ZN(
        n13801) );
  AOI22_X1 U13484 ( .A1(n13628), .A2(n13801), .B1(n11005), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10577) );
  XOR2_X1 U13485 ( .A(n10606), .B(n10607), .Z(n13870) );
  AOI22_X1 U13486 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10585) );
  AOI22_X1 U13487 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10584) );
  AOI22_X1 U13488 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10583) );
  AOI22_X1 U13489 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10582) );
  NAND4_X1 U13490 ( .A1(n10585), .A2(n10584), .A3(n10583), .A4(n10582), .ZN(
        n10591) );
  AOI22_X1 U13491 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U13492 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10588) );
  AOI22_X1 U13493 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10587) );
  AOI22_X1 U13494 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10586) );
  NAND4_X1 U13495 ( .A1(n10589), .A2(n10588), .A3(n10587), .A4(n10586), .ZN(
        n10590) );
  OAI21_X1 U13496 ( .B1(n10591), .B2(n10590), .A(n10684), .ZN(n10594) );
  NAND2_X1 U13497 ( .A1(n11006), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n10593) );
  NAND2_X1 U13498 ( .A1(n11005), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10592) );
  NAND3_X1 U13499 ( .A1(n10594), .A2(n10593), .A3(n10592), .ZN(n10595) );
  AOI22_X1 U13500 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10599) );
  AOI22_X1 U13501 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9676), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10598) );
  AOI22_X1 U13502 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10250), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10597) );
  AOI22_X1 U13503 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10596) );
  NAND4_X1 U13504 ( .A1(n10599), .A2(n10598), .A3(n10597), .A4(n10596), .ZN(
        n10605) );
  AOI22_X1 U13505 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U13506 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10602) );
  AOI22_X1 U13507 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10601) );
  AOI22_X1 U13508 ( .A1(n10979), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10600) );
  NAND4_X1 U13509 ( .A1(n10603), .A2(n10602), .A3(n10601), .A4(n10600), .ZN(
        n10604) );
  NOR2_X1 U13510 ( .A1(n10605), .A2(n10604), .ZN(n10611) );
  XNOR2_X1 U13511 ( .A(n10612), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14718) );
  NAND2_X1 U13512 ( .A1(n14718), .A2(n13628), .ZN(n10609) );
  AOI22_X1 U13513 ( .A1(n11006), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n11005), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10608) );
  OAI211_X1 U13514 ( .C1(n10611), .C2(n10610), .A(n10609), .B(n10608), .ZN(
        n13825) );
  INV_X1 U13515 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10615) );
  OAI21_X1 U13516 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n10613), .A(
        n10630), .ZN(n16061) );
  NAND2_X1 U13517 ( .A1(n16061), .A2(n13628), .ZN(n10614) );
  OAI21_X1 U13518 ( .B1(n10615), .B2(n10689), .A(n10614), .ZN(n10616) );
  AOI21_X1 U13519 ( .B1(n10428), .B2(P1_EAX_REG_11__SCAN_IN), .A(n10616), .ZN(
        n10617) );
  AOI22_X1 U13520 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10621) );
  AOI22_X1 U13521 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U13522 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13523 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10618) );
  NAND4_X1 U13524 ( .A1(n10621), .A2(n10620), .A3(n10619), .A4(n10618), .ZN(
        n10627) );
  AOI22_X1 U13525 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10956), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10625) );
  AOI22_X1 U13526 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10624) );
  AOI22_X1 U13527 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10623) );
  AOI22_X1 U13528 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10622) );
  NAND4_X1 U13529 ( .A1(n10625), .A2(n10624), .A3(n10623), .A4(n10622), .ZN(
        n10626) );
  OR2_X1 U13530 ( .A1(n10627), .A2(n10626), .ZN(n10628) );
  AND2_X1 U13531 ( .A1(n10684), .A2(n10628), .ZN(n13967) );
  XOR2_X1 U13532 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n10645), .Z(
        n16015) );
  AOI22_X1 U13533 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10634) );
  AOI22_X1 U13534 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10633) );
  AOI22_X1 U13535 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10632) );
  AOI22_X1 U13536 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10631) );
  NAND4_X1 U13537 ( .A1(n10634), .A2(n10633), .A3(n10632), .A4(n10631), .ZN(
        n10640) );
  AOI22_X1 U13538 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10956), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10638) );
  AOI22_X1 U13539 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10637) );
  AOI22_X1 U13540 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10636) );
  AOI22_X1 U13541 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10635) );
  NAND4_X1 U13542 ( .A1(n10638), .A2(n10637), .A3(n10636), .A4(n10635), .ZN(
        n10639) );
  OAI21_X1 U13543 ( .B1(n10640), .B2(n10639), .A(n10684), .ZN(n10643) );
  NAND2_X1 U13544 ( .A1(n11006), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n10642) );
  NAND2_X1 U13545 ( .A1(n11005), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10641) );
  AND3_X1 U13546 ( .A1(n10643), .A2(n10642), .A3(n10641), .ZN(n10644) );
  OAI21_X1 U13547 ( .B1(n16015), .B2(n11004), .A(n10644), .ZN(n14003) );
  XNOR2_X1 U13548 ( .A(n10660), .B(n10659), .ZN(n14997) );
  AOI22_X1 U13549 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10956), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10649) );
  AOI22_X1 U13550 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10648) );
  AOI22_X1 U13551 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10647) );
  AOI22_X1 U13552 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10646) );
  NAND4_X1 U13553 ( .A1(n10649), .A2(n10648), .A3(n10647), .A4(n10646), .ZN(
        n10655) );
  AOI22_X1 U13554 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U13555 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U13556 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10651) );
  AOI22_X1 U13557 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10650) );
  NAND4_X1 U13558 ( .A1(n10653), .A2(n10652), .A3(n10651), .A4(n10650), .ZN(
        n10654) );
  OAI21_X1 U13559 ( .B1(n10655), .B2(n10654), .A(n10684), .ZN(n10657) );
  NAND2_X1 U13560 ( .A1(n10428), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n10656) );
  OAI211_X1 U13561 ( .C1(n10689), .C2(n10659), .A(n10657), .B(n10656), .ZN(
        n10658) );
  AOI21_X1 U13562 ( .B1(n14997), .B2(n10426), .A(n10658), .ZN(n14702) );
  INV_X1 U13563 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16005) );
  XNOR2_X1 U13564 ( .A(n16005), .B(n10675), .ZN(n16043) );
  AOI22_X1 U13565 ( .A1(n10987), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10664) );
  AOI22_X1 U13566 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10663) );
  AOI22_X1 U13567 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10662) );
  AOI22_X1 U13568 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10661) );
  NAND4_X1 U13569 ( .A1(n10664), .A2(n10663), .A3(n10662), .A4(n10661), .ZN(
        n10670) );
  AOI22_X1 U13570 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U13571 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9676), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U13572 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10666) );
  AOI22_X1 U13573 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10665) );
  NAND4_X1 U13574 ( .A1(n10668), .A2(n10667), .A3(n10666), .A4(n10665), .ZN(
        n10669) );
  OAI21_X1 U13575 ( .B1(n10670), .B2(n10669), .A(n10684), .ZN(n10673) );
  NAND2_X1 U13576 ( .A1(n10428), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n10672) );
  NAND2_X1 U13577 ( .A1(n11005), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10671) );
  AND3_X1 U13578 ( .A1(n10673), .A2(n10672), .A3(n10671), .ZN(n10674) );
  OAI21_X1 U13579 ( .B1(n16043), .B2(n11004), .A(n10674), .ZN(n14771) );
  XNOR2_X1 U13580 ( .A(n10705), .B(n14696), .ZN(n14988) );
  AOI22_X1 U13581 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10987), .B1(
        n10956), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U13582 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n10938), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10678) );
  AOI22_X1 U13583 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10677) );
  AOI22_X1 U13584 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10676) );
  NAND4_X1 U13585 ( .A1(n10679), .A2(n10678), .A3(n10677), .A4(n10676), .ZN(
        n10686) );
  AOI22_X1 U13586 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10986), .B1(
        n9674), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U13587 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U13588 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U13589 ( .A1(n9668), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n9666), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10680) );
  NAND4_X1 U13590 ( .A1(n10683), .A2(n10682), .A3(n10681), .A4(n10680), .ZN(
        n10685) );
  OAI21_X1 U13591 ( .B1(n10686), .B2(n10685), .A(n10684), .ZN(n10688) );
  NAND2_X1 U13592 ( .A1(n11006), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n10687) );
  OAI211_X1 U13593 ( .C1(n10689), .C2(n14696), .A(n10688), .B(n10687), .ZN(
        n10690) );
  AOI21_X1 U13594 ( .B1(n14988), .B2(n10426), .A(n10690), .ZN(n14690) );
  AOI22_X1 U13595 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9674), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10694) );
  AOI22_X1 U13596 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U13597 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U13598 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10691) );
  NAND4_X1 U13599 ( .A1(n10694), .A2(n10693), .A3(n10692), .A4(n10691), .ZN(
        n10700) );
  AOI22_X1 U13600 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10956), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U13601 ( .A1(n10987), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10697) );
  AOI22_X1 U13602 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10696) );
  AOI22_X1 U13603 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10695) );
  NAND4_X1 U13604 ( .A1(n10698), .A2(n10697), .A3(n10696), .A4(n10695), .ZN(
        n10699) );
  NOR2_X1 U13605 ( .A1(n10700), .A2(n10699), .ZN(n10704) );
  INV_X1 U13606 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21034) );
  OAI21_X1 U13607 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n21034), .A(
        n20837), .ZN(n10701) );
  INV_X1 U13608 ( .A(n10701), .ZN(n10702) );
  AOI21_X1 U13609 ( .B1(n10428), .B2(P1_EAX_REG_16__SCAN_IN), .A(n10702), .ZN(
        n10703) );
  OAI21_X1 U13610 ( .B1(n11001), .B2(n10704), .A(n10703), .ZN(n10708) );
  OAI21_X1 U13611 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n10706), .A(
        n10720), .ZN(n16037) );
  OR2_X1 U13612 ( .A1(n11004), .A2(n16037), .ZN(n10707) );
  NAND2_X1 U13613 ( .A1(n10708), .A2(n10707), .ZN(n14766) );
  INV_X1 U13614 ( .A(n14766), .ZN(n10709) );
  AOI22_X1 U13615 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10713) );
  AOI22_X1 U13616 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13617 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13618 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10710) );
  NAND4_X1 U13619 ( .A1(n10713), .A2(n10712), .A3(n10711), .A4(n10710), .ZN(
        n10719) );
  AOI22_X1 U13620 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9676), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U13621 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10980), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13622 ( .A1(n10979), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10715) );
  AOI22_X1 U13623 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10714) );
  NAND4_X1 U13624 ( .A1(n10717), .A2(n10716), .A3(n10715), .A4(n10714), .ZN(
        n10718) );
  OR2_X1 U13625 ( .A1(n10719), .A2(n10718), .ZN(n10723) );
  INV_X1 U13626 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14834) );
  XNOR2_X1 U13627 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n10738), .ZN(
        n14976) );
  AOI22_X1 U13628 ( .A1(n13628), .A2(n14976), .B1(n11005), .B2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10721) );
  OAI21_X1 U13629 ( .B1(n10905), .B2(n14834), .A(n10721), .ZN(n10722) );
  AOI22_X1 U13630 ( .A1(n10987), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10727) );
  AOI22_X1 U13631 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U13632 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10725) );
  AOI22_X1 U13633 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10724) );
  NAND4_X1 U13634 ( .A1(n10727), .A2(n10726), .A3(n10725), .A4(n10724), .ZN(
        n10733) );
  AOI22_X1 U13635 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U13636 ( .A1(n10979), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10730) );
  AOI22_X1 U13637 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10980), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10729) );
  AOI22_X1 U13638 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10728) );
  NAND4_X1 U13639 ( .A1(n10731), .A2(n10730), .A3(n10729), .A4(n10728), .ZN(
        n10732) );
  NOR2_X1 U13640 ( .A1(n10733), .A2(n10732), .ZN(n10737) );
  OAI21_X1 U13641 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n21034), .A(
        n20837), .ZN(n10734) );
  INV_X1 U13642 ( .A(n10734), .ZN(n10735) );
  AOI21_X1 U13643 ( .B1(n10428), .B2(P1_EAX_REG_18__SCAN_IN), .A(n10735), .ZN(
        n10736) );
  OAI21_X1 U13644 ( .B1(n11001), .B2(n10737), .A(n10736), .ZN(n10744) );
  INV_X1 U13645 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10741) );
  INV_X1 U13646 ( .A(n10739), .ZN(n10740) );
  NAND2_X1 U13647 ( .A1(n10741), .A2(n10740), .ZN(n10742) );
  AND2_X1 U13648 ( .A1(n10775), .A2(n10742), .ZN(n14962) );
  NAND2_X1 U13649 ( .A1(n14962), .A2(n10426), .ZN(n10743) );
  AOI22_X1 U13650 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10748) );
  AOI22_X1 U13651 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U13652 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10746) );
  AOI22_X1 U13653 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10745) );
  NAND4_X1 U13654 ( .A1(n10748), .A2(n10747), .A3(n10746), .A4(n10745), .ZN(
        n10754) );
  AOI22_X1 U13655 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9676), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10752) );
  AOI22_X1 U13656 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10751) );
  AOI22_X1 U13657 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10750) );
  AOI22_X1 U13658 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10749) );
  NAND4_X1 U13659 ( .A1(n10752), .A2(n10751), .A3(n10750), .A4(n10749), .ZN(
        n10753) );
  NOR2_X1 U13660 ( .A1(n10754), .A2(n10753), .ZN(n10757) );
  INV_X1 U13661 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10774) );
  AOI21_X1 U13662 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n10774), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10755) );
  AOI21_X1 U13663 ( .B1(n10428), .B2(P1_EAX_REG_19__SCAN_IN), .A(n10755), .ZN(
        n10756) );
  OAI21_X1 U13664 ( .B1(n11001), .B2(n10757), .A(n10756), .ZN(n10759) );
  XNOR2_X1 U13665 ( .A(n10775), .B(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14950) );
  NAND2_X1 U13666 ( .A1(n14950), .A2(n10426), .ZN(n10758) );
  AOI22_X1 U13667 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9676), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10763) );
  AOI22_X1 U13668 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U13669 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10761) );
  AOI22_X1 U13670 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10760) );
  NAND4_X1 U13671 ( .A1(n10763), .A2(n10762), .A3(n10761), .A4(n10760), .ZN(
        n10769) );
  AOI22_X1 U13672 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10767) );
  AOI22_X1 U13673 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10766) );
  AOI22_X1 U13674 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10980), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10765) );
  AOI22_X1 U13675 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10764) );
  NAND4_X1 U13676 ( .A1(n10767), .A2(n10766), .A3(n10765), .A4(n10764), .ZN(
        n10768) );
  NOR2_X1 U13677 ( .A1(n10769), .A2(n10768), .ZN(n10773) );
  NAND2_X1 U13678 ( .A1(n20837), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10770) );
  NAND2_X1 U13679 ( .A1(n11004), .A2(n10770), .ZN(n10771) );
  AOI21_X1 U13680 ( .B1(n10428), .B2(P1_EAX_REG_20__SCAN_IN), .A(n10771), .ZN(
        n10772) );
  OAI21_X1 U13681 ( .B1(n11001), .B2(n10773), .A(n10772), .ZN(n10780) );
  INV_X1 U13682 ( .A(n10776), .ZN(n10777) );
  INV_X1 U13683 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14638) );
  NAND2_X1 U13684 ( .A1(n10777), .A2(n14638), .ZN(n10778) );
  NAND2_X1 U13685 ( .A1(n10812), .A2(n10778), .ZN(n14943) );
  OR2_X1 U13686 ( .A1(n14943), .A2(n11004), .ZN(n10779) );
  NAND2_X1 U13687 ( .A1(n10780), .A2(n10779), .ZN(n14637) );
  AOI22_X1 U13688 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10785) );
  AOI22_X1 U13689 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9676), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10784) );
  AOI22_X1 U13690 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10783) );
  AOI22_X1 U13691 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10980), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10782) );
  NAND4_X1 U13692 ( .A1(n10785), .A2(n10784), .A3(n10783), .A4(n10782), .ZN(
        n10791) );
  AOI22_X1 U13693 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U13694 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10788) );
  AOI22_X1 U13695 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10787) );
  AOI22_X1 U13696 ( .A1(n10979), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10786) );
  NAND4_X1 U13697 ( .A1(n10789), .A2(n10788), .A3(n10787), .A4(n10786), .ZN(
        n10790) );
  NOR2_X1 U13698 ( .A1(n10791), .A2(n10790), .ZN(n10795) );
  NAND2_X1 U13699 ( .A1(n20837), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10792) );
  NAND2_X1 U13700 ( .A1(n11004), .A2(n10792), .ZN(n10793) );
  AOI21_X1 U13701 ( .B1(n10428), .B2(P1_EAX_REG_21__SCAN_IN), .A(n10793), .ZN(
        n10794) );
  OAI21_X1 U13702 ( .B1(n11001), .B2(n10795), .A(n10794), .ZN(n10797) );
  XNOR2_X1 U13703 ( .A(n10812), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14933) );
  NAND2_X1 U13704 ( .A1(n14933), .A2(n10426), .ZN(n10796) );
  NAND2_X1 U13705 ( .A1(n10797), .A2(n10796), .ZN(n14626) );
  AOI22_X1 U13706 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10956), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10801) );
  AOI22_X1 U13707 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10800) );
  AOI22_X1 U13708 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10799) );
  AOI22_X1 U13709 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10798) );
  NAND4_X1 U13710 ( .A1(n10801), .A2(n10800), .A3(n10799), .A4(n10798), .ZN(
        n10807) );
  AOI22_X1 U13711 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10805) );
  AOI22_X1 U13712 ( .A1(n10987), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10804) );
  AOI22_X1 U13713 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10980), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U13714 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10802) );
  NAND4_X1 U13715 ( .A1(n10805), .A2(n10804), .A3(n10803), .A4(n10802), .ZN(
        n10806) );
  NOR2_X1 U13716 ( .A1(n10807), .A2(n10806), .ZN(n10811) );
  NAND2_X1 U13717 ( .A1(n20837), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10808) );
  NAND2_X1 U13718 ( .A1(n11004), .A2(n10808), .ZN(n10809) );
  AOI21_X1 U13719 ( .B1(n10428), .B2(P1_EAX_REG_22__SCAN_IN), .A(n10809), .ZN(
        n10810) );
  OAI21_X1 U13720 ( .B1(n11001), .B2(n10811), .A(n10810), .ZN(n10819) );
  INV_X1 U13721 ( .A(n10814), .ZN(n10816) );
  INV_X1 U13722 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10815) );
  NAND2_X1 U13723 ( .A1(n10816), .A2(n10815), .ZN(n10817) );
  NAND2_X1 U13724 ( .A1(n10876), .A2(n10817), .ZN(n14926) );
  AOI22_X1 U13725 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U13726 ( .A1(n10987), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U13727 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U13728 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10821) );
  NAND4_X1 U13729 ( .A1(n10824), .A2(n10823), .A3(n10822), .A4(n10821), .ZN(
        n10830) );
  AOI22_X1 U13730 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U13731 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10957), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U13732 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10826) );
  AOI22_X1 U13733 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10825) );
  NAND4_X1 U13734 ( .A1(n10828), .A2(n10827), .A3(n10826), .A4(n10825), .ZN(
        n10829) );
  NOR2_X1 U13735 ( .A1(n10830), .A2(n10829), .ZN(n10850) );
  AOI22_X1 U13736 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n10956), .B1(
        n9676), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10835) );
  AOI22_X1 U13737 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10987), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10834) );
  AOI22_X1 U13738 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10833) );
  AOI22_X1 U13739 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10832) );
  NAND4_X1 U13740 ( .A1(n10835), .A2(n10834), .A3(n10833), .A4(n10832), .ZN(
        n10842) );
  AOI22_X1 U13741 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10962), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U13742 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n10986), .B1(
        n9674), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10839) );
  AOI22_X1 U13743 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U13744 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n9666), .B1(
        n10980), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10837) );
  NAND4_X1 U13745 ( .A1(n10840), .A2(n10839), .A3(n10838), .A4(n10837), .ZN(
        n10841) );
  NOR2_X1 U13746 ( .A1(n10842), .A2(n10841), .ZN(n10849) );
  XOR2_X1 U13747 ( .A(n10850), .B(n10849), .Z(n10843) );
  NAND2_X1 U13748 ( .A1(n10843), .A2(n10970), .ZN(n10848) );
  NAND2_X1 U13749 ( .A1(n20837), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10844) );
  NAND2_X1 U13750 ( .A1(n11004), .A2(n10844), .ZN(n10845) );
  AOI21_X1 U13751 ( .B1(n10428), .B2(P1_EAX_REG_23__SCAN_IN), .A(n10845), .ZN(
        n10847) );
  XNOR2_X1 U13752 ( .A(n10876), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14597) );
  NOR2_X1 U13753 ( .A1(n10850), .A2(n10849), .ZN(n10882) );
  AOI22_X1 U13754 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U13755 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U13756 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10852) );
  AOI22_X1 U13757 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10851) );
  NAND4_X1 U13758 ( .A1(n10854), .A2(n10853), .A3(n10852), .A4(n10851), .ZN(
        n10860) );
  AOI22_X1 U13759 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U13760 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10831), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U13761 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10856) );
  AOI22_X1 U13762 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10855) );
  NAND4_X1 U13763 ( .A1(n10858), .A2(n10857), .A3(n10856), .A4(n10855), .ZN(
        n10859) );
  OR2_X1 U13764 ( .A1(n10860), .A2(n10859), .ZN(n10880) );
  NAND2_X1 U13765 ( .A1(n10882), .A2(n10880), .ZN(n10891) );
  AOI22_X1 U13766 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10864) );
  AOI22_X1 U13767 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10863) );
  AOI22_X1 U13768 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U13769 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10861) );
  NAND4_X1 U13770 ( .A1(n10864), .A2(n10863), .A3(n10862), .A4(n10861), .ZN(
        n10870) );
  AOI22_X1 U13771 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9676), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10868) );
  AOI22_X1 U13772 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10867) );
  AOI22_X1 U13773 ( .A1(n10987), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U13774 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10250), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10865) );
  NAND4_X1 U13775 ( .A1(n10868), .A2(n10867), .A3(n10866), .A4(n10865), .ZN(
        n10869) );
  NOR2_X1 U13776 ( .A1(n10870), .A2(n10869), .ZN(n10892) );
  XOR2_X1 U13777 ( .A(n10891), .B(n10892), .Z(n10871) );
  NAND2_X1 U13778 ( .A1(n10871), .A2(n10970), .ZN(n10875) );
  NAND2_X1 U13779 ( .A1(n20837), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10872) );
  NAND2_X1 U13780 ( .A1(n11004), .A2(n10872), .ZN(n10873) );
  AOI21_X1 U13781 ( .B1(n10428), .B2(P1_EAX_REG_25__SCAN_IN), .A(n10873), .ZN(
        n10874) );
  NAND2_X1 U13782 ( .A1(n10875), .A2(n10874), .ZN(n10879) );
  XNOR2_X1 U13783 ( .A(n10909), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14896) );
  NAND2_X1 U13784 ( .A1(n14896), .A2(n10426), .ZN(n10878) );
  NAND2_X1 U13785 ( .A1(n10879), .A2(n10878), .ZN(n14572) );
  INV_X1 U13786 ( .A(n10880), .ZN(n10881) );
  XNOR2_X1 U13787 ( .A(n10882), .B(n10881), .ZN(n10885) );
  INV_X1 U13788 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14803) );
  NAND2_X1 U13789 ( .A1(n20837), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10883) );
  OAI211_X1 U13790 ( .C1(n10905), .C2(n14803), .A(n11004), .B(n10883), .ZN(
        n10884) );
  AOI21_X1 U13791 ( .B1(n10885), .B2(n10970), .A(n10884), .ZN(n10890) );
  INV_X1 U13792 ( .A(n10886), .ZN(n10887) );
  INV_X1 U13793 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14588) );
  NAND2_X1 U13794 ( .A1(n10887), .A2(n14588), .ZN(n10888) );
  NAND2_X1 U13795 ( .A1(n10909), .A2(n10888), .ZN(n14909) );
  NOR2_X1 U13796 ( .A1(n14909), .A2(n11004), .ZN(n10889) );
  NOR2_X1 U13797 ( .A1(n10892), .A2(n10891), .ZN(n10915) );
  AOI22_X1 U13798 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10896) );
  AOI22_X1 U13799 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U13800 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U13801 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10820), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10893) );
  NAND4_X1 U13802 ( .A1(n10896), .A2(n10895), .A3(n10894), .A4(n10893), .ZN(
        n10902) );
  AOI22_X1 U13803 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10900) );
  AOI22_X1 U13804 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10899) );
  AOI22_X1 U13805 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10898) );
  AOI22_X1 U13806 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10897) );
  NAND4_X1 U13807 ( .A1(n10900), .A2(n10899), .A3(n10898), .A4(n10897), .ZN(
        n10901) );
  OR2_X1 U13808 ( .A1(n10902), .A2(n10901), .ZN(n10914) );
  INV_X1 U13809 ( .A(n10914), .ZN(n10903) );
  XNOR2_X1 U13810 ( .A(n10915), .B(n10903), .ZN(n10907) );
  INV_X1 U13811 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14794) );
  NAND2_X1 U13812 ( .A1(n20837), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10904) );
  OAI211_X1 U13813 ( .C1(n10905), .C2(n14794), .A(n11004), .B(n10904), .ZN(
        n10906) );
  AOI21_X1 U13814 ( .B1(n10907), .B2(n10970), .A(n10906), .ZN(n10913) );
  INV_X1 U13815 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10908) );
  INV_X1 U13816 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14561) );
  NAND2_X1 U13817 ( .A1(n10910), .A2(n14561), .ZN(n10911) );
  NAND2_X1 U13818 ( .A1(n10931), .A2(n10911), .ZN(n14888) );
  NOR2_X1 U13819 ( .A1(n14888), .A2(n11004), .ZN(n10912) );
  NAND2_X1 U13820 ( .A1(n10915), .A2(n10914), .ZN(n10936) );
  AOI22_X1 U13821 ( .A1(n10979), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10919) );
  AOI22_X1 U13822 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10250), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10918) );
  AOI22_X1 U13823 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U13824 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10916) );
  NAND4_X1 U13825 ( .A1(n10919), .A2(n10918), .A3(n10917), .A4(n10916), .ZN(
        n10925) );
  AOI22_X1 U13826 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U13827 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10986), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U13828 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10921) );
  AOI22_X1 U13829 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9666), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10920) );
  NAND4_X1 U13830 ( .A1(n10923), .A2(n10922), .A3(n10921), .A4(n10920), .ZN(
        n10924) );
  NOR2_X1 U13831 ( .A1(n10925), .A2(n10924), .ZN(n10937) );
  XOR2_X1 U13832 ( .A(n10936), .B(n10937), .Z(n10926) );
  NAND2_X1 U13833 ( .A1(n10926), .A2(n10970), .ZN(n10929) );
  INV_X1 U13834 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10930) );
  NOR2_X1 U13835 ( .A1(n10930), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10927) );
  AOI211_X1 U13836 ( .C1(n10428), .C2(P1_EAX_REG_27__SCAN_IN), .A(n10426), .B(
        n10927), .ZN(n10928) );
  XNOR2_X1 U13837 ( .A(n10931), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14877) );
  AOI22_X1 U13838 ( .A1(n10929), .A2(n10928), .B1(n13628), .B2(n14877), .ZN(
        n14546) );
  INV_X1 U13839 ( .A(n10932), .ZN(n10934) );
  INV_X1 U13840 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10933) );
  NAND2_X1 U13841 ( .A1(n10934), .A2(n10933), .ZN(n10935) );
  NAND2_X1 U13842 ( .A1(n10976), .A2(n10935), .ZN(n14870) );
  NOR2_X1 U13843 ( .A1(n10937), .A2(n10936), .ZN(n10954) );
  AOI22_X1 U13844 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10987), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U13845 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U13846 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U13847 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10939) );
  NAND4_X1 U13848 ( .A1(n10942), .A2(n10941), .A3(n10940), .A4(n10939), .ZN(
        n10948) );
  AOI22_X1 U13849 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10946) );
  AOI22_X1 U13850 ( .A1(n10986), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10945) );
  AOI22_X1 U13851 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U13852 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10943) );
  NAND4_X1 U13853 ( .A1(n10946), .A2(n10945), .A3(n10944), .A4(n10943), .ZN(
        n10947) );
  OR2_X1 U13854 ( .A1(n10948), .A2(n10947), .ZN(n10953) );
  XNOR2_X1 U13855 ( .A(n10954), .B(n10953), .ZN(n10951) );
  AOI21_X1 U13856 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20837), .A(
        n13628), .ZN(n10950) );
  NAND2_X1 U13857 ( .A1(n11006), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n10949) );
  OAI211_X1 U13858 ( .C1(n10951), .C2(n11001), .A(n10950), .B(n10949), .ZN(
        n10952) );
  OAI21_X1 U13859 ( .B1(n11004), .B2(n14870), .A(n10952), .ZN(n12834) );
  NAND2_X1 U13860 ( .A1(n10954), .A2(n10953), .ZN(n10995) );
  AOI22_X1 U13861 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10986), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10961) );
  AOI22_X1 U13862 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U13863 ( .A1(n10957), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U13864 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10958) );
  NAND4_X1 U13865 ( .A1(n10961), .A2(n10960), .A3(n10959), .A4(n10958), .ZN(
        n10969) );
  AOI22_X1 U13866 ( .A1(n10962), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10967) );
  AOI22_X1 U13867 ( .A1(n9674), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10966) );
  AOI22_X1 U13868 ( .A1(n10987), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10965) );
  AOI22_X1 U13869 ( .A1(n10980), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10964) );
  NAND4_X1 U13870 ( .A1(n10967), .A2(n10966), .A3(n10965), .A4(n10964), .ZN(
        n10968) );
  NOR2_X1 U13871 ( .A1(n10969), .A2(n10968), .ZN(n10996) );
  XOR2_X1 U13872 ( .A(n10995), .B(n10996), .Z(n10971) );
  NAND2_X1 U13873 ( .A1(n10971), .A2(n10970), .ZN(n10974) );
  INV_X1 U13874 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10975) );
  NOR2_X1 U13875 ( .A1(n10975), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10972) );
  AOI211_X1 U13876 ( .C1(n10428), .C2(P1_EAX_REG_29__SCAN_IN), .A(n10426), .B(
        n10972), .ZN(n10973) );
  XNOR2_X1 U13877 ( .A(n10976), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14528) );
  INV_X1 U13878 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14515) );
  XNOR2_X1 U13879 ( .A(n12253), .B(n14515), .ZN(n14860) );
  AOI22_X1 U13880 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n9674), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10985) );
  AOI22_X1 U13881 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10979), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10984) );
  AOI22_X1 U13882 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10955), .B1(
        n10980), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10983) );
  AOI22_X1 U13883 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10982) );
  NAND4_X1 U13884 ( .A1(n10985), .A2(n10984), .A3(n10983), .A4(n10982), .ZN(
        n10994) );
  AOI22_X1 U13885 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n10962), .B1(
        n10986), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10992) );
  AOI22_X1 U13886 ( .A1(n10987), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10957), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10991) );
  AOI22_X1 U13887 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10990) );
  AOI22_X1 U13888 ( .A1(n9676), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10988), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10989) );
  NAND4_X1 U13889 ( .A1(n10992), .A2(n10991), .A3(n10990), .A4(n10989), .ZN(
        n10993) );
  NOR2_X1 U13890 ( .A1(n10994), .A2(n10993), .ZN(n10998) );
  NOR2_X1 U13891 ( .A1(n10996), .A2(n10995), .ZN(n10997) );
  XOR2_X1 U13892 ( .A(n10998), .B(n10997), .Z(n11002) );
  AOI21_X1 U13893 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20837), .A(
        n13628), .ZN(n11000) );
  NAND2_X1 U13894 ( .A1(n11006), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n10999) );
  OAI211_X1 U13895 ( .C1(n11002), .C2(n11001), .A(n11000), .B(n10999), .ZN(
        n11003) );
  OAI21_X1 U13896 ( .B1(n11004), .B2(n14860), .A(n11003), .ZN(n11088) );
  AOI22_X1 U13897 ( .A1(n11006), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n11005), .ZN(n11007) );
  NAND2_X1 U13898 ( .A1(n10183), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11009) );
  NAND2_X1 U13899 ( .A1(n11010), .A2(n11009), .ZN(n11021) );
  XNOR2_X1 U13900 ( .A(n9920), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11016) );
  INV_X1 U13901 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20236) );
  NOR2_X1 U13902 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20236), .ZN(
        n11012) );
  NAND2_X1 U13903 ( .A1(n11061), .A2(n11045), .ZN(n11054) );
  NAND2_X1 U13904 ( .A1(n11061), .A2(n11024), .ZN(n11052) );
  NAND3_X1 U13905 ( .A1(n16175), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n11013), .ZN(n11059) );
  INV_X1 U13906 ( .A(n11045), .ZN(n11049) );
  AOI21_X1 U13907 ( .B1(n11016), .B2(n11015), .A(n11014), .ZN(n11017) );
  INV_X1 U13908 ( .A(n11017), .ZN(n11056) );
  OR2_X1 U13909 ( .A1(n13632), .A2(n14160), .ZN(n11018) );
  NAND2_X1 U13910 ( .A1(n11018), .A2(n13310), .ZN(n11041) );
  XNOR2_X1 U13911 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11019) );
  XNOR2_X1 U13912 ( .A(n11020), .B(n11019), .ZN(n11058) );
  NAND2_X1 U13913 ( .A1(n11021), .A2(n11026), .ZN(n11022) );
  NAND2_X1 U13914 ( .A1(n11023), .A2(n11022), .ZN(n11057) );
  INV_X1 U13915 ( .A(n11036), .ZN(n11025) );
  NOR2_X1 U13916 ( .A1(n11057), .A2(n11025), .ZN(n11031) );
  OAI21_X1 U13917 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20692), .A(
        n11026), .ZN(n11027) );
  NOR2_X1 U13918 ( .A1(n11040), .A2(n11027), .ZN(n11030) );
  INV_X1 U13919 ( .A(n11027), .ZN(n11028) );
  OAI211_X1 U13920 ( .C1(n13632), .C2(n12247), .A(n11041), .B(n11028), .ZN(
        n11029) );
  OAI21_X1 U13921 ( .B1(n11045), .B2(n11030), .A(n11029), .ZN(n11033) );
  AND2_X1 U13922 ( .A1(n11031), .A2(n11033), .ZN(n11039) );
  OAI21_X1 U13923 ( .B1(n11040), .B2(n11058), .A(n11041), .ZN(n11032) );
  AOI21_X1 U13924 ( .B1(n11046), .B2(n11058), .A(n11032), .ZN(n11038) );
  INV_X1 U13925 ( .A(n11057), .ZN(n11035) );
  NOR2_X1 U13926 ( .A1(n11036), .A2(n11033), .ZN(n11034) );
  AOI211_X1 U13927 ( .C1(n11036), .C2(n20258), .A(n11035), .B(n11034), .ZN(
        n11037) );
  OAI33_X1 U13928 ( .A1(n11041), .A2(n11040), .A3(n11058), .B1(n11039), .B2(
        n11038), .B3(n11037), .ZN(n11044) );
  NAND2_X1 U13929 ( .A1(n11042), .A2(n11056), .ZN(n11043) );
  AOI22_X1 U13930 ( .A1(n11045), .A2(n11056), .B1(n11044), .B2(n11043), .ZN(
        n11048) );
  NOR2_X1 U13931 ( .A1(n11046), .A2(n11059), .ZN(n11047) );
  OAI22_X1 U13932 ( .A1(n11059), .A2(n11049), .B1(n11048), .B2(n11047), .ZN(
        n11050) );
  AOI21_X1 U13933 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20914), .A(
        n11050), .ZN(n11051) );
  NAND2_X1 U13934 ( .A1(n11052), .A2(n11051), .ZN(n11053) );
  INV_X1 U13935 ( .A(n10306), .ZN(n15164) );
  NOR2_X1 U13936 ( .A1(n14482), .A2(n13169), .ZN(n11055) );
  NAND2_X1 U13937 ( .A1(n15164), .A2(n11055), .ZN(n14471) );
  NOR3_X1 U13938 ( .A1(n11058), .A2(n11057), .A3(n11056), .ZN(n11060) );
  OAI21_X1 U13939 ( .B1(n11061), .B2(n11060), .A(n11059), .ZN(n14475) );
  AND2_X1 U13940 ( .A1(n14475), .A2(n11062), .ZN(n14480) );
  NAND2_X1 U13941 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20918) );
  NAND3_X1 U13942 ( .A1(n14480), .A2(n13310), .A3(n20918), .ZN(n11063) );
  INV_X1 U13943 ( .A(n11065), .ZN(n11066) );
  NAND2_X1 U13944 ( .A1(n11066), .A2(n20918), .ZN(n11067) );
  INV_X1 U13945 ( .A(n13330), .ZN(n13178) );
  INV_X1 U13946 ( .A(n20289), .ZN(n14161) );
  NAND3_X1 U13947 ( .A1(n14161), .A2(n13329), .A3(n20280), .ZN(n11090) );
  OAI22_X1 U13948 ( .A1(n14483), .A2(n11067), .B1(n13178), .B2(n11090), .ZN(
        n11068) );
  OR2_X1 U13949 ( .A1(n14849), .A2(n13311), .ZN(n11082) );
  NOR4_X1 U13950 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n11073) );
  NOR4_X1 U13951 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n11072) );
  NOR4_X1 U13952 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n11071) );
  NOR4_X1 U13953 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n11070) );
  AND4_X1 U13954 ( .A1(n11073), .A2(n11072), .A3(n11071), .A4(n11070), .ZN(
        n11078) );
  NOR4_X1 U13955 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n11076) );
  NOR4_X1 U13956 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n11075) );
  NOR4_X1 U13957 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n11074) );
  INV_X1 U13958 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20858) );
  AND4_X1 U13959 ( .A1(n11076), .A2(n11075), .A3(n11074), .A4(n20858), .ZN(
        n11077) );
  NAND2_X1 U13960 ( .A1(n11078), .A2(n11077), .ZN(n11079) );
  AND2_X2 U13961 ( .A1(n11079), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20238)
         );
  AOI22_X1 U13962 ( .A1(n11080), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14849), .ZN(n11081) );
  INV_X1 U13963 ( .A(n11081), .ZN(n11085) );
  INV_X1 U13964 ( .A(n11082), .ZN(n11083) );
  NAND2_X1 U13965 ( .A1(n11083), .A2(n20238), .ZN(n14823) );
  INV_X1 U13966 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20287) );
  NOR2_X1 U13967 ( .A1(n14823), .A2(n20287), .ZN(n11084) );
  NOR2_X1 U13968 ( .A1(n11085), .A2(n11084), .ZN(n11086) );
  NAND2_X1 U13969 ( .A1(n11087), .A2(n11086), .ZN(P1_U2873) );
  AND2_X1 U13970 ( .A1(n9636), .A2(n10299), .ZN(n11089) );
  NAND2_X1 U13971 ( .A1(n14483), .A2(n14474), .ZN(n11093) );
  INV_X1 U13972 ( .A(n11090), .ZN(n11091) );
  NAND4_X1 U13973 ( .A1(n11091), .A2(n10304), .A3(n9636), .A4(n13165), .ZN(
        n11092) );
  OR2_X2 U13974 ( .A1(n14769), .A2(n14161), .ZN(n14779) );
  INV_X1 U13975 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n11095) );
  NAND2_X1 U13976 ( .A1(n9636), .A2(n11095), .ZN(n11096) );
  OAI211_X1 U13977 ( .C1(n11180), .C2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n11096), .B(n11155), .ZN(n11097) );
  NAND2_X1 U13978 ( .A1(n11162), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11102) );
  INV_X1 U13979 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n11100) );
  NAND2_X1 U13980 ( .A1(n11155), .A2(n11100), .ZN(n11101) );
  NAND2_X1 U13981 ( .A1(n11102), .A2(n11101), .ZN(n13082) );
  MUX2_X1 U13982 ( .A(n11184), .B(n11162), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n11104) );
  NAND2_X1 U13983 ( .A1(n14492), .A2(n11180), .ZN(n11137) );
  NAND2_X1 U13984 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14492), .ZN(
        n11103) );
  NAND3_X1 U13985 ( .A1(n11104), .A2(n11137), .A3(n11103), .ZN(n13303) );
  MUX2_X1 U13986 ( .A(n11175), .B(n11155), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n11106) );
  INV_X1 U13987 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20197) );
  NAND2_X1 U13988 ( .A1(n11176), .A2(n20197), .ZN(n11105) );
  NAND2_X1 U13989 ( .A1(n13471), .A2(n13470), .ZN(n13469) );
  MUX2_X1 U13990 ( .A(n11184), .B(n11162), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n11108) );
  INV_X1 U13991 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20188) );
  OR2_X1 U13992 ( .A1(n20188), .A2(n9658), .ZN(n11107) );
  AND3_X1 U13993 ( .A1(n11108), .A2(n11137), .A3(n11107), .ZN(n13380) );
  OR2_X1 U13994 ( .A1(n11175), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n11112) );
  INV_X1 U13995 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16169) );
  INV_X1 U13996 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n11109) );
  NAND2_X1 U13997 ( .A1(n9636), .A2(n11109), .ZN(n11110) );
  OAI211_X1 U13998 ( .C1(n14490), .C2(n16169), .A(n11110), .B(n11162), .ZN(
        n11111) );
  NAND2_X1 U13999 ( .A1(n11112), .A2(n11111), .ZN(n13367) );
  INV_X1 U14000 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16148) );
  MUX2_X1 U14001 ( .A(n11184), .B(n11162), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n11114) );
  OAI211_X1 U14002 ( .C1(n9658), .C2(n16148), .A(n11114), .B(n11137), .ZN(
        n13657) );
  OR2_X1 U14003 ( .A1(n11175), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n11117) );
  INV_X1 U14004 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16157) );
  INV_X1 U14005 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13660) );
  NAND2_X1 U14006 ( .A1(n9658), .A2(n13660), .ZN(n11115) );
  OAI211_X1 U14007 ( .C1(n14490), .C2(n16157), .A(n11115), .B(n11162), .ZN(
        n11116) );
  NAND2_X1 U14008 ( .A1(n13657), .A2(n13656), .ZN(n11118) );
  NOR2_X2 U14009 ( .A1(n13366), .A2(n11118), .ZN(n13696) );
  MUX2_X1 U14010 ( .A(n11184), .B(n11162), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n11120) );
  INV_X1 U14011 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16151) );
  OR2_X1 U14012 ( .A1(n16151), .A2(n9658), .ZN(n11119) );
  NAND3_X1 U14013 ( .A1(n11120), .A2(n11137), .A3(n11119), .ZN(n13695) );
  OR2_X1 U14014 ( .A1(n11175), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n11123) );
  INV_X1 U14015 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16139) );
  INV_X1 U14016 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20025) );
  NAND2_X1 U14017 ( .A1(n9658), .A2(n20025), .ZN(n11121) );
  OAI211_X1 U14018 ( .C1(n14490), .C2(n16139), .A(n11121), .B(n11162), .ZN(
        n11122) );
  NAND2_X1 U14019 ( .A1(n11123), .A2(n11122), .ZN(n13747) );
  OR2_X1 U14020 ( .A1(n11184), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n11128) );
  INV_X1 U14021 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n11125) );
  NAND2_X1 U14022 ( .A1(n9658), .A2(n11125), .ZN(n11126) );
  OAI211_X1 U14023 ( .C1(n11180), .C2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n11126), .B(n11155), .ZN(n11127) );
  MUX2_X1 U14024 ( .A(n11175), .B(n11155), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n11130) );
  INV_X1 U14025 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16116) );
  NAND2_X1 U14026 ( .A1(n11176), .A2(n16116), .ZN(n11129) );
  MUX2_X1 U14027 ( .A(n11184), .B(n11162), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n11132) );
  NAND2_X1 U14028 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14492), .ZN(
        n11131) );
  NAND3_X1 U14029 ( .A1(n11132), .A2(n11137), .A3(n11131), .ZN(n14006) );
  INV_X1 U14030 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n11133) );
  MUX2_X1 U14031 ( .A(n11155), .B(n11175), .S(n11133), .Z(n11135) );
  NAND2_X1 U14032 ( .A1(n11176), .A2(n12230), .ZN(n11134) );
  NAND2_X1 U14033 ( .A1(n11135), .A2(n11134), .ZN(n14707) );
  OR2_X2 U14034 ( .A1(n14708), .A2(n14707), .ZN(n14773) );
  MUX2_X1 U14035 ( .A(n11184), .B(n11162), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n11138) );
  INV_X1 U14036 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16114) );
  OR2_X1 U14037 ( .A1(n16114), .A2(n9658), .ZN(n11136) );
  AND3_X1 U14038 ( .A1(n11138), .A2(n11137), .A3(n11136), .ZN(n14772) );
  OR2_X2 U14039 ( .A1(n14773), .A2(n14772), .ZN(n14775) );
  MUX2_X1 U14040 ( .A(n11175), .B(n11155), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n11140) );
  INV_X1 U14041 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14042) );
  NAND2_X1 U14042 ( .A1(n11176), .A2(n14042), .ZN(n11139) );
  NAND2_X1 U14043 ( .A1(n11140), .A2(n11139), .ZN(n14692) );
  OR2_X1 U14044 ( .A1(n11184), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n11143) );
  INV_X1 U14045 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n16000) );
  NAND2_X1 U14046 ( .A1(n9658), .A2(n16000), .ZN(n11141) );
  OAI211_X1 U14047 ( .C1(n11180), .C2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11141), .B(n11155), .ZN(n11142) );
  NAND2_X1 U14048 ( .A1(n11143), .A2(n11142), .ZN(n14030) );
  OR2_X1 U14049 ( .A1(n11175), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n11146) );
  INV_X1 U14050 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14974) );
  INV_X1 U14051 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14681) );
  NAND2_X1 U14052 ( .A1(n9658), .A2(n14681), .ZN(n11144) );
  OAI211_X1 U14053 ( .C1(n14490), .C2(n14974), .A(n11144), .B(n11162), .ZN(
        n11145) );
  NAND2_X1 U14054 ( .A1(n11146), .A2(n11145), .ZN(n14675) );
  OR2_X1 U14055 ( .A1(n11184), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n11149) );
  INV_X1 U14056 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14666) );
  NAND2_X1 U14057 ( .A1(n9658), .A2(n14666), .ZN(n11147) );
  OAI211_X1 U14058 ( .C1(n11180), .C2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n11147), .B(n11155), .ZN(n11148) );
  AND2_X1 U14059 ( .A1(n11149), .A2(n11148), .ZN(n14663) );
  OR2_X1 U14060 ( .A1(n11175), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n11152) );
  INV_X1 U14061 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15138) );
  INV_X1 U14062 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14758) );
  NAND2_X1 U14063 ( .A1(n9658), .A2(n14758), .ZN(n11150) );
  OAI211_X1 U14064 ( .C1(n14490), .C2(n15138), .A(n11150), .B(n11162), .ZN(
        n11151) );
  AND2_X1 U14065 ( .A1(n11152), .A2(n11151), .ZN(n14650) );
  MUX2_X1 U14066 ( .A(n11184), .B(n11162), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n11154) );
  INV_X1 U14067 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15123) );
  OR2_X1 U14068 ( .A1(n9636), .A2(n15123), .ZN(n11153) );
  NAND2_X1 U14069 ( .A1(n11154), .A2(n11153), .ZN(n14640) );
  MUX2_X1 U14070 ( .A(n11175), .B(n11155), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n11157) );
  INV_X1 U14071 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12239) );
  NAND2_X1 U14072 ( .A1(n11176), .A2(n12239), .ZN(n11156) );
  NAND2_X1 U14073 ( .A1(n11157), .A2(n11156), .ZN(n14629) );
  OR2_X1 U14074 ( .A1(n11184), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n11161) );
  INV_X1 U14075 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n11158) );
  NAND2_X1 U14076 ( .A1(n9658), .A2(n11158), .ZN(n11159) );
  OAI211_X1 U14077 ( .C1(n11180), .C2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n11159), .B(n11155), .ZN(n11160) );
  AND2_X1 U14078 ( .A1(n11161), .A2(n11160), .ZN(n14612) );
  OR2_X1 U14079 ( .A1(n11175), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n11165) );
  INV_X1 U14080 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15092) );
  INV_X1 U14081 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14754) );
  NAND2_X1 U14082 ( .A1(n9658), .A2(n14754), .ZN(n11163) );
  OAI211_X1 U14083 ( .C1(n14490), .C2(n15092), .A(n11163), .B(n11162), .ZN(
        n11164) );
  AND2_X1 U14084 ( .A1(n11165), .A2(n11164), .ZN(n14599) );
  OR2_X1 U14085 ( .A1(n11184), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n11168) );
  INV_X1 U14086 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14753) );
  NAND2_X1 U14087 ( .A1(n9658), .A2(n14753), .ZN(n11166) );
  OAI211_X1 U14088 ( .C1(n11180), .C2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11166), .B(n11155), .ZN(n11167) );
  NAND2_X1 U14089 ( .A1(n11168), .A2(n11167), .ZN(n14587) );
  MUX2_X1 U14090 ( .A(n11175), .B(n11155), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n11170) );
  INV_X1 U14091 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15068) );
  NAND2_X1 U14092 ( .A1(n11176), .A2(n15068), .ZN(n11169) );
  NAND2_X1 U14093 ( .A1(n11170), .A2(n11169), .ZN(n14575) );
  OR2_X1 U14094 ( .A1(n11184), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n11174) );
  INV_X1 U14095 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n11171) );
  NAND2_X1 U14096 ( .A1(n9658), .A2(n11171), .ZN(n11172) );
  OAI211_X1 U14097 ( .C1(n11180), .C2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11172), .B(n11155), .ZN(n11173) );
  AND2_X1 U14098 ( .A1(n11174), .A2(n11173), .ZN(n14560) );
  MUX2_X1 U14099 ( .A(n11175), .B(n11155), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n11178) );
  INV_X1 U14100 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14865) );
  NAND2_X1 U14101 ( .A1(n11176), .A2(n14865), .ZN(n11177) );
  NAND2_X1 U14102 ( .A1(n11178), .A2(n11177), .ZN(n14547) );
  OR2_X1 U14103 ( .A1(n11184), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n11182) );
  INV_X1 U14104 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14540) );
  NAND2_X1 U14105 ( .A1(n9658), .A2(n14540), .ZN(n11179) );
  OAI211_X1 U14106 ( .C1(n11180), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11179), .B(n11155), .ZN(n11181) );
  NAND2_X1 U14107 ( .A1(n11182), .A2(n11181), .ZN(n12835) );
  AND2_X2 U14108 ( .A1(n14549), .A2(n12835), .ZN(n14166) );
  INV_X1 U14109 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14531) );
  NAND2_X1 U14110 ( .A1(n9658), .A2(n14531), .ZN(n11183) );
  OAI21_X1 U14111 ( .B1(n14491), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11183), .ZN(n11187) );
  OR2_X1 U14112 ( .A1(n11187), .A2(n14490), .ZN(n11186) );
  OR2_X1 U14113 ( .A1(n11184), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n11185) );
  NAND2_X1 U14114 ( .A1(n11186), .A2(n11185), .ZN(n14165) );
  AND2_X2 U14115 ( .A1(n14166), .A2(n14165), .ZN(n14488) );
  INV_X1 U14116 ( .A(n14166), .ZN(n11188) );
  INV_X1 U14117 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15018) );
  OR2_X1 U14118 ( .A1(n9658), .A2(n15018), .ZN(n11190) );
  NAND2_X1 U14119 ( .A1(n14491), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n11189) );
  NAND2_X1 U14120 ( .A1(n11190), .A2(n11189), .ZN(n14489) );
  INV_X1 U14121 ( .A(n14517), .ZN(n11195) );
  INV_X1 U14122 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n11192) );
  BUF_X4 U14123 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n15832) );
  XNOR2_X1 U14124 ( .A(n15832), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11203) );
  NAND2_X1 U14125 ( .A1(n11203), .A2(n11204), .ZN(n11205) );
  NAND2_X1 U14126 ( .A1(n19956), .A2(n15832), .ZN(n11197) );
  NAND2_X1 U14127 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19946), .ZN(
        n11198) );
  NAND2_X1 U14128 ( .A1(n11208), .A2(n11198), .ZN(n11200) );
  INV_X2 U14129 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11223) );
  NAND2_X1 U14130 ( .A1(n11223), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11199) );
  INV_X1 U14131 ( .A(n11206), .ZN(n11201) );
  NAND3_X1 U14132 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n11211), .A3(
        n15903), .ZN(n11978) );
  INV_X1 U14133 ( .A(n11203), .ZN(n11962) );
  INV_X1 U14134 ( .A(n11204), .ZN(n11215) );
  NAND2_X1 U14135 ( .A1(n11962), .A2(n11215), .ZN(n11277) );
  AND2_X1 U14136 ( .A1(n11277), .A2(n11205), .ZN(n11964) );
  XNOR2_X1 U14137 ( .A(n11207), .B(n11206), .ZN(n11976) );
  INV_X1 U14138 ( .A(n11208), .ZN(n11210) );
  MUX2_X1 U14139 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n19946), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11209) );
  XNOR2_X1 U14140 ( .A(n11210), .B(n11209), .ZN(n11970) );
  AND2_X1 U14141 ( .A1(n11976), .A2(n11970), .ZN(n11216) );
  AND3_X1 U14142 ( .A1(n11978), .A2(n11964), .A3(n11216), .ZN(n11213) );
  INV_X1 U14143 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15986) );
  NOR2_X1 U14144 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15986), .ZN(
        n11212) );
  NAND2_X1 U14145 ( .A1(n13761), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11214) );
  NAND2_X1 U14146 ( .A1(n11215), .A2(n11214), .ZN(n11963) );
  INV_X1 U14147 ( .A(n11963), .ZN(n11262) );
  AND3_X1 U14148 ( .A1(n11978), .A2(n11262), .A3(n11216), .ZN(n11217) );
  OAI21_X1 U14149 ( .B1(n16357), .B2(n11217), .A(n11444), .ZN(n11220) );
  AOI21_X1 U14150 ( .B1(n11221), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16364) );
  NAND2_X1 U14151 ( .A1(n14303), .A2(n16364), .ZN(n11219) );
  NOR2_X1 U14152 ( .A1(n11444), .A2(P2_FLUSH_REG_SCAN_IN), .ZN(n11218) );
  NAND2_X1 U14153 ( .A1(n11219), .A2(n11218), .ZN(n19957) );
  AOI22_X1 U14154 ( .A1(n14399), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11229) );
  AOI22_X1 U14155 ( .A1(n11312), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9653), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11227) );
  AND2_X4 U14156 ( .A1(n11222), .A2(n15832), .ZN(n14437) );
  AND2_X4 U14157 ( .A1(n15829), .A2(n11223), .ZN(n11374) );
  AOI22_X1 U14158 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9651), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11226) );
  NOR2_X2 U14159 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11224) );
  NAND2_X2 U14160 ( .A1(n11224), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11317) );
  INV_X2 U14161 ( .A(n11317), .ZN(n11367) );
  AOI22_X1 U14162 ( .A1(n14440), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11225) );
  AOI22_X1 U14163 ( .A1(n11312), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14436), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11233) );
  AOI22_X1 U14164 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14399), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11232) );
  AOI22_X1 U14165 ( .A1(n9651), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9655), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11231) );
  AOI22_X1 U14166 ( .A1(n14440), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11230) );
  NAND2_X1 U14167 ( .A1(n19968), .A2(n19989), .ZN(n11307) );
  AND2_X2 U14168 ( .A1(n11312), .A2(n16338), .ZN(n14287) );
  AOI22_X1 U14169 ( .A1(n11288), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11240) );
  INV_X1 U14170 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19256) );
  NAND2_X2 U14172 ( .A1(n9653), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14289) );
  INV_X1 U14173 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11235) );
  OAI22_X1 U14174 ( .A1(n19256), .A2(n14290), .B1(n14289), .B2(n11235), .ZN(
        n11236) );
  INV_X1 U14175 ( .A(n11236), .ZN(n11239) );
  NAND2_X1 U14176 ( .A1(n11374), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11539) );
  AOI22_X1 U14177 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14293), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11238) );
  AND2_X2 U14178 ( .A1(n14440), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11531) );
  AOI22_X1 U14179 ( .A1(n11531), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11237) );
  NAND4_X1 U14180 ( .A1(n11240), .A2(n11239), .A3(n11238), .A4(n11237), .ZN(
        n11249) );
  AND2_X2 U14181 ( .A1(n14440), .A2(n16338), .ZN(n14299) );
  AOI22_X1 U14182 ( .A1(n14300), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11247) );
  CLKBUF_X3 U14183 ( .A(n14437), .Z(n14417) );
  AND2_X2 U14184 ( .A1(n14417), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11530) );
  OR2_X1 U14185 ( .A1(n11317), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12378) );
  AOI22_X1 U14186 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14301), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11246) );
  INV_X1 U14187 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11242) );
  INV_X1 U14188 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11241) );
  OAI22_X1 U14189 ( .A1(n14305), .A2(n11242), .B1(n14303), .B2(n11241), .ZN(
        n11243) );
  INV_X1 U14190 ( .A(n11243), .ZN(n11245) );
  AOI22_X1 U14191 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14307), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11244) );
  NAND4_X1 U14192 ( .A1(n11247), .A2(n11246), .A3(n11245), .A4(n11244), .ZN(
        n11248) );
  AOI22_X1 U14193 ( .A1(n11312), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14436), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11253) );
  AOI22_X1 U14194 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11374), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11252) );
  AOI22_X1 U14195 ( .A1(n14399), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9637), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11251) );
  AOI22_X1 U14196 ( .A1(n14440), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11250) );
  NAND4_X1 U14197 ( .A1(n11253), .A2(n11252), .A3(n11251), .A4(n11250), .ZN(
        n11254) );
  NAND2_X1 U14198 ( .A1(n11254), .A2(n16338), .ZN(n11261) );
  AOI22_X1 U14199 ( .A1(n11312), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9654), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11258) );
  AOI22_X1 U14200 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9651), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11257) );
  AOI22_X1 U14201 ( .A1(n14440), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11256) );
  AOI22_X1 U14202 ( .A1(n14399), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9657), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11255) );
  NAND4_X1 U14203 ( .A1(n11258), .A2(n11257), .A3(n11256), .A4(n11255), .ZN(
        n11259) );
  MUX2_X1 U14204 ( .A(n12292), .B(n11262), .S(n12811), .Z(n11671) );
  AOI22_X1 U14205 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11288), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11267) );
  INV_X1 U14206 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19264) );
  INV_X1 U14207 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12379) );
  OAI22_X1 U14208 ( .A1(n19264), .A2(n14290), .B1(n14289), .B2(n12379), .ZN(
        n11263) );
  INV_X1 U14209 ( .A(n11263), .ZN(n11266) );
  AOI22_X1 U14210 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14293), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11265) );
  AOI22_X1 U14211 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n11531), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11264) );
  NAND4_X1 U14212 ( .A1(n11267), .A2(n11266), .A3(n11265), .A4(n11264), .ZN(
        n11275) );
  AOI22_X1 U14213 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n14300), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11273) );
  AOI22_X1 U14214 ( .A1(n12466), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12465), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11272) );
  AOI22_X1 U14215 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n14307), .ZN(n11271) );
  INV_X1 U14216 ( .A(n11530), .ZN(n11295) );
  INV_X1 U14217 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13913) );
  INV_X1 U14218 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11268) );
  OAI22_X1 U14219 ( .A1(n11295), .A2(n13913), .B1(n12378), .B2(n11268), .ZN(
        n11269) );
  INV_X1 U14220 ( .A(n11269), .ZN(n11270) );
  NAND4_X1 U14221 ( .A1(n11273), .A2(n11272), .A3(n11271), .A4(n11270), .ZN(
        n11274) );
  INV_X1 U14222 ( .A(n11426), .ZN(n19971) );
  NAND2_X1 U14223 ( .A1(n11547), .A2(n19971), .ZN(n11276) );
  NAND2_X1 U14224 ( .A1(n12811), .A2(n11970), .ZN(n11973) );
  AOI21_X1 U14225 ( .B1(n11671), .B2(n11277), .A(n11650), .ZN(n11304) );
  AOI22_X1 U14226 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11288), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11281) );
  AOI22_X1 U14227 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12459), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11280) );
  AOI22_X1 U14228 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n14293), .B1(
        n14294), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11279) );
  AOI22_X1 U14229 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11531), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11278) );
  NAND4_X1 U14230 ( .A1(n11281), .A2(n11280), .A3(n11279), .A4(n11278), .ZN(
        n11287) );
  AOI22_X1 U14231 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n14307), .ZN(n11285) );
  AOI22_X1 U14232 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n14299), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11284) );
  AOI22_X1 U14233 ( .A1(n12466), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12465), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11283) );
  AOI22_X1 U14234 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14301), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11282) );
  NAND4_X1 U14235 ( .A1(n11285), .A2(n11284), .A3(n11283), .A4(n11282), .ZN(
        n11286) );
  MUX2_X1 U14236 ( .A(n11978), .B(n12324), .S(n19971), .Z(n11655) );
  AOI22_X1 U14237 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11288), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11293) );
  INV_X1 U14238 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19269) );
  INV_X1 U14239 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12395) );
  OAI22_X1 U14240 ( .A1(n19269), .A2(n14290), .B1(n14289), .B2(n12395), .ZN(
        n11289) );
  INV_X1 U14241 ( .A(n11289), .ZN(n11292) );
  AOI22_X1 U14242 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14293), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11291) );
  AOI22_X1 U14243 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n11531), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11290) );
  NAND4_X1 U14244 ( .A1(n11293), .A2(n11292), .A3(n11291), .A4(n11290), .ZN(
        n11302) );
  AOI22_X1 U14245 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n14300), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11300) );
  AOI22_X1 U14246 ( .A1(n12466), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12465), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11299) );
  AOI22_X1 U14247 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n14307), .ZN(n11298) );
  INV_X1 U14248 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13976) );
  INV_X1 U14249 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11294) );
  OAI22_X1 U14250 ( .A1(n11295), .A2(n13976), .B1(n12378), .B2(n11294), .ZN(
        n11296) );
  INV_X1 U14251 ( .A(n11296), .ZN(n11297) );
  NAND4_X1 U14252 ( .A1(n11300), .A2(n11299), .A3(n11298), .A4(n11297), .ZN(
        n11301) );
  MUX2_X1 U14253 ( .A(n12319), .B(n11976), .S(n12811), .Z(n11649) );
  NAND2_X1 U14254 ( .A1(n11655), .A2(n11649), .ZN(n11961) );
  INV_X1 U14255 ( .A(n11984), .ZN(n11303) );
  OAI21_X1 U14256 ( .B1(n11304), .B2(n11961), .A(n11303), .ZN(n19969) );
  AND2_X1 U14257 ( .A1(n11551), .A2(n11388), .ZN(n19970) );
  INV_X1 U14258 ( .A(n19970), .ZN(n12288) );
  NAND2_X1 U14259 ( .A1(n11307), .A2(n11306), .ZN(n11384) );
  AOI22_X1 U14260 ( .A1(n11312), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9654), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11311) );
  AOI22_X1 U14261 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11374), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11310) );
  AOI22_X1 U14262 ( .A1(n14399), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9637), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11309) );
  AOI22_X1 U14263 ( .A1(n14440), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11308) );
  AOI22_X1 U14264 ( .A1(n11312), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14436), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11314) );
  AOI22_X1 U14265 ( .A1(n14440), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11313) );
  AOI22_X1 U14266 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11374), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11316) );
  AOI22_X1 U14267 ( .A1(n9648), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(n9637), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11315) );
  AOI22_X1 U14268 ( .A1(n11312), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9654), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U14269 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11374), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11320) );
  AOI22_X1 U14270 ( .A1(n14399), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9657), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11319) );
  INV_X4 U14271 ( .A(n11317), .ZN(n14272) );
  AOI22_X1 U14272 ( .A1(n14440), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11318) );
  AOI22_X1 U14273 ( .A1(n11312), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14436), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14274 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11374), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14275 ( .A1(n9648), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(n9637), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U14276 ( .A1(n14440), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11323) );
  NAND2_X4 U14277 ( .A1(n11329), .A2(n11328), .ZN(n11413) );
  AOI22_X1 U14278 ( .A1(n11312), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14436), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11334) );
  AOI22_X1 U14279 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9651), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14280 ( .A1(n14399), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9637), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14281 ( .A1(n14440), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11331) );
  NAND4_X1 U14282 ( .A1(n11334), .A2(n11333), .A3(n11332), .A4(n11331), .ZN(
        n11335) );
  AOI22_X1 U14283 ( .A1(n11312), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9654), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11339) );
  AOI22_X1 U14284 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11374), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11338) );
  AOI22_X1 U14285 ( .A1(n14399), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11337) );
  AOI22_X1 U14286 ( .A1(n14440), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11336) );
  NAND4_X1 U14287 ( .A1(n11339), .A2(n11338), .A3(n11337), .A4(n11336), .ZN(
        n11340) );
  NAND2_X1 U14288 ( .A1(n11340), .A2(n16338), .ZN(n11341) );
  AND3_X2 U14289 ( .A1(n11390), .A2(n11413), .A3(n19265), .ZN(n11399) );
  AOI22_X1 U14290 ( .A1(n11312), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14436), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11346) );
  AOI22_X1 U14291 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9651), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11345) );
  AOI22_X1 U14292 ( .A1(n14399), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9655), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11344) );
  AOI22_X1 U14293 ( .A1(n14440), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11343) );
  NAND4_X1 U14294 ( .A1(n11346), .A2(n11345), .A3(n11344), .A4(n11343), .ZN(
        n11347) );
  AOI22_X1 U14295 ( .A1(n11312), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9653), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11351) );
  AOI22_X1 U14296 ( .A1(n14440), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U14297 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11374), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11349) );
  AOI22_X1 U14298 ( .A1(n9648), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9637), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11348) );
  NAND4_X1 U14299 ( .A1(n11351), .A2(n11350), .A3(n11349), .A4(n11348), .ZN(
        n11352) );
  NAND2_X1 U14300 ( .A1(n11352), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11353) );
  AOI22_X1 U14301 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11312), .B1(
        n9654), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14302 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11374), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14303 ( .A1(n14440), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U14304 ( .A1(n9648), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n9657), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11355) );
  NAND4_X1 U14305 ( .A1(n11358), .A2(n11357), .A3(n11356), .A4(n11355), .ZN(
        n11359) );
  NAND2_X1 U14306 ( .A1(n11359), .A2(n16338), .ZN(n11366) );
  AOI22_X1 U14307 ( .A1(n11312), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14436), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14308 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11374), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U14309 ( .A1(n14440), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11361) );
  AOI22_X1 U14310 ( .A1(n14399), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11360) );
  NAND4_X1 U14311 ( .A1(n11363), .A2(n11362), .A3(n11361), .A4(n11360), .ZN(
        n11364) );
  NAND2_X1 U14312 ( .A1(n11364), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11365) );
  AOI22_X1 U14313 ( .A1(n14440), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11367), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U14314 ( .A1(n9648), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9656), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11368) );
  AOI22_X1 U14315 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11374), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11372) );
  AOI22_X1 U14316 ( .A1(n11312), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9653), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11371) );
  NAND3_X1 U14317 ( .A1(n9714), .A2(n11372), .A3(n11371), .ZN(n11380) );
  AOI22_X1 U14318 ( .A1(n9648), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n9655), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11373) );
  AOI22_X1 U14319 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9651), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U14320 ( .A1(n14440), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11377) );
  AOI22_X1 U14321 ( .A1(n11312), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9654), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11376) );
  NAND4_X1 U14322 ( .A1(n10164), .A2(n11378), .A3(n11377), .A4(n11376), .ZN(
        n11379) );
  NAND2_X2 U14323 ( .A1(n11380), .A2(n11379), .ZN(n11417) );
  NOR2_X1 U14324 ( .A1(n13264), .A2(n11417), .ZN(n11381) );
  NAND2_X1 U14326 ( .A1(n11444), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12817) );
  INV_X1 U14327 ( .A(n12817), .ZN(n11382) );
  NAND2_X1 U14328 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n11382), .ZN(n19845) );
  NOR2_X1 U14329 ( .A1(n11397), .A2(n19845), .ZN(n11383) );
  AND2_X1 U14330 ( .A1(n12283), .A2(n19971), .ZN(n16297) );
  INV_X1 U14331 ( .A(n16297), .ZN(n11993) );
  NAND2_X1 U14332 ( .A1(n9634), .A2(n11387), .ZN(n11386) );
  NAND2_X1 U14333 ( .A1(n12969), .A2(n11417), .ZN(n11385) );
  NAND2_X1 U14334 ( .A1(n11455), .A2(n16366), .ZN(n11396) );
  NAND2_X1 U14335 ( .A1(n11420), .A2(n11413), .ZN(n11394) );
  INV_X2 U14336 ( .A(n11417), .ZN(n11389) );
  NAND4_X1 U14337 ( .A1(n11391), .A2(n11418), .A3(n11390), .A4(n11389), .ZN(
        n11392) );
  NOR2_X2 U14338 ( .A1(n11392), .A2(n13264), .ZN(n11410) );
  NOR2_X1 U14339 ( .A1(n11410), .A2(n11388), .ZN(n11393) );
  NAND2_X1 U14340 ( .A1(n11396), .A2(n12519), .ZN(n11404) );
  NAND3_X1 U14341 ( .A1(n11397), .A2(n11413), .A3(n19989), .ZN(n11402) );
  NAND2_X1 U14342 ( .A1(n11398), .A2(n11417), .ZN(n12295) );
  AND2_X2 U14343 ( .A1(n11400), .A2(n11399), .ZN(n11428) );
  INV_X1 U14344 ( .A(n11428), .ZN(n11401) );
  NAND2_X1 U14345 ( .A1(n11402), .A2(n11401), .ZN(n12508) );
  NAND2_X1 U14346 ( .A1(n11388), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19986) );
  NOR2_X1 U14347 ( .A1(n12508), .A2(n19986), .ZN(n11403) );
  AOI21_X2 U14348 ( .B1(n11404), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11403), 
        .ZN(n11452) );
  INV_X1 U14349 ( .A(n12266), .ZN(n12290) );
  INV_X1 U14350 ( .A(n12271), .ZN(n11405) );
  NAND2_X1 U14351 ( .A1(n11406), .A2(n11418), .ZN(n11407) );
  NAND2_X1 U14352 ( .A1(n11454), .A2(n11429), .ZN(n11408) );
  NAND2_X1 U14353 ( .A1(n19987), .A2(n11444), .ZN(n19979) );
  NOR2_X1 U14354 ( .A1(n19979), .A2(n19938), .ZN(n11409) );
  AOI21_X1 U14355 ( .B1(n11466), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11409), .ZN(n11435) );
  NAND2_X1 U14356 ( .A1(n11428), .A2(n11388), .ZN(n11411) );
  NAND2_X1 U14357 ( .A1(n11410), .A2(n16366), .ZN(n12264) );
  AND2_X2 U14358 ( .A1(n11411), .A2(n12264), .ZN(n12509) );
  NAND2_X1 U14359 ( .A1(n16366), .A2(n11412), .ZN(n11416) );
  INV_X1 U14360 ( .A(n11416), .ZN(n11966) );
  INV_X1 U14361 ( .A(n13264), .ZN(n11414) );
  NAND3_X1 U14362 ( .A1(n12514), .A2(n19275), .A3(n11414), .ZN(n11415) );
  NAND2_X1 U14363 ( .A1(n11449), .A2(n11551), .ZN(n11424) );
  NAND3_X1 U14364 ( .A1(n12515), .A2(n19288), .A3(n11387), .ZN(n11423) );
  NOR2_X2 U14365 ( .A1(n11423), .A2(n11422), .ZN(n12507) );
  NAND2_X1 U14366 ( .A1(n12507), .A2(n12525), .ZN(n15828) );
  INV_X1 U14367 ( .A(n12525), .ZN(n11425) );
  INV_X1 U14368 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n11430) );
  INV_X1 U14369 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12785) );
  OAI22_X1 U14370 ( .A1(n11858), .A2(n11430), .B1(n11444), .B2(n12785), .ZN(
        n11431) );
  AOI21_X1 U14371 ( .B1(n11463), .B2(P2_EBX_REG_3__SCAN_IN), .A(n11431), .ZN(
        n11432) );
  NAND2_X1 U14372 ( .A1(n11433), .A2(n11432), .ZN(n11436) );
  INV_X1 U14373 ( .A(n11436), .ZN(n11434) );
  INV_X1 U14374 ( .A(n11435), .ZN(n11437) );
  NAND2_X1 U14375 ( .A1(n11466), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11439) );
  AOI21_X1 U14376 ( .B1(n19987), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11438) );
  INV_X1 U14377 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13141) );
  INV_X1 U14378 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n11440) );
  INV_X1 U14379 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14464) );
  OAI22_X1 U14380 ( .A1(n11858), .A2(n11440), .B1(n11444), .B2(n14464), .ZN(
        n11441) );
  AOI21_X1 U14381 ( .B1(n11463), .B2(P2_EBX_REG_2__SCAN_IN), .A(n11441), .ZN(
        n11442) );
  INV_X1 U14382 ( .A(n11856), .ZN(n11443) );
  NAND2_X1 U14383 ( .A1(n11443), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11448) );
  INV_X1 U14384 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n11445) );
  OAI22_X1 U14385 ( .A1(n11858), .A2(n11445), .B1(n11444), .B2(n13808), .ZN(
        n11446) );
  AOI21_X1 U14386 ( .B1(n11463), .B2(P2_EBX_REG_1__SCAN_IN), .A(n11446), .ZN(
        n11447) );
  AND2_X2 U14387 ( .A1(n11448), .A2(n11447), .ZN(n11475) );
  NAND2_X1 U14388 ( .A1(n13762), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11450) );
  OAI21_X1 U14389 ( .B1(n19956), .B2(n19979), .A(n11450), .ZN(n11451) );
  AOI21_X2 U14390 ( .B1(n11466), .B2(n15832), .A(n11451), .ZN(n11470) );
  INV_X1 U14391 ( .A(n11470), .ZN(n11476) );
  INV_X1 U14392 ( .A(n11856), .ZN(n11453) );
  NAND2_X1 U14393 ( .A1(n11453), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11461) );
  INV_X1 U14394 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n11457) );
  NAND2_X1 U14395 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11456) );
  OAI211_X1 U14396 ( .C1(n11858), .C2(n11457), .A(n19979), .B(n11456), .ZN(
        n11458) );
  AOI21_X1 U14397 ( .B1(n11463), .B2(P2_EBX_REG_0__SCAN_IN), .A(n11458), .ZN(
        n11459) );
  NAND2_X1 U14398 ( .A1(n12525), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11462) );
  NOR2_X1 U14399 ( .A1(n11462), .A2(n12811), .ZN(n11465) );
  OAI21_X1 U14400 ( .B1(n11466), .B2(n11465), .A(n11464), .ZN(n11469) );
  OAI22_X1 U14401 ( .A1(n15828), .A2(n19987), .B1(n19966), .B2(n19979), .ZN(
        n11467) );
  INV_X1 U14402 ( .A(n11467), .ZN(n11468) );
  NAND2_X1 U14403 ( .A1(n11469), .A2(n11468), .ZN(n11472) );
  NAND2_X2 U14404 ( .A1(n11475), .A2(n11470), .ZN(n11486) );
  OR2_X1 U14405 ( .A1(n11472), .A2(n11471), .ZN(n11473) );
  BUF_X2 U14406 ( .A(n11474), .Z(n11494) );
  XNOR2_X2 U14407 ( .A(n11494), .B(n11485), .ZN(n11496) );
  NAND2_X1 U14408 ( .A1(n11486), .A2(n11482), .ZN(n11479) );
  INV_X1 U14409 ( .A(n11475), .ZN(n11477) );
  NAND2_X1 U14410 ( .A1(n11477), .A2(n11476), .ZN(n11484) );
  NAND2_X1 U14411 ( .A1(n11484), .A2(n11849), .ZN(n11478) );
  NAND2_X1 U14412 ( .A1(n11484), .A2(n11482), .ZN(n11481) );
  NAND2_X1 U14413 ( .A1(n11486), .A2(n11849), .ZN(n11480) );
  AOI21_X2 U14414 ( .B1(n11481), .B2(n11480), .A(n11483), .ZN(n11492) );
  NAND3_X1 U14415 ( .A1(n11488), .A2(n11485), .A3(n11484), .ZN(n11491) );
  INV_X1 U14416 ( .A(n11485), .ZN(n11487) );
  NAND2_X1 U14417 ( .A1(n11487), .A2(n11486), .ZN(n11489) );
  OR2_X2 U14418 ( .A1(n11489), .A2(n11488), .ZN(n11490) );
  OAI211_X4 U14419 ( .C1(n11493), .C2(n11492), .A(n11491), .B(n11490), .ZN(
        n13115) );
  AND2_X2 U14420 ( .A1(n11501), .A2(n11497), .ZN(n19250) );
  INV_X1 U14421 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19259) );
  AND2_X1 U14422 ( .A1(n11494), .A2(n15823), .ZN(n11509) );
  INV_X1 U14423 ( .A(n19771), .ZN(n11495) );
  INV_X1 U14424 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12360) );
  INV_X1 U14425 ( .A(n11498), .ZN(n11499) );
  NOR2_X1 U14426 ( .A1(n11500), .A2(n11499), .ZN(n11528) );
  AND2_X2 U14427 ( .A1(n11501), .A2(n13680), .ZN(n11503) );
  AND2_X2 U14428 ( .A1(n11503), .A2(n11502), .ZN(n11572) );
  AOI22_X1 U14429 ( .A1(n11572), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11557), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11506) );
  AND2_X2 U14430 ( .A1(n11503), .A2(n11496), .ZN(n11562) );
  AND2_X1 U14431 ( .A1(n11506), .A2(n11505), .ZN(n11527) );
  NAND2_X1 U14432 ( .A1(n13115), .A2(n11509), .ZN(n11507) );
  NAND2_X1 U14433 ( .A1(n11566), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11514) );
  NAND2_X1 U14434 ( .A1(n11553), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11513) );
  INV_X1 U14435 ( .A(n11509), .ZN(n11510) );
  NOR2_X1 U14436 ( .A1(n13115), .A2(n11510), .ZN(n11511) );
  NAND2_X1 U14437 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11512) );
  INV_X1 U14438 ( .A(n11494), .ZN(n11515) );
  INV_X1 U14439 ( .A(n11520), .ZN(n11516) );
  NOR2_X1 U14440 ( .A1(n13115), .A2(n11516), .ZN(n11517) );
  NAND2_X1 U14441 ( .A1(n13115), .A2(n11520), .ZN(n11518) );
  NOR2_X1 U14442 ( .A1(n11518), .A2(n15859), .ZN(n11568) );
  AOI22_X1 U14443 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11565), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11524) );
  NAND2_X1 U14444 ( .A1(n19613), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11523) );
  AOI22_X1 U14445 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n11555), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11522) );
  INV_X1 U14446 ( .A(n12292), .ZN(n13072) );
  AOI22_X1 U14447 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n14293), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11529) );
  OAI21_X1 U14448 ( .B1(n19259), .B2(n14290), .A(n11529), .ZN(n11537) );
  AOI22_X1 U14449 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12466), .B1(
        n14308), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U14450 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n12465), .B1(
        n11288), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11534) );
  AOI22_X1 U14451 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14452 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n14287), .B1(
        n11531), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11532) );
  NAND4_X1 U14453 ( .A1(n11535), .A2(n11534), .A3(n11533), .A4(n11532), .ZN(
        n11536) );
  AOI211_X1 U14454 ( .C1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .C2(n14307), .A(
        n11537), .B(n11536), .ZN(n11545) );
  INV_X1 U14455 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11538) );
  OAI22_X1 U14456 ( .A1(n12360), .A2(n14289), .B1(n11539), .B2(n11538), .ZN(
        n11543) );
  INV_X1 U14457 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11541) );
  INV_X1 U14458 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11540) );
  OAI22_X1 U14459 ( .A1(n11541), .A2(n12408), .B1(n12378), .B2(n11540), .ZN(
        n11542) );
  NOR2_X1 U14460 ( .A1(n11543), .A2(n11542), .ZN(n11544) );
  NOR2_X1 U14461 ( .A1(n13072), .A2(n12302), .ZN(n11546) );
  NAND2_X1 U14462 ( .A1(n11551), .A2(n11546), .ZN(n11803) );
  NAND2_X1 U14463 ( .A1(n11803), .A2(n12311), .ZN(n11548) );
  AOI22_X1 U14464 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n11566), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11550) );
  INV_X1 U14465 ( .A(n14355), .ZN(n11551) );
  NAND2_X1 U14466 ( .A1(n12319), .A2(n11551), .ZN(n11552) );
  INV_X1 U14467 ( .A(n11660), .ZN(n11588) );
  AOI22_X1 U14468 ( .A1(n19338), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11553), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U14469 ( .A1(n19250), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11554), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11560) );
  AOI22_X1 U14470 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n11555), .B1(
        n11556), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11559) );
  NAND2_X1 U14471 ( .A1(n11557), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11558) );
  AOI22_X1 U14472 ( .A1(n11562), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U14473 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19771), .B1(
        n19613), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11571) );
  AOI22_X1 U14474 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n11565), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14475 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n11567), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11569) );
  AND3_X1 U14476 ( .A1(n11571), .A2(n11570), .A3(n11569), .ZN(n11574) );
  NAND2_X1 U14477 ( .A1(n11572), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11573) );
  AOI22_X1 U14478 ( .A1(n11288), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14479 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12459), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14480 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14293), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U14481 ( .A1(n14301), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11576) );
  NAND4_X1 U14482 ( .A1(n11579), .A2(n11578), .A3(n11577), .A4(n11576), .ZN(
        n11585) );
  AOI22_X1 U14483 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11531), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14484 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14485 ( .A1(n12466), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11581) );
  AOI22_X1 U14486 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14307), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11580) );
  NAND4_X1 U14487 ( .A1(n11583), .A2(n11582), .A3(n11581), .A4(n11580), .ZN(
        n11584) );
  INV_X1 U14488 ( .A(n11656), .ZN(n11586) );
  NAND2_X1 U14489 ( .A1(n11586), .A2(n11551), .ZN(n11587) );
  NAND2_X1 U14490 ( .A1(n11572), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11592) );
  AOI22_X1 U14491 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11566), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11591) );
  AOI22_X1 U14492 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11567), .B1(
        n11565), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11590) );
  AOI22_X1 U14493 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19771), .B1(
        n19613), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11589) );
  INV_X1 U14494 ( .A(n19338), .ZN(n11595) );
  INV_X1 U14495 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14254) );
  INV_X1 U14496 ( .A(n11554), .ZN(n11594) );
  INV_X1 U14497 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11593) );
  OAI22_X1 U14498 ( .A1(n11595), .A2(n14254), .B1(n11594), .B2(n11593), .ZN(
        n11600) );
  INV_X1 U14499 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11598) );
  INV_X1 U14500 ( .A(n11556), .ZN(n19550) );
  INV_X1 U14501 ( .A(n11555), .ZN(n11597) );
  INV_X1 U14502 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11596) );
  OAI22_X1 U14503 ( .A1(n11598), .A2(n19550), .B1(n11597), .B2(n11596), .ZN(
        n11599) );
  NOR2_X1 U14504 ( .A1(n11600), .A2(n11599), .ZN(n11605) );
  INV_X1 U14505 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19286) );
  INV_X1 U14506 ( .A(n11553), .ZN(n11601) );
  INV_X1 U14507 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12448) );
  OAI22_X1 U14508 ( .A1(n19245), .A2(n19286), .B1(n11601), .B2(n12448), .ZN(
        n11602) );
  AOI21_X1 U14509 ( .B1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n11562), .A(
        n11602), .ZN(n11604) );
  AOI22_X1 U14510 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n11557), .B1(
        n11564), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11603) );
  NAND4_X1 U14511 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(
        n11618) );
  AOI22_X1 U14512 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n14293), .B1(
        n14294), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U14513 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11288), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U14514 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12459), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11608) );
  AOI22_X1 U14515 ( .A1(n12466), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11531), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11607) );
  NAND4_X1 U14516 ( .A1(n11610), .A2(n11609), .A3(n11608), .A4(n11607), .ZN(
        n11616) );
  AOI22_X1 U14517 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14308), .B1(
        n11530), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11614) );
  AOI22_X1 U14518 ( .A1(n14300), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n14307), .ZN(n11613) );
  AOI22_X1 U14519 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n12465), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11612) );
  AOI22_X1 U14520 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n14299), .B1(
        n14301), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11611) );
  NAND4_X1 U14521 ( .A1(n11614), .A2(n11613), .A3(n11612), .A4(n11611), .ZN(
        n11615) );
  NAND2_X1 U14522 ( .A1(n11647), .A2(n11551), .ZN(n11617) );
  INV_X1 U14523 ( .A(n11816), .ZN(n11619) );
  NAND2_X1 U14524 ( .A1(n11620), .A2(n11816), .ZN(n11621) );
  INV_X1 U14525 ( .A(n14308), .ZN(n11624) );
  INV_X1 U14526 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11623) );
  INV_X1 U14527 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11622) );
  OAI22_X1 U14528 ( .A1(n11624), .A2(n11623), .B1(n12378), .B2(n11622), .ZN(
        n11630) );
  INV_X1 U14529 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11628) );
  INV_X1 U14530 ( .A(n11625), .ZN(n11627) );
  INV_X1 U14531 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11626) );
  OAI22_X1 U14532 ( .A1(n11628), .A2(n12408), .B1(n11627), .B2(n11626), .ZN(
        n11629) );
  NOR2_X1 U14533 ( .A1(n11630), .A2(n11629), .ZN(n11646) );
  NAND2_X1 U14534 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11634) );
  NAND2_X1 U14535 ( .A1(n11288), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11633) );
  NAND2_X1 U14536 ( .A1(n12459), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11632) );
  NAND2_X1 U14537 ( .A1(n14287), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11631) );
  NAND2_X1 U14538 ( .A1(n12466), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11638) );
  NAND2_X1 U14539 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11637) );
  NAND2_X1 U14540 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n14307), .ZN(
        n11636) );
  NAND2_X1 U14541 ( .A1(n14299), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11635) );
  NAND2_X1 U14542 ( .A1(n14293), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11642) );
  NAND2_X1 U14543 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11641) );
  NAND2_X1 U14544 ( .A1(n11531), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11640) );
  NAND2_X1 U14545 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11639) );
  NAND4_X1 U14546 ( .A1(n11646), .A2(n11645), .A3(n11644), .A4(n11643), .ZN(
        n11683) );
  MUX2_X1 U14547 ( .A(n11647), .B(P2_EBX_REG_6__SCAN_IN), .S(n19275), .Z(
        n11658) );
  INV_X1 U14548 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n11648) );
  MUX2_X1 U14549 ( .A(n11649), .B(n11648), .S(n19275), .Z(n11668) );
  INV_X1 U14550 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n14219) );
  MUX2_X1 U14551 ( .A(n14219), .B(n11650), .S(n9632), .Z(n11667) );
  NAND2_X1 U14552 ( .A1(n11668), .A2(n11667), .ZN(n11653) );
  INV_X1 U14553 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n11651) );
  INV_X1 U14554 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13044) );
  NAND2_X1 U14555 ( .A1(n11651), .A2(n13044), .ZN(n11652) );
  MUX2_X2 U14556 ( .A(n11652), .B(n12302), .S(n9632), .Z(n11673) );
  INV_X1 U14557 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n11654) );
  MUX2_X1 U14558 ( .A(n11655), .B(n11654), .S(n19275), .Z(n11677) );
  NAND2_X1 U14559 ( .A1(n9632), .A2(n11656), .ZN(n12328) );
  INV_X1 U14560 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13206) );
  NAND2_X1 U14561 ( .A1(n19275), .A2(n13206), .ZN(n11657) );
  AOI21_X1 U14562 ( .B1(n11658), .B2(n11661), .A(n11691), .ZN(n19098) );
  XNOR2_X1 U14563 ( .A(n11681), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13928) );
  INV_X1 U14564 ( .A(n11661), .ZN(n11662) );
  AOI21_X1 U14565 ( .B1(n11664), .B2(n11663), .A(n11662), .ZN(n19114) );
  INV_X1 U14566 ( .A(n11667), .ZN(n11670) );
  NOR2_X1 U14567 ( .A1(n11673), .A2(n11670), .ZN(n11669) );
  OAI21_X1 U14568 ( .B1(n11669), .B2(n11668), .A(n9946), .ZN(n13543) );
  OAI21_X2 U14569 ( .B1(n13487), .B2(n11790), .A(n13543), .ZN(n13484) );
  XNOR2_X1 U14570 ( .A(n11673), .B(n11670), .ZN(n13677) );
  MUX2_X1 U14571 ( .A(n11671), .B(P2_EBX_REG_0__SCAN_IN), .S(n19275), .Z(
        n19130) );
  NAND2_X1 U14572 ( .A1(n19130), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13070) );
  NAND3_X1 U14573 ( .A1(n19275), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n11672) );
  NAND2_X1 U14574 ( .A1(n11673), .A2(n11672), .ZN(n13807) );
  NOR2_X1 U14575 ( .A1(n13070), .A2(n13807), .ZN(n11674) );
  NAND2_X1 U14576 ( .A1(n13070), .A2(n13807), .ZN(n13046) );
  OAI21_X1 U14577 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n11674), .A(
        n13046), .ZN(n13152) );
  XNOR2_X1 U14578 ( .A(n13677), .B(n13141), .ZN(n13151) );
  OR2_X1 U14579 ( .A1(n13152), .A2(n13151), .ZN(n14466) );
  OAI21_X1 U14580 ( .B1(n13677), .B2(n13141), .A(n14466), .ZN(n13485) );
  INV_X1 U14581 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13500) );
  NAND2_X1 U14582 ( .A1(n13484), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11675) );
  NAND2_X1 U14583 ( .A1(n11676), .A2(n11675), .ZN(n13595) );
  XNOR2_X1 U14584 ( .A(n11678), .B(n11677), .ZN(n13563) );
  XNOR2_X1 U14585 ( .A(n13563), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13596) );
  INV_X1 U14586 ( .A(n13563), .ZN(n11679) );
  INV_X1 U14587 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13789) );
  INV_X1 U14588 ( .A(n11681), .ZN(n11682) );
  INV_X1 U14589 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13273) );
  MUX2_X1 U14590 ( .A(n11683), .B(n13273), .S(n19275), .Z(n11689) );
  INV_X1 U14591 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n13353) );
  NAND2_X1 U14592 ( .A1(n11687), .A2(n13353), .ZN(n11685) );
  NAND2_X1 U14593 ( .A1(n19275), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11686) );
  NOR2_X1 U14594 ( .A1(n11687), .A2(n11686), .ZN(n11688) );
  OR2_X1 U14595 ( .A1(n11695), .A2(n11688), .ZN(n13594) );
  NAND2_X1 U14596 ( .A1(n11790), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11826) );
  NOR2_X1 U14597 ( .A1(n13594), .A2(n11826), .ZN(n16280) );
  INV_X1 U14598 ( .A(n11689), .ZN(n11690) );
  XNOR2_X1 U14599 ( .A(n11691), .B(n11690), .ZN(n13607) );
  NOR2_X1 U14600 ( .A1(n16280), .A2(n16278), .ZN(n11693) );
  INV_X1 U14601 ( .A(n13594), .ZN(n11692) );
  AOI21_X1 U14602 ( .B1(n11692), .B2(n11790), .A(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16281) );
  NOR2_X1 U14603 ( .A1(n13607), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13944) );
  AND2_X1 U14604 ( .A1(n19275), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11694) );
  XNOR2_X1 U14605 ( .A(n11695), .B(n11694), .ZN(n19090) );
  NAND2_X1 U14606 ( .A1(n19090), .A2(n11790), .ZN(n11700) );
  INV_X1 U14607 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15810) );
  NAND2_X1 U14608 ( .A1(n11700), .A2(n15810), .ZN(n15551) );
  INV_X1 U14609 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n13360) );
  INV_X1 U14610 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13519) );
  INV_X1 U14611 ( .A(n11792), .ZN(n11699) );
  NAND2_X1 U14612 ( .A1(n19275), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11696) );
  NOR2_X1 U14613 ( .A1(n11697), .A2(n11696), .ZN(n11698) );
  OR3_X1 U14614 ( .A1(n11706), .A2(n11699), .A3(n11698), .ZN(n13582) );
  INV_X1 U14615 ( .A(n13582), .ZN(n11702) );
  AOI21_X1 U14616 ( .B1(n11702), .B2(n11790), .A(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16269) );
  AND2_X1 U14617 ( .A1(n11790), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11701) );
  INV_X1 U14618 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11704) );
  INV_X1 U14619 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n11705) );
  OR3_X1 U14620 ( .A1(n11706), .A2(n11705), .A3(n9632), .ZN(n11708) );
  INV_X1 U14621 ( .A(n11710), .ZN(n11707) );
  NAND2_X1 U14622 ( .A1(n11708), .A2(n11707), .ZN(n19079) );
  NOR2_X1 U14623 ( .A1(n19079), .A2(n15461), .ZN(n15795) );
  NAND2_X1 U14624 ( .A1(n19275), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11709) );
  AND2_X1 U14625 ( .A1(n19275), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11711) );
  OR2_X2 U14626 ( .A1(n11726), .A2(n11711), .ZN(n11729) );
  AND2_X1 U14627 ( .A1(n19275), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11728) );
  NAND2_X2 U14628 ( .A1(n11713), .A2(n11712), .ZN(n11731) );
  INV_X1 U14629 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n11717) );
  INV_X1 U14630 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11714) );
  NAND2_X1 U14631 ( .A1(n11717), .A2(n11714), .ZN(n11715) );
  AND2_X1 U14632 ( .A1(n19275), .A2(n11715), .ZN(n11716) );
  NOR2_X4 U14633 ( .A1(n11731), .A2(n11716), .ZN(n11741) );
  INV_X1 U14634 ( .A(n11741), .ZN(n11720) );
  INV_X1 U14635 ( .A(n11731), .ZN(n11718) );
  NAND2_X1 U14636 ( .A1(n11718), .A2(n11717), .ZN(n11722) );
  NAND3_X1 U14637 ( .A1(n11722), .A2(P2_EBX_REG_19__SCAN_IN), .A3(n19275), 
        .ZN(n11719) );
  NAND2_X1 U14638 ( .A1(n11720), .A2(n11719), .ZN(n19006) );
  INV_X1 U14639 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15684) );
  NAND2_X1 U14640 ( .A1(n11747), .A2(n15684), .ZN(n15492) );
  NAND2_X1 U14641 ( .A1(n11731), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11721) );
  MUX2_X1 U14642 ( .A(n11721), .B(n11731), .S(n9632), .Z(n11723) );
  NAND2_X1 U14643 ( .A1(n11723), .A2(n11722), .ZN(n15227) );
  INV_X1 U14644 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15696) );
  OAI21_X1 U14645 ( .B1(n15227), .B2(n15461), .A(n15696), .ZN(n15493) );
  AND2_X1 U14646 ( .A1(n15492), .A2(n15493), .ZN(n15478) );
  AND2_X1 U14647 ( .A1(n19275), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11724) );
  XNOR2_X1 U14648 ( .A(n11741), .B(n11724), .ZN(n18987) );
  NAND2_X1 U14649 ( .A1(n18987), .A2(n11790), .ZN(n11753) );
  INV_X1 U14650 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15673) );
  NAND2_X1 U14651 ( .A1(n11753), .A2(n15673), .ZN(n15481) );
  AND2_X1 U14652 ( .A1(n15478), .A2(n15481), .ZN(n15467) );
  NAND3_X1 U14653 ( .A1(n11726), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n19275), 
        .ZN(n11725) );
  OAI211_X1 U14654 ( .C1(n11726), .C2(P2_EBX_REG_16__SCAN_IN), .A(n11725), .B(
        n11792), .ZN(n19025) );
  OR2_X1 U14655 ( .A1(n19025), .A2(n15461), .ZN(n11727) );
  XNOR2_X1 U14656 ( .A(n11727), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15528) );
  NAND2_X1 U14657 ( .A1(n11729), .A2(n11728), .ZN(n11730) );
  NAND2_X1 U14658 ( .A1(n19021), .A2(n11790), .ZN(n11748) );
  INV_X1 U14659 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15508) );
  AND2_X1 U14660 ( .A1(n11748), .A2(n15508), .ZN(n15518) );
  XNOR2_X1 U14661 ( .A(n11732), .B(n9751), .ZN(n12855) );
  AOI21_X1 U14662 ( .B1(n12855), .B2(n11790), .A(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15538) );
  XNOR2_X1 U14663 ( .A(n11733), .B(n9742), .ZN(n19040) );
  AOI21_X1 U14664 ( .B1(n19040), .B2(n11790), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15463) );
  XNOR2_X1 U14665 ( .A(n11734), .B(n10172), .ZN(n19053) );
  NAND2_X1 U14666 ( .A1(n19053), .A2(n11790), .ZN(n11735) );
  INV_X1 U14667 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15769) );
  NAND2_X1 U14668 ( .A1(n11735), .A2(n15769), .ZN(n15761) );
  NAND3_X1 U14669 ( .A1(n19275), .A2(P2_EBX_REG_12__SCAN_IN), .A3(n11736), 
        .ZN(n11737) );
  NAND2_X1 U14670 ( .A1(n11734), .A2(n11737), .ZN(n19064) );
  OR2_X1 U14671 ( .A1(n19064), .A2(n15461), .ZN(n11738) );
  NAND2_X1 U14672 ( .A1(n11738), .A2(n11704), .ZN(n15777) );
  NAND2_X1 U14673 ( .A1(n15761), .A2(n15777), .ZN(n11739) );
  NOR4_X1 U14674 ( .A1(n15518), .A2(n15538), .A3(n15463), .A4(n11739), .ZN(
        n11745) );
  INV_X1 U14675 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n11740) );
  NAND3_X1 U14676 ( .A1(n11743), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n19275), 
        .ZN(n11742) );
  AND2_X1 U14677 ( .A1(n11742), .A2(n11792), .ZN(n11744) );
  INV_X1 U14678 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15473) );
  OAI21_X1 U14679 ( .B1(n18976), .B2(n15461), .A(n15473), .ZN(n15468) );
  NAND4_X1 U14680 ( .A1(n15467), .A2(n15528), .A3(n11745), .A4(n15468), .ZN(
        n11746) );
  INV_X1 U14681 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15721) );
  OR3_X1 U14682 ( .A1(n19025), .A2(n15461), .A3(n15721), .ZN(n15464) );
  INV_X1 U14683 ( .A(n12855), .ZN(n11749) );
  INV_X1 U14684 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15543) );
  INV_X1 U14685 ( .A(n19053), .ZN(n11750) );
  AND2_X1 U14686 ( .A1(n11790), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11751) );
  NAND2_X1 U14687 ( .A1(n19040), .A2(n11751), .ZN(n15741) );
  NAND4_X1 U14688 ( .A1(n15464), .A2(n15539), .A3(n15760), .A4(n15741), .ZN(
        n11752) );
  INV_X1 U14689 ( .A(n11753), .ZN(n11754) );
  NAND2_X1 U14690 ( .A1(n11790), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11755) );
  AND2_X1 U14691 ( .A1(n19275), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11758) );
  AOI21_X2 U14692 ( .B1(n11757), .B2(n11792), .A(n11758), .ZN(n11760) );
  AOI21_X1 U14693 ( .B1(n11758), .B2(n11757), .A(n11760), .ZN(n12892) );
  AOI21_X1 U14694 ( .B1(n12892), .B2(n11790), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15451) );
  NAND3_X1 U14695 ( .A1(n12892), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n11790), .ZN(n15449) );
  NAND2_X1 U14696 ( .A1(n19275), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11759) );
  AND2_X2 U14697 ( .A1(n11760), .A2(n11759), .ZN(n11766) );
  NOR2_X1 U14698 ( .A1(n11760), .A2(n11759), .ZN(n11761) );
  OR2_X1 U14699 ( .A1(n11766), .A2(n11761), .ZN(n12869) );
  XNOR2_X1 U14700 ( .A(n11762), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15439) );
  INV_X1 U14701 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15633) );
  NAND2_X1 U14702 ( .A1(n19275), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11763) );
  MUX2_X1 U14703 ( .A(n11763), .B(P2_EBX_REG_24__SCAN_IN), .S(n11766), .Z(
        n11764) );
  NAND2_X1 U14704 ( .A1(n11764), .A2(n11792), .ZN(n16216) );
  NOR2_X1 U14705 ( .A1(n16216), .A2(n15461), .ZN(n15429) );
  INV_X1 U14706 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15619) );
  NAND2_X1 U14707 ( .A1(n11792), .A2(n11790), .ZN(n11782) );
  INV_X1 U14708 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15607) );
  NAND2_X1 U14709 ( .A1(n11782), .A2(n15607), .ZN(n15417) );
  INV_X1 U14710 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n15270) );
  OR2_X2 U14711 ( .A1(n15208), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11768) );
  AND2_X1 U14712 ( .A1(n19275), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11767) );
  AOI21_X1 U14713 ( .B1(n11768), .B2(n11767), .A(n11770), .ZN(n16205) );
  AND2_X1 U14714 ( .A1(n16205), .A2(n11790), .ZN(n11769) );
  NAND3_X1 U14715 ( .A1(n16205), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n11790), .ZN(n11783) );
  OAI21_X1 U14716 ( .B1(n11769), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11783), .ZN(n15408) );
  NAND2_X1 U14717 ( .A1(n19275), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11771) );
  INV_X1 U14718 ( .A(n11771), .ZN(n11772) );
  NAND2_X1 U14719 ( .A1(n11772), .A2(n9707), .ZN(n11773) );
  NAND2_X1 U14720 ( .A1(n11775), .A2(n11773), .ZN(n12880) );
  INV_X1 U14721 ( .A(n11775), .ZN(n11777) );
  AND2_X1 U14722 ( .A1(n19275), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11774) );
  INV_X1 U14723 ( .A(n11774), .ZN(n11776) );
  OAI21_X1 U14724 ( .B1(n11777), .B2(n11776), .A(n11786), .ZN(n15199) );
  NOR2_X2 U14725 ( .A1(n15199), .A2(n15461), .ZN(n14196) );
  OAI21_X1 U14726 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n14196), .ZN(n11778) );
  INV_X1 U14727 ( .A(n14196), .ZN(n11779) );
  INV_X1 U14728 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15564) );
  NAND2_X1 U14729 ( .A1(n11779), .A2(n15564), .ZN(n11780) );
  OR2_X1 U14730 ( .A1(n11782), .A2(n15607), .ZN(n15418) );
  NAND2_X1 U14731 ( .A1(n19275), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11784) );
  XOR2_X1 U14732 ( .A(n11784), .B(n11786), .Z(n11789) );
  INV_X1 U14733 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12287) );
  OAI21_X1 U14734 ( .B1(n11789), .B2(n15461), .A(n12287), .ZN(n12260) );
  INV_X1 U14735 ( .A(n11784), .ZN(n11785) );
  NAND2_X1 U14736 ( .A1(n19275), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11787) );
  XNOR2_X1 U14737 ( .A(n11791), .B(n11787), .ZN(n12813) );
  AOI21_X1 U14738 ( .B1(n12813), .B2(n11790), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14185) );
  AND2_X1 U14739 ( .A1(n11790), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11788) );
  NAND2_X1 U14740 ( .A1(n12813), .A2(n11788), .ZN(n14183) );
  INV_X1 U14741 ( .A(n11789), .ZN(n16197) );
  NAND3_X1 U14742 ( .A1(n16197), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11790), .ZN(n14181) );
  OAI21_X1 U14743 ( .B1(n11791), .B2(P2_EBX_REG_30__SCAN_IN), .A(n19275), .ZN(
        n11793) );
  NAND2_X1 U14744 ( .A1(n11793), .A2(n11792), .ZN(n16183) );
  NOR2_X1 U14745 ( .A1(n16183), .A2(n15461), .ZN(n11794) );
  XOR2_X1 U14746 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11794), .Z(
        n11795) );
  XNOR2_X1 U14747 ( .A(n11796), .B(n11795), .ZN(n14180) );
  NAND2_X1 U14748 ( .A1(n11797), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13778) );
  NAND2_X1 U14749 ( .A1(n13072), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13071) );
  INV_X1 U14750 ( .A(n13071), .ZN(n11799) );
  INV_X1 U14751 ( .A(n12302), .ZN(n11798) );
  NAND2_X1 U14752 ( .A1(n11799), .A2(n11798), .ZN(n11802) );
  NOR2_X1 U14753 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n12292), .ZN(
        n11800) );
  XNOR2_X1 U14754 ( .A(n11798), .B(n11800), .ZN(n13048) );
  NAND2_X1 U14755 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13048), .ZN(
        n11801) );
  NAND2_X1 U14756 ( .A1(n11802), .A2(n11801), .ZN(n11804) );
  XNOR2_X1 U14757 ( .A(n13141), .B(n11804), .ZN(n13155) );
  XNOR2_X1 U14758 ( .A(n11803), .B(n12311), .ZN(n13153) );
  NAND2_X1 U14759 ( .A1(n13155), .A2(n13153), .ZN(n11806) );
  NAND2_X1 U14760 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11804), .ZN(
        n11805) );
  NAND2_X1 U14761 ( .A1(n11806), .A2(n11805), .ZN(n11807) );
  XNOR2_X1 U14762 ( .A(n11807), .B(n13500), .ZN(n13488) );
  NAND2_X1 U14763 ( .A1(n11807), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11808) );
  XNOR2_X1 U14764 ( .A(n11809), .B(n12324), .ZN(n11811) );
  INV_X1 U14765 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13788) );
  NAND2_X1 U14766 ( .A1(n13597), .A2(n13788), .ZN(n11814) );
  INV_X1 U14767 ( .A(n11810), .ZN(n11813) );
  INV_X1 U14768 ( .A(n11811), .ZN(n11812) );
  NAND2_X1 U14769 ( .A1(n11813), .A2(n11812), .ZN(n13598) );
  INV_X1 U14770 ( .A(n11797), .ZN(n11815) );
  NAND2_X1 U14771 ( .A1(n11815), .A2(n13789), .ZN(n13777) );
  INV_X1 U14772 ( .A(n13778), .ZN(n13781) );
  NAND2_X1 U14773 ( .A1(n13782), .A2(n13778), .ZN(n11820) );
  NAND2_X1 U14774 ( .A1(n11820), .A2(n11819), .ZN(n11821) );
  BUF_X1 U14775 ( .A(n11822), .Z(n11823) );
  INV_X1 U14776 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16336) );
  NAND2_X1 U14777 ( .A1(n13951), .A2(n11825), .ZN(n11831) );
  NAND3_X1 U14778 ( .A1(n16287), .A2(n16285), .A3(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11829) );
  INV_X1 U14779 ( .A(n11823), .ZN(n11828) );
  INV_X1 U14780 ( .A(n11826), .ZN(n11827) );
  NAND2_X1 U14781 ( .A1(n11828), .A2(n11827), .ZN(n16284) );
  NAND2_X1 U14782 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15808) );
  INV_X1 U14783 ( .A(n15808), .ZN(n11832) );
  AND2_X1 U14784 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15754) );
  AND3_X1 U14785 ( .A1(n15754), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15534) );
  AND2_X1 U14786 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n15534), .ZN(
        n11833) );
  OR2_X1 U14787 ( .A1(n15508), .A2(n15696), .ZN(n15501) );
  INV_X1 U14788 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15641) );
  INV_X1 U14789 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15414) );
  NAND2_X1 U14790 ( .A1(n14188), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11837) );
  XNOR2_X1 U14791 ( .A(n11837), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14177) );
  NAND2_X1 U14792 ( .A1(n12283), .A2(n11388), .ZN(n12916) );
  NOR2_X2 U14793 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19939) );
  NOR2_X1 U14794 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18952) );
  OR2_X1 U14795 ( .A1(n19939), .A2(n18952), .ZN(n19947) );
  NAND2_X1 U14796 ( .A1(n19947), .A2(n19987), .ZN(n11838) );
  NAND2_X1 U14797 ( .A1(n19987), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13114) );
  INV_X1 U14798 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19643) );
  NAND2_X1 U14799 ( .A1(n19643), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11839) );
  NAND2_X1 U14800 ( .A1(n13114), .A2(n11839), .ZN(n13109) );
  NOR2_X1 U14801 ( .A1(n11841), .A2(n15557), .ZN(n11842) );
  INV_X1 U14802 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11843) );
  INV_X1 U14803 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15545) );
  INV_X1 U14804 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11844) );
  OR2_X1 U14805 ( .A1(n11844), .A2(n15521), .ZN(n11845) );
  INV_X1 U14806 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15499) );
  NAND2_X1 U14807 ( .A1(n12771), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12772) );
  INV_X1 U14808 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15441) );
  NAND2_X1 U14809 ( .A1(n12793), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12769) );
  INV_X1 U14810 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15422) );
  NOR2_X2 U14811 ( .A1(n12769), .A2(n15422), .ZN(n12766) );
  INV_X1 U14812 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12767) );
  NAND2_X1 U14813 ( .A1(n12766), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12764) );
  INV_X1 U14814 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15399) );
  INV_X1 U14815 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11847) );
  NAND2_X1 U14816 ( .A1(n11850), .A2(n11849), .ZN(n11851) );
  NAND2_X1 U14817 ( .A1(n11852), .A2(n11851), .ZN(n11855) );
  BUF_X1 U14818 ( .A(n11856), .Z(n11857) );
  OR2_X1 U14819 ( .A1(n11857), .A2(n13788), .ZN(n11863) );
  INV_X1 U14820 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11860) );
  INV_X1 U14821 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11859) );
  OAI22_X1 U14822 ( .A1(n11957), .A2(n11860), .B1(n11444), .B2(n11859), .ZN(
        n11861) );
  AOI21_X1 U14823 ( .B1(n11897), .B2(P2_EBX_REG_4__SCAN_IN), .A(n11861), .ZN(
        n11862) );
  NAND2_X1 U14824 ( .A1(n11863), .A2(n11862), .ZN(n13211) );
  OR2_X1 U14825 ( .A1(n11857), .A2(n13789), .ZN(n11867) );
  INV_X1 U14826 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n11864) );
  OAI22_X1 U14827 ( .A1(n11957), .A2(n11864), .B1(n11444), .B2(n16309), .ZN(
        n11865) );
  AOI21_X1 U14828 ( .B1(n11897), .B2(P2_EBX_REG_5__SCAN_IN), .A(n11865), .ZN(
        n11866) );
  INV_X1 U14829 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13932) );
  OR2_X1 U14830 ( .A1(n11857), .A2(n13932), .ZN(n11872) );
  INV_X1 U14831 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n11869) );
  INV_X1 U14832 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11868) );
  OAI22_X1 U14833 ( .A1(n11957), .A2(n11869), .B1(n11444), .B2(n11868), .ZN(
        n11870) );
  AOI21_X1 U14834 ( .B1(n11897), .B2(P2_EBX_REG_6__SCAN_IN), .A(n11870), .ZN(
        n11871) );
  NAND2_X1 U14835 ( .A1(n11872), .A2(n11871), .ZN(n13221) );
  AOI22_X1 U14836 ( .A1(n11873), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11874) );
  OAI21_X1 U14837 ( .B1(n11900), .B2(n13273), .A(n11874), .ZN(n11875) );
  AOI21_X1 U14838 ( .B1(n11453), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n11875), .ZN(n13272) );
  OR2_X1 U14839 ( .A1(n11857), .A2(n16336), .ZN(n11878) );
  INV_X1 U14840 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n13590) );
  OAI22_X1 U14841 ( .A1(n11957), .A2(n13590), .B1(n11444), .B2(n11841), .ZN(
        n11876) );
  AOI21_X1 U14842 ( .B1(n11897), .B2(P2_EBX_REG_8__SCAN_IN), .A(n11876), .ZN(
        n11877) );
  NAND2_X1 U14843 ( .A1(n11878), .A2(n11877), .ZN(n13349) );
  NAND2_X1 U14844 ( .A1(n13271), .A2(n13349), .ZN(n13355) );
  OR2_X1 U14845 ( .A1(n11857), .A2(n15810), .ZN(n11882) );
  INV_X1 U14846 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n11879) );
  OAI22_X1 U14847 ( .A1(n11957), .A2(n11879), .B1(n11444), .B2(n15557), .ZN(
        n11880) );
  AOI21_X1 U14848 ( .B1(n11897), .B2(P2_EBX_REG_9__SCAN_IN), .A(n11880), .ZN(
        n11881) );
  INV_X1 U14849 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11883) );
  OR2_X1 U14850 ( .A1(n11857), .A2(n11883), .ZN(n11887) );
  INV_X1 U14851 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n13578) );
  INV_X1 U14852 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11884) );
  OAI22_X1 U14853 ( .A1(n11957), .A2(n13578), .B1(n11444), .B2(n11884), .ZN(
        n11885) );
  AOI21_X1 U14854 ( .B1(n11897), .B2(P2_EBX_REG_10__SCAN_IN), .A(n11885), .ZN(
        n11886) );
  NAND2_X1 U14855 ( .A1(n11887), .A2(n11886), .ZN(n13515) );
  INV_X1 U14856 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15802) );
  OR2_X1 U14857 ( .A1(n11857), .A2(n15802), .ZN(n11891) );
  INV_X1 U14858 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n11888) );
  OAI22_X1 U14859 ( .A1(n11957), .A2(n11888), .B1(n11444), .B2(n19074), .ZN(
        n11889) );
  AOI21_X1 U14860 ( .B1(n11897), .B2(P2_EBX_REG_11__SCAN_IN), .A(n11889), .ZN(
        n11890) );
  OR2_X1 U14861 ( .A1(n11857), .A2(n11704), .ZN(n11894) );
  INV_X1 U14862 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n12425) );
  OAI22_X1 U14863 ( .A1(n11957), .A2(n12425), .B1(n11444), .B2(n11843), .ZN(
        n11892) );
  AOI21_X1 U14864 ( .B1(n11897), .B2(P2_EBX_REG_12__SCAN_IN), .A(n11892), .ZN(
        n11893) );
  NAND2_X1 U14865 ( .A1(n11894), .A2(n11893), .ZN(n13665) );
  OR2_X1 U14866 ( .A1(n11857), .A2(n15769), .ZN(n11899) );
  INV_X1 U14867 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n11895) );
  OAI22_X1 U14868 ( .A1(n11957), .A2(n11895), .B1(n11444), .B2(n16253), .ZN(
        n11896) );
  AOI21_X1 U14869 ( .B1(n11897), .B2(P2_EBX_REG_13__SCAN_IN), .A(n11896), .ZN(
        n11898) );
  NAND2_X1 U14870 ( .A1(n11899), .A2(n11898), .ZN(n13685) );
  NAND2_X1 U14871 ( .A1(n13664), .A2(n13685), .ZN(n13684) );
  INV_X1 U14872 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15753) );
  OR2_X1 U14873 ( .A1(n11857), .A2(n15753), .ZN(n11905) );
  INV_X1 U14874 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n11902) );
  INV_X1 U14875 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11901) );
  OAI22_X1 U14876 ( .A1(n11957), .A2(n11902), .B1(n11444), .B2(n11901), .ZN(
        n11903) );
  AOI21_X1 U14877 ( .B1(n11897), .B2(P2_EBX_REG_14__SCAN_IN), .A(n11903), .ZN(
        n11904) );
  OR2_X1 U14878 ( .A1(n11857), .A2(n15543), .ZN(n11908) );
  INV_X1 U14879 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19888) );
  OAI22_X1 U14880 ( .A1(n11957), .A2(n19888), .B1(n11444), .B2(n15545), .ZN(
        n11906) );
  AOI21_X1 U14881 ( .B1(n11897), .B2(P2_EBX_REG_15__SCAN_IN), .A(n11906), .ZN(
        n11907) );
  OR2_X1 U14882 ( .A1(n11857), .A2(n15721), .ZN(n11911) );
  INV_X1 U14883 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19890) );
  INV_X1 U14884 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n19024) );
  OAI22_X1 U14885 ( .A1(n11957), .A2(n19890), .B1(n11444), .B2(n19024), .ZN(
        n11909) );
  AOI21_X1 U14886 ( .B1(n11897), .B2(P2_EBX_REG_16__SCAN_IN), .A(n11909), .ZN(
        n11910) );
  OR2_X1 U14887 ( .A1(n11857), .A2(n15508), .ZN(n11914) );
  INV_X1 U14888 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19892) );
  OAI22_X1 U14889 ( .A1(n11957), .A2(n19892), .B1(n11444), .B2(n15521), .ZN(
        n11912) );
  AOI21_X1 U14890 ( .B1(n11897), .B2(P2_EBX_REG_17__SCAN_IN), .A(n11912), .ZN(
        n11913) );
  NAND2_X1 U14891 ( .A1(n11914), .A2(n11913), .ZN(n13892) );
  OR2_X1 U14892 ( .A1(n11857), .A2(n15696), .ZN(n11917) );
  INV_X1 U14893 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15223) );
  OAI22_X1 U14894 ( .A1(n11957), .A2(n15223), .B1(n11444), .B2(n11844), .ZN(
        n11915) );
  AOI21_X1 U14895 ( .B1(n11897), .B2(P2_EBX_REG_18__SCAN_IN), .A(n11915), .ZN(
        n11916) );
  OR2_X1 U14896 ( .A1(n11857), .A2(n15684), .ZN(n11920) );
  INV_X1 U14897 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19895) );
  OAI22_X1 U14898 ( .A1(n11957), .A2(n19895), .B1(n11444), .B2(n15499), .ZN(
        n11918) );
  AOI21_X1 U14899 ( .B1(n11897), .B2(P2_EBX_REG_19__SCAN_IN), .A(n11918), .ZN(
        n11919) );
  OR2_X1 U14900 ( .A1(n11857), .A2(n15673), .ZN(n11924) );
  INV_X1 U14901 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n15485) );
  INV_X1 U14902 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11921) );
  OAI22_X1 U14903 ( .A1(n11957), .A2(n15485), .B1(n11444), .B2(n11921), .ZN(
        n11922) );
  AOI21_X1 U14904 ( .B1(n11897), .B2(P2_EBX_REG_20__SCAN_IN), .A(n11922), .ZN(
        n11923) );
  NAND2_X1 U14905 ( .A1(n11924), .A2(n11923), .ZN(n15299) );
  OR2_X1 U14906 ( .A1(n11857), .A2(n15473), .ZN(n11927) );
  INV_X1 U14907 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19898) );
  OAI22_X1 U14908 ( .A1(n11957), .A2(n19898), .B1(n11444), .B2(n11846), .ZN(
        n11925) );
  AOI21_X1 U14909 ( .B1(n11897), .B2(P2_EBX_REG_21__SCAN_IN), .A(n11925), .ZN(
        n11926) );
  NAND2_X1 U14910 ( .A1(n11927), .A2(n11926), .ZN(n15290) );
  OR2_X1 U14911 ( .A1(n11857), .A2(n15641), .ZN(n11931) );
  INV_X1 U14912 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19900) );
  INV_X1 U14913 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11928) );
  OAI22_X1 U14914 ( .A1(n11957), .A2(n19900), .B1(n11444), .B2(n11928), .ZN(
        n11929) );
  AOI21_X1 U14915 ( .B1(n11897), .B2(P2_EBX_REG_22__SCAN_IN), .A(n11929), .ZN(
        n11930) );
  OR2_X1 U14916 ( .A1(n11857), .A2(n15633), .ZN(n11934) );
  INV_X1 U14917 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19902) );
  OAI22_X1 U14918 ( .A1(n11957), .A2(n19902), .B1(n11444), .B2(n15441), .ZN(
        n11932) );
  AOI21_X1 U14919 ( .B1(n11897), .B2(P2_EBX_REG_23__SCAN_IN), .A(n11932), .ZN(
        n11933) );
  OR2_X1 U14920 ( .A1(n11857), .A2(n15619), .ZN(n11938) );
  INV_X1 U14921 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n11935) );
  INV_X1 U14922 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15433) );
  OAI22_X1 U14923 ( .A1(n11957), .A2(n11935), .B1(n11444), .B2(n15433), .ZN(
        n11936) );
  AOI21_X1 U14924 ( .B1(n11897), .B2(P2_EBX_REG_24__SCAN_IN), .A(n11936), .ZN(
        n11937) );
  NAND2_X1 U14925 ( .A1(n11938), .A2(n11937), .ZN(n15266) );
  OR2_X1 U14926 ( .A1(n11857), .A2(n15607), .ZN(n11941) );
  INV_X1 U14927 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19905) );
  OAI22_X1 U14928 ( .A1(n11957), .A2(n19905), .B1(n11444), .B2(n15422), .ZN(
        n11939) );
  AOI21_X1 U14929 ( .B1(n11897), .B2(P2_EBX_REG_25__SCAN_IN), .A(n11939), .ZN(
        n11940) );
  NAND2_X1 U14930 ( .A1(n11941), .A2(n11940), .ZN(n15211) );
  OR2_X1 U14931 ( .A1(n11857), .A2(n15414), .ZN(n11944) );
  INV_X1 U14932 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19907) );
  OAI22_X1 U14933 ( .A1(n11957), .A2(n19907), .B1(n11444), .B2(n12767), .ZN(
        n11942) );
  AOI21_X1 U14934 ( .B1(n11897), .B2(P2_EBX_REG_26__SCAN_IN), .A(n11942), .ZN(
        n11943) );
  INV_X1 U14935 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12555) );
  OR2_X1 U14936 ( .A1(n11857), .A2(n12555), .ZN(n11947) );
  INV_X1 U14937 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19910) );
  OAI22_X1 U14938 ( .A1(n11957), .A2(n19910), .B1(n11444), .B2(n15399), .ZN(
        n11945) );
  AOI21_X1 U14939 ( .B1(n11897), .B2(P2_EBX_REG_27__SCAN_IN), .A(n11945), .ZN(
        n11946) );
  OR2_X1 U14940 ( .A1(n11857), .A2(n15564), .ZN(n11950) );
  INV_X1 U14941 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19911) );
  INV_X1 U14942 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14202) );
  OAI22_X1 U14943 ( .A1(n11957), .A2(n19911), .B1(n11444), .B2(n14202), .ZN(
        n11948) );
  AOI21_X1 U14944 ( .B1(n11897), .B2(P2_EBX_REG_28__SCAN_IN), .A(n11948), .ZN(
        n11949) );
  NAND2_X1 U14945 ( .A1(n11950), .A2(n11949), .ZN(n14197) );
  OR2_X1 U14946 ( .A1(n11857), .A2(n12287), .ZN(n11953) );
  INV_X1 U14947 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19913) );
  INV_X1 U14948 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15389) );
  OAI22_X1 U14949 ( .A1(n11957), .A2(n19913), .B1(n11444), .B2(n15389), .ZN(
        n11951) );
  AOI21_X1 U14950 ( .B1(n11897), .B2(P2_EBX_REG_29__SCAN_IN), .A(n11951), .ZN(
        n11952) );
  AND2_X1 U14951 ( .A1(n11953), .A2(n11952), .ZN(n12551) );
  INV_X1 U14952 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14208) );
  OR2_X1 U14953 ( .A1(n11857), .A2(n14208), .ZN(n11956) );
  INV_X1 U14954 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19917) );
  INV_X1 U14955 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14189) );
  OAI22_X1 U14956 ( .A1(n11957), .A2(n19917), .B1(n11444), .B2(n14189), .ZN(
        n11954) );
  AOI21_X1 U14957 ( .B1(n11897), .B2(P2_EBX_REG_30__SCAN_IN), .A(n11954), .ZN(
        n11955) );
  AND2_X1 U14958 ( .A1(n11956), .A2(n11955), .ZN(n12807) );
  INV_X1 U14959 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12762) );
  AOI22_X1 U14960 ( .A1(n11873), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11959) );
  NAND2_X1 U14961 ( .A1(n11897), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n11958) );
  OAI211_X1 U14962 ( .C1(n11857), .C2(n12762), .A(n11959), .B(n11958), .ZN(
        n11960) );
  NAND2_X1 U14963 ( .A1(n11961), .A2(n12811), .ZN(n11982) );
  NOR2_X1 U14964 ( .A1(n11963), .A2(n11962), .ZN(n11969) );
  NAND2_X1 U14965 ( .A1(n11551), .A2(n11963), .ZN(n11965) );
  NAND3_X1 U14966 ( .A1(n11965), .A2(n16366), .A3(n11964), .ZN(n11968) );
  NAND2_X1 U14967 ( .A1(n11966), .A2(n11970), .ZN(n11967) );
  OAI211_X1 U14968 ( .C1(n12811), .C2(n11969), .A(n11968), .B(n11967), .ZN(
        n11975) );
  INV_X1 U14969 ( .A(n19986), .ZN(n13026) );
  INV_X1 U14970 ( .A(n11970), .ZN(n11971) );
  OAI21_X1 U14971 ( .B1(n13026), .B2(n11551), .A(n11971), .ZN(n11972) );
  NAND2_X1 U14972 ( .A1(n11973), .A2(n11972), .ZN(n11974) );
  NAND2_X1 U14973 ( .A1(n11975), .A2(n11974), .ZN(n11977) );
  NAND2_X1 U14974 ( .A1(n11977), .A2(n11976), .ZN(n11981) );
  NOR2_X1 U14975 ( .A1(n11978), .A2(n12811), .ZN(n11979) );
  AOI21_X1 U14976 ( .B1(n11982), .B2(n11981), .A(n11980), .ZN(n11983) );
  MUX2_X1 U14977 ( .A(n11983), .B(n15903), .S(n19987), .Z(n12263) );
  AOI21_X1 U14978 ( .B1(n19769), .B2(n11444), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19984) );
  NAND2_X1 U14979 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19958) );
  NAND2_X1 U14980 ( .A1(n19984), .A2(n19958), .ZN(n11986) );
  NAND2_X1 U14981 ( .A1(n16186), .A2(n16306), .ZN(n11990) );
  INV_X1 U14982 ( .A(n19979), .ZN(n11987) );
  AND2_X1 U14983 ( .A1(n11987), .A2(n19939), .ZN(n11988) );
  INV_X2 U14984 ( .A(n11988), .ZN(n19113) );
  INV_X1 U14985 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19920) );
  NOR2_X1 U14986 ( .A1(n19113), .A2(n19920), .ZN(n14172) );
  AOI21_X1 U14987 ( .B1(n19231), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14172), .ZN(n11989) );
  OAI211_X1 U14988 ( .C1(n19240), .C2(n12763), .A(n11990), .B(n11989), .ZN(
        n11991) );
  AOI21_X1 U14989 ( .B1(n14177), .B2(n19236), .A(n11991), .ZN(n11992) );
  OAI21_X1 U14990 ( .B1(n11993), .B2(n14180), .A(n11992), .ZN(P2_U2983) );
  INV_X1 U14991 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16593) );
  NAND2_X1 U14992 ( .A1(n17816), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16801) );
  NOR2_X2 U14993 ( .A1(n17739), .A2(n17740), .ZN(n17711) );
  INV_X1 U14994 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17662) );
  INV_X1 U14995 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17622) );
  INV_X1 U14996 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17908) );
  NAND2_X1 U14997 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17606) );
  INV_X1 U14998 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11998) );
  INV_X1 U14999 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17565) );
  INV_X1 U15000 ( .A(n12722), .ZN(n11995) );
  XNOR2_X1 U15001 ( .A(n9893), .B(n12001), .ZN(n16574) );
  AOI21_X1 U15002 ( .B1(n16593), .B2(n11995), .A(n12001), .ZN(n16587) );
  OAI21_X1 U15003 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n11996), .A(
        n12011), .ZN(n17582) );
  INV_X1 U15004 ( .A(n17582), .ZN(n16606) );
  AOI21_X1 U15005 ( .B1(n11998), .B2(n11997), .A(n11996), .ZN(n17584) );
  INV_X1 U15006 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17616) );
  AOI22_X1 U15007 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n12009), .B1(
        n11999), .B2(n17616), .ZN(n17612) );
  INV_X1 U15008 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17639) );
  INV_X1 U15009 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17651) );
  NOR3_X1 U15010 ( .A1(n17908), .A2(n17698), .A3(n17699), .ZN(n17675) );
  NAND3_X1 U15011 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A3(n17675), .ZN(n17635) );
  INV_X1 U15012 ( .A(n17635), .ZN(n16693) );
  NAND2_X1 U15013 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16693), .ZN(
        n12002) );
  OR2_X1 U15014 ( .A1(n17651), .A2(n12002), .ZN(n12000) );
  NOR2_X1 U15015 ( .A1(n17908), .A2(n17623), .ZN(n12006) );
  AOI21_X1 U15016 ( .B1(n17639), .B2(n12000), .A(n12006), .ZN(n17642) );
  OAI21_X1 U15017 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n16693), .A(
        n12002), .ZN(n17666) );
  INV_X1 U15018 ( .A(n17666), .ZN(n16685) );
  INV_X1 U15019 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16863) );
  NOR2_X1 U15020 ( .A1(n16685), .A2(n16684), .ZN(n16683) );
  NOR2_X1 U15021 ( .A1(n16683), .A2(n16862), .ZN(n16673) );
  INV_X1 U15022 ( .A(n16673), .ZN(n12004) );
  XOR2_X1 U15023 ( .A(n17651), .B(n12002), .Z(n17654) );
  NAND2_X1 U15024 ( .A1(n12004), .A2(n12003), .ZN(n16671) );
  INV_X1 U15025 ( .A(n16862), .ZN(n12005) );
  NOR2_X1 U15026 ( .A1(n17642), .A2(n16663), .ZN(n16662) );
  NOR2_X1 U15027 ( .A1(n16662), .A2(n16862), .ZN(n16651) );
  INV_X1 U15028 ( .A(n16651), .ZN(n12008) );
  INV_X1 U15029 ( .A(n12006), .ZN(n17596) );
  AOI21_X1 U15030 ( .B1(n17622), .B2(n17596), .A(n12009), .ZN(n17625) );
  INV_X1 U15031 ( .A(n17625), .ZN(n12007) );
  NAND2_X1 U15032 ( .A1(n12008), .A2(n12007), .ZN(n16649) );
  NOR2_X1 U15033 ( .A1(n17612), .A2(n16641), .ZN(n16640) );
  NOR2_X1 U15034 ( .A1(n16640), .A2(n16862), .ZN(n16630) );
  INV_X1 U15035 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16632) );
  NAND2_X1 U15036 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n12009), .ZN(
        n12010) );
  AOI21_X1 U15037 ( .B1(n16632), .B2(n12010), .A(n17562), .ZN(n17597) );
  NOR2_X1 U15038 ( .A1(n17584), .A2(n16619), .ZN(n16618) );
  NOR2_X1 U15039 ( .A1(n16618), .A2(n16862), .ZN(n16605) );
  NOR2_X1 U15040 ( .A1(n16606), .A2(n16605), .ZN(n16604) );
  OR2_X1 U15041 ( .A1(n16604), .A2(n16862), .ZN(n16596) );
  AOI21_X1 U15042 ( .B1(n17565), .B2(n12011), .A(n12722), .ZN(n17554) );
  INV_X1 U15043 ( .A(n17554), .ZN(n12012) );
  NAND2_X1 U15044 ( .A1(n16596), .A2(n12012), .ZN(n16597) );
  NOR2_X1 U15045 ( .A1(n16587), .A2(n16586), .ZN(n16585) );
  NOR2_X1 U15046 ( .A1(n16585), .A2(n16862), .ZN(n16573) );
  INV_X1 U15047 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18253) );
  INV_X1 U15048 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18783) );
  INV_X1 U15049 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18931) );
  NAND4_X1 U15050 ( .A1(n18253), .A2(n18783), .A3(n18931), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n16913) );
  NOR2_X1 U15051 ( .A1(n16862), .A2(n16913), .ZN(n16768) );
  INV_X1 U15052 ( .A(n16768), .ZN(n12013) );
  NOR3_X1 U15053 ( .A1(n16574), .A2(n16573), .A3(n12013), .ZN(n12152) );
  INV_X2 U15054 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12014) );
  INV_X4 U15055 ( .A(n17208), .ZN(n17230) );
  INV_X1 U15056 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12016) );
  NAND2_X2 U15057 ( .A1(n18897), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12020) );
  AOI22_X1 U15058 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17225), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12015) );
  OAI21_X1 U15059 ( .B1(n17241), .B2(n12016), .A(n12015), .ZN(n12032) );
  AOI22_X1 U15060 ( .A1(n17202), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12030) );
  OR2_X2 U15061 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12017), .ZN(
        n17163) );
  INV_X4 U15062 ( .A(n17163), .ZN(n17228) );
  OAI22_X1 U15063 ( .A1(n17205), .A2(n17207), .B1(n17184), .B2(n18516), .ZN(
        n12028) );
  INV_X2 U15064 ( .A(n12643), .ZN(n12100) );
  AOI22_X1 U15065 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12026) );
  INV_X4 U15066 ( .A(n17099), .ZN(n17229) );
  INV_X2 U15067 ( .A(n12562), .ZN(n17223) );
  AOI22_X1 U15068 ( .A1(n17229), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12025) );
  NOR2_X2 U15069 ( .A1(n12023), .A2(n18897), .ZN(n18712) );
  AOI22_X1 U15070 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17209), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12024) );
  NAND3_X1 U15071 ( .A1(n12026), .A2(n12025), .A3(n12024), .ZN(n12027) );
  OAI211_X1 U15072 ( .C1(n17227), .C2(n18601), .A(n12030), .B(n12029), .ZN(
        n12031) );
  AOI211_X4 U15073 ( .C1(n17230), .C2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n12032), .B(n12031), .ZN(n18932) );
  INV_X1 U15074 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17234) );
  INV_X1 U15075 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17240) );
  AOI22_X1 U15076 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12035) );
  INV_X2 U15077 ( .A(n17035), .ZN(n17224) );
  AOI22_X1 U15078 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12034) );
  OAI211_X1 U15079 ( .C1(n17235), .C2(n17240), .A(n12035), .B(n12034), .ZN(
        n12041) );
  INV_X2 U15080 ( .A(n12086), .ZN(n17148) );
  AOI22_X1 U15081 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12039) );
  AOI22_X1 U15082 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12038) );
  INV_X2 U15083 ( .A(n9699), .ZN(n17225) );
  AOI22_X1 U15084 ( .A1(n17225), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17161), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12037) );
  NAND2_X1 U15085 ( .A1(n17204), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12036) );
  NAND4_X1 U15086 ( .A1(n12039), .A2(n12038), .A3(n12037), .A4(n12036), .ZN(
        n12040) );
  INV_X1 U15087 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17116) );
  AOI22_X1 U15088 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12044) );
  OAI21_X1 U15089 ( .B1(n12608), .B2(n17116), .A(n12044), .ZN(n12052) );
  INV_X1 U15090 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15091 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12049) );
  INV_X1 U15092 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17115) );
  INV_X1 U15093 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16969) );
  OAI22_X1 U15094 ( .A1(n17035), .A2(n17115), .B1(n17205), .B2(n16969), .ZN(
        n12047) );
  AOI22_X1 U15095 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12046) );
  INV_X2 U15096 ( .A(n17217), .ZN(n17186) );
  AOI22_X1 U15097 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17209), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12045) );
  OAI211_X1 U15098 ( .C1(n17227), .C2(n12050), .A(n12049), .B(n12048), .ZN(
        n12051) );
  INV_X1 U15099 ( .A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17166) );
  AOI22_X1 U15100 ( .A1(n17225), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12053) );
  OAI21_X1 U15101 ( .B1(n17217), .B2(n17166), .A(n12053), .ZN(n12062) );
  INV_X1 U15102 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14082) );
  AOI22_X1 U15103 ( .A1(n17204), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12060) );
  INV_X1 U15104 ( .A(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17162) );
  AOI22_X1 U15105 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17209), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12054) );
  OAI21_X1 U15106 ( .B1(n17099), .B2(n17162), .A(n12054), .ZN(n12058) );
  INV_X1 U15107 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14083) );
  AOI22_X1 U15108 ( .A1(n17202), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15863), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12056) );
  AOI22_X1 U15109 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12055) );
  OAI211_X1 U15110 ( .C1(n17167), .C2(n14083), .A(n12056), .B(n12055), .ZN(
        n12057) );
  AOI211_X1 U15111 ( .C1(n12616), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n12058), .B(n12057), .ZN(n12059) );
  OAI211_X1 U15112 ( .C1(n17241), .C2(n14082), .A(n12060), .B(n12059), .ZN(
        n12061) );
  AOI211_X4 U15113 ( .C1(n17230), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n12062), .B(n12061), .ZN(n18277) );
  INV_X1 U15114 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17022) );
  OAI22_X1 U15115 ( .A1(n17227), .A2(n15873), .B1(n17167), .B2(n17022), .ZN(
        n12067) );
  INV_X2 U15116 ( .A(n17114), .ZN(n15863) );
  AOI22_X1 U15117 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15863), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U15118 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U15119 ( .A1(n12616), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17209), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12063) );
  NAND3_X1 U15120 ( .A1(n12065), .A2(n12064), .A3(n12063), .ZN(n12066) );
  AOI211_X1 U15121 ( .C1(n17101), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n12067), .B(n12066), .ZN(n12075) );
  INV_X1 U15122 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14070) );
  AOI22_X1 U15123 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(n9652), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12068) );
  OAI21_X1 U15124 ( .B1(n9699), .B2(n14070), .A(n12068), .ZN(n12069) );
  INV_X1 U15125 ( .A(n12069), .ZN(n12074) );
  AOI22_X1 U15126 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12073) );
  INV_X1 U15127 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17034) );
  INV_X1 U15128 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17183) );
  AOI22_X1 U15129 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12076) );
  OAI21_X1 U15130 ( .B1(n17241), .B2(n17183), .A(n12076), .ZN(n12085) );
  INV_X1 U15131 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17276) );
  AOI22_X1 U15132 ( .A1(n17225), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12083) );
  INV_X1 U15133 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17071) );
  OAI22_X1 U15134 ( .A1(n17227), .A2(n18605), .B1(n17205), .B2(n17071), .ZN(
        n12081) );
  AOI22_X1 U15135 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15136 ( .A1(n17202), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15137 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17209), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12077) );
  NAND3_X1 U15138 ( .A1(n12079), .A2(n12078), .A3(n12077), .ZN(n12080) );
  AOI211_X1 U15139 ( .C1(n9635), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n12081), .B(n12080), .ZN(n12082) );
  OAI211_X1 U15140 ( .C1(n12562), .C2(n17276), .A(n12083), .B(n12082), .ZN(
        n12084) );
  AOI211_X4 U15141 ( .C1(n17142), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n12085), .B(n12084), .ZN(n18273) );
  INV_X1 U15142 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17040) );
  AOI22_X1 U15143 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12087) );
  OAI21_X1 U15144 ( .B1(n12608), .B2(n17040), .A(n12087), .ZN(n12098) );
  INV_X1 U15145 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17145) );
  AOI22_X1 U15146 ( .A1(n17225), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17204), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12096) );
  INV_X1 U15147 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14133) );
  INV_X1 U15148 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17041) );
  OAI22_X1 U15149 ( .A1(n17205), .A2(n14133), .B1(n12100), .B2(n17041), .ZN(
        n12094) );
  AOI22_X1 U15150 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15863), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U15151 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U15152 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17209), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12090) );
  NAND3_X1 U15153 ( .A1(n12092), .A2(n12091), .A3(n12090), .ZN(n12093) );
  AOI211_X1 U15154 ( .C1(n17228), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n12094), .B(n12093), .ZN(n12095) );
  OAI211_X1 U15155 ( .C1(n17208), .C2(n17145), .A(n12096), .B(n12095), .ZN(
        n12097) );
  AOI211_X2 U15156 ( .C1(n17101), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n12098), .B(n12097), .ZN(n18281) );
  AOI22_X1 U15157 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15863), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12099) );
  OAI21_X1 U15158 ( .B1(n12562), .B2(n17256), .A(n12099), .ZN(n12109) );
  AOI22_X1 U15159 ( .A1(n17225), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12107) );
  AOI22_X1 U15160 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U15161 ( .A1(n12616), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17209), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12105) );
  INV_X1 U15162 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16949) );
  INV_X1 U15163 ( .A(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17007) );
  OAI22_X1 U15164 ( .A1(n17227), .A2(n16949), .B1(n12100), .B2(n17007), .ZN(
        n12103) );
  INV_X1 U15165 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16958) );
  AOI22_X1 U15166 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12101) );
  OAI21_X1 U15167 ( .B1(n17167), .B2(n16958), .A(n12101), .ZN(n12102) );
  AOI211_X1 U15168 ( .C1(n17229), .C2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n12103), .B(n12102), .ZN(n12104) );
  NAND4_X1 U15169 ( .A1(n12107), .A2(n12106), .A3(n12105), .A4(n12104), .ZN(
        n12108) );
  INV_X1 U15170 ( .A(n9649), .ZN(n17292) );
  NAND2_X1 U15171 ( .A1(n12110), .A2(n17292), .ZN(n12113) );
  NOR2_X2 U15172 ( .A1(n17485), .A2(n15889), .ZN(n16555) );
  NAND2_X1 U15173 ( .A1(n18273), .A2(n12110), .ZN(n15911) );
  NAND2_X1 U15174 ( .A1(n12110), .A2(n9649), .ZN(n15992) );
  INV_X1 U15175 ( .A(n15992), .ZN(n18739) );
  NOR2_X1 U15176 ( .A1(n17291), .A2(n18739), .ZN(n15991) );
  NAND2_X1 U15177 ( .A1(n18932), .A2(n18267), .ZN(n12111) );
  AOI21_X1 U15178 ( .B1(n15911), .B2(n12112), .A(n15893), .ZN(n12121) );
  AOI21_X1 U15179 ( .B1(n18294), .B2(n12113), .A(n18281), .ZN(n12119) );
  NOR2_X1 U15180 ( .A1(n18932), .A2(n18267), .ZN(n12114) );
  INV_X1 U15181 ( .A(n18273), .ZN(n15908) );
  NOR2_X1 U15182 ( .A1(n12114), .A2(n15908), .ZN(n12718) );
  OAI21_X1 U15183 ( .B1(n15908), .B2(n18267), .A(n15992), .ZN(n12115) );
  OAI21_X1 U15184 ( .B1(n15906), .B2(n12116), .A(n12115), .ZN(n12117) );
  OAI21_X1 U15185 ( .B1(n15906), .B2(n12718), .A(n12117), .ZN(n12118) );
  AOI211_X2 U15186 ( .C1(n18277), .C2(n12120), .A(n12119), .B(n12118), .ZN(
        n15890) );
  OAI21_X1 U15187 ( .B1(n18277), .B2(n12121), .A(n15890), .ZN(n12712) );
  NOR2_X2 U15188 ( .A1(n12122), .A2(n12712), .ZN(n18720) );
  NAND2_X1 U15189 ( .A1(n17292), .A2(n18286), .ZN(n12717) );
  INV_X1 U15190 ( .A(n14064), .ZN(n12123) );
  NAND3_X1 U15191 ( .A1(n12124), .A2(n18932), .A3(n12123), .ZN(n12125) );
  INV_X2 U15192 ( .A(n15898), .ZN(n18730) );
  NAND3_X1 U15193 ( .A1(n18905), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18781) );
  NAND2_X1 U15194 ( .A1(n18539), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12706) );
  AOI22_X1 U15195 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n18743), .B2(n12023), .ZN(
        n12710) );
  XNOR2_X1 U15196 ( .A(n12706), .B(n12710), .ZN(n12137) );
  AOI22_X1 U15197 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18761), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18897), .ZN(n12132) );
  NAND2_X1 U15198 ( .A1(n12132), .A2(n12133), .ZN(n12129) );
  OAI21_X1 U15199 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18897), .A(
        n12129), .ZN(n12130) );
  OAI22_X1 U15200 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18763), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12130), .ZN(n12134) );
  NOR2_X1 U15201 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18763), .ZN(
        n12131) );
  NAND2_X1 U15202 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12130), .ZN(
        n12135) );
  AOI22_X1 U15203 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12134), .B1(
        n12131), .B2(n12135), .ZN(n12707) );
  XOR2_X1 U15204 ( .A(n12133), .B(n12132), .Z(n12714) );
  NAND2_X1 U15205 ( .A1(n12707), .A2(n12714), .ZN(n12708) );
  AOI21_X1 U15206 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12135), .A(
        n12134), .ZN(n12136) );
  AOI21_X1 U15207 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18763), .A(
        n12136), .ZN(n12709) );
  INV_X1 U15208 ( .A(n18943), .ZN(n18946) );
  NAND2_X1 U15209 ( .A1(n18905), .A2(n18883), .ZN(n18892) );
  NOR2_X1 U15210 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18892), .ZN(n18944) );
  AOI21_X1 U15211 ( .B1(n18905), .B2(n18653), .A(n18783), .ZN(n18777) );
  INV_X1 U15212 ( .A(n18777), .ZN(n12138) );
  OAI21_X1 U15213 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18944), .A(n12138), 
        .ZN(n12139) );
  INV_X1 U15214 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18807) );
  NOR2_X2 U15215 ( .A1(n18799), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18870) );
  NOR2_X1 U15216 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18793) );
  INV_X1 U15217 ( .A(n18793), .ZN(n16551) );
  NAND3_X1 U15218 ( .A1(n18807), .A2(n18873), .A3(n16551), .ZN(n18930) );
  NAND2_X1 U15219 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n18933) );
  INV_X1 U15220 ( .A(n18933), .ZN(n18785) );
  AOI211_X1 U15221 ( .C1(n18930), .C2(n18932), .A(n18785), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n12141) );
  INV_X1 U15222 ( .A(n12141), .ZN(n18776) );
  NOR2_X1 U15223 ( .A1(n16929), .A2(n16884), .ZN(n16692) );
  INV_X1 U15224 ( .A(n16692), .ZN(n16935) );
  INV_X1 U15225 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18866) );
  INV_X1 U15226 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18863) );
  INV_X1 U15227 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18860) );
  INV_X1 U15228 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18856) );
  INV_X1 U15229 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18849) );
  INV_X1 U15230 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18837) );
  INV_X1 U15231 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18832) );
  INV_X1 U15232 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18828) );
  INV_X1 U15233 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18824) );
  INV_X1 U15234 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18818) );
  INV_X1 U15235 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18816) );
  NAND3_X1 U15236 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16883) );
  NOR3_X1 U15237 ( .A1(n18818), .A2(n18816), .A3(n16883), .ZN(n16840) );
  NAND3_X1 U15238 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .A3(n16840), .ZN(n16831) );
  NOR2_X1 U15239 ( .A1(n18824), .A2(n16831), .ZN(n16806) );
  NAND2_X1 U15240 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16806), .ZN(n16803) );
  NOR2_X1 U15241 ( .A1(n18828), .A2(n16803), .ZN(n16788) );
  NAND2_X1 U15242 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16788), .ZN(n16783) );
  NOR2_X1 U15243 ( .A1(n18832), .A2(n16783), .ZN(n16765) );
  NAND2_X1 U15244 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16765), .ZN(n16717) );
  NOR2_X1 U15245 ( .A1(n18837), .A2(n16717), .ZN(n16753) );
  NAND4_X1 U15246 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16753), .A3(
        P3_REIP_REG_16__SCAN_IN), .A4(P3_REIP_REG_15__SCAN_IN), .ZN(n16681) );
  NAND2_X1 U15247 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16703) );
  NOR3_X1 U15248 ( .A1(n18849), .A2(n16681), .A3(n16703), .ZN(n16652) );
  NAND4_X1 U15249 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16652), .A3(
        P3_REIP_REG_22__SCAN_IN), .A4(P3_REIP_REG_21__SCAN_IN), .ZN(n16648) );
  NOR2_X1 U15250 ( .A1(n18856), .A2(n16648), .ZN(n16631) );
  NAND2_X1 U15251 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16631), .ZN(n16626) );
  NOR2_X1 U15252 ( .A1(n18860), .A2(n16626), .ZN(n16615) );
  NAND2_X1 U15253 ( .A1(n16884), .A2(n16615), .ZN(n16608) );
  NOR3_X1 U15254 ( .A1(n18866), .A2(n18863), .A3(n16608), .ZN(n16582) );
  NAND2_X1 U15255 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16582), .ZN(n12142) );
  NAND2_X1 U15256 ( .A1(n16935), .A2(n12142), .ZN(n16575) );
  INV_X1 U15257 ( .A(n16575), .ZN(n16590) );
  NOR2_X1 U15258 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n12142), .ZN(n16577) );
  OAI21_X1 U15259 ( .B1(n16590), .B2(n16577), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n12140) );
  AOI211_X4 U15260 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n15987), .A(n12141), .B(
        n12145), .ZN(n16891) );
  INV_X1 U15261 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18872) );
  NOR3_X1 U15262 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18872), .A3(n12142), 
        .ZN(n12143) );
  AOI21_X1 U15263 ( .B1(n16891), .B2(P3_EBX_REG_31__SCAN_IN), .A(n12143), .ZN(
        n12150) );
  NAND2_X1 U15264 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n15987), .ZN(n12144) );
  AOI211_X4 U15265 ( .C1(n18931), .C2(n18933), .A(n12145), .B(n12144), .ZN(
        n16901) );
  NOR3_X1 U15266 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16907) );
  INV_X1 U15267 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17267) );
  NAND2_X1 U15268 ( .A1(n16907), .A2(n17267), .ZN(n16900) );
  NOR2_X1 U15269 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16900), .ZN(n16878) );
  INV_X1 U15270 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16870) );
  NAND2_X1 U15271 ( .A1(n16878), .A2(n16870), .ZN(n16869) );
  NOR2_X1 U15272 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16869), .ZN(n16849) );
  INV_X1 U15273 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16846) );
  NAND2_X1 U15274 ( .A1(n16849), .A2(n16846), .ZN(n16845) );
  NOR2_X1 U15275 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16845), .ZN(n16816) );
  INV_X1 U15276 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n12146) );
  NAND2_X1 U15277 ( .A1(n16816), .A2(n12146), .ZN(n16808) );
  INV_X1 U15278 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16797) );
  NAND2_X1 U15279 ( .A1(n16807), .A2(n16797), .ZN(n16796) );
  INV_X1 U15280 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16772) );
  NAND2_X1 U15281 ( .A1(n16778), .A2(n16772), .ZN(n16769) );
  INV_X1 U15282 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16746) );
  NAND2_X1 U15283 ( .A1(n16754), .A2(n16746), .ZN(n16744) );
  INV_X1 U15284 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16721) );
  NAND2_X1 U15285 ( .A1(n16733), .A2(n16721), .ZN(n16719) );
  INV_X1 U15286 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16702) );
  NAND2_X1 U15287 ( .A1(n16707), .A2(n16702), .ZN(n16701) );
  INV_X1 U15288 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17038) );
  NAND2_X1 U15289 ( .A1(n16686), .A2(n17038), .ZN(n16678) );
  NOR2_X1 U15290 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16678), .ZN(n16664) );
  INV_X1 U15291 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16657) );
  NAND2_X1 U15292 ( .A1(n16664), .A2(n16657), .ZN(n16656) );
  NOR2_X1 U15293 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16656), .ZN(n16627) );
  INV_X1 U15294 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16984) );
  NAND2_X1 U15295 ( .A1(n16627), .A2(n16984), .ZN(n16617) );
  NOR2_X1 U15296 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16617), .ZN(n16616) );
  INV_X1 U15297 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16982) );
  NAND2_X1 U15298 ( .A1(n16616), .A2(n16982), .ZN(n16611) );
  NOR2_X1 U15299 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16611), .ZN(n16595) );
  INV_X1 U15300 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16944) );
  NAND2_X1 U15301 ( .A1(n16595), .A2(n16944), .ZN(n16572) );
  NOR2_X1 U15302 ( .A1(n16933), .A2(n16572), .ZN(n16579) );
  INV_X1 U15303 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n12148) );
  NOR2_X1 U15304 ( .A1(n16885), .A2(n9894), .ZN(n12147) );
  NAND3_X1 U15305 ( .A1(n12140), .A2(n12150), .A3(n12149), .ZN(n12151) );
  AND3_X1 U15306 ( .A1(n20914), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n12153) );
  NOR2_X1 U15307 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n12248) );
  NAND2_X1 U15308 ( .A1(n12153), .A2(n20783), .ZN(n16049) );
  INV_X1 U15309 ( .A(n12214), .ZN(n12176) );
  NAND2_X1 U15310 ( .A1(n13632), .A2(n20267), .ZN(n12166) );
  OAI21_X1 U15311 ( .B1(n13246), .B2(n12157), .A(n12166), .ZN(n12154) );
  INV_X1 U15312 ( .A(n12154), .ZN(n12155) );
  NAND2_X1 U15313 ( .A1(n12156), .A2(n20258), .ZN(n12162) );
  NAND2_X1 U15314 ( .A1(n12157), .A2(n12158), .ZN(n12174) );
  OAI21_X1 U15315 ( .B1(n12158), .B2(n12157), .A(n12174), .ZN(n12159) );
  OAI211_X1 U15316 ( .C1(n12159), .C2(n13246), .A(n10299), .B(n14160), .ZN(
        n12160) );
  INV_X1 U15317 ( .A(n12160), .ZN(n12161) );
  NAND2_X1 U15318 ( .A1(n12162), .A2(n12161), .ZN(n12164) );
  NAND2_X1 U15319 ( .A1(n13286), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20221) );
  INV_X1 U15320 ( .A(n12163), .ZN(n13062) );
  NAND2_X1 U15321 ( .A1(n13062), .A2(n12164), .ZN(n12165) );
  INV_X1 U15322 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20204) );
  OR2_X1 U15323 ( .A1(n20240), .A2(n12176), .ZN(n12170) );
  XNOR2_X1 U15324 ( .A(n12174), .B(n12173), .ZN(n12168) );
  INV_X1 U15325 ( .A(n12166), .ZN(n12167) );
  AOI21_X1 U15326 ( .B1(n12168), .B2(n20910), .A(n12167), .ZN(n12169) );
  NAND2_X1 U15327 ( .A1(n12170), .A2(n12169), .ZN(n13292) );
  NAND2_X1 U15328 ( .A1(n13293), .A2(n13292), .ZN(n13291) );
  NAND2_X1 U15329 ( .A1(n12171), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12172) );
  NAND2_X1 U15330 ( .A1(n13291), .A2(n12172), .ZN(n13370) );
  NAND2_X1 U15331 ( .A1(n12174), .A2(n12173), .ZN(n12181) );
  XNOR2_X1 U15332 ( .A(n12181), .B(n12180), .ZN(n12175) );
  XNOR2_X1 U15333 ( .A(n12177), .B(n20197), .ZN(n13371) );
  NAND2_X1 U15334 ( .A1(n13370), .A2(n13371), .ZN(n13369) );
  NAND2_X1 U15335 ( .A1(n9644), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12178) );
  NAND2_X1 U15336 ( .A1(n13369), .A2(n12178), .ZN(n20171) );
  NAND2_X1 U15337 ( .A1(n12179), .A2(n12214), .ZN(n12184) );
  NAND2_X1 U15338 ( .A1(n12181), .A2(n12180), .ZN(n12190) );
  XNOR2_X1 U15339 ( .A(n12190), .B(n12188), .ZN(n12182) );
  NAND2_X1 U15340 ( .A1(n12182), .A2(n20910), .ZN(n12183) );
  NAND2_X1 U15341 ( .A1(n12184), .A2(n12183), .ZN(n12185) );
  XNOR2_X1 U15342 ( .A(n12185), .B(n20188), .ZN(n20170) );
  NAND2_X1 U15343 ( .A1(n20171), .A2(n20170), .ZN(n20169) );
  NAND2_X1 U15344 ( .A1(n12185), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12186) );
  NAND2_X1 U15345 ( .A1(n20169), .A2(n12186), .ZN(n16075) );
  NAND2_X1 U15346 ( .A1(n12187), .A2(n12214), .ZN(n12193) );
  INV_X1 U15347 ( .A(n12188), .ZN(n12189) );
  OR2_X1 U15348 ( .A1(n12190), .A2(n12189), .ZN(n12197) );
  XNOR2_X1 U15349 ( .A(n12197), .B(n12198), .ZN(n12191) );
  NAND2_X1 U15350 ( .A1(n12191), .A2(n20910), .ZN(n12192) );
  NAND2_X1 U15351 ( .A1(n12193), .A2(n12192), .ZN(n12194) );
  XNOR2_X1 U15352 ( .A(n12194), .B(n16169), .ZN(n16074) );
  NAND2_X1 U15353 ( .A1(n16075), .A2(n16074), .ZN(n16073) );
  NAND2_X1 U15354 ( .A1(n12194), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12195) );
  NAND2_X1 U15355 ( .A1(n16073), .A2(n12195), .ZN(n16069) );
  NAND2_X1 U15356 ( .A1(n12196), .A2(n12214), .ZN(n12202) );
  INV_X1 U15357 ( .A(n12197), .ZN(n12199) );
  NAND2_X1 U15358 ( .A1(n12199), .A2(n12198), .ZN(n12206) );
  XNOR2_X1 U15359 ( .A(n12206), .B(n12207), .ZN(n12200) );
  NAND2_X1 U15360 ( .A1(n12200), .A2(n20910), .ZN(n12201) );
  NAND2_X1 U15361 ( .A1(n12202), .A2(n12201), .ZN(n12203) );
  XNOR2_X1 U15362 ( .A(n12203), .B(n16148), .ZN(n16068) );
  NAND2_X1 U15363 ( .A1(n16069), .A2(n16068), .ZN(n16067) );
  NAND2_X1 U15364 ( .A1(n12203), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12204) );
  NAND2_X1 U15365 ( .A1(n12205), .A2(n12214), .ZN(n12211) );
  INV_X1 U15366 ( .A(n12206), .ZN(n12208) );
  NAND2_X1 U15367 ( .A1(n12208), .A2(n12207), .ZN(n12221) );
  XNOR2_X1 U15368 ( .A(n12221), .B(n12219), .ZN(n12209) );
  NAND2_X1 U15369 ( .A1(n12209), .A2(n20910), .ZN(n12210) );
  NAND2_X1 U15370 ( .A1(n12211), .A2(n12210), .ZN(n16062) );
  OR2_X1 U15371 ( .A1(n16062), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12212) );
  NAND2_X1 U15372 ( .A1(n16062), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12213) );
  NAND2_X1 U15373 ( .A1(n12214), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12216) );
  NOR2_X1 U15374 ( .A1(n12216), .A2(n12215), .ZN(n12217) );
  NAND2_X1 U15375 ( .A1(n20910), .A2(n12219), .ZN(n12220) );
  OR2_X1 U15376 ( .A1(n12221), .A2(n12220), .ZN(n12222) );
  NAND2_X1 U15377 ( .A1(n9673), .A2(n12222), .ZN(n13797) );
  AND2_X1 U15378 ( .A1(n13797), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12223) );
  NAND2_X1 U15379 ( .A1(n12224), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12225) );
  NAND2_X1 U15380 ( .A1(n14972), .A2(n16139), .ZN(n12226) );
  XNOR2_X1 U15381 ( .A(n9672), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14995) );
  INV_X1 U15382 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12227) );
  NAND2_X1 U15383 ( .A1(n9672), .A2(n12227), .ZN(n14992) );
  NAND2_X1 U15384 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12228) );
  NAND2_X1 U15385 ( .A1(n9673), .A2(n12228), .ZN(n14010) );
  AND2_X1 U15386 ( .A1(n14992), .A2(n14010), .ZN(n12229) );
  INV_X1 U15387 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12230) );
  NAND2_X1 U15388 ( .A1(n16114), .A2(n12230), .ZN(n12231) );
  NAND2_X1 U15389 ( .A1(n12224), .A2(n12231), .ZN(n12234) );
  XNOR2_X1 U15390 ( .A(n9672), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14033) );
  NAND2_X1 U15391 ( .A1(n9673), .A2(n14042), .ZN(n14980) );
  NAND2_X1 U15392 ( .A1(n14033), .A2(n14980), .ZN(n12232) );
  AOI21_X1 U15393 ( .B1(n14031), .B2(n12234), .A(n12232), .ZN(n14967) );
  OAI21_X1 U15394 ( .B1(n12224), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n14967), .ZN(n12238) );
  INV_X1 U15395 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16133) );
  NAND2_X1 U15396 ( .A1(n16133), .A2(n16116), .ZN(n12233) );
  NAND2_X1 U15397 ( .A1(n12224), .A2(n12233), .ZN(n14011) );
  NAND2_X1 U15398 ( .A1(n12224), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14013) );
  NAND2_X1 U15399 ( .A1(n14011), .A2(n14013), .ZN(n16038) );
  INV_X1 U15400 ( .A(n12234), .ZN(n12235) );
  NOR2_X1 U15401 ( .A1(n14972), .A2(n14042), .ZN(n14982) );
  NOR2_X1 U15402 ( .A1(n14983), .A2(n14982), .ZN(n14032) );
  OAI21_X1 U15403 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(n12224), .ZN(n12236) );
  XNOR2_X1 U15404 ( .A(n14972), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14963) );
  NAND2_X1 U15405 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15105) );
  NAND2_X1 U15406 ( .A1(n14922), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12241) );
  NAND2_X1 U15407 ( .A1(n15123), .A2(n15138), .ZN(n12240) );
  INV_X1 U15408 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14905) );
  NAND4_X2 U15409 ( .A1(n14914), .A2(n15068), .A3(n14905), .A4(n15092), .ZN(
        n14883) );
  NAND2_X1 U15410 ( .A1(n12241), .A2(n14972), .ZN(n14892) );
  NOR2_X1 U15411 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15045) );
  AND2_X1 U15412 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15044) );
  NAND3_X1 U15413 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15061) );
  INV_X1 U15414 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15037) );
  NAND2_X1 U15415 ( .A1(n12224), .A2(n15037), .ZN(n14857) );
  INV_X1 U15416 ( .A(n14874), .ZN(n12244) );
  NAND2_X1 U15417 ( .A1(n14972), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14149) );
  INV_X1 U15418 ( .A(n15044), .ZN(n15011) );
  OR2_X1 U15419 ( .A1(n14149), .A2(n15011), .ZN(n12243) );
  INV_X1 U15420 ( .A(n12245), .ZN(n13171) );
  NAND2_X1 U15421 ( .A1(n10306), .A2(n13632), .ZN(n12246) );
  NAND3_X1 U15422 ( .A1(n13171), .A2(n10299), .A3(n12246), .ZN(n13189) );
  OR2_X1 U15423 ( .A1(n13189), .A2(n12247), .ZN(n14472) );
  INV_X1 U15424 ( .A(n20000), .ZN(n13227) );
  INV_X1 U15425 ( .A(n12248), .ZN(n20781) );
  NAND2_X1 U15426 ( .A1(n20781), .A2(n12250), .ZN(n20917) );
  NAND2_X1 U15427 ( .A1(n20917), .A2(n20914), .ZN(n12249) );
  INV_X2 U15428 ( .A(n13067), .ZN(n20168) );
  OR2_X1 U15429 ( .A1(n12250), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20064) );
  INV_X1 U15430 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21032) );
  NOR2_X1 U15431 ( .A1(n20225), .A2(n21032), .ZN(n15020) );
  NAND2_X1 U15432 ( .A1(n20914), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12252) );
  NAND2_X1 U15433 ( .A1(n21034), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12251) );
  AND2_X1 U15434 ( .A1(n12252), .A2(n12251), .ZN(n13066) );
  OR2_X2 U15435 ( .A1(n20168), .A2(n13066), .ZN(n20178) );
  INV_X1 U15436 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12254) );
  INV_X1 U15437 ( .A(n13641), .ZN(n12256) );
  NOR2_X1 U15438 ( .A1(n20178), .A2(n12256), .ZN(n12257) );
  AOI211_X1 U15439 ( .C1(n20168), .C2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15020), .B(n12257), .ZN(n12258) );
  OR2_X1 U15440 ( .A1(n16363), .A2(n11551), .ZN(n13024) );
  INV_X1 U15441 ( .A(n13024), .ZN(n12261) );
  NOR2_X1 U15442 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19863) );
  AOI211_X1 U15443 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n19863), .ZN(n19988) );
  INV_X1 U15444 ( .A(n19988), .ZN(n19859) );
  NAND2_X1 U15445 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19985) );
  INV_X1 U15446 ( .A(n19985), .ZN(n19867) );
  NOR2_X1 U15447 ( .A1(n19859), .A2(n19867), .ZN(n12914) );
  NAND2_X1 U15448 ( .A1(n12261), .A2(n12914), .ZN(n13749) );
  INV_X1 U15449 ( .A(n16357), .ZN(n12904) );
  NAND2_X1 U15450 ( .A1(n11551), .A2(n12917), .ZN(n12262) );
  AOI21_X1 U15451 ( .B1(n13749), .B2(n12262), .A(n11413), .ZN(n12282) );
  OAI211_X1 U15452 ( .C1(n12263), .C2(n11388), .A(n13024), .B(n11387), .ZN(
        n12280) );
  NAND2_X1 U15453 ( .A1(n12266), .A2(n11387), .ZN(n12267) );
  NAND2_X1 U15454 ( .A1(n12267), .A2(n11413), .ZN(n12268) );
  NAND2_X1 U15455 ( .A1(n12265), .A2(n12268), .ZN(n12275) );
  NAND2_X1 U15456 ( .A1(n11387), .A2(n11551), .ZN(n12512) );
  NAND2_X1 U15457 ( .A1(n12512), .A2(n16366), .ZN(n12269) );
  NAND2_X1 U15458 ( .A1(n12269), .A2(n19288), .ZN(n12270) );
  AOI21_X1 U15459 ( .B1(n12270), .B2(n11413), .A(n12525), .ZN(n12274) );
  NAND2_X1 U15460 ( .A1(n12271), .A2(n19288), .ZN(n12272) );
  NAND2_X1 U15461 ( .A1(n12272), .A2(n19970), .ZN(n12522) );
  NAND4_X1 U15462 ( .A1(n12275), .A2(n12274), .A3(n12522), .A4(n12273), .ZN(
        n12513) );
  INV_X1 U15463 ( .A(n12914), .ZN(n12276) );
  NOR2_X1 U15464 ( .A1(n16357), .A2(n12276), .ZN(n12277) );
  AND2_X1 U15465 ( .A1(n16386), .A2(n12277), .ZN(n12278) );
  NOR2_X1 U15466 ( .A1(n12513), .A2(n12278), .ZN(n13752) );
  NAND3_X1 U15467 ( .A1(n16386), .A2(n19989), .A3(n12917), .ZN(n12279) );
  NAND3_X1 U15468 ( .A1(n12280), .A2(n13752), .A3(n12279), .ZN(n12281) );
  OAI21_X1 U15469 ( .B1(n12282), .B2(n12281), .A(n13262), .ZN(n12285) );
  INV_X1 U15470 ( .A(n12283), .ZN(n12284) );
  NAND2_X2 U15471 ( .A1(n12285), .A2(n12284), .ZN(n12554) );
  NOR2_X1 U15472 ( .A1(n11397), .A2(n12811), .ZN(n12286) );
  NAND2_X2 U15473 ( .A1(n12554), .A2(n12286), .ZN(n16320) );
  AOI21_X1 U15474 ( .B1(n12287), .B2(n14203), .A(n14188), .ZN(n15393) );
  NOR2_X1 U15475 ( .A1(n11397), .A2(n12288), .ZN(n12289) );
  AND2_X2 U15476 ( .A1(n12554), .A2(n12289), .ZN(n16328) );
  NAND2_X1 U15477 ( .A1(n12290), .A2(n14168), .ZN(n12310) );
  NAND2_X1 U15478 ( .A1(n12473), .A2(n12292), .ZN(n12294) );
  MUX2_X1 U15479 ( .A(n19288), .B(n19966), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12293) );
  NAND3_X1 U15480 ( .A1(n12310), .A2(n12294), .A3(n12293), .ZN(n13074) );
  INV_X1 U15481 ( .A(n12295), .ZN(n12296) );
  NAND2_X1 U15482 ( .A1(n12314), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12299) );
  INV_X1 U15483 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13020) );
  OAI21_X1 U15484 ( .B1(n19288), .B2(n13020), .A(n19645), .ZN(n12297) );
  AOI21_X1 U15485 ( .B1(n14168), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12297), .ZN(n12298) );
  NAND2_X1 U15486 ( .A1(n12299), .A2(n12298), .ZN(n13073) );
  NAND2_X1 U15487 ( .A1(n12314), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12301) );
  AOI22_X1 U15488 ( .A1(n12503), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n14168), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12300) );
  NAND2_X1 U15489 ( .A1(n12301), .A2(n12300), .ZN(n12306) );
  OR2_X1 U15490 ( .A1(n12302), .A2(n12336), .ZN(n12305) );
  NAND2_X1 U15491 ( .A1(n12266), .A2(n19288), .ZN(n12303) );
  MUX2_X1 U15492 ( .A(n12303), .B(n19956), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12304) );
  NAND2_X1 U15493 ( .A1(n12305), .A2(n12304), .ZN(n13049) );
  NOR2_X1 U15494 ( .A1(n13050), .A2(n13049), .ZN(n12308) );
  NOR2_X1 U15495 ( .A1(n13076), .A2(n12306), .ZN(n12307) );
  NOR2_X2 U15496 ( .A1(n12308), .A2(n12307), .ZN(n12313) );
  NAND2_X1 U15497 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12309) );
  OAI211_X1 U15498 ( .C1(n12336), .C2(n12311), .A(n12310), .B(n12309), .ZN(
        n12312) );
  NOR2_X1 U15499 ( .A1(n12313), .A2(n12312), .ZN(n12318) );
  XNOR2_X1 U15500 ( .A(n12313), .B(n12312), .ZN(n13144) );
  NAND2_X1 U15501 ( .A1(n12314), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U15502 ( .A1(n12503), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n14168), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12316) );
  NAND2_X1 U15503 ( .A1(n12317), .A2(n12316), .ZN(n13143) );
  NOR2_X1 U15504 ( .A1(n13144), .A2(n13143), .ZN(n13145) );
  NAND2_X1 U15505 ( .A1(n12314), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12323) );
  NAND2_X1 U15506 ( .A1(n12473), .A2(n12319), .ZN(n12322) );
  AOI22_X1 U15507 ( .A1(n14168), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12321) );
  NAND2_X1 U15508 ( .A1(n12503), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12320) );
  NAND2_X1 U15509 ( .A1(n12314), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12327) );
  NAND2_X1 U15510 ( .A1(n12473), .A2(n12324), .ZN(n12326) );
  AOI22_X1 U15511 ( .A1(n12503), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n14168), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12325) );
  INV_X1 U15512 ( .A(n12328), .ZN(n12329) );
  AOI22_X1 U15513 ( .A1(n12314), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n12329), 
        .B2(n12974), .ZN(n12331) );
  AOI22_X1 U15514 ( .A1(n12315), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n14168), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12330) );
  NAND2_X1 U15515 ( .A1(n12331), .A2(n12330), .ZN(n13784) );
  NAND2_X1 U15516 ( .A1(n12473), .A2(n12332), .ZN(n13267) );
  NAND2_X1 U15517 ( .A1(n13783), .A2(n13267), .ZN(n12335) );
  NAND2_X1 U15518 ( .A1(n12314), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12334) );
  AOI22_X1 U15519 ( .A1(n12315), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n14168), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12333) );
  NAND2_X1 U15520 ( .A1(n12334), .A2(n12333), .ZN(n13266) );
  NAND2_X1 U15521 ( .A1(n12335), .A2(n13266), .ZN(n13270) );
  NAND2_X1 U15522 ( .A1(n12314), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U15523 ( .A1(n12315), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n14168), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12337) );
  NAND2_X1 U15524 ( .A1(n12338), .A2(n12337), .ZN(n13257) );
  NAND2_X1 U15525 ( .A1(n12314), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12354) );
  AOI22_X1 U15526 ( .A1(n12466), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11531), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12343) );
  AOI22_X1 U15527 ( .A1(n11288), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12342) );
  INV_X1 U15528 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13830) );
  OAI22_X1 U15529 ( .A1(n14290), .A2(n13830), .B1(n14289), .B2(n19256), .ZN(
        n12339) );
  INV_X1 U15530 ( .A(n12339), .ZN(n12341) );
  AOI22_X1 U15531 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14293), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12340) );
  NAND4_X1 U15532 ( .A1(n12343), .A2(n12342), .A3(n12341), .A4(n12340), .ZN(
        n12351) );
  AOI22_X1 U15533 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11530), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12349) );
  INV_X1 U15534 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12344) );
  INV_X1 U15535 ( .A(n14245), .ZN(n12415) );
  INV_X1 U15536 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13831) );
  OAI22_X1 U15537 ( .A1(n12408), .A2(n12344), .B1(n12415), .B2(n13831), .ZN(
        n12345) );
  INV_X1 U15538 ( .A(n12345), .ZN(n12348) );
  AOI22_X1 U15539 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U15540 ( .A1(n14301), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12346) );
  NAND4_X1 U15541 ( .A1(n12349), .A2(n12348), .A3(n12347), .A4(n12346), .ZN(
        n12350) );
  NAND2_X1 U15542 ( .A1(n12473), .A2(n13348), .ZN(n12353) );
  AOI22_X1 U15543 ( .A1(n12315), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n14168), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12352) );
  AOI22_X1 U15544 ( .A1(n12314), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n12315), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n12370) );
  AOI22_X1 U15545 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11288), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12359) );
  INV_X1 U15546 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13875) );
  OAI22_X1 U15547 ( .A1(n13875), .A2(n14290), .B1(n14289), .B2(n19259), .ZN(
        n12355) );
  INV_X1 U15548 ( .A(n12355), .ZN(n12358) );
  AOI22_X1 U15549 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14293), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12357) );
  AOI22_X1 U15550 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11531), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12356) );
  NAND4_X1 U15551 ( .A1(n12359), .A2(n12358), .A3(n12357), .A4(n12356), .ZN(
        n12368) );
  AOI22_X1 U15552 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n14300), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12366) );
  AOI22_X1 U15553 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14301), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12365) );
  INV_X1 U15554 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12361) );
  OAI22_X1 U15555 ( .A1(n14305), .A2(n12361), .B1(n14303), .B2(n12360), .ZN(
        n12362) );
  INV_X1 U15556 ( .A(n12362), .ZN(n12364) );
  AOI22_X1 U15557 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n14307), .ZN(n12363) );
  NAND4_X1 U15558 ( .A1(n12366), .A2(n12365), .A3(n12364), .A4(n12363), .ZN(
        n12367) );
  AOI22_X1 U15559 ( .A1(n12473), .A2(n13354), .B1(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n14168), .ZN(n12369) );
  NAND2_X1 U15560 ( .A1(n12370), .A2(n12369), .ZN(n13276) );
  AOI22_X1 U15561 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14293), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12374) );
  AOI22_X1 U15562 ( .A1(n12459), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12373) );
  AOI22_X1 U15563 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11288), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12372) );
  AOI22_X1 U15564 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n14300), .B1(
        n11531), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12371) );
  NAND4_X1 U15565 ( .A1(n12374), .A2(n12373), .A3(n12372), .A4(n12371), .ZN(
        n12386) );
  AOI22_X1 U15566 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12384) );
  AOI22_X1 U15567 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12383) );
  INV_X1 U15568 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12375) );
  INV_X1 U15569 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13907) );
  OAI22_X1 U15570 ( .A1(n14305), .A2(n12375), .B1(n13907), .B2(n12415), .ZN(
        n12376) );
  INV_X1 U15571 ( .A(n12376), .ZN(n12382) );
  INV_X1 U15572 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12377) );
  OAI22_X1 U15573 ( .A1(n12379), .A2(n14303), .B1(n12378), .B2(n12377), .ZN(
        n12380) );
  INV_X1 U15574 ( .A(n12380), .ZN(n12381) );
  NAND4_X1 U15575 ( .A1(n12384), .A2(n12383), .A3(n12382), .A4(n12381), .ZN(
        n12385) );
  NOR2_X1 U15576 ( .A1(n12386), .A2(n12385), .ZN(n13510) );
  INV_X1 U15577 ( .A(n13510), .ZN(n12389) );
  AOI22_X1 U15578 ( .A1(n12315), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12387) );
  OAI21_X1 U15579 ( .B1(n12476), .B2(n13578), .A(n12387), .ZN(n12388) );
  AOI21_X1 U15580 ( .B1(n12473), .B2(n12389), .A(n12388), .ZN(n13572) );
  NAND2_X1 U15581 ( .A1(n12314), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12406) );
  AOI22_X1 U15582 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n11288), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12394) );
  INV_X1 U15583 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13969) );
  OAI22_X1 U15584 ( .A1(n13969), .A2(n14290), .B1(n14289), .B2(n19269), .ZN(
        n12390) );
  INV_X1 U15585 ( .A(n12390), .ZN(n12393) );
  AOI22_X1 U15586 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14293), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12392) );
  AOI22_X1 U15587 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n11531), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12391) );
  NAND4_X1 U15588 ( .A1(n12394), .A2(n12393), .A3(n12392), .A4(n12391), .ZN(
        n12403) );
  AOI22_X1 U15589 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n14300), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12401) );
  AOI22_X1 U15590 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14301), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12400) );
  INV_X1 U15591 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12396) );
  OAI22_X1 U15592 ( .A1(n14305), .A2(n12396), .B1(n14303), .B2(n12395), .ZN(
        n12397) );
  INV_X1 U15593 ( .A(n12397), .ZN(n12399) );
  AOI22_X1 U15594 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n14307), .ZN(n12398) );
  NAND4_X1 U15595 ( .A1(n12401), .A2(n12400), .A3(n12399), .A4(n12398), .ZN(
        n12402) );
  NAND2_X1 U15596 ( .A1(n12473), .A2(n13620), .ZN(n12405) );
  AOI22_X1 U15597 ( .A1(n12315), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12404) );
  NAND3_X1 U15598 ( .A1(n12406), .A2(n12405), .A3(n12404), .ZN(n13278) );
  AOI22_X1 U15599 ( .A1(n12459), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11288), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U15600 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12413) );
  AOI22_X1 U15601 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14293), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12412) );
  INV_X1 U15602 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12409) );
  INV_X1 U15603 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12407) );
  OAI22_X1 U15604 ( .A1(n12409), .A2(n12408), .B1(n14303), .B2(n12407), .ZN(
        n12410) );
  INV_X1 U15605 ( .A(n12410), .ZN(n12411) );
  NAND4_X1 U15606 ( .A1(n12414), .A2(n12413), .A3(n12412), .A4(n12411), .ZN(
        n12423) );
  AOI22_X1 U15607 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11531), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U15608 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12420) );
  AOI22_X1 U15609 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n14301), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12419) );
  INV_X1 U15610 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12416) );
  INV_X1 U15611 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14237) );
  OAI22_X1 U15612 ( .A1(n14305), .A2(n12416), .B1(n14237), .B2(n12415), .ZN(
        n12417) );
  INV_X1 U15613 ( .A(n12417), .ZN(n12418) );
  NAND4_X1 U15614 ( .A1(n12421), .A2(n12420), .A3(n12419), .A4(n12418), .ZN(
        n12422) );
  AOI22_X1 U15615 ( .A1(n12315), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12424) );
  OAI21_X1 U15616 ( .B1(n12476), .B2(n12425), .A(n12424), .ZN(n12426) );
  AOI21_X1 U15617 ( .B1(n12473), .B2(n13667), .A(n12426), .ZN(n15784) );
  AOI22_X1 U15618 ( .A1(n12314), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n12315), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n12442) );
  AOI22_X1 U15619 ( .A1(n11288), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12431) );
  INV_X1 U15620 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14221) );
  INV_X1 U15621 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13216) );
  OAI22_X1 U15622 ( .A1(n14290), .A2(n14221), .B1(n14289), .B2(n13216), .ZN(
        n12427) );
  INV_X1 U15623 ( .A(n12427), .ZN(n12430) );
  AOI22_X1 U15624 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14293), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12429) );
  AOI22_X1 U15625 ( .A1(n11531), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12428) );
  NAND4_X1 U15626 ( .A1(n12431), .A2(n12430), .A3(n12429), .A4(n12428), .ZN(
        n12440) );
  AOI22_X1 U15627 ( .A1(n14300), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U15628 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14301), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12437) );
  INV_X1 U15629 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12433) );
  INV_X1 U15630 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12432) );
  OAI22_X1 U15631 ( .A1(n14305), .A2(n12433), .B1(n14303), .B2(n12432), .ZN(
        n12434) );
  INV_X1 U15632 ( .A(n12434), .ZN(n12436) );
  AOI22_X1 U15633 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14307), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12435) );
  NAND4_X1 U15634 ( .A1(n12438), .A2(n12437), .A3(n12436), .A4(n12435), .ZN(
        n12439) );
  AOI22_X1 U15635 ( .A1(n12473), .A2(n13709), .B1(n14168), .B2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12441) );
  NAND2_X1 U15636 ( .A1(n12442), .A2(n12441), .ZN(n13506) );
  NAND2_X1 U15637 ( .A1(n12314), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U15638 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n14287), .B1(
        n11288), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12446) );
  AOI22_X1 U15639 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12459), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12445) );
  AOI22_X1 U15640 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n14293), .B1(
        n14294), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12444) );
  AOI22_X1 U15641 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n11531), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12443) );
  NAND4_X1 U15642 ( .A1(n12446), .A2(n12445), .A3(n12444), .A4(n12443), .ZN(
        n12455) );
  AOI22_X1 U15643 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n14245), .ZN(n12453) );
  AOI22_X1 U15644 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14299), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12452) );
  INV_X1 U15645 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12447) );
  OAI22_X1 U15646 ( .A1(n14305), .A2(n12448), .B1(n14303), .B2(n12447), .ZN(
        n12449) );
  INV_X1 U15647 ( .A(n12449), .ZN(n12451) );
  AOI22_X1 U15648 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14301), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12450) );
  NAND4_X1 U15649 ( .A1(n12453), .A2(n12452), .A3(n12451), .A4(n12450), .ZN(
        n12454) );
  OR2_X1 U15650 ( .A1(n12455), .A2(n12454), .ZN(n13710) );
  NAND2_X1 U15651 ( .A1(n12473), .A2(n13710), .ZN(n12457) );
  AOI22_X1 U15652 ( .A1(n12315), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12456) );
  AOI22_X1 U15653 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n11288), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U15654 ( .A1(n12460), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12459), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12463) );
  AOI22_X1 U15655 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n14293), .B1(
        n14294), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12462) );
  AOI22_X1 U15656 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n11531), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12461) );
  NAND4_X1 U15657 ( .A1(n12464), .A2(n12463), .A3(n12462), .A4(n12461), .ZN(
        n12472) );
  AOI22_X1 U15658 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n14307), .ZN(n12470) );
  AOI22_X1 U15659 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14299), .B1(
        n14300), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12469) );
  AOI22_X1 U15660 ( .A1(n12466), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12465), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12468) );
  AOI22_X1 U15661 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14301), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12467) );
  NAND4_X1 U15662 ( .A1(n12470), .A2(n12469), .A3(n12468), .A4(n12467), .ZN(
        n12471) );
  NAND2_X1 U15663 ( .A1(n12473), .A2(n13819), .ZN(n12475) );
  AOI22_X1 U15664 ( .A1(n12503), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12474) );
  OAI211_X1 U15665 ( .C1(n12476), .C2(n19888), .A(n12475), .B(n12474), .ZN(
        n12859) );
  NAND2_X1 U15666 ( .A1(n12314), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U15667 ( .A1(n12503), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12477) );
  AND2_X1 U15668 ( .A1(n12478), .A2(n12477), .ZN(n13861) );
  NAND2_X1 U15669 ( .A1(n12314), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12480) );
  AOI22_X1 U15670 ( .A1(n12503), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12479) );
  NAND2_X1 U15671 ( .A1(n12314), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U15672 ( .A1(n12503), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12481) );
  NAND2_X1 U15673 ( .A1(n12482), .A2(n12481), .ZN(n15219) );
  NAND2_X1 U15674 ( .A1(n12314), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12484) );
  AOI22_X1 U15675 ( .A1(n12503), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12483) );
  NAND2_X1 U15676 ( .A1(n12484), .A2(n12483), .ZN(n13991) );
  NAND2_X1 U15677 ( .A1(n12314), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12486) );
  AOI22_X1 U15678 ( .A1(n12503), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12485) );
  AND2_X1 U15679 ( .A1(n12486), .A2(n12485), .ZN(n15664) );
  NAND2_X1 U15680 ( .A1(n12314), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12488) );
  AOI22_X1 U15681 ( .A1(n12503), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12487) );
  AND2_X1 U15682 ( .A1(n12488), .A2(n12487), .ZN(n15378) );
  NAND2_X1 U15683 ( .A1(n12314), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12490) );
  AOI22_X1 U15684 ( .A1(n12503), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12489) );
  AND2_X1 U15685 ( .A1(n12490), .A2(n12489), .ZN(n12897) );
  NAND2_X1 U15686 ( .A1(n12314), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12492) );
  AOI22_X1 U15687 ( .A1(n12503), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12491) );
  NAND2_X1 U15688 ( .A1(n12492), .A2(n12491), .ZN(n12870) );
  NAND2_X1 U15689 ( .A1(n12314), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12494) );
  AOI22_X1 U15690 ( .A1(n12503), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12493) );
  AND2_X1 U15691 ( .A1(n12494), .A2(n12493), .ZN(n15353) );
  NAND2_X1 U15692 ( .A1(n12314), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12496) );
  AOI22_X1 U15693 ( .A1(n12503), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12495) );
  AND2_X1 U15694 ( .A1(n12496), .A2(n12495), .ZN(n15203) );
  NAND2_X1 U15695 ( .A1(n12314), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12498) );
  AOI22_X1 U15696 ( .A1(n12503), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12497) );
  NAND2_X1 U15697 ( .A1(n12498), .A2(n12497), .ZN(n15336) );
  NAND2_X1 U15698 ( .A1(n12314), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12500) );
  AOI22_X1 U15699 ( .A1(n12503), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12499) );
  NAND2_X1 U15700 ( .A1(n12500), .A2(n12499), .ZN(n12882) );
  NAND2_X1 U15701 ( .A1(n12314), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12502) );
  AOI22_X1 U15702 ( .A1(n12503), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12501) );
  AND2_X1 U15703 ( .A1(n12502), .A2(n12501), .ZN(n15189) );
  NAND2_X1 U15704 ( .A1(n12314), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12505) );
  AOI22_X1 U15705 ( .A1(n12503), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n14168), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12504) );
  NAND2_X1 U15706 ( .A1(n9716), .A2(n9764), .ZN(n12506) );
  NAND2_X1 U15707 ( .A1(n12805), .A2(n12506), .ZN(n16203) );
  AND2_X1 U15708 ( .A1(n12508), .A2(n12507), .ZN(n15835) );
  NOR2_X1 U15709 ( .A1(n12509), .A2(n11551), .ZN(n12510) );
  OR2_X1 U15710 ( .A1(n15835), .A2(n12510), .ZN(n12511) );
  INV_X1 U15711 ( .A(n15836), .ZN(n16359) );
  NAND2_X1 U15712 ( .A1(n12554), .A2(n16359), .ZN(n13149) );
  AND2_X1 U15713 ( .A1(n12514), .A2(n12524), .ZN(n13263) );
  OAI22_X1 U15714 ( .A1(n12913), .A2(n12516), .B1(n16366), .B2(n11413), .ZN(
        n12517) );
  INV_X1 U15715 ( .A(n12517), .ZN(n12518) );
  NAND2_X1 U15716 ( .A1(n12519), .A2(n12518), .ZN(n12520) );
  NOR2_X1 U15717 ( .A1(n13263), .A2(n12520), .ZN(n12529) );
  NAND2_X1 U15718 ( .A1(n12521), .A2(n19989), .ZN(n13759) );
  NAND2_X1 U15719 ( .A1(n13759), .A2(n12522), .ZN(n12523) );
  NAND2_X1 U15720 ( .A1(n12523), .A2(n19265), .ZN(n12528) );
  OAI21_X1 U15721 ( .B1(n12524), .B2(n10155), .A(n12913), .ZN(n12526) );
  NAND2_X1 U15722 ( .A1(n12526), .A2(n12525), .ZN(n12527) );
  AND3_X1 U15723 ( .A1(n12529), .A2(n12528), .A3(n12527), .ZN(n15840) );
  NAND2_X1 U15724 ( .A1(n15840), .A2(n9732), .ZN(n12530) );
  NAND2_X1 U15725 ( .A1(n12554), .A2(n12530), .ZN(n15706) );
  NAND2_X2 U15726 ( .A1(n13149), .A2(n15706), .ZN(n15798) );
  INV_X1 U15727 ( .A(n13149), .ZN(n15705) );
  NAND2_X1 U15728 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13051) );
  NOR2_X1 U15729 ( .A1(n13141), .A2(n13051), .ZN(n13147) );
  NAND2_X1 U15730 ( .A1(n13141), .A2(n13051), .ZN(n13161) );
  OAI21_X1 U15731 ( .B1(n15705), .B2(n13147), .A(n13161), .ZN(n13499) );
  NOR3_X2 U15732 ( .A1(n15710), .A2(n13500), .A3(n13499), .ZN(n13957) );
  INV_X1 U15733 ( .A(n13957), .ZN(n13787) );
  INV_X1 U15734 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16323) );
  NOR2_X1 U15735 ( .A1(n13789), .A2(n13788), .ZN(n13956) );
  NAND2_X1 U15736 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13956), .ZN(
        n13929) );
  OR3_X1 U15737 ( .A1(n16323), .A2(n16336), .A3(n13929), .ZN(n12531) );
  NAND3_X1 U15738 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12534) );
  NOR2_X2 U15739 ( .A1(n15797), .A2(n12534), .ZN(n15766) );
  AND2_X1 U15740 ( .A1(n15754), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12536) );
  NAND2_X1 U15741 ( .A1(n15766), .A2(n12536), .ZN(n15731) );
  AND3_X1 U15742 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15697) );
  NAND2_X1 U15743 ( .A1(n15697), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12539) );
  NOR2_X2 U15744 ( .A1(n15731), .A2(n12539), .ZN(n15685) );
  AND2_X1 U15745 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12541) );
  NAND2_X1 U15746 ( .A1(n15685), .A2(n12541), .ZN(n15653) );
  NAND2_X1 U15747 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15626) );
  OR2_X2 U15748 ( .A1(n15648), .A2(n15626), .ZN(n15614) );
  NOR2_X2 U15749 ( .A1(n15614), .A2(n15619), .ZN(n15608) );
  NOR2_X1 U15750 ( .A1(n15607), .A2(n15414), .ZN(n12546) );
  NAND2_X1 U15751 ( .A1(n15608), .A2(n12546), .ZN(n15570) );
  OR2_X1 U15752 ( .A1(n15570), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15584) );
  INV_X1 U15753 ( .A(n13161), .ZN(n13497) );
  OR3_X1 U15754 ( .A1(n13497), .A2(n13500), .A3(n12531), .ZN(n12532) );
  AND2_X1 U15755 ( .A1(n15798), .A2(n12532), .ZN(n12533) );
  OR2_X1 U15756 ( .A1(n15706), .A2(n13147), .ZN(n13140) );
  OR2_X1 U15757 ( .A1(n12554), .A2(n11988), .ZN(n13142) );
  NAND2_X1 U15758 ( .A1(n13140), .A2(n13142), .ZN(n13496) );
  OR2_X1 U15759 ( .A1(n12533), .A2(n13496), .ZN(n15813) );
  AND2_X1 U15760 ( .A1(n15798), .A2(n12534), .ZN(n12535) );
  NOR2_X1 U15761 ( .A1(n15813), .A2(n12535), .ZN(n15787) );
  INV_X1 U15762 ( .A(n12536), .ZN(n12537) );
  NAND2_X1 U15763 ( .A1(n15798), .A2(n12537), .ZN(n12538) );
  NAND2_X1 U15764 ( .A1(n15787), .A2(n12538), .ZN(n15734) );
  OR2_X1 U15765 ( .A1(n15734), .A2(n15798), .ZN(n12547) );
  OR2_X1 U15766 ( .A1(n15734), .A2(n12539), .ZN(n12540) );
  NAND2_X1 U15767 ( .A1(n12547), .A2(n12540), .ZN(n15691) );
  INV_X1 U15768 ( .A(n12541), .ZN(n12542) );
  AOI21_X1 U15769 ( .B1(n15798), .B2(n12542), .A(n15473), .ZN(n12543) );
  NAND2_X1 U15770 ( .A1(n15691), .A2(n12543), .ZN(n15654) );
  NAND2_X1 U15771 ( .A1(n15654), .A2(n12547), .ZN(n15642) );
  NAND3_X1 U15772 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12544) );
  NAND2_X1 U15773 ( .A1(n12547), .A2(n12544), .ZN(n12545) );
  NAND2_X1 U15774 ( .A1(n15642), .A2(n12545), .ZN(n15615) );
  INV_X1 U15775 ( .A(n12546), .ZN(n15594) );
  AND2_X1 U15776 ( .A1(n12547), .A2(n15594), .ZN(n12548) );
  INV_X1 U15777 ( .A(n15583), .ZN(n12549) );
  AND2_X1 U15778 ( .A1(n15584), .A2(n12549), .ZN(n15563) );
  OAI21_X1 U15779 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n15570), .A(
        n15563), .ZN(n12558) );
  NAND2_X1 U15780 ( .A1(n12550), .A2(n12551), .ZN(n12552) );
  NAND2_X1 U15781 ( .A1(n12554), .A2(n12553), .ZN(n15811) );
  OR4_X1 U15782 ( .A1(n15564), .A2(n12555), .A3(n15570), .A4(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12556) );
  NAND2_X1 U15783 ( .A1(n15544), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15388) );
  OAI211_X1 U15784 ( .C1(n16199), .C2(n15811), .A(n12556), .B(n15388), .ZN(
        n12557) );
  OAI21_X1 U15785 ( .B1(n16203), .B2(n15816), .A(n12559), .ZN(n12560) );
  AOI21_X1 U15786 ( .B1(n15393), .B2(n16328), .A(n12560), .ZN(n12561) );
  OAI21_X1 U15787 ( .B1(n15395), .B2(n16320), .A(n12561), .ZN(P2_U3017) );
  INV_X1 U15788 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17113) );
  INV_X2 U15789 ( .A(n12562), .ZN(n17020) );
  AOI22_X1 U15790 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12573) );
  INV_X1 U15791 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12565) );
  AOI22_X1 U15792 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17225), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U15793 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12563) );
  OAI211_X1 U15794 ( .C1(n17167), .C2(n12565), .A(n12564), .B(n12563), .ZN(
        n12571) );
  AOI22_X1 U15795 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12569) );
  AOI22_X1 U15796 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12568) );
  AOI22_X1 U15797 ( .A1(n17204), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12567) );
  NAND2_X1 U15798 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12566) );
  NAND4_X1 U15799 ( .A1(n12569), .A2(n12568), .A3(n12567), .A4(n12566), .ZN(
        n12570) );
  INV_X1 U15800 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17025) );
  AOI22_X1 U15801 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15863), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12574) );
  OAI21_X1 U15802 ( .B1(n12562), .B2(n17025), .A(n12574), .ZN(n12583) );
  AOI22_X1 U15803 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12581) );
  INV_X1 U15804 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17029) );
  INV_X1 U15805 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18529) );
  OAI22_X1 U15806 ( .A1(n12608), .A2(n17029), .B1(n17167), .B2(n18529), .ZN(
        n12579) );
  AOI22_X1 U15807 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17231), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12577) );
  AOI22_X1 U15808 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12576) );
  AOI22_X1 U15809 ( .A1(n12616), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17209), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12575) );
  NAND3_X1 U15810 ( .A1(n12577), .A2(n12576), .A3(n12575), .ZN(n12578) );
  AOI211_X1 U15811 ( .C1(n17204), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n12579), .B(n12578), .ZN(n12580) );
  OAI211_X1 U15812 ( .C1(n17241), .C2(n15873), .A(n12581), .B(n12580), .ZN(
        n12582) );
  INV_X1 U15813 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17171) );
  INV_X1 U15814 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18522) );
  OAI22_X1 U15815 ( .A1(n17227), .A2(n17171), .B1(n17167), .B2(n18522), .ZN(
        n12588) );
  AOI22_X1 U15816 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12586) );
  AOI22_X1 U15817 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U15818 ( .A1(n12616), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17209), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12584) );
  NAND3_X1 U15819 ( .A1(n12586), .A2(n12585), .A3(n12584), .ZN(n12587) );
  AOI211_X1 U15820 ( .C1(n17225), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n12588), .B(n12587), .ZN(n12595) );
  INV_X1 U15821 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17269) );
  AOI22_X1 U15822 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12589) );
  OAI21_X1 U15823 ( .B1(n17208), .B2(n17269), .A(n12589), .ZN(n12593) );
  AOI22_X1 U15824 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15863), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12591) );
  NAND2_X1 U15825 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12590) );
  NAND3_X1 U15826 ( .A1(n12591), .A2(n10166), .A3(n12590), .ZN(n12592) );
  INV_X1 U15827 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17197) );
  AOI22_X1 U15828 ( .A1(n12596), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12599) );
  AOI22_X1 U15829 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12597), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12598) );
  OAI211_X1 U15830 ( .C1(n17235), .C2(n17197), .A(n12599), .B(n12598), .ZN(
        n12600) );
  INV_X1 U15831 ( .A(n12600), .ZN(n12606) );
  AOI22_X1 U15832 ( .A1(n17204), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12605) );
  INV_X2 U15833 ( .A(n9699), .ZN(n17181) );
  AOI22_X1 U15834 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12601), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12604) );
  AOI22_X1 U15835 ( .A1(n12643), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12603) );
  NAND2_X1 U15836 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12602) );
  AOI22_X1 U15837 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12607) );
  INV_X1 U15838 ( .A(n17434), .ZN(n12621) );
  AOI22_X1 U15839 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12612) );
  AOI22_X1 U15840 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12611) );
  AOI22_X1 U15841 ( .A1(n9631), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17229), .ZN(n12610) );
  NAND2_X1 U15842 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17209), .ZN(
        n12609) );
  AOI22_X1 U15843 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17020), .ZN(n12614) );
  AOI22_X1 U15844 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n9652), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n12643), .ZN(n12613) );
  OAI211_X1 U15845 ( .C1(n18516), .C2(n17167), .A(n12614), .B(n12613), .ZN(
        n12615) );
  AOI22_X1 U15846 ( .A1(n12601), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n12597), .ZN(n12619) );
  INV_X1 U15847 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17093) );
  NAND2_X1 U15848 ( .A1(n12621), .A2(n12725), .ZN(n12660) );
  AOI22_X1 U15849 ( .A1(n17202), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U15850 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12630) );
  AOI22_X1 U15851 ( .A1(n12616), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17209), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12629) );
  INV_X1 U15852 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17266) );
  INV_X1 U15853 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18525) );
  OAI22_X1 U15854 ( .A1(n17208), .A2(n17266), .B1(n17167), .B2(n18525), .ZN(
        n12627) );
  AOI22_X1 U15855 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12625) );
  AOI22_X1 U15856 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17225), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12624) );
  AOI22_X1 U15857 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12623) );
  NAND2_X1 U15858 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12622) );
  NAND4_X1 U15859 ( .A1(n12625), .A2(n12624), .A3(n12623), .A4(n12622), .ZN(
        n12626) );
  AOI211_X1 U15860 ( .C1(n9631), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n12627), .B(n12626), .ZN(n12628) );
  NAND4_X1 U15861 ( .A1(n12631), .A2(n12630), .A3(n12629), .A4(n12628), .ZN(
        n12663) );
  NAND2_X1 U15862 ( .A1(n12664), .A2(n12663), .ZN(n12667) );
  INV_X1 U15863 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U15864 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17204), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12641) );
  INV_X1 U15865 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18532) );
  AOI22_X1 U15866 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12633) );
  AOI22_X1 U15867 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9633), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12632) );
  OAI211_X1 U15868 ( .C1(n17167), .C2(n18532), .A(n12633), .B(n12632), .ZN(
        n12639) );
  AOI22_X1 U15869 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12637) );
  AOI22_X1 U15870 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12636) );
  AOI22_X1 U15871 ( .A1(n17202), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12635) );
  NAND2_X1 U15872 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12634) );
  NAND4_X1 U15873 ( .A1(n12637), .A2(n12636), .A3(n12635), .A4(n12634), .ZN(
        n12638) );
  AOI211_X1 U15874 ( .C1(n12616), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n12639), .B(n12638), .ZN(n12640) );
  OAI211_X1 U15875 ( .C1(n17217), .C2(n17131), .A(n12641), .B(n12640), .ZN(
        n12671) );
  XNOR2_X1 U15876 ( .A(n12658), .B(n12642), .ZN(n17892) );
  INV_X1 U15877 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18890) );
  XNOR2_X1 U15878 ( .A(n18890), .B(n12725), .ZN(n17904) );
  AOI22_X1 U15879 ( .A1(n12643), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12648) );
  AOI22_X1 U15880 ( .A1(n12601), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15863), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12647) );
  AOI22_X1 U15881 ( .A1(n17204), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12646) );
  NAND2_X1 U15882 ( .A1(n12616), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12645) );
  AOI22_X1 U15883 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12655) );
  INV_X1 U15884 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17226) );
  AOI22_X1 U15885 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12650) );
  AOI22_X1 U15886 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12649) );
  OAI211_X1 U15887 ( .C1(n17235), .C2(n17226), .A(n12650), .B(n12649), .ZN(
        n12651) );
  INV_X1 U15888 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18597) );
  NAND2_X1 U15889 ( .A1(n17911), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17910) );
  NOR2_X1 U15890 ( .A1(n17904), .A2(n17910), .ZN(n17903) );
  NOR2_X1 U15891 ( .A1(n12725), .A2(n18890), .ZN(n12657) );
  NOR2_X1 U15892 ( .A1(n17903), .A2(n12657), .ZN(n17893) );
  NOR2_X1 U15893 ( .A1(n17892), .A2(n17893), .ZN(n17891) );
  NOR2_X1 U15894 ( .A1(n12642), .A2(n12658), .ZN(n12659) );
  XNOR2_X1 U15895 ( .A(n17429), .B(n12660), .ZN(n12661) );
  INV_X1 U15896 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18216) );
  XNOR2_X1 U15897 ( .A(n12662), .B(n12661), .ZN(n17885) );
  INV_X1 U15898 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18207) );
  XNOR2_X1 U15899 ( .A(n17426), .B(n12664), .ZN(n12665) );
  XNOR2_X1 U15900 ( .A(n17422), .B(n12667), .ZN(n12668) );
  XNOR2_X1 U15901 ( .A(n12669), .B(n12668), .ZN(n17861) );
  INV_X1 U15902 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18189) );
  NOR2_X2 U15903 ( .A1(n17861), .A2(n18189), .ZN(n17860) );
  NOR2_X1 U15904 ( .A1(n12669), .A2(n12668), .ZN(n12670) );
  INV_X1 U15905 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17851) );
  INV_X1 U15906 ( .A(n12671), .ZN(n17419) );
  XNOR2_X1 U15907 ( .A(n17419), .B(n12672), .ZN(n12673) );
  XOR2_X1 U15908 ( .A(n17851), .B(n12673), .Z(n17846) );
  OAI21_X1 U15909 ( .B1(n12674), .B2(n16437), .A(n17815), .ZN(n12675) );
  INV_X1 U15910 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18175) );
  OR2_X2 U15911 ( .A1(n17842), .A2(n18175), .ZN(n17840) );
  NOR2_X1 U15912 ( .A1(n17815), .A2(n17827), .ZN(n17814) );
  NOR2_X1 U15913 ( .A1(n17814), .A2(n12678), .ZN(n17728) );
  INV_X1 U15914 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18146) );
  NOR2_X1 U15915 ( .A1(n18146), .A2(n18134), .ZN(n18126) );
  INV_X1 U15916 ( .A(n18126), .ZN(n18095) );
  INV_X1 U15917 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18093) );
  NOR2_X1 U15918 ( .A1(n18095), .A2(n18093), .ZN(n18114) );
  NAND2_X1 U15919 ( .A1(n18114), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18108) );
  NAND2_X1 U15920 ( .A1(n18075), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18060) );
  INV_X1 U15921 ( .A(n18060), .ZN(n18078) );
  NAND2_X1 U15922 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18078), .ZN(
        n18049) );
  INV_X1 U15923 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18074) );
  NOR2_X1 U15924 ( .A1(n18049), .A2(n18074), .ZN(n16442) );
  NOR2_X1 U15925 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17798) );
  INV_X1 U15926 ( .A(n17798), .ZN(n17799) );
  NOR2_X1 U15927 ( .A1(n17799), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12677) );
  INV_X1 U15928 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18083) );
  INV_X1 U15929 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18092) );
  INV_X1 U15930 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18076) );
  NAND4_X1 U15931 ( .A1(n18083), .A2(n18092), .A3(n18076), .A4(n18074), .ZN(
        n12679) );
  INV_X1 U15932 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18053) );
  INV_X1 U15933 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18029) );
  NAND2_X1 U15934 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17693) );
  INV_X1 U15935 ( .A(n17693), .ZN(n18028) );
  NAND2_X1 U15936 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17999) );
  INV_X1 U15937 ( .A(n17999), .ZN(n17980) );
  NAND3_X1 U15938 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n17980), .ZN(n17645) );
  INV_X1 U15939 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17992) );
  NOR2_X1 U15940 ( .A1(n17645), .A2(n17992), .ZN(n12689) );
  NAND2_X1 U15941 ( .A1(n18028), .A2(n12689), .ZN(n17968) );
  INV_X1 U15942 ( .A(n17968), .ZN(n15920) );
  NAND2_X1 U15943 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n15920), .ZN(
        n17618) );
  INV_X1 U15944 ( .A(n17618), .ZN(n12685) );
  INV_X1 U15945 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18021) );
  NAND2_X1 U15946 ( .A1(n17690), .A2(n18021), .ZN(n12686) );
  INV_X1 U15947 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18000) );
  NAND2_X1 U15948 ( .A1(n18028), .A2(n17709), .ZN(n17655) );
  INV_X1 U15949 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17631) );
  INV_X1 U15950 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17939) );
  NAND2_X1 U15951 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17924) );
  AND2_X1 U15952 ( .A1(n10022), .A2(n17924), .ZN(n12691) );
  NOR2_X2 U15953 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n12692), .ZN(
        n17572) );
  INV_X1 U15954 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17555) );
  NAND2_X1 U15955 ( .A1(n17572), .A2(n17555), .ZN(n12694) );
  NOR2_X2 U15956 ( .A1(n17574), .A2(n17815), .ZN(n16433) );
  INV_X1 U15957 ( .A(n16433), .ZN(n12693) );
  NAND2_X1 U15958 ( .A1(n12694), .A2(n12693), .ZN(n12695) );
  NOR2_X1 U15959 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17815), .ZN(
        n16447) );
  AOI21_X1 U15960 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17815), .A(
        n16447), .ZN(n17558) );
  INV_X1 U15961 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17918) );
  NOR2_X1 U15962 ( .A1(n17918), .A2(n17555), .ZN(n15924) );
  AND2_X1 U15963 ( .A1(n15924), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16404) );
  NAND2_X1 U15964 ( .A1(n16404), .A2(n16433), .ZN(n12699) );
  INV_X1 U15965 ( .A(n12699), .ZN(n12696) );
  INV_X1 U15966 ( .A(n15973), .ZN(n12705) );
  INV_X1 U15967 ( .A(n12701), .ZN(n12698) );
  INV_X1 U15968 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18891) );
  AOI22_X1 U15969 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n10022), .B1(
        n17815), .B2(n18891), .ZN(n12702) );
  NAND2_X1 U15970 ( .A1(n12698), .A2(n12702), .ZN(n12704) );
  INV_X1 U15971 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16422) );
  OAI21_X1 U15972 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16422), .A(
        n12699), .ZN(n12700) );
  OAI22_X1 U15973 ( .A1(n12701), .A2(n12700), .B1(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18891), .ZN(n12703) );
  OAI22_X1 U15974 ( .A1(n12705), .A2(n12704), .B1(n12703), .B2(n12702), .ZN(
        n16432) );
  INV_X1 U15975 ( .A(n18781), .ZN(n18927) );
  OAI211_X1 U15976 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18539), .A(
        n12707), .B(n12706), .ZN(n12715) );
  OAI211_X1 U15977 ( .C1(n12710), .C2(n12715), .A(n12709), .B(n12708), .ZN(
        n15914) );
  NAND2_X1 U15978 ( .A1(n9649), .A2(n15905), .ZN(n18715) );
  NOR2_X1 U15979 ( .A1(n12711), .A2(n15888), .ZN(n12713) );
  INV_X1 U15980 ( .A(n12714), .ZN(n12716) );
  INV_X1 U15981 ( .A(n16553), .ZN(n18755) );
  OAI21_X1 U15982 ( .B1(n12716), .B2(n12715), .A(n18755), .ZN(n15916) );
  NAND2_X1 U15983 ( .A1(n18273), .A2(n15987), .ZN(n15909) );
  NOR2_X1 U15984 ( .A1(n9649), .A2(n15909), .ZN(n15917) );
  NAND2_X1 U15985 ( .A1(n12718), .A2(n12717), .ZN(n12719) );
  INV_X1 U15986 ( .A(n16437), .ZN(n17415) );
  NAND2_X1 U15987 ( .A1(n18253), .A2(n18883), .ZN(n16549) );
  NAND2_X1 U15988 ( .A1(n18892), .A2(n16549), .ZN(n15878) );
  INV_X1 U15989 ( .A(n15878), .ZN(n18926) );
  NOR2_X1 U15990 ( .A1(n18905), .A2(n18931), .ZN(n17820) );
  INV_X1 U15991 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18869) );
  NOR2_X1 U15992 ( .A1(n18869), .A2(n18140), .ZN(n16427) );
  NOR2_X1 U15993 ( .A1(n17605), .A2(n17606), .ZN(n17583) );
  NAND2_X1 U15994 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17583), .ZN(
        n17564) );
  INV_X1 U15995 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16607) );
  NOR2_X1 U15996 ( .A1(n17564), .A2(n16607), .ZN(n17566) );
  NAND2_X1 U15997 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17566), .ZN(
        n16413) );
  NOR2_X1 U15998 ( .A1(n16593), .A2(n16413), .ZN(n12721) );
  NAND2_X1 U15999 ( .A1(n18783), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18791) );
  NOR2_X1 U16000 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18883), .ZN(
        n18909) );
  NOR2_X1 U16001 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18935) );
  AOI21_X1 U16002 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n18935), .ZN(n18788) );
  NAND3_X1 U16003 ( .A1(n18253), .A2(n18883), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18508) );
  NAND2_X1 U16004 ( .A1(n12721), .A2(n17748), .ZN(n16401) );
  XNOR2_X1 U16005 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12723) );
  NOR2_X1 U16006 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17665), .ZN(
        n16410) );
  OR2_X1 U16007 ( .A1(n18592), .A2(n12721), .ZN(n16414) );
  OAI211_X1 U16008 ( .C1(n12722), .C2(n18791), .A(n16414), .B(n17912), .ZN(
        n16409) );
  NOR2_X1 U16009 ( .A1(n16410), .A2(n16409), .ZN(n16400) );
  OAI22_X1 U16010 ( .A1(n16401), .A2(n12723), .B1(n16400), .B2(n9894), .ZN(
        n12724) );
  AOI211_X1 U16011 ( .C1(n17770), .C2(n12005), .A(n16427), .B(n12724), .ZN(
        n12760) );
  NAND3_X1 U16012 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n18891), .ZN(n16424) );
  NAND2_X1 U16013 ( .A1(n17911), .A2(n12725), .ZN(n12730) );
  NAND2_X1 U16014 ( .A1(n17434), .A2(n12730), .ZN(n12729) );
  INV_X1 U16015 ( .A(n17429), .ZN(n12728) );
  NAND2_X1 U16016 ( .A1(n12729), .A2(n12728), .ZN(n12739) );
  NOR2_X1 U16017 ( .A1(n17426), .A2(n12739), .ZN(n12727) );
  INV_X1 U16018 ( .A(n17422), .ZN(n12726) );
  NAND2_X1 U16019 ( .A1(n12727), .A2(n12726), .ZN(n12744) );
  NOR2_X1 U16020 ( .A1(n17419), .A2(n12744), .ZN(n12748) );
  NAND2_X1 U16021 ( .A1(n12748), .A2(n16437), .ZN(n12749) );
  XNOR2_X1 U16022 ( .A(n12727), .B(n17422), .ZN(n12742) );
  XNOR2_X1 U16023 ( .A(n12729), .B(n12728), .ZN(n12737) );
  NOR2_X1 U16024 ( .A1(n12737), .A2(n18216), .ZN(n12738) );
  XOR2_X1 U16025 ( .A(n17434), .B(n12730), .Z(n12731) );
  NOR2_X1 U16026 ( .A1(n12731), .A2(n12642), .ZN(n12736) );
  XOR2_X1 U16027 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12731), .Z(
        n17895) );
  INV_X1 U16028 ( .A(n17911), .ZN(n12733) );
  OAI21_X1 U16029 ( .B1(n18890), .B2(n17445), .A(n12733), .ZN(n12734) );
  NAND2_X1 U16030 ( .A1(n18890), .A2(n17445), .ZN(n12732) );
  OAI221_X1 U16031 ( .B1(n12734), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C1(
        n17445), .C2(n12733), .A(n12732), .ZN(n17894) );
  NOR2_X1 U16032 ( .A1(n17895), .A2(n17894), .ZN(n12735) );
  NOR2_X1 U16033 ( .A1(n12736), .A2(n12735), .ZN(n17883) );
  XOR2_X1 U16034 ( .A(n12737), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n17882) );
  NOR2_X1 U16035 ( .A1(n17883), .A2(n17882), .ZN(n17881) );
  NOR2_X1 U16036 ( .A1(n12738), .A2(n17881), .ZN(n12740) );
  NOR2_X1 U16037 ( .A1(n12740), .A2(n18207), .ZN(n12741) );
  XNOR2_X1 U16038 ( .A(n12739), .B(n17426), .ZN(n17872) );
  XOR2_X1 U16039 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n12740), .Z(
        n17871) );
  NOR2_X1 U16040 ( .A1(n17872), .A2(n17871), .ZN(n17870) );
  XOR2_X1 U16041 ( .A(n18189), .B(n12742), .Z(n17858) );
  XNOR2_X1 U16042 ( .A(n12744), .B(n17419), .ZN(n12746) );
  NOR2_X1 U16043 ( .A1(n12745), .A2(n12746), .ZN(n12747) );
  XNOR2_X1 U16044 ( .A(n12746), .B(n12745), .ZN(n17852) );
  XNOR2_X1 U16045 ( .A(n12748), .B(n16437), .ZN(n12751) );
  NAND2_X1 U16046 ( .A1(n12750), .A2(n12751), .ZN(n17837) );
  NAND2_X1 U16047 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17837), .ZN(
        n12753) );
  NOR2_X1 U16048 ( .A1(n12749), .A2(n12753), .ZN(n12755) );
  INV_X1 U16049 ( .A(n12749), .ZN(n12754) );
  OR2_X1 U16050 ( .A1(n12751), .A2(n12750), .ZN(n17838) );
  OAI21_X1 U16051 ( .B1(n12754), .B2(n12753), .A(n17838), .ZN(n12752) );
  AOI21_X1 U16052 ( .B1(n12754), .B2(n12753), .A(n12752), .ZN(n17826) );
  NAND2_X1 U16053 ( .A1(n17955), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17600) );
  NAND2_X1 U16054 ( .A1(n17920), .A2(n15924), .ZN(n16439) );
  NAND2_X1 U16055 ( .A1(n17920), .A2(n16404), .ZN(n16398) );
  OAI21_X1 U16056 ( .B1(n16422), .B2(n16398), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12756) );
  OAI21_X1 U16057 ( .B1(n16424), .B2(n16439), .A(n12756), .ZN(n16429) );
  INV_X1 U16058 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17960) );
  NOR2_X1 U16059 ( .A1(n17631), .A2(n17960), .ZN(n17942) );
  INV_X1 U16060 ( .A(n17942), .ZN(n17923) );
  NOR2_X1 U16061 ( .A1(n17924), .A2(n17923), .ZN(n15927) );
  NAND2_X1 U16062 ( .A1(n15920), .A2(n15927), .ZN(n17917) );
  NAND2_X1 U16063 ( .A1(n15924), .A2(n17919), .ZN(n16438) );
  NAND2_X1 U16064 ( .A1(n16404), .A2(n17919), .ZN(n16397) );
  OAI21_X1 U16065 ( .B1(n16422), .B2(n16397), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12758) );
  OAI21_X1 U16066 ( .B1(n16424), .B2(n16438), .A(n12758), .ZN(n16428) );
  AOI22_X1 U16067 ( .A1(n17902), .A2(n16429), .B1(n17828), .B2(n16428), .ZN(
        n12759) );
  OAI21_X1 U16068 ( .B1(n16432), .B2(n17831), .A(n12761), .ZN(P3_U2799) );
  AOI21_X1 U16069 ( .B1(n15399), .B2(n12764), .A(n12765), .ZN(n15397) );
  NAND2_X1 U16070 ( .A1(n12770), .A2(n12767), .ZN(n12768) );
  NAND2_X1 U16071 ( .A1(n12764), .A2(n12768), .ZN(n15410) );
  INV_X1 U16072 ( .A(n15410), .ZN(n16210) );
  AOI21_X1 U16073 ( .B1(n15422), .B2(n12769), .A(n12766), .ZN(n15425) );
  OAI21_X1 U16074 ( .B1(n12771), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n12772), .ZN(n15456) );
  INV_X1 U16075 ( .A(n15456), .ZN(n12891) );
  AOI21_X1 U16076 ( .B1(n9688), .B2(n11846), .A(n12771), .ZN(n18982) );
  OAI21_X1 U16077 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12773), .A(
        n9688), .ZN(n15487) );
  INV_X1 U16078 ( .A(n15487), .ZN(n18993) );
  AOI21_X1 U16079 ( .B1(n15499), .B2(n9687), .A(n12773), .ZN(n19001) );
  NOR2_X1 U16080 ( .A1(n15521), .A2(n12774), .ZN(n12792) );
  OAI21_X1 U16081 ( .B1(n12792), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n9687), .ZN(n12775) );
  INV_X1 U16082 ( .A(n12775), .ZN(n15512) );
  AOI21_X1 U16083 ( .B1(n12776), .B2(n15545), .A(n12777), .ZN(n15547) );
  AOI21_X1 U16084 ( .B1(n16253), .B2(n12789), .A(n12778), .ZN(n19051) );
  NOR2_X1 U16085 ( .A1(n19074), .A2(n12779), .ZN(n12790) );
  AOI21_X1 U16086 ( .B1(n19074), .B2(n12779), .A(n12790), .ZN(n19084) );
  NAND2_X1 U16087 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n12780), .ZN(
        n12787) );
  AOI21_X1 U16088 ( .B1(n15557), .B2(n12787), .A(n12788), .ZN(n19088) );
  INV_X1 U16089 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13947) );
  NAND2_X1 U16090 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n12781), .ZN(
        n12786) );
  AOI21_X1 U16091 ( .B1(n13947), .B2(n12786), .A(n12780), .ZN(n13950) );
  AOI21_X1 U16092 ( .B1(n16309), .B2(n12782), .A(n12781), .ZN(n19120) );
  AOI21_X1 U16093 ( .B1(n12785), .B2(n12783), .A(n12784), .ZN(n13538) );
  OAI22_X1 U16094 ( .A1(n19987), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19146) );
  INV_X1 U16095 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13808) );
  OAI22_X1 U16096 ( .A1(n19987), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13808), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13768) );
  AND2_X1 U16097 ( .A1(n19146), .A2(n13768), .ZN(n13671) );
  OAI21_X1 U16098 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12783), .ZN(n14461) );
  NAND2_X1 U16099 ( .A1(n13671), .A2(n14461), .ZN(n13536) );
  NOR2_X1 U16100 ( .A1(n13538), .A2(n13536), .ZN(n13557) );
  OAI21_X1 U16101 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12784), .A(
        n12782), .ZN(n19239) );
  NAND2_X1 U16102 ( .A1(n13557), .A2(n19239), .ZN(n19118) );
  NOR2_X1 U16103 ( .A1(n19120), .A2(n19118), .ZN(n19104) );
  OAI21_X1 U16104 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12781), .A(
        n12786), .ZN(n19106) );
  NAND2_X1 U16105 ( .A1(n19104), .A2(n19106), .ZN(n13608) );
  NOR2_X1 U16106 ( .A1(n13950), .A2(n13608), .ZN(n13586) );
  OAI21_X1 U16107 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12780), .A(
        n12787), .ZN(n16293) );
  NAND2_X1 U16108 ( .A1(n13586), .A2(n16293), .ZN(n19087) );
  NOR2_X1 U16109 ( .A1(n19088), .A2(n19087), .ZN(n13574) );
  OAI21_X1 U16110 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12788), .A(
        n12779), .ZN(n16277) );
  NAND2_X1 U16111 ( .A1(n13574), .A2(n16277), .ZN(n19072) );
  NOR2_X1 U16112 ( .A1(n19084), .A2(n19072), .ZN(n19071) );
  OAI21_X1 U16113 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12790), .A(
        n12789), .ZN(n19061) );
  NAND2_X1 U16114 ( .A1(n19071), .A2(n19061), .ZN(n19050) );
  NOR2_X1 U16115 ( .A1(n19051), .A2(n19050), .ZN(n19037) );
  OAI21_X1 U16116 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n12778), .A(
        n12776), .ZN(n19038) );
  NAND2_X1 U16117 ( .A1(n19037), .A2(n19038), .ZN(n12854) );
  NOR2_X1 U16118 ( .A1(n15547), .A2(n12854), .ZN(n19027) );
  OAI21_X1 U16119 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12777), .A(
        n12774), .ZN(n19029) );
  AOI21_X1 U16120 ( .B1(n12774), .B2(n15521), .A(n12792), .ZN(n19017) );
  NOR2_X1 U16121 ( .A1(n19105), .A2(n15228), .ZN(n18999) );
  NOR2_X1 U16122 ( .A1(n19001), .A2(n18999), .ZN(n19000) );
  NOR2_X1 U16123 ( .A1(n19105), .A2(n19000), .ZN(n18991) );
  NOR2_X1 U16124 ( .A1(n18993), .A2(n18991), .ZN(n18992) );
  NOR2_X1 U16125 ( .A1(n19105), .A2(n12890), .ZN(n12866) );
  AOI21_X1 U16126 ( .B1(n15441), .B2(n12772), .A(n12793), .ZN(n15444) );
  OR2_X1 U16127 ( .A1(n12866), .A2(n15444), .ZN(n12867) );
  INV_X1 U16128 ( .A(n19105), .ZN(n12794) );
  NAND2_X1 U16129 ( .A1(n12867), .A2(n12794), .ZN(n16221) );
  OR2_X1 U16130 ( .A1(n12793), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12795) );
  AND2_X1 U16131 ( .A1(n12769), .A2(n12795), .ZN(n16223) );
  INV_X1 U16132 ( .A(n16223), .ZN(n12796) );
  NOR2_X1 U16133 ( .A1(n19105), .A2(n16209), .ZN(n12878) );
  NOR2_X1 U16134 ( .A1(n15397), .A2(n12878), .ZN(n12879) );
  NOR2_X1 U16135 ( .A1(n19105), .A2(n12879), .ZN(n15192) );
  INV_X1 U16136 ( .A(n12765), .ZN(n12798) );
  AOI21_X1 U16137 ( .B1(n14202), .B2(n12798), .A(n12797), .ZN(n15195) );
  NOR2_X1 U16138 ( .A1(n12797), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12800) );
  XNOR2_X1 U16139 ( .A(n12799), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16187) );
  XNOR2_X1 U16140 ( .A(n12801), .B(n16187), .ZN(n12832) );
  NAND4_X1 U16141 ( .A1(n19769), .A2(n19987), .A3(n19643), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19851) );
  INV_X1 U16142 ( .A(n12805), .ZN(n12803) );
  AOI222_X1 U16143 ( .A1(n12314), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n12503), 
        .B2(P2_EAX_REG_30__SCAN_IN), .C1(n14168), .C2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12804) );
  INV_X1 U16144 ( .A(n12804), .ZN(n12802) );
  NOR2_X1 U16145 ( .A1(n16357), .A2(n12509), .ZN(n13259) );
  AND3_X1 U16146 ( .A1(n19970), .A2(n19643), .A3(n12914), .ZN(n16385) );
  NAND2_X1 U16147 ( .A1(n12808), .A2(n12807), .ZN(n12810) );
  NOR2_X1 U16148 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19867), .ZN(n12814) );
  INV_X1 U16149 ( .A(n12814), .ZN(n12825) );
  NOR2_X1 U16150 ( .A1(n12811), .A2(n12825), .ZN(n12812) );
  INV_X1 U16151 ( .A(n12813), .ZN(n12822) );
  INV_X1 U16152 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n15234) );
  NOR2_X1 U16153 ( .A1(n12814), .A2(n15234), .ZN(n12815) );
  AND2_X1 U16154 ( .A1(n19971), .A2(n12815), .ZN(n12816) );
  NAND2_X1 U16155 ( .A1(n19980), .A2(n12816), .ZN(n19101) );
  NOR3_X1 U16156 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n12817), .A3(n19645), 
        .ZN(n16380) );
  INV_X1 U16157 ( .A(n16380), .ZN(n12818) );
  NAND2_X1 U16158 ( .A1(n19851), .A2(n12818), .ZN(n12819) );
  OR2_X1 U16159 ( .A1(n15544), .A2(n12819), .ZN(n12820) );
  NAND2_X1 U16160 ( .A1(n19133), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19073) );
  INV_X2 U16161 ( .A(n19073), .ZN(n19142) );
  AOI22_X1 U16162 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(n19076), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n19142), .ZN(n12821) );
  OAI21_X1 U16163 ( .B1(n12822), .B2(n19101), .A(n12821), .ZN(n12828) );
  AND2_X1 U16164 ( .A1(n16386), .A2(n13262), .ZN(n12919) );
  NAND2_X1 U16165 ( .A1(n12919), .A2(n11388), .ZN(n12823) );
  NAND2_X1 U16166 ( .A1(n12914), .A2(n19643), .ZN(n12824) );
  AND2_X1 U16167 ( .A1(n12963), .A2(n12824), .ZN(n16185) );
  AND3_X1 U16168 ( .A1(n12905), .A2(n15234), .A3(n12825), .ZN(n12826) );
  OR2_X2 U16169 ( .A1(n16185), .A2(n12826), .ZN(n19135) );
  AND2_X1 U16170 ( .A1(n19135), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12827) );
  OAI21_X1 U16171 ( .B1(n12832), .B2(n19851), .A(n12831), .ZN(P2_U2825) );
  AOI21_X1 U16172 ( .B1(n12834), .B2(n12833), .A(n14153), .ZN(n14872) );
  INV_X1 U16173 ( .A(n14872), .ZN(n14789) );
  NOR2_X1 U16174 ( .A1(n14549), .A2(n12835), .ZN(n12836) );
  NOR2_X1 U16175 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12840) );
  NOR4_X1 U16176 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12839) );
  NAND4_X1 U16177 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12840), .A4(n12839), .ZN(n12852) );
  NOR2_X1 U16178 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12852), .ZN(n16529)
         );
  INV_X1 U16179 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21028) );
  INV_X1 U16180 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n20979) );
  NOR4_X1 U16181 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), .A3(
        n21028), .A4(n20979), .ZN(n12842) );
  NOR4_X1 U16182 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n12841)
         );
  NAND3_X1 U16183 ( .A1(n20238), .A2(n12842), .A3(n12841), .ZN(U214) );
  NOR4_X1 U16184 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12846) );
  NOR4_X1 U16185 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12845) );
  NOR4_X1 U16186 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12844) );
  NOR4_X1 U16187 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12843) );
  NAND4_X1 U16188 ( .A1(n12846), .A2(n12845), .A3(n12844), .A4(n12843), .ZN(
        n12851) );
  NOR4_X1 U16189 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12849) );
  NOR4_X1 U16190 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12848) );
  NOR4_X1 U16191 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12847) );
  INV_X1 U16192 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19875) );
  NAND4_X1 U16193 ( .A1(n12849), .A2(n12848), .A3(n12847), .A4(n19875), .ZN(
        n12850) );
  NOR2_X1 U16194 ( .A1(n13854), .A2(n12852), .ZN(n16453) );
  NAND2_X1 U16195 ( .A1(n16453), .A2(U214), .ZN(U212) );
  INV_X1 U16196 ( .A(n19851), .ZN(n19123) );
  NAND2_X1 U16197 ( .A1(n19123), .A2(n12794), .ZN(n19145) );
  AOI211_X1 U16198 ( .C1(n15547), .C2(n12854), .A(n19027), .B(n19145), .ZN(
        n12865) );
  INV_X1 U16199 ( .A(n19135), .ZN(n19100) );
  INV_X1 U16200 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n13824) );
  OAI22_X1 U16201 ( .A1(n19100), .A2(n13824), .B1(n15545), .B2(n19073), .ZN(
        n12864) );
  NOR2_X1 U16202 ( .A1(n19851), .A2(n12794), .ZN(n19141) );
  AOI22_X1 U16203 ( .A1(n12855), .A2(n19131), .B1(n19141), .B2(n15547), .ZN(
        n12856) );
  OAI211_X1 U16204 ( .C1(n19888), .C2(n19133), .A(n12856), .B(n19113), .ZN(
        n12863) );
  OAI21_X1 U16205 ( .B1(n12857), .B2(n12859), .A(n12858), .ZN(n15736) );
  NAND2_X1 U16206 ( .A1(n13714), .A2(n12860), .ZN(n12861) );
  NAND2_X1 U16207 ( .A1(n13849), .A2(n12861), .ZN(n15730) );
  OAI22_X1 U16208 ( .A1(n15736), .A2(n19127), .B1(n19137), .B2(n15730), .ZN(
        n12862) );
  OR4_X1 U16209 ( .A1(n12865), .A2(n12864), .A3(n12863), .A4(n12862), .ZN(
        P2_U2840) );
  INV_X1 U16210 ( .A(n12867), .ZN(n12868) );
  AOI211_X1 U16211 ( .C1(n15444), .C2(n12866), .A(n12868), .B(n19851), .ZN(
        n12877) );
  OAI22_X1 U16212 ( .A1(n12869), .A2(n19101), .B1(n19902), .B2(n19133), .ZN(
        n12876) );
  INV_X1 U16213 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n15279) );
  OAI22_X1 U16214 ( .A1(n19100), .A2(n15279), .B1(n15441), .B2(n19073), .ZN(
        n12875) );
  OR2_X1 U16215 ( .A1(n12895), .A2(n12870), .ZN(n12871) );
  AND2_X1 U16216 ( .A1(n12871), .A2(n15354), .ZN(n15635) );
  INV_X1 U16217 ( .A(n15635), .ZN(n15368) );
  AND2_X1 U16218 ( .A1(n9695), .A2(n12872), .ZN(n12873) );
  OR2_X1 U16219 ( .A1(n12873), .A2(n15267), .ZN(n15629) );
  OAI22_X1 U16220 ( .A1(n15368), .A2(n19127), .B1(n19137), .B2(n15629), .ZN(
        n12874) );
  OR4_X1 U16221 ( .A1(n12877), .A2(n12876), .A3(n12875), .A4(n12874), .ZN(
        P2_U2832) );
  AOI211_X1 U16222 ( .C1(n15397), .C2(n12878), .A(n12879), .B(n19851), .ZN(
        n12889) );
  OAI22_X1 U16223 ( .A1(n12880), .A2(n19101), .B1(n19910), .B2(n19133), .ZN(
        n12888) );
  AOI22_X1 U16224 ( .A1(n19135), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n19142), .ZN(n12881) );
  INV_X1 U16225 ( .A(n12881), .ZN(n12887) );
  OAI21_X1 U16226 ( .B1(n15334), .B2(n12882), .A(n15190), .ZN(n15586) );
  AOI21_X1 U16227 ( .B1(n12885), .B2(n12883), .A(n12884), .ZN(n15404) );
  INV_X1 U16228 ( .A(n15404), .ZN(n15581) );
  OAI22_X1 U16229 ( .A1(n15586), .A2(n19127), .B1(n15581), .B2(n19137), .ZN(
        n12886) );
  OR4_X1 U16230 ( .A1(n12889), .A2(n12888), .A3(n12887), .A4(n12886), .ZN(
        P2_U2828) );
  AOI211_X1 U16231 ( .C1(n12891), .C2(n9746), .A(n12890), .B(n19851), .ZN(
        n12903) );
  INV_X1 U16232 ( .A(n12892), .ZN(n12893) );
  OAI22_X1 U16233 ( .A1(n12893), .A2(n19101), .B1(n19073), .B2(n11928), .ZN(
        n12902) );
  AOI22_X1 U16234 ( .A1(n19135), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19076), .ZN(n12894) );
  INV_X1 U16235 ( .A(n12894), .ZN(n12901) );
  AOI21_X1 U16236 ( .B1(n12897), .B2(n12896), .A(n12895), .ZN(n15640) );
  INV_X1 U16237 ( .A(n15640), .ZN(n15373) );
  NAND2_X1 U16238 ( .A1(n9736), .A2(n12898), .ZN(n12899) );
  AND2_X1 U16239 ( .A1(n9695), .A2(n12899), .ZN(n15645) );
  INV_X1 U16240 ( .A(n15645), .ZN(n15283) );
  OAI22_X1 U16241 ( .A1(n15373), .A2(n19127), .B1(n19137), .B2(n15283), .ZN(
        n12900) );
  OR4_X1 U16242 ( .A1(n12903), .A2(n12902), .A3(n12901), .A4(n12900), .ZN(
        P2_U2833) );
  NOR2_X1 U16243 ( .A1(n12265), .A2(n19845), .ZN(n13021) );
  NAND2_X1 U16244 ( .A1(n12904), .A2(n13021), .ZN(n13683) );
  INV_X1 U16245 ( .A(n13683), .ZN(n19140) );
  INV_X1 U16246 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12908) );
  INV_X1 U16247 ( .A(n12905), .ZN(n12907) );
  INV_X1 U16248 ( .A(n19939), .ZN(n19719) );
  NOR2_X1 U16249 ( .A1(n19719), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12909) );
  INV_X1 U16250 ( .A(n12909), .ZN(n12906) );
  OAI211_X1 U16251 ( .C1(n19140), .C2(n12908), .A(n12907), .B(n12906), .ZN(
        P2_U2814) );
  INV_X1 U16252 ( .A(n12913), .ZN(n12912) );
  INV_X1 U16253 ( .A(n19980), .ZN(n12911) );
  OAI21_X1 U16254 ( .B1(n12909), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n12911), 
        .ZN(n12910) );
  OAI21_X1 U16255 ( .B1(n12912), .B2(n12911), .A(n12910), .ZN(P2_U3612) );
  AND2_X1 U16256 ( .A1(n12913), .A2(n19985), .ZN(n13258) );
  NOR2_X1 U16257 ( .A1(n13258), .A2(n12914), .ZN(n12915) );
  NAND2_X1 U16258 ( .A1(n13259), .A2(n12915), .ZN(n16371) );
  AND2_X1 U16259 ( .A1(n16371), .A2(n13262), .ZN(n19978) );
  INV_X1 U16260 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n15985) );
  OAI21_X1 U16261 ( .B1(n19978), .B2(n15985), .A(n12916), .ZN(P2_U2819) );
  AND2_X1 U16262 ( .A1(n11388), .A2(n12917), .ZN(n12918) );
  NAND2_X1 U16263 ( .A1(n12919), .A2(n12918), .ZN(n12920) );
  INV_X1 U16264 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n12922) );
  NOR2_X1 U16265 ( .A1(n12920), .A2(n11551), .ZN(n13006) );
  INV_X1 U16266 ( .A(n13006), .ZN(n12967) );
  AOI22_X1 U16267 ( .A1(n13853), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13854), .ZN(n19290) );
  NOR2_X1 U16268 ( .A1(n12967), .A2(n19290), .ZN(n12940) );
  AOI21_X1 U16269 ( .B1(n12963), .B2(P2_EAX_REG_23__SCAN_IN), .A(n12940), .ZN(
        n12921) );
  OAI21_X1 U16270 ( .B1(n12982), .B2(n12922), .A(n12921), .ZN(P2_U2959) );
  INV_X1 U16271 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n12924) );
  AOI22_X1 U16272 ( .A1(n13853), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13854), .ZN(n19266) );
  NOR2_X1 U16273 ( .A1(n12967), .A2(n19266), .ZN(n12931) );
  AOI21_X1 U16274 ( .B1(P2_EAX_REG_3__SCAN_IN), .B2(n12963), .A(n12931), .ZN(
        n12923) );
  OAI21_X1 U16275 ( .B1(n12982), .B2(n12924), .A(n12923), .ZN(P2_U2970) );
  INV_X1 U16276 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n12926) );
  OAI22_X1 U16277 ( .A1(n13854), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13853), .ZN(n19270) );
  NOR2_X1 U16278 ( .A1(n12967), .A2(n19270), .ZN(n12937) );
  AOI21_X1 U16279 ( .B1(P2_EAX_REG_4__SCAN_IN), .B2(n12963), .A(n12937), .ZN(
        n12925) );
  OAI21_X1 U16280 ( .B1(n12982), .B2(n12926), .A(n12925), .ZN(P2_U2971) );
  INV_X1 U16281 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n12928) );
  AOI22_X1 U16282 ( .A1(n13853), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13854), .ZN(n19280) );
  NOR2_X1 U16283 ( .A1(n12967), .A2(n19280), .ZN(n12943) );
  AOI21_X1 U16284 ( .B1(n12963), .B2(P2_EAX_REG_6__SCAN_IN), .A(n12943), .ZN(
        n12927) );
  OAI21_X1 U16285 ( .B1(n12982), .B2(n12928), .A(n12927), .ZN(P2_U2973) );
  INV_X1 U16286 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n12930) );
  AOI22_X1 U16287 ( .A1(n13853), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13854), .ZN(n19276) );
  NOR2_X1 U16288 ( .A1(n12967), .A2(n19276), .ZN(n12934) );
  AOI21_X1 U16289 ( .B1(P2_EAX_REG_5__SCAN_IN), .B2(n12963), .A(n12934), .ZN(
        n12929) );
  OAI21_X1 U16290 ( .B1(n12982), .B2(n12930), .A(n12929), .ZN(P2_U2972) );
  INV_X1 U16291 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n12933) );
  AOI21_X1 U16292 ( .B1(n12963), .B2(P2_EAX_REG_19__SCAN_IN), .A(n12931), .ZN(
        n12932) );
  OAI21_X1 U16293 ( .B1(n12982), .B2(n12933), .A(n12932), .ZN(P2_U2955) );
  INV_X1 U16294 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n12936) );
  AOI21_X1 U16295 ( .B1(n12963), .B2(P2_EAX_REG_21__SCAN_IN), .A(n12934), .ZN(
        n12935) );
  OAI21_X1 U16296 ( .B1(n12982), .B2(n12936), .A(n12935), .ZN(P2_U2957) );
  INV_X1 U16297 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n12939) );
  AOI21_X1 U16298 ( .B1(n12963), .B2(P2_EAX_REG_20__SCAN_IN), .A(n12937), .ZN(
        n12938) );
  OAI21_X1 U16299 ( .B1(n12982), .B2(n12939), .A(n12938), .ZN(P2_U2956) );
  INV_X1 U16300 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n12942) );
  AOI21_X1 U16301 ( .B1(n12963), .B2(P2_EAX_REG_7__SCAN_IN), .A(n12940), .ZN(
        n12941) );
  OAI21_X1 U16302 ( .B1(n12982), .B2(n12942), .A(n12941), .ZN(P2_U2974) );
  INV_X1 U16303 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n12945) );
  AOI21_X1 U16304 ( .B1(n12963), .B2(P2_EAX_REG_22__SCAN_IN), .A(n12943), .ZN(
        n12944) );
  OAI21_X1 U16305 ( .B1(n12982), .B2(n12945), .A(n12944), .ZN(P2_U2958) );
  INV_X1 U16306 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n12949) );
  INV_X1 U16307 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16478) );
  OR2_X1 U16308 ( .A1(n13854), .A2(n16478), .ZN(n12947) );
  NAND2_X1 U16309 ( .A1(n13003), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12946) );
  NAND2_X1 U16310 ( .A1(n12947), .A2(n12946), .ZN(n15315) );
  NAND2_X1 U16311 ( .A1(n13006), .A2(n15315), .ZN(n13008) );
  NAND2_X1 U16312 ( .A1(n12963), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n12948) );
  OAI211_X1 U16313 ( .C1(n12982), .C2(n12949), .A(n13008), .B(n12948), .ZN(
        P2_U2980) );
  INV_X1 U16314 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n12953) );
  INV_X1 U16315 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16486) );
  OR2_X1 U16316 ( .A1(n13854), .A2(n16486), .ZN(n12951) );
  NAND2_X1 U16317 ( .A1(n13854), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12950) );
  NAND2_X1 U16318 ( .A1(n12951), .A2(n12950), .ZN(n15343) );
  NAND2_X1 U16319 ( .A1(n13006), .A2(n15343), .ZN(n13001) );
  NAND2_X1 U16320 ( .A1(n12963), .A2(P2_EAX_REG_9__SCAN_IN), .ZN(n12952) );
  OAI211_X1 U16321 ( .C1(n12982), .C2(n12953), .A(n13001), .B(n12952), .ZN(
        P2_U2976) );
  INV_X1 U16322 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n12956) );
  AOI22_X1 U16323 ( .A1(n13853), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13854), .ZN(n19187) );
  INV_X1 U16324 ( .A(n19187), .ZN(n12954) );
  NAND2_X1 U16325 ( .A1(n13006), .A2(n12954), .ZN(n13015) );
  NAND2_X1 U16326 ( .A1(n12963), .A2(P2_EAX_REG_1__SCAN_IN), .ZN(n12955) );
  OAI211_X1 U16327 ( .C1(n12982), .C2(n12956), .A(n13015), .B(n12955), .ZN(
        P2_U2968) );
  INV_X1 U16328 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n12958) );
  OAI22_X1 U16329 ( .A1(n13854), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13853), .ZN(n19261) );
  INV_X1 U16330 ( .A(n19261), .ZN(n16234) );
  NAND2_X1 U16331 ( .A1(n13006), .A2(n16234), .ZN(n13010) );
  NAND2_X1 U16332 ( .A1(n12963), .A2(P2_EAX_REG_2__SCAN_IN), .ZN(n12957) );
  OAI211_X1 U16333 ( .C1(n12982), .C2(n12958), .A(n13010), .B(n12957), .ZN(
        P2_U2969) );
  INV_X1 U16334 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n12960) );
  AOI22_X1 U16335 ( .A1(n13853), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13854), .ZN(n19248) );
  INV_X1 U16336 ( .A(n19248), .ZN(n13856) );
  NAND2_X1 U16337 ( .A1(n13006), .A2(n13856), .ZN(n13018) );
  NAND2_X1 U16338 ( .A1(n12963), .A2(P2_EAX_REG_16__SCAN_IN), .ZN(n12959) );
  OAI211_X1 U16339 ( .C1(n12982), .C2(n12960), .A(n13018), .B(n12959), .ZN(
        P2_U2952) );
  INV_X1 U16340 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n12965) );
  INV_X1 U16341 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16482) );
  OR2_X1 U16342 ( .A1(n13854), .A2(n16482), .ZN(n12962) );
  NAND2_X1 U16343 ( .A1(n13854), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12961) );
  NAND2_X1 U16344 ( .A1(n12962), .A2(n12961), .ZN(n15327) );
  NAND2_X1 U16345 ( .A1(n13006), .A2(n15327), .ZN(n12997) );
  NAND2_X1 U16346 ( .A1(n12963), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n12964) );
  OAI211_X1 U16347 ( .C1(n12982), .C2(n12965), .A(n12997), .B(n12964), .ZN(
        P2_U2978) );
  INV_X1 U16348 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12968) );
  AOI22_X1 U16349 ( .A1(n13853), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13854), .ZN(n13570) );
  INV_X1 U16350 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12966) );
  OAI222_X1 U16351 ( .A1(n12968), .A2(n12982), .B1(n12967), .B2(n13570), .C1(
        n12966), .C2(n13022), .ZN(P2_U2982) );
  NAND2_X1 U16352 ( .A1(n19279), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12970) );
  AOI22_X1 U16353 ( .A1(n13126), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19939), .B2(n19966), .ZN(n12971) );
  INV_X1 U16354 ( .A(n15826), .ZN(n12976) );
  NOR2_X1 U16355 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12973) );
  NOR2_X1 U16356 ( .A1(n19279), .A2(n19987), .ZN(n13041) );
  OAI21_X1 U16357 ( .B1(n12974), .B2(n12973), .A(n13041), .ZN(n12975) );
  NAND2_X1 U16358 ( .A1(n16363), .A2(n15835), .ZN(n13753) );
  NAND2_X1 U16359 ( .A1(n13753), .A2(n9732), .ZN(n12977) );
  MUX2_X1 U16360 ( .A(n19138), .B(n11651), .S(n15269), .Z(n12979) );
  OAI21_X1 U16361 ( .B1(n19961), .B2(n15312), .A(n12979), .ZN(P2_U2887) );
  NAND2_X1 U16362 ( .A1(n14480), .A2(n20000), .ZN(n13038) );
  AND2_X1 U16363 ( .A1(n20783), .A2(n16181), .ZN(n20003) );
  AOI21_X1 U16364 ( .B1(n13038), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n20003), 
        .ZN(n12981) );
  NAND2_X1 U16365 ( .A1(n13248), .A2(n12981), .ZN(P1_U2801) );
  INV_X1 U16366 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19208) );
  NAND2_X1 U16367 ( .A1(n13017), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12985) );
  INV_X1 U16368 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16484) );
  OR2_X1 U16369 ( .A1(n13854), .A2(n16484), .ZN(n12984) );
  NAND2_X1 U16370 ( .A1(n13003), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12983) );
  NAND2_X1 U16371 ( .A1(n12984), .A2(n12983), .ZN(n19159) );
  NAND2_X1 U16372 ( .A1(n13006), .A2(n19159), .ZN(n12989) );
  OAI211_X1 U16373 ( .C1(n19208), .C2(n13022), .A(n12985), .B(n12989), .ZN(
        P2_U2977) );
  INV_X1 U16374 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19204) );
  NAND2_X1 U16375 ( .A1(n13017), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12988) );
  INV_X1 U16376 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16480) );
  OR2_X1 U16377 ( .A1(n13854), .A2(n16480), .ZN(n12987) );
  NAND2_X1 U16378 ( .A1(n13854), .A2(BUF2_REG_12__SCAN_IN), .ZN(n12986) );
  NAND2_X1 U16379 ( .A1(n12987), .A2(n12986), .ZN(n19155) );
  NAND2_X1 U16380 ( .A1(n13006), .A2(n19155), .ZN(n12999) );
  OAI211_X1 U16381 ( .C1(n19204), .C2(n13022), .A(n12988), .B(n12999), .ZN(
        P2_U2979) );
  INV_X1 U16382 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13091) );
  NAND2_X1 U16383 ( .A1(n13017), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12990) );
  OAI211_X1 U16384 ( .C1(n13091), .C2(n13022), .A(n12990), .B(n12989), .ZN(
        P2_U2962) );
  INV_X1 U16385 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19200) );
  NAND2_X1 U16386 ( .A1(n13017), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n12994) );
  INV_X1 U16387 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n12991) );
  OR2_X1 U16388 ( .A1(n13003), .A2(n12991), .ZN(n12993) );
  NAND2_X1 U16389 ( .A1(n13003), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12992) );
  NAND2_X1 U16390 ( .A1(n12993), .A2(n12992), .ZN(n19152) );
  NAND2_X1 U16391 ( .A1(n13006), .A2(n19152), .ZN(n12995) );
  OAI211_X1 U16392 ( .C1(n19200), .C2(n13022), .A(n12994), .B(n12995), .ZN(
        P2_U2981) );
  INV_X1 U16393 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13028) );
  NAND2_X1 U16394 ( .A1(n13017), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12996) );
  OAI211_X1 U16395 ( .C1(n13028), .C2(n13022), .A(n12996), .B(n12995), .ZN(
        P2_U2966) );
  INV_X1 U16396 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13030) );
  NAND2_X1 U16397 ( .A1(n13017), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n12998) );
  OAI211_X1 U16398 ( .C1(n13022), .C2(n13030), .A(n12998), .B(n12997), .ZN(
        P2_U2963) );
  INV_X1 U16399 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13037) );
  NAND2_X1 U16400 ( .A1(n13017), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13000) );
  OAI211_X1 U16401 ( .C1(n13037), .C2(n13022), .A(n13000), .B(n12999), .ZN(
        P2_U2964) );
  INV_X1 U16402 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13035) );
  NAND2_X1 U16403 ( .A1(n13017), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13002) );
  OAI211_X1 U16404 ( .C1(n13022), .C2(n13035), .A(n13002), .B(n13001), .ZN(
        P2_U2961) );
  INV_X1 U16405 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13033) );
  NAND2_X1 U16406 ( .A1(n13017), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13007) );
  INV_X1 U16407 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16488) );
  OR2_X1 U16408 ( .A1(n13854), .A2(n16488), .ZN(n13005) );
  NAND2_X1 U16409 ( .A1(n13003), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13004) );
  NAND2_X1 U16410 ( .A1(n13005), .A2(n13004), .ZN(n19163) );
  NAND2_X1 U16411 ( .A1(n13006), .A2(n19163), .ZN(n13013) );
  OAI211_X1 U16412 ( .C1(n13033), .C2(n13022), .A(n13007), .B(n13013), .ZN(
        P2_U2960) );
  INV_X1 U16413 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13096) );
  NAND2_X1 U16414 ( .A1(n13017), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13009) );
  OAI211_X1 U16415 ( .C1(n13022), .C2(n13096), .A(n13009), .B(n13008), .ZN(
        P2_U2965) );
  INV_X1 U16416 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13012) );
  NAND2_X1 U16417 ( .A1(n13017), .A2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13011) );
  OAI211_X1 U16418 ( .C1(n13022), .C2(n13012), .A(n13011), .B(n13010), .ZN(
        P2_U2954) );
  INV_X1 U16419 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19213) );
  NAND2_X1 U16420 ( .A1(n13017), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13014) );
  OAI211_X1 U16421 ( .C1(n19213), .C2(n13022), .A(n13014), .B(n13013), .ZN(
        P2_U2975) );
  INV_X1 U16422 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13899) );
  NAND2_X1 U16423 ( .A1(n13017), .A2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13016) );
  OAI211_X1 U16424 ( .C1(n13022), .C2(n13899), .A(n13016), .B(n13015), .ZN(
        P2_U2953) );
  NAND2_X1 U16425 ( .A1(n13017), .A2(P2_LWORD_REG_0__SCAN_IN), .ZN(n13019) );
  OAI211_X1 U16426 ( .C1(n13020), .C2(n13022), .A(n13019), .B(n13018), .ZN(
        P2_U2967) );
  INV_X1 U16427 ( .A(n13021), .ZN(n13023) );
  OAI21_X1 U16428 ( .B1(n13024), .B2(n13023), .A(n13022), .ZN(n13025) );
  NAND2_X1 U16429 ( .A1(n19197), .A2(n13026), .ZN(n13095) );
  NOR2_X1 U16430 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19958), .ZN(n13089) );
  AOI22_X1 U16431 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n19211), .B1(n19982), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13027) );
  OAI21_X1 U16432 ( .B1(n13028), .B2(n13095), .A(n13027), .ZN(P2_U2921) );
  AOI22_X1 U16433 ( .A1(n13089), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13029) );
  OAI21_X1 U16434 ( .B1(n13030), .B2(n13095), .A(n13029), .ZN(P2_U2924) );
  INV_X1 U16435 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15361) );
  AOI22_X1 U16436 ( .A1(n13089), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13031) );
  OAI21_X1 U16437 ( .B1(n15361), .B2(n13095), .A(n13031), .ZN(P2_U2928) );
  AOI22_X1 U16438 ( .A1(n13089), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13032) );
  OAI21_X1 U16439 ( .B1(n13033), .B2(n13095), .A(n13032), .ZN(P2_U2927) );
  AOI22_X1 U16440 ( .A1(n13089), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13034) );
  OAI21_X1 U16441 ( .B1(n13035), .B2(n13095), .A(n13034), .ZN(P2_U2926) );
  AOI22_X1 U16442 ( .A1(n19982), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13036) );
  OAI21_X1 U16443 ( .B1(n13037), .B2(n13095), .A(n13036), .ZN(P2_U2923) );
  NOR2_X1 U16444 ( .A1(n20003), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n13040)
         );
  OAI21_X1 U16445 ( .B1(n14484), .B2(n14490), .A(n20916), .ZN(n13039) );
  OAI21_X1 U16446 ( .B1(n13040), .B2(n20916), .A(n13039), .ZN(P1_U3487) );
  NAND2_X1 U16447 ( .A1(n14393), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13119) );
  NAND2_X1 U16448 ( .A1(n13126), .A2(n15832), .ZN(n13042) );
  XNOR2_X1 U16449 ( .A(n19966), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19404) );
  NAND2_X1 U16450 ( .A1(n19404), .A2(n19939), .ZN(n19580) );
  NAND2_X1 U16451 ( .A1(n13042), .A2(n19580), .ZN(n13043) );
  MUX2_X1 U16452 ( .A(n13044), .B(n11502), .S(n15302), .Z(n13045) );
  OAI21_X1 U16453 ( .B1(n19949), .B2(n15312), .A(n13045), .ZN(P2_U2886) );
  INV_X1 U16454 ( .A(n16320), .ZN(n16332) );
  OAI21_X1 U16455 ( .B1(n13807), .B2(n13070), .A(n13046), .ZN(n13047) );
  INV_X1 U16456 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13769) );
  XOR2_X1 U16457 ( .A(n13047), .B(n13769), .Z(n13101) );
  NAND2_X1 U16458 ( .A1(n15544), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13099) );
  OAI21_X1 U16459 ( .B1(n13142), .B2(n13769), .A(n13099), .ZN(n13055) );
  XOR2_X1 U16460 ( .A(n13048), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n13097) );
  XNOR2_X1 U16461 ( .A(n13050), .B(n13049), .ZN(n19954) );
  AOI22_X1 U16462 ( .A1(n16328), .A2(n13097), .B1(n16324), .B2(n19954), .ZN(
        n13053) );
  OAI211_X1 U16463 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n15798), .B(n13051), .ZN(n13052) );
  NAND2_X1 U16464 ( .A1(n13053), .A2(n13052), .ZN(n13054) );
  AOI211_X1 U16465 ( .C1(n16332), .C2(n13101), .A(n13055), .B(n13054), .ZN(
        n13056) );
  OAI21_X1 U16466 ( .B1(n11502), .B2(n15811), .A(n13056), .ZN(P2_U3045) );
  INV_X1 U16467 ( .A(n13057), .ZN(n13060) );
  OAI21_X1 U16468 ( .B1(n13060), .B2(n13059), .A(n13058), .ZN(n14745) );
  INV_X1 U16469 ( .A(n13061), .ZN(n13063) );
  AOI21_X1 U16470 ( .B1(n13063), .B2(n15169), .A(n13062), .ZN(n13308) );
  INV_X1 U16471 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13064) );
  NOR2_X1 U16472 ( .A1(n20225), .A2(n13064), .ZN(n13343) );
  INV_X1 U16473 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13065) );
  AOI21_X1 U16474 ( .B1(n13067), .B2(n13066), .A(n13065), .ZN(n13068) );
  AOI211_X1 U16475 ( .C1(n13308), .C2(n20174), .A(n13343), .B(n13068), .ZN(
        n13069) );
  OAI21_X1 U16476 ( .B1(n16049), .B2(n14745), .A(n13069), .ZN(P1_U2999) );
  OAI21_X1 U16477 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19130), .A(
        n13070), .ZN(n13106) );
  INV_X1 U16478 ( .A(n13106), .ZN(n13079) );
  NAND2_X1 U16479 ( .A1(n15544), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13105) );
  OAI21_X1 U16480 ( .B1(n15811), .B2(n19138), .A(n13105), .ZN(n13078) );
  OAI21_X1 U16481 ( .B1(n13072), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13071), .ZN(n13104) );
  NOR2_X1 U16482 ( .A1(n13074), .A2(n13073), .ZN(n13075) );
  OR2_X1 U16483 ( .A1(n13076), .A2(n13075), .ZN(n19128) );
  OAI22_X1 U16484 ( .A1(n13104), .A2(n15804), .B1(n15816), .B2(n19128), .ZN(
        n13077) );
  AOI211_X1 U16485 ( .C1(n16332), .C2(n13079), .A(n13078), .B(n13077), .ZN(
        n13081) );
  MUX2_X1 U16486 ( .A(n15710), .B(n13142), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13080) );
  NAND2_X1 U16487 ( .A1(n13081), .A2(n13080), .ZN(P2_U3046) );
  OAI21_X1 U16488 ( .B1(n14491), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13082), .ZN(n14741) );
  OAI222_X1 U16489 ( .A1(n14741), .A2(n14777), .B1(n11100), .B2(n14778), .C1(
        n14745), .C2(n14779), .ZN(P1_U2872) );
  AOI22_X1 U16490 ( .A1(n13089), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13083) );
  OAI21_X1 U16491 ( .B1(n13012), .B2(n13095), .A(n13083), .ZN(P2_U2933) );
  INV_X1 U16492 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13993) );
  AOI22_X1 U16493 ( .A1(n13089), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13084) );
  OAI21_X1 U16494 ( .B1(n13993), .B2(n13095), .A(n13084), .ZN(P2_U2932) );
  INV_X1 U16495 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n15372) );
  AOI22_X1 U16496 ( .A1(n13089), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13085) );
  OAI21_X1 U16497 ( .B1(n15372), .B2(n13095), .A(n13085), .ZN(P2_U2929) );
  INV_X1 U16498 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13087) );
  AOI22_X1 U16499 ( .A1(n13089), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13086) );
  OAI21_X1 U16500 ( .B1(n13087), .B2(n13095), .A(n13086), .ZN(P2_U2931) );
  INV_X1 U16501 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15379) );
  AOI22_X1 U16502 ( .A1(n13089), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13088) );
  OAI21_X1 U16503 ( .B1(n15379), .B2(n13095), .A(n13088), .ZN(P2_U2930) );
  AOI22_X1 U16504 ( .A1(n13089), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13090) );
  OAI21_X1 U16505 ( .B1(n13091), .B2(n13095), .A(n13090), .ZN(P2_U2925) );
  AOI22_X1 U16506 ( .A1(n19982), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13092) );
  OAI21_X1 U16507 ( .B1(n13899), .B2(n13095), .A(n13092), .ZN(P2_U2934) );
  INV_X1 U16508 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13859) );
  AOI22_X1 U16509 ( .A1(n19982), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13093) );
  OAI21_X1 U16510 ( .B1(n13859), .B2(n13095), .A(n13093), .ZN(P2_U2935) );
  AOI22_X1 U16511 ( .A1(n19982), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13094) );
  OAI21_X1 U16512 ( .B1(n13096), .B2(n13095), .A(n13094), .ZN(P2_U2922) );
  NAND2_X1 U16513 ( .A1(n19236), .A2(n13097), .ZN(n13098) );
  OAI211_X1 U16514 ( .C1(n16310), .C2(n13808), .A(n13099), .B(n13098), .ZN(
        n13100) );
  AOI21_X1 U16515 ( .B1(n16301), .B2(n13808), .A(n13100), .ZN(n13103) );
  NAND2_X1 U16516 ( .A1(n13101), .A2(n16297), .ZN(n13102) );
  OAI211_X1 U16517 ( .C1(n11502), .C2(n13736), .A(n13103), .B(n13102), .ZN(
        P2_U3013) );
  INV_X1 U16518 ( .A(n13104), .ZN(n13108) );
  OAI21_X1 U16519 ( .B1(n11993), .B2(n13106), .A(n13105), .ZN(n13107) );
  AOI21_X1 U16520 ( .B1(n19236), .B2(n13108), .A(n13107), .ZN(n13111) );
  OAI21_X1 U16521 ( .B1(n19231), .B2(n13109), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13110) );
  OAI211_X1 U16522 ( .C1(n19138), .C2(n13736), .A(n13111), .B(n13110), .ZN(
        P2_U3014) );
  NAND2_X1 U16523 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19609) );
  NAND2_X1 U16524 ( .A1(n19609), .A2(n19946), .ZN(n13112) );
  NOR2_X1 U16525 ( .A1(n19946), .A2(n19956), .ZN(n19715) );
  NAND2_X1 U16526 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19715), .ZN(
        n19243) );
  AND2_X1 U16527 ( .A1(n13112), .A2(n19243), .ZN(n19403) );
  AOI22_X1 U16528 ( .A1(n13126), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19939), .B2(n19403), .ZN(n13113) );
  AND2_X1 U16529 ( .A1(n14393), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13116) );
  NAND2_X1 U16530 ( .A1(n13117), .A2(n13116), .ZN(n13124) );
  OR2_X1 U16531 ( .A1(n13117), .A2(n13116), .ZN(n13118) );
  INV_X1 U16532 ( .A(n13119), .ZN(n13120) );
  NOR2_X1 U16533 ( .A1(n15826), .A2(n13120), .ZN(n13121) );
  NAND2_X1 U16534 ( .A1(n13520), .A2(n13521), .ZN(n13125) );
  NAND2_X1 U16535 ( .A1(n13125), .A2(n13124), .ZN(n13136) );
  NAND2_X1 U16536 ( .A1(n13126), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13130) );
  NAND2_X1 U16537 ( .A1(n19243), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13128) );
  NAND2_X1 U16538 ( .A1(n19715), .A2(n19938), .ZN(n19493) );
  INV_X1 U16539 ( .A(n19493), .ZN(n13127) );
  NAND2_X1 U16540 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13127), .ZN(
        n19524) );
  NAND2_X1 U16541 ( .A1(n13128), .A2(n19524), .ZN(n13129) );
  NAND2_X1 U16542 ( .A1(n19939), .A2(n13129), .ZN(n19655) );
  NAND2_X1 U16543 ( .A1(n13130), .A2(n19655), .ZN(n13131) );
  NAND2_X1 U16544 ( .A1(n14393), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13133) );
  NAND2_X1 U16545 ( .A1(n13134), .A2(n13133), .ZN(n13135) );
  MUX2_X1 U16546 ( .A(n13138), .B(n11648), .S(n15269), .Z(n13139) );
  OAI21_X1 U16547 ( .B1(n19934), .B2(n15312), .A(n13139), .ZN(P2_U2884) );
  OAI21_X1 U16548 ( .B1(n13142), .B2(n13141), .A(n13140), .ZN(n13160) );
  NAND2_X1 U16549 ( .A1(n13144), .A2(n13143), .ZN(n13146) );
  AND2_X1 U16550 ( .A1(n13146), .A2(n9957), .ZN(n13718) );
  INV_X1 U16551 ( .A(n13718), .ZN(n19944) );
  INV_X1 U16552 ( .A(n13147), .ZN(n13148) );
  NAND2_X1 U16553 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(n15544), .ZN(n14462) );
  OAI221_X1 U16554 ( .B1(n13149), .B2(n13161), .C1(n13149), .C2(n13148), .A(
        n14462), .ZN(n13150) );
  AOI21_X1 U16555 ( .B1(n19944), .B2(n16324), .A(n13150), .ZN(n13158) );
  NAND2_X1 U16556 ( .A1(n13152), .A2(n13151), .ZN(n14465) );
  AND2_X1 U16557 ( .A1(n14466), .A2(n14465), .ZN(n13156) );
  INV_X1 U16558 ( .A(n13153), .ZN(n13154) );
  XNOR2_X1 U16559 ( .A(n13155), .B(n13154), .ZN(n14469) );
  AOI22_X1 U16560 ( .A1(n16332), .A2(n13156), .B1(n16328), .B2(n14469), .ZN(
        n13157) );
  OAI211_X1 U16561 ( .C1(n15841), .C2(n15811), .A(n13158), .B(n13157), .ZN(
        n13159) );
  AOI21_X1 U16562 ( .B1(n13161), .B2(n13160), .A(n13159), .ZN(n13162) );
  INV_X1 U16563 ( .A(n13162), .ZN(P2_U3044) );
  INV_X1 U16564 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20525) );
  NAND2_X1 U16565 ( .A1(n13163), .A2(n20258), .ZN(n13318) );
  AND3_X1 U16566 ( .A1(n13164), .A2(n20244), .A3(n13318), .ZN(n13188) );
  INV_X1 U16567 ( .A(n13165), .ZN(n13417) );
  AOI21_X1 U16568 ( .B1(n10318), .B2(n20263), .A(n14161), .ZN(n13166) );
  AND2_X1 U16569 ( .A1(n13167), .A2(n20258), .ZN(n13168) );
  NOR2_X1 U16570 ( .A1(n13188), .A2(n13168), .ZN(n13175) );
  AOI22_X1 U16571 ( .A1(n14491), .A2(n13169), .B1(n20244), .B2(n20263), .ZN(
        n13170) );
  OAI21_X1 U16572 ( .B1(n13171), .B2(n11155), .A(n13170), .ZN(n13172) );
  INV_X1 U16573 ( .A(n13172), .ZN(n13174) );
  NAND2_X1 U16574 ( .A1(n10307), .A2(n14484), .ZN(n13173) );
  AND3_X1 U16575 ( .A1(n13175), .A2(n13174), .A3(n13173), .ZN(n13335) );
  NAND2_X1 U16576 ( .A1(n13178), .A2(n13336), .ZN(n13179) );
  NOR2_X1 U16577 ( .A1(n13177), .A2(n13179), .ZN(n13180) );
  NAND3_X1 U16578 ( .A1(n13335), .A2(n13176), .A3(n13180), .ZN(n13439) );
  AOI22_X1 U16579 ( .A1(n10445), .A2(n13439), .B1(n15164), .B2(n13182), .ZN(
        n15936) );
  OAI22_X1 U16580 ( .A1(n15936), .A2(n15184), .B1(n16181), .B2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13181) );
  AOI21_X1 U16581 ( .B1(n15968), .B2(n13182), .A(n13181), .ZN(n13199) );
  AND2_X1 U16582 ( .A1(n11062), .A2(n20258), .ZN(n15166) );
  INV_X1 U16583 ( .A(n13183), .ZN(n13184) );
  INV_X1 U16584 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20847) );
  NAND2_X1 U16585 ( .A1(n13184), .A2(n20847), .ZN(n15981) );
  INV_X1 U16586 ( .A(n15981), .ZN(n13185) );
  NAND2_X1 U16587 ( .A1(n15166), .A2(n13185), .ZN(n13226) );
  OR2_X1 U16588 ( .A1(n9636), .A2(n13185), .ZN(n14485) );
  NAND2_X1 U16589 ( .A1(n13177), .A2(n14485), .ZN(n13186) );
  INV_X1 U16590 ( .A(n20918), .ZN(n15980) );
  AOI21_X1 U16591 ( .B1(n13226), .B2(n13186), .A(n15980), .ZN(n13187) );
  MUX2_X1 U16592 ( .A(n13187), .B(n14474), .S(n14483), .Z(n13194) );
  NOR2_X1 U16593 ( .A1(n13189), .A2(n13188), .ZN(n13190) );
  NOR2_X1 U16594 ( .A1(n11062), .A2(n13190), .ZN(n13319) );
  NAND2_X1 U16595 ( .A1(n13632), .A2(n20258), .ZN(n13643) );
  NOR2_X1 U16596 ( .A1(n13643), .A2(n20263), .ZN(n13191) );
  OR2_X1 U16597 ( .A1(n13319), .A2(n13191), .ZN(n13192) );
  NAND2_X1 U16598 ( .A1(n15939), .A2(n20000), .ZN(n13197) );
  NAND2_X1 U16599 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16177) );
  INV_X1 U16600 ( .A(n16177), .ZN(n13447) );
  NAND2_X1 U16601 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13447), .ZN(n16182) );
  INV_X1 U16602 ( .A(n16182), .ZN(n13195) );
  NAND2_X1 U16603 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13195), .ZN(n13196) );
  NAND2_X1 U16604 ( .A1(n13197), .A2(n13196), .ZN(n16171) );
  AOI21_X1 U16605 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20914), .A(n16171), 
        .ZN(n15173) );
  AND2_X1 U16606 ( .A1(n15166), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15937) );
  AOI22_X1 U16607 ( .A1(n15937), .A2(n16172), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15173), .ZN(n13198) );
  OAI21_X1 U16608 ( .B1(n13199), .B2(n15173), .A(n13198), .ZN(P1_U3474) );
  NAND2_X1 U16609 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19279), .ZN(
        n13200) );
  XOR2_X1 U16610 ( .A(n13217), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13208)
         );
  NAND2_X1 U16611 ( .A1(n13203), .A2(n13212), .ZN(n13205) );
  AND2_X1 U16612 ( .A1(n13205), .A2(n10051), .ZN(n19121) );
  INV_X1 U16613 ( .A(n19121), .ZN(n13786) );
  MUX2_X1 U16614 ( .A(n13786), .B(n13206), .S(n15269), .Z(n13207) );
  OAI21_X1 U16615 ( .B1(n13208), .B2(n15312), .A(n13207), .ZN(P2_U2882) );
  OAI21_X1 U16616 ( .B1(n13210), .B2(n13209), .A(n13217), .ZN(n19168) );
  OR2_X1 U16617 ( .A1(n9762), .A2(n13211), .ZN(n13213) );
  AND2_X1 U16618 ( .A1(n13213), .A2(n13212), .ZN(n13602) );
  INV_X1 U16619 ( .A(n13602), .ZN(n19232) );
  NOR2_X1 U16620 ( .A1(n19232), .A2(n15309), .ZN(n13214) );
  AOI21_X1 U16621 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n15309), .A(n13214), .ZN(
        n13215) );
  OAI21_X1 U16622 ( .B1(n19168), .B2(n15312), .A(n13215), .ZN(P2_U2883) );
  INV_X1 U16623 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19099) );
  NOR2_X1 U16624 ( .A1(n13217), .A2(n13216), .ZN(n13220) );
  INV_X1 U16625 ( .A(n13218), .ZN(n13219) );
  OAI211_X1 U16626 ( .C1(n13220), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15298), .B(n13347), .ZN(n13225) );
  INV_X1 U16627 ( .A(n15269), .ZN(n15305) );
  OR2_X1 U16628 ( .A1(n13221), .A2(n13204), .ZN(n13223) );
  NAND2_X1 U16629 ( .A1(n13223), .A2(n13222), .ZN(n16294) );
  INV_X1 U16630 ( .A(n16294), .ZN(n19108) );
  NAND2_X1 U16631 ( .A1(n15305), .A2(n19108), .ZN(n13224) );
  OAI211_X1 U16632 ( .C1(n15302), .C2(n19099), .A(n13225), .B(n13224), .ZN(
        P2_U2881) );
  NAND2_X1 U16633 ( .A1(n13177), .A2(n20910), .ZN(n13332) );
  OR2_X1 U16634 ( .A1(n13332), .A2(n15981), .ZN(n15961) );
  AND2_X1 U16635 ( .A1(n13226), .A2(n15961), .ZN(n13228) );
  NOR2_X1 U16636 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16177), .ZN(n20125) );
  NOR2_X4 U16637 ( .A1(n13229), .A2(n20919), .ZN(n15983) );
  AOI22_X1 U16638 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13230) );
  OAI21_X1 U16639 ( .B1(n14803), .B2(n13555), .A(n13230), .ZN(P1_U2912) );
  INV_X1 U16640 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13232) );
  AOI22_X1 U16641 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13231) );
  OAI21_X1 U16642 ( .B1(n13232), .B2(n13555), .A(n13231), .ZN(P1_U2908) );
  INV_X1 U16643 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14830) );
  AOI22_X1 U16644 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20125), .B1(n15983), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13233) );
  OAI21_X1 U16645 ( .B1(n14830), .B2(n13555), .A(n13233), .ZN(P1_U2918) );
  INV_X1 U16646 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13235) );
  AOI22_X1 U16647 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13234) );
  OAI21_X1 U16648 ( .B1(n13235), .B2(n13555), .A(n13234), .ZN(P1_U2909) );
  INV_X1 U16649 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13237) );
  AOI22_X1 U16650 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13236) );
  OAI21_X1 U16651 ( .B1(n13237), .B2(n13555), .A(n13236), .ZN(P1_U2907) );
  INV_X1 U16652 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14839) );
  AOI22_X1 U16653 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20125), .B1(n15983), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13238) );
  OAI21_X1 U16654 ( .B1(n14839), .B2(n13555), .A(n13238), .ZN(P1_U2920) );
  INV_X1 U16655 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13240) );
  AOI22_X1 U16656 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13239) );
  OAI21_X1 U16657 ( .B1(n13240), .B2(n13555), .A(n13239), .ZN(P1_U2911) );
  AOI22_X1 U16658 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20125), .B1(n15983), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13241) );
  OAI21_X1 U16659 ( .B1(n14834), .B2(n13555), .A(n13241), .ZN(P1_U2919) );
  INV_X1 U16660 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13243) );
  AOI22_X1 U16661 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13242) );
  OAI21_X1 U16662 ( .B1(n13243), .B2(n13555), .A(n13242), .ZN(P1_U2917) );
  INV_X1 U16663 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13245) );
  AOI22_X1 U16664 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13244) );
  OAI21_X1 U16665 ( .B1(n13245), .B2(n13555), .A(n13244), .ZN(P1_U2913) );
  AND2_X1 U16666 ( .A1(n13246), .A2(n15980), .ZN(n13247) );
  OR2_X1 U16667 ( .A1(n20135), .A2(n20258), .ZN(n13386) );
  INV_X1 U16668 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13252) );
  NAND2_X1 U16669 ( .A1(n13452), .A2(n20258), .ZN(n13387) );
  INV_X1 U16670 ( .A(DATAI_15_), .ZN(n13250) );
  INV_X1 U16671 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13249) );
  MUX2_X1 U16672 ( .A(n13250), .B(n13249), .S(n20238), .Z(n14846) );
  INV_X1 U16673 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13251) );
  OAI222_X1 U16674 ( .A1(n13386), .A2(n13252), .B1(n13387), .B2(n14846), .C1(
        n13251), .C2(n13452), .ZN(P1_U2967) );
  OAI21_X1 U16675 ( .B1(n13254), .B2(n13253), .A(n13296), .ZN(n13651) );
  XNOR2_X1 U16676 ( .A(n13648), .B(n9658), .ZN(n20227) );
  AOI22_X1 U16677 ( .A1(n11194), .A2(n20227), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n14769), .ZN(n13255) );
  OAI21_X1 U16678 ( .B1(n13651), .B2(n14779), .A(n13255), .ZN(P1_U2871) );
  XOR2_X1 U16679 ( .A(n13257), .B(n13256), .Z(n13961) );
  INV_X1 U16680 ( .A(n13961), .ZN(n13265) );
  OR2_X1 U16681 ( .A1(n16363), .A2(n15836), .ZN(n13261) );
  NAND2_X1 U16682 ( .A1(n13259), .A2(n13258), .ZN(n13260) );
  OAI21_X4 U16683 ( .B1(n13755), .B2(n13263), .A(n13262), .ZN(n19188) );
  OR2_X1 U16684 ( .A1(n19188), .A2(n19288), .ZN(n16237) );
  AND2_X1 U16685 ( .A1(n19183), .A2(n16237), .ZN(n19174) );
  INV_X1 U16686 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19215) );
  OR2_X1 U16687 ( .A1(n19188), .A2(n12295), .ZN(n15381) );
  OR2_X1 U16688 ( .A1(n19188), .A2(n13264), .ZN(n13855) );
  OAI222_X1 U16689 ( .A1(n13265), .A2(n19174), .B1(n15380), .B2(n19215), .C1(
        n19196), .C2(n19290), .ZN(P2_U2912) );
  INV_X1 U16690 ( .A(n13266), .ZN(n13268) );
  NAND3_X1 U16691 ( .A1(n13783), .A2(n13268), .A3(n13267), .ZN(n13269) );
  NAND2_X1 U16692 ( .A1(n13270), .A2(n13269), .ZN(n19112) );
  INV_X1 U16693 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19217) );
  OAI222_X1 U16694 ( .A1(n19112), .A2(n19174), .B1(n15380), .B2(n19217), .C1(
        n19196), .C2(n19280), .ZN(P2_U2913) );
  XOR2_X1 U16695 ( .A(n13347), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13275)
         );
  AOI21_X1 U16696 ( .B1(n13272), .B2(n13222), .A(n13271), .ZN(n13613) );
  INV_X1 U16697 ( .A(n13613), .ZN(n13955) );
  MUX2_X1 U16698 ( .A(n13273), .B(n13955), .S(n15302), .Z(n13274) );
  OAI21_X1 U16699 ( .B1(n13275), .B2(n15312), .A(n13274), .ZN(P2_U2880) );
  INV_X1 U16700 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19210) );
  INV_X1 U16701 ( .A(n15343), .ZN(n13277) );
  OAI21_X1 U16702 ( .B1(n13583), .B2(n13276), .A(n13573), .ZN(n19093) );
  OAI222_X1 U16703 ( .A1(n15380), .A2(n19210), .B1(n13277), .B2(n19196), .C1(
        n19093), .C2(n19174), .ZN(P2_U2910) );
  OAI21_X1 U16704 ( .B1(n13278), .B2(n13571), .A(n15783), .ZN(n19078) );
  INV_X1 U16705 ( .A(n15327), .ZN(n13279) );
  INV_X1 U16706 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19206) );
  OAI222_X1 U16707 ( .A1(n19078), .A2(n19174), .B1(n13279), .B2(n19196), .C1(
        n19206), .C2(n15380), .ZN(P2_U2908) );
  NAND2_X1 U16708 ( .A1(n13280), .A2(n20289), .ZN(n13281) );
  INV_X1 U16709 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20124) );
  NAND2_X1 U16710 ( .A1(n20237), .A2(DATAI_1_), .ZN(n13283) );
  NAND2_X1 U16711 ( .A1(n20238), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13282) );
  AND2_X1 U16712 ( .A1(n13283), .A2(n13282), .ZN(n20259) );
  OAI222_X1 U16713 ( .A1(n14848), .A2(n13651), .B1(n14853), .B2(n20124), .C1(
        n14852), .C2(n20259), .ZN(P1_U2903) );
  INV_X1 U16714 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20128) );
  NAND2_X1 U16715 ( .A1(n20237), .A2(DATAI_0_), .ZN(n13285) );
  NAND2_X1 U16716 ( .A1(n20238), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13284) );
  AND2_X1 U16717 ( .A1(n13285), .A2(n13284), .ZN(n20251) );
  OAI222_X1 U16718 ( .A1(n14848), .A2(n14745), .B1(n14853), .B2(n20128), .C1(
        n14852), .C2(n20251), .ZN(P1_U2904) );
  NOR2_X1 U16719 ( .A1(n13286), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20223) );
  NOR2_X1 U16720 ( .A1(n20223), .A2(n20007), .ZN(n13289) );
  INV_X2 U16721 ( .A(n20064), .ZN(n20167) );
  AOI22_X1 U16722 ( .A1(n20168), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20167), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13287) );
  OAI21_X1 U16723 ( .B1(n20178), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13287), .ZN(n13288) );
  AOI21_X1 U16724 ( .B1(n13289), .B2(n20221), .A(n13288), .ZN(n13290) );
  OAI21_X1 U16725 ( .B1(n16049), .B2(n13651), .A(n13290), .ZN(P1_U2998) );
  OAI21_X1 U16726 ( .B1(n13293), .B2(n13292), .A(n13291), .ZN(n20203) );
  INV_X1 U16727 ( .A(n13294), .ZN(n13295) );
  AOI21_X1 U16728 ( .B1(n13297), .B2(n13296), .A(n13295), .ZN(n14728) );
  NAND2_X1 U16729 ( .A1(n20167), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n20200) );
  NAND2_X1 U16730 ( .A1(n20168), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13298) );
  OAI211_X1 U16731 ( .C1(n20178), .C2(n14729), .A(n20200), .B(n13298), .ZN(
        n13299) );
  AOI21_X1 U16732 ( .B1(n14728), .B2(n20239), .A(n13299), .ZN(n13300) );
  OAI21_X1 U16733 ( .B1(n20007), .B2(n20203), .A(n13300), .ZN(P1_U2997) );
  INV_X1 U16734 ( .A(n14728), .ZN(n13306) );
  INV_X1 U16735 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20122) );
  NAND2_X1 U16736 ( .A1(n20237), .A2(DATAI_2_), .ZN(n13302) );
  NAND2_X1 U16737 ( .A1(n20238), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13301) );
  AND2_X1 U16738 ( .A1(n13302), .A2(n13301), .ZN(n20264) );
  OAI222_X1 U16739 ( .A1(n14848), .A2(n13306), .B1(n14853), .B2(n20122), .C1(
        n14852), .C2(n20264), .ZN(P1_U2902) );
  NOR2_X1 U16740 ( .A1(n13304), .A2(n13303), .ZN(n13305) );
  OR2_X1 U16741 ( .A1(n13471), .A2(n13305), .ZN(n20199) );
  INV_X1 U16742 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13307) );
  OAI222_X1 U16743 ( .A1(n20199), .A2(n14777), .B1(n14778), .B2(n13307), .C1(
        n13306), .C2(n14779), .ZN(P1_U2870) );
  INV_X1 U16744 ( .A(n13308), .ZN(n13346) );
  AOI21_X1 U16745 ( .B1(n20258), .B2(n15981), .A(n15980), .ZN(n13309) );
  NAND2_X1 U16746 ( .A1(n14475), .A2(n13309), .ZN(n13317) );
  NAND2_X1 U16747 ( .A1(n13310), .A2(n15981), .ZN(n13633) );
  AND2_X1 U16748 ( .A1(n13633), .A2(n20918), .ZN(n13313) );
  NAND2_X1 U16749 ( .A1(n20244), .A2(n13311), .ZN(n13312) );
  AOI21_X1 U16750 ( .B1(n13177), .B2(n13313), .A(n13312), .ZN(n13314) );
  OR2_X1 U16751 ( .A1(n14483), .A2(n13314), .ZN(n13316) );
  MUX2_X1 U16752 ( .A(n13317), .B(n13316), .S(n13315), .Z(n13322) );
  INV_X1 U16753 ( .A(n13318), .ZN(n13320) );
  AOI21_X1 U16754 ( .B1(n14483), .B2(n13320), .A(n13319), .ZN(n13321) );
  NAND2_X1 U16755 ( .A1(n13322), .A2(n13321), .ZN(n13323) );
  OAI211_X1 U16756 ( .C1(n13329), .C2(n13324), .A(n14472), .B(n14471), .ZN(
        n13326) );
  OR2_X1 U16757 ( .A1(n13326), .A2(n13325), .ZN(n13327) );
  NAND3_X1 U16758 ( .A1(n13330), .A2(n13329), .A3(n13328), .ZN(n13331) );
  NAND2_X1 U16759 ( .A1(n13332), .A2(n13331), .ZN(n13333) );
  AND2_X2 U16760 ( .A1(n13340), .A2(n13333), .ZN(n20228) );
  INV_X1 U16761 ( .A(n14741), .ZN(n13344) );
  INV_X1 U16762 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15169) );
  OAI211_X1 U16763 ( .C1(n13336), .C2(n20244), .A(n13335), .B(n13334), .ZN(
        n13337) );
  NAND2_X1 U16764 ( .A1(n13340), .A2(n13337), .ZN(n15098) );
  NOR2_X1 U16765 ( .A1(n15098), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13339) );
  NOR2_X1 U16766 ( .A1(n13340), .A2(n20167), .ZN(n13338) );
  AOI21_X1 U16767 ( .B1(n20209), .B2(n15169), .A(n20214), .ZN(n20232) );
  NAND2_X1 U16768 ( .A1(n13340), .A2(n15166), .ZN(n15100) );
  NOR2_X1 U16769 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20209), .ZN(
        n13341) );
  AOI22_X1 U16770 ( .A1(n20232), .A2(n15100), .B1(n15098), .B2(n13341), .ZN(
        n13342) );
  AOI211_X1 U16771 ( .C1(n20228), .C2(n13344), .A(n13343), .B(n13342), .ZN(
        n13345) );
  OAI21_X1 U16772 ( .B1(n13346), .B2(n20222), .A(n13345), .ZN(P1_U3031) );
  INV_X1 U16773 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14302) );
  OAI211_X1 U16774 ( .C1(n9760), .C2(n13348), .A(n13508), .B(n15298), .ZN(
        n13352) );
  OR2_X1 U16775 ( .A1(n13349), .A2(n13271), .ZN(n13350) );
  AND2_X1 U16776 ( .A1(n13350), .A2(n13355), .ZN(n16330) );
  NAND2_X1 U16777 ( .A1(n15302), .A2(n16330), .ZN(n13351) );
  OAI211_X1 U16778 ( .C1(n15302), .C2(n13353), .A(n13352), .B(n13351), .ZN(
        P2_U2879) );
  INV_X1 U16779 ( .A(n13354), .ZN(n13511) );
  XNOR2_X1 U16780 ( .A(n13508), .B(n13511), .ZN(n13362) );
  NAND2_X1 U16781 ( .A1(n13356), .A2(n13355), .ZN(n13359) );
  INV_X1 U16782 ( .A(n13357), .ZN(n13358) );
  NAND2_X1 U16783 ( .A1(n13359), .A2(n13358), .ZN(n19092) );
  MUX2_X1 U16784 ( .A(n19092), .B(n13360), .S(n15269), .Z(n13361) );
  OAI21_X1 U16785 ( .B1(n13362), .B2(n15312), .A(n13361), .ZN(P2_U2878) );
  OAI21_X1 U16786 ( .B1(n13363), .B2(n13365), .A(n13364), .ZN(n16077) );
  INV_X1 U16787 ( .A(n13366), .ZN(n13658) );
  AOI21_X1 U16788 ( .B1(n13367), .B2(n13382), .A(n13658), .ZN(n20063) );
  AOI22_X1 U16789 ( .A1(n20063), .A2(n11194), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n14769), .ZN(n13368) );
  OAI21_X1 U16790 ( .B1(n16077), .B2(n14779), .A(n13368), .ZN(P1_U2867) );
  OAI21_X1 U16791 ( .B1(n13371), .B2(n13370), .A(n13369), .ZN(n20192) );
  XOR2_X1 U16792 ( .A(n13372), .B(n13373), .Z(n20100) );
  NAND2_X1 U16793 ( .A1(n20167), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n20189) );
  NAND2_X1 U16794 ( .A1(n20168), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13374) );
  OAI211_X1 U16795 ( .C1(n20178), .C2(n20090), .A(n20189), .B(n13374), .ZN(
        n13375) );
  AOI21_X1 U16796 ( .B1(n20100), .B2(n20239), .A(n13375), .ZN(n13376) );
  OAI21_X1 U16797 ( .B1(n20007), .B2(n20192), .A(n13376), .ZN(P1_U2996) );
  AND2_X1 U16798 ( .A1(n13378), .A2(n13377), .ZN(n13379) );
  OR2_X1 U16799 ( .A1(n13363), .A2(n13379), .ZN(n20076) );
  INV_X1 U16800 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13383) );
  NAND2_X1 U16801 ( .A1(n13469), .A2(n13380), .ZN(n13381) );
  NAND2_X1 U16802 ( .A1(n13382), .A2(n13381), .ZN(n20181) );
  OAI222_X1 U16803 ( .A1(n20076), .A2(n14779), .B1(n14778), .B2(n13383), .C1(
        n20181), .C2(n14777), .ZN(P1_U2868) );
  INV_X1 U16804 ( .A(n20100), .ZN(n13472) );
  INV_X1 U16805 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20120) );
  NAND2_X1 U16806 ( .A1(n20237), .A2(DATAI_3_), .ZN(n13385) );
  NAND2_X1 U16807 ( .A1(n20238), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13384) );
  AND2_X1 U16808 ( .A1(n13385), .A2(n13384), .ZN(n20268) );
  OAI222_X1 U16809 ( .A1(n14848), .A2(n13472), .B1(n14853), .B2(n20120), .C1(
        n14852), .C2(n20268), .ZN(P1_U2901) );
  AOI22_X1 U16810 ( .A1(n20164), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20159), .ZN(n13389) );
  INV_X1 U16811 ( .A(n20264), .ZN(n13388) );
  NAND2_X1 U16812 ( .A1(n20149), .A2(n13388), .ZN(n13461) );
  NAND2_X1 U16813 ( .A1(n13389), .A2(n13461), .ZN(P1_U2954) );
  AOI22_X1 U16814 ( .A1(n20164), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20159), .ZN(n13393) );
  INV_X1 U16815 ( .A(DATAI_6_), .ZN(n13391) );
  INV_X1 U16816 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n13390) );
  MUX2_X1 U16817 ( .A(n13391), .B(n13390), .S(n20238), .Z(n20281) );
  INV_X1 U16818 ( .A(n20281), .ZN(n13392) );
  NAND2_X1 U16819 ( .A1(n20149), .A2(n13392), .ZN(n13457) );
  NAND2_X1 U16820 ( .A1(n13393), .A2(n13457), .ZN(P1_U2958) );
  AOI22_X1 U16821 ( .A1(n20164), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20159), .ZN(n13395) );
  INV_X1 U16822 ( .A(n20268), .ZN(n13394) );
  NAND2_X1 U16823 ( .A1(n20149), .A2(n13394), .ZN(n13465) );
  NAND2_X1 U16824 ( .A1(n13395), .A2(n13465), .ZN(P1_U2955) );
  AOI22_X1 U16825 ( .A1(n20164), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20159), .ZN(n13399) );
  INV_X1 U16826 ( .A(DATAI_7_), .ZN(n13397) );
  INV_X1 U16827 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n13396) );
  MUX2_X1 U16828 ( .A(n13397), .B(n13396), .S(n20238), .Z(n20292) );
  INV_X1 U16829 ( .A(n20292), .ZN(n13398) );
  NAND2_X1 U16830 ( .A1(n20149), .A2(n13398), .ZN(n13463) );
  NAND2_X1 U16831 ( .A1(n13399), .A2(n13463), .ZN(P1_U2959) );
  AOI22_X1 U16832 ( .A1(n20164), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20159), .ZN(n13403) );
  INV_X1 U16833 ( .A(DATAI_5_), .ZN(n13401) );
  INV_X1 U16834 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n13400) );
  MUX2_X1 U16835 ( .A(n13401), .B(n13400), .S(n20238), .Z(n20276) );
  INV_X1 U16836 ( .A(n20276), .ZN(n13402) );
  NAND2_X1 U16837 ( .A1(n20149), .A2(n13402), .ZN(n13467) );
  NAND2_X1 U16838 ( .A1(n13403), .A2(n13467), .ZN(P1_U2957) );
  AOI22_X1 U16839 ( .A1(n20164), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20159), .ZN(n13406) );
  INV_X1 U16840 ( .A(DATAI_4_), .ZN(n13405) );
  NAND2_X1 U16841 ( .A1(n20238), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13404) );
  OAI21_X1 U16842 ( .B1(n20238), .B2(n13405), .A(n13404), .ZN(n14819) );
  NAND2_X1 U16843 ( .A1(n20149), .A2(n14819), .ZN(n13453) );
  NAND2_X1 U16844 ( .A1(n13406), .A2(n13453), .ZN(P1_U2956) );
  AOI22_X1 U16845 ( .A1(n20164), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20135), .ZN(n13408) );
  INV_X1 U16846 ( .A(n20251), .ZN(n13407) );
  NAND2_X1 U16847 ( .A1(n20149), .A2(n13407), .ZN(n13459) );
  NAND2_X1 U16848 ( .A1(n13408), .A2(n13459), .ZN(P1_U2952) );
  AOI22_X1 U16849 ( .A1(n20164), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20135), .ZN(n13410) );
  INV_X1 U16850 ( .A(n20259), .ZN(n13409) );
  NAND2_X1 U16851 ( .A1(n20149), .A2(n13409), .ZN(n13455) );
  NAND2_X1 U16852 ( .A1(n13410), .A2(n13455), .ZN(P1_U2953) );
  INV_X1 U16853 ( .A(n20401), .ZN(n20650) );
  NOR2_X1 U16854 ( .A1(n10454), .A2(n20650), .ZN(n13411) );
  XOR2_X1 U16855 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n13411), .Z(
        n20077) );
  INV_X1 U16856 ( .A(n20077), .ZN(n13412) );
  NOR2_X1 U16857 ( .A1(n13412), .A2(n13176), .ZN(n16173) );
  NAND2_X1 U16858 ( .A1(n15939), .A2(n16181), .ZN(n13414) );
  OAI21_X1 U16859 ( .B1(n16175), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13414), .ZN(
        n13413) );
  OAI21_X1 U16860 ( .B1(n16173), .B2(n13414), .A(n13413), .ZN(n15958) );
  INV_X1 U16861 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20008) );
  INV_X1 U16862 ( .A(n13439), .ZN(n15168) );
  NOR2_X1 U16863 ( .A1(n13439), .A2(n13417), .ZN(n13428) );
  XNOR2_X1 U16864 ( .A(n15163), .B(n10184), .ZN(n15175) );
  INV_X1 U16865 ( .A(n15166), .ZN(n13420) );
  XNOR2_X1 U16866 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13419) );
  INV_X1 U16867 ( .A(n14471), .ZN(n13418) );
  NOR2_X1 U16868 ( .A1(n14474), .A2(n13418), .ZN(n13430) );
  OAI22_X1 U16869 ( .A1(n13420), .A2(n13419), .B1(n15175), .B2(n13430), .ZN(
        n13421) );
  AOI21_X1 U16870 ( .B1(n13428), .B2(n15175), .A(n13421), .ZN(n13422) );
  OAI21_X1 U16871 ( .B1(n13416), .B2(n15168), .A(n13422), .ZN(n15179) );
  MUX2_X1 U16872 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n15179), .S(
        n15939), .Z(n15946) );
  NOR2_X1 U16873 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n16181), .ZN(n13441) );
  AOI22_X1 U16874 ( .A1(n15946), .A2(n16181), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n13441), .ZN(n13443) );
  NOR2_X1 U16875 ( .A1(n15163), .A2(n9920), .ZN(n13426) );
  NOR2_X1 U16876 ( .A1(n13426), .A2(n13425), .ZN(n13427) );
  NAND2_X1 U16877 ( .A1(n10382), .A2(n13427), .ZN(n15183) );
  NAND2_X1 U16878 ( .A1(n13428), .A2(n15183), .ZN(n13437) );
  XNOR2_X1 U16879 ( .A(n13429), .B(n9920), .ZN(n13435) );
  INV_X1 U16880 ( .A(n13430), .ZN(n13434) );
  MUX2_X1 U16881 ( .A(n10193), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15163), .Z(n13432) );
  NOR2_X1 U16882 ( .A1(n13432), .A2(n13431), .ZN(n13433) );
  AOI22_X1 U16883 ( .A1(n15166), .A2(n13435), .B1(n13434), .B2(n13433), .ZN(
        n13436) );
  NAND2_X1 U16884 ( .A1(n13437), .A2(n13436), .ZN(n13438) );
  AOI21_X1 U16885 ( .B1(n13423), .B2(n13439), .A(n13438), .ZN(n15185) );
  MUX2_X1 U16886 ( .A(n9920), .B(n15185), .S(n15939), .Z(n13440) );
  AOI22_X1 U16887 ( .A1(n13441), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n16181), .B2(n15949), .ZN(n13442) );
  NOR2_X1 U16888 ( .A1(n13443), .A2(n13442), .ZN(n15956) );
  INV_X1 U16889 ( .A(n10190), .ZN(n13444) );
  NAND2_X1 U16890 ( .A1(n15956), .A2(n13444), .ZN(n13446) );
  AND3_X1 U16891 ( .A1(n15958), .A2(n20008), .A3(n13446), .ZN(n13445) );
  NAND2_X1 U16892 ( .A1(n20837), .A2(n16181), .ZN(n20913) );
  INV_X1 U16893 ( .A(n20913), .ZN(n15967) );
  INV_X1 U16894 ( .A(n20299), .ZN(n20406) );
  NAND3_X1 U16895 ( .A1(n15958), .A2(n13447), .A3(n13446), .ZN(n15971) );
  INV_X1 U16896 ( .A(n15971), .ZN(n13450) );
  INV_X1 U16897 ( .A(n10445), .ZN(n14739) );
  NAND2_X1 U16898 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20525), .ZN(n15158) );
  INV_X1 U16899 ( .A(n15158), .ZN(n13448) );
  OAI22_X1 U16900 ( .A1(n20326), .A2(n20781), .B1(n14739), .B2(n13448), .ZN(
        n13449) );
  OAI21_X1 U16901 ( .B1(n13450), .B2(n13449), .A(n20235), .ZN(n13451) );
  OAI21_X1 U16902 ( .B1(n20235), .B2(n20692), .A(n13451), .ZN(P1_U3478) );
  AOI22_X1 U16903 ( .A1(n20164), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20135), .ZN(n13454) );
  NAND2_X1 U16904 ( .A1(n13454), .A2(n13453), .ZN(P1_U2941) );
  AOI22_X1 U16905 ( .A1(n20164), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20159), .ZN(n13456) );
  NAND2_X1 U16906 ( .A1(n13456), .A2(n13455), .ZN(P1_U2938) );
  AOI22_X1 U16907 ( .A1(n20164), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20159), .ZN(n13458) );
  NAND2_X1 U16908 ( .A1(n13458), .A2(n13457), .ZN(P1_U2943) );
  AOI22_X1 U16909 ( .A1(n20164), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20159), .ZN(n13460) );
  NAND2_X1 U16910 ( .A1(n13460), .A2(n13459), .ZN(P1_U2937) );
  AOI22_X1 U16911 ( .A1(n20164), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20159), .ZN(n13462) );
  NAND2_X1 U16912 ( .A1(n13462), .A2(n13461), .ZN(P1_U2939) );
  AOI22_X1 U16913 ( .A1(n20164), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20159), .ZN(n13464) );
  NAND2_X1 U16914 ( .A1(n13464), .A2(n13463), .ZN(P1_U2944) );
  AOI22_X1 U16915 ( .A1(n20164), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20159), .ZN(n13466) );
  NAND2_X1 U16916 ( .A1(n13466), .A2(n13465), .ZN(P1_U2940) );
  AOI22_X1 U16917 ( .A1(n20164), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20159), .ZN(n13468) );
  NAND2_X1 U16918 ( .A1(n13468), .A2(n13467), .ZN(P1_U2942) );
  INV_X1 U16919 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20116) );
  OAI222_X1 U16920 ( .A1(n14848), .A2(n16077), .B1(n14853), .B2(n20116), .C1(
        n14852), .C2(n20276), .ZN(P1_U2899) );
  OAI21_X1 U16921 ( .B1(n13471), .B2(n13470), .A(n13469), .ZN(n20087) );
  INV_X1 U16922 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13473) );
  OAI222_X1 U16923 ( .A1(n20087), .A2(n14777), .B1(n13473), .B2(n14778), .C1(
        n13472), .C2(n14779), .ZN(P1_U2869) );
  INV_X1 U16924 ( .A(n20235), .ZN(n13483) );
  INV_X1 U16925 ( .A(n9677), .ZN(n13475) );
  OR2_X1 U16926 ( .A1(n9677), .A2(n21034), .ZN(n20548) );
  OAI21_X1 U16927 ( .B1(n13475), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20548), 
        .ZN(n13477) );
  AOI22_X1 U16928 ( .A1(n13477), .A2(n20783), .B1(n9665), .B2(n15158), .ZN(
        n13479) );
  NAND2_X1 U16929 ( .A1(n13483), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13478) );
  OAI21_X1 U16930 ( .B1(n13483), .B2(n13479), .A(n13478), .ZN(P1_U3477) );
  NAND2_X1 U16931 ( .A1(n9677), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20777) );
  XNOR2_X1 U16932 ( .A(n15155), .B(n20777), .ZN(n13480) );
  INV_X1 U16933 ( .A(n13416), .ZN(n20247) );
  AOI22_X1 U16934 ( .A1(n13480), .A2(n20783), .B1(n20247), .B2(n15158), .ZN(
        n13482) );
  NAND2_X1 U16935 ( .A1(n13483), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13481) );
  OAI21_X1 U16936 ( .B1(n13483), .B2(n13482), .A(n13481), .ZN(P1_U3476) );
  XNOR2_X1 U16937 ( .A(n13485), .B(n13500), .ZN(n13486) );
  XNOR2_X1 U16938 ( .A(n13484), .B(n13486), .ZN(n13505) );
  XNOR2_X1 U16939 ( .A(n13487), .B(n13488), .ZN(n13503) );
  NOR2_X1 U16940 ( .A1(n19113), .A2(n11430), .ZN(n13494) );
  NOR2_X1 U16941 ( .A1(n16310), .A2(n12785), .ZN(n13489) );
  AOI211_X1 U16942 ( .C1(n13538), .C2(n16301), .A(n13494), .B(n13489), .ZN(
        n13490) );
  OAI21_X1 U16943 ( .B1(n13138), .B2(n13736), .A(n13490), .ZN(n13491) );
  AOI21_X1 U16944 ( .B1(n13503), .B2(n19236), .A(n13491), .ZN(n13492) );
  OAI21_X1 U16945 ( .B1(n13505), .B2(n11993), .A(n13492), .ZN(P2_U3011) );
  XNOR2_X1 U16946 ( .A(n13493), .B(n9763), .ZN(n19936) );
  INV_X1 U16947 ( .A(n19936), .ZN(n13719) );
  AOI21_X1 U16948 ( .B1(n16331), .B2(n15859), .A(n13494), .ZN(n13495) );
  OAI21_X1 U16949 ( .B1(n13719), .B2(n15816), .A(n13495), .ZN(n13502) );
  AOI21_X1 U16950 ( .B1(n15705), .B2(n13497), .A(n13496), .ZN(n13600) );
  NAND2_X1 U16951 ( .A1(n13500), .A2(n15798), .ZN(n13498) );
  OAI22_X1 U16952 ( .A1(n13600), .A2(n13500), .B1(n13499), .B2(n13498), .ZN(
        n13501) );
  AOI211_X1 U16953 ( .C1(n13503), .C2(n16328), .A(n13502), .B(n13501), .ZN(
        n13504) );
  OAI21_X1 U16954 ( .B1(n13505), .B2(n16320), .A(n13504), .ZN(P2_U3043) );
  INV_X1 U16955 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19202) );
  INV_X1 U16956 ( .A(n15315), .ZN(n13507) );
  OAI21_X1 U16957 ( .B1(n15782), .B2(n13506), .A(n15748), .ZN(n19056) );
  OAI222_X1 U16958 ( .A1(n15380), .A2(n19202), .B1(n13507), .B2(n19196), .C1(
        n19056), .C2(n19174), .ZN(P2_U2906) );
  OAI21_X1 U16959 ( .B1(n13508), .B2(n13511), .A(n13510), .ZN(n13514) );
  NAND3_X1 U16960 ( .A1(n13514), .A2(n15298), .A3(n13618), .ZN(n13518) );
  OR2_X1 U16961 ( .A1(n13515), .A2(n13357), .ZN(n13516) );
  AND2_X1 U16962 ( .A1(n13516), .A2(n9756), .ZN(n16316) );
  NAND2_X1 U16963 ( .A1(n15302), .A2(n16316), .ZN(n13517) );
  OAI211_X1 U16964 ( .C1(n15302), .C2(n13519), .A(n13518), .B(n13517), .ZN(
        P2_U2877) );
  XNOR2_X1 U16965 ( .A(n19942), .B(n13718), .ZN(n13526) );
  INV_X1 U16966 ( .A(n19954), .ZN(n13522) );
  NAND2_X1 U16967 ( .A1(n19949), .A2(n13522), .ZN(n13523) );
  OAI21_X1 U16968 ( .B1(n19949), .B2(n13522), .A(n13523), .ZN(n19182) );
  NOR2_X1 U16969 ( .A1(n19961), .A2(n19128), .ZN(n19190) );
  NOR2_X1 U16970 ( .A1(n19182), .A2(n19190), .ZN(n19181) );
  INV_X1 U16971 ( .A(n13523), .ZN(n13524) );
  NOR2_X1 U16972 ( .A1(n19181), .A2(n13524), .ZN(n13525) );
  NOR2_X1 U16973 ( .A1(n13525), .A2(n13526), .ZN(n13717) );
  AOI21_X1 U16974 ( .B1(n13526), .B2(n13525), .A(n13717), .ZN(n13529) );
  AOI22_X1 U16975 ( .A1(n19167), .A2(n16234), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19188), .ZN(n13528) );
  NAND2_X1 U16976 ( .A1(n19944), .A2(n19189), .ZN(n13527) );
  OAI211_X1 U16977 ( .C1(n13529), .C2(n19183), .A(n13528), .B(n13527), .ZN(
        P2_U2917) );
  INV_X1 U16978 ( .A(n13531), .ZN(n13532) );
  NAND2_X1 U16979 ( .A1(n13364), .A2(n13532), .ZN(n13533) );
  AND2_X1 U16980 ( .A1(n13530), .A2(n13533), .ZN(n20059) );
  INV_X1 U16981 ( .A(n20059), .ZN(n13535) );
  INV_X1 U16982 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n13534) );
  XNOR2_X1 U16983 ( .A(n13658), .B(n13657), .ZN(n16159) );
  OAI222_X1 U16984 ( .A1(n14779), .A2(n13535), .B1(n13534), .B2(n14778), .C1(
        n14777), .C2(n16159), .ZN(P1_U2866) );
  OAI222_X1 U16985 ( .A1(n14848), .A2(n13535), .B1(n14853), .B2(n10546), .C1(
        n14852), .C2(n20281), .ZN(P1_U2898) );
  NAND2_X1 U16986 ( .A1(n12794), .A2(n13536), .ZN(n13537) );
  XNOR2_X1 U16987 ( .A(n13538), .B(n13537), .ZN(n13539) );
  NAND2_X1 U16988 ( .A1(n13539), .A2(n19123), .ZN(n13546) );
  OAI22_X1 U16989 ( .A1(n19100), .A2(n11648), .B1(n19127), .B2(n13719), .ZN(
        n13541) );
  NOR2_X1 U16990 ( .A1(n19133), .A2(n11430), .ZN(n13540) );
  AOI211_X1 U16991 ( .C1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .C2(n19142), .A(
        n13541), .B(n13540), .ZN(n13542) );
  OAI21_X1 U16992 ( .B1(n13543), .B2(n19101), .A(n13542), .ZN(n13544) );
  AOI21_X1 U16993 ( .B1(n15859), .B2(n19122), .A(n13544), .ZN(n13545) );
  OAI211_X1 U16994 ( .C1(n13683), .C2(n19934), .A(n13546), .B(n13545), .ZN(
        P2_U2852) );
  INV_X1 U16995 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13548) );
  AOI22_X1 U16996 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13547) );
  OAI21_X1 U16997 ( .B1(n13548), .B2(n13555), .A(n13547), .ZN(P1_U2916) );
  INV_X1 U16998 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13550) );
  AOI22_X1 U16999 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13549) );
  OAI21_X1 U17000 ( .B1(n13550), .B2(n13555), .A(n13549), .ZN(P1_U2914) );
  INV_X1 U17001 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13552) );
  AOI22_X1 U17002 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13551) );
  OAI21_X1 U17003 ( .B1(n13552), .B2(n13555), .A(n13551), .ZN(P1_U2915) );
  AOI22_X1 U17004 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13553) );
  OAI21_X1 U17005 ( .B1(n14794), .B2(n13555), .A(n13553), .ZN(P1_U2910) );
  INV_X1 U17006 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13556) );
  AOI22_X1 U17007 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20919), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n15983), .ZN(n13554) );
  OAI21_X1 U17008 ( .B1(n13556), .B2(n13555), .A(n13554), .ZN(P1_U2906) );
  INV_X1 U17009 ( .A(n19239), .ZN(n13560) );
  NOR2_X1 U17010 ( .A1(n19105), .A2(n13557), .ZN(n13559) );
  AOI21_X1 U17011 ( .B1(n13560), .B2(n13559), .A(n19851), .ZN(n13558) );
  OAI21_X1 U17012 ( .B1(n13560), .B2(n13559), .A(n13558), .ZN(n13569) );
  OAI21_X1 U17013 ( .B1(n19133), .B2(n11860), .A(n19113), .ZN(n13561) );
  AOI21_X1 U17014 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n19135), .A(n13561), .ZN(
        n13562) );
  OAI21_X1 U17015 ( .B1(n13563), .B2(n19101), .A(n13562), .ZN(n13567) );
  XNOR2_X1 U17016 ( .A(n13565), .B(n13564), .ZN(n13722) );
  OAI22_X1 U17017 ( .A1(n11859), .A2(n19073), .B1(n19127), .B2(n13722), .ZN(
        n13566) );
  AOI211_X1 U17018 ( .C1(n13602), .C2(n19122), .A(n13567), .B(n13566), .ZN(
        n13568) );
  OAI211_X1 U17019 ( .C1(n19168), .C2(n13683), .A(n13569), .B(n13568), .ZN(
        P2_U2851) );
  INV_X1 U17020 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20118) );
  INV_X1 U17021 ( .A(n14819), .ZN(n20272) );
  OAI222_X1 U17022 ( .A1(n20076), .A2(n14848), .B1(n20118), .B2(n14853), .C1(
        n14852), .C2(n20272), .ZN(P1_U2900) );
  OAI222_X1 U17023 ( .A1(n15736), .A2(n19174), .B1(n15380), .B2(n12966), .C1(
        n13570), .C2(n19196), .ZN(P2_U2904) );
  AOI21_X1 U17024 ( .B1(n13573), .B2(n13572), .A(n13571), .ZN(n19158) );
  NOR2_X1 U17025 ( .A1(n19105), .A2(n13574), .ZN(n13575) );
  XNOR2_X1 U17026 ( .A(n13575), .B(n16277), .ZN(n13576) );
  AOI22_X1 U17027 ( .A1(n19129), .A2(n19158), .B1(n19123), .B2(n13576), .ZN(
        n13581) );
  AOI22_X1 U17028 ( .A1(P2_EBX_REG_10__SCAN_IN), .A2(n19135), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19142), .ZN(n13577) );
  OAI211_X1 U17029 ( .C1(n19133), .C2(n13578), .A(n13577), .B(n19113), .ZN(
        n13579) );
  AOI21_X1 U17030 ( .B1(n16316), .B2(n19122), .A(n13579), .ZN(n13580) );
  OAI211_X1 U17031 ( .C1(n13582), .C2(n19101), .A(n13581), .B(n13580), .ZN(
        P2_U2845) );
  AOI21_X1 U17032 ( .B1(n13585), .B2(n13584), .A(n13583), .ZN(n19162) );
  NOR2_X1 U17033 ( .A1(n19105), .A2(n13586), .ZN(n13587) );
  XNOR2_X1 U17034 ( .A(n13587), .B(n16293), .ZN(n13588) );
  AOI22_X1 U17035 ( .A1(n19129), .A2(n19162), .B1(n19123), .B2(n13588), .ZN(
        n13593) );
  AOI22_X1 U17036 ( .A1(P2_EBX_REG_8__SCAN_IN), .A2(n19135), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19142), .ZN(n13589) );
  OAI211_X1 U17037 ( .C1(n19133), .C2(n13590), .A(n13589), .B(n19113), .ZN(
        n13591) );
  AOI21_X1 U17038 ( .B1(n16330), .B2(n19122), .A(n13591), .ZN(n13592) );
  OAI211_X1 U17039 ( .C1(n13594), .C2(n19101), .A(n13593), .B(n13592), .ZN(
        P2_U2847) );
  XNOR2_X1 U17040 ( .A(n13595), .B(n13596), .ZN(n19233) );
  NAND2_X1 U17041 ( .A1(n13598), .A2(n13597), .ZN(n13599) );
  XNOR2_X1 U17042 ( .A(n13599), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19235) );
  OAI21_X1 U17043 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15710), .A(
        n13600), .ZN(n13931) );
  NOR2_X1 U17044 ( .A1(n11860), .A2(n19113), .ZN(n13601) );
  AOI221_X1 U17045 ( .B1(n13957), .B2(n13788), .C1(n13931), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n13601), .ZN(n13604) );
  NAND2_X1 U17046 ( .A1(n13602), .A2(n16331), .ZN(n13603) );
  OAI211_X1 U17047 ( .C1(n15816), .C2(n13722), .A(n13604), .B(n13603), .ZN(
        n13605) );
  AOI21_X1 U17048 ( .B1(n16328), .B2(n19235), .A(n13605), .ZN(n13606) );
  OAI21_X1 U17049 ( .B1(n19233), .B2(n16320), .A(n13606), .ZN(P2_U3042) );
  INV_X1 U17050 ( .A(n13607), .ZN(n13616) );
  NAND2_X1 U17051 ( .A1(n12794), .A2(n13608), .ZN(n13609) );
  XNOR2_X1 U17052 ( .A(n13950), .B(n13609), .ZN(n13610) );
  AOI22_X1 U17053 ( .A1(n19129), .A2(n13961), .B1(n19123), .B2(n13610), .ZN(
        n13615) );
  INV_X1 U17054 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19879) );
  AOI22_X1 U17055 ( .A1(P2_EBX_REG_7__SCAN_IN), .A2(n19135), .B1(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19142), .ZN(n13611) );
  OAI211_X1 U17056 ( .C1(n19133), .C2(n19879), .A(n13611), .B(n19113), .ZN(
        n13612) );
  AOI21_X1 U17057 ( .B1(n13613), .B2(n19122), .A(n13612), .ZN(n13614) );
  OAI211_X1 U17058 ( .C1(n13616), .C2(n19101), .A(n13615), .B(n13614), .ZN(
        P2_U2848) );
  INV_X1 U17059 ( .A(n13618), .ZN(n13621) );
  INV_X1 U17060 ( .A(n13668), .ZN(n13619) );
  OAI211_X1 U17061 ( .C1(n13621), .C2(n13620), .A(n13619), .B(n15298), .ZN(
        n13626) );
  AND2_X1 U17062 ( .A1(n9756), .A2(n13622), .ZN(n13624) );
  NAND2_X1 U17063 ( .A1(n10163), .A2(n15305), .ZN(n13625) );
  OAI211_X1 U17064 ( .C1(n15305), .C2(n11705), .A(n13626), .B(n13625), .ZN(
        P2_U2876) );
  NAND2_X1 U17065 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n15967), .ZN(n15963) );
  AND2_X1 U17066 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20914), .ZN(n13627) );
  NAND2_X1 U17067 ( .A1(n13628), .A2(n13627), .ZN(n13629) );
  OAI211_X1 U17068 ( .C1(n15963), .C2(n20914), .A(n20225), .B(n13629), .ZN(
        n13630) );
  OAI21_X1 U17069 ( .B1(n13644), .B2(n14482), .A(n20029), .ZN(n20099) );
  INV_X1 U17070 ( .A(n20099), .ZN(n14746) );
  AND2_X1 U17071 ( .A1(n20918), .A2(n21034), .ZN(n13637) );
  AND2_X1 U17072 ( .A1(n13633), .A2(n13637), .ZN(n13635) );
  INV_X1 U17073 ( .A(n20044), .ZN(n20051) );
  INV_X1 U17074 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20855) );
  NAND2_X1 U17075 ( .A1(n20258), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13638) );
  INV_X1 U17076 ( .A(n13638), .ZN(n13634) );
  NOR2_X1 U17077 ( .A1(n13635), .A2(n13634), .ZN(n13636) );
  AOI22_X1 U17078 ( .A1(n20051), .A2(n20855), .B1(n20088), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13650) );
  NOR2_X1 U17079 ( .A1(n13638), .A2(n13637), .ZN(n13639) );
  NOR2_X1 U17080 ( .A1(n13641), .A2(n16181), .ZN(n13642) );
  NOR2_X1 U17081 ( .A1(n13644), .A2(n13643), .ZN(n20094) );
  NAND2_X1 U17082 ( .A1(n9665), .A2(n20094), .ZN(n13646) );
  INV_X1 U17083 ( .A(n14727), .ZN(n14498) );
  AOI22_X1 U17084 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n14498), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13645) );
  OAI211_X1 U17085 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20078), .A(
        n13646), .B(n13645), .ZN(n13647) );
  AOI21_X1 U17086 ( .B1(n20089), .B2(n13648), .A(n13647), .ZN(n13649) );
  OAI211_X1 U17087 ( .C1(n13651), .C2(n14746), .A(n13650), .B(n13649), .ZN(
        P1_U2839) );
  NAND2_X1 U17088 ( .A1(n13530), .A2(n13653), .ZN(n13654) );
  AND2_X1 U17089 ( .A1(n13652), .A2(n13654), .ZN(n20046) );
  INV_X1 U17090 ( .A(n20046), .ZN(n13655) );
  OAI222_X1 U17091 ( .A1(n14848), .A2(n13655), .B1(n14853), .B2(n10564), .C1(
        n14852), .C2(n20292), .ZN(P1_U2897) );
  AOI21_X1 U17092 ( .B1(n13658), .B2(n13657), .A(n13656), .ZN(n13659) );
  OR2_X1 U17093 ( .A1(n13659), .A2(n13696), .ZN(n16152) );
  OAI22_X1 U17094 ( .A1(n16152), .A2(n14777), .B1(n13660), .B2(n14778), .ZN(
        n13661) );
  AOI21_X1 U17095 ( .B1(n20046), .B2(n13662), .A(n13661), .ZN(n13663) );
  INV_X1 U17096 ( .A(n13663), .ZN(P1_U2865) );
  NOR2_X1 U17097 ( .A1(n13623), .A2(n13665), .ZN(n13666) );
  OR2_X1 U17098 ( .A1(n13664), .A2(n13666), .ZN(n16255) );
  OAI211_X1 U17099 ( .C1(n13668), .C2(n13667), .A(n13708), .B(n15298), .ZN(
        n13670) );
  NAND2_X1 U17100 ( .A1(n15269), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13669) );
  OAI211_X1 U17101 ( .C1(n16255), .C2(n15269), .A(n13670), .B(n13669), .ZN(
        P2_U2875) );
  INV_X1 U17102 ( .A(n14461), .ZN(n13673) );
  NOR2_X1 U17103 ( .A1(n19105), .A2(n13671), .ZN(n13767) );
  INV_X1 U17104 ( .A(n13767), .ZN(n13672) );
  AOI221_X1 U17105 ( .B1(n13673), .B2(n13767), .C1(n14461), .C2(n13672), .A(
        n19851), .ZN(n13674) );
  INV_X1 U17106 ( .A(n13674), .ZN(n13682) );
  AOI22_X1 U17107 ( .A1(P2_EBX_REG_2__SCAN_IN), .A2(n19135), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n19076), .ZN(n13676) );
  NAND2_X1 U17108 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19142), .ZN(
        n13675) );
  OAI211_X1 U17109 ( .C1(n13677), .C2(n19101), .A(n13676), .B(n13675), .ZN(
        n13679) );
  NOR2_X1 U17110 ( .A1(n13718), .A2(n19127), .ZN(n13678) );
  AOI211_X1 U17111 ( .C1(n19122), .C2(n13680), .A(n13679), .B(n13678), .ZN(
        n13681) );
  OAI211_X1 U17112 ( .C1(n19942), .C2(n13683), .A(n13682), .B(n13681), .ZN(
        P2_U2853) );
  XOR2_X1 U17113 ( .A(n13708), .B(n13709), .Z(n13689) );
  INV_X1 U17114 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n13687) );
  OR2_X1 U17115 ( .A1(n13664), .A2(n13685), .ZN(n13686) );
  AND2_X1 U17116 ( .A1(n13684), .A2(n13686), .ZN(n16250) );
  INV_X1 U17117 ( .A(n16250), .ZN(n19055) );
  MUX2_X1 U17118 ( .A(n13687), .B(n19055), .S(n15302), .Z(n13688) );
  OAI21_X1 U17119 ( .B1(n13689), .B2(n15312), .A(n13688), .ZN(P2_U2874) );
  INV_X1 U17120 ( .A(n13691), .ZN(n13692) );
  AOI21_X1 U17121 ( .B1(n13693), .B2(n13652), .A(n13692), .ZN(n13803) );
  INV_X1 U17122 ( .A(n13803), .ZN(n13706) );
  INV_X1 U17123 ( .A(n13801), .ZN(n13702) );
  INV_X1 U17124 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20866) );
  NAND2_X1 U17125 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n14726) );
  NAND2_X1 U17126 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .ZN(n20052) );
  NAND2_X1 U17127 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20041) );
  NOR3_X1 U17128 ( .A1(n14726), .A2(n20052), .A3(n20041), .ZN(n20039) );
  NAND2_X1 U17129 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20039), .ZN(n13699) );
  NOR2_X1 U17130 ( .A1(n20866), .A2(n13699), .ZN(n14495) );
  INV_X1 U17131 ( .A(n14495), .ZN(n14704) );
  NAND2_X1 U17132 ( .A1(n20044), .A2(n14727), .ZN(n20042) );
  OAI21_X1 U17133 ( .B1(n14498), .B2(n14704), .A(n20042), .ZN(n20026) );
  AOI22_X1 U17134 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n20091), .B1(
        P1_EBX_REG_8__SCAN_IN), .B2(n20088), .ZN(n13694) );
  OAI211_X1 U17135 ( .C1(n20026), .C2(n20866), .A(n13694), .B(n20064), .ZN(
        n13701) );
  OR2_X1 U17136 ( .A1(n13696), .A2(n13695), .ZN(n13697) );
  NAND2_X1 U17137 ( .A1(n13746), .A2(n13697), .ZN(n16145) );
  NAND2_X1 U17138 ( .A1(n20051), .A2(n14704), .ZN(n13698) );
  OAI22_X1 U17139 ( .A1(n20086), .A2(n16145), .B1(n13699), .B2(n13698), .ZN(
        n13700) );
  AOI211_X1 U17140 ( .C1(n20093), .C2(n13702), .A(n13701), .B(n13700), .ZN(
        n13703) );
  OAI21_X1 U17141 ( .B1(n13706), .B2(n20029), .A(n13703), .ZN(P1_U2832) );
  INV_X1 U17142 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13704) );
  OAI222_X1 U17143 ( .A1(n13706), .A2(n14779), .B1(n14778), .B2(n13704), .C1(
        n16145), .C2(n14777), .ZN(P1_U2864) );
  INV_X1 U17144 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13705) );
  INV_X1 U17145 ( .A(DATAI_8_), .ZN(n21119) );
  MUX2_X1 U17146 ( .A(n21119), .B(n16488), .S(n20238), .Z(n20129) );
  OAI222_X1 U17147 ( .A1(n13706), .A2(n14848), .B1(n13705), .B2(n14853), .C1(
        n14852), .C2(n20129), .ZN(P1_U2896) );
  INV_X1 U17148 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n19042) );
  INV_X1 U17149 ( .A(n13709), .ZN(n13707) );
  NOR2_X1 U17150 ( .A1(n13708), .A2(n13707), .ZN(n13711) );
  OAI211_X1 U17151 ( .C1(n13711), .C2(n13710), .A(n15298), .B(n13817), .ZN(
        n13716) );
  NAND2_X1 U17152 ( .A1(n13684), .A2(n13712), .ZN(n13713) );
  AND2_X1 U17153 ( .A1(n13714), .A2(n13713), .ZN(n19044) );
  NAND2_X1 U17154 ( .A1(n19044), .A2(n15302), .ZN(n13715) );
  OAI211_X1 U17155 ( .C1(n15302), .C2(n19042), .A(n13716), .B(n13715), .ZN(
        P2_U2873) );
  AOI21_X1 U17156 ( .B1(n13718), .B2(n19942), .A(n13717), .ZN(n19176) );
  XNOR2_X1 U17157 ( .A(n13719), .B(n19934), .ZN(n19177) );
  NOR2_X1 U17158 ( .A1(n19176), .A2(n19177), .ZN(n19175) );
  INV_X1 U17159 ( .A(n19934), .ZN(n13720) );
  NOR2_X1 U17160 ( .A1(n13720), .A2(n19936), .ZN(n13721) );
  OAI21_X1 U17161 ( .B1(n19175), .B2(n13721), .A(n13722), .ZN(n19170) );
  XOR2_X1 U17162 ( .A(n19168), .B(n19170), .Z(n13726) );
  INV_X1 U17163 ( .A(n13722), .ZN(n13723) );
  AOI22_X1 U17164 ( .A1(n19189), .A2(n13723), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19188), .ZN(n13725) );
  INV_X1 U17165 ( .A(n19270), .ZN(n16229) );
  NAND2_X1 U17166 ( .A1(n19167), .A2(n16229), .ZN(n13724) );
  OAI211_X1 U17167 ( .C1(n13726), .C2(n19183), .A(n13725), .B(n13724), .ZN(
        P2_U2915) );
  NOR2_X1 U17168 ( .A1(n19934), .A2(n19643), .ZN(n19777) );
  NAND2_X1 U17169 ( .A1(n19777), .A2(n10178), .ZN(n13727) );
  NAND3_X1 U17170 ( .A1(n19956), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19646) );
  NAND2_X1 U17171 ( .A1(n13727), .A2(n19646), .ZN(n13732) );
  NOR2_X1 U17172 ( .A1(n19966), .A2(n19646), .ZN(n19718) );
  INV_X1 U17173 ( .A(n19718), .ZN(n19707) );
  NAND2_X1 U17174 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19707), .ZN(n13728) );
  NOR2_X1 U17175 ( .A1(n11555), .A2(n13728), .ZN(n13735) );
  NAND2_X1 U17176 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19707), .ZN(n13729) );
  NAND2_X1 U17177 ( .A1(n19781), .A2(n13729), .ZN(n13730) );
  NOR2_X1 U17178 ( .A1(n13735), .A2(n13730), .ZN(n13731) );
  NAND2_X1 U17179 ( .A1(n13732), .A2(n13731), .ZN(n19711) );
  INV_X1 U17180 ( .A(n19711), .ZN(n19686) );
  INV_X1 U17181 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13741) );
  INV_X1 U17182 ( .A(n19646), .ZN(n13733) );
  AOI21_X1 U17183 ( .B1(n19645), .B2(n13733), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13734) );
  OR2_X1 U17184 ( .A1(n13735), .A2(n13734), .ZN(n19708) );
  INV_X1 U17185 ( .A(n19708), .ZN(n13739) );
  NOR2_X2 U17186 ( .A1(n19187), .A2(n19466), .ZN(n19732) );
  NAND2_X1 U17187 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19781), .ZN(n19274) );
  NOR2_X2 U17188 ( .A1(n11551), .A2(n19274), .ZN(n19730) );
  INV_X1 U17189 ( .A(n19730), .ZN(n19788) );
  AOI22_X1 U17190 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19292), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19291), .ZN(n19735) );
  INV_X1 U17191 ( .A(n19703), .ZN(n19710) );
  AOI22_X1 U17192 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19292), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19291), .ZN(n19794) );
  INV_X1 U17193 ( .A(n19794), .ZN(n19731) );
  AOI22_X1 U17194 ( .A1(n19745), .A2(n19791), .B1(n19710), .B2(n19731), .ZN(
        n13737) );
  OAI21_X1 U17195 ( .B1(n19788), .B2(n19707), .A(n13737), .ZN(n13738) );
  AOI21_X1 U17196 ( .B1(n13739), .B2(n19732), .A(n13738), .ZN(n13740) );
  OAI21_X1 U17197 ( .B1(n19686), .B2(n13741), .A(n13740), .ZN(P2_U3153) );
  AND2_X1 U17198 ( .A1(n13691), .A2(n13742), .ZN(n13744) );
  OR2_X1 U17199 ( .A1(n13744), .A2(n13743), .ZN(n20030) );
  INV_X1 U17200 ( .A(n13827), .ZN(n13745) );
  AOI21_X1 U17201 ( .B1(n13747), .B2(n13746), .A(n13745), .ZN(n20024) );
  AOI22_X1 U17202 ( .A1(n20024), .A2(n11194), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n14769), .ZN(n13748) );
  OAI21_X1 U17203 ( .B1(n20030), .B2(n14779), .A(n13748), .ZN(P1_U2863) );
  NOR2_X1 U17204 ( .A1(n19987), .A2(n19958), .ZN(n16382) );
  INV_X1 U17205 ( .A(n13749), .ZN(n13751) );
  INV_X1 U17206 ( .A(n12265), .ZN(n13750) );
  NAND2_X1 U17207 ( .A1(n13751), .A2(n13750), .ZN(n13757) );
  NAND2_X1 U17208 ( .A1(n13753), .A2(n13752), .ZN(n13754) );
  NOR2_X1 U17209 ( .A1(n13755), .A2(n13754), .ZN(n13756) );
  OAI22_X1 U17210 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19645), .B1(n16374), 
        .B2(n19845), .ZN(n13758) );
  AOI21_X1 U17211 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16382), .A(n13758), .ZN(
        n15860) );
  INV_X1 U17212 ( .A(n15840), .ZN(n15858) );
  NAND2_X1 U17213 ( .A1(n11496), .A2(n15858), .ZN(n13766) );
  INV_X1 U17214 ( .A(n12507), .ZN(n13760) );
  NAND2_X1 U17215 ( .A1(n13760), .A2(n13759), .ZN(n15821) );
  XNOR2_X1 U17216 ( .A(n13761), .B(n15832), .ZN(n13764) );
  AOI22_X1 U17217 ( .A1(n15821), .A2(n13764), .B1(n13763), .B2(n15848), .ZN(
        n13765) );
  NAND2_X1 U17218 ( .A1(n13766), .A2(n13765), .ZN(n16343) );
  INV_X1 U17219 ( .A(n16388), .ZN(n13772) );
  OAI21_X1 U17220 ( .B1(n19146), .B2(n13768), .A(n13767), .ZN(n13816) );
  OAI21_X1 U17221 ( .B1(n12794), .B2(n13769), .A(n13816), .ZN(n15843) );
  INV_X1 U17222 ( .A(n15843), .ZN(n13771) );
  INV_X1 U17223 ( .A(n19146), .ZN(n13770) );
  AOI22_X1 U17224 ( .A1(n19105), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n13770), .B2(n12794), .ZN(n15824) );
  NOR2_X1 U17225 ( .A1(n15824), .A2(n11444), .ZN(n15842) );
  AOI222_X1 U17226 ( .A1(n16343), .A2(n18952), .B1(n13772), .B2(n19952), .C1(
        n13771), .C2(n15842), .ZN(n13774) );
  NAND2_X1 U17227 ( .A1(n15860), .A2(n15832), .ZN(n13773) );
  OAI21_X1 U17228 ( .B1(n15860), .B2(n13774), .A(n13773), .ZN(P2_U3600) );
  XNOR2_X1 U17229 ( .A(n9642), .B(n13775), .ZN(n16304) );
  AND2_X1 U17230 ( .A1(n13778), .A2(n13777), .ZN(n13779) );
  OAI22_X1 U17231 ( .A1(n13782), .A2(n13781), .B1(n13780), .B2(n13779), .ZN(
        n16302) );
  INV_X1 U17232 ( .A(n16302), .ZN(n13795) );
  OAI21_X1 U17233 ( .B1(n13785), .B2(n13784), .A(n13783), .ZN(n19173) );
  OAI22_X1 U17234 ( .A1(n19173), .A2(n15816), .B1(n15811), .B2(n13786), .ZN(
        n13794) );
  NOR2_X1 U17235 ( .A1(n11864), .A2(n19113), .ZN(n13791) );
  AOI211_X1 U17236 ( .C1(n13789), .C2(n13788), .A(n13956), .B(n13787), .ZN(
        n13790) );
  AOI211_X1 U17237 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n13931), .A(
        n13791), .B(n13790), .ZN(n13792) );
  INV_X1 U17238 ( .A(n13792), .ZN(n13793) );
  AOI211_X1 U17239 ( .C1(n13795), .C2(n16328), .A(n13794), .B(n13793), .ZN(
        n13796) );
  OAI21_X1 U17240 ( .B1(n16320), .B2(n16304), .A(n13796), .ZN(P2_U3041) );
  XNOR2_X1 U17241 ( .A(n13797), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13798) );
  XNOR2_X1 U17242 ( .A(n13799), .B(n13798), .ZN(n16147) );
  INV_X1 U17243 ( .A(n16147), .ZN(n13805) );
  AOI22_X1 U17244 ( .A1(n20168), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20167), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13800) );
  OAI21_X1 U17245 ( .B1(n20178), .B2(n13801), .A(n13800), .ZN(n13802) );
  AOI21_X1 U17246 ( .B1(n13803), .B2(n20239), .A(n13802), .ZN(n13804) );
  OAI21_X1 U17247 ( .B1(n13805), .B2(n20007), .A(n13804), .ZN(P1_U2991) );
  INV_X1 U17248 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n13806) );
  INV_X1 U17249 ( .A(DATAI_9_), .ZN(n21017) );
  MUX2_X1 U17250 ( .A(n21017), .B(n16486), .S(n20238), .Z(n20132) );
  OAI222_X1 U17251 ( .A1(n20030), .A2(n14848), .B1(n13806), .B2(n14853), .C1(
        n14852), .C2(n20132), .ZN(P1_U2895) );
  NOR2_X1 U17252 ( .A1(n19101), .A2(n13807), .ZN(n13812) );
  AOI22_X1 U17253 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(n19135), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19142), .ZN(n13810) );
  NAND2_X1 U17254 ( .A1(n19141), .A2(n13808), .ZN(n13809) );
  OAI211_X1 U17255 ( .C1(n19133), .C2(n11445), .A(n13810), .B(n13809), .ZN(
        n13811) );
  AOI211_X1 U17256 ( .C1(n19954), .C2(n19129), .A(n13812), .B(n13811), .ZN(
        n13813) );
  OAI21_X1 U17257 ( .B1(n11502), .B2(n19137), .A(n13813), .ZN(n13814) );
  AOI21_X1 U17258 ( .B1(n19952), .B2(n19140), .A(n13814), .ZN(n13815) );
  OAI21_X1 U17259 ( .B1(n13816), .B2(n19851), .A(n13815), .ZN(P2_U2854) );
  INV_X1 U17260 ( .A(n13817), .ZN(n13820) );
  INV_X1 U17261 ( .A(n13845), .ZN(n13818) );
  OAI211_X1 U17262 ( .C1(n13820), .C2(n13819), .A(n13818), .B(n15298), .ZN(
        n13823) );
  INV_X1 U17263 ( .A(n15730), .ZN(n13821) );
  NAND2_X1 U17264 ( .A1(n13821), .A2(n15305), .ZN(n13822) );
  OAI211_X1 U17265 ( .C1(n15302), .C2(n13824), .A(n13823), .B(n13822), .ZN(
        P2_U2872) );
  XOR2_X1 U17266 ( .A(n13825), .B(n13743), .Z(n14061) );
  INV_X1 U17267 ( .A(n14061), .ZN(n14725) );
  AND2_X1 U17268 ( .A1(n13827), .A2(n13826), .ZN(n13828) );
  NOR2_X1 U17269 ( .A1(n9749), .A2(n13828), .ZN(n16129) );
  AOI22_X1 U17270 ( .A1(n16129), .A2(n11194), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14769), .ZN(n13829) );
  OAI21_X1 U17271 ( .B1(n14725), .B2(n14779), .A(n13829), .ZN(P1_U2862) );
  AOI22_X1 U17272 ( .A1(n11288), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13836) );
  OAI22_X1 U17273 ( .A1(n14290), .A2(n13831), .B1(n14289), .B2(n13830), .ZN(
        n13832) );
  INV_X1 U17274 ( .A(n13832), .ZN(n13835) );
  AOI22_X1 U17275 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14293), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13834) );
  AOI22_X1 U17276 ( .A1(n11531), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13833) );
  NAND4_X1 U17277 ( .A1(n13836), .A2(n13835), .A3(n13834), .A4(n13833), .ZN(
        n13844) );
  AOI22_X1 U17278 ( .A1(n14300), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13842) );
  AOI22_X1 U17279 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14301), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13841) );
  INV_X1 U17280 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13837) );
  OAI22_X1 U17281 ( .A1(n14305), .A2(n13837), .B1(n14303), .B2(n19256), .ZN(
        n13838) );
  INV_X1 U17282 ( .A(n13838), .ZN(n13840) );
  AOI22_X1 U17283 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14307), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13839) );
  NAND4_X1 U17284 ( .A1(n13842), .A2(n13841), .A3(n13840), .A4(n13839), .ZN(
        n13843) );
  OR2_X1 U17285 ( .A1(n13844), .A2(n13843), .ZN(n13846) );
  NOR2_X1 U17286 ( .A1(n13845), .A2(n13846), .ZN(n13847) );
  OR2_X1 U17287 ( .A1(n15287), .A2(n13847), .ZN(n13865) );
  AND2_X1 U17288 ( .A1(n13849), .A2(n13848), .ZN(n13850) );
  OR2_X1 U17289 ( .A1(n13850), .A2(n13893), .ZN(n19030) );
  NOR2_X1 U17290 ( .A1(n19030), .A2(n15309), .ZN(n13851) );
  AOI21_X1 U17291 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n15309), .A(n13851), .ZN(
        n13852) );
  OAI21_X1 U17292 ( .B1(n13865), .B2(n15312), .A(n13852), .ZN(P2_U2871) );
  NOR2_X2 U17293 ( .A1(n13855), .A2(n13853), .ZN(n19147) );
  NAND2_X1 U17294 ( .A1(n19149), .A2(BUF1_REG_16__SCAN_IN), .ZN(n13858) );
  NAND2_X1 U17295 ( .A1(n16235), .A2(n13856), .ZN(n13857) );
  OAI211_X1 U17296 ( .C1(n15380), .C2(n13859), .A(n13858), .B(n13857), .ZN(
        n13863) );
  INV_X1 U17297 ( .A(n13897), .ZN(n13860) );
  AOI21_X1 U17298 ( .B1(n13861), .B2(n12858), .A(n13860), .ZN(n15725) );
  INV_X1 U17299 ( .A(n15725), .ZN(n19031) );
  NOR2_X1 U17300 ( .A1(n19031), .A2(n16237), .ZN(n13862) );
  AOI211_X1 U17301 ( .C1(n19147), .C2(BUF2_REG_16__SCAN_IN), .A(n13863), .B(
        n13862), .ZN(n13864) );
  OAI21_X1 U17302 ( .B1(n19183), .B2(n13865), .A(n13864), .ZN(P2_U2903) );
  INV_X1 U17303 ( .A(DATAI_10_), .ZN(n21087) );
  MUX2_X1 U17304 ( .A(n21087), .B(n16484), .S(n20238), .Z(n20136) );
  INV_X1 U17305 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13866) );
  OAI222_X1 U17306 ( .A1(n14852), .A2(n20136), .B1(n14848), .B2(n14725), .C1(
        n13866), .C2(n14853), .ZN(P1_U2894) );
  XNOR2_X1 U17307 ( .A(n9672), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13867) );
  XNOR2_X1 U17308 ( .A(n13868), .B(n13867), .ZN(n16136) );
  INV_X1 U17309 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n13869) );
  NOR2_X1 U17310 ( .A1(n20225), .A2(n13869), .ZN(n16134) );
  AOI21_X1 U17311 ( .B1(n20168), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16134), .ZN(n13872) );
  INV_X1 U17312 ( .A(n20178), .ZN(n16044) );
  NAND2_X1 U17313 ( .A1(n16044), .A2(n13870), .ZN(n13871) );
  OAI211_X1 U17314 ( .C1(n20030), .C2(n16049), .A(n13872), .B(n13871), .ZN(
        n13873) );
  AOI21_X1 U17315 ( .B1(n16136), .B2(n20174), .A(n13873), .ZN(n13874) );
  INV_X1 U17316 ( .A(n13874), .ZN(P1_U2990) );
  AOI22_X1 U17317 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n14287), .B1(
        n11288), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13881) );
  INV_X1 U17318 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13876) );
  OAI22_X1 U17319 ( .A1(n13876), .A2(n14290), .B1(n14289), .B2(n13875), .ZN(
        n13877) );
  INV_X1 U17320 ( .A(n13877), .ZN(n13880) );
  AOI22_X1 U17321 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14293), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13879) );
  AOI22_X1 U17322 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11531), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13878) );
  NAND4_X1 U17323 ( .A1(n13881), .A2(n13880), .A3(n13879), .A4(n13878), .ZN(
        n13889) );
  AOI22_X1 U17324 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n14300), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13887) );
  AOI22_X1 U17325 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14301), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13886) );
  INV_X1 U17326 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13882) );
  OAI22_X1 U17327 ( .A1(n14305), .A2(n13882), .B1(n14303), .B2(n19259), .ZN(
        n13883) );
  INV_X1 U17328 ( .A(n13883), .ZN(n13885) );
  AOI22_X1 U17329 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n14307), .ZN(n13884) );
  NAND4_X1 U17330 ( .A1(n13887), .A2(n13886), .A3(n13885), .A4(n13884), .ZN(
        n13888) );
  OR2_X1 U17331 ( .A1(n13889), .A2(n13888), .ZN(n13985) );
  NAND2_X1 U17332 ( .A1(n15287), .A2(n13985), .ZN(n13921) );
  OR2_X1 U17333 ( .A1(n15287), .A2(n13985), .ZN(n13890) );
  NAND2_X1 U17334 ( .A1(n13921), .A2(n13890), .ZN(n13905) );
  OR2_X1 U17335 ( .A1(n13893), .A2(n13892), .ZN(n13894) );
  NAND2_X1 U17336 ( .A1(n13891), .A2(n13894), .ZN(n19015) );
  NOR2_X1 U17337 ( .A1(n19015), .A2(n15309), .ZN(n13895) );
  AOI21_X1 U17338 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n15309), .A(n13895), .ZN(
        n13896) );
  OAI21_X1 U17339 ( .B1(n13905), .B2(n15312), .A(n13896), .ZN(P2_U2870) );
  AOI21_X1 U17340 ( .B1(n13898), .B2(n13897), .A(n15220), .ZN(n19011) );
  INV_X1 U17341 ( .A(n19147), .ZN(n15384) );
  INV_X1 U17342 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n13902) );
  OAI22_X1 U17343 ( .A1(n19187), .A2(n15381), .B1(n15380), .B2(n13899), .ZN(
        n13900) );
  AOI21_X1 U17344 ( .B1(n19149), .B2(BUF1_REG_17__SCAN_IN), .A(n13900), .ZN(
        n13901) );
  OAI21_X1 U17345 ( .B1(n15384), .B2(n13902), .A(n13901), .ZN(n13903) );
  AOI21_X1 U17346 ( .B1(n19011), .B2(n19189), .A(n13903), .ZN(n13904) );
  OAI21_X1 U17347 ( .B1(n19183), .B2(n13905), .A(n13904), .ZN(P2_U2902) );
  AOI22_X1 U17348 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n14287), .B1(
        n11288), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13912) );
  INV_X1 U17349 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13906) );
  OAI22_X1 U17350 ( .A1(n13907), .A2(n14290), .B1(n14289), .B2(n13906), .ZN(
        n13908) );
  INV_X1 U17351 ( .A(n13908), .ZN(n13911) );
  AOI22_X1 U17352 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14293), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13910) );
  AOI22_X1 U17353 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n11531), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13909) );
  NAND4_X1 U17354 ( .A1(n13912), .A2(n13911), .A3(n13910), .A4(n13909), .ZN(
        n13920) );
  AOI22_X1 U17355 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n14300), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13918) );
  AOI22_X1 U17356 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14301), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13917) );
  OAI22_X1 U17357 ( .A1(n14305), .A2(n13913), .B1(n14303), .B2(n19264), .ZN(
        n13914) );
  INV_X1 U17358 ( .A(n13914), .ZN(n13916) );
  AOI22_X1 U17359 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__2__SCAN_IN), .B2(n14307), .ZN(n13915) );
  NAND4_X1 U17360 ( .A1(n13918), .A2(n13917), .A3(n13916), .A4(n13915), .ZN(
        n13919) );
  NOR2_X1 U17361 ( .A1(n13920), .A2(n13919), .ZN(n13984) );
  NAND2_X1 U17362 ( .A1(n13921), .A2(n13984), .ZN(n13922) );
  NAND2_X1 U17363 ( .A1(n13988), .A2(n13922), .ZN(n16236) );
  NAND2_X1 U17364 ( .A1(n15269), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n13926) );
  NAND2_X1 U17365 ( .A1(n13891), .A2(n13923), .ZN(n13924) );
  NAND2_X1 U17366 ( .A1(n9694), .A2(n13924), .ZN(n15693) );
  INV_X1 U17367 ( .A(n15693), .ZN(n15225) );
  NAND2_X1 U17368 ( .A1(n15225), .A2(n15302), .ZN(n13925) );
  OAI211_X1 U17369 ( .C1(n16236), .C2(n15312), .A(n13926), .B(n13925), .ZN(
        P2_U2869) );
  XOR2_X1 U17370 ( .A(n13928), .B(n13927), .Z(n16298) );
  INV_X1 U17371 ( .A(n16298), .ZN(n13943) );
  AND2_X1 U17372 ( .A1(n15798), .A2(n13929), .ZN(n13930) );
  NOR2_X1 U17373 ( .A1(n13931), .A2(n13930), .ZN(n16337) );
  INV_X1 U17374 ( .A(n16337), .ZN(n13941) );
  AND2_X1 U17375 ( .A1(n13957), .A2(n13956), .ZN(n13933) );
  NAND2_X1 U17376 ( .A1(n13933), .A2(n13932), .ZN(n13936) );
  NOR2_X1 U17377 ( .A1(n11869), .A2(n19113), .ZN(n13934) );
  AOI21_X1 U17378 ( .B1(n16331), .B2(n19108), .A(n13934), .ZN(n13935) );
  OAI211_X1 U17379 ( .C1(n15816), .C2(n19112), .A(n13936), .B(n13935), .ZN(
        n13940) );
  OAI21_X1 U17380 ( .B1(n13938), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13937), .ZN(n16295) );
  NOR2_X1 U17381 ( .A1(n16295), .A2(n15804), .ZN(n13939) );
  AOI211_X1 U17382 ( .C1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n13941), .A(
        n13940), .B(n13939), .ZN(n13942) );
  OAI21_X1 U17383 ( .B1(n16320), .B2(n13943), .A(n13942), .ZN(P2_U3040) );
  NOR2_X1 U17384 ( .A1(n9710), .A2(n13944), .ZN(n16279) );
  INV_X1 U17385 ( .A(n16279), .ZN(n13946) );
  OAI21_X1 U17386 ( .B1(n16278), .B2(n13944), .A(n9710), .ZN(n13945) );
  OAI21_X1 U17387 ( .B1(n13946), .B2(n16278), .A(n13945), .ZN(n13966) );
  NOR2_X1 U17388 ( .A1(n13955), .A2(n13736), .ZN(n13949) );
  OAI22_X1 U17389 ( .A1(n16310), .A2(n13947), .B1(n19879), .B2(n19113), .ZN(
        n13948) );
  AOI211_X1 U17390 ( .C1(n16301), .C2(n13950), .A(n13949), .B(n13948), .ZN(
        n13954) );
  XNOR2_X1 U17391 ( .A(n16288), .B(n16287), .ZN(n13952) );
  NOR2_X1 U17392 ( .A1(n13952), .A2(n16323), .ZN(n16286) );
  INV_X1 U17393 ( .A(n16286), .ZN(n13963) );
  NAND2_X1 U17394 ( .A1(n13952), .A2(n16323), .ZN(n13962) );
  NAND3_X1 U17395 ( .A1(n13963), .A2(n19236), .A3(n13962), .ZN(n13953) );
  OAI211_X1 U17396 ( .C1(n13966), .C2(n11993), .A(n13954), .B(n13953), .ZN(
        P2_U3007) );
  NOR2_X1 U17397 ( .A1(n15811), .A2(n13955), .ZN(n13960) );
  NAND3_X1 U17398 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13957), .A3(
        n13956), .ZN(n16322) );
  NAND2_X1 U17399 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n15544), .ZN(n13958) );
  OAI221_X1 U17400 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16322), .C1(
        n16323), .C2(n16337), .A(n13958), .ZN(n13959) );
  AOI211_X1 U17401 ( .C1(n16324), .C2(n13961), .A(n13960), .B(n13959), .ZN(
        n13965) );
  NAND3_X1 U17402 ( .A1(n13963), .A2(n16328), .A3(n13962), .ZN(n13964) );
  OAI211_X1 U17403 ( .C1(n13966), .C2(n16320), .A(n13965), .B(n13964), .ZN(
        P2_U3039) );
  OAI21_X1 U17404 ( .B1(n9682), .B2(n13967), .A(n9743), .ZN(n16030) );
  INV_X1 U17405 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n13968) );
  INV_X1 U17406 ( .A(DATAI_11_), .ZN(n21047) );
  MUX2_X1 U17407 ( .A(n21047), .B(n16482), .S(n20238), .Z(n20139) );
  OAI222_X1 U17408 ( .A1(n16030), .A2(n14848), .B1(n13968), .B2(n14853), .C1(
        n14852), .C2(n20139), .ZN(P1_U2893) );
  AOI22_X1 U17409 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n14287), .B1(
        n11288), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13975) );
  INV_X1 U17410 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13970) );
  OAI22_X1 U17411 ( .A1(n13970), .A2(n14290), .B1(n14289), .B2(n13969), .ZN(
        n13971) );
  INV_X1 U17412 ( .A(n13971), .ZN(n13974) );
  AOI22_X1 U17413 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14293), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13973) );
  AOI22_X1 U17414 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n11531), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13972) );
  NAND4_X1 U17415 ( .A1(n13975), .A2(n13974), .A3(n13973), .A4(n13972), .ZN(
        n13983) );
  AOI22_X1 U17416 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n14300), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13981) );
  AOI22_X1 U17417 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14301), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13980) );
  OAI22_X1 U17418 ( .A1(n14305), .A2(n13976), .B1(n14303), .B2(n19269), .ZN(
        n13977) );
  INV_X1 U17419 ( .A(n13977), .ZN(n13979) );
  AOI22_X1 U17420 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__3__SCAN_IN), .B2(n14245), .ZN(n13978) );
  NAND4_X1 U17421 ( .A1(n13981), .A2(n13980), .A3(n13979), .A4(n13978), .ZN(
        n13982) );
  NOR2_X1 U17422 ( .A1(n13983), .A2(n13982), .ZN(n13987) );
  NOR2_X1 U17423 ( .A1(n13987), .A2(n13984), .ZN(n13986) );
  AND2_X1 U17424 ( .A1(n13986), .A2(n13985), .ZN(n14252) );
  NAND2_X1 U17425 ( .A1(n15287), .A2(n14252), .ZN(n15295) );
  NAND2_X1 U17426 ( .A1(n13988), .A2(n13987), .ZN(n13989) );
  NAND2_X1 U17427 ( .A1(n15295), .A2(n13989), .ZN(n15313) );
  OR2_X1 U17428 ( .A1(n13990), .A2(n13991), .ZN(n13992) );
  NAND2_X1 U17429 ( .A1(n15665), .A2(n13992), .ZN(n19010) );
  INV_X1 U17430 ( .A(n19010), .ZN(n13998) );
  INV_X1 U17431 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n13996) );
  OAI22_X1 U17432 ( .A1(n19266), .A2(n15381), .B1(n15380), .B2(n13993), .ZN(
        n13994) );
  AOI21_X1 U17433 ( .B1(n19149), .B2(BUF1_REG_19__SCAN_IN), .A(n13994), .ZN(
        n13995) );
  OAI21_X1 U17434 ( .B1(n15384), .B2(n13996), .A(n13995), .ZN(n13997) );
  AOI21_X1 U17435 ( .B1(n13998), .B2(n19189), .A(n13997), .ZN(n13999) );
  OAI21_X1 U17436 ( .B1(n19183), .B2(n15313), .A(n13999), .ZN(P2_U2900) );
  NOR2_X1 U17437 ( .A1(n9749), .A2(n14000), .ZN(n14001) );
  OR2_X1 U17438 ( .A1(n14007), .A2(n14001), .ZN(n16118) );
  INV_X1 U17439 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n16023) );
  OAI222_X1 U17440 ( .A1(n16118), .A2(n14777), .B1(n16023), .B2(n14778), .C1(
        n16030), .C2(n14779), .ZN(P1_U2861) );
  OR2_X1 U17441 ( .A1(n14004), .A2(n14003), .ZN(n14005) );
  NAND2_X1 U17442 ( .A1(n14002), .A2(n14005), .ZN(n16050) );
  XOR2_X1 U17443 ( .A(n14007), .B(n14006), .Z(n16014) );
  AOI22_X1 U17444 ( .A1(n16014), .A2(n11194), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n14769), .ZN(n14008) );
  OAI21_X1 U17445 ( .B1(n16050), .B2(n14779), .A(n14008), .ZN(P1_U2860) );
  INV_X1 U17446 ( .A(n14009), .ZN(n14969) );
  AND2_X1 U17447 ( .A1(n14969), .A2(n14010), .ZN(n14993) );
  INV_X1 U17448 ( .A(n14011), .ZN(n14012) );
  NOR2_X1 U17449 ( .A1(n14993), .A2(n14012), .ZN(n14015) );
  NAND2_X1 U17450 ( .A1(n14013), .A2(n14992), .ZN(n14014) );
  XNOR2_X1 U17451 ( .A(n14015), .B(n14014), .ZN(n16054) );
  AOI22_X1 U17452 ( .A1(n16014), .A2(n20228), .B1(n20167), .B2(
        P1_REIP_REG_12__SCAN_IN), .ZN(n14028) );
  NAND3_X1 U17453 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16130) );
  NOR3_X1 U17454 ( .A1(n16133), .A2(n16139), .A3(n16130), .ZN(n16117) );
  INV_X1 U17455 ( .A(n16117), .ZN(n14020) );
  NOR2_X1 U17456 ( .A1(n16116), .A2(n14020), .ZN(n14035) );
  INV_X1 U17457 ( .A(n14035), .ZN(n14016) );
  NAND2_X1 U17458 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20185) );
  NOR2_X1 U17459 ( .A1(n16169), .A2(n20185), .ZN(n14019) );
  AOI21_X1 U17460 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20208) );
  INV_X1 U17461 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20233) );
  NAND2_X1 U17462 ( .A1(n15169), .A2(n15100), .ZN(n20219) );
  NAND2_X1 U17463 ( .A1(n16142), .A2(n20219), .ZN(n14017) );
  NOR2_X1 U17464 ( .A1(n20233), .A2(n14017), .ZN(n20205) );
  NAND2_X1 U17465 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n20205), .ZN(
        n16144) );
  NAND2_X1 U17466 ( .A1(n14019), .A2(n20193), .ZN(n16164) );
  NOR2_X1 U17467 ( .A1(n14016), .A2(n16164), .ZN(n14025) );
  INV_X1 U17468 ( .A(n14017), .ZN(n14046) );
  INV_X1 U17469 ( .A(n14019), .ZN(n14018) );
  NOR2_X1 U17470 ( .A1(n20208), .A2(n14018), .ZN(n16126) );
  AND2_X1 U17471 ( .A1(n14035), .A2(n16126), .ZN(n14022) );
  NAND3_X1 U17472 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n14019), .ZN(n14037) );
  AOI221_X1 U17473 ( .B1(n14037), .B2(n16142), .C1(n14020), .C2(n16142), .A(
        n20214), .ZN(n14021) );
  OAI21_X1 U17474 ( .B1(n14022), .B2(n20210), .A(n14021), .ZN(n16120) );
  AOI21_X1 U17475 ( .B1(n14046), .B2(n16116), .A(n16120), .ZN(n14023) );
  INV_X1 U17476 ( .A(n14023), .ZN(n14024) );
  MUX2_X1 U17477 ( .A(n14025), .B(n14024), .S(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n14026) );
  INV_X1 U17478 ( .A(n14026), .ZN(n14027) );
  OAI211_X1 U17479 ( .C1(n16054), .C2(n20222), .A(n14028), .B(n14027), .ZN(
        P1_U3019) );
  INV_X1 U17480 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14029) );
  INV_X1 U17481 ( .A(DATAI_12_), .ZN(n21062) );
  MUX2_X1 U17482 ( .A(n21062), .B(n16480), .S(n20238), .Z(n20142) );
  OAI222_X1 U17483 ( .A1(n16050), .A2(n14848), .B1(n14029), .B2(n14853), .C1(
        n14852), .C2(n20142), .ZN(P1_U2892) );
  OAI21_X1 U17484 ( .B1(n14691), .B2(n14030), .A(n14676), .ZN(n14767) );
  NOR2_X1 U17485 ( .A1(n9643), .A2(n14031), .ZN(n14984) );
  INV_X1 U17486 ( .A(n14032), .ZN(n14968) );
  OAI21_X1 U17487 ( .B1(n14984), .B2(n14968), .A(n14980), .ZN(n14034) );
  XNOR2_X1 U17488 ( .A(n14034), .B(n14033), .ZN(n16033) );
  NAND2_X1 U17489 ( .A1(n16033), .A2(n20206), .ZN(n14053) );
  NAND2_X1 U17490 ( .A1(n20220), .A2(n16114), .ZN(n14040) );
  NAND2_X1 U17491 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14035), .ZN(
        n16107) );
  INV_X1 U17492 ( .A(n16126), .ZN(n16127) );
  OR2_X1 U17493 ( .A1(n16107), .A2(n16127), .ZN(n15095) );
  NOR2_X1 U17494 ( .A1(n12230), .A2(n15095), .ZN(n14047) );
  INV_X1 U17495 ( .A(n14047), .ZN(n14036) );
  NAND2_X1 U17496 ( .A1(n20209), .A2(n14036), .ZN(n14039) );
  NOR2_X1 U17497 ( .A1(n14037), .A2(n16107), .ZN(n15145) );
  NAND2_X1 U17498 ( .A1(n15145), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14044) );
  AOI21_X1 U17499 ( .B1(n16142), .B2(n14044), .A(n20214), .ZN(n14038) );
  NAND2_X1 U17500 ( .A1(n14040), .A2(n16115), .ZN(n16100) );
  INV_X1 U17501 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14041) );
  NOR2_X1 U17502 ( .A1(n14042), .A2(n14041), .ZN(n16092) );
  AOI21_X1 U17503 ( .B1(n14042), .B2(n14041), .A(n16092), .ZN(n14043) );
  INV_X1 U17504 ( .A(n14043), .ZN(n14050) );
  INV_X1 U17505 ( .A(n14044), .ZN(n14045) );
  NAND2_X1 U17506 ( .A1(n14046), .A2(n14045), .ZN(n15078) );
  NAND2_X1 U17507 ( .A1(n20209), .A2(n14047), .ZN(n14048) );
  NAND2_X1 U17508 ( .A1(n15078), .A2(n14048), .ZN(n15016) );
  NAND2_X1 U17509 ( .A1(n15016), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16106) );
  INV_X1 U17510 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14049) );
  OAI22_X1 U17511 ( .A1(n14050), .A2(n16106), .B1(n20225), .B2(n14049), .ZN(
        n14051) );
  AOI21_X1 U17512 ( .B1(n16100), .B2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n14051), .ZN(n14052) );
  OAI211_X1 U17513 ( .C1(n20182), .C2(n14767), .A(n14053), .B(n14052), .ZN(
        P1_U3015) );
  NAND2_X1 U17514 ( .A1(n14056), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14055) );
  XNOR2_X1 U17515 ( .A(n9643), .B(n16133), .ZN(n14054) );
  MUX2_X1 U17516 ( .A(n14055), .B(n14054), .S(n9673), .Z(n14058) );
  NOR3_X1 U17517 ( .A1(n14056), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n14972), .ZN(n16055) );
  INV_X1 U17518 ( .A(n16055), .ZN(n14057) );
  NAND2_X1 U17519 ( .A1(n14058), .A2(n14057), .ZN(n16128) );
  INV_X1 U17520 ( .A(n16128), .ZN(n14063) );
  AOI22_X1 U17521 ( .A1(n20168), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20167), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14059) );
  OAI21_X1 U17522 ( .B1(n20178), .B2(n14718), .A(n14059), .ZN(n14060) );
  AOI21_X1 U17523 ( .B1(n14061), .B2(n20239), .A(n14060), .ZN(n14062) );
  OAI21_X1 U17524 ( .B1(n14063), .B2(n20007), .A(n14062), .ZN(P1_U2989) );
  NAND2_X1 U17525 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16940) );
  INV_X1 U17526 ( .A(n16940), .ZN(n14069) );
  INV_X1 U17527 ( .A(n15914), .ZN(n18752) );
  NOR4_X4 U17528 ( .A1(n18932), .A2(n14066), .A3(n15988), .A4(n18781), .ZN(
        n17285) );
  NOR2_X1 U17529 ( .A1(n18294), .A2(n14067), .ZN(n17281) );
  INV_X1 U17530 ( .A(n17281), .ZN(n17279) );
  INV_X1 U17531 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n16734) );
  INV_X1 U17532 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n16854) );
  INV_X1 U17533 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n16909) );
  INV_X1 U17534 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17284) );
  INV_X1 U17535 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17278) );
  NOR2_X1 U17536 ( .A1(n17284), .A2(n17278), .ZN(n17273) );
  INV_X1 U17537 ( .A(n17273), .ZN(n16925) );
  NOR2_X1 U17538 ( .A1(n16909), .A2(n16925), .ZN(n17261) );
  NAND3_X1 U17539 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17261), .ZN(n17263) );
  NAND2_X1 U17540 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17250), .ZN(n17177) );
  NAND4_X1 U17541 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(n14068), .ZN(n17178) );
  NOR3_X2 U17542 ( .A1(n16734), .A2(n16746), .A3(n17127), .ZN(n17095) );
  NAND2_X1 U17543 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17095), .ZN(n17094) );
  NAND3_X1 U17544 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .ZN(n16942) );
  NOR2_X2 U17545 ( .A1(n17004), .A2(n16942), .ZN(n17003) );
  NAND2_X1 U17546 ( .A1(n17274), .A2(n16985), .ZN(n16987) );
  OAI21_X1 U17547 ( .B1(n14069), .B2(n17279), .A(n16987), .ZN(n16979) );
  OAI22_X1 U17548 ( .A1(n17227), .A2(n17025), .B1(n17035), .B2(n14070), .ZN(
        n14080) );
  AOI22_X1 U17549 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14078) );
  AOI22_X1 U17550 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(n9652), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14077) );
  AOI22_X1 U17551 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14071) );
  OAI21_X1 U17552 ( .B1(n17163), .B2(n17022), .A(n14071), .ZN(n14075) );
  AOI22_X1 U17553 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14073) );
  AOI22_X1 U17554 ( .A1(n17225), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14072) );
  OAI211_X1 U17555 ( .C1(n17167), .C2(n15873), .A(n14073), .B(n14072), .ZN(
        n14074) );
  AOI211_X1 U17556 ( .C1(n12616), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n14075), .B(n14074), .ZN(n14076) );
  NAND3_X1 U17557 ( .A1(n14078), .A2(n14077), .A3(n14076), .ZN(n14079) );
  AOI211_X1 U17558 ( .C1(n17231), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n14080), .B(n14079), .ZN(n14144) );
  AOI22_X1 U17559 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14081) );
  OAI21_X1 U17560 ( .B1(n12100), .B2(n14082), .A(n14081), .ZN(n14092) );
  INV_X1 U17561 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17056) );
  AOI22_X1 U17562 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9630), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14090) );
  OAI22_X1 U17563 ( .A1(n9699), .A2(n18522), .B1(n17163), .B2(n14083), .ZN(
        n14088) );
  AOI22_X1 U17564 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14086) );
  AOI22_X1 U17565 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14085) );
  AOI22_X1 U17566 ( .A1(n12616), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17209), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14084) );
  NAND3_X1 U17567 ( .A1(n14086), .A2(n14085), .A3(n14084), .ZN(n14087) );
  AOI211_X1 U17568 ( .C1(n17101), .C2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A(
        n14088), .B(n14087), .ZN(n14089) );
  OAI211_X1 U17569 ( .C1(n17227), .C2(n17056), .A(n14090), .B(n14089), .ZN(
        n14091) );
  AOI211_X1 U17570 ( .C1(n17142), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n14092), .B(n14091), .ZN(n16983) );
  AOI22_X1 U17571 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17202), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14093) );
  OAI21_X1 U17572 ( .B1(n9699), .B2(n18516), .A(n14093), .ZN(n14102) );
  INV_X1 U17573 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17206) );
  AOI22_X1 U17574 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17231), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14100) );
  OAI22_X1 U17575 ( .A1(n17227), .A2(n17207), .B1(n18601), .B2(n17167), .ZN(
        n14098) );
  AOI22_X1 U17576 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17223), .ZN(n14096) );
  AOI22_X1 U17577 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n9633), .ZN(n14095) );
  AOI22_X1 U17578 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17209), .B1(
        n12616), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14094) );
  NAND3_X1 U17579 ( .A1(n14096), .A2(n14095), .A3(n14094), .ZN(n14097) );
  AOI211_X1 U17580 ( .C1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .C2(n17185), .A(
        n14098), .B(n14097), .ZN(n14099) );
  OAI211_X1 U17581 ( .C1(n17208), .C2(n17206), .A(n14100), .B(n14099), .ZN(
        n14101) );
  AOI211_X1 U17582 ( .C1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .C2(n17229), .A(
        n14102), .B(n14101), .ZN(n16995) );
  INV_X1 U17583 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18513) );
  AOI22_X1 U17584 ( .A1(n17204), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14112) );
  AOI22_X1 U17585 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15863), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14104) );
  AOI22_X1 U17586 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14103) );
  OAI211_X1 U17587 ( .C1(n17167), .C2(n18597), .A(n14104), .B(n14103), .ZN(
        n14110) );
  AOI22_X1 U17588 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14108) );
  AOI22_X1 U17589 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14107) );
  AOI22_X1 U17590 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14106) );
  NAND2_X1 U17591 ( .A1(n12616), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n14105) );
  NAND4_X1 U17592 ( .A1(n14108), .A2(n14107), .A3(n14106), .A4(n14105), .ZN(
        n14109) );
  AOI211_X1 U17593 ( .C1(n17209), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n14110), .B(n14109), .ZN(n14111) );
  OAI211_X1 U17594 ( .C1(n9699), .C2(n18513), .A(n14112), .B(n14111), .ZN(
        n17000) );
  AOI22_X1 U17595 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9630), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14122) );
  AOI22_X1 U17596 ( .A1(n17225), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14114) );
  AOI22_X1 U17597 ( .A1(n17229), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14113) );
  OAI211_X1 U17598 ( .C1(n17235), .C2(n16969), .A(n14114), .B(n14113), .ZN(
        n14120) );
  AOI22_X1 U17599 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14118) );
  AOI22_X1 U17600 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14117) );
  AOI22_X1 U17601 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n15863), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14116) );
  NAND2_X1 U17602 ( .A1(n17204), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14115) );
  NAND4_X1 U17603 ( .A1(n14118), .A2(n14117), .A3(n14116), .A4(n14115), .ZN(
        n14119) );
  AOI211_X1 U17604 ( .C1(n12616), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n14120), .B(n14119), .ZN(n14121) );
  OAI211_X1 U17605 ( .C1(n12608), .C2(n17113), .A(n14122), .B(n14121), .ZN(
        n17001) );
  NAND2_X1 U17606 ( .A1(n17000), .A2(n17001), .ZN(n16999) );
  NOR2_X1 U17607 ( .A1(n16995), .A2(n16999), .ZN(n16992) );
  AOI22_X1 U17608 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17209), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14132) );
  AOI22_X1 U17609 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15863), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14124) );
  AOI22_X1 U17610 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14123) );
  OAI211_X1 U17611 ( .C1(n17167), .C2(n18605), .A(n14124), .B(n14123), .ZN(
        n14130) );
  AOI22_X1 U17612 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17225), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14128) );
  AOI22_X1 U17613 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14127) );
  AOI22_X1 U17614 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14126) );
  NAND2_X1 U17615 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n14125) );
  NAND4_X1 U17616 ( .A1(n14128), .A2(n14127), .A3(n14126), .A4(n14125), .ZN(
        n14129) );
  AOI211_X1 U17617 ( .C1(n12616), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n14130), .B(n14129), .ZN(n14131) );
  OAI211_X1 U17618 ( .C1(n17227), .C2(n17071), .A(n14132), .B(n14131), .ZN(
        n16991) );
  NAND2_X1 U17619 ( .A1(n16992), .A2(n16991), .ZN(n16990) );
  NOR2_X1 U17620 ( .A1(n16983), .A2(n16990), .ZN(n17312) );
  AOI22_X1 U17621 ( .A1(n17225), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14143) );
  AOI22_X1 U17622 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14142) );
  AOI22_X1 U17623 ( .A1(n12616), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9630), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14141) );
  OAI22_X1 U17624 ( .A1(n17217), .A2(n17145), .B1(n17227), .B2(n14133), .ZN(
        n14139) );
  AOI22_X1 U17625 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n15863), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14137) );
  AOI22_X1 U17626 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14136) );
  AOI22_X1 U17627 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14135) );
  NAND2_X1 U17628 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n14134) );
  NAND4_X1 U17629 ( .A1(n14137), .A2(n14136), .A3(n14135), .A4(n14134), .ZN(
        n14138) );
  AOI211_X1 U17630 ( .C1(n17229), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n14139), .B(n14138), .ZN(n14140) );
  NAND4_X1 U17631 ( .A1(n14143), .A2(n14142), .A3(n14141), .A4(n14140), .ZN(
        n17311) );
  NAND2_X1 U17632 ( .A1(n17312), .A2(n17311), .ZN(n17310) );
  NOR2_X1 U17633 ( .A1(n14144), .A2(n17310), .ZN(n16976) );
  AOI21_X1 U17634 ( .B1(n14144), .B2(n17310), .A(n16976), .ZN(n17304) );
  AOI22_X1 U17635 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16979), .B1(n17282), 
        .B2(n17304), .ZN(n14148) );
  INV_X1 U17636 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14146) );
  INV_X1 U17637 ( .A(n16985), .ZN(n14145) );
  NAND3_X1 U17638 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14146), .A3(n14145), 
        .ZN(n14147) );
  NAND2_X1 U17639 ( .A1(n14148), .A2(n14147), .ZN(P3_U2675) );
  NAND2_X1 U17640 ( .A1(n14857), .A2(n14149), .ZN(n14151) );
  INV_X1 U17641 ( .A(n14159), .ZN(n14526) );
  INV_X1 U17642 ( .A(n14528), .ZN(n14156) );
  INV_X1 U17643 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21052) );
  NOR2_X1 U17644 ( .A1(n20225), .A2(n21052), .ZN(n15034) );
  AOI21_X1 U17645 ( .B1(n20168), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15034), .ZN(n14155) );
  OAI21_X1 U17646 ( .B1(n20178), .B2(n14156), .A(n14155), .ZN(n14157) );
  OAI21_X1 U17647 ( .B1(n20007), .B2(n15042), .A(n14158), .ZN(P1_U2970) );
  NOR3_X1 U17648 ( .A1(n14849), .A2(n14161), .A3(n14160), .ZN(n14820) );
  INV_X1 U17649 ( .A(DATAI_13_), .ZN(n21050) );
  MUX2_X1 U17650 ( .A(n21050), .B(n16478), .S(n20238), .Z(n20145) );
  OAI22_X1 U17651 ( .A1(n14840), .A2(n20145), .B1(n14853), .B2(n13237), .ZN(
        n14162) );
  AOI21_X1 U17652 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n14842), .A(n14162), .ZN(
        n14164) );
  NAND2_X1 U17653 ( .A1(n11080), .A2(DATAI_29_), .ZN(n14163) );
  OAI211_X1 U17654 ( .C1(n14159), .C2(n14848), .A(n14164), .B(n14163), .ZN(
        P1_U2875) );
  NOR2_X1 U17655 ( .A1(n14166), .A2(n14165), .ZN(n14167) );
  OAI222_X1 U17656 ( .A1(n14159), .A2(n14779), .B1(n14531), .B2(n14778), .C1(
        n14527), .C2(n14777), .ZN(P1_U2843) );
  AOI222_X1 U17657 ( .A1(n12314), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12503), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n14168), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14169) );
  NAND3_X1 U17658 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14207) );
  AND2_X1 U17659 ( .A1(n15798), .A2(n14207), .ZN(n14171) );
  NOR2_X1 U17660 ( .A1(n15583), .A2(n14171), .ZN(n14209) );
  OAI21_X1 U17661 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15710), .A(
        n14209), .ZN(n14173) );
  AOI21_X1 U17662 ( .B1(n14173), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n14172), .ZN(n14174) );
  INV_X1 U17663 ( .A(n14174), .ZN(n14175) );
  NAND2_X1 U17664 ( .A1(n14177), .A2(n16328), .ZN(n14178) );
  OAI211_X1 U17665 ( .C1(n14180), .C2(n16320), .A(n14179), .B(n14178), .ZN(
        P2_U3015) );
  NAND2_X1 U17666 ( .A1(n14182), .A2(n14181), .ZN(n14187) );
  INV_X1 U17667 ( .A(n14183), .ZN(n14184) );
  NOR2_X1 U17668 ( .A1(n14185), .A2(n14184), .ZN(n14186) );
  XNOR2_X1 U17669 ( .A(n14187), .B(n14186), .ZN(n14218) );
  XNOR2_X1 U17670 ( .A(n14188), .B(n14208), .ZN(n14215) );
  INV_X1 U17671 ( .A(n16187), .ZN(n14191) );
  NAND2_X1 U17672 ( .A1(n15544), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n14211) );
  OAI21_X1 U17673 ( .B1(n16310), .B2(n14189), .A(n14211), .ZN(n14190) );
  AOI21_X1 U17674 ( .B1(n16301), .B2(n14191), .A(n14190), .ZN(n14192) );
  OAI21_X1 U17675 ( .B1(n14457), .B2(n13736), .A(n14192), .ZN(n14193) );
  AOI21_X1 U17676 ( .B1(n14215), .B2(n19236), .A(n14193), .ZN(n14194) );
  OAI21_X1 U17677 ( .B1(n14218), .B2(n11993), .A(n14194), .ZN(P2_U2984) );
  INV_X1 U17678 ( .A(n12884), .ZN(n14199) );
  INV_X1 U17679 ( .A(n14197), .ZN(n14198) );
  NAND2_X1 U17680 ( .A1(n14199), .A2(n14198), .ZN(n14200) );
  NAND2_X1 U17681 ( .A1(n16301), .A2(n15195), .ZN(n14201) );
  NAND2_X1 U17682 ( .A1(n15544), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15565) );
  OAI211_X1 U17683 ( .C1(n16310), .C2(n14202), .A(n14201), .B(n15565), .ZN(
        n14205) );
  OAI21_X1 U17684 ( .B1(n15400), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14203), .ZN(n15562) );
  NOR2_X1 U17685 ( .A1(n15562), .A2(n16303), .ZN(n14204) );
  AOI211_X1 U17686 ( .C1(n16306), .C2(n15567), .A(n14205), .B(n14204), .ZN(
        n14206) );
  OAI21_X1 U17687 ( .B1(n15578), .B2(n11993), .A(n14206), .ZN(P2_U2986) );
  OR2_X1 U17688 ( .A1(n14209), .A2(n14208), .ZN(n14210) );
  OAI211_X1 U17689 ( .C1(n14457), .C2(n15811), .A(n14211), .B(n14210), .ZN(
        n14212) );
  INV_X1 U17690 ( .A(n14212), .ZN(n14213) );
  INV_X1 U17691 ( .A(n14214), .ZN(n14217) );
  NAND2_X1 U17692 ( .A1(n14215), .A2(n16328), .ZN(n14216) );
  OAI211_X1 U17693 ( .C1(n14218), .C2(n16320), .A(n14217), .B(n14216), .ZN(
        P2_U3016) );
  MUX2_X1 U17694 ( .A(n15841), .B(n14219), .S(n15269), .Z(n14220) );
  OAI21_X1 U17695 ( .B1(n19942), .B2(n15312), .A(n14220), .ZN(P2_U2885) );
  AOI22_X1 U17696 ( .A1(n11288), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14287), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14227) );
  INV_X1 U17697 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14222) );
  OAI22_X1 U17698 ( .A1(n14290), .A2(n14222), .B1(n14289), .B2(n14221), .ZN(
        n14223) );
  INV_X1 U17699 ( .A(n14223), .ZN(n14226) );
  AOI22_X1 U17700 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14293), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14225) );
  AOI22_X1 U17701 ( .A1(n11531), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14224) );
  NAND4_X1 U17702 ( .A1(n14227), .A2(n14226), .A3(n14225), .A4(n14224), .ZN(
        n14235) );
  AOI22_X1 U17703 ( .A1(n14300), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14233) );
  AOI22_X1 U17704 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14301), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14232) );
  INV_X1 U17705 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14228) );
  OAI22_X1 U17706 ( .A1(n14305), .A2(n14228), .B1(n14303), .B2(n13216), .ZN(
        n14229) );
  INV_X1 U17707 ( .A(n14229), .ZN(n14231) );
  AOI22_X1 U17708 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14307), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14230) );
  NAND4_X1 U17709 ( .A1(n14233), .A2(n14232), .A3(n14231), .A4(n14230), .ZN(
        n14234) );
  OR2_X1 U17710 ( .A1(n14235), .A2(n14234), .ZN(n15289) );
  AOI22_X1 U17711 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n14287), .B1(
        n11288), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14242) );
  INV_X1 U17712 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14236) );
  OAI22_X1 U17713 ( .A1(n14237), .A2(n14290), .B1(n14289), .B2(n14236), .ZN(
        n14238) );
  INV_X1 U17714 ( .A(n14238), .ZN(n14241) );
  AOI22_X1 U17715 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14293), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14240) );
  AOI22_X1 U17716 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11531), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14239) );
  NAND4_X1 U17717 ( .A1(n14242), .A2(n14241), .A3(n14240), .A4(n14239), .ZN(
        n14251) );
  AOI22_X1 U17718 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n14300), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14249) );
  AOI22_X1 U17719 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14301), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14248) );
  INV_X1 U17720 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14243) );
  INV_X1 U17721 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19273) );
  OAI22_X1 U17722 ( .A1(n14305), .A2(n14243), .B1(n14303), .B2(n19273), .ZN(
        n14244) );
  INV_X1 U17723 ( .A(n14244), .ZN(n14247) );
  AOI22_X1 U17724 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .B2(n14245), .ZN(n14246) );
  NAND4_X1 U17725 ( .A1(n14249), .A2(n14248), .A3(n14247), .A4(n14246), .ZN(
        n14250) );
  OR2_X1 U17726 ( .A1(n14251), .A2(n14250), .ZN(n15293) );
  AND2_X1 U17727 ( .A1(n15293), .A2(n14252), .ZN(n15286) );
  AND2_X1 U17728 ( .A1(n15289), .A2(n15286), .ZN(n15280) );
  AOI22_X1 U17729 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n14287), .B1(
        n11288), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14260) );
  INV_X1 U17730 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14253) );
  OAI22_X1 U17731 ( .A1(n14254), .A2(n14290), .B1(n14289), .B2(n14253), .ZN(
        n14255) );
  INV_X1 U17732 ( .A(n14255), .ZN(n14259) );
  AOI22_X1 U17733 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14293), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14258) );
  AOI22_X1 U17734 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n11531), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14257) );
  NAND4_X1 U17735 ( .A1(n14260), .A2(n14259), .A3(n14258), .A4(n14257), .ZN(
        n14268) );
  AOI22_X1 U17736 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n14300), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14266) );
  AOI22_X1 U17737 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14301), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14265) );
  INV_X1 U17738 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14261) );
  OAI22_X1 U17739 ( .A1(n14305), .A2(n14261), .B1(n14303), .B2(n19286), .ZN(
        n14262) );
  INV_X1 U17740 ( .A(n14262), .ZN(n14264) );
  AOI22_X1 U17741 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n14307), .ZN(n14263) );
  NAND4_X1 U17742 ( .A1(n14266), .A2(n14265), .A3(n14264), .A4(n14263), .ZN(
        n14267) );
  OR2_X1 U17743 ( .A1(n14268), .A2(n14267), .ZN(n15281) );
  AND2_X1 U17744 ( .A1(n15280), .A2(n15281), .ZN(n14269) );
  NAND2_X1 U17745 ( .A1(n14270), .A2(n14269), .ZN(n14317) );
  AOI22_X1 U17746 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9637), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14274) );
  AOI22_X1 U17747 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14273) );
  AND2_X1 U17748 ( .A1(n14274), .A2(n14273), .ZN(n14277) );
  AOI22_X1 U17749 ( .A1(n9648), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9651), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14276) );
  AOI22_X1 U17750 ( .A1(n11375), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9653), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14275) );
  XNOR2_X1 U17751 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14441) );
  NAND4_X1 U17752 ( .A1(n14277), .A2(n14276), .A3(n14275), .A4(n14441), .ZN(
        n14286) );
  AOI22_X1 U17753 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14399), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14284) );
  NAND2_X1 U17754 ( .A1(n11374), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n14281) );
  NAND2_X1 U17755 ( .A1(n11375), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n14280) );
  NAND2_X1 U17756 ( .A1(n14436), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n14279) );
  NAND2_X1 U17757 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n14278) );
  AND4_X1 U17758 ( .A1(n14281), .A2(n14280), .A3(n14279), .A4(n14278), .ZN(
        n14283) );
  INV_X1 U17759 ( .A(n14441), .ZN(n14433) );
  AOI22_X1 U17760 ( .A1(n9637), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14282) );
  NAND4_X1 U17761 ( .A1(n14284), .A2(n14283), .A3(n14433), .A4(n14282), .ZN(
        n14285) );
  NAND2_X1 U17762 ( .A1(n14286), .A2(n14285), .ZN(n14337) );
  NOR2_X1 U17763 ( .A1(n11551), .A2(n14337), .ZN(n14316) );
  AOI22_X1 U17764 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n14287), .B1(
        n11288), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14298) );
  INV_X1 U17765 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14291) );
  INV_X1 U17766 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14288) );
  OAI22_X1 U17767 ( .A1(n14291), .A2(n14290), .B1(n14289), .B2(n14288), .ZN(
        n14292) );
  INV_X1 U17768 ( .A(n14292), .ZN(n14297) );
  AOI22_X1 U17769 ( .A1(n14294), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14293), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14296) );
  AOI22_X1 U17770 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n11531), .B1(
        n11625), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14295) );
  NAND4_X1 U17771 ( .A1(n14298), .A2(n14297), .A3(n14296), .A4(n14295), .ZN(
        n14314) );
  AOI22_X1 U17772 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n14300), .B1(
        n14299), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14312) );
  AOI22_X1 U17773 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14301), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14311) );
  INV_X1 U17774 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14304) );
  OAI22_X1 U17775 ( .A1(n14305), .A2(n14304), .B1(n14303), .B2(n14302), .ZN(
        n14306) );
  INV_X1 U17776 ( .A(n14306), .ZN(n14310) );
  AOI22_X1 U17777 ( .A1(n14308), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n14307), .ZN(n14309) );
  NAND4_X1 U17778 ( .A1(n14312), .A2(n14311), .A3(n14310), .A4(n14309), .ZN(
        n14313) );
  OR2_X1 U17779 ( .A1(n14314), .A2(n14313), .ZN(n14333) );
  INV_X1 U17780 ( .A(n14333), .ZN(n14315) );
  XNOR2_X1 U17781 ( .A(n14316), .B(n14315), .ZN(n14335) );
  XNOR2_X1 U17782 ( .A(n14317), .B(n14335), .ZN(n15273) );
  INV_X1 U17783 ( .A(n14337), .ZN(n14332) );
  AND2_X1 U17784 ( .A1(n11551), .A2(n14332), .ZN(n15272) );
  INV_X1 U17785 ( .A(n14317), .ZN(n14318) );
  AOI22_X1 U17786 ( .A1(n9647), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(n9656), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14321) );
  AOI22_X1 U17787 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14320) );
  AND2_X1 U17788 ( .A1(n14321), .A2(n14320), .ZN(n14324) );
  AOI22_X1 U17789 ( .A1(n14417), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9651), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14323) );
  AOI22_X1 U17790 ( .A1(n11375), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n14436), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14322) );
  NAND4_X1 U17791 ( .A1(n14324), .A2(n14323), .A3(n14322), .A4(n14441), .ZN(
        n14331) );
  AOI22_X1 U17792 ( .A1(n9647), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9655), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14326) );
  AOI22_X1 U17793 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14325) );
  AND2_X1 U17794 ( .A1(n14326), .A2(n14325), .ZN(n14329) );
  AOI22_X1 U17795 ( .A1(n14417), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11374), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14328) );
  AOI22_X1 U17796 ( .A1(n11375), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14436), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14327) );
  NAND4_X1 U17797 ( .A1(n14329), .A2(n14433), .A3(n14328), .A4(n14327), .ZN(
        n14330) );
  AND2_X1 U17798 ( .A1(n14331), .A2(n14330), .ZN(n14336) );
  AND2_X1 U17799 ( .A1(n14333), .A2(n14332), .ZN(n14334) );
  NAND2_X1 U17800 ( .A1(n14334), .A2(n14336), .ZN(n14339) );
  OAI211_X1 U17801 ( .C1(n14336), .C2(n14334), .A(n14393), .B(n14339), .ZN(
        n15262) );
  INV_X1 U17802 ( .A(n14335), .ZN(n14338) );
  NAND2_X1 U17803 ( .A1(n11551), .A2(n14336), .ZN(n15265) );
  INV_X1 U17804 ( .A(n14339), .ZN(n14352) );
  AOI22_X1 U17805 ( .A1(n9647), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n9657), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14341) );
  AOI22_X1 U17806 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14340) );
  AND2_X1 U17807 ( .A1(n14341), .A2(n14340), .ZN(n14344) );
  AOI22_X1 U17808 ( .A1(n14417), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9651), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14343) );
  AOI22_X1 U17809 ( .A1(n11375), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9654), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14342) );
  NAND4_X1 U17810 ( .A1(n14344), .A2(n14343), .A3(n14342), .A4(n14441), .ZN(
        n14351) );
  AOI22_X1 U17811 ( .A1(n9647), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9637), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14346) );
  AOI22_X1 U17812 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14345) );
  AND2_X1 U17813 ( .A1(n14346), .A2(n14345), .ZN(n14349) );
  AOI22_X1 U17814 ( .A1(n14417), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9651), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14348) );
  AOI22_X1 U17815 ( .A1(n11375), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14436), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14347) );
  NAND4_X1 U17816 ( .A1(n14349), .A2(n14433), .A3(n14348), .A4(n14347), .ZN(
        n14350) );
  AND2_X1 U17817 ( .A1(n14351), .A2(n14350), .ZN(n14353) );
  NAND2_X1 U17818 ( .A1(n14352), .A2(n14353), .ZN(n14374) );
  OAI211_X1 U17819 ( .C1(n14352), .C2(n14353), .A(n14393), .B(n14374), .ZN(
        n14357) );
  INV_X1 U17820 ( .A(n14353), .ZN(n14354) );
  NOR2_X1 U17821 ( .A1(n14355), .A2(n14354), .ZN(n15258) );
  INV_X1 U17822 ( .A(n14356), .ZN(n14359) );
  NAND2_X2 U17823 ( .A1(n15257), .A2(n14360), .ZN(n14378) );
  AOI22_X1 U17824 ( .A1(n9647), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9655), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14362) );
  AOI22_X1 U17825 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14361) );
  AND2_X1 U17826 ( .A1(n14362), .A2(n14361), .ZN(n14365) );
  AOI22_X1 U17827 ( .A1(n14417), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9651), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14364) );
  AOI22_X1 U17828 ( .A1(n11375), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9653), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14363) );
  NAND4_X1 U17829 ( .A1(n14365), .A2(n14364), .A3(n14363), .A4(n14441), .ZN(
        n14372) );
  AOI22_X1 U17830 ( .A1(n9647), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9637), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14367) );
  AOI22_X1 U17831 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14366) );
  AND2_X1 U17832 ( .A1(n14367), .A2(n14366), .ZN(n14370) );
  AOI22_X1 U17833 ( .A1(n14417), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11374), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14369) );
  AOI22_X1 U17834 ( .A1(n11375), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9654), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14368) );
  NAND4_X1 U17835 ( .A1(n14370), .A2(n14433), .A3(n14369), .A4(n14368), .ZN(
        n14371) );
  NAND2_X1 U17836 ( .A1(n14372), .A2(n14371), .ZN(n14376) );
  INV_X1 U17837 ( .A(n14393), .ZN(n14373) );
  AOI21_X1 U17838 ( .B1(n14374), .B2(n14376), .A(n14373), .ZN(n14375) );
  OR2_X1 U17839 ( .A1(n14374), .A2(n14376), .ZN(n14380) );
  XNOR2_X2 U17840 ( .A(n14378), .B(n9757), .ZN(n15254) );
  INV_X1 U17841 ( .A(n14376), .ZN(n14377) );
  NAND2_X1 U17842 ( .A1(n11551), .A2(n14377), .ZN(n15253) );
  INV_X1 U17843 ( .A(n14380), .ZN(n14394) );
  AOI22_X1 U17844 ( .A1(n9647), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(n9657), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14382) );
  AOI22_X1 U17845 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14381) );
  AND2_X1 U17846 ( .A1(n14382), .A2(n14381), .ZN(n14385) );
  AOI22_X1 U17847 ( .A1(n14417), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9651), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14384) );
  AOI22_X1 U17848 ( .A1(n11375), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9654), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14383) );
  NAND4_X1 U17849 ( .A1(n14385), .A2(n14384), .A3(n14383), .A4(n14441), .ZN(
        n14392) );
  AOI22_X1 U17850 ( .A1(n9647), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14387) );
  AOI22_X1 U17851 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14386) );
  AND2_X1 U17852 ( .A1(n14387), .A2(n14386), .ZN(n14390) );
  AOI22_X1 U17853 ( .A1(n14417), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11374), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14389) );
  AOI22_X1 U17854 ( .A1(n11375), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9654), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14388) );
  NAND4_X1 U17855 ( .A1(n14390), .A2(n14433), .A3(n14389), .A4(n14388), .ZN(
        n14391) );
  AND2_X1 U17856 ( .A1(n14392), .A2(n14391), .ZN(n14396) );
  NAND2_X1 U17857 ( .A1(n14394), .A2(n14396), .ZN(n15240) );
  OAI211_X1 U17858 ( .C1(n14394), .C2(n14396), .A(n15240), .B(n14393), .ZN(
        n14395) );
  INV_X1 U17859 ( .A(n14396), .ZN(n14397) );
  NOR2_X1 U17860 ( .A1(n19989), .A2(n14397), .ZN(n15246) );
  NAND2_X1 U17861 ( .A1(n15247), .A2(n15246), .ZN(n15245) );
  AOI22_X1 U17862 ( .A1(n9647), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(n9637), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14401) );
  AOI22_X1 U17863 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14400) );
  AND2_X1 U17864 ( .A1(n14401), .A2(n14400), .ZN(n14404) );
  AOI22_X1 U17865 ( .A1(n14417), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11374), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14403) );
  AOI22_X1 U17866 ( .A1(n11375), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14436), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14402) );
  NAND4_X1 U17867 ( .A1(n14404), .A2(n14403), .A3(n14402), .A4(n14441), .ZN(
        n14411) );
  AOI22_X1 U17868 ( .A1(n9647), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9637), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14406) );
  AOI22_X1 U17869 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14405) );
  AND2_X1 U17870 ( .A1(n14406), .A2(n14405), .ZN(n14409) );
  AOI22_X1 U17871 ( .A1(n14417), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11374), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14408) );
  AOI22_X1 U17872 ( .A1(n11375), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9653), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14407) );
  NAND4_X1 U17873 ( .A1(n14409), .A2(n14433), .A3(n14408), .A4(n14407), .ZN(
        n14410) );
  NAND2_X1 U17874 ( .A1(n14411), .A2(n14410), .ZN(n14425) );
  AOI21_X2 U17875 ( .B1(n15245), .B2(n10126), .A(n14425), .ZN(n15236) );
  AOI22_X1 U17876 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n9655), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14413) );
  AOI22_X1 U17877 ( .A1(n9647), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14412) );
  AND2_X1 U17878 ( .A1(n14413), .A2(n14412), .ZN(n14416) );
  AOI22_X1 U17879 ( .A1(n14417), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11374), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14415) );
  AOI22_X1 U17880 ( .A1(n11375), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9654), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14414) );
  NAND4_X1 U17881 ( .A1(n14416), .A2(n14415), .A3(n14414), .A4(n14441), .ZN(
        n14424) );
  AOI22_X1 U17882 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9656), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14419) );
  AOI22_X1 U17883 ( .A1(n14417), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14418) );
  AND2_X1 U17884 ( .A1(n14419), .A2(n14418), .ZN(n14422) );
  AOI22_X1 U17885 ( .A1(n9647), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9651), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14421) );
  AOI22_X1 U17886 ( .A1(n11375), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14436), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14420) );
  NAND4_X1 U17887 ( .A1(n14422), .A2(n14433), .A3(n14421), .A4(n14420), .ZN(
        n14423) );
  NAND2_X1 U17888 ( .A1(n14424), .A2(n14423), .ZN(n14428) );
  INV_X1 U17889 ( .A(n14425), .ZN(n15241) );
  NAND2_X1 U17890 ( .A1(n19989), .A2(n15241), .ZN(n14426) );
  OR2_X1 U17891 ( .A1(n15240), .A2(n14426), .ZN(n14427) );
  NOR2_X1 U17892 ( .A1(n14427), .A2(n14428), .ZN(n14429) );
  AOI21_X1 U17893 ( .B1(n14428), .B2(n14427), .A(n14429), .ZN(n15235) );
  NAND2_X1 U17894 ( .A1(n15236), .A2(n15235), .ZN(n15237) );
  INV_X1 U17895 ( .A(n14429), .ZN(n14430) );
  AOI22_X1 U17896 ( .A1(n11375), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9654), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14432) );
  AOI22_X1 U17897 ( .A1(n9647), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11374), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14431) );
  NAND2_X1 U17898 ( .A1(n14432), .A2(n14431), .ZN(n14447) );
  AOI22_X1 U17899 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9661), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14435) );
  AOI22_X1 U17900 ( .A1(n9637), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14434) );
  NAND3_X1 U17901 ( .A1(n14435), .A2(n14434), .A3(n14433), .ZN(n14446) );
  AOI22_X1 U17902 ( .A1(n11375), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9653), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14439) );
  AOI22_X1 U17903 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9651), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14438) );
  NAND2_X1 U17904 ( .A1(n14439), .A2(n14438), .ZN(n14445) );
  AOI22_X1 U17905 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n9657), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14443) );
  AOI22_X1 U17906 ( .A1(n9647), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14272), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14442) );
  NAND3_X1 U17907 ( .A1(n14443), .A2(n14442), .A3(n14441), .ZN(n14444) );
  OAI22_X1 U17908 ( .A1(n14447), .A2(n14446), .B1(n14445), .B2(n14444), .ZN(
        n14448) );
  INV_X1 U17909 ( .A(n14448), .ZN(n14449) );
  INV_X1 U17910 ( .A(n19149), .ZN(n15346) );
  INV_X1 U17911 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n14783) );
  AOI22_X1 U17912 ( .A1(n16235), .A2(n19152), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n19188), .ZN(n14453) );
  NAND2_X1 U17913 ( .A1(n19147), .A2(BUF2_REG_30__SCAN_IN), .ZN(n14452) );
  OAI211_X1 U17914 ( .C1(n15346), .C2(n14783), .A(n14453), .B(n14452), .ZN(
        n14454) );
  AOI21_X1 U17915 ( .B1(n14455), .B2(n19189), .A(n14454), .ZN(n14456) );
  OAI21_X1 U17916 ( .B1(n14460), .B2(n19183), .A(n14456), .ZN(P2_U2889) );
  NOR2_X1 U17917 ( .A1(n14457), .A2(n15309), .ZN(n14458) );
  AOI21_X1 U17918 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n15269), .A(n14458), .ZN(
        n14459) );
  OAI21_X1 U17919 ( .B1(n14460), .B2(n15312), .A(n14459), .ZN(P2_U2857) );
  NAND2_X1 U17920 ( .A1(n16301), .A2(n13673), .ZN(n14463) );
  OAI211_X1 U17921 ( .C1(n16310), .C2(n14464), .A(n14463), .B(n14462), .ZN(
        n14468) );
  AND3_X1 U17922 ( .A1(n14466), .A2(n14465), .A3(n16297), .ZN(n14467) );
  AOI211_X1 U17923 ( .C1(n14469), .C2(n19236), .A(n14468), .B(n14467), .ZN(
        n14470) );
  OAI21_X1 U17924 ( .B1(n15841), .B2(n13736), .A(n14470), .ZN(P2_U3012) );
  NAND3_X1 U17925 ( .A1(n14472), .A2(n12980), .A3(n14471), .ZN(n14473) );
  MUX2_X1 U17926 ( .A(n14474), .B(n14473), .S(n14483), .Z(n14478) );
  INV_X1 U17927 ( .A(n11062), .ZN(n14476) );
  NOR2_X1 U17928 ( .A1(n14476), .A2(n14475), .ZN(n14477) );
  OR2_X1 U17929 ( .A1(n14478), .A2(n14477), .ZN(n15955) );
  INV_X1 U17930 ( .A(n12980), .ZN(n14479) );
  NOR2_X1 U17931 ( .A1(n14480), .A2(n14479), .ZN(n14481) );
  AOI21_X1 U17932 ( .B1(n14483), .B2(n14482), .A(n14481), .ZN(n20001) );
  OR2_X1 U17933 ( .A1(n14485), .A2(n14484), .ZN(n20912) );
  NAND2_X1 U17934 ( .A1(n20912), .A2(n20918), .ZN(n14486) );
  NAND2_X1 U17935 ( .A1(n20001), .A2(n14486), .ZN(n15953) );
  AND2_X1 U17936 ( .A1(n15953), .A2(n20000), .ZN(n20009) );
  MUX2_X1 U17937 ( .A(P1_MORE_REG_SCAN_IN), .B(n15955), .S(n20009), .Z(
        P1_U3484) );
  INV_X1 U17938 ( .A(n14487), .ZN(n14514) );
  MUX2_X1 U17939 ( .A(n14490), .B(n14489), .S(n14488), .Z(n14494) );
  AOI22_X1 U17940 ( .A1(n14492), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(n14491), .ZN(n14493) );
  XNOR2_X1 U17941 ( .A(n14494), .B(n14493), .ZN(n15022) );
  INV_X1 U17942 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14684) );
  INV_X1 U17943 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20873) );
  NAND4_X1 U17944 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(P1_REIP_REG_10__SCAN_IN), .A4(P1_REIP_REG_9__SCAN_IN), .ZN(n14705)
         );
  NOR2_X1 U17945 ( .A1(n20873), .A2(n14705), .ZN(n16006) );
  NAND3_X1 U17946 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n14495), .A3(n16006), 
        .ZN(n14497) );
  NAND3_X1 U17947 ( .A1(n15995), .A2(P1_REIP_REG_16__SCAN_IN), .A3(
        P1_REIP_REG_15__SCAN_IN), .ZN(n14683) );
  NAND2_X1 U17948 ( .A1(n14653), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14656) );
  INV_X1 U17949 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n14951) );
  NAND2_X1 U17950 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n14496) );
  NAND2_X1 U17951 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14566) );
  INV_X1 U17952 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21019) );
  NOR2_X1 U17953 ( .A1(n14566), .A2(n21019), .ZN(n14504) );
  NAND2_X1 U17954 ( .A1(n14565), .A2(n14504), .ZN(n14555) );
  NAND2_X1 U17955 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n14507) );
  NAND2_X1 U17956 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14509) );
  NOR3_X1 U17957 ( .A1(n14535), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14509), 
        .ZN(n14512) );
  NOR2_X1 U17958 ( .A1(n14498), .A2(n14497), .ZN(n14694) );
  NAND4_X1 U17959 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .A4(n14694), .ZN(n14499) );
  NAND2_X1 U17960 ( .A1(n20042), .A2(n14499), .ZN(n14682) );
  NAND3_X1 U17961 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(P1_REIP_REG_20__SCAN_IN), .ZN(n14500) );
  NAND2_X1 U17962 ( .A1(n20042), .A2(n14500), .ZN(n14501) );
  NAND2_X1 U17963 ( .A1(n14682), .A2(n14501), .ZN(n14644) );
  NAND3_X1 U17964 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(P1_REIP_REG_21__SCAN_IN), .ZN(n14502) );
  AND2_X1 U17965 ( .A1(n20042), .A2(n14502), .ZN(n14503) );
  INV_X1 U17966 ( .A(n14504), .ZN(n14505) );
  AND2_X1 U17967 ( .A1(n20042), .A2(n14505), .ZN(n14506) );
  NOR2_X1 U17968 ( .A1(n14604), .A2(n14506), .ZN(n14564) );
  NAND2_X1 U17969 ( .A1(n20042), .A2(n14507), .ZN(n14508) );
  NAND2_X1 U17970 ( .A1(n14564), .A2(n14508), .ZN(n14536) );
  AOI21_X1 U17971 ( .B1(n14509), .B2(n20042), .A(n14536), .ZN(n14521) );
  AOI22_X1 U17972 ( .A1(n20088), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20091), .ZN(n14510) );
  OAI21_X1 U17973 ( .B1(n14521), .B2(n21032), .A(n14510), .ZN(n14511) );
  AOI211_X1 U17974 ( .C1(n15022), .C2(n20089), .A(n14512), .B(n14511), .ZN(
        n14513) );
  OAI21_X1 U17975 ( .B1(n14514), .B2(n20029), .A(n14513), .ZN(P1_U2809) );
  INV_X1 U17976 ( .A(n20088), .ZN(n14519) );
  OAI22_X1 U17977 ( .A1(n20067), .A2(n14515), .B1(n14860), .B2(n20078), .ZN(
        n14516) );
  INV_X1 U17978 ( .A(n14516), .ZN(n14518) );
  INV_X1 U17979 ( .A(n14520), .ZN(n14525) );
  NOR2_X1 U17980 ( .A1(n14535), .A2(n21052), .ZN(n14523) );
  INV_X1 U17981 ( .A(n14521), .ZN(n14522) );
  OAI21_X1 U17982 ( .B1(n14523), .B2(P1_REIP_REG_30__SCAN_IN), .A(n14522), 
        .ZN(n14524) );
  OAI211_X1 U17983 ( .C1(n14863), .C2(n20029), .A(n14525), .B(n14524), .ZN(
        P1_U2810) );
  NAND2_X1 U17984 ( .A1(n14526), .A2(n20058), .ZN(n14534) );
  INV_X1 U17985 ( .A(n14527), .ZN(n15040) );
  NAND2_X1 U17986 ( .A1(n14536), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14530) );
  AOI22_X1 U17987 ( .A1(n20093), .A2(n14528), .B1(n20091), .B2(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14529) );
  OAI211_X1 U17988 ( .C1(n14531), .C2(n14519), .A(n14530), .B(n14529), .ZN(
        n14532) );
  AOI21_X1 U17989 ( .B1(n15040), .B2(n20089), .A(n14532), .ZN(n14533) );
  OAI211_X1 U17990 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(n14535), .A(n14534), 
        .B(n14533), .ZN(P1_U2811) );
  INV_X1 U17991 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21065) );
  NAND2_X1 U17992 ( .A1(n21065), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14544) );
  NAND2_X1 U17993 ( .A1(n14872), .A2(n20058), .ZN(n14543) );
  NAND2_X1 U17994 ( .A1(n14536), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14539) );
  INV_X1 U17995 ( .A(n14870), .ZN(n14537) );
  AOI22_X1 U17996 ( .A1(n20093), .A2(n14537), .B1(n20091), .B2(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14538) );
  OAI211_X1 U17997 ( .C1(n14540), .C2(n14519), .A(n14539), .B(n14538), .ZN(
        n14541) );
  AOI21_X1 U17998 ( .B1(n10171), .B2(n20089), .A(n14541), .ZN(n14542) );
  OAI211_X1 U17999 ( .C1(n14555), .C2(n14544), .A(n14543), .B(n14542), .ZN(
        P1_U2812) );
  OAI21_X1 U18000 ( .B1(n14545), .B2(n14546), .A(n12833), .ZN(n14793) );
  INV_X1 U18001 ( .A(n14793), .ZN(n14881) );
  NAND2_X1 U18002 ( .A1(n14881), .A2(n20058), .ZN(n14554) );
  AND2_X1 U18003 ( .A1(n14558), .A2(n14547), .ZN(n14548) );
  NOR2_X1 U18004 ( .A1(n14549), .A2(n14548), .ZN(n15056) );
  INV_X1 U18005 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21060) );
  AOI22_X1 U18006 ( .A1(n20093), .A2(n14877), .B1(n20091), .B2(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14551) );
  NAND2_X1 U18007 ( .A1(n20088), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n14550) );
  OAI211_X1 U18008 ( .C1(n14564), .C2(n21060), .A(n14551), .B(n14550), .ZN(
        n14552) );
  AOI21_X1 U18009 ( .B1(n15056), .B2(n20089), .A(n14552), .ZN(n14553) );
  OAI211_X1 U18010 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14555), .A(n14554), 
        .B(n14553), .ZN(P1_U2813) );
  AOI21_X1 U18011 ( .B1(n14557), .B2(n14556), .A(n14545), .ZN(n14890) );
  INV_X1 U18012 ( .A(n14890), .ZN(n14798) );
  INV_X1 U18013 ( .A(n14558), .ZN(n14559) );
  AOI21_X1 U18014 ( .B1(n14560), .B2(n14573), .A(n14559), .ZN(n15060) );
  OAI22_X1 U18015 ( .A1(n20067), .A2(n14561), .B1(n14888), .B2(n20078), .ZN(
        n14562) );
  AOI21_X1 U18016 ( .B1(n20088), .B2(P1_EBX_REG_26__SCAN_IN), .A(n14562), .ZN(
        n14563) );
  OAI21_X1 U18017 ( .B1(n14564), .B2(n21019), .A(n14563), .ZN(n14568) );
  INV_X1 U18018 ( .A(n14565), .ZN(n14580) );
  NOR3_X1 U18019 ( .A1(n14580), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n14566), 
        .ZN(n14567) );
  AOI211_X1 U18020 ( .C1(n15060), .C2(n20089), .A(n14568), .B(n14567), .ZN(
        n14569) );
  OAI21_X1 U18021 ( .B1(n14798), .B2(n20029), .A(n14569), .ZN(P1_U2814) );
  OR2_X1 U18022 ( .A1(n14570), .A2(n14585), .ZN(n14583) );
  INV_X1 U18023 ( .A(n14556), .ZN(n14571) );
  INV_X1 U18024 ( .A(n14573), .ZN(n14574) );
  AOI21_X1 U18025 ( .B1(n14575), .B2(n14586), .A(n14574), .ZN(n15067) );
  INV_X1 U18026 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14577) );
  AOI22_X1 U18027 ( .A1(n20093), .A2(n14896), .B1(n20091), .B2(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14576) );
  OAI21_X1 U18028 ( .B1(n14519), .B2(n14577), .A(n14576), .ZN(n14579) );
  INV_X1 U18029 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14907) );
  NOR3_X1 U18030 ( .A1(n14580), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n14907), 
        .ZN(n14578) );
  AOI211_X1 U18031 ( .C1(n15067), .C2(n20089), .A(n14579), .B(n14578), .ZN(
        n14582) );
  NOR2_X1 U18032 ( .A1(n14580), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14592) );
  OAI21_X1 U18033 ( .B1(n14592), .B2(n14604), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14581) );
  OAI211_X1 U18034 ( .C1(n14802), .C2(n20029), .A(n14582), .B(n14581), .ZN(
        P1_U2815) );
  INV_X1 U18035 ( .A(n14583), .ZN(n14584) );
  AOI21_X1 U18036 ( .B1(n14585), .B2(n14570), .A(n14584), .ZN(n14911) );
  INV_X1 U18037 ( .A(n14911), .ZN(n14807) );
  OAI21_X1 U18038 ( .B1(n14601), .B2(n14587), .A(n14586), .ZN(n14752) );
  INV_X1 U18039 ( .A(n14752), .ZN(n15075) );
  INV_X1 U18040 ( .A(n14604), .ZN(n14591) );
  OAI22_X1 U18041 ( .A1(n20067), .A2(n14588), .B1(n14909), .B2(n20078), .ZN(
        n14589) );
  AOI21_X1 U18042 ( .B1(n20088), .B2(P1_EBX_REG_24__SCAN_IN), .A(n14589), .ZN(
        n14590) );
  OAI21_X1 U18043 ( .B1(n14591), .B2(n14907), .A(n14590), .ZN(n14593) );
  AOI211_X1 U18044 ( .C1(n15075), .C2(n20089), .A(n14593), .B(n14592), .ZN(
        n14594) );
  OAI21_X1 U18045 ( .B1(n14807), .B2(n20029), .A(n14594), .ZN(P1_U2816) );
  OAI21_X1 U18046 ( .B1(n14595), .B2(n14596), .A(n14570), .ZN(n14915) );
  INV_X1 U18047 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14598) );
  INV_X1 U18048 ( .A(n14597), .ZN(n14918) );
  OAI22_X1 U18049 ( .A1(n20067), .A2(n14598), .B1(n14918), .B2(n20078), .ZN(
        n14603) );
  NOR2_X1 U18050 ( .A1(n14614), .A2(n14599), .ZN(n14600) );
  OR2_X1 U18051 ( .A1(n14601), .A2(n14600), .ZN(n15088) );
  NOR2_X1 U18052 ( .A1(n15088), .A2(n20086), .ZN(n14602) );
  AOI211_X1 U18053 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n20088), .A(n14603), .B(
        n14602), .ZN(n14607) );
  OAI21_X1 U18054 ( .B1(n14605), .B2(P1_REIP_REG_23__SCAN_IN), .A(n14604), 
        .ZN(n14606) );
  OAI211_X1 U18055 ( .C1(n14915), .C2(n20029), .A(n14607), .B(n14606), .ZN(
        P1_U2817) );
  INV_X1 U18056 ( .A(n14608), .ZN(n14611) );
  INV_X1 U18057 ( .A(n14609), .ZN(n14610) );
  AOI21_X1 U18058 ( .B1(n14611), .B2(n14610), .A(n14595), .ZN(n14928) );
  NAND2_X1 U18059 ( .A1(n14928), .A2(n20058), .ZN(n14624) );
  AND2_X1 U18060 ( .A1(n14627), .A2(n14612), .ZN(n14613) );
  NOR2_X1 U18061 ( .A1(n14614), .A2(n14613), .ZN(n15109) );
  NAND2_X1 U18062 ( .A1(n20088), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n14617) );
  INV_X1 U18063 ( .A(n14926), .ZN(n14615) );
  AOI22_X1 U18064 ( .A1(n20093), .A2(n14615), .B1(n20091), .B2(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14616) );
  NAND2_X1 U18065 ( .A1(n14617), .A2(n14616), .ZN(n14618) );
  AOI21_X1 U18066 ( .B1(n15109), .B2(n20089), .A(n14618), .ZN(n14623) );
  INV_X1 U18067 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20994) );
  NAND2_X1 U18068 ( .A1(n20994), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n14619) );
  NOR2_X1 U18069 ( .A1(n14643), .A2(n14619), .ZN(n14633) );
  OAI21_X1 U18070 ( .B1(n14633), .B2(n14644), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14622) );
  INV_X1 U18071 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21059) );
  NAND2_X1 U18072 ( .A1(n14620), .A2(n21059), .ZN(n14621) );
  NAND4_X1 U18073 ( .A1(n14624), .A2(n14623), .A3(n14622), .A4(n14621), .ZN(
        P1_U2818) );
  AOI21_X1 U18074 ( .B1(n14626), .B2(n14625), .A(n14609), .ZN(n14937) );
  INV_X1 U18075 ( .A(n14937), .ZN(n14818) );
  INV_X1 U18076 ( .A(n14627), .ZN(n14628) );
  AOI21_X1 U18077 ( .B1(n14629), .B2(n14639), .A(n14628), .ZN(n15117) );
  INV_X1 U18078 ( .A(n14644), .ZN(n14632) );
  AOI22_X1 U18079 ( .A1(n20093), .A2(n14933), .B1(n20091), .B2(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14631) );
  NAND2_X1 U18080 ( .A1(n20088), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n14630) );
  OAI211_X1 U18081 ( .C1(n14632), .C2(n20994), .A(n14631), .B(n14630), .ZN(
        n14634) );
  AOI211_X1 U18082 ( .C1(n15117), .C2(n20089), .A(n14634), .B(n14633), .ZN(
        n14635) );
  OAI21_X1 U18083 ( .B1(n14818), .B2(n20029), .A(n14635), .ZN(P1_U2819) );
  XOR2_X1 U18084 ( .A(n14637), .B(n14636), .Z(n14945) );
  OAI22_X1 U18085 ( .A1(n20067), .A2(n14638), .B1(n14943), .B2(n20078), .ZN(
        n14642) );
  OAI21_X1 U18086 ( .B1(n14652), .B2(n14640), .A(n14639), .ZN(n15121) );
  NOR2_X1 U18087 ( .A1(n15121), .A2(n20086), .ZN(n14641) );
  AOI211_X1 U18088 ( .C1(n20088), .C2(P1_EBX_REG_20__SCAN_IN), .A(n14642), .B(
        n14641), .ZN(n14647) );
  INV_X1 U18089 ( .A(n14643), .ZN(n14645) );
  OAI21_X1 U18090 ( .B1(n14645), .B2(P1_REIP_REG_20__SCAN_IN), .A(n14644), 
        .ZN(n14646) );
  OAI211_X1 U18091 ( .C1(n14826), .C2(n20029), .A(n14647), .B(n14646), .ZN(
        P1_U2820) );
  OAI21_X1 U18092 ( .B1(n14648), .B2(n14649), .A(n14636), .ZN(n14949) );
  NOR2_X1 U18093 ( .A1(n14665), .A2(n14650), .ZN(n14651) );
  OR2_X1 U18094 ( .A1(n14652), .A2(n14651), .ZN(n14759) );
  INV_X1 U18095 ( .A(n14759), .ZN(n15140) );
  INV_X1 U18096 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n14958) );
  NAND2_X1 U18097 ( .A1(n14653), .A2(n14958), .ZN(n14668) );
  AOI21_X1 U18098 ( .B1(n14682), .B2(n14668), .A(n14951), .ZN(n14658) );
  AOI21_X1 U18099 ( .B1(n20091), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n20167), .ZN(n14655) );
  AOI22_X1 U18100 ( .A1(n20088), .A2(P1_EBX_REG_19__SCAN_IN), .B1(n14950), 
        .B2(n20093), .ZN(n14654) );
  OAI211_X1 U18101 ( .C1(P1_REIP_REG_19__SCAN_IN), .C2(n14656), .A(n14655), 
        .B(n14654), .ZN(n14657) );
  AOI211_X1 U18102 ( .C1(n15140), .C2(n20089), .A(n14658), .B(n14657), .ZN(
        n14659) );
  OAI21_X1 U18103 ( .B1(n14949), .B2(n20029), .A(n14659), .ZN(P1_U2821) );
  INV_X1 U18104 ( .A(n14648), .ZN(n14661) );
  OAI21_X1 U18105 ( .B1(n14662), .B2(n14660), .A(n14661), .ZN(n14959) );
  AND2_X1 U18106 ( .A1(n14678), .A2(n14663), .ZN(n14664) );
  NOR2_X1 U18107 ( .A1(n14665), .A2(n14664), .ZN(n16086) );
  INV_X1 U18108 ( .A(n14962), .ZN(n14670) );
  OAI22_X1 U18109 ( .A1(n14666), .A2(n14519), .B1(n14682), .B2(n14958), .ZN(
        n14667) );
  AOI211_X1 U18110 ( .C1(n20091), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20167), .B(n14667), .ZN(n14669) );
  OAI211_X1 U18111 ( .C1(n20078), .C2(n14670), .A(n14669), .B(n14668), .ZN(
        n14671) );
  AOI21_X1 U18112 ( .B1(n16086), .B2(n20089), .A(n14671), .ZN(n14672) );
  OAI21_X1 U18113 ( .B1(n14959), .B2(n20029), .A(n14672), .ZN(P1_U2822) );
  AOI21_X1 U18114 ( .B1(n14674), .B2(n14673), .A(n14660), .ZN(n14978) );
  INV_X1 U18115 ( .A(n14978), .ZN(n14838) );
  NAND2_X1 U18116 ( .A1(n14676), .A2(n14675), .ZN(n14677) );
  AND2_X1 U18117 ( .A1(n14678), .A2(n14677), .ZN(n16094) );
  NOR2_X1 U18118 ( .A1(n20078), .A2(n14976), .ZN(n14679) );
  AOI211_X1 U18119 ( .C1(n20091), .C2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n20167), .B(n14679), .ZN(n14680) );
  OAI21_X1 U18120 ( .B1(n14681), .B2(n14519), .A(n14680), .ZN(n14686) );
  AOI21_X1 U18121 ( .B1(n14684), .B2(n14683), .A(n14682), .ZN(n14685) );
  AOI211_X1 U18122 ( .C1(n16094), .C2(n20089), .A(n14686), .B(n14685), .ZN(
        n14687) );
  OAI21_X1 U18123 ( .B1(n14838), .B2(n20029), .A(n14687), .ZN(P1_U2823) );
  INV_X1 U18124 ( .A(n14689), .ZN(n14765) );
  AOI21_X1 U18125 ( .B1(n14690), .B2(n14688), .A(n14689), .ZN(n14990) );
  INV_X1 U18126 ( .A(n14990), .ZN(n14847) );
  AOI21_X1 U18127 ( .B1(n14775), .B2(n14692), .A(n14691), .ZN(n16102) );
  INV_X1 U18128 ( .A(n20042), .ZN(n14693) );
  OR2_X1 U18129 ( .A1(n14694), .A2(n14693), .ZN(n16007) );
  INV_X1 U18130 ( .A(n16007), .ZN(n15997) );
  AOI22_X1 U18131 ( .A1(n20088), .A2(P1_EBX_REG_15__SCAN_IN), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n15997), .ZN(n14695) );
  OAI211_X1 U18132 ( .C1(n20067), .C2(n14696), .A(n14695), .B(n20064), .ZN(
        n14698) );
  NOR2_X1 U18133 ( .A1(n20078), .A2(n14988), .ZN(n14697) );
  AOI211_X1 U18134 ( .C1(n16102), .C2(n20089), .A(n14698), .B(n14697), .ZN(
        n14700) );
  INV_X1 U18135 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20875) );
  AND2_X1 U18136 ( .A1(n20875), .A2(n15995), .ZN(n15996) );
  INV_X1 U18137 ( .A(n15996), .ZN(n14699) );
  OAI211_X1 U18138 ( .C1(n14847), .C2(n20029), .A(n14700), .B(n14699), .ZN(
        P1_U2825) );
  AOI21_X1 U18139 ( .B1(n14702), .B2(n14002), .A(n14701), .ZN(n14999) );
  INV_X1 U18140 ( .A(n14999), .ZN(n14855) );
  INV_X1 U18141 ( .A(n14705), .ZN(n14703) );
  OAI21_X1 U18142 ( .B1(n14703), .B2(n20044), .A(n20026), .ZN(n16018) );
  NOR2_X1 U18143 ( .A1(n20044), .A2(n14704), .ZN(n20023) );
  NAND2_X1 U18144 ( .A1(n20023), .A2(n20873), .ZN(n14706) );
  NOR2_X1 U18145 ( .A1(n14706), .A2(n14705), .ZN(n14714) );
  NAND2_X1 U18146 ( .A1(n14708), .A2(n14707), .ZN(n14709) );
  NAND2_X1 U18147 ( .A1(n14773), .A2(n14709), .ZN(n15143) );
  NAND2_X1 U18148 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14710) );
  OAI211_X1 U18149 ( .C1(n14997), .C2(n20078), .A(n14710), .B(n20064), .ZN(
        n14711) );
  AOI21_X1 U18150 ( .B1(n20088), .B2(P1_EBX_REG_13__SCAN_IN), .A(n14711), .ZN(
        n14712) );
  OAI21_X1 U18151 ( .B1(n15143), .B2(n20086), .A(n14712), .ZN(n14713) );
  AOI211_X1 U18152 ( .C1(n16018), .C2(P1_REIP_REG_13__SCAN_IN), .A(n14714), 
        .B(n14713), .ZN(n14715) );
  OAI21_X1 U18153 ( .B1(n14855), .B2(n20029), .A(n14715), .ZN(P1_U2827) );
  INV_X1 U18154 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14716) );
  NOR2_X1 U18155 ( .A1(n14716), .A2(n13869), .ZN(n16017) );
  OAI21_X1 U18156 ( .B1(n16017), .B2(n20044), .A(n20026), .ZN(n16027) );
  INV_X1 U18157 ( .A(n16129), .ZN(n14722) );
  NAND3_X1 U18158 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n20023), .A3(n14716), 
        .ZN(n14721) );
  AOI21_X1 U18159 ( .B1(n20091), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20167), .ZN(n14717) );
  OAI21_X1 U18160 ( .B1(n20078), .B2(n14718), .A(n14717), .ZN(n14719) );
  AOI21_X1 U18161 ( .B1(n20088), .B2(P1_EBX_REG_10__SCAN_IN), .A(n14719), .ZN(
        n14720) );
  OAI211_X1 U18162 ( .C1(n20086), .C2(n14722), .A(n14721), .B(n14720), .ZN(
        n14723) );
  AOI21_X1 U18163 ( .B1(n16027), .B2(P1_REIP_REG_10__SCAN_IN), .A(n14723), 
        .ZN(n14724) );
  OAI21_X1 U18164 ( .B1(n14725), .B2(n20029), .A(n14724), .ZN(P1_U2830) );
  AOI21_X1 U18165 ( .B1(n20051), .B2(P1_REIP_REG_1__SCAN_IN), .A(
        P1_REIP_REG_2__SCAN_IN), .ZN(n14736) );
  INV_X1 U18166 ( .A(n14726), .ZN(n20050) );
  NAND2_X1 U18167 ( .A1(n20050), .A2(n14727), .ZN(n20043) );
  NAND2_X1 U18168 ( .A1(n20042), .A2(n20043), .ZN(n20103) );
  NAND2_X1 U18169 ( .A1(n14728), .A2(n20099), .ZN(n14735) );
  INV_X1 U18170 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14730) );
  OAI22_X1 U18171 ( .A1(n20067), .A2(n14730), .B1(n14729), .B2(n20078), .ZN(
        n14731) );
  AOI21_X1 U18172 ( .B1(P1_EBX_REG_2__SCAN_IN), .B2(n20088), .A(n14731), .ZN(
        n14732) );
  OAI21_X1 U18173 ( .B1(n20086), .B2(n20199), .A(n14732), .ZN(n14733) );
  AOI21_X1 U18174 ( .B1(n20247), .B2(n20094), .A(n14733), .ZN(n14734) );
  OAI211_X1 U18175 ( .C1(n14736), .C2(n20103), .A(n14735), .B(n14734), .ZN(
        P1_U2838) );
  INV_X1 U18176 ( .A(n20094), .ZN(n14740) );
  NAND2_X1 U18177 ( .A1(n20088), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n14738) );
  OAI21_X1 U18178 ( .B1(n20093), .B2(n20091), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14737) );
  OAI211_X1 U18179 ( .C1(n14740), .C2(n14739), .A(n14738), .B(n14737), .ZN(
        n14743) );
  NOR2_X1 U18180 ( .A1(n20086), .A2(n14741), .ZN(n14742) );
  AOI211_X1 U18181 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(n20042), .A(n14743), .B(
        n14742), .ZN(n14744) );
  OAI21_X1 U18182 ( .B1(n14746), .B2(n14745), .A(n14744), .ZN(P1_U2840) );
  INV_X1 U18183 ( .A(n15022), .ZN(n14748) );
  INV_X1 U18184 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14747) );
  OAI22_X1 U18185 ( .A1(n14748), .A2(n14777), .B1(n14778), .B2(n14747), .ZN(
        P1_U2841) );
  AOI22_X1 U18186 ( .A1(n15056), .A2(n11194), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n14769), .ZN(n14749) );
  OAI21_X1 U18187 ( .B1(n14793), .B2(n14779), .A(n14749), .ZN(P1_U2845) );
  AOI22_X1 U18188 ( .A1(n15060), .A2(n11194), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n14769), .ZN(n14750) );
  OAI21_X1 U18189 ( .B1(n14798), .B2(n14779), .A(n14750), .ZN(P1_U2846) );
  AOI22_X1 U18190 ( .A1(n15067), .A2(n11194), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(n14769), .ZN(n14751) );
  OAI21_X1 U18191 ( .B1(n14802), .B2(n14779), .A(n14751), .ZN(P1_U2847) );
  OAI222_X1 U18192 ( .A1(n14807), .A2(n14779), .B1(n14753), .B2(n14778), .C1(
        n14752), .C2(n14777), .ZN(P1_U2848) );
  OAI222_X1 U18193 ( .A1(n14915), .A2(n14779), .B1(n14754), .B2(n14778), .C1(
        n15088), .C2(n14777), .ZN(P1_U2849) );
  INV_X1 U18194 ( .A(n14928), .ZN(n14814) );
  AOI22_X1 U18195 ( .A1(n15109), .A2(n11194), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n14769), .ZN(n14755) );
  OAI21_X1 U18196 ( .B1(n14814), .B2(n14779), .A(n14755), .ZN(P1_U2850) );
  AOI22_X1 U18197 ( .A1(n15117), .A2(n11194), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n14769), .ZN(n14756) );
  OAI21_X1 U18198 ( .B1(n14818), .B2(n14779), .A(n14756), .ZN(P1_U2851) );
  INV_X1 U18199 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14757) );
  OAI222_X1 U18200 ( .A1(n14826), .A2(n14779), .B1(n14778), .B2(n14757), .C1(
        n15121), .C2(n14777), .ZN(P1_U2852) );
  OAI22_X1 U18201 ( .A1(n14759), .A2(n14777), .B1(n14758), .B2(n14778), .ZN(
        n14760) );
  INV_X1 U18202 ( .A(n14760), .ZN(n14761) );
  OAI21_X1 U18203 ( .B1(n14949), .B2(n14779), .A(n14761), .ZN(P1_U2853) );
  AOI22_X1 U18204 ( .A1(n16086), .A2(n11194), .B1(P1_EBX_REG_18__SCAN_IN), 
        .B2(n14769), .ZN(n14762) );
  OAI21_X1 U18205 ( .B1(n14959), .B2(n14779), .A(n14762), .ZN(P1_U2854) );
  AOI22_X1 U18206 ( .A1(n16094), .A2(n11194), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14769), .ZN(n14763) );
  OAI21_X1 U18207 ( .B1(n14838), .B2(n14779), .A(n14763), .ZN(P1_U2855) );
  INV_X1 U18208 ( .A(n14673), .ZN(n14764) );
  AOI21_X1 U18209 ( .B1(n14766), .B2(n14765), .A(n14764), .ZN(n16034) );
  INV_X1 U18210 ( .A(n16034), .ZN(n14845) );
  INV_X1 U18211 ( .A(n14767), .ZN(n16002) );
  AOI22_X1 U18212 ( .A1(n16002), .A2(n11194), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n14769), .ZN(n14768) );
  OAI21_X1 U18213 ( .B1(n14845), .B2(n14779), .A(n14768), .ZN(P1_U2856) );
  AOI22_X1 U18214 ( .A1(n16102), .A2(n11194), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n14769), .ZN(n14770) );
  OAI21_X1 U18215 ( .B1(n14847), .B2(n14779), .A(n14770), .ZN(P1_U2857) );
  OAI21_X1 U18216 ( .B1(n14701), .B2(n14771), .A(n14688), .ZN(n16011) );
  INV_X1 U18217 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14776) );
  NAND2_X1 U18218 ( .A1(n14773), .A2(n14772), .ZN(n14774) );
  NAND2_X1 U18219 ( .A1(n14775), .A2(n14774), .ZN(n16108) );
  OAI222_X1 U18220 ( .A1(n16011), .A2(n14779), .B1(n14776), .B2(n14778), .C1(
        n16108), .C2(n14777), .ZN(P1_U2858) );
  OAI222_X1 U18221 ( .A1(n14855), .A2(n14779), .B1(n14778), .B2(n11133), .C1(
        n15143), .C2(n14777), .ZN(P1_U2859) );
  INV_X1 U18222 ( .A(DATAI_14_), .ZN(n14781) );
  NAND2_X1 U18223 ( .A1(n20238), .A2(BUF1_REG_14__SCAN_IN), .ZN(n14780) );
  OAI21_X1 U18224 ( .B1(n20238), .B2(n14781), .A(n14780), .ZN(n20148) );
  AOI22_X1 U18225 ( .A1(n14820), .A2(n20148), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n14849), .ZN(n14782) );
  OAI21_X1 U18226 ( .B1(n14783), .B2(n14823), .A(n14782), .ZN(n14784) );
  AOI21_X1 U18227 ( .B1(n11080), .B2(DATAI_30_), .A(n14784), .ZN(n14785) );
  OAI21_X1 U18228 ( .B1(n14863), .B2(n14848), .A(n14785), .ZN(P1_U2874) );
  OAI22_X1 U18229 ( .A1(n14840), .A2(n20142), .B1(n14853), .B2(n13232), .ZN(
        n14786) );
  AOI21_X1 U18230 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n14842), .A(n14786), .ZN(
        n14788) );
  NAND2_X1 U18231 ( .A1(n11080), .A2(DATAI_28_), .ZN(n14787) );
  OAI211_X1 U18232 ( .C1(n14789), .C2(n14848), .A(n14788), .B(n14787), .ZN(
        P1_U2876) );
  OAI22_X1 U18233 ( .A1(n14840), .A2(n20139), .B1(n14853), .B2(n13235), .ZN(
        n14790) );
  AOI21_X1 U18234 ( .B1(BUF1_REG_27__SCAN_IN), .B2(n14842), .A(n14790), .ZN(
        n14792) );
  NAND2_X1 U18235 ( .A1(n11080), .A2(DATAI_27_), .ZN(n14791) );
  OAI211_X1 U18236 ( .C1(n14793), .C2(n14848), .A(n14792), .B(n14791), .ZN(
        P1_U2877) );
  OAI22_X1 U18237 ( .A1(n14840), .A2(n20136), .B1(n14853), .B2(n14794), .ZN(
        n14795) );
  AOI21_X1 U18238 ( .B1(BUF1_REG_26__SCAN_IN), .B2(n14842), .A(n14795), .ZN(
        n14797) );
  NAND2_X1 U18239 ( .A1(n11080), .A2(DATAI_26_), .ZN(n14796) );
  OAI211_X1 U18240 ( .C1(n14798), .C2(n14848), .A(n14797), .B(n14796), .ZN(
        P1_U2878) );
  OAI22_X1 U18241 ( .A1(n14840), .A2(n20132), .B1(n14853), .B2(n13240), .ZN(
        n14799) );
  AOI21_X1 U18242 ( .B1(n14842), .B2(BUF1_REG_25__SCAN_IN), .A(n14799), .ZN(
        n14801) );
  NAND2_X1 U18243 ( .A1(n11080), .A2(DATAI_25_), .ZN(n14800) );
  OAI211_X1 U18244 ( .C1(n14802), .C2(n14848), .A(n14801), .B(n14800), .ZN(
        P1_U2879) );
  OAI22_X1 U18245 ( .A1(n14840), .A2(n20129), .B1(n14853), .B2(n14803), .ZN(
        n14804) );
  AOI21_X1 U18246 ( .B1(n14842), .B2(BUF1_REG_24__SCAN_IN), .A(n14804), .ZN(
        n14806) );
  NAND2_X1 U18247 ( .A1(n11080), .A2(DATAI_24_), .ZN(n14805) );
  OAI211_X1 U18248 ( .C1(n14807), .C2(n14848), .A(n14806), .B(n14805), .ZN(
        P1_U2880) );
  OAI22_X1 U18249 ( .A1(n14840), .A2(n20292), .B1(n14853), .B2(n13245), .ZN(
        n14808) );
  AOI21_X1 U18250 ( .B1(n14842), .B2(BUF1_REG_23__SCAN_IN), .A(n14808), .ZN(
        n14810) );
  NAND2_X1 U18251 ( .A1(n11080), .A2(DATAI_23_), .ZN(n14809) );
  OAI211_X1 U18252 ( .C1(n14915), .C2(n14848), .A(n14810), .B(n14809), .ZN(
        P1_U2881) );
  OAI22_X1 U18253 ( .A1(n14840), .A2(n20281), .B1(n14853), .B2(n13550), .ZN(
        n14811) );
  AOI21_X1 U18254 ( .B1(n14842), .B2(BUF1_REG_22__SCAN_IN), .A(n14811), .ZN(
        n14813) );
  NAND2_X1 U18255 ( .A1(n11080), .A2(DATAI_22_), .ZN(n14812) );
  OAI211_X1 U18256 ( .C1(n14814), .C2(n14848), .A(n14813), .B(n14812), .ZN(
        P1_U2882) );
  OAI22_X1 U18257 ( .A1(n14840), .A2(n20276), .B1(n14853), .B2(n13552), .ZN(
        n14815) );
  AOI21_X1 U18258 ( .B1(n14842), .B2(BUF1_REG_21__SCAN_IN), .A(n14815), .ZN(
        n14817) );
  NAND2_X1 U18259 ( .A1(n11080), .A2(DATAI_21_), .ZN(n14816) );
  OAI211_X1 U18260 ( .C1(n14818), .C2(n14848), .A(n14817), .B(n14816), .ZN(
        P1_U2883) );
  INV_X1 U18261 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n14822) );
  AOI22_X1 U18262 ( .A1(n14820), .A2(n14819), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n14849), .ZN(n14821) );
  OAI21_X1 U18263 ( .B1(n14823), .B2(n14822), .A(n14821), .ZN(n14824) );
  AOI21_X1 U18264 ( .B1(n11080), .B2(DATAI_20_), .A(n14824), .ZN(n14825) );
  OAI21_X1 U18265 ( .B1(n14826), .B2(n14848), .A(n14825), .ZN(P1_U2884) );
  OAI22_X1 U18266 ( .A1(n14840), .A2(n20268), .B1(n14853), .B2(n13243), .ZN(
        n14827) );
  AOI21_X1 U18267 ( .B1(n14842), .B2(BUF1_REG_19__SCAN_IN), .A(n14827), .ZN(
        n14829) );
  NAND2_X1 U18268 ( .A1(n11080), .A2(DATAI_19_), .ZN(n14828) );
  OAI211_X1 U18269 ( .C1(n14949), .C2(n14848), .A(n14829), .B(n14828), .ZN(
        P1_U2885) );
  OAI22_X1 U18270 ( .A1(n14840), .A2(n20264), .B1(n14853), .B2(n14830), .ZN(
        n14831) );
  AOI21_X1 U18271 ( .B1(n14842), .B2(BUF1_REG_18__SCAN_IN), .A(n14831), .ZN(
        n14833) );
  NAND2_X1 U18272 ( .A1(n11080), .A2(DATAI_18_), .ZN(n14832) );
  OAI211_X1 U18273 ( .C1(n14959), .C2(n14848), .A(n14833), .B(n14832), .ZN(
        P1_U2886) );
  OAI22_X1 U18274 ( .A1(n14840), .A2(n20259), .B1(n14853), .B2(n14834), .ZN(
        n14835) );
  AOI21_X1 U18275 ( .B1(n14842), .B2(BUF1_REG_17__SCAN_IN), .A(n14835), .ZN(
        n14837) );
  NAND2_X1 U18276 ( .A1(n11080), .A2(DATAI_17_), .ZN(n14836) );
  OAI211_X1 U18277 ( .C1(n14838), .C2(n14848), .A(n14837), .B(n14836), .ZN(
        P1_U2887) );
  OAI22_X1 U18278 ( .A1(n14840), .A2(n20251), .B1(n14853), .B2(n14839), .ZN(
        n14841) );
  AOI21_X1 U18279 ( .B1(n14842), .B2(BUF1_REG_16__SCAN_IN), .A(n14841), .ZN(
        n14844) );
  NAND2_X1 U18280 ( .A1(n11080), .A2(DATAI_16_), .ZN(n14843) );
  OAI211_X1 U18281 ( .C1(n14845), .C2(n14848), .A(n14844), .B(n14843), .ZN(
        P1_U2888) );
  OAI222_X1 U18282 ( .A1(n14848), .A2(n14847), .B1(n14853), .B2(n13252), .C1(
        n14852), .C2(n14846), .ZN(P1_U2889) );
  INV_X1 U18283 ( .A(n14852), .ZN(n14850) );
  AOI22_X1 U18284 ( .A1(n14850), .A2(n20148), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14849), .ZN(n14851) );
  OAI21_X1 U18285 ( .B1(n16011), .B2(n14848), .A(n14851), .ZN(P1_U2890) );
  INV_X1 U18286 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14854) );
  OAI222_X1 U18287 ( .A1(n14855), .A2(n14848), .B1(n14854), .B2(n14853), .C1(
        n14852), .C2(n20145), .ZN(P1_U2891) );
  NAND2_X1 U18288 ( .A1(n20167), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15030) );
  NAND2_X1 U18289 ( .A1(n20168), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14859) );
  OAI211_X1 U18290 ( .C1(n20178), .C2(n14860), .A(n15030), .B(n14859), .ZN(
        n14861) );
  AOI21_X1 U18291 ( .B1(n15032), .B2(n20174), .A(n14861), .ZN(n14862) );
  OAI21_X1 U18292 ( .B1(n14863), .B2(n16049), .A(n14862), .ZN(P1_U2969) );
  NAND2_X1 U18293 ( .A1(n14972), .A2(n15061), .ZN(n14884) );
  NAND2_X1 U18294 ( .A1(n14884), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14864) );
  OAI22_X1 U18295 ( .A1(n14883), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n14914), .B2(n14864), .ZN(n14867) );
  MUX2_X1 U18296 ( .A(n14865), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n9673), .Z(n14866) );
  NAND2_X1 U18297 ( .A1(n14867), .A2(n14866), .ZN(n14868) );
  XOR2_X1 U18298 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n14868), .Z(
        n15050) );
  NOR2_X1 U18299 ( .A1(n20225), .A2(n21065), .ZN(n15047) );
  AOI21_X1 U18300 ( .B1(n20168), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15047), .ZN(n14869) );
  OAI21_X1 U18301 ( .B1(n20178), .B2(n14870), .A(n14869), .ZN(n14871) );
  AOI21_X1 U18302 ( .B1(n14872), .B2(n20239), .A(n14871), .ZN(n14873) );
  OAI21_X1 U18303 ( .B1(n20007), .B2(n15050), .A(n14873), .ZN(P1_U2971) );
  MUX2_X1 U18304 ( .A(n14875), .B(n14874), .S(n9672), .Z(n14876) );
  XNOR2_X1 U18305 ( .A(n14876), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15058) );
  INV_X1 U18306 ( .A(n14877), .ZN(n14879) );
  NOR2_X1 U18307 ( .A1(n20225), .A2(n21060), .ZN(n15051) );
  AOI21_X1 U18308 ( .B1(n20168), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15051), .ZN(n14878) );
  OAI21_X1 U18309 ( .B1(n20178), .B2(n14879), .A(n14878), .ZN(n14880) );
  AOI21_X1 U18310 ( .B1(n14881), .B2(n20239), .A(n14880), .ZN(n14882) );
  OAI21_X1 U18311 ( .B1(n20007), .B2(n15058), .A(n14882), .ZN(P1_U2972) );
  OAI21_X1 U18312 ( .B1(n12224), .B2(n14914), .A(n14883), .ZN(n14885) );
  NAND2_X1 U18313 ( .A1(n14885), .A2(n14884), .ZN(n14886) );
  XOR2_X1 U18314 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n14886), .Z(
        n15065) );
  NOR2_X1 U18315 ( .A1(n20225), .A2(n21019), .ZN(n15059) );
  AOI21_X1 U18316 ( .B1(n20168), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15059), .ZN(n14887) );
  OAI21_X1 U18317 ( .B1(n20178), .B2(n14888), .A(n14887), .ZN(n14889) );
  AOI21_X1 U18318 ( .B1(n14890), .B2(n20239), .A(n14889), .ZN(n14891) );
  OAI21_X1 U18319 ( .B1(n20007), .B2(n15065), .A(n14891), .ZN(P1_U2973) );
  NAND2_X1 U18320 ( .A1(n14892), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14903) );
  NAND2_X1 U18321 ( .A1(n14914), .A2(n15092), .ZN(n14893) );
  MUX2_X1 U18322 ( .A(n14893), .B(n14905), .S(n14972), .Z(n14894) );
  AOI21_X1 U18323 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14903), .A(
        n14894), .ZN(n14895) );
  XNOR2_X1 U18324 ( .A(n14895), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15073) );
  INV_X1 U18325 ( .A(n14896), .ZN(n14899) );
  INV_X1 U18326 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n14897) );
  NOR2_X1 U18327 ( .A1(n20225), .A2(n14897), .ZN(n15066) );
  AOI21_X1 U18328 ( .B1(n20168), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15066), .ZN(n14898) );
  OAI21_X1 U18329 ( .B1(n20178), .B2(n14899), .A(n14898), .ZN(n14900) );
  AOI21_X1 U18330 ( .B1(n14901), .B2(n20239), .A(n14900), .ZN(n14902) );
  OAI21_X1 U18331 ( .B1(n20007), .B2(n15073), .A(n14902), .ZN(P1_U2974) );
  NAND2_X1 U18332 ( .A1(n14914), .A2(n14903), .ZN(n14904) );
  MUX2_X1 U18333 ( .A(n14904), .B(n14903), .S(n14972), .Z(n14906) );
  XNOR2_X1 U18334 ( .A(n14906), .B(n14905), .ZN(n15084) );
  NOR2_X1 U18335 ( .A1(n20225), .A2(n14907), .ZN(n15074) );
  AOI21_X1 U18336 ( .B1(n20168), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15074), .ZN(n14908) );
  OAI21_X1 U18337 ( .B1(n20178), .B2(n14909), .A(n14908), .ZN(n14910) );
  AOI21_X1 U18338 ( .B1(n14911), .B2(n20239), .A(n14910), .ZN(n14912) );
  OAI21_X1 U18339 ( .B1(n20007), .B2(n15084), .A(n14912), .ZN(P1_U2975) );
  XNOR2_X1 U18340 ( .A(n9672), .B(n15092), .ZN(n14913) );
  XNOR2_X1 U18341 ( .A(n14914), .B(n14913), .ZN(n15089) );
  INV_X1 U18342 ( .A(n14915), .ZN(n14920) );
  INV_X1 U18343 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14916) );
  NOR2_X1 U18344 ( .A1(n20225), .A2(n14916), .ZN(n15085) );
  AOI21_X1 U18345 ( .B1(n20168), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15085), .ZN(n14917) );
  OAI21_X1 U18346 ( .B1(n20178), .B2(n14918), .A(n14917), .ZN(n14919) );
  AOI21_X1 U18347 ( .B1(n14920), .B2(n20239), .A(n14919), .ZN(n14921) );
  OAI21_X1 U18348 ( .B1(n15089), .B2(n20007), .A(n14921), .ZN(P1_U2976) );
  NAND2_X1 U18349 ( .A1(n14923), .A2(n14922), .ZN(n14924) );
  XOR2_X1 U18350 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n14924), .Z(
        n15112) );
  NOR2_X1 U18351 ( .A1(n20225), .A2(n21059), .ZN(n15108) );
  AOI21_X1 U18352 ( .B1(n20168), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15108), .ZN(n14925) );
  OAI21_X1 U18353 ( .B1(n20178), .B2(n14926), .A(n14925), .ZN(n14927) );
  AOI21_X1 U18354 ( .B1(n14928), .B2(n20239), .A(n14927), .ZN(n14929) );
  OAI21_X1 U18355 ( .B1(n20007), .B2(n15112), .A(n14929), .ZN(P1_U2977) );
  INV_X1 U18356 ( .A(n16082), .ZN(n14930) );
  NAND3_X1 U18357 ( .A1(n14930), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n9673), .ZN(n14939) );
  OAI22_X1 U18358 ( .A1(n14939), .A2(n15123), .B1(n14972), .B2(n14931), .ZN(
        n14932) );
  XNOR2_X1 U18359 ( .A(n14932), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15120) );
  INV_X1 U18360 ( .A(n14933), .ZN(n14935) );
  NOR2_X1 U18361 ( .A1(n20225), .A2(n20994), .ZN(n15115) );
  AOI21_X1 U18362 ( .B1(n20168), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15115), .ZN(n14934) );
  OAI21_X1 U18363 ( .B1(n20178), .B2(n14935), .A(n14934), .ZN(n14936) );
  AOI21_X1 U18364 ( .B1(n14937), .B2(n20239), .A(n14936), .ZN(n14938) );
  OAI21_X1 U18365 ( .B1(n15120), .B2(n20007), .A(n14938), .ZN(P1_U2978) );
  NOR2_X1 U18366 ( .A1(n14972), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14947) );
  NAND2_X1 U18367 ( .A1(n14947), .A2(n15138), .ZN(n14940) );
  OAI21_X1 U18368 ( .B1(n9671), .B2(n14940), .A(n14939), .ZN(n14941) );
  XNOR2_X1 U18369 ( .A(n14941), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15132) );
  INV_X1 U18370 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20985) );
  NOR2_X1 U18371 ( .A1(n20225), .A2(n20985), .ZN(n15128) );
  AOI21_X1 U18372 ( .B1(n20168), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15128), .ZN(n14942) );
  OAI21_X1 U18373 ( .B1(n20178), .B2(n14943), .A(n14942), .ZN(n14944) );
  AOI21_X1 U18374 ( .B1(n14945), .B2(n20239), .A(n14944), .ZN(n14946) );
  OAI21_X1 U18375 ( .B1(n15132), .B2(n20007), .A(n14946), .ZN(P1_U2979) );
  MUX2_X1 U18376 ( .A(n9673), .B(n14947), .S(n16082), .Z(n14948) );
  XNOR2_X1 U18377 ( .A(n14948), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15142) );
  INV_X1 U18378 ( .A(n14949), .ZN(n14955) );
  INV_X1 U18379 ( .A(n14950), .ZN(n14953) );
  NOR2_X1 U18380 ( .A1(n20225), .A2(n14951), .ZN(n15133) );
  AOI21_X1 U18381 ( .B1(n20168), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15133), .ZN(n14952) );
  OAI21_X1 U18382 ( .B1(n20178), .B2(n14953), .A(n14952), .ZN(n14954) );
  AOI21_X1 U18383 ( .B1(n14955), .B2(n20239), .A(n14954), .ZN(n14956) );
  OAI21_X1 U18384 ( .B1(n20007), .B2(n15142), .A(n14956), .ZN(P1_U2980) );
  NAND2_X1 U18385 ( .A1(n20168), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14957) );
  OAI21_X1 U18386 ( .B1(n14958), .B2(n20225), .A(n14957), .ZN(n14961) );
  NOR2_X1 U18387 ( .A1(n14959), .A2(n16049), .ZN(n14960) );
  AOI211_X1 U18388 ( .C1(n16044), .C2(n14962), .A(n14961), .B(n14960), .ZN(
        n14966) );
  OR2_X1 U18389 ( .A1(n9671), .A2(n14963), .ZN(n16083) );
  NAND3_X1 U18390 ( .A1(n16083), .A2(n16082), .A3(n20174), .ZN(n14965) );
  NAND2_X1 U18391 ( .A1(n14966), .A2(n14965), .ZN(P1_U2981) );
  NOR2_X1 U18392 ( .A1(n14972), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14971) );
  OAI21_X1 U18393 ( .B1(n14969), .B2(n14968), .A(n14967), .ZN(n14970) );
  MUX2_X1 U18394 ( .A(n14972), .B(n14971), .S(n14970), .Z(n14973) );
  XOR2_X1 U18395 ( .A(n14974), .B(n14973), .Z(n16093) );
  AOI22_X1 U18396 ( .A1(n20168), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20167), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n14975) );
  OAI21_X1 U18397 ( .B1(n20178), .B2(n14976), .A(n14975), .ZN(n14977) );
  AOI21_X1 U18398 ( .B1(n14978), .B2(n20239), .A(n14977), .ZN(n14979) );
  OAI21_X1 U18399 ( .B1(n16093), .B2(n20007), .A(n14979), .ZN(P1_U2982) );
  INV_X1 U18400 ( .A(n14980), .ZN(n14981) );
  NOR2_X1 U18401 ( .A1(n14982), .A2(n14981), .ZN(n14986) );
  NOR2_X1 U18402 ( .A1(n14984), .A2(n14983), .ZN(n14985) );
  XOR2_X1 U18403 ( .A(n14986), .B(n14985), .Z(n16101) );
  AOI22_X1 U18404 ( .A1(n20168), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20167), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n14987) );
  OAI21_X1 U18405 ( .B1(n20178), .B2(n14988), .A(n14987), .ZN(n14989) );
  AOI21_X1 U18406 ( .B1(n14990), .B2(n20239), .A(n14989), .ZN(n14991) );
  OAI21_X1 U18407 ( .B1(n16101), .B2(n20007), .A(n14991), .ZN(P1_U2984) );
  OAI21_X1 U18408 ( .B1(n14993), .B2(n16038), .A(n14992), .ZN(n14994) );
  XOR2_X1 U18409 ( .A(n14995), .B(n14994), .Z(n15153) );
  AOI22_X1 U18410 ( .A1(n20168), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n20167), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14996) );
  OAI21_X1 U18411 ( .B1(n20178), .B2(n14997), .A(n14996), .ZN(n14998) );
  AOI21_X1 U18412 ( .B1(n14999), .B2(n20239), .A(n14998), .ZN(n15000) );
  OAI21_X1 U18413 ( .B1(n15153), .B2(n20007), .A(n15000), .ZN(P1_U2986) );
  INV_X1 U18414 ( .A(n20220), .ZN(n15012) );
  INV_X1 U18415 ( .A(n20214), .ZN(n15001) );
  NAND2_X1 U18416 ( .A1(n15012), .A2(n15001), .ZN(n15004) );
  NAND2_X1 U18417 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n16092), .ZN(
        n16090) );
  NAND2_X1 U18418 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15002) );
  NOR2_X1 U18419 ( .A1(n16090), .A2(n15002), .ZN(n15101) );
  NAND2_X1 U18420 ( .A1(n16115), .A2(n15101), .ZN(n15003) );
  NAND2_X1 U18421 ( .A1(n15004), .A2(n15003), .ZN(n15137) );
  NAND2_X1 U18422 ( .A1(n15004), .A2(n15105), .ZN(n15005) );
  NAND2_X1 U18423 ( .A1(n15137), .A2(n15005), .ZN(n15116) );
  NAND2_X1 U18424 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15013) );
  AND2_X1 U18425 ( .A1(n20220), .A2(n15013), .ZN(n15006) );
  NOR2_X1 U18426 ( .A1(n15086), .A2(n20220), .ZN(n15009) );
  INV_X1 U18427 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15170) );
  NOR2_X1 U18428 ( .A1(n15009), .A2(n15170), .ZN(n15021) );
  INV_X1 U18429 ( .A(n15009), .ZN(n15010) );
  AND2_X1 U18430 ( .A1(n20209), .A2(n15092), .ZN(n15007) );
  OR2_X1 U18431 ( .A1(n15086), .A2(n15007), .ZN(n15076) );
  AND2_X1 U18432 ( .A1(n20220), .A2(n15061), .ZN(n15008) );
  NOR2_X1 U18433 ( .A1(n15076), .A2(n15008), .ZN(n15070) );
  AOI21_X1 U18434 ( .B1(n15070), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15009), .ZN(n15052) );
  AOI21_X1 U18435 ( .B1(n15011), .B2(n15010), .A(n15052), .ZN(n15038) );
  OAI211_X1 U18436 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15012), .A(
        n15038), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15027) );
  NOR2_X1 U18437 ( .A1(n15105), .A2(n15013), .ZN(n15014) );
  AND2_X1 U18438 ( .A1(n15101), .A2(n15014), .ZN(n15015) );
  NAND2_X1 U18439 ( .A1(n15016), .A2(n15015), .ZN(n15079) );
  INV_X1 U18440 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15017) );
  NOR3_X1 U18441 ( .A1(n15079), .A2(n15017), .A3(n15061), .ZN(n15043) );
  NAND3_X1 U18442 ( .A1(n15043), .A2(n15044), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15026) );
  NOR3_X1 U18443 ( .A1(n15026), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15018), .ZN(n15019) );
  AOI211_X1 U18444 ( .C1(n15021), .C2(n15027), .A(n15020), .B(n15019), .ZN(
        n15024) );
  NAND2_X1 U18445 ( .A1(n15022), .A2(n20228), .ZN(n15023) );
  INV_X1 U18446 ( .A(n15026), .ZN(n15028) );
  OAI21_X1 U18447 ( .B1(n15028), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n15027), .ZN(n15029) );
  OAI211_X1 U18448 ( .C1(n14517), .C2(n20182), .A(n15030), .B(n15029), .ZN(
        n15031) );
  AOI21_X1 U18449 ( .B1(n15032), .B2(n20206), .A(n15031), .ZN(n15033) );
  INV_X1 U18450 ( .A(n15033), .ZN(P1_U3001) );
  NAND3_X1 U18451 ( .A1(n15043), .A2(n15044), .A3(n15037), .ZN(n15036) );
  INV_X1 U18452 ( .A(n15034), .ZN(n15035) );
  OAI211_X1 U18453 ( .C1(n15038), .C2(n15037), .A(n15036), .B(n15035), .ZN(
        n15039) );
  AOI21_X1 U18454 ( .B1(n15040), .B2(n20228), .A(n15039), .ZN(n15041) );
  OAI21_X1 U18455 ( .B1(n15042), .B2(n20222), .A(n15041), .ZN(P1_U3002) );
  INV_X1 U18456 ( .A(n15043), .ZN(n15054) );
  NOR3_X1 U18457 ( .A1(n15054), .A2(n15045), .A3(n15044), .ZN(n15046) );
  AOI211_X1 U18458 ( .C1(n15052), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15047), .B(n15046), .ZN(n15049) );
  NAND2_X1 U18459 ( .A1(n10171), .A2(n20228), .ZN(n15048) );
  OAI211_X1 U18460 ( .C1(n15050), .C2(n20222), .A(n15049), .B(n15048), .ZN(
        P1_U3003) );
  AOI21_X1 U18461 ( .B1(n15052), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15051), .ZN(n15053) );
  OAI21_X1 U18462 ( .B1(n15054), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15053), .ZN(n15055) );
  AOI21_X1 U18463 ( .B1(n15056), .B2(n20228), .A(n15055), .ZN(n15057) );
  OAI21_X1 U18464 ( .B1(n15058), .B2(n20222), .A(n15057), .ZN(P1_U3004) );
  AOI21_X1 U18465 ( .B1(n15060), .B2(n20228), .A(n15059), .ZN(n15064) );
  INV_X1 U18466 ( .A(n15079), .ZN(n15093) );
  NAND2_X1 U18467 ( .A1(n15093), .A2(n9780), .ZN(n15062) );
  MUX2_X1 U18468 ( .A(n15062), .B(n15070), .S(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n15063) );
  OAI211_X1 U18469 ( .C1(n15065), .C2(n20222), .A(n15064), .B(n15063), .ZN(
        P1_U3005) );
  AOI21_X1 U18470 ( .B1(n15067), .B2(n20228), .A(n15066), .ZN(n15072) );
  NAND3_X1 U18471 ( .A1(n15093), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15069) );
  MUX2_X1 U18472 ( .A(n15070), .B(n15069), .S(n15068), .Z(n15071) );
  OAI211_X1 U18473 ( .C1(n15073), .C2(n20222), .A(n15072), .B(n15071), .ZN(
        P1_U3006) );
  AOI21_X1 U18474 ( .B1(n15075), .B2(n20228), .A(n15074), .ZN(n15083) );
  INV_X1 U18475 ( .A(n15076), .ZN(n15077) );
  OAI21_X1 U18476 ( .B1(n15078), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15077), .ZN(n15081) );
  NOR3_X1 U18477 ( .A1(n15079), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15092), .ZN(n15080) );
  AOI21_X1 U18478 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15081), .A(
        n15080), .ZN(n15082) );
  OAI211_X1 U18479 ( .C1(n15084), .C2(n20222), .A(n15083), .B(n15082), .ZN(
        P1_U3007) );
  AOI21_X1 U18480 ( .B1(n15086), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15085), .ZN(n15087) );
  OAI21_X1 U18481 ( .B1(n15088), .B2(n20182), .A(n15087), .ZN(n15091) );
  NOR2_X1 U18482 ( .A1(n15089), .A2(n20222), .ZN(n15090) );
  AOI211_X1 U18483 ( .C1(n15093), .C2(n15092), .A(n15091), .B(n15090), .ZN(
        n15094) );
  INV_X1 U18484 ( .A(n15094), .ZN(P1_U3008) );
  INV_X1 U18485 ( .A(n15095), .ZN(n15096) );
  NAND2_X1 U18486 ( .A1(n20209), .A2(n15096), .ZN(n15104) );
  NAND2_X1 U18487 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15145), .ZN(
        n15097) );
  OR2_X1 U18488 ( .A1(n15098), .A2(n15097), .ZN(n15099) );
  NAND2_X1 U18489 ( .A1(n15104), .A2(n15099), .ZN(n15144) );
  INV_X1 U18490 ( .A(n15100), .ZN(n15146) );
  OR2_X1 U18491 ( .A1(n15144), .A2(n15146), .ZN(n15122) );
  INV_X1 U18492 ( .A(n15145), .ZN(n15103) );
  NAND2_X1 U18493 ( .A1(n15101), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15102) );
  AOI21_X1 U18494 ( .B1(n15104), .B2(n15103), .A(n15102), .ZN(n15134) );
  NAND3_X1 U18495 ( .A1(n15122), .A2(n15134), .A3(n10044), .ZN(n15113) );
  XNOR2_X1 U18496 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15106) );
  NOR2_X1 U18497 ( .A1(n15113), .A2(n15106), .ZN(n15107) );
  AOI211_X1 U18498 ( .C1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n15116), .A(
        n15108), .B(n15107), .ZN(n15111) );
  NAND2_X1 U18499 ( .A1(n15109), .A2(n20228), .ZN(n15110) );
  OAI211_X1 U18500 ( .C1(n15112), .C2(n20222), .A(n15111), .B(n15110), .ZN(
        P1_U3009) );
  NOR2_X1 U18501 ( .A1(n15113), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15114) );
  AOI211_X1 U18502 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15116), .A(
        n15115), .B(n15114), .ZN(n15119) );
  NAND2_X1 U18503 ( .A1(n15117), .A2(n20228), .ZN(n15118) );
  OAI211_X1 U18504 ( .C1(n15120), .C2(n20222), .A(n15119), .B(n15118), .ZN(
        P1_U3010) );
  NOR2_X1 U18505 ( .A1(n15121), .A2(n20182), .ZN(n15130) );
  INV_X1 U18506 ( .A(n15122), .ZN(n15125) );
  NOR2_X1 U18507 ( .A1(n15125), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15135) );
  INV_X1 U18508 ( .A(n15135), .ZN(n15124) );
  AOI21_X1 U18509 ( .B1(n15124), .B2(n15137), .A(n15123), .ZN(n15129) );
  INV_X1 U18510 ( .A(n15134), .ZN(n15126) );
  NOR4_X1 U18511 ( .A1(n15126), .A2(n15125), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A4(n15138), .ZN(n15127) );
  NOR4_X1 U18512 ( .A1(n15130), .A2(n15129), .A3(n15128), .A4(n15127), .ZN(
        n15131) );
  OAI21_X1 U18513 ( .B1(n15132), .B2(n20222), .A(n15131), .ZN(P1_U3011) );
  AOI21_X1 U18514 ( .B1(n15135), .B2(n15134), .A(n15133), .ZN(n15136) );
  OAI21_X1 U18515 ( .B1(n15138), .B2(n15137), .A(n15136), .ZN(n15139) );
  AOI21_X1 U18516 ( .B1(n15140), .B2(n20228), .A(n15139), .ZN(n15141) );
  OAI21_X1 U18517 ( .B1(n15142), .B2(n20222), .A(n15141), .ZN(P1_U3012) );
  INV_X1 U18518 ( .A(n15143), .ZN(n15151) );
  NOR2_X1 U18519 ( .A1(n16115), .A2(n12230), .ZN(n15150) );
  AOI21_X1 U18520 ( .B1(n15146), .B2(n15145), .A(n15144), .ZN(n15148) );
  NAND2_X1 U18521 ( .A1(n20167), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15147) );
  OAI21_X1 U18522 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15148), .A(
        n15147), .ZN(n15149) );
  AOI211_X1 U18523 ( .C1(n15151), .C2(n20228), .A(n15150), .B(n15149), .ZN(
        n15152) );
  OAI21_X1 U18524 ( .B1(n15153), .B2(n20222), .A(n15152), .ZN(P1_U3018) );
  INV_X1 U18525 ( .A(n20622), .ZN(n20618) );
  INV_X1 U18526 ( .A(n20777), .ZN(n20368) );
  AND3_X1 U18527 ( .A1(n20490), .A2(n20783), .A3(n20368), .ZN(n20497) );
  INV_X1 U18528 ( .A(n20548), .ZN(n15157) );
  AND3_X1 U18529 ( .A1(n20720), .A2(n20783), .A3(n15157), .ZN(n20696) );
  NOR2_X1 U18530 ( .A1(n20497), .A2(n20696), .ZN(n15161) );
  INV_X1 U18531 ( .A(n15154), .ZN(n15159) );
  NOR2_X1 U18532 ( .A1(n20781), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20328) );
  AOI22_X1 U18533 ( .A1(n15159), .A2(n20328), .B1(n15158), .B2(n13423), .ZN(
        n15160) );
  OAI211_X1 U18534 ( .C1(n20781), .C2(n20618), .A(n15161), .B(n15160), .ZN(
        n15162) );
  MUX2_X1 U18535 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n15162), .S(
        n20235), .Z(P1_U3475) );
  NOR2_X1 U18536 ( .A1(n10190), .A2(n15163), .ZN(n15165) );
  INV_X1 U18537 ( .A(n15165), .ZN(n15172) );
  AOI22_X1 U18538 ( .A1(n15166), .A2(n10183), .B1(n15165), .B2(n15164), .ZN(
        n15167) );
  OAI21_X1 U18539 ( .B1(n20651), .B2(n15168), .A(n15167), .ZN(n15940) );
  NOR2_X1 U18540 ( .A1(n16181), .A2(n15169), .ZN(n15178) );
  OAI22_X1 U18541 ( .A1(n15170), .A2(n20233), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15176) );
  AOI22_X1 U18542 ( .A1(n15940), .A2(n16172), .B1(n15178), .B2(n15176), .ZN(
        n15171) );
  OAI21_X1 U18543 ( .B1(n15187), .B2(n15172), .A(n15171), .ZN(n15174) );
  INV_X1 U18544 ( .A(n15173), .ZN(n16176) );
  MUX2_X1 U18545 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15174), .S(
        n16176), .Z(P1_U3473) );
  INV_X1 U18546 ( .A(n15175), .ZN(n15181) );
  INV_X1 U18547 ( .A(n15176), .ZN(n15177) );
  AOI22_X1 U18548 ( .A1(n15179), .A2(n16172), .B1(n15178), .B2(n15177), .ZN(
        n15180) );
  OAI21_X1 U18549 ( .B1(n15187), .B2(n15181), .A(n15180), .ZN(n15182) );
  MUX2_X1 U18550 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n15182), .S(
        n16176), .Z(P1_U3472) );
  INV_X1 U18551 ( .A(n15183), .ZN(n15186) );
  OAI22_X1 U18552 ( .A1(n15187), .A2(n15186), .B1(n15185), .B2(n15184), .ZN(
        n15188) );
  MUX2_X1 U18553 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15188), .S(
        n16176), .Z(P1_U3469) );
  NAND2_X1 U18554 ( .A1(n15190), .A2(n15189), .ZN(n15191) );
  NAND2_X1 U18555 ( .A1(n9716), .A2(n15191), .ZN(n15574) );
  INV_X1 U18556 ( .A(n15193), .ZN(n15194) );
  AOI211_X1 U18557 ( .C1(n15195), .C2(n15192), .A(n15194), .B(n19851), .ZN(
        n15196) );
  INV_X1 U18558 ( .A(n15196), .ZN(n15202) );
  NAND2_X1 U18559 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n19135), .ZN(n15198) );
  AOI22_X1 U18560 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19142), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19076), .ZN(n15197) );
  OAI211_X1 U18561 ( .C1(n15199), .C2(n19101), .A(n15198), .B(n15197), .ZN(
        n15200) );
  AOI21_X1 U18562 ( .B1(n15567), .B2(n19122), .A(n15200), .ZN(n15201) );
  OAI211_X1 U18563 ( .C1(n15574), .C2(n19127), .A(n15202), .B(n15201), .ZN(
        P2_U2827) );
  AND2_X1 U18564 ( .A1(n15356), .A2(n15203), .ZN(n15204) );
  OR2_X1 U18565 ( .A1(n15204), .A2(n15337), .ZN(n15604) );
  AOI211_X1 U18566 ( .C1(n15205), .C2(n15425), .A(n15206), .B(n19851), .ZN(
        n15207) );
  INV_X1 U18567 ( .A(n15207), .ZN(n15218) );
  XOR2_X1 U18568 ( .A(P2_EBX_REG_25__SCAN_IN), .B(n15208), .Z(n15216) );
  OR2_X1 U18569 ( .A1(n15210), .A2(n15211), .ZN(n15212) );
  NAND2_X1 U18570 ( .A1(n15209), .A2(n15212), .ZN(n15603) );
  AOI22_X1 U18571 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19142), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19076), .ZN(n15214) );
  NAND2_X1 U18572 ( .A1(n19135), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n15213) );
  OAI211_X1 U18573 ( .C1(n15603), .C2(n19137), .A(n15214), .B(n15213), .ZN(
        n15215) );
  AOI21_X1 U18574 ( .B1(n15216), .B2(n19131), .A(n15215), .ZN(n15217) );
  OAI211_X1 U18575 ( .C1(n15604), .C2(n19127), .A(n15218), .B(n15217), .ZN(
        P2_U2830) );
  NOR2_X1 U18576 ( .A1(n15220), .A2(n15219), .ZN(n15221) );
  OR2_X1 U18577 ( .A1(n13990), .A2(n15221), .ZN(n16238) );
  INV_X1 U18578 ( .A(n16238), .ZN(n15231) );
  AOI22_X1 U18579 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(n19135), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19142), .ZN(n15222) );
  OAI211_X1 U18580 ( .C1(n19133), .C2(n15223), .A(n15222), .B(n19113), .ZN(
        n15224) );
  AOI21_X1 U18581 ( .B1(n15225), .B2(n19122), .A(n15224), .ZN(n15226) );
  OAI21_X1 U18582 ( .B1(n15227), .B2(n19101), .A(n15226), .ZN(n15230) );
  AOI211_X1 U18583 ( .C1(n15512), .C2(n9994), .A(n15228), .B(n19851), .ZN(
        n15229) );
  AOI211_X1 U18584 ( .C1(n19129), .C2(n15231), .A(n15230), .B(n15229), .ZN(
        n15232) );
  INV_X1 U18585 ( .A(n15232), .ZN(P2_U2837) );
  NAND2_X1 U18586 ( .A1(n16186), .A2(n15305), .ZN(n15233) );
  OAI21_X1 U18587 ( .B1(n15302), .B2(n15234), .A(n15233), .ZN(P2_U2856) );
  OR2_X1 U18588 ( .A1(n15236), .A2(n15235), .ZN(n15314) );
  NAND3_X1 U18589 ( .A1(n15314), .A2(n15237), .A3(n15298), .ZN(n15239) );
  NAND2_X1 U18590 ( .A1(n15269), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15238) );
  OAI211_X1 U18591 ( .C1(n15269), .C2(n16199), .A(n15239), .B(n15238), .ZN(
        P2_U2858) );
  NAND2_X1 U18592 ( .A1(n10126), .A2(n15240), .ZN(n15242) );
  XNOR2_X1 U18593 ( .A(n15242), .B(n15241), .ZN(n15326) );
  NAND2_X1 U18594 ( .A1(n15269), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15244) );
  NAND2_X1 U18595 ( .A1(n15567), .A2(n15302), .ZN(n15243) );
  OAI211_X1 U18596 ( .C1(n15326), .C2(n15312), .A(n15244), .B(n15243), .ZN(
        P2_U2859) );
  OAI21_X1 U18597 ( .B1(n15247), .B2(n15246), .A(n15245), .ZN(n15333) );
  NAND2_X1 U18598 ( .A1(n15269), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15249) );
  NAND2_X1 U18599 ( .A1(n15404), .A2(n15302), .ZN(n15248) );
  OAI211_X1 U18600 ( .C1(n15333), .C2(n15312), .A(n15249), .B(n15248), .ZN(
        P2_U2860) );
  INV_X1 U18601 ( .A(n12883), .ZN(n15250) );
  AOI21_X1 U18602 ( .B1(n15251), .B2(n15209), .A(n15250), .ZN(n16207) );
  INV_X1 U18603 ( .A(n16207), .ZN(n15592) );
  AOI21_X1 U18604 ( .B1(n15254), .B2(n15253), .A(n15252), .ZN(n15338) );
  NAND2_X1 U18605 ( .A1(n15338), .A2(n15298), .ZN(n15256) );
  NAND2_X1 U18606 ( .A1(n15269), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15255) );
  OAI211_X1 U18607 ( .C1(n15592), .C2(n15269), .A(n15256), .B(n15255), .ZN(
        P2_U2861) );
  OAI21_X1 U18608 ( .B1(n15259), .B2(n15258), .A(n15257), .ZN(n15350) );
  NOR2_X1 U18609 ( .A1(n15603), .A2(n15309), .ZN(n15260) );
  AOI21_X1 U18610 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n15269), .A(n15260), .ZN(
        n15261) );
  OAI21_X1 U18611 ( .B1(n15350), .B2(n15312), .A(n15261), .ZN(P2_U2862) );
  AOI21_X1 U18612 ( .B1(n15263), .B2(n15262), .A(n9715), .ZN(n15264) );
  XOR2_X1 U18613 ( .A(n15265), .B(n15264), .Z(n15360) );
  NOR2_X1 U18614 ( .A1(n15267), .A2(n15266), .ZN(n15268) );
  OR2_X1 U18615 ( .A1(n15210), .A2(n15268), .ZN(n16218) );
  MUX2_X1 U18616 ( .A(n16218), .B(n15270), .S(n15269), .Z(n15271) );
  OAI21_X1 U18617 ( .B1(n15360), .B2(n15312), .A(n15271), .ZN(P2_U2863) );
  NOR2_X1 U18618 ( .A1(n15273), .A2(n15272), .ZN(n15275) );
  NOR2_X1 U18619 ( .A1(n15275), .A2(n15274), .ZN(n15365) );
  NAND2_X1 U18620 ( .A1(n15365), .A2(n15298), .ZN(n15278) );
  INV_X1 U18621 ( .A(n15629), .ZN(n15276) );
  NAND2_X1 U18622 ( .A1(n15276), .A2(n15302), .ZN(n15277) );
  OAI211_X1 U18623 ( .C1(n15302), .C2(n15279), .A(n15278), .B(n15277), .ZN(
        P2_U2864) );
  NAND2_X1 U18624 ( .A1(n15287), .A2(n15280), .ZN(n15288) );
  INV_X1 U18625 ( .A(n15288), .ZN(n15282) );
  OAI21_X1 U18626 ( .B1(n15282), .B2(n15281), .A(n14317), .ZN(n15377) );
  NOR2_X1 U18627 ( .A1(n15283), .A2(n15309), .ZN(n15284) );
  AOI21_X1 U18628 ( .B1(P2_EBX_REG_22__SCAN_IN), .B2(n15269), .A(n15284), .ZN(
        n15285) );
  OAI21_X1 U18629 ( .B1(n15377), .B2(n15312), .A(n15285), .ZN(P2_U2865) );
  AND2_X1 U18630 ( .A1(n15287), .A2(n15286), .ZN(n15297) );
  OAI21_X1 U18631 ( .B1(n15297), .B2(n15289), .A(n15288), .ZN(n15387) );
  OAI21_X1 U18632 ( .B1(n15301), .B2(n15290), .A(n9736), .ZN(n15658) );
  NOR2_X1 U18633 ( .A1(n15658), .A2(n15309), .ZN(n15291) );
  AOI21_X1 U18634 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n15269), .A(n15291), .ZN(
        n15292) );
  OAI21_X1 U18635 ( .B1(n15387), .B2(n15312), .A(n15292), .ZN(P2_U2866) );
  INV_X1 U18636 ( .A(n15293), .ZN(n15294) );
  AND2_X1 U18637 ( .A1(n15295), .A2(n15294), .ZN(n15296) );
  NOR2_X1 U18638 ( .A1(n15297), .A2(n15296), .ZN(n16230) );
  NAND2_X1 U18639 ( .A1(n16230), .A2(n15298), .ZN(n15304) );
  NOR2_X1 U18640 ( .A1(n15307), .A2(n15299), .ZN(n15300) );
  OR2_X1 U18641 ( .A1(n15301), .A2(n15300), .ZN(n18988) );
  NAND2_X1 U18642 ( .A1(n15670), .A2(n15302), .ZN(n15303) );
  OAI211_X1 U18643 ( .C1(n15305), .C2(n11740), .A(n15304), .B(n15303), .ZN(
        P2_U2867) );
  AND2_X1 U18644 ( .A1(n9694), .A2(n15306), .ZN(n15308) );
  OR2_X1 U18645 ( .A1(n15308), .A2(n15307), .ZN(n15497) );
  NOR2_X1 U18646 ( .A1(n15497), .A2(n15309), .ZN(n15310) );
  AOI21_X1 U18647 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n15269), .A(n15310), .ZN(
        n15311) );
  OAI21_X1 U18648 ( .B1(n15313), .B2(n15312), .A(n15311), .ZN(P2_U2868) );
  INV_X1 U18649 ( .A(n19183), .ZN(n19191) );
  NAND3_X1 U18650 ( .A1(n15314), .A2(n15237), .A3(n19191), .ZN(n15320) );
  INV_X1 U18651 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n15317) );
  AOI22_X1 U18652 ( .A1(n16235), .A2(n15315), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n19188), .ZN(n15316) );
  OAI21_X1 U18653 ( .B1(n15346), .B2(n15317), .A(n15316), .ZN(n15318) );
  AOI21_X1 U18654 ( .B1(n19147), .B2(BUF2_REG_29__SCAN_IN), .A(n15318), .ZN(
        n15319) );
  OAI211_X1 U18655 ( .C1(n16237), .C2(n16203), .A(n15320), .B(n15319), .ZN(
        P2_U2890) );
  INV_X1 U18656 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n15322) );
  AOI22_X1 U18657 ( .A1(n16235), .A2(n19155), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n19188), .ZN(n15321) );
  OAI21_X1 U18658 ( .B1(n15346), .B2(n15322), .A(n15321), .ZN(n15324) );
  NOR2_X1 U18659 ( .A1(n15574), .A2(n16237), .ZN(n15323) );
  AOI211_X1 U18660 ( .C1(n19147), .C2(BUF2_REG_28__SCAN_IN), .A(n15324), .B(
        n15323), .ZN(n15325) );
  OAI21_X1 U18661 ( .B1(n15326), .B2(n19183), .A(n15325), .ZN(P2_U2891) );
  INV_X1 U18662 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n15329) );
  AOI22_X1 U18663 ( .A1(n16235), .A2(n15327), .B1(P2_EAX_REG_27__SCAN_IN), 
        .B2(n19188), .ZN(n15328) );
  OAI21_X1 U18664 ( .B1(n15346), .B2(n15329), .A(n15328), .ZN(n15331) );
  NOR2_X1 U18665 ( .A1(n15586), .A2(n16237), .ZN(n15330) );
  AOI211_X1 U18666 ( .C1(n19147), .C2(BUF2_REG_27__SCAN_IN), .A(n15331), .B(
        n15330), .ZN(n15332) );
  OAI21_X1 U18667 ( .B1(n15333), .B2(n19183), .A(n15332), .ZN(P2_U2892) );
  INV_X1 U18668 ( .A(n15334), .ZN(n15335) );
  OAI21_X1 U18669 ( .B1(n15337), .B2(n15336), .A(n15335), .ZN(n16206) );
  NAND2_X1 U18670 ( .A1(n15338), .A2(n19191), .ZN(n15342) );
  AOI22_X1 U18671 ( .A1(n16235), .A2(n19159), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n19188), .ZN(n15339) );
  OAI21_X1 U18672 ( .B1(n15346), .B2(n20262), .A(n15339), .ZN(n15340) );
  AOI21_X1 U18673 ( .B1(n19147), .B2(BUF2_REG_26__SCAN_IN), .A(n15340), .ZN(
        n15341) );
  OAI211_X1 U18674 ( .C1(n16206), .C2(n16237), .A(n15342), .B(n15341), .ZN(
        P2_U2893) );
  INV_X1 U18675 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n15345) );
  AOI22_X1 U18676 ( .A1(n16235), .A2(n15343), .B1(P2_EAX_REG_25__SCAN_IN), 
        .B2(n19188), .ZN(n15344) );
  OAI21_X1 U18677 ( .B1(n15346), .B2(n15345), .A(n15344), .ZN(n15348) );
  NOR2_X1 U18678 ( .A1(n15604), .A2(n16237), .ZN(n15347) );
  AOI211_X1 U18679 ( .C1(n19147), .C2(BUF2_REG_25__SCAN_IN), .A(n15348), .B(
        n15347), .ZN(n15349) );
  OAI21_X1 U18680 ( .B1(n19183), .B2(n15350), .A(n15349), .ZN(P2_U2894) );
  NAND2_X1 U18681 ( .A1(n19149), .A2(BUF1_REG_24__SCAN_IN), .ZN(n15352) );
  AOI22_X1 U18682 ( .A1(n16235), .A2(n19163), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n19188), .ZN(n15351) );
  NAND2_X1 U18683 ( .A1(n15352), .A2(n15351), .ZN(n15358) );
  NAND2_X1 U18684 ( .A1(n15354), .A2(n15353), .ZN(n15355) );
  NAND2_X1 U18685 ( .A1(n15356), .A2(n15355), .ZN(n16219) );
  NOR2_X1 U18686 ( .A1(n16219), .A2(n16237), .ZN(n15357) );
  AOI211_X1 U18687 ( .C1(n19147), .C2(BUF2_REG_24__SCAN_IN), .A(n15358), .B(
        n15357), .ZN(n15359) );
  OAI21_X1 U18688 ( .B1(n15360), .B2(n19183), .A(n15359), .ZN(P2_U2895) );
  OAI22_X1 U18689 ( .A1(n19290), .A2(n15381), .B1(n15380), .B2(n15361), .ZN(
        n15364) );
  INV_X1 U18690 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n15362) );
  NOR2_X1 U18691 ( .A1(n15384), .A2(n15362), .ZN(n15363) );
  AOI211_X1 U18692 ( .C1(BUF1_REG_23__SCAN_IN), .C2(n19149), .A(n15364), .B(
        n15363), .ZN(n15367) );
  NAND2_X1 U18693 ( .A1(n15365), .A2(n19191), .ZN(n15366) );
  OAI211_X1 U18694 ( .C1(n15368), .C2(n16237), .A(n15367), .B(n15366), .ZN(
        P2_U2896) );
  NAND2_X1 U18695 ( .A1(n19149), .A2(BUF1_REG_22__SCAN_IN), .ZN(n15371) );
  INV_X1 U18696 ( .A(n19280), .ZN(n15369) );
  NAND2_X1 U18697 ( .A1(n16235), .A2(n15369), .ZN(n15370) );
  OAI211_X1 U18698 ( .C1(n15380), .C2(n15372), .A(n15371), .B(n15370), .ZN(
        n15375) );
  NOR2_X1 U18699 ( .A1(n15373), .A2(n16237), .ZN(n15374) );
  AOI211_X1 U18700 ( .C1(n19147), .C2(BUF2_REG_22__SCAN_IN), .A(n15375), .B(
        n15374), .ZN(n15376) );
  OAI21_X1 U18701 ( .B1(n19183), .B2(n15377), .A(n15376), .ZN(P2_U2897) );
  XOR2_X1 U18702 ( .A(n15378), .B(n15667), .Z(n18984) );
  OAI22_X1 U18703 ( .A1(n19276), .A2(n15381), .B1(n15380), .B2(n15379), .ZN(
        n15382) );
  AOI21_X1 U18704 ( .B1(n19149), .B2(BUF1_REG_21__SCAN_IN), .A(n15382), .ZN(
        n15383) );
  OAI21_X1 U18705 ( .B1(n15384), .B2(n18284), .A(n15383), .ZN(n15385) );
  AOI21_X1 U18706 ( .B1(n18984), .B2(n19189), .A(n15385), .ZN(n15386) );
  OAI21_X1 U18707 ( .B1(n19183), .B2(n15387), .A(n15386), .ZN(P2_U2898) );
  OAI21_X1 U18708 ( .B1(n16310), .B2(n15389), .A(n15388), .ZN(n15390) );
  AOI21_X1 U18709 ( .B1(n16301), .B2(n10160), .A(n15390), .ZN(n15391) );
  OAI21_X1 U18710 ( .B1(n16199), .B2(n13736), .A(n15391), .ZN(n15392) );
  AOI21_X1 U18711 ( .B1(n15393), .B2(n19236), .A(n15392), .ZN(n15394) );
  OAI21_X1 U18712 ( .B1(n15395), .B2(n11993), .A(n15394), .ZN(P2_U2985) );
  XNOR2_X1 U18713 ( .A(n15396), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15590) );
  NAND2_X1 U18714 ( .A1(n16301), .A2(n15397), .ZN(n15398) );
  NAND2_X1 U18715 ( .A1(n15544), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15580) );
  OAI211_X1 U18716 ( .C1(n16310), .C2(n15399), .A(n15398), .B(n15580), .ZN(
        n15403) );
  INV_X1 U18717 ( .A(n15400), .ZN(n15401) );
  NOR2_X1 U18718 ( .A1(n15579), .A2(n16303), .ZN(n15402) );
  OAI21_X1 U18719 ( .B1(n15590), .B2(n11993), .A(n15405), .ZN(P2_U2987) );
  NAND2_X1 U18720 ( .A1(n15406), .A2(n15418), .ZN(n15407) );
  XOR2_X1 U18721 ( .A(n15408), .B(n15407), .Z(n15600) );
  NAND2_X1 U18722 ( .A1(n15544), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15591) );
  NAND2_X1 U18723 ( .A1(n19231), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15409) );
  OAI211_X1 U18724 ( .C1(n19240), .C2(n15410), .A(n15591), .B(n15409), .ZN(
        n15411) );
  AOI21_X1 U18725 ( .B1(n16207), .B2(n16306), .A(n15411), .ZN(n15416) );
  AOI21_X1 U18726 ( .B1(n15414), .B2(n15412), .A(n15413), .ZN(n15598) );
  NAND2_X1 U18727 ( .A1(n15598), .A2(n19236), .ZN(n15415) );
  OAI211_X1 U18728 ( .C1(n15600), .C2(n11993), .A(n15416), .B(n15415), .ZN(
        P2_U2988) );
  INV_X1 U18729 ( .A(n15418), .ZN(n15421) );
  AND2_X1 U18730 ( .A1(n15418), .A2(n15417), .ZN(n15419) );
  OAI22_X1 U18731 ( .A1(n15406), .A2(n15421), .B1(n15420), .B2(n15419), .ZN(
        n15612) );
  NAND2_X1 U18732 ( .A1(n15544), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15602) );
  OAI21_X1 U18733 ( .B1(n16310), .B2(n15422), .A(n15602), .ZN(n15424) );
  NOR2_X1 U18734 ( .A1(n15603), .A2(n13736), .ZN(n15423) );
  AOI211_X1 U18735 ( .C1(n16301), .C2(n15425), .A(n15424), .B(n15423), .ZN(
        n15428) );
  NAND2_X1 U18736 ( .A1(n15426), .A2(n15607), .ZN(n15609) );
  NAND3_X1 U18737 ( .A1(n15412), .A2(n19236), .A3(n15609), .ZN(n15427) );
  OAI211_X1 U18738 ( .C1(n15612), .C2(n11993), .A(n15428), .B(n15427), .ZN(
        P2_U2989) );
  XNOR2_X1 U18739 ( .A(n15429), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15430) );
  XNOR2_X1 U18740 ( .A(n15431), .B(n15430), .ZN(n15625) );
  INV_X1 U18741 ( .A(n16218), .ZN(n15437) );
  NAND2_X1 U18742 ( .A1(n16301), .A2(n16223), .ZN(n15432) );
  NAND2_X1 U18743 ( .A1(n15544), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15617) );
  OAI211_X1 U18744 ( .C1(n16310), .C2(n15433), .A(n15432), .B(n15617), .ZN(
        n15436) );
  OAI21_X1 U18745 ( .B1(n15434), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15426), .ZN(n15613) );
  NOR2_X1 U18746 ( .A1(n15613), .A2(n16303), .ZN(n15435) );
  AOI211_X1 U18747 ( .C1(n16306), .C2(n15437), .A(n15436), .B(n15435), .ZN(
        n15438) );
  OAI21_X1 U18748 ( .B1(n15625), .B2(n11993), .A(n15438), .ZN(P2_U2990) );
  XNOR2_X1 U18749 ( .A(n9640), .B(n15439), .ZN(n15639) );
  NAND2_X1 U18750 ( .A1(n15544), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15628) );
  OAI21_X1 U18751 ( .B1(n16310), .B2(n15441), .A(n15628), .ZN(n15443) );
  NOR2_X1 U18752 ( .A1(n15629), .A2(n13736), .ZN(n15442) );
  AOI211_X1 U18753 ( .C1(n16301), .C2(n15444), .A(n15443), .B(n15442), .ZN(
        n15447) );
  AOI21_X1 U18754 ( .B1(n15633), .B2(n15445), .A(n15434), .ZN(n15636) );
  NAND2_X1 U18755 ( .A1(n15636), .A2(n19236), .ZN(n15446) );
  OAI211_X1 U18756 ( .C1(n15639), .C2(n11993), .A(n15447), .B(n15446), .ZN(
        P2_U2991) );
  OAI21_X1 U18757 ( .B1(n10037), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15445), .ZN(n15652) );
  INV_X1 U18758 ( .A(n15449), .ZN(n15450) );
  NOR2_X1 U18759 ( .A1(n15451), .A2(n15450), .ZN(n15452) );
  XNOR2_X1 U18760 ( .A(n15453), .B(n15452), .ZN(n15650) );
  NAND2_X1 U18761 ( .A1(n15645), .A2(n16306), .ZN(n15455) );
  NOR2_X1 U18762 ( .A1(n19113), .A2(n19900), .ZN(n15644) );
  AOI21_X1 U18763 ( .B1(n19231), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15644), .ZN(n15454) );
  OAI211_X1 U18764 ( .C1(n19240), .C2(n15456), .A(n15455), .B(n15454), .ZN(
        n15457) );
  AOI21_X1 U18765 ( .B1(n15650), .B2(n16297), .A(n15457), .ZN(n15458) );
  OAI21_X1 U18766 ( .B1(n16303), .B2(n15652), .A(n15458), .ZN(P2_U2992) );
  NOR2_X1 U18767 ( .A1(n15460), .A2(n15459), .ZN(n15780) );
  NOR3_X1 U18768 ( .A1(n19064), .A2(n15461), .A3(n11704), .ZN(n15779) );
  INV_X1 U18769 ( .A(n15761), .ZN(n15462) );
  INV_X1 U18770 ( .A(n15463), .ZN(n15742) );
  INV_X1 U18771 ( .A(n15464), .ZN(n15465) );
  NAND2_X1 U18772 ( .A1(n9953), .A2(n15468), .ZN(n15469) );
  XNOR2_X1 U18773 ( .A(n15470), .B(n15469), .ZN(n15663) );
  INV_X1 U18774 ( .A(n15658), .ZN(n18979) );
  NAND2_X1 U18775 ( .A1(n16301), .A2(n18982), .ZN(n15471) );
  NAND2_X1 U18776 ( .A1(n15544), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15656) );
  OAI211_X1 U18777 ( .C1(n16310), .C2(n11846), .A(n15471), .B(n15656), .ZN(
        n15476) );
  NAND2_X1 U18778 ( .A1(n15472), .A2(n15473), .ZN(n15474) );
  NAND2_X1 U18779 ( .A1(n15448), .A2(n15474), .ZN(n15659) );
  NOR2_X1 U18780 ( .A1(n15659), .A2(n16303), .ZN(n15475) );
  AOI211_X1 U18781 ( .C1(n18979), .C2(n16306), .A(n15476), .B(n15475), .ZN(
        n15477) );
  OAI21_X1 U18782 ( .B1(n15663), .B2(n11993), .A(n15477), .ZN(P2_U2993) );
  NAND2_X1 U18783 ( .A1(n15479), .A2(n15478), .ZN(n15484) );
  INV_X1 U18784 ( .A(n15480), .ZN(n15482) );
  NAND2_X1 U18785 ( .A1(n15482), .A2(n15481), .ZN(n15483) );
  XNOR2_X1 U18786 ( .A(n15484), .B(n15483), .ZN(n15678) );
  NOR2_X1 U18787 ( .A1(n19113), .A2(n15485), .ZN(n15669) );
  AOI21_X1 U18788 ( .B1(n19231), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15669), .ZN(n15486) );
  OAI21_X1 U18789 ( .B1(n19240), .B2(n15487), .A(n15486), .ZN(n15490) );
  OAI21_X1 U18790 ( .B1(n15680), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15472), .ZN(n15674) );
  NOR2_X1 U18791 ( .A1(n15674), .A2(n16303), .ZN(n15489) );
  AOI211_X1 U18792 ( .C1(n16306), .C2(n15670), .A(n15490), .B(n15489), .ZN(
        n15491) );
  OAI21_X1 U18793 ( .B1(n15678), .B2(n11993), .A(n15491), .ZN(P2_U2994) );
  NAND2_X1 U18794 ( .A1(n9733), .A2(n15492), .ZN(n15496) );
  INV_X1 U18795 ( .A(n15493), .ZN(n15506) );
  XOR2_X1 U18796 ( .A(n15496), .B(n15495), .Z(n15690) );
  NAND2_X1 U18797 ( .A1(n16301), .A2(n19001), .ZN(n15498) );
  NAND2_X1 U18798 ( .A1(n15544), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15682) );
  OAI211_X1 U18799 ( .C1(n16310), .C2(n15499), .A(n15498), .B(n15682), .ZN(
        n15503) );
  NOR2_X1 U18800 ( .A1(n15500), .A2(n15501), .ZN(n15509) );
  NOR2_X1 U18801 ( .A1(n15509), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15679) );
  NOR3_X1 U18802 ( .A1(n15679), .A2(n15680), .A3(n16303), .ZN(n15502) );
  AOI211_X1 U18803 ( .C1(n16306), .C2(n19004), .A(n15503), .B(n15502), .ZN(
        n15504) );
  OAI21_X1 U18804 ( .B1(n15690), .B2(n11993), .A(n15504), .ZN(P2_U2995) );
  NOR2_X1 U18805 ( .A1(n15506), .A2(n15505), .ZN(n15507) );
  XNOR2_X1 U18806 ( .A(n15519), .B(n15507), .ZN(n15704) );
  OR2_X1 U18807 ( .A1(n15500), .A2(n15508), .ZN(n15510) );
  AOI21_X1 U18808 ( .B1(n15696), .B2(n15510), .A(n15509), .ZN(n15702) );
  NAND2_X1 U18809 ( .A1(n15544), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n15692) );
  OAI21_X1 U18810 ( .B1(n16310), .B2(n11844), .A(n15692), .ZN(n15511) );
  AOI21_X1 U18811 ( .B1(n16301), .B2(n15512), .A(n15511), .ZN(n15513) );
  OAI21_X1 U18812 ( .B1(n15693), .B2(n13736), .A(n15513), .ZN(n15514) );
  AOI21_X1 U18813 ( .B1(n15702), .B2(n19236), .A(n15514), .ZN(n15515) );
  OAI21_X1 U18814 ( .B1(n15704), .B2(n11993), .A(n15515), .ZN(P2_U2996) );
  OAI22_X1 U18815 ( .A1(n15519), .A2(n15518), .B1(n15517), .B2(n15516), .ZN(
        n15520) );
  INV_X1 U18816 ( .A(n15520), .ZN(n15718) );
  XNOR2_X1 U18817 ( .A(n15500), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15525) );
  NAND2_X1 U18818 ( .A1(n15544), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15711) );
  OAI21_X1 U18819 ( .B1(n16310), .B2(n15521), .A(n15711), .ZN(n15522) );
  AOI21_X1 U18820 ( .B1(n16301), .B2(n19017), .A(n15522), .ZN(n15523) );
  OAI21_X1 U18821 ( .B1(n19015), .B2(n13736), .A(n15523), .ZN(n15524) );
  AOI21_X1 U18822 ( .B1(n15525), .B2(n19236), .A(n15524), .ZN(n15526) );
  OAI21_X1 U18823 ( .B1(n15718), .B2(n11993), .A(n15526), .ZN(P2_U2997) );
  XOR2_X1 U18824 ( .A(n15528), .B(n15527), .Z(n15719) );
  INV_X1 U18825 ( .A(n15719), .ZN(n15537) );
  INV_X1 U18826 ( .A(n19030), .ZN(n15531) );
  NAND2_X1 U18827 ( .A1(n15544), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15720) );
  NAND2_X1 U18828 ( .A1(n19231), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15529) );
  OAI211_X1 U18829 ( .C1(n19240), .C2(n19029), .A(n15720), .B(n15529), .ZN(
        n15530) );
  AOI21_X1 U18830 ( .B1(n15531), .B2(n16306), .A(n15530), .ZN(n15536) );
  OAI211_X1 U18831 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15542), .A(
        n15500), .B(n19236), .ZN(n15535) );
  OAI211_X1 U18832 ( .C1(n15537), .C2(n11993), .A(n15536), .B(n15535), .ZN(
        P2_U2998) );
  NAND2_X1 U18833 ( .A1(n9897), .A2(n15539), .ZN(n15540) );
  XNOR2_X1 U18834 ( .A(n15541), .B(n15540), .ZN(n15740) );
  NAND2_X1 U18835 ( .A1(n16257), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15765) );
  AOI21_X1 U18836 ( .B1(n15746), .B2(n15543), .A(n15542), .ZN(n15738) );
  NAND2_X1 U18837 ( .A1(n15544), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n15729) );
  OAI21_X1 U18838 ( .B1(n16310), .B2(n15545), .A(n15729), .ZN(n15546) );
  AOI21_X1 U18839 ( .B1(n16301), .B2(n15547), .A(n15546), .ZN(n15548) );
  OAI21_X1 U18840 ( .B1(n15730), .B2(n13736), .A(n15548), .ZN(n15549) );
  AOI21_X1 U18841 ( .B1(n15738), .B2(n19236), .A(n15549), .ZN(n15550) );
  OAI21_X1 U18842 ( .B1(n15740), .B2(n11993), .A(n15550), .ZN(P2_U2999) );
  NAND2_X1 U18843 ( .A1(n16268), .A2(n15551), .ZN(n15552) );
  XOR2_X1 U18844 ( .A(n15552), .B(n9706), .Z(n15820) );
  INV_X1 U18845 ( .A(n15553), .ZN(n15556) );
  INV_X1 U18846 ( .A(n15554), .ZN(n15555) );
  AOI21_X1 U18847 ( .B1(n15556), .B2(n15810), .A(n15555), .ZN(n15818) );
  OAI22_X1 U18848 ( .A1(n16310), .A2(n15557), .B1(n11879), .B2(n19113), .ZN(
        n15560) );
  INV_X1 U18849 ( .A(n19088), .ZN(n15558) );
  OAI22_X1 U18850 ( .A1(n13736), .A2(n19092), .B1(n19240), .B2(n15558), .ZN(
        n15559) );
  AOI211_X1 U18851 ( .C1(n15818), .C2(n19236), .A(n15560), .B(n15559), .ZN(
        n15561) );
  OAI21_X1 U18852 ( .B1(n15820), .B2(n11993), .A(n15561), .ZN(P2_U3005) );
  INV_X1 U18853 ( .A(n15562), .ZN(n15576) );
  INV_X1 U18854 ( .A(n15563), .ZN(n15572) );
  NAND2_X1 U18855 ( .A1(n15564), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15569) );
  INV_X1 U18856 ( .A(n15565), .ZN(n15566) );
  AOI21_X1 U18857 ( .B1(n15567), .B2(n16331), .A(n15566), .ZN(n15568) );
  OAI21_X1 U18858 ( .B1(n15570), .B2(n15569), .A(n15568), .ZN(n15571) );
  AOI21_X1 U18859 ( .B1(n15572), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15571), .ZN(n15573) );
  OAI21_X1 U18860 ( .B1(n15574), .B2(n15816), .A(n15573), .ZN(n15575) );
  AOI21_X1 U18861 ( .B1(n15576), .B2(n16328), .A(n15575), .ZN(n15577) );
  OAI21_X1 U18862 ( .B1(n15578), .B2(n16320), .A(n15577), .ZN(P2_U3018) );
  INV_X1 U18863 ( .A(n15579), .ZN(n15588) );
  OAI21_X1 U18864 ( .B1(n15581), .B2(n15811), .A(n15580), .ZN(n15582) );
  AOI21_X1 U18865 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15583), .A(
        n15582), .ZN(n15585) );
  OAI211_X1 U18866 ( .C1(n15586), .C2(n15816), .A(n15585), .B(n15584), .ZN(
        n15587) );
  AOI21_X1 U18867 ( .B1(n15588), .B2(n16328), .A(n15587), .ZN(n15589) );
  OAI21_X1 U18868 ( .B1(n15590), .B2(n16320), .A(n15589), .ZN(P2_U3019) );
  OAI21_X1 U18869 ( .B1(n15592), .B2(n15811), .A(n15591), .ZN(n15593) );
  AOI21_X1 U18870 ( .B1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n15615), .A(
        n15593), .ZN(n15596) );
  OAI211_X1 U18871 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n15608), .B(n15594), .ZN(
        n15595) );
  OAI211_X1 U18872 ( .C1(n16206), .C2(n15816), .A(n15596), .B(n15595), .ZN(
        n15597) );
  AOI21_X1 U18873 ( .B1(n15598), .B2(n16328), .A(n15597), .ZN(n15599) );
  OAI21_X1 U18874 ( .B1(n15600), .B2(n16320), .A(n15599), .ZN(P2_U3020) );
  NAND2_X1 U18875 ( .A1(n15615), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15601) );
  OAI211_X1 U18876 ( .C1(n15603), .C2(n15811), .A(n15602), .B(n15601), .ZN(
        n15606) );
  NOR2_X1 U18877 ( .A1(n15604), .A2(n15816), .ZN(n15605) );
  AOI211_X1 U18878 ( .C1(n15608), .C2(n15607), .A(n15606), .B(n15605), .ZN(
        n15611) );
  NAND3_X1 U18879 ( .A1(n15412), .A2(n16328), .A3(n15609), .ZN(n15610) );
  OAI211_X1 U18880 ( .C1(n15612), .C2(n16320), .A(n15611), .B(n15610), .ZN(
        P2_U3021) );
  INV_X1 U18881 ( .A(n15613), .ZN(n15623) );
  INV_X1 U18882 ( .A(n15614), .ZN(n15620) );
  NAND2_X1 U18883 ( .A1(n15615), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15616) );
  OAI211_X1 U18884 ( .C1(n16218), .C2(n15811), .A(n15617), .B(n15616), .ZN(
        n15618) );
  AOI21_X1 U18885 ( .B1(n15620), .B2(n15619), .A(n15618), .ZN(n15621) );
  OAI21_X1 U18886 ( .B1(n16219), .B2(n15816), .A(n15621), .ZN(n15622) );
  AOI21_X1 U18887 ( .B1(n15623), .B2(n16328), .A(n15622), .ZN(n15624) );
  OAI21_X1 U18888 ( .B1(n15625), .B2(n16320), .A(n15624), .ZN(P2_U3022) );
  INV_X1 U18889 ( .A(n15648), .ZN(n15627) );
  OAI211_X1 U18890 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15627), .B(n15626), .ZN(
        n15632) );
  OAI21_X1 U18891 ( .B1(n15629), .B2(n15811), .A(n15628), .ZN(n15630) );
  INV_X1 U18892 ( .A(n15630), .ZN(n15631) );
  OAI211_X1 U18893 ( .C1(n15642), .C2(n15633), .A(n15632), .B(n15631), .ZN(
        n15634) );
  AOI21_X1 U18894 ( .B1(n15635), .B2(n16324), .A(n15634), .ZN(n15638) );
  NAND2_X1 U18895 ( .A1(n15636), .A2(n16328), .ZN(n15637) );
  OAI211_X1 U18896 ( .C1(n15639), .C2(n16320), .A(n15638), .B(n15637), .ZN(
        P2_U3023) );
  NAND2_X1 U18897 ( .A1(n15640), .A2(n16324), .ZN(n15647) );
  NOR2_X1 U18898 ( .A1(n15642), .A2(n15641), .ZN(n15643) );
  AOI211_X1 U18899 ( .C1(n15645), .C2(n16331), .A(n15644), .B(n15643), .ZN(
        n15646) );
  OAI211_X1 U18900 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n15648), .A(
        n15647), .B(n15646), .ZN(n15649) );
  AOI21_X1 U18901 ( .B1(n15650), .B2(n16332), .A(n15649), .ZN(n15651) );
  OAI21_X1 U18902 ( .B1(n15804), .B2(n15652), .A(n15651), .ZN(P2_U3024) );
  INV_X1 U18903 ( .A(n15653), .ZN(n15655) );
  OAI21_X1 U18904 ( .B1(n15655), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15654), .ZN(n15657) );
  OAI211_X1 U18905 ( .C1(n15811), .C2(n15658), .A(n15657), .B(n15656), .ZN(
        n15661) );
  NOR2_X1 U18906 ( .A1(n15659), .A2(n15804), .ZN(n15660) );
  AOI211_X1 U18907 ( .C1(n16324), .C2(n18984), .A(n15661), .B(n15660), .ZN(
        n15662) );
  OAI21_X1 U18908 ( .B1(n15663), .B2(n16320), .A(n15662), .ZN(P2_U3025) );
  NAND2_X1 U18909 ( .A1(n15665), .A2(n15664), .ZN(n15666) );
  AND2_X1 U18910 ( .A1(n15667), .A2(n15666), .ZN(n18990) );
  XNOR2_X1 U18911 ( .A(n15673), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15668) );
  NAND2_X1 U18912 ( .A1(n15685), .A2(n15668), .ZN(n15672) );
  AOI21_X1 U18913 ( .B1(n15670), .B2(n16331), .A(n15669), .ZN(n15671) );
  OAI211_X1 U18914 ( .C1(n15691), .C2(n15673), .A(n15672), .B(n15671), .ZN(
        n15676) );
  NOR2_X1 U18915 ( .A1(n15674), .A2(n15804), .ZN(n15675) );
  AOI211_X1 U18916 ( .C1(n16324), .C2(n18990), .A(n15676), .B(n15675), .ZN(
        n15677) );
  OAI21_X1 U18917 ( .B1(n15678), .B2(n16320), .A(n15677), .ZN(P2_U3026) );
  OR3_X1 U18918 ( .A1(n15680), .A2(n15679), .A3(n15804), .ZN(n15687) );
  NAND2_X1 U18919 ( .A1(n19004), .A2(n16331), .ZN(n15681) );
  OAI211_X1 U18920 ( .C1(n15691), .C2(n15684), .A(n15682), .B(n15681), .ZN(
        n15683) );
  AOI21_X1 U18921 ( .B1(n15685), .B2(n15684), .A(n15683), .ZN(n15686) );
  OAI211_X1 U18922 ( .C1(n15816), .C2(n19010), .A(n15687), .B(n15686), .ZN(
        n15688) );
  INV_X1 U18923 ( .A(n15688), .ZN(n15689) );
  OAI21_X1 U18924 ( .B1(n15690), .B2(n16320), .A(n15689), .ZN(P2_U3027) );
  INV_X1 U18925 ( .A(n15691), .ZN(n15695) );
  OAI21_X1 U18926 ( .B1(n15693), .B2(n15811), .A(n15692), .ZN(n15694) );
  AOI21_X1 U18927 ( .B1(n15695), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15694), .ZN(n15700) );
  INV_X1 U18928 ( .A(n15731), .ZN(n15698) );
  NAND3_X1 U18929 ( .A1(n15698), .A2(n15697), .A3(n15696), .ZN(n15699) );
  OAI211_X1 U18930 ( .C1(n16238), .C2(n15816), .A(n15700), .B(n15699), .ZN(
        n15701) );
  AOI21_X1 U18931 ( .B1(n15702), .B2(n16328), .A(n15701), .ZN(n15703) );
  OAI21_X1 U18932 ( .B1(n15704), .B2(n16320), .A(n15703), .ZN(P2_U3028) );
  OR2_X1 U18933 ( .A1(n15705), .A2(n16328), .ZN(n15709) );
  NOR2_X1 U18934 ( .A1(n15706), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15707) );
  OR2_X1 U18935 ( .A1(n15734), .A2(n15707), .ZN(n15708) );
  AOI21_X1 U18936 ( .B1(n15500), .B2(n15709), .A(n15708), .ZN(n15722) );
  OAI21_X1 U18937 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15710), .A(
        n15722), .ZN(n15716) );
  NAND2_X1 U18938 ( .A1(n19011), .A2(n16324), .ZN(n15712) );
  OAI211_X1 U18939 ( .C1(n19015), .C2(n15811), .A(n15712), .B(n15711), .ZN(
        n15715) );
  OAI21_X1 U18940 ( .B1(n15746), .B2(n15804), .A(n15731), .ZN(n15713) );
  NAND2_X1 U18941 ( .A1(n15713), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15728) );
  NOR3_X1 U18942 ( .A1(n15728), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15721), .ZN(n15714) );
  AOI211_X1 U18943 ( .C1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n15716), .A(
        n15715), .B(n15714), .ZN(n15717) );
  OAI21_X1 U18944 ( .B1(n15718), .B2(n16320), .A(n15717), .ZN(P2_U3029) );
  NAND2_X1 U18945 ( .A1(n15719), .A2(n16332), .ZN(n15727) );
  OAI21_X1 U18946 ( .B1(n19030), .B2(n15811), .A(n15720), .ZN(n15724) );
  NOR2_X1 U18947 ( .A1(n15722), .A2(n15721), .ZN(n15723) );
  AOI211_X1 U18948 ( .C1(n16324), .C2(n15725), .A(n15724), .B(n15723), .ZN(
        n15726) );
  OAI211_X1 U18949 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15728), .A(
        n15727), .B(n15726), .ZN(P2_U3030) );
  OAI21_X1 U18950 ( .B1(n15811), .B2(n15730), .A(n15729), .ZN(n15733) );
  NOR2_X1 U18951 ( .A1(n15731), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15732) );
  AOI211_X1 U18952 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15734), .A(
        n15733), .B(n15732), .ZN(n15735) );
  OAI21_X1 U18953 ( .B1(n15816), .B2(n15736), .A(n15735), .ZN(n15737) );
  AOI21_X1 U18954 ( .B1(n15738), .B2(n16328), .A(n15737), .ZN(n15739) );
  OAI21_X1 U18955 ( .B1(n15740), .B2(n16320), .A(n15739), .ZN(P2_U3031) );
  NAND2_X1 U18956 ( .A1(n15742), .A2(n15741), .ZN(n15743) );
  XNOR2_X1 U18957 ( .A(n15744), .B(n15743), .ZN(n16244) );
  INV_X1 U18958 ( .A(n16244), .ZN(n15759) );
  NAND2_X1 U18959 ( .A1(n15765), .A2(n15753), .ZN(n15745) );
  AND2_X1 U18960 ( .A1(n15748), .A2(n15747), .ZN(n15749) );
  OR2_X1 U18961 ( .A1(n15749), .A2(n12857), .ZN(n19154) );
  NAND2_X1 U18962 ( .A1(n15766), .A2(n11704), .ZN(n15785) );
  NAND2_X1 U18963 ( .A1(n15787), .A2(n15785), .ZN(n15767) );
  AOI21_X1 U18964 ( .B1(n15766), .B2(n15769), .A(n15767), .ZN(n15751) );
  NAND2_X1 U18965 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n11988), .ZN(n15750) );
  OAI21_X1 U18966 ( .B1(n15753), .B2(n15751), .A(n15750), .ZN(n15752) );
  AOI21_X1 U18967 ( .B1(n16331), .B2(n19044), .A(n15752), .ZN(n15756) );
  NAND3_X1 U18968 ( .A1(n15766), .A2(n15754), .A3(n15753), .ZN(n15755) );
  OAI211_X1 U18969 ( .C1(n19154), .C2(n15816), .A(n15756), .B(n15755), .ZN(
        n15757) );
  AOI21_X1 U18970 ( .B1(n16243), .B2(n16328), .A(n15757), .ZN(n15758) );
  OAI21_X1 U18971 ( .B1(n15759), .B2(n16320), .A(n15758), .ZN(P2_U3032) );
  NAND2_X1 U18972 ( .A1(n15761), .A2(n15760), .ZN(n15762) );
  XNOR2_X1 U18973 ( .A(n15763), .B(n15762), .ZN(n16248) );
  OR2_X1 U18974 ( .A1(n16257), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15764) );
  NAND2_X1 U18975 ( .A1(n15765), .A2(n15764), .ZN(n16247) );
  INV_X1 U18976 ( .A(n16247), .ZN(n15775) );
  NOR2_X1 U18977 ( .A1(n11895), .A2(n19113), .ZN(n15772) );
  NAND2_X1 U18978 ( .A1(n15766), .A2(n15769), .ZN(n15770) );
  INV_X1 U18979 ( .A(n15767), .ZN(n15768) );
  OAI22_X1 U18980 ( .A1(n15770), .A2(n11704), .B1(n15769), .B2(n15768), .ZN(
        n15771) );
  AOI211_X1 U18981 ( .C1(n16331), .C2(n16250), .A(n15772), .B(n15771), .ZN(
        n15773) );
  OAI21_X1 U18982 ( .B1(n19056), .B2(n15816), .A(n15773), .ZN(n15774) );
  AOI21_X1 U18983 ( .B1(n15775), .B2(n16328), .A(n15774), .ZN(n15776) );
  OAI21_X1 U18984 ( .B1(n16248), .B2(n16320), .A(n15776), .ZN(P2_U3033) );
  INV_X1 U18985 ( .A(n15777), .ZN(n15778) );
  NOR2_X1 U18986 ( .A1(n15779), .A2(n15778), .ZN(n15781) );
  XOR2_X1 U18987 ( .A(n15781), .B(n9646), .Z(n16259) );
  INV_X1 U18988 ( .A(n16259), .ZN(n15793) );
  INV_X1 U18989 ( .A(n16255), .ZN(n19067) );
  AOI21_X1 U18990 ( .B1(n15784), .B2(n15783), .A(n15782), .ZN(n19066) );
  INV_X1 U18991 ( .A(n19066), .ZN(n19157) );
  NAND2_X1 U18992 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n11988), .ZN(n15786) );
  OAI211_X1 U18993 ( .C1(n15816), .C2(n19157), .A(n15786), .B(n15785), .ZN(
        n15789) );
  NOR2_X1 U18994 ( .A1(n15787), .A2(n11704), .ZN(n15788) );
  AOI211_X1 U18995 ( .C1(n19067), .C2(n16331), .A(n15789), .B(n15788), .ZN(
        n15792) );
  INV_X1 U18996 ( .A(n16257), .ZN(n15790) );
  NAND2_X1 U18997 ( .A1(n15533), .A2(n11704), .ZN(n16254) );
  NAND3_X1 U18998 ( .A1(n15790), .A2(n16328), .A3(n16254), .ZN(n15791) );
  OAI211_X1 U18999 ( .C1(n15793), .C2(n16320), .A(n15792), .B(n15791), .ZN(
        P2_U3034) );
  XOR2_X1 U19000 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n15795), .Z(
        n15796) );
  XNOR2_X1 U19001 ( .A(n9641), .B(n15796), .ZN(n16263) );
  AOI211_X1 U19002 ( .C1(n15802), .C2(n11883), .A(n15810), .B(n15797), .ZN(
        n15807) );
  AOI21_X1 U19003 ( .B1(n15810), .B2(n15798), .A(n15813), .ZN(n16313) );
  NOR2_X1 U19004 ( .A1(n11888), .A2(n19113), .ZN(n15800) );
  NOR2_X1 U19005 ( .A1(n15816), .A2(n19078), .ZN(n15799) );
  AOI211_X1 U19006 ( .C1(n10163), .C2(n16331), .A(n15800), .B(n15799), .ZN(
        n15801) );
  OAI21_X1 U19007 ( .B1(n16313), .B2(n15802), .A(n15801), .ZN(n15806) );
  OR2_X1 U19008 ( .A1(n15554), .A2(n11883), .ZN(n16273) );
  INV_X1 U19009 ( .A(n16273), .ZN(n15803) );
  OAI21_X1 U19010 ( .B1(n15803), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15533), .ZN(n16262) );
  NOR2_X1 U19011 ( .A1(n16262), .A2(n15804), .ZN(n15805) );
  AOI211_X1 U19012 ( .C1(n15808), .C2(n15807), .A(n15806), .B(n15805), .ZN(
        n15809) );
  OAI21_X1 U19013 ( .B1(n16263), .B2(n16320), .A(n15809), .ZN(P2_U3035) );
  NAND2_X1 U19014 ( .A1(n16311), .A2(n15810), .ZN(n15815) );
  OAI22_X1 U19015 ( .A1(n15811), .A2(n19092), .B1(n11879), .B2(n19113), .ZN(
        n15812) );
  AOI21_X1 U19016 ( .B1(n15813), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15812), .ZN(n15814) );
  OAI211_X1 U19017 ( .C1(n19093), .C2(n15816), .A(n15815), .B(n15814), .ZN(
        n15817) );
  AOI21_X1 U19018 ( .B1(n15818), .B2(n16328), .A(n15817), .ZN(n15819) );
  OAI21_X1 U19019 ( .B1(n15820), .B2(n16320), .A(n15819), .ZN(P2_U3037) );
  INV_X1 U19020 ( .A(n18952), .ZN(n19929) );
  MUX2_X1 U19021 ( .A(n15821), .B(n15848), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15822) );
  AOI21_X1 U19022 ( .B1(n15823), .B2(n15858), .A(n15822), .ZN(n16341) );
  INV_X1 U19023 ( .A(n15824), .ZN(n15825) );
  OAI222_X1 U19024 ( .A1(n16388), .A2(n15826), .B1(n19929), .B2(n16341), .C1(
        n11444), .C2(n15825), .ZN(n15827) );
  INV_X1 U19025 ( .A(n15860), .ZN(n15904) );
  MUX2_X1 U19026 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n15827), .S(
        n15904), .Z(P2_U3601) );
  AOI21_X1 U19027 ( .B1(n9732), .B2(n15828), .A(n11375), .ZN(n15852) );
  INV_X1 U19028 ( .A(n15829), .ZN(n15830) );
  NAND2_X1 U19029 ( .A1(n15830), .A2(n11223), .ZN(n15846) );
  INV_X1 U19030 ( .A(n11221), .ZN(n15831) );
  NAND2_X1 U19031 ( .A1(n15848), .A2(n15831), .ZN(n15854) );
  NOR2_X1 U19032 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n15832), .ZN(
        n15833) );
  NOR2_X1 U19033 ( .A1(n15854), .A2(n15833), .ZN(n15834) );
  AOI21_X1 U19034 ( .B1(n15852), .B2(n15846), .A(n15834), .ZN(n15839) );
  INV_X1 U19035 ( .A(n15846), .ZN(n15851) );
  INV_X1 U19036 ( .A(n15835), .ZN(n16362) );
  NAND2_X1 U19037 ( .A1(n16362), .A2(n15836), .ZN(n15847) );
  OAI21_X1 U19038 ( .B1(n11375), .B2(n15851), .A(n15847), .ZN(n15838) );
  OAI211_X1 U19039 ( .C1(n15841), .C2(n15840), .A(n15839), .B(n15838), .ZN(
        n16356) );
  AOI22_X1 U19040 ( .A1(n16356), .A2(n18952), .B1(n15843), .B2(n15842), .ZN(
        n15844) );
  OAI21_X1 U19041 ( .B1(n19942), .B2(n16388), .A(n15844), .ZN(n15845) );
  MUX2_X1 U19042 ( .A(n15845), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15860), .Z(P2_U3599) );
  NAND2_X1 U19043 ( .A1(n15847), .A2(n15846), .ZN(n15850) );
  AOI21_X1 U19044 ( .B1(n15848), .B2(n11221), .A(n11375), .ZN(n15849) );
  NAND2_X1 U19045 ( .A1(n15850), .A2(n15849), .ZN(n15856) );
  INV_X1 U19046 ( .A(n15852), .ZN(n15853) );
  NAND3_X1 U19047 ( .A1(n15846), .A2(n15854), .A3(n15853), .ZN(n15855) );
  MUX2_X1 U19048 ( .A(n15856), .B(n15855), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15857) );
  AOI21_X1 U19049 ( .B1(n15859), .B2(n15858), .A(n15857), .ZN(n16351) );
  OAI22_X1 U19050 ( .A1(n19934), .A2(n16388), .B1(n16351), .B2(n19929), .ZN(
        n15861) );
  MUX2_X1 U19051 ( .A(n15861), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15860), .Z(P2_U3596) );
  NAND2_X1 U19052 ( .A1(n17274), .A2(P3_EBX_REG_13__SCAN_IN), .ZN(n15876) );
  AOI22_X1 U19053 ( .A1(n17225), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15872) );
  AOI22_X1 U19054 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15862) );
  OAI21_X1 U19055 ( .B1(n17099), .B2(n17022), .A(n15862), .ZN(n15870) );
  AOI22_X1 U19056 ( .A1(n9631), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9630), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15868) );
  INV_X1 U19057 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17260) );
  AOI22_X1 U19058 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15865) );
  AOI22_X1 U19059 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15863), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15864) );
  OAI211_X1 U19060 ( .C1(n17235), .C2(n17260), .A(n15865), .B(n15864), .ZN(
        n15866) );
  AOI21_X1 U19061 ( .B1(n12616), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n15866), .ZN(n15867) );
  OAI211_X1 U19062 ( .C1(n17035), .C2(n17029), .A(n15868), .B(n15867), .ZN(
        n15869) );
  AOI211_X1 U19063 ( .C1(n17142), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n15870), .B(n15869), .ZN(n15871) );
  OAI211_X1 U19064 ( .C1(n17217), .C2(n15873), .A(n15872), .B(n15871), .ZN(
        n17387) );
  NOR2_X1 U19065 ( .A1(n18294), .A2(n15874), .ZN(n17160) );
  AOI22_X1 U19066 ( .A1(n17282), .A2(n17387), .B1(n17160), .B2(n16772), .ZN(
        n15875) );
  OAI21_X1 U19067 ( .B1(n15877), .B2(n15876), .A(n15875), .ZN(P3_U2690) );
  INV_X1 U19068 ( .A(n17820), .ZN(n17750) );
  NAND2_X1 U19069 ( .A1(n15878), .A2(n17750), .ZN(n15882) );
  NAND2_X1 U19070 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18264) );
  NAND3_X1 U19071 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18881)
         );
  AOI21_X1 U19072 ( .B1(n18712), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15899) );
  NAND2_X1 U19073 ( .A1(n15899), .A2(n17227), .ZN(n18254) );
  INV_X1 U19074 ( .A(n18254), .ZN(n15879) );
  INV_X1 U19075 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18255) );
  OR2_X1 U19076 ( .A1(n18255), .A2(n18881), .ZN(n15897) );
  OAI211_X1 U19077 ( .C1(n18881), .C2(n15879), .A(n18345), .B(n15897), .ZN(
        n18261) );
  INV_X1 U19078 ( .A(n18261), .ZN(n15884) );
  AOI21_X1 U19079 ( .B1(n15882), .B2(n18264), .A(n15884), .ZN(n15885) );
  INV_X1 U19080 ( .A(n15885), .ZN(n15881) );
  INV_X1 U19081 ( .A(n18508), .ZN(n18626) );
  NOR2_X1 U19082 ( .A1(n18883), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18256) );
  INV_X1 U19083 ( .A(n18256), .ZN(n18302) );
  NAND2_X1 U19084 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18302), .ZN(
        n18344) );
  NOR3_X1 U19085 ( .A1(n18626), .A2(n15884), .A3(n18344), .ZN(n15880) );
  AOI21_X1 U19086 ( .B1(n18743), .B2(n15881), .A(n15880), .ZN(P3_U2864) );
  NOR2_X1 U19087 ( .A1(n18761), .A2(n18743), .ZN(n18434) );
  AOI22_X1 U19088 ( .A1(n18434), .A2(n18302), .B1(n18883), .B2(n15882), .ZN(
        n15883) );
  NOR2_X1 U19089 ( .A1(n15884), .A2(n15883), .ZN(n18260) );
  AOI22_X1 U19090 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n15885), .B1(
        n18626), .B2(n18261), .ZN(n18259) );
  AOI22_X1 U19091 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18260), .B1(
        n18259), .B2(n18761), .ZN(P3_U2865) );
  NOR2_X1 U19092 ( .A1(n15886), .A2(n18730), .ZN(n15887) );
  NOR3_X4 U19093 ( .A1(n18785), .A2(n15887), .A3(n16553), .ZN(n15990) );
  NAND2_X1 U19094 ( .A1(n18755), .A2(n18933), .ZN(n15894) );
  INV_X1 U19095 ( .A(n18930), .ZN(n15907) );
  AOI21_X1 U19096 ( .B1(n15891), .B2(n15890), .A(n15889), .ZN(n15892) );
  NOR2_X1 U19097 ( .A1(n15893), .A2(n15892), .ZN(n15913) );
  OAI21_X1 U19098 ( .B1(n15894), .B2(n17446), .A(n15913), .ZN(n15895) );
  AOI211_X4 U19099 ( .C1(n15896), .C2(n18752), .A(n15990), .B(n15895), .ZN(
        n18766) );
  NAND2_X1 U19100 ( .A1(n18783), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18266) );
  INV_X1 U19101 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16879) );
  INV_X1 U19102 ( .A(n18892), .ZN(n18902) );
  NOR2_X1 U19103 ( .A1(n15899), .A2(n15898), .ZN(n18765) );
  NAND3_X1 U19104 ( .A1(n18910), .A2(n18902), .A3(n18765), .ZN(n15900) );
  OAI21_X1 U19105 ( .B1(n18910), .B2(n16879), .A(n15900), .ZN(P3_U3284) );
  NOR4_X1 U19106 ( .A1(n12265), .A2(n16364), .A3(n19989), .A4(n19929), .ZN(
        n15901) );
  NAND2_X1 U19107 ( .A1(n15904), .A2(n15901), .ZN(n15902) );
  OAI21_X1 U19108 ( .B1(n15904), .B2(n15903), .A(n15902), .ZN(P2_U3595) );
  INV_X1 U19109 ( .A(n16438), .ZN(n15926) );
  AOI21_X1 U19110 ( .B1(n18273), .B2(n15906), .A(n15905), .ZN(n15915) );
  AOI21_X1 U19111 ( .B1(n18932), .B2(n15908), .A(n15907), .ZN(n15910) );
  AOI21_X1 U19112 ( .B1(n15910), .B2(n15909), .A(n18785), .ZN(n16554) );
  NAND3_X1 U19113 ( .A1(n18755), .A2(n16554), .A3(n15911), .ZN(n15912) );
  OAI211_X1 U19114 ( .C1(n15915), .C2(n15914), .A(n15913), .B(n15912), .ZN(
        n15918) );
  INV_X1 U19115 ( .A(n15916), .ZN(n18756) );
  NOR2_X1 U19116 ( .A1(n16437), .A2(n18240), .ZN(n18166) );
  NAND2_X1 U19117 ( .A1(n18750), .A2(n18243), .ZN(n18230) );
  NOR2_X1 U19118 ( .A1(n12642), .A2(n18890), .ZN(n18197) );
  INV_X1 U19119 ( .A(n18197), .ZN(n15919) );
  NAND3_X1 U19120 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18032) );
  NOR2_X1 U19121 ( .A1(n15919), .A2(n18032), .ZN(n18157) );
  NAND2_X1 U19122 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18162) );
  NOR2_X1 U19123 ( .A1(n10018), .A2(n18162), .ZN(n18033) );
  NAND2_X1 U19124 ( .A1(n18157), .A2(n18033), .ZN(n18094) );
  NOR2_X1 U19125 ( .A1(n18035), .A2(n18094), .ZN(n18024) );
  NOR2_X1 U19126 ( .A1(n17693), .A2(n17645), .ZN(n17984) );
  NAND2_X1 U19127 ( .A1(n18024), .A2(n17984), .ZN(n17921) );
  NOR2_X1 U19128 ( .A1(n17992), .A2(n17921), .ZN(n17922) );
  INV_X1 U19129 ( .A(n17922), .ZN(n15923) );
  INV_X1 U19130 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18251) );
  OAI21_X1 U19131 ( .B1(n18251), .B2(n18890), .A(n12642), .ZN(n18031) );
  INV_X1 U19132 ( .A(n18031), .ZN(n18195) );
  NOR2_X1 U19133 ( .A1(n18195), .A2(n18032), .ZN(n18156) );
  NAND2_X1 U19134 ( .A1(n18033), .A2(n18156), .ZN(n18047) );
  NOR2_X1 U19135 ( .A1(n18035), .A2(n18047), .ZN(n17975) );
  AND2_X1 U19136 ( .A1(n15920), .A2(n17975), .ZN(n17958) );
  NOR2_X1 U19137 ( .A1(n18251), .A2(n18094), .ZN(n18107) );
  NAND2_X1 U19138 ( .A1(n16442), .A2(n18107), .ZN(n18045) );
  NOR2_X1 U19139 ( .A1(n17968), .A2(n18045), .ZN(n15921) );
  AOI22_X1 U19140 ( .A1(n18751), .A2(n17958), .B1(n15921), .B2(n18738), .ZN(
        n15922) );
  OAI21_X1 U19141 ( .B1(n18740), .B2(n15923), .A(n15922), .ZN(n17941) );
  NAND4_X1 U19142 ( .A1(n15927), .A2(n15924), .A3(n18243), .A4(n17941), .ZN(
        n16423) );
  OAI21_X1 U19143 ( .B1(n18230), .B2(n16439), .A(n16423), .ZN(n15925) );
  AOI21_X1 U19144 ( .B1(n15926), .B2(n18166), .A(n15925), .ZN(n15975) );
  INV_X1 U19145 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16419) );
  NOR3_X1 U19146 ( .A1(n17918), .A2(n17917), .A3(n18045), .ZN(n15930) );
  AOI21_X1 U19147 ( .B1(n15927), .B2(n17922), .A(n18740), .ZN(n15928) );
  NOR2_X1 U19148 ( .A1(n17968), .A2(n17923), .ZN(n17598) );
  AOI21_X1 U19149 ( .B1(n17975), .B2(n17598), .A(n18721), .ZN(n17940) );
  AOI211_X1 U19150 ( .C1(n18751), .C2(n17924), .A(n15928), .B(n17940), .ZN(
        n15929) );
  INV_X2 U19151 ( .A(n18140), .ZN(n18071) );
  NOR2_X2 U19152 ( .A1(n18071), .A2(n18243), .ZN(n18242) );
  OAI211_X1 U19153 ( .C1(n18128), .C2(n15930), .A(n15929), .B(n18233), .ZN(
        n16434) );
  INV_X1 U19154 ( .A(n18200), .ZN(n18052) );
  OAI22_X1 U19155 ( .A1(n18138), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n18052), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15932) );
  AOI22_X1 U19156 ( .A1(n16397), .A2(n18166), .B1(n16398), .B2(n18246), .ZN(
        n15931) );
  INV_X1 U19157 ( .A(n15931), .ZN(n15977) );
  AOI221_X1 U19158 ( .B1(n16434), .B2(n18140), .C1(n15932), .C2(n18140), .A(
        n15977), .ZN(n15935) );
  XOR2_X1 U19159 ( .A(n16419), .B(n15933), .Z(n16417) );
  AOI22_X1 U19160 ( .A1(n18071), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n18151), 
        .B2(n16417), .ZN(n15934) );
  OAI221_X1 U19161 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15975), 
        .C1(n16419), .C2(n15935), .A(n15934), .ZN(P3_U2833) );
  INV_X1 U19162 ( .A(n15946), .ZN(n15948) );
  INV_X1 U19163 ( .A(n15936), .ZN(n15938) );
  NOR3_X1 U19164 ( .A1(n15938), .A2(n15937), .A3(n20692), .ZN(n15943) );
  INV_X1 U19165 ( .A(n15939), .ZN(n15942) );
  INV_X1 U19166 ( .A(n15940), .ZN(n15941) );
  OAI22_X1 U19167 ( .A1(n15943), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n15942), .B2(n15941), .ZN(n15945) );
  NAND2_X1 U19168 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n15943), .ZN(
        n15944) );
  OAI211_X1 U19169 ( .C1(n15946), .C2(n20646), .A(n15945), .B(n15944), .ZN(
        n15947) );
  OAI21_X1 U19170 ( .B1(n15948), .B2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n15947), .ZN(n15950) );
  AOI222_X1 U19171 ( .A1(n15950), .A2(n20645), .B1(n15950), .B2(n15949), .C1(
        n20645), .C2(n15949), .ZN(n15959) );
  INV_X1 U19172 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n21069) );
  AND2_X1 U19173 ( .A1(n20008), .A2(n21069), .ZN(n15952) );
  OAI21_X1 U19174 ( .B1(n15953), .B2(n15952), .A(n15951), .ZN(n15954) );
  NOR3_X1 U19175 ( .A1(n15956), .A2(n15955), .A3(n15954), .ZN(n15957) );
  OAI211_X1 U19176 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n15959), .A(
        n15958), .B(n15957), .ZN(n15964) );
  NOR3_X1 U19177 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20837), .A3(n20918), 
        .ZN(n15962) );
  NAND2_X1 U19178 ( .A1(n21034), .A2(n20918), .ZN(n15960) );
  OAI22_X1 U19179 ( .A1(n15965), .A2(n15962), .B1(n15961), .B2(n15960), .ZN(
        n16179) );
  AOI221_X1 U19180 ( .B1(n20914), .B2(n16181), .C1(n15964), .C2(n16181), .A(
        n16179), .ZN(n15966) );
  NOR2_X1 U19181 ( .A1(n15966), .A2(n20914), .ZN(n20836) );
  OAI211_X1 U19182 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20918), .A(n20836), 
        .B(n15963), .ZN(n16180) );
  AOI21_X1 U19183 ( .B1(n15965), .B2(n15964), .A(n16180), .ZN(n15972) );
  AOI21_X1 U19184 ( .B1(n15968), .B2(n15967), .A(n15966), .ZN(n15969) );
  INV_X1 U19185 ( .A(n15969), .ZN(n15970) );
  AOI22_X1 U19186 ( .A1(n15972), .A2(n15971), .B1(n20914), .B2(n15970), .ZN(
        P1_U3161) );
  OAI21_X1 U19187 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15974), .A(
        n15973), .ZN(n16407) );
  NAND2_X1 U19188 ( .A1(n18200), .A2(n18243), .ZN(n18234) );
  NAND2_X1 U19189 ( .A1(n18140), .A2(n16434), .ZN(n15976) );
  OAI21_X1 U19190 ( .B1(n16404), .B2(n18234), .A(n15976), .ZN(n16421) );
  NOR2_X1 U19191 ( .A1(n16421), .A2(n15977), .ZN(n15978) );
  MUX2_X1 U19192 ( .A(n10152), .B(n15978), .S(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(n15979) );
  NAND2_X1 U19193 ( .A1(n18071), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16399) );
  OAI211_X1 U19194 ( .C1(n18170), .C2(n16407), .A(n15979), .B(n16399), .ZN(
        P3_U2832) );
  INV_X1 U19195 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20853) );
  INV_X1 U19196 ( .A(HOLD), .ZN(n21063) );
  NOR2_X1 U19197 ( .A1(n20853), .A2(n21063), .ZN(n20842) );
  AOI22_X1 U19198 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15982) );
  NAND2_X1 U19199 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n15980), .ZN(n20840) );
  OAI211_X1 U19200 ( .C1(n20842), .C2(n15982), .A(n15981), .B(n20840), .ZN(
        P1_U3195) );
  AND2_X1 U19201 ( .A1(n15983), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NAND2_X1 U19202 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19769), .ZN(n19844) );
  NOR2_X1 U19203 ( .A1(n19985), .A2(n19844), .ZN(n16381) );
  AOI221_X1 U19204 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .C1(P2_STATE2_REG_0__SCAN_IN), .C2(
        P2_STATE2_REG_1__SCAN_IN), .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n15984)
         );
  NOR3_X1 U19205 ( .A1(n16381), .A2(n16382), .A3(n15984), .ZN(P2_U3178) );
  INV_X1 U19206 ( .A(n16382), .ZN(n16396) );
  OAI221_X1 U19207 ( .B1(n15985), .B2(n16396), .C1(n19968), .C2(n16396), .A(
        n19466), .ZN(n19965) );
  NOR2_X1 U19208 ( .A1(n15986), .A2(n19965), .ZN(P2_U3047) );
  OAI21_X2 U19209 ( .B1(n15990), .B2(n15989), .A(n18927), .ZN(n17438) );
  NOR2_X1 U19210 ( .A1(n18294), .A2(n17438), .ZN(n17441) );
  INV_X1 U19211 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17517) );
  INV_X1 U19212 ( .A(n17438), .ZN(n15994) );
  AOI22_X1 U19213 ( .A1(n17439), .A2(BUF2_REG_0__SCAN_IN), .B1(n17409), .B2(
        n17911), .ZN(n15993) );
  OAI221_X1 U19214 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17414), .C1(n17517), 
        .C2(n15994), .A(n15993), .ZN(P3_U2735) );
  NAND3_X1 U19215 ( .A1(n15995), .A2(P1_REIP_REG_15__SCAN_IN), .A3(n14049), 
        .ZN(n15999) );
  OAI21_X1 U19216 ( .B1(n15997), .B2(n15996), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n15998) );
  OAI211_X1 U19217 ( .C1(n16000), .C2(n14519), .A(n15999), .B(n15998), .ZN(
        n16001) );
  AOI211_X1 U19218 ( .C1(n20091), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20167), .B(n16001), .ZN(n16004) );
  AOI22_X1 U19219 ( .A1(n16034), .A2(n20058), .B1(n20089), .B2(n16002), .ZN(
        n16003) );
  OAI211_X1 U19220 ( .C1(n16037), .C2(n20078), .A(n16004), .B(n16003), .ZN(
        P1_U2824) );
  OAI21_X1 U19221 ( .B1(n20067), .B2(n16005), .A(n20064), .ZN(n16010) );
  AOI21_X1 U19222 ( .B1(n16006), .B2(n20023), .A(P1_REIP_REG_14__SCAN_IN), 
        .ZN(n16008) );
  NOR2_X1 U19223 ( .A1(n16008), .A2(n16007), .ZN(n16009) );
  AOI211_X1 U19224 ( .C1(P1_EBX_REG_14__SCAN_IN), .C2(n20088), .A(n16010), .B(
        n16009), .ZN(n16013) );
  INV_X1 U19225 ( .A(n16011), .ZN(n16045) );
  AOI22_X1 U19226 ( .A1(n16045), .A2(n20058), .B1(n20093), .B2(n16043), .ZN(
        n16012) );
  OAI211_X1 U19227 ( .C1(n20086), .C2(n16108), .A(n16013), .B(n16012), .ZN(
        P1_U2826) );
  AOI22_X1 U19228 ( .A1(n20088), .A2(P1_EBX_REG_12__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n20091), .ZN(n16022) );
  AOI21_X1 U19229 ( .B1(n20089), .B2(n16014), .A(n20167), .ZN(n16021) );
  INV_X1 U19230 ( .A(n16015), .ZN(n16048) );
  OAI22_X1 U19231 ( .A1(n16050), .A2(n20029), .B1(n20078), .B2(n16048), .ZN(
        n16016) );
  INV_X1 U19232 ( .A(n16016), .ZN(n16020) );
  AND2_X1 U19233 ( .A1(n16017), .A2(n20023), .ZN(n16029) );
  OAI221_X1 U19234 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(P1_REIP_REG_11__SCAN_IN), .C1(P1_REIP_REG_12__SCAN_IN), .C2(n16029), .A(n16018), .ZN(n16019) );
  NAND4_X1 U19235 ( .A1(n16022), .A2(n16021), .A3(n16020), .A4(n16019), .ZN(
        P1_U2828) );
  INV_X1 U19236 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n16028) );
  OAI22_X1 U19237 ( .A1(n16118), .A2(n20086), .B1(n14519), .B2(n16023), .ZN(
        n16024) );
  INV_X1 U19238 ( .A(n16024), .ZN(n16025) );
  OAI211_X1 U19239 ( .C1(n20067), .C2(n10615), .A(n16025), .B(n20064), .ZN(
        n16026) );
  AOI221_X1 U19240 ( .B1(n16029), .B2(n16028), .C1(n16027), .C2(
        P1_REIP_REG_11__SCAN_IN), .A(n16026), .ZN(n16032) );
  INV_X1 U19241 ( .A(n16030), .ZN(n16058) );
  NAND2_X1 U19242 ( .A1(n16058), .A2(n20058), .ZN(n16031) );
  OAI211_X1 U19243 ( .C1(n20078), .C2(n16061), .A(n16032), .B(n16031), .ZN(
        P1_U2829) );
  AOI22_X1 U19244 ( .A1(n20168), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20167), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16036) );
  AOI22_X1 U19245 ( .A1(n16034), .A2(n20239), .B1(n20174), .B2(n16033), .ZN(
        n16035) );
  OAI211_X1 U19246 ( .C1(n20178), .C2(n16037), .A(n16036), .B(n16035), .ZN(
        P1_U2983) );
  INV_X1 U19247 ( .A(n16038), .ZN(n16039) );
  AOI21_X1 U19248 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n12224), .A(
        n16040), .ZN(n16042) );
  XNOR2_X1 U19249 ( .A(n9672), .B(n16114), .ZN(n16041) );
  XNOR2_X1 U19250 ( .A(n16042), .B(n16041), .ZN(n16109) );
  AOI22_X1 U19251 ( .A1(n20168), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20167), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16047) );
  AOI22_X1 U19252 ( .A1(n16045), .A2(n20239), .B1(n16044), .B2(n16043), .ZN(
        n16046) );
  OAI211_X1 U19253 ( .C1(n16109), .C2(n20007), .A(n16047), .B(n16046), .ZN(
        P1_U2985) );
  AOI22_X1 U19254 ( .A1(n20168), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20167), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16053) );
  OAI22_X1 U19255 ( .A1(n16050), .A2(n16049), .B1(n20178), .B2(n16048), .ZN(
        n16051) );
  INV_X1 U19256 ( .A(n16051), .ZN(n16052) );
  OAI211_X1 U19257 ( .C1(n16054), .C2(n20007), .A(n16053), .B(n16052), .ZN(
        P1_U2987) );
  AOI22_X1 U19258 ( .A1(n20168), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20167), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16060) );
  NOR3_X1 U19259 ( .A1(n9643), .A2(n12224), .A3(n16133), .ZN(n16056) );
  NOR2_X1 U19260 ( .A1(n16056), .A2(n16055), .ZN(n16057) );
  XNOR2_X1 U19261 ( .A(n16057), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16121) );
  AOI22_X1 U19262 ( .A1(n16121), .A2(n20174), .B1(n20239), .B2(n16058), .ZN(
        n16059) );
  OAI211_X1 U19263 ( .C1(n20178), .C2(n16061), .A(n16060), .B(n16059), .ZN(
        P1_U2988) );
  AOI22_X1 U19264 ( .A1(n20168), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20167), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16066) );
  XNOR2_X1 U19265 ( .A(n16062), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16063) );
  XNOR2_X1 U19266 ( .A(n16064), .B(n16063), .ZN(n16154) );
  AOI22_X1 U19267 ( .A1(n16154), .A2(n20174), .B1(n20239), .B2(n20046), .ZN(
        n16065) );
  OAI211_X1 U19268 ( .C1(n20178), .C2(n20049), .A(n16066), .B(n16065), .ZN(
        P1_U2992) );
  AOI22_X1 U19269 ( .A1(n20168), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20167), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16072) );
  OAI21_X1 U19270 ( .B1(n16069), .B2(n16068), .A(n16067), .ZN(n16070) );
  INV_X1 U19271 ( .A(n16070), .ZN(n16161) );
  AOI22_X1 U19272 ( .A1(n16161), .A2(n20174), .B1(n20239), .B2(n20059), .ZN(
        n16071) );
  OAI211_X1 U19273 ( .C1(n20178), .C2(n20062), .A(n16072), .B(n16071), .ZN(
        P1_U2993) );
  AOI22_X1 U19274 ( .A1(n20168), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20167), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16079) );
  OAI21_X1 U19275 ( .B1(n16075), .B2(n16074), .A(n16073), .ZN(n16076) );
  INV_X1 U19276 ( .A(n16076), .ZN(n16166) );
  INV_X1 U19277 ( .A(n16077), .ZN(n20071) );
  AOI22_X1 U19278 ( .A1(n16166), .A2(n20174), .B1(n20239), .B2(n20071), .ZN(
        n16078) );
  OAI211_X1 U19279 ( .C1(n20178), .C2(n20074), .A(n16079), .B(n16078), .ZN(
        P1_U2994) );
  INV_X1 U19280 ( .A(n16106), .ZN(n16091) );
  INV_X1 U19281 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16081) );
  NAND2_X1 U19282 ( .A1(n16091), .A2(n16081), .ZN(n16089) );
  AND2_X1 U19283 ( .A1(n20220), .A2(n16090), .ZN(n16080) );
  NOR2_X1 U19284 ( .A1(n16100), .A2(n16080), .ZN(n16099) );
  NOR2_X1 U19285 ( .A1(n16099), .A2(n16081), .ZN(n16085) );
  AND3_X1 U19286 ( .A1(n16083), .A2(n16082), .A3(n20206), .ZN(n16084) );
  AOI211_X1 U19287 ( .C1(n20228), .C2(n16086), .A(n16085), .B(n16084), .ZN(
        n16088) );
  NAND2_X1 U19288 ( .A1(n20167), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n16087) );
  OAI211_X1 U19289 ( .C1(n16090), .C2(n16089), .A(n16088), .B(n16087), .ZN(
        P1_U3013) );
  AOI21_X1 U19290 ( .B1(n16092), .B2(n16091), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16098) );
  INV_X1 U19291 ( .A(n16093), .ZN(n16095) );
  AOI22_X1 U19292 ( .A1(n16095), .A2(n20206), .B1(n20228), .B2(n16094), .ZN(
        n16097) );
  NAND2_X1 U19293 ( .A1(n20167), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16096) );
  OAI211_X1 U19294 ( .C1(n16099), .C2(n16098), .A(n16097), .B(n16096), .ZN(
        P1_U3014) );
  AOI22_X1 U19295 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16100), .B1(
        n20167), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16105) );
  INV_X1 U19296 ( .A(n16101), .ZN(n16103) );
  AOI22_X1 U19297 ( .A1(n16103), .A2(n20206), .B1(n20228), .B2(n16102), .ZN(
        n16104) );
  OAI211_X1 U19298 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16106), .A(
        n16105), .B(n16104), .ZN(P1_U3016) );
  NOR4_X1 U19299 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n12230), .A3(
        n16107), .A4(n16164), .ZN(n16111) );
  OAI22_X1 U19300 ( .A1(n16109), .A2(n20222), .B1(n20182), .B2(n16108), .ZN(
        n16110) );
  NOR2_X1 U19301 ( .A1(n16111), .A2(n16110), .ZN(n16113) );
  NAND2_X1 U19302 ( .A1(n20167), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n16112) );
  OAI211_X1 U19303 ( .C1(n16115), .C2(n16114), .A(n16113), .B(n16112), .ZN(
        P1_U3017) );
  NAND2_X1 U19304 ( .A1(n16117), .A2(n16116), .ZN(n16124) );
  OAI22_X1 U19305 ( .A1(n16118), .A2(n20182), .B1(n20225), .B2(n16028), .ZN(
        n16119) );
  INV_X1 U19306 ( .A(n16119), .ZN(n16123) );
  AOI22_X1 U19307 ( .A1(n16121), .A2(n20206), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16120), .ZN(n16122) );
  OAI211_X1 U19308 ( .C1(n16164), .C2(n16124), .A(n16123), .B(n16122), .ZN(
        P1_U3020) );
  NAND2_X1 U19309 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16125) );
  AOI21_X1 U19310 ( .B1(n16142), .B2(n16125), .A(n20214), .ZN(n20179) );
  OAI21_X1 U19311 ( .B1(n16126), .B2(n20210), .A(n20179), .ZN(n16141) );
  AOI221_X1 U19312 ( .B1(n16130), .B2(n20220), .C1(n16127), .C2(n20220), .A(
        n16141), .ZN(n16140) );
  AOI222_X1 U19313 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n20167), .B1(n20228), 
        .B2(n16129), .C1(n16128), .C2(n20206), .ZN(n16132) );
  NOR2_X1 U19314 ( .A1(n16130), .A2(n16164), .ZN(n16135) );
  OAI221_X1 U19315 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n16133), .C2(n16139), .A(
        n16135), .ZN(n16131) );
  OAI211_X1 U19316 ( .C1(n16140), .C2(n16133), .A(n16132), .B(n16131), .ZN(
        P1_U3021) );
  AOI21_X1 U19317 ( .B1(n20024), .B2(n20228), .A(n16134), .ZN(n16138) );
  AOI22_X1 U19318 ( .A1(n16136), .A2(n20206), .B1(n16135), .B2(n16139), .ZN(
        n16137) );
  OAI211_X1 U19319 ( .C1(n16140), .C2(n16139), .A(n16138), .B(n16137), .ZN(
        P1_U3022) );
  NOR2_X1 U19320 ( .A1(n20185), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16165) );
  INV_X1 U19321 ( .A(n16165), .ZN(n16143) );
  AOI21_X1 U19322 ( .B1(n16142), .B2(n20185), .A(n16141), .ZN(n16170) );
  OAI21_X1 U19323 ( .B1(n16144), .B2(n16143), .A(n16170), .ZN(n16160) );
  AOI21_X1 U19324 ( .B1(n16148), .B2(n20220), .A(n16160), .ZN(n16158) );
  OAI22_X1 U19325 ( .A1(n20182), .A2(n16145), .B1(n20866), .B2(n20225), .ZN(
        n16146) );
  AOI21_X1 U19326 ( .B1(n16147), .B2(n20206), .A(n16146), .ZN(n16150) );
  NOR2_X1 U19327 ( .A1(n16148), .A2(n16164), .ZN(n16153) );
  OAI221_X1 U19328 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16151), .C2(n16157), .A(
        n16153), .ZN(n16149) );
  OAI211_X1 U19329 ( .C1(n16158), .C2(n16151), .A(n16150), .B(n16149), .ZN(
        P1_U3023) );
  INV_X1 U19330 ( .A(n16152), .ZN(n20035) );
  AOI22_X1 U19331 ( .A1(n20035), .A2(n20228), .B1(n20167), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16156) );
  AOI22_X1 U19332 ( .A1(n16154), .A2(n20206), .B1(n16157), .B2(n16153), .ZN(
        n16155) );
  OAI211_X1 U19333 ( .C1(n16158), .C2(n16157), .A(n16156), .B(n16155), .ZN(
        P1_U3024) );
  INV_X1 U19334 ( .A(n16159), .ZN(n20053) );
  AOI22_X1 U19335 ( .A1(n20053), .A2(n20228), .B1(n20167), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16163) );
  AOI22_X1 U19336 ( .A1(n16161), .A2(n20206), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16160), .ZN(n16162) );
  OAI211_X1 U19337 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16164), .A(
        n16163), .B(n16162), .ZN(P1_U3025) );
  AOI22_X1 U19338 ( .A1(n20063), .A2(n20228), .B1(n20167), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n16168) );
  AOI22_X1 U19339 ( .A1(n16166), .A2(n20206), .B1(n16165), .B2(n20193), .ZN(
        n16167) );
  OAI211_X1 U19340 ( .C1(n16170), .C2(n16169), .A(n16168), .B(n16167), .ZN(
        P1_U3026) );
  NAND3_X1 U19341 ( .A1(n16173), .A2(n16172), .A3(n16171), .ZN(n16174) );
  OAI21_X1 U19342 ( .B1(n16176), .B2(n16175), .A(n16174), .ZN(P1_U3468) );
  OAI221_X1 U19343 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n20914), .C2(n20918), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n20838) );
  NAND2_X1 U19344 ( .A1(n16177), .A2(n20838), .ZN(n16178) );
  AOI22_X1 U19345 ( .A1(n16181), .A2(n16180), .B1(n16179), .B2(n16178), .ZN(
        P1_U3162) );
  OAI21_X1 U19346 ( .B1(n20836), .B2(n20525), .A(n16182), .ZN(P1_U3466) );
  INV_X1 U19347 ( .A(n16183), .ZN(n16184) );
  AOI22_X1 U19348 ( .A1(n16184), .A2(n19131), .B1(P2_REIP_REG_31__SCAN_IN), 
        .B2(n19076), .ZN(n16192) );
  AOI22_X1 U19349 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n19142), .B1(
        P2_EBX_REG_31__SCAN_IN), .B2(n16185), .ZN(n16191) );
  AOI22_X1 U19350 ( .A1(n19148), .A2(n19129), .B1(n19122), .B2(n16186), .ZN(
        n16190) );
  NAND4_X1 U19351 ( .A1(n19123), .A2(n16188), .A3(n16187), .A4(n12794), .ZN(
        n16189) );
  NAND4_X1 U19352 ( .A1(n16192), .A2(n16191), .A3(n16190), .A4(n16189), .ZN(
        P2_U2824) );
  AOI22_X1 U19353 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n19135), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19142), .ZN(n16195) );
  OAI21_X1 U19354 ( .B1(n19133), .B2(n19913), .A(n16195), .ZN(n16196) );
  AOI21_X1 U19355 ( .B1(n16197), .B2(n19131), .A(n16196), .ZN(n16198) );
  OAI21_X1 U19356 ( .B1(n16199), .B2(n19137), .A(n16198), .ZN(n16200) );
  AOI21_X1 U19357 ( .B1(n16193), .B2(n16201), .A(n16200), .ZN(n16202) );
  OAI21_X1 U19358 ( .B1(n16203), .B2(n19127), .A(n16202), .ZN(P2_U2826) );
  NOR2_X1 U19359 ( .A1(n19133), .A2(n19907), .ZN(n16204) );
  AOI21_X1 U19360 ( .B1(n16205), .B2(n19131), .A(n16204), .ZN(n16215) );
  AOI22_X1 U19361 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n19135), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19142), .ZN(n16214) );
  INV_X1 U19362 ( .A(n16206), .ZN(n16208) );
  AOI22_X1 U19363 ( .A1(n16208), .A2(n19129), .B1(n19122), .B2(n16207), .ZN(
        n16213) );
  AOI21_X1 U19364 ( .B1(n16210), .B2(n9678), .A(n16209), .ZN(n16211) );
  NAND2_X1 U19365 ( .A1(n19123), .A2(n16211), .ZN(n16212) );
  NAND4_X1 U19366 ( .A1(n16215), .A2(n16214), .A3(n16213), .A4(n16212), .ZN(
        P2_U2829) );
  INV_X1 U19367 ( .A(n16216), .ZN(n16217) );
  AOI22_X1 U19368 ( .A1(n16217), .A2(n19131), .B1(P2_REIP_REG_24__SCAN_IN), 
        .B2(n19076), .ZN(n16228) );
  AOI22_X1 U19369 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n19135), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19142), .ZN(n16227) );
  OAI22_X1 U19370 ( .A1(n16219), .A2(n19127), .B1(n19137), .B2(n16218), .ZN(
        n16220) );
  INV_X1 U19371 ( .A(n16220), .ZN(n16226) );
  INV_X1 U19372 ( .A(n16221), .ZN(n16222) );
  AOI21_X1 U19373 ( .B1(n16223), .B2(n16222), .A(n9679), .ZN(n16224) );
  NAND2_X1 U19374 ( .A1(n19123), .A2(n16224), .ZN(n16225) );
  NAND4_X1 U19375 ( .A1(n16228), .A2(n16227), .A3(n16226), .A4(n16225), .ZN(
        P2_U2831) );
  AOI22_X1 U19376 ( .A1(n16235), .A2(n16229), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19188), .ZN(n16233) );
  AOI22_X1 U19377 ( .A1(n19147), .A2(BUF2_REG_20__SCAN_IN), .B1(n19149), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16232) );
  AOI22_X1 U19378 ( .A1(n18990), .A2(n19189), .B1(n19191), .B2(n16230), .ZN(
        n16231) );
  NAND3_X1 U19379 ( .A1(n16233), .A2(n16232), .A3(n16231), .ZN(P2_U2899) );
  AOI22_X1 U19380 ( .A1(n16235), .A2(n16234), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19188), .ZN(n16242) );
  AOI22_X1 U19381 ( .A1(n19147), .A2(BUF2_REG_18__SCAN_IN), .B1(n19149), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16241) );
  OAI22_X1 U19382 ( .A1(n16238), .A2(n16237), .B1(n19183), .B2(n16236), .ZN(
        n16239) );
  INV_X1 U19383 ( .A(n16239), .ZN(n16240) );
  NAND3_X1 U19384 ( .A1(n16242), .A2(n16241), .A3(n16240), .ZN(P2_U2901) );
  AOI22_X1 U19385 ( .A1(n19231), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n11988), .ZN(n16246) );
  AOI222_X1 U19386 ( .A1(n16244), .A2(n16297), .B1(n19236), .B2(n16243), .C1(
        n16306), .C2(n19044), .ZN(n16245) );
  OAI211_X1 U19387 ( .C1(n19240), .C2(n19038), .A(n16246), .B(n16245), .ZN(
        P2_U3000) );
  AOI22_X1 U19388 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n15544), .B1(n16301), 
        .B2(n19051), .ZN(n16252) );
  OAI22_X1 U19389 ( .A1(n16248), .A2(n11993), .B1(n16303), .B2(n16247), .ZN(
        n16249) );
  AOI21_X1 U19390 ( .B1(n16306), .B2(n16250), .A(n16249), .ZN(n16251) );
  OAI211_X1 U19391 ( .C1(n16310), .C2(n16253), .A(n16252), .B(n16251), .ZN(
        P2_U3001) );
  AOI22_X1 U19392 ( .A1(n19231), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n11988), .ZN(n16261) );
  NAND2_X1 U19393 ( .A1(n16254), .A2(n19236), .ZN(n16256) );
  OAI22_X1 U19394 ( .A1(n16257), .A2(n16256), .B1(n13736), .B2(n16255), .ZN(
        n16258) );
  AOI21_X1 U19395 ( .B1(n16259), .B2(n16297), .A(n16258), .ZN(n16260) );
  OAI211_X1 U19396 ( .C1(n19240), .C2(n19061), .A(n16261), .B(n16260), .ZN(
        P2_U3002) );
  AOI22_X1 U19397 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n11988), .B1(n16301), 
        .B2(n19084), .ZN(n16266) );
  OAI22_X1 U19398 ( .A1(n16263), .A2(n11993), .B1(n16303), .B2(n16262), .ZN(
        n16264) );
  AOI21_X1 U19399 ( .B1(n16306), .B2(n10163), .A(n16264), .ZN(n16265) );
  OAI211_X1 U19400 ( .C1(n16310), .C2(n19074), .A(n16266), .B(n16265), .ZN(
        P2_U3003) );
  AOI22_X1 U19401 ( .A1(n19231), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n11988), .ZN(n16276) );
  NAND2_X1 U19402 ( .A1(n16267), .A2(n16268), .ZN(n16271) );
  NOR2_X1 U19403 ( .A1(n16269), .A2(n10174), .ZN(n16270) );
  XNOR2_X1 U19404 ( .A(n16271), .B(n16270), .ZN(n16321) );
  INV_X1 U19405 ( .A(n16321), .ZN(n16274) );
  NAND2_X1 U19406 ( .A1(n15554), .A2(n11883), .ZN(n16272) );
  AOI222_X1 U19407 ( .A1(n16274), .A2(n16297), .B1(n16306), .B2(n16316), .C1(
        n19236), .C2(n16317), .ZN(n16275) );
  OAI211_X1 U19408 ( .C1(n19240), .C2(n16277), .A(n16276), .B(n16275), .ZN(
        P2_U3004) );
  AOI22_X1 U19409 ( .A1(n19231), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n11988), .ZN(n16292) );
  NOR2_X1 U19410 ( .A1(n16279), .A2(n16278), .ZN(n16283) );
  NOR2_X1 U19411 ( .A1(n16281), .A2(n16280), .ZN(n16282) );
  XNOR2_X1 U19412 ( .A(n16283), .B(n16282), .ZN(n16333) );
  NAND2_X1 U19413 ( .A1(n16285), .A2(n16284), .ZN(n16290) );
  AOI21_X1 U19414 ( .B1(n16288), .B2(n16287), .A(n16286), .ZN(n16289) );
  XOR2_X1 U19415 ( .A(n16290), .B(n16289), .Z(n16329) );
  AOI222_X1 U19416 ( .A1(n16333), .A2(n16297), .B1(n16306), .B2(n16330), .C1(
        n16329), .C2(n19236), .ZN(n16291) );
  OAI211_X1 U19417 ( .C1(n19240), .C2(n16293), .A(n16292), .B(n16291), .ZN(
        P2_U3006) );
  AOI22_X1 U19418 ( .A1(n19231), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n11988), .ZN(n16300) );
  OAI22_X1 U19419 ( .A1(n16295), .A2(n16303), .B1(n13736), .B2(n16294), .ZN(
        n16296) );
  AOI21_X1 U19420 ( .B1(n16298), .B2(n16297), .A(n16296), .ZN(n16299) );
  OAI211_X1 U19421 ( .C1(n19240), .C2(n19106), .A(n16300), .B(n16299), .ZN(
        P2_U3008) );
  AOI22_X1 U19422 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n11988), .B1(n16301), 
        .B2(n19120), .ZN(n16308) );
  OAI22_X1 U19423 ( .A1(n16304), .A2(n11993), .B1(n16303), .B2(n16302), .ZN(
        n16305) );
  AOI21_X1 U19424 ( .B1(n16306), .B2(n19121), .A(n16305), .ZN(n16307) );
  OAI211_X1 U19425 ( .C1(n16310), .C2(n16309), .A(n16308), .B(n16307), .ZN(
        P2_U3009) );
  NAND2_X1 U19426 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16311), .ZN(
        n16314) );
  NAND2_X1 U19427 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n15544), .ZN(n16312) );
  OAI221_X1 U19428 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16314), 
        .C1(n11883), .C2(n16313), .A(n16312), .ZN(n16315) );
  AOI21_X1 U19429 ( .B1(n16324), .B2(n19158), .A(n16315), .ZN(n16319) );
  AOI22_X1 U19430 ( .A1(n16317), .A2(n16328), .B1(n16331), .B2(n16316), .ZN(
        n16318) );
  OAI211_X1 U19431 ( .C1(n16321), .C2(n16320), .A(n16319), .B(n16318), .ZN(
        P2_U3036) );
  AOI221_X1 U19432 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C1(n16323), .C2(n16336), .A(
        n16322), .ZN(n16327) );
  NAND2_X1 U19433 ( .A1(n16324), .A2(n19162), .ZN(n16325) );
  OAI21_X1 U19434 ( .B1(n13590), .B2(n19113), .A(n16325), .ZN(n16326) );
  NOR2_X1 U19435 ( .A1(n16327), .A2(n16326), .ZN(n16335) );
  AOI222_X1 U19436 ( .A1(n16333), .A2(n16332), .B1(n16331), .B2(n16330), .C1(
        n16329), .C2(n16328), .ZN(n16334) );
  OAI211_X1 U19437 ( .C1(n16337), .C2(n16336), .A(n16335), .B(n16334), .ZN(
        P2_U3038) );
  INV_X1 U19438 ( .A(n16374), .ZN(n16346) );
  NAND2_X1 U19439 ( .A1(n16351), .A2(n16346), .ZN(n16340) );
  NAND2_X1 U19440 ( .A1(n16374), .A2(n16338), .ZN(n16339) );
  NAND2_X1 U19441 ( .A1(n16340), .A2(n16339), .ZN(n16377) );
  NAND2_X1 U19442 ( .A1(n16343), .A2(n19956), .ZN(n16342) );
  NAND3_X1 U19443 ( .A1(n16342), .A2(n16341), .A3(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n16345) );
  OR2_X1 U19444 ( .A1(n16343), .A2(n19956), .ZN(n16344) );
  NAND2_X1 U19445 ( .A1(n16345), .A2(n16344), .ZN(n16350) );
  NAND2_X1 U19446 ( .A1(n16350), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n16347) );
  NAND3_X1 U19447 ( .A1(n16347), .A2(n16346), .A3(n16356), .ZN(n16348) );
  NAND2_X1 U19448 ( .A1(n16377), .A2(n16348), .ZN(n16349) );
  NAND2_X1 U19449 ( .A1(n16349), .A2(n19938), .ZN(n16354) );
  AOI211_X1 U19450 ( .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n16351), .A(
        n16374), .B(n16350), .ZN(n16352) );
  NAND2_X1 U19451 ( .A1(n16352), .A2(n19946), .ZN(n16353) );
  NAND2_X1 U19452 ( .A1(n16354), .A2(n16353), .ZN(n16379) );
  NAND2_X1 U19453 ( .A1(n16374), .A2(n11223), .ZN(n16355) );
  OAI21_X1 U19454 ( .B1(n16356), .B2(n16374), .A(n16355), .ZN(n16376) );
  INV_X1 U19455 ( .A(n12509), .ZN(n16358) );
  NAND2_X1 U19456 ( .A1(n16358), .A2(n16357), .ZN(n16361) );
  NAND2_X1 U19457 ( .A1(n16363), .A2(n16359), .ZN(n16360) );
  OAI211_X1 U19458 ( .C1(n16363), .C2(n16362), .A(n16361), .B(n16360), .ZN(
        n19975) );
  NOR2_X1 U19459 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n16370) );
  INV_X1 U19460 ( .A(n16364), .ZN(n16365) );
  NAND2_X1 U19461 ( .A1(n11551), .A2(n16365), .ZN(n16367) );
  OAI22_X1 U19462 ( .A1(n12265), .A2(n16367), .B1(n16366), .B2(n11397), .ZN(
        n16368) );
  INV_X1 U19463 ( .A(n16368), .ZN(n16369) );
  OAI21_X1 U19464 ( .B1(n16371), .B2(n16370), .A(n16369), .ZN(n16372) );
  OR2_X1 U19465 ( .A1(n19975), .A2(n16372), .ZN(n16373) );
  AOI21_X1 U19466 ( .B1(n16374), .B2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16373), .ZN(n16375) );
  OAI21_X1 U19467 ( .B1(n16377), .B2(n16376), .A(n16375), .ZN(n16378) );
  AOI21_X1 U19468 ( .B1(n16379), .B2(n15986), .A(n16378), .ZN(n16394) );
  AOI211_X1 U19469 ( .C1(n19968), .C2(n16382), .A(n16381), .B(n16380), .ZN(
        n16393) );
  NAND2_X1 U19470 ( .A1(n16394), .A2(n11444), .ZN(n16383) );
  NAND2_X1 U19471 ( .A1(n16383), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16387) );
  NAND2_X1 U19472 ( .A1(n19979), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16384) );
  AOI21_X1 U19473 ( .B1(n16386), .B2(n16385), .A(n16384), .ZN(n16390) );
  AND2_X1 U19474 ( .A1(n16387), .A2(n16390), .ZN(n16395) );
  AOI21_X1 U19475 ( .B1(n16388), .B2(n19987), .A(n19984), .ZN(n16389) );
  AOI21_X1 U19476 ( .B1(n16390), .B2(n19867), .A(n16389), .ZN(n16391) );
  AOI21_X1 U19477 ( .B1(n16395), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16391), 
        .ZN(n16392) );
  OAI211_X1 U19478 ( .C1(n16394), .C2(n19845), .A(n16393), .B(n16392), .ZN(
        P2_U3176) );
  OAI221_X1 U19479 ( .B1(n19645), .B2(P2_STATE2_REG_0__SCAN_IN), .C1(n19645), 
        .C2(n19848), .A(n16396), .ZN(P2_U3593) );
  NAND2_X1 U19480 ( .A1(n17828), .A2(n16397), .ZN(n16420) );
  NAND2_X1 U19481 ( .A1(n17902), .A2(n16398), .ZN(n16408) );
  AOI21_X1 U19482 ( .B1(n16420), .B2(n16408), .A(n16422), .ZN(n16403) );
  OAI221_X1 U19483 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16401), .C1(
        n9893), .C2(n16400), .A(n16399), .ZN(n16402) );
  AOI211_X1 U19484 ( .C1(n17770), .C2(n16574), .A(n16403), .B(n16402), .ZN(
        n16406) );
  NAND3_X1 U19485 ( .A1(n16404), .A2(n17571), .A3(n16422), .ZN(n16405) );
  OAI211_X1 U19486 ( .C1(n16407), .C2(n17831), .A(n16406), .B(n16405), .ZN(
        P3_U2800) );
  AOI21_X1 U19487 ( .B1(n16439), .B2(n16419), .A(n16408), .ZN(n16416) );
  AOI22_X1 U19488 ( .A1(n18071), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16409), .ZN(n16412) );
  OAI21_X1 U19489 ( .B1(n16410), .B2(n17770), .A(n16587), .ZN(n16411) );
  OAI211_X1 U19490 ( .C1(n16414), .C2(n16413), .A(n16412), .B(n16411), .ZN(
        n16415) );
  AOI211_X1 U19491 ( .C1(n17810), .C2(n16417), .A(n16416), .B(n16415), .ZN(
        n16418) );
  OAI221_X1 U19492 ( .B1(n16420), .B2(n16419), .C1(n16420), .C2(n16438), .A(
        n16418), .ZN(P3_U2801) );
  INV_X1 U19493 ( .A(n18234), .ZN(n18160) );
  AOI21_X1 U19494 ( .B1(n18160), .B2(n16422), .A(n16421), .ZN(n16425) );
  OAI22_X1 U19495 ( .A1(n16425), .A2(n18891), .B1(n16424), .B2(n16423), .ZN(
        n16426) );
  AOI211_X1 U19496 ( .C1(n18166), .C2(n16428), .A(n16427), .B(n16426), .ZN(
        n16431) );
  NAND2_X1 U19497 ( .A1(n18246), .A2(n16429), .ZN(n16430) );
  OAI211_X1 U19498 ( .C1(n16432), .C2(n18170), .A(n16431), .B(n16430), .ZN(
        P3_U2831) );
  NAND2_X1 U19499 ( .A1(n17558), .A2(n17572), .ZN(n16450) );
  AOI21_X1 U19500 ( .B1(n10022), .B2(n17574), .A(n17572), .ZN(n17557) );
  INV_X1 U19501 ( .A(n17556), .ZN(n16436) );
  INV_X1 U19502 ( .A(n18138), .ZN(n18050) );
  OR2_X1 U19503 ( .A1(n16434), .A2(n10153), .ZN(n16435) );
  NOR2_X1 U19504 ( .A1(n18757), .A2(n16437), .ZN(n18101) );
  AOI22_X1 U19505 ( .A1(n18750), .A2(n16439), .B1(n18101), .B2(n16438), .ZN(
        n16440) );
  NAND2_X1 U19506 ( .A1(n16441), .A2(n16440), .ZN(n16446) );
  INV_X1 U19507 ( .A(n18101), .ZN(n18120) );
  OAI22_X1 U19508 ( .A1(n18123), .A2(n18097), .B1(n17782), .B2(n18120), .ZN(
        n18030) );
  OAI21_X1 U19509 ( .B1(n18128), .B2(n18251), .A(n18740), .ZN(n18218) );
  NOR3_X1 U19510 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17918), .A3(
        n17917), .ZN(n17561) );
  NOR2_X1 U19511 ( .A1(n18140), .A2(n18866), .ZN(n17553) );
  INV_X1 U19512 ( .A(n16443), .ZN(n16444) );
  AOI21_X1 U19513 ( .B1(n16446), .B2(n16445), .A(n16444), .ZN(n16449) );
  NAND3_X1 U19514 ( .A1(n16447), .A2(n18248), .A3(n17557), .ZN(n16448) );
  OAI211_X1 U19515 ( .C1(n18170), .C2(n16450), .A(n16449), .B(n16448), .ZN(
        P3_U2834) );
  NOR3_X1 U19516 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16452) );
  NOR4_X1 U19517 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16451) );
  INV_X2 U19518 ( .A(n16539), .ZN(U215) );
  NAND4_X1 U19519 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16452), .A3(n16451), .A4(
        U215), .ZN(U213) );
  INV_X1 U19520 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16542) );
  INV_X1 U19521 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16541) );
  OAI222_X1 U19522 ( .A1(U212), .A2(n16542), .B1(n16503), .B2(n20287), .C1(
        U214), .C2(n16541), .ZN(U216) );
  INV_X2 U19523 ( .A(U212), .ZN(n16501) );
  AOI22_X1 U19524 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n16500), .ZN(n16454) );
  OAI21_X1 U19525 ( .B1(n14783), .B2(n16503), .A(n16454), .ZN(U217) );
  AOI22_X1 U19526 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16500), .ZN(n16455) );
  OAI21_X1 U19527 ( .B1(n15317), .B2(n16503), .A(n16455), .ZN(U218) );
  AOI22_X1 U19528 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16500), .ZN(n16456) );
  OAI21_X1 U19529 ( .B1(n15322), .B2(n16503), .A(n16456), .ZN(U219) );
  AOI22_X1 U19530 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16500), .ZN(n16457) );
  OAI21_X1 U19531 ( .B1(n15329), .B2(n16503), .A(n16457), .ZN(U220) );
  INV_X1 U19532 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20262) );
  AOI22_X1 U19533 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16500), .ZN(n16458) );
  OAI21_X1 U19534 ( .B1(n20262), .B2(n16503), .A(n16458), .ZN(U221) );
  AOI22_X1 U19535 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16500), .ZN(n16459) );
  OAI21_X1 U19536 ( .B1(n15345), .B2(n16503), .A(n16459), .ZN(U222) );
  INV_X1 U19537 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16461) );
  AOI22_X1 U19538 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16500), .ZN(n16460) );
  OAI21_X1 U19539 ( .B1(n16461), .B2(n16503), .A(n16460), .ZN(U223) );
  INV_X1 U19540 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16463) );
  AOI22_X1 U19541 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16500), .ZN(n16462) );
  OAI21_X1 U19542 ( .B1(n16463), .B2(n16503), .A(n16462), .ZN(U224) );
  INV_X1 U19543 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20279) );
  AOI22_X1 U19544 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16500), .ZN(n16464) );
  OAI21_X1 U19545 ( .B1(n20279), .B2(n16503), .A(n16464), .ZN(U225) );
  INV_X1 U19546 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16466) );
  AOI22_X1 U19547 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16500), .ZN(n16465) );
  OAI21_X1 U19548 ( .B1(n16466), .B2(n16503), .A(n16465), .ZN(U226) );
  AOI22_X1 U19549 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16500), .ZN(n16467) );
  OAI21_X1 U19550 ( .B1(n14822), .B2(n16503), .A(n16467), .ZN(U227) );
  INV_X1 U19551 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16469) );
  AOI22_X1 U19552 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16500), .ZN(n16468) );
  OAI21_X1 U19553 ( .B1(n16469), .B2(n16503), .A(n16468), .ZN(U228) );
  INV_X1 U19554 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16471) );
  AOI22_X1 U19555 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16500), .ZN(n16470) );
  OAI21_X1 U19556 ( .B1(n16471), .B2(n16503), .A(n16470), .ZN(U229) );
  INV_X1 U19557 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20257) );
  AOI22_X1 U19558 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16500), .ZN(n16472) );
  OAI21_X1 U19559 ( .B1(n20257), .B2(n16503), .A(n16472), .ZN(U230) );
  INV_X1 U19560 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16474) );
  AOI22_X1 U19561 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16500), .ZN(n16473) );
  OAI21_X1 U19562 ( .B1(n16474), .B2(n16503), .A(n16473), .ZN(U231) );
  AOI22_X1 U19563 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16500), .ZN(n16475) );
  OAI21_X1 U19564 ( .B1(n13249), .B2(n16503), .A(n16475), .ZN(U232) );
  AOI22_X1 U19565 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16500), .ZN(n16476) );
  OAI21_X1 U19566 ( .B1(n12991), .B2(n16503), .A(n16476), .ZN(U233) );
  AOI22_X1 U19567 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16500), .ZN(n16477) );
  OAI21_X1 U19568 ( .B1(n16478), .B2(n16503), .A(n16477), .ZN(U234) );
  AOI22_X1 U19569 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16500), .ZN(n16479) );
  OAI21_X1 U19570 ( .B1(n16480), .B2(n16503), .A(n16479), .ZN(U235) );
  AOI22_X1 U19571 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16500), .ZN(n16481) );
  OAI21_X1 U19572 ( .B1(n16482), .B2(n16503), .A(n16481), .ZN(U236) );
  AOI22_X1 U19573 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16500), .ZN(n16483) );
  OAI21_X1 U19574 ( .B1(n16484), .B2(n16503), .A(n16483), .ZN(U237) );
  AOI22_X1 U19575 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16500), .ZN(n16485) );
  OAI21_X1 U19576 ( .B1(n16486), .B2(n16503), .A(n16485), .ZN(U238) );
  AOI22_X1 U19577 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16500), .ZN(n16487) );
  OAI21_X1 U19578 ( .B1(n16488), .B2(n16503), .A(n16487), .ZN(U239) );
  AOI22_X1 U19579 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16500), .ZN(n16489) );
  OAI21_X1 U19580 ( .B1(n13396), .B2(n16503), .A(n16489), .ZN(U240) );
  AOI22_X1 U19581 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16500), .ZN(n16490) );
  OAI21_X1 U19582 ( .B1(n13390), .B2(n16503), .A(n16490), .ZN(U241) );
  AOI22_X1 U19583 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16500), .ZN(n16491) );
  OAI21_X1 U19584 ( .B1(n13400), .B2(n16503), .A(n16491), .ZN(U242) );
  INV_X1 U19585 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16493) );
  AOI22_X1 U19586 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16500), .ZN(n16492) );
  OAI21_X1 U19587 ( .B1(n16493), .B2(n16503), .A(n16492), .ZN(U243) );
  INV_X1 U19588 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16495) );
  AOI22_X1 U19589 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16500), .ZN(n16494) );
  OAI21_X1 U19590 ( .B1(n16495), .B2(n16503), .A(n16494), .ZN(U244) );
  INV_X1 U19591 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16497) );
  AOI22_X1 U19592 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16500), .ZN(n16496) );
  OAI21_X1 U19593 ( .B1(n16497), .B2(n16503), .A(n16496), .ZN(U245) );
  INV_X1 U19594 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16499) );
  AOI22_X1 U19595 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16500), .ZN(n16498) );
  OAI21_X1 U19596 ( .B1(n16499), .B2(n16503), .A(n16498), .ZN(U246) );
  INV_X1 U19597 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16504) );
  AOI22_X1 U19598 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n16501), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16500), .ZN(n16502) );
  OAI21_X1 U19599 ( .B1(n16504), .B2(n16503), .A(n16502), .ZN(U247) );
  OAI22_X1 U19600 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16539), .ZN(n16505) );
  INV_X1 U19601 ( .A(n16505), .ZN(U251) );
  OAI22_X1 U19602 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16539), .ZN(n16506) );
  INV_X1 U19603 ( .A(n16506), .ZN(U252) );
  OAI22_X1 U19604 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16539), .ZN(n16507) );
  INV_X1 U19605 ( .A(n16507), .ZN(U253) );
  OAI22_X1 U19606 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16539), .ZN(n16508) );
  INV_X1 U19607 ( .A(n16508), .ZN(U254) );
  OAI22_X1 U19608 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16539), .ZN(n16509) );
  INV_X1 U19609 ( .A(n16509), .ZN(U255) );
  OAI22_X1 U19610 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16539), .ZN(n16510) );
  INV_X1 U19611 ( .A(n16510), .ZN(U256) );
  OAI22_X1 U19612 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16539), .ZN(n16511) );
  INV_X1 U19613 ( .A(n16511), .ZN(U257) );
  OAI22_X1 U19614 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16539), .ZN(n16512) );
  INV_X1 U19615 ( .A(n16512), .ZN(U258) );
  OAI22_X1 U19616 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16539), .ZN(n16513) );
  INV_X1 U19617 ( .A(n16513), .ZN(U259) );
  OAI22_X1 U19618 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16529), .ZN(n16514) );
  INV_X1 U19619 ( .A(n16514), .ZN(U260) );
  INV_X1 U19620 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16516) );
  INV_X1 U19621 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n16515) );
  AOI22_X1 U19622 ( .A1(n16539), .A2(n16516), .B1(n16515), .B2(U215), .ZN(U261) );
  OAI22_X1 U19623 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16529), .ZN(n16517) );
  INV_X1 U19624 ( .A(n16517), .ZN(U262) );
  OAI22_X1 U19625 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16539), .ZN(n16518) );
  INV_X1 U19626 ( .A(n16518), .ZN(U263) );
  OAI22_X1 U19627 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16529), .ZN(n16519) );
  INV_X1 U19628 ( .A(n16519), .ZN(U264) );
  OAI22_X1 U19629 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16539), .ZN(n16520) );
  INV_X1 U19630 ( .A(n16520), .ZN(U265) );
  OAI22_X1 U19631 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16539), .ZN(n16521) );
  INV_X1 U19632 ( .A(n16521), .ZN(U266) );
  OAI22_X1 U19633 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16529), .ZN(n16522) );
  INV_X1 U19634 ( .A(n16522), .ZN(U267) );
  OAI22_X1 U19635 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16529), .ZN(n16523) );
  INV_X1 U19636 ( .A(n16523), .ZN(U268) );
  OAI22_X1 U19637 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16529), .ZN(n16524) );
  INV_X1 U19638 ( .A(n16524), .ZN(U269) );
  OAI22_X1 U19639 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16529), .ZN(n16525) );
  INV_X1 U19640 ( .A(n16525), .ZN(U270) );
  OAI22_X1 U19641 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16529), .ZN(n16526) );
  INV_X1 U19642 ( .A(n16526), .ZN(U271) );
  OAI22_X1 U19643 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16529), .ZN(n16527) );
  INV_X1 U19644 ( .A(n16527), .ZN(U272) );
  OAI22_X1 U19645 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16539), .ZN(n16528) );
  INV_X1 U19646 ( .A(n16528), .ZN(U273) );
  OAI22_X1 U19647 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16529), .ZN(n16530) );
  INV_X1 U19648 ( .A(n16530), .ZN(U274) );
  OAI22_X1 U19649 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16539), .ZN(n16531) );
  INV_X1 U19650 ( .A(n16531), .ZN(U275) );
  OAI22_X1 U19651 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16539), .ZN(n16532) );
  INV_X1 U19652 ( .A(n16532), .ZN(U276) );
  OAI22_X1 U19653 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16539), .ZN(n16533) );
  INV_X1 U19654 ( .A(n16533), .ZN(U277) );
  OAI22_X1 U19655 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16539), .ZN(n16534) );
  INV_X1 U19656 ( .A(n16534), .ZN(U278) );
  OAI22_X1 U19657 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16539), .ZN(n16535) );
  INV_X1 U19658 ( .A(n16535), .ZN(U279) );
  OAI22_X1 U19659 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16539), .ZN(n16536) );
  INV_X1 U19660 ( .A(n16536), .ZN(U280) );
  OAI22_X1 U19661 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16539), .ZN(n16537) );
  INV_X1 U19662 ( .A(n16537), .ZN(U281) );
  INV_X1 U19663 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18298) );
  AOI22_X1 U19664 ( .A1(n16539), .A2(n16542), .B1(n18298), .B2(U215), .ZN(U282) );
  INV_X1 U19665 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16540) );
  AOI222_X1 U19666 ( .A1(n16542), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16541), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n16540), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16543) );
  INV_X2 U19667 ( .A(n16545), .ZN(n16544) );
  INV_X1 U19668 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18829) );
  INV_X1 U19669 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19883) );
  AOI22_X1 U19670 ( .A1(n16544), .A2(n18829), .B1(n19883), .B2(n16545), .ZN(
        U347) );
  INV_X1 U19671 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18827) );
  INV_X1 U19672 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19882) );
  AOI22_X1 U19673 ( .A1(n16544), .A2(n18827), .B1(n19882), .B2(n16545), .ZN(
        U348) );
  INV_X1 U19674 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18825) );
  INV_X1 U19675 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19881) );
  AOI22_X1 U19676 ( .A1(n16544), .A2(n18825), .B1(n19881), .B2(n16545), .ZN(
        U349) );
  INV_X1 U19677 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18823) );
  INV_X1 U19678 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19880) );
  AOI22_X1 U19679 ( .A1(n16544), .A2(n18823), .B1(n19880), .B2(n16545), .ZN(
        U350) );
  INV_X1 U19680 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18821) );
  INV_X1 U19681 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19878) );
  AOI22_X1 U19682 ( .A1(n16544), .A2(n18821), .B1(n19878), .B2(n16545), .ZN(
        U351) );
  INV_X1 U19683 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18819) );
  INV_X1 U19684 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19877) );
  AOI22_X1 U19685 ( .A1(n16544), .A2(n18819), .B1(n19877), .B2(n16545), .ZN(
        U352) );
  INV_X1 U19686 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18817) );
  INV_X1 U19687 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19876) );
  AOI22_X1 U19688 ( .A1(n16544), .A2(n18817), .B1(n19876), .B2(n16545), .ZN(
        U353) );
  INV_X1 U19689 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18815) );
  AOI22_X1 U19690 ( .A1(n16544), .A2(n18815), .B1(n19875), .B2(n16545), .ZN(
        U354) );
  INV_X1 U19691 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18868) );
  INV_X1 U19692 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19914) );
  AOI22_X1 U19693 ( .A1(n16544), .A2(n18868), .B1(n19914), .B2(n16545), .ZN(
        U356) );
  INV_X1 U19694 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18865) );
  INV_X1 U19695 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19912) );
  AOI22_X1 U19696 ( .A1(n16544), .A2(n18865), .B1(n19912), .B2(n16545), .ZN(
        U357) );
  INV_X1 U19697 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18864) );
  INV_X1 U19698 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19909) );
  AOI22_X1 U19699 ( .A1(n16544), .A2(n18864), .B1(n19909), .B2(n16545), .ZN(
        U358) );
  INV_X1 U19700 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18861) );
  INV_X1 U19701 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19908) );
  AOI22_X1 U19702 ( .A1(n16544), .A2(n18861), .B1(n19908), .B2(n16545), .ZN(
        U359) );
  INV_X1 U19703 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18859) );
  INV_X1 U19704 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19906) );
  AOI22_X1 U19705 ( .A1(n16544), .A2(n18859), .B1(n19906), .B2(n16545), .ZN(
        U360) );
  INV_X1 U19706 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18857) );
  INV_X1 U19707 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19904) );
  AOI22_X1 U19708 ( .A1(n16544), .A2(n18857), .B1(n19904), .B2(n16545), .ZN(
        U361) );
  INV_X1 U19709 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18855) );
  INV_X1 U19710 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19903) );
  AOI22_X1 U19711 ( .A1(n16544), .A2(n18855), .B1(n19903), .B2(n16545), .ZN(
        U362) );
  INV_X1 U19712 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18853) );
  INV_X1 U19713 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19901) );
  AOI22_X1 U19714 ( .A1(n16544), .A2(n18853), .B1(n19901), .B2(n16545), .ZN(
        U363) );
  INV_X1 U19715 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18851) );
  INV_X1 U19716 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19899) );
  AOI22_X1 U19717 ( .A1(n16544), .A2(n18851), .B1(n19899), .B2(n16545), .ZN(
        U364) );
  INV_X1 U19718 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18813) );
  INV_X1 U19719 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19874) );
  AOI22_X1 U19720 ( .A1(n16544), .A2(n18813), .B1(n19874), .B2(n16545), .ZN(
        U365) );
  INV_X1 U19721 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18848) );
  INV_X1 U19722 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19897) );
  AOI22_X1 U19723 ( .A1(n16544), .A2(n18848), .B1(n19897), .B2(n16545), .ZN(
        U366) );
  INV_X1 U19724 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18847) );
  INV_X1 U19725 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19896) );
  AOI22_X1 U19726 ( .A1(n16544), .A2(n18847), .B1(n19896), .B2(n16545), .ZN(
        U367) );
  INV_X1 U19727 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18845) );
  INV_X1 U19728 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19894) );
  AOI22_X1 U19729 ( .A1(n16544), .A2(n18845), .B1(n19894), .B2(n16545), .ZN(
        U368) );
  INV_X1 U19730 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18842) );
  INV_X1 U19731 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19893) );
  AOI22_X1 U19732 ( .A1(n16544), .A2(n18842), .B1(n19893), .B2(n16545), .ZN(
        U369) );
  INV_X1 U19733 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18841) );
  INV_X1 U19734 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19891) );
  AOI22_X1 U19735 ( .A1(n16544), .A2(n18841), .B1(n19891), .B2(n16545), .ZN(
        U370) );
  INV_X1 U19736 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18839) );
  INV_X1 U19737 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19889) );
  AOI22_X1 U19738 ( .A1(n16544), .A2(n18839), .B1(n19889), .B2(n16545), .ZN(
        U371) );
  INV_X1 U19739 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18836) );
  INV_X1 U19740 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19887) );
  AOI22_X1 U19741 ( .A1(n16544), .A2(n18836), .B1(n19887), .B2(n16545), .ZN(
        U372) );
  INV_X1 U19742 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18835) );
  INV_X1 U19743 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19886) );
  AOI22_X1 U19744 ( .A1(n16544), .A2(n18835), .B1(n19886), .B2(n16545), .ZN(
        U373) );
  INV_X1 U19745 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18833) );
  INV_X1 U19746 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19885) );
  AOI22_X1 U19747 ( .A1(n16544), .A2(n18833), .B1(n19885), .B2(n16545), .ZN(
        U374) );
  INV_X1 U19748 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18831) );
  INV_X1 U19749 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19884) );
  AOI22_X1 U19750 ( .A1(n16544), .A2(n18831), .B1(n19884), .B2(n16545), .ZN(
        U375) );
  INV_X1 U19751 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18810) );
  INV_X1 U19752 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19873) );
  AOI22_X1 U19753 ( .A1(n16544), .A2(n18810), .B1(n19873), .B2(n16545), .ZN(
        U376) );
  INV_X1 U19754 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16546) );
  NOR2_X1 U19755 ( .A1(n18799), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18798) );
  OAI22_X1 U19756 ( .A1(n18807), .A2(n18798), .B1(n18799), .B2(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18792) );
  OAI21_X1 U19757 ( .B1(n18807), .B2(n16546), .A(n18879), .ZN(P3_U2633) );
  NAND2_X1 U19758 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18905), .ZN(n16548) );
  OAI21_X1 U19759 ( .B1(n16555), .B2(n17483), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16547) );
  OAI21_X1 U19760 ( .B1(n16549), .B2(n16548), .A(n16547), .ZN(P3_U2634) );
  INV_X1 U19761 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18809) );
  AOI21_X1 U19762 ( .B1(n18807), .B2(n18809), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16550) );
  AOI22_X1 U19763 ( .A1(n18870), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16550), 
        .B2(n18941), .ZN(P3_U2635) );
  INV_X1 U19764 ( .A(BS16), .ZN(n21029) );
  AOI21_X1 U19765 ( .B1(n16551), .B2(n21029), .A(n18879), .ZN(n18878) );
  AOI21_X1 U19766 ( .B1(n18879), .B2(P3_STATEBS16_REG_SCAN_IN), .A(n18878), 
        .ZN(n16552) );
  INV_X1 U19767 ( .A(n16552), .ZN(P3_U2636) );
  NOR3_X1 U19768 ( .A1(n16555), .A2(n16554), .A3(n16553), .ZN(n18767) );
  NOR2_X1 U19769 ( .A1(n18767), .A2(n18781), .ZN(n18924) );
  OAI21_X1 U19770 ( .B1(n18924), .B2(n18255), .A(n16556), .ZN(P3_U2637) );
  NOR4_X1 U19771 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16560) );
  NOR4_X1 U19772 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16559) );
  NOR4_X1 U19773 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16558) );
  NOR4_X1 U19774 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16557) );
  NAND4_X1 U19775 ( .A1(n16560), .A2(n16559), .A3(n16558), .A4(n16557), .ZN(
        n16566) );
  NOR4_X1 U19776 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16564) );
  AOI211_X1 U19777 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16563) );
  NOR4_X1 U19778 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16562) );
  NOR4_X1 U19779 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16561) );
  NAND4_X1 U19780 ( .A1(n16564), .A2(n16563), .A3(n16562), .A4(n16561), .ZN(
        n16565) );
  NOR2_X1 U19781 ( .A1(n16566), .A2(n16565), .ZN(n18922) );
  INV_X1 U19782 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16568) );
  NOR3_X1 U19783 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16569) );
  OAI21_X1 U19784 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16569), .A(n18922), .ZN(
        n16567) );
  OAI21_X1 U19785 ( .B1(n18922), .B2(n16568), .A(n16567), .ZN(P3_U2638) );
  INV_X1 U19786 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16571) );
  NOR2_X1 U19787 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18916) );
  OAI21_X1 U19788 ( .B1(n16569), .B2(n18916), .A(n18922), .ZN(n16570) );
  OAI21_X1 U19789 ( .B1(n18922), .B2(n16571), .A(n16570), .ZN(P3_U2639) );
  NAND2_X1 U19790 ( .A1(n16901), .A2(n16572), .ZN(n16583) );
  XOR2_X1 U19791 ( .A(n16574), .B(n16573), .Z(n16578) );
  INV_X1 U19792 ( .A(n16913), .ZN(n18784) );
  OAI22_X1 U19793 ( .A1(n9893), .A2(n16885), .B1(n18872), .B2(n16575), .ZN(
        n16576) );
  OAI21_X1 U19794 ( .B1(n16891), .B2(n16579), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16580) );
  OAI211_X1 U19795 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16583), .A(n16581), .B(
        n16580), .ZN(P3_U2641) );
  INV_X1 U19796 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18867) );
  AOI22_X1 U19797 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16891), .B1(n16582), 
        .B2(n18867), .ZN(n16592) );
  INV_X1 U19798 ( .A(n16595), .ZN(n16584) );
  AOI21_X1 U19799 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16584), .A(n16583), .ZN(
        n16589) );
  AOI211_X1 U19800 ( .C1(n16587), .C2(n16586), .A(n16585), .B(n16913), .ZN(
        n16588) );
  AOI211_X1 U19801 ( .C1(n16590), .C2(P3_REIP_REG_29__SCAN_IN), .A(n16589), 
        .B(n16588), .ZN(n16591) );
  OAI211_X1 U19802 ( .C1(n16593), .C2(n16885), .A(n16592), .B(n16591), .ZN(
        P3_U2642) );
  AOI221_X1 U19803 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(P3_REIP_REG_27__SCAN_IN), .C1(n18866), .C2(n18863), .A(n16608), .ZN(n16594) );
  AOI21_X1 U19804 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n16891), .A(n16594), .ZN(
        n16603) );
  OAI21_X1 U19805 ( .B1(n16615), .B2(n16924), .A(n16937), .ZN(n16622) );
  AOI211_X1 U19806 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16611), .A(n16595), .B(
        n16933), .ZN(n16601) );
  INV_X1 U19807 ( .A(n16596), .ZN(n16599) );
  INV_X1 U19808 ( .A(n16597), .ZN(n16598) );
  AOI211_X1 U19809 ( .C1(n17554), .C2(n16599), .A(n16598), .B(n16913), .ZN(
        n16600) );
  AOI211_X1 U19810 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16622), .A(n16601), 
        .B(n16600), .ZN(n16602) );
  OAI211_X1 U19811 ( .C1(n17565), .C2(n16885), .A(n16603), .B(n16602), .ZN(
        P3_U2643) );
  INV_X1 U19812 ( .A(n16622), .ZN(n16614) );
  AOI211_X1 U19813 ( .C1(n16606), .C2(n16605), .A(n16604), .B(n16913), .ZN(
        n16610) );
  OAI22_X1 U19814 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16608), .B1(n16607), 
        .B2(n16885), .ZN(n16609) );
  AOI211_X1 U19815 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16891), .A(n16610), .B(
        n16609), .ZN(n16613) );
  OAI211_X1 U19816 ( .C1(n16616), .C2(n16982), .A(n16901), .B(n16611), .ZN(
        n16612) );
  OAI211_X1 U19817 ( .C1(n16614), .C2(n18863), .A(n16613), .B(n16612), .ZN(
        P3_U2644) );
  OR2_X1 U19818 ( .A1(n16615), .A2(n16924), .ZN(n16625) );
  AOI22_X1 U19819 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16922), .B1(
        n16891), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16624) );
  AOI211_X1 U19820 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16617), .A(n16616), .B(
        n16933), .ZN(n16621) );
  AOI211_X1 U19821 ( .C1(n17584), .C2(n16619), .A(n16618), .B(n16913), .ZN(
        n16620) );
  AOI211_X1 U19822 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16622), .A(n16621), 
        .B(n16620), .ZN(n16623) );
  OAI211_X1 U19823 ( .C1(n16626), .C2(n16625), .A(n16624), .B(n16623), .ZN(
        P3_U2645) );
  OR2_X1 U19824 ( .A1(n16933), .A2(n16627), .ZN(n16639) );
  AOI21_X1 U19825 ( .B1(n16901), .B2(n16627), .A(n16891), .ZN(n16638) );
  AOI21_X1 U19826 ( .B1(n16884), .B2(n16648), .A(n16929), .ZN(n16660) );
  OAI21_X1 U19827 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n16924), .A(n16660), 
        .ZN(n16636) );
  INV_X1 U19828 ( .A(n16628), .ZN(n16629) );
  AOI211_X1 U19829 ( .C1(n17597), .C2(n16630), .A(n16629), .B(n16913), .ZN(
        n16635) );
  NAND2_X1 U19830 ( .A1(n16884), .A2(n16631), .ZN(n16633) );
  OAI22_X1 U19831 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16633), .B1(n16632), 
        .B2(n16885), .ZN(n16634) );
  AOI211_X1 U19832 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16636), .A(n16635), 
        .B(n16634), .ZN(n16637) );
  OAI221_X1 U19833 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n16639), .C1(n16984), 
        .C2(n16638), .A(n16637), .ZN(P3_U2646) );
  NAND2_X1 U19834 ( .A1(n16884), .A2(n18856), .ZN(n16647) );
  AOI22_X1 U19835 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16922), .B1(
        n16891), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n16646) );
  INV_X1 U19836 ( .A(n16660), .ZN(n16644) );
  AOI21_X1 U19837 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16656), .A(n16639), .ZN(
        n16643) );
  AOI211_X1 U19838 ( .C1(n17612), .C2(n16641), .A(n16640), .B(n16913), .ZN(
        n16642) );
  AOI211_X1 U19839 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16644), .A(n16643), 
        .B(n16642), .ZN(n16645) );
  OAI211_X1 U19840 ( .C1(n16648), .C2(n16647), .A(n16646), .B(n16645), .ZN(
        P3_U2647) );
  INV_X1 U19841 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18854) );
  INV_X1 U19842 ( .A(n16649), .ZN(n16650) );
  AOI211_X1 U19843 ( .C1(n17625), .C2(n16651), .A(n16650), .B(n16913), .ZN(
        n16655) );
  NAND2_X1 U19844 ( .A1(n16884), .A2(n16652), .ZN(n16665) );
  NAND3_X1 U19845 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .A3(n16661), .ZN(n16653) );
  OAI22_X1 U19846 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16653), .B1(n17622), 
        .B2(n16885), .ZN(n16654) );
  AOI211_X1 U19847 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n16891), .A(n16655), .B(
        n16654), .ZN(n16659) );
  OAI211_X1 U19848 ( .C1(n16664), .C2(n16657), .A(n16901), .B(n16656), .ZN(
        n16658) );
  OAI211_X1 U19849 ( .C1(n16660), .C2(n18854), .A(n16659), .B(n16658), .ZN(
        P3_U2648) );
  INV_X1 U19850 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18852) );
  NOR2_X1 U19851 ( .A1(n16692), .A2(n16661), .ZN(n16677) );
  INV_X1 U19852 ( .A(n16677), .ZN(n16691) );
  INV_X1 U19853 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18850) );
  NAND2_X1 U19854 ( .A1(n16661), .A2(n18850), .ZN(n16674) );
  AOI211_X1 U19855 ( .C1(n17642), .C2(n16663), .A(n16662), .B(n16913), .ZN(
        n16669) );
  AOI211_X1 U19856 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16678), .A(n16664), .B(
        n16933), .ZN(n16668) );
  NOR3_X1 U19857 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n18850), .A3(n16665), 
        .ZN(n16667) );
  INV_X1 U19858 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16998) );
  OAI22_X1 U19859 ( .A1(n17639), .A2(n16885), .B1(n16934), .B2(n16998), .ZN(
        n16666) );
  NOR4_X1 U19860 ( .A1(n16669), .A2(n16668), .A3(n16667), .A4(n16666), .ZN(
        n16670) );
  OAI221_X1 U19861 ( .B1(n18852), .B2(n16691), .C1(n18852), .C2(n16674), .A(
        n16670), .ZN(P3_U2649) );
  INV_X1 U19862 ( .A(n16671), .ZN(n16672) );
  AOI211_X1 U19863 ( .C1(n17654), .C2(n16673), .A(n16672), .B(n16913), .ZN(
        n16676) );
  OAI21_X1 U19864 ( .B1(n17038), .B2(n16934), .A(n16674), .ZN(n16675) );
  AOI211_X1 U19865 ( .C1(n16677), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16676), 
        .B(n16675), .ZN(n16680) );
  OAI211_X1 U19866 ( .C1(n16686), .C2(n17038), .A(n16901), .B(n16678), .ZN(
        n16679) );
  OAI211_X1 U19867 ( .C1(n16885), .C2(n17651), .A(n16680), .B(n16679), .ZN(
        P3_U2650) );
  NOR2_X1 U19868 ( .A1(n16924), .A2(n16681), .ZN(n16709) );
  NOR2_X1 U19869 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16703), .ZN(n16682) );
  AOI22_X1 U19870 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16922), .B1(
        n16709), .B2(n16682), .ZN(n16690) );
  AOI211_X1 U19871 ( .C1(n16685), .C2(n16684), .A(n16683), .B(n16913), .ZN(
        n16688) );
  AOI211_X1 U19872 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16701), .A(n16686), .B(
        n16933), .ZN(n16687) );
  AOI211_X1 U19873 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16891), .A(n16688), .B(
        n16687), .ZN(n16689) );
  OAI211_X1 U19874 ( .C1(n18849), .C2(n16691), .A(n16690), .B(n16689), .ZN(
        P3_U2651) );
  NOR2_X1 U19875 ( .A1(n16692), .A2(n16709), .ZN(n16716) );
  INV_X1 U19876 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16698) );
  NAND2_X1 U19877 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17675), .ZN(
        n16711) );
  AOI21_X1 U19878 ( .B1(n16698), .B2(n16711), .A(n16693), .ZN(n16694) );
  INV_X1 U19879 ( .A(n16694), .ZN(n17676) );
  NAND2_X1 U19880 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16695), .ZN(
        n17752) );
  INV_X1 U19881 ( .A(n17752), .ZN(n16790) );
  NAND2_X1 U19882 ( .A1(n17749), .A2(n16790), .ZN(n16764) );
  NOR2_X1 U19883 ( .A1(n17740), .A2(n16764), .ZN(n17712) );
  NAND2_X1 U19884 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17712), .ZN(
        n16741) );
  OR2_X1 U19885 ( .A1(n16741), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16731) );
  OAI21_X1 U19886 ( .B1(n16711), .B2(n16731), .A(n12005), .ZN(n16697) );
  OAI21_X1 U19887 ( .B1(n17676), .B2(n16697), .A(n18784), .ZN(n16696) );
  AOI21_X1 U19888 ( .B1(n17676), .B2(n16697), .A(n16696), .ZN(n16700) );
  OAI22_X1 U19889 ( .A1(n16698), .A2(n16885), .B1(n16934), .B2(n16702), .ZN(
        n16699) );
  AOI211_X1 U19890 ( .C1(n16716), .C2(P3_REIP_REG_19__SCAN_IN), .A(n16700), 
        .B(n16699), .ZN(n16706) );
  OAI211_X1 U19891 ( .C1(n16707), .C2(n16702), .A(n16901), .B(n16701), .ZN(
        n16705) );
  OAI211_X1 U19892 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16709), .B(n16703), .ZN(n16704) );
  NAND4_X1 U19893 ( .A1(n16706), .A2(n18140), .A3(n16705), .A4(n16704), .ZN(
        P3_U2652) );
  AOI22_X1 U19894 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16922), .B1(
        n16891), .B2(P3_EBX_REG_18__SCAN_IN), .ZN(n16715) );
  INV_X1 U19895 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18844) );
  AOI211_X1 U19896 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16719), .A(n16707), .B(
        n16933), .ZN(n16708) );
  AOI211_X1 U19897 ( .C1(n16709), .C2(n18844), .A(n18071), .B(n16708), .ZN(
        n16714) );
  NAND2_X1 U19898 ( .A1(n16863), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16914) );
  INV_X1 U19899 ( .A(n16914), .ZN(n16877) );
  AOI21_X1 U19900 ( .B1(n16710), .B2(n16877), .A(n16862), .ZN(n16726) );
  OAI21_X1 U19901 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17675), .A(
        n16711), .ZN(n17685) );
  XNOR2_X1 U19902 ( .A(n16726), .B(n17685), .ZN(n16712) );
  AOI22_X1 U19903 ( .A1(n18784), .A2(n16712), .B1(P3_REIP_REG_18__SCAN_IN), 
        .B2(n16716), .ZN(n16713) );
  NAND3_X1 U19904 ( .A1(n16715), .A2(n16714), .A3(n16713), .ZN(P3_U2653) );
  INV_X1 U19905 ( .A(n16716), .ZN(n16729) );
  INV_X1 U19906 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18843) );
  NAND2_X1 U19907 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16718) );
  NOR2_X1 U19908 ( .A1(n16924), .A2(n16717), .ZN(n16757) );
  NAND2_X1 U19909 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16757), .ZN(n16742) );
  NOR3_X1 U19910 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16718), .A3(n16742), 
        .ZN(n16723) );
  OAI211_X1 U19911 ( .C1(n16733), .C2(n16721), .A(n16901), .B(n16719), .ZN(
        n16720) );
  OAI211_X1 U19912 ( .C1(n16934), .C2(n16721), .A(n18140), .B(n16720), .ZN(
        n16722) );
  AOI211_X1 U19913 ( .C1(n16922), .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16723), .B(n16722), .ZN(n16728) );
  NOR2_X1 U19914 ( .A1(n17908), .A2(n17698), .ZN(n16730) );
  INV_X1 U19915 ( .A(n16730), .ZN(n16724) );
  AOI21_X1 U19916 ( .B1(n17699), .B2(n16724), .A(n17675), .ZN(n17702) );
  NOR2_X1 U19917 ( .A1(n16913), .A2(n12005), .ZN(n16882) );
  AOI221_X1 U19918 ( .B1(n17698), .B2(n17702), .C1(n16914), .C2(n17702), .A(
        n16913), .ZN(n16725) );
  OAI22_X1 U19919 ( .A1(n17702), .A2(n16726), .B1(n16882), .B2(n16725), .ZN(
        n16727) );
  OAI211_X1 U19920 ( .C1(n16729), .C2(n18843), .A(n16728), .B(n16727), .ZN(
        P3_U2654) );
  INV_X1 U19921 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16735) );
  AOI21_X1 U19922 ( .B1(n16735), .B2(n16741), .A(n16730), .ZN(n17713) );
  NAND2_X1 U19923 ( .A1(n16768), .A2(n16731), .ZN(n16751) );
  OAI21_X1 U19924 ( .B1(n16753), .B2(n16924), .A(n16937), .ZN(n16759) );
  AOI21_X1 U19925 ( .B1(n12005), .B2(n16731), .A(n16913), .ZN(n16732) );
  AOI22_X1 U19926 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n16759), .B1(n17713), 
        .B2(n16732), .ZN(n16740) );
  INV_X1 U19927 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18840) );
  INV_X1 U19928 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18838) );
  AOI221_X1 U19929 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(P3_REIP_REG_15__SCAN_IN), .C1(n18840), .C2(n18838), .A(n16742), .ZN(n16738) );
  AOI211_X1 U19930 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16744), .A(n16733), .B(
        n16933), .ZN(n16737) );
  OAI22_X1 U19931 ( .A1(n16735), .A2(n16885), .B1(n16934), .B2(n16734), .ZN(
        n16736) );
  NOR4_X1 U19932 ( .A1(n18071), .A2(n16738), .A3(n16737), .A4(n16736), .ZN(
        n16739) );
  OAI211_X1 U19933 ( .C1(n17713), .C2(n16751), .A(n16740), .B(n16739), .ZN(
        P3_U2655) );
  OAI21_X1 U19934 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17712), .A(
        n16741), .ZN(n17723) );
  INV_X1 U19935 ( .A(n17723), .ZN(n16752) );
  NOR2_X1 U19936 ( .A1(n16862), .A2(n16863), .ZN(n16923) );
  NOR2_X1 U19937 ( .A1(n16923), .A2(n16913), .ZN(n16853) );
  OAI21_X1 U19938 ( .B1(n17712), .B2(n16862), .A(n16853), .ZN(n16750) );
  INV_X1 U19939 ( .A(n16759), .ZN(n16743) );
  AOI22_X1 U19940 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16743), .B1(n16742), 
        .B2(n18838), .ZN(n16748) );
  OAI211_X1 U19941 ( .C1(n16754), .C2(n16746), .A(n16901), .B(n16744), .ZN(
        n16745) );
  OAI211_X1 U19942 ( .C1(n16934), .C2(n16746), .A(n18140), .B(n16745), .ZN(
        n16747) );
  AOI211_X1 U19943 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16922), .A(
        n16748), .B(n16747), .ZN(n16749) );
  OAI221_X1 U19944 ( .B1(n16752), .B2(n16751), .C1(n17723), .C2(n16750), .A(
        n16749), .ZN(P3_U2656) );
  AOI22_X1 U19945 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16922), .B1(
        n16891), .B2(P3_EBX_REG_14__SCAN_IN), .ZN(n16763) );
  INV_X1 U19946 ( .A(n16753), .ZN(n16756) );
  AOI211_X1 U19947 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16769), .A(n16754), .B(
        n16933), .ZN(n16755) );
  AOI211_X1 U19948 ( .C1(n16757), .C2(n16756), .A(n18071), .B(n16755), .ZN(
        n16762) );
  AOI21_X1 U19949 ( .B1(n17740), .B2(n16764), .A(n17712), .ZN(n17742) );
  NAND3_X1 U19950 ( .A1(n17749), .A2(n16790), .A3(n16863), .ZN(n16767) );
  NAND2_X1 U19951 ( .A1(n12005), .A2(n16767), .ZN(n16758) );
  XNOR2_X1 U19952 ( .A(n17742), .B(n16758), .ZN(n16760) );
  AOI22_X1 U19953 ( .A1(n18784), .A2(n16760), .B1(P3_REIP_REG_14__SCAN_IN), 
        .B2(n16759), .ZN(n16761) );
  NAND3_X1 U19954 ( .A1(n16763), .A2(n16762), .A3(n16761), .ZN(P3_U2657) );
  NOR2_X1 U19955 ( .A1(n17766), .A2(n17752), .ZN(n16780) );
  OAI21_X1 U19956 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16780), .A(
        n16764), .ZN(n17753) );
  OAI21_X1 U19957 ( .B1(n16780), .B2(n16862), .A(n16853), .ZN(n16777) );
  AOI21_X1 U19958 ( .B1(n16884), .B2(n16783), .A(n16929), .ZN(n16793) );
  OAI21_X1 U19959 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n16924), .A(n16793), 
        .ZN(n16775) );
  INV_X1 U19960 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18834) );
  NAND3_X1 U19961 ( .A1(n16884), .A2(n16765), .A3(n18834), .ZN(n16766) );
  OAI211_X1 U19962 ( .C1(n17755), .C2(n16885), .A(n18140), .B(n16766), .ZN(
        n16774) );
  NAND3_X1 U19963 ( .A1(n16768), .A2(n17753), .A3(n16767), .ZN(n16771) );
  OAI211_X1 U19964 ( .C1(n16778), .C2(n16772), .A(n16901), .B(n16769), .ZN(
        n16770) );
  OAI211_X1 U19965 ( .C1(n16772), .C2(n16934), .A(n16771), .B(n16770), .ZN(
        n16773) );
  AOI211_X1 U19966 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16775), .A(n16774), 
        .B(n16773), .ZN(n16776) );
  OAI21_X1 U19967 ( .B1(n17753), .B2(n16777), .A(n16776), .ZN(P3_U2658) );
  AOI211_X1 U19968 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16796), .A(n16778), .B(
        n16933), .ZN(n16779) );
  AOI21_X1 U19969 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n16891), .A(n16779), .ZN(
        n16787) );
  AOI21_X1 U19970 ( .B1(n17766), .B2(n17752), .A(n16780), .ZN(n17769) );
  OAI21_X1 U19971 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17752), .A(
        n12005), .ZN(n16781) );
  XNOR2_X1 U19972 ( .A(n17769), .B(n16781), .ZN(n16785) );
  NAND2_X1 U19973 ( .A1(n16884), .A2(n18832), .ZN(n16782) );
  OAI22_X1 U19974 ( .A1(n17766), .A2(n16885), .B1(n16783), .B2(n16782), .ZN(
        n16784) );
  AOI211_X1 U19975 ( .C1(n18784), .C2(n16785), .A(n18071), .B(n16784), .ZN(
        n16786) );
  OAI211_X1 U19976 ( .C1(n18832), .C2(n16793), .A(n16787), .B(n16786), .ZN(
        P3_U2659) );
  AOI21_X1 U19977 ( .B1(n16884), .B2(n16788), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16794) );
  OR2_X1 U19978 ( .A1(n17908), .A2(n16789), .ZN(n16802) );
  AOI21_X1 U19979 ( .B1(n16800), .B2(n16802), .A(n16790), .ZN(n17781) );
  OAI21_X1 U19980 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16802), .A(
        n12005), .ZN(n16791) );
  XOR2_X1 U19981 ( .A(n17781), .B(n16791), .Z(n16792) );
  OAI22_X1 U19982 ( .A1(n16794), .A2(n16793), .B1(n16913), .B2(n16792), .ZN(
        n16795) );
  AOI211_X1 U19983 ( .C1(n16891), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18071), .B(
        n16795), .ZN(n16799) );
  OAI211_X1 U19984 ( .C1(n16807), .C2(n16797), .A(n16901), .B(n16796), .ZN(
        n16798) );
  OAI211_X1 U19985 ( .C1(n16885), .C2(n16800), .A(n16799), .B(n16798), .ZN(
        P3_U2660) );
  OR2_X1 U19986 ( .A1(n17819), .A2(n17834), .ZN(n17817) );
  NOR3_X1 U19987 ( .A1(n17821), .A2(n17817), .A3(n16914), .ZN(n16818) );
  AOI21_X1 U19988 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16818), .A(
        n16862), .ZN(n16817) );
  NAND2_X1 U19989 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17853), .ZN(
        n16864) );
  INV_X1 U19990 ( .A(n16864), .ZN(n16852) );
  NAND2_X1 U19991 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16852), .ZN(
        n16851) );
  NOR2_X1 U19992 ( .A1(n16801), .A2(n16851), .ZN(n16814) );
  OAI21_X1 U19993 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16814), .A(
        n16802), .ZN(n17790) );
  XOR2_X1 U19994 ( .A(n16817), .B(n17790), .Z(n16813) );
  NOR3_X1 U19995 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n16924), .A3(n16803), 
        .ZN(n16804) );
  AOI211_X1 U19996 ( .C1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n16922), .A(
        n18071), .B(n16804), .ZN(n16812) );
  OAI21_X1 U19997 ( .B1(n16924), .B2(n16806), .A(n16937), .ZN(n16805) );
  INV_X1 U19998 ( .A(n16805), .ZN(n16836) );
  INV_X1 U19999 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18826) );
  NAND3_X1 U20000 ( .A1(n16884), .A2(n16806), .A3(n18826), .ZN(n16823) );
  AOI21_X1 U20001 ( .B1(n16836), .B2(n16823), .A(n18828), .ZN(n16810) );
  AOI211_X1 U20002 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16808), .A(n16807), .B(
        n16933), .ZN(n16809) );
  AOI211_X1 U20003 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16891), .A(n16810), .B(
        n16809), .ZN(n16811) );
  OAI211_X1 U20004 ( .C1(n16913), .C2(n16813), .A(n16812), .B(n16811), .ZN(
        P3_U2661) );
  OR2_X1 U20005 ( .A1(n16933), .A2(n16816), .ZN(n16825) );
  INV_X1 U20006 ( .A(n16851), .ZN(n16838) );
  AND2_X1 U20007 ( .A1(n17816), .A2(n16838), .ZN(n16827) );
  INV_X1 U20008 ( .A(n16814), .ZN(n16815) );
  OAI21_X1 U20009 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16827), .A(
        n16815), .ZN(n17806) );
  INV_X1 U20010 ( .A(n16882), .ZN(n16921) );
  OAI21_X1 U20011 ( .B1(n17806), .B2(n16921), .A(n18140), .ZN(n16822) );
  OAI221_X1 U20012 ( .B1(n16891), .B2(n16901), .C1(n16891), .C2(n16816), .A(
        P3_EBX_REG_9__SCAN_IN), .ZN(n16820) );
  OAI211_X1 U20013 ( .C1(n16818), .C2(n17806), .A(n18784), .B(n16817), .ZN(
        n16819) );
  OAI211_X1 U20014 ( .C1(n16836), .C2(n18826), .A(n16820), .B(n16819), .ZN(
        n16821) );
  AOI211_X1 U20015 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n16922), .A(
        n16822), .B(n16821), .ZN(n16824) );
  OAI211_X1 U20016 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n16825), .A(n16824), .B(
        n16823), .ZN(P3_U2662) );
  AOI21_X1 U20017 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n16845), .A(n16825), .ZN(
        n16826) );
  AOI211_X1 U20018 ( .C1(n16891), .C2(P3_EBX_REG_8__SCAN_IN), .A(n18071), .B(
        n16826), .ZN(n16835) );
  NAND2_X1 U20019 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16838), .ZN(
        n16837) );
  AOI21_X1 U20020 ( .B1(n17821), .B2(n16837), .A(n16827), .ZN(n17824) );
  NOR2_X1 U20021 ( .A1(n17817), .A2(n16914), .ZN(n16828) );
  NOR2_X1 U20022 ( .A1(n16828), .A2(n16862), .ZN(n16830) );
  OAI21_X1 U20023 ( .B1(n17824), .B2(n16830), .A(n18784), .ZN(n16829) );
  AOI21_X1 U20024 ( .B1(n17824), .B2(n16830), .A(n16829), .ZN(n16833) );
  NOR3_X1 U20025 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16924), .A3(n16831), .ZN(
        n16832) );
  AOI211_X1 U20026 ( .C1(n16922), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16833), .B(n16832), .ZN(n16834) );
  OAI211_X1 U20027 ( .C1(n18824), .C2(n16836), .A(n16835), .B(n16834), .ZN(
        P3_U2663) );
  OAI21_X1 U20028 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16838), .A(
        n16837), .ZN(n17845) );
  AOI21_X1 U20029 ( .B1(n16838), .B2(n16863), .A(n16862), .ZN(n16857) );
  XNOR2_X1 U20030 ( .A(n17845), .B(n16857), .ZN(n16844) );
  NAND2_X1 U20031 ( .A1(n16884), .A2(n16840), .ZN(n16839) );
  NAND2_X1 U20032 ( .A1(n16935), .A2(n16839), .ZN(n16866) );
  INV_X1 U20033 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18820) );
  NAND3_X1 U20034 ( .A1(n16884), .A2(n16840), .A3(n18820), .ZN(n16859) );
  INV_X1 U20035 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18822) );
  AOI21_X1 U20036 ( .B1(n16866), .B2(n16859), .A(n18822), .ZN(n16843) );
  NAND4_X1 U20037 ( .A1(n16884), .A2(P3_REIP_REG_6__SCAN_IN), .A3(n16840), 
        .A4(n18822), .ZN(n16841) );
  OAI211_X1 U20038 ( .C1(n16934), .C2(n16846), .A(n18140), .B(n16841), .ZN(
        n16842) );
  AOI211_X1 U20039 ( .C1(n18784), .C2(n16844), .A(n16843), .B(n16842), .ZN(
        n16848) );
  OAI211_X1 U20040 ( .C1(n16849), .C2(n16846), .A(n16901), .B(n16845), .ZN(
        n16847) );
  OAI211_X1 U20041 ( .C1(n16885), .C2(n17834), .A(n16848), .B(n16847), .ZN(
        P3_U2664) );
  AOI211_X1 U20042 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16869), .A(n16849), .B(
        n16933), .ZN(n16850) );
  NOR2_X1 U20043 ( .A1(n18071), .A2(n16850), .ZN(n16861) );
  OAI21_X1 U20044 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16852), .A(
        n16851), .ZN(n17856) );
  INV_X1 U20045 ( .A(n16853), .ZN(n16932) );
  AOI211_X1 U20046 ( .C1(n12005), .C2(n16864), .A(n17856), .B(n16932), .ZN(
        n16856) );
  OAI22_X1 U20047 ( .A1(n16934), .A2(n16854), .B1(n18820), .B2(n16866), .ZN(
        n16855) );
  AOI211_X1 U20048 ( .C1(n16922), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16856), .B(n16855), .ZN(n16860) );
  NAND3_X1 U20049 ( .A1(n18784), .A2(n17856), .A3(n16857), .ZN(n16858) );
  NAND4_X1 U20050 ( .A1(n16861), .A2(n16860), .A3(n16859), .A4(n16858), .ZN(
        P3_U2665) );
  NOR2_X1 U20051 ( .A1(n16924), .A2(n16883), .ZN(n16887) );
  AOI21_X1 U20052 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n16887), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n16867) );
  NOR3_X1 U20053 ( .A1(n17908), .A2(n17873), .A3(n17880), .ZN(n16873) );
  AOI21_X1 U20054 ( .B1(n16873), .B2(n16863), .A(n16862), .ZN(n16875) );
  OAI21_X1 U20055 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16873), .A(
        n16864), .ZN(n17867) );
  XOR2_X1 U20056 ( .A(n16875), .B(n17867), .Z(n16865) );
  OAI22_X1 U20057 ( .A1(n16867), .A2(n16866), .B1(n16913), .B2(n16865), .ZN(
        n16868) );
  AOI211_X1 U20058 ( .C1(n16891), .C2(P3_EBX_REG_5__SCAN_IN), .A(n18071), .B(
        n16868), .ZN(n16872) );
  OAI211_X1 U20059 ( .C1(n16878), .C2(n16870), .A(n16901), .B(n16869), .ZN(
        n16871) );
  OAI211_X1 U20060 ( .C1(n16885), .C2(n17862), .A(n16872), .B(n16871), .ZN(
        P3_U2666) );
  NOR2_X1 U20061 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17873), .ZN(
        n16876) );
  OR2_X1 U20062 ( .A1(n17908), .A2(n17873), .ZN(n16895) );
  AOI21_X1 U20063 ( .B1(n17880), .B2(n16895), .A(n16873), .ZN(n17877) );
  INV_X1 U20064 ( .A(n17877), .ZN(n16874) );
  AOI22_X1 U20065 ( .A1(n16877), .A2(n16876), .B1(n16875), .B2(n16874), .ZN(
        n16890) );
  AOI211_X1 U20066 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16900), .A(n16878), .B(
        n16933), .ZN(n16881) );
  NOR2_X1 U20067 ( .A1(n18267), .A2(n18946), .ZN(n16893) );
  OAI221_X1 U20068 ( .B1(n18948), .B2(n17208), .C1(n18948), .C2(n16879), .A(
        n18140), .ZN(n16880) );
  AOI211_X1 U20069 ( .C1(n16882), .C2(n17877), .A(n16881), .B(n16880), .ZN(
        n16889) );
  NAND2_X1 U20070 ( .A1(n16884), .A2(n16883), .ZN(n16892) );
  NAND2_X1 U20071 ( .A1(n16937), .A2(n16892), .ZN(n16898) );
  INV_X1 U20072 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n17262) );
  OAI22_X1 U20073 ( .A1(n17880), .A2(n16885), .B1(n16934), .B2(n17262), .ZN(
        n16886) );
  AOI221_X1 U20074 ( .B1(n16887), .B2(n18816), .C1(n16898), .C2(
        P3_REIP_REG_4__SCAN_IN), .A(n16886), .ZN(n16888) );
  OAI211_X1 U20075 ( .C1(n16890), .C2(n16913), .A(n16889), .B(n16888), .ZN(
        P3_U2667) );
  AOI22_X1 U20076 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n16922), .B1(
        n16891), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n16905) );
  INV_X1 U20077 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18811) );
  INV_X1 U20078 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18812) );
  NOR2_X1 U20079 ( .A1(n18811), .A2(n18812), .ZN(n16916) );
  INV_X1 U20080 ( .A(n16892), .ZN(n16894) );
  NAND2_X1 U20081 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18712), .ZN(
        n18716) );
  AOI21_X1 U20082 ( .B1(n12014), .B2(n18716), .A(n17230), .ZN(n18886) );
  AOI22_X1 U20083 ( .A1(n16916), .A2(n16894), .B1(n16893), .B2(n18886), .ZN(
        n16904) );
  INV_X1 U20084 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17900) );
  NOR2_X1 U20085 ( .A1(n17908), .A2(n17900), .ZN(n16906) );
  OAI21_X1 U20086 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n16906), .A(
        n16895), .ZN(n16896) );
  INV_X1 U20087 ( .A(n16896), .ZN(n17886) );
  INV_X1 U20088 ( .A(n16906), .ZN(n16897) );
  OAI21_X1 U20089 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16897), .A(
        n12005), .ZN(n16912) );
  XNOR2_X1 U20090 ( .A(n17886), .B(n16912), .ZN(n16899) );
  AOI22_X1 U20091 ( .A1(n18784), .A2(n16899), .B1(P3_REIP_REG_3__SCAN_IN), 
        .B2(n16898), .ZN(n16903) );
  OAI211_X1 U20092 ( .C1(n16907), .C2(n17267), .A(n16901), .B(n16900), .ZN(
        n16902) );
  NAND4_X1 U20093 ( .A1(n16905), .A2(n16904), .A3(n16903), .A4(n16902), .ZN(
        P3_U2668) );
  AOI21_X1 U20094 ( .B1(n17908), .B2(n17900), .A(n16906), .ZN(n16915) );
  INV_X1 U20095 ( .A(n16915), .ZN(n17896) );
  NAND2_X1 U20096 ( .A1(n17284), .A2(n17278), .ZN(n16908) );
  AOI211_X1 U20097 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16908), .A(n16907), .B(
        n16933), .ZN(n16911) );
  NAND2_X1 U20098 ( .A1(n18728), .A2(n18897), .ZN(n18718) );
  INV_X1 U20099 ( .A(n18718), .ZN(n18722) );
  AOI21_X1 U20100 ( .B1(n18712), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n18722), .ZN(n18895) );
  INV_X1 U20101 ( .A(n18895), .ZN(n18736) );
  OAI22_X1 U20102 ( .A1(n16934), .A2(n16909), .B1(n18736), .B2(n18948), .ZN(
        n16910) );
  AOI211_X1 U20103 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(n16929), .A(n16911), .B(
        n16910), .ZN(n16920) );
  AOI211_X1 U20104 ( .C1(n16915), .C2(n16914), .A(n16913), .B(n16912), .ZN(
        n16918) );
  AOI211_X1 U20105 ( .C1(n18811), .C2(n18812), .A(n16916), .B(n16924), .ZN(
        n16917) );
  AOI211_X1 U20106 ( .C1(n16922), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n16918), .B(n16917), .ZN(n16919) );
  OAI211_X1 U20107 ( .C1(n17896), .C2(n16921), .A(n16920), .B(n16919), .ZN(
        P3_U2669) );
  AOI21_X1 U20108 ( .B1(n16923), .B2(n18784), .A(n16922), .ZN(n16931) );
  OAI22_X1 U20109 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16924), .B1(n16934), 
        .B2(n17278), .ZN(n16928) );
  OAI21_X1 U20110 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n16925), .ZN(n17280) );
  NAND2_X1 U20111 ( .A1(n18728), .A2(n16926), .ZN(n18898) );
  OAI22_X1 U20112 ( .A1(n16933), .A2(n17280), .B1(n18898), .B2(n18948), .ZN(
        n16927) );
  AOI211_X1 U20113 ( .C1(n16929), .C2(P3_REIP_REG_1__SCAN_IN), .A(n16928), .B(
        n16927), .ZN(n16930) );
  OAI221_X1 U20114 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16932), .C1(
        n17908), .C2(n16931), .A(n16930), .ZN(P3_U2670) );
  NAND2_X1 U20115 ( .A1(n16934), .A2(n16933), .ZN(n16936) );
  AOI22_X1 U20116 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n16936), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n16935), .ZN(n16939) );
  NAND3_X1 U20117 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18892), .A3(
        n16937), .ZN(n16938) );
  OAI211_X1 U20118 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18948), .A(
        n16939), .B(n16938), .ZN(P3_U2671) );
  INV_X1 U20119 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17019) );
  NAND3_X1 U20120 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_24__SCAN_IN), .ZN(n16941) );
  NOR3_X1 U20121 ( .A1(n16942), .A2(n16941), .A3(n16940), .ZN(n16978) );
  INV_X1 U20122 ( .A(n16978), .ZN(n16943) );
  NOR4_X1 U20123 ( .A1(n16944), .A2(n17019), .A3(n17065), .A4(n16943), .ZN(
        n16972) );
  NAND2_X1 U20124 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16972), .ZN(n16971) );
  INV_X1 U20125 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n16946) );
  INV_X1 U20126 ( .A(n16971), .ZN(n16945) );
  OAI33_X1 U20127 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n16971), .A3(n18294), 
        .B1(n16946), .B2(n17282), .B3(n16945), .ZN(P3_U2672) );
  AOI22_X1 U20128 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16957) );
  AOI22_X1 U20129 ( .A1(n17202), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16948) );
  AOI22_X1 U20130 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16947) );
  OAI211_X1 U20131 ( .C1(n17167), .C2(n16949), .A(n16948), .B(n16947), .ZN(
        n16955) );
  AOI22_X1 U20132 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16953) );
  AOI22_X1 U20133 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16952) );
  AOI22_X1 U20134 ( .A1(n17204), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16951) );
  NAND2_X1 U20135 ( .A1(n17209), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n16950) );
  NAND4_X1 U20136 ( .A1(n16953), .A2(n16952), .A3(n16951), .A4(n16950), .ZN(
        n16954) );
  AOI211_X1 U20137 ( .C1(n12616), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n16955), .B(n16954), .ZN(n16956) );
  OAI211_X1 U20138 ( .C1(n17163), .C2(n16958), .A(n16957), .B(n16956), .ZN(
        n16975) );
  NAND2_X1 U20139 ( .A1(n16976), .A2(n16975), .ZN(n16974) );
  AOI22_X1 U20140 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12616), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16968) );
  AOI22_X1 U20141 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16960) );
  AOI22_X1 U20142 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16959) );
  OAI211_X1 U20143 ( .C1(n17235), .C2(n17115), .A(n16960), .B(n16959), .ZN(
        n16966) );
  AOI22_X1 U20144 ( .A1(n17202), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16964) );
  AOI22_X1 U20145 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16963) );
  AOI22_X1 U20146 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17161), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16962) );
  NAND2_X1 U20147 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n16961) );
  NAND4_X1 U20148 ( .A1(n16964), .A2(n16963), .A3(n16962), .A4(n16961), .ZN(
        n16965) );
  AOI211_X1 U20149 ( .C1(n9630), .C2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n16966), .B(n16965), .ZN(n16967) );
  OAI211_X1 U20150 ( .C1(n17227), .C2(n16969), .A(n16968), .B(n16967), .ZN(
        n16970) );
  XOR2_X1 U20151 ( .A(n16974), .B(n16970), .Z(n17299) );
  OAI211_X1 U20152 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16972), .A(n16971), .B(
        n17274), .ZN(n16973) );
  OAI21_X1 U20153 ( .B1(n17299), .B2(n17274), .A(n16973), .ZN(P3_U2673) );
  OAI21_X1 U20154 ( .B1(n16976), .B2(n16975), .A(n16974), .ZN(n17303) );
  NOR2_X1 U20155 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17004), .ZN(n16977) );
  AOI22_X1 U20156 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16979), .B1(n16978), 
        .B2(n16977), .ZN(n16980) );
  OAI21_X1 U20157 ( .B1(n17303), .B2(n17274), .A(n16980), .ZN(P3_U2674) );
  OAI211_X1 U20158 ( .C1(n17312), .C2(n17311), .A(n17282), .B(n17310), .ZN(
        n16981) );
  OAI221_X1 U20159 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n16985), .C1(n16982), 
        .C2(n16987), .A(n16981), .ZN(P3_U2676) );
  INV_X1 U20160 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16988) );
  AOI21_X1 U20161 ( .B1(n16983), .B2(n16990), .A(n17312), .ZN(n17317) );
  NAND2_X1 U20162 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17003), .ZN(n16989) );
  NOR2_X1 U20163 ( .A1(n16984), .A2(n16989), .ZN(n16994) );
  AOI22_X1 U20164 ( .A1(n17282), .A2(n17317), .B1(n16994), .B2(n16985), .ZN(
        n16986) );
  OAI21_X1 U20165 ( .B1(n16988), .B2(n16987), .A(n16986), .ZN(P3_U2677) );
  INV_X1 U20166 ( .A(n16989), .ZN(n16997) );
  AOI21_X1 U20167 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17274), .A(n16997), .ZN(
        n16993) );
  OAI21_X1 U20168 ( .B1(n16992), .B2(n16991), .A(n16990), .ZN(n17326) );
  OAI22_X1 U20169 ( .A1(n16994), .A2(n16993), .B1(n17274), .B2(n17326), .ZN(
        P3_U2678) );
  AOI21_X1 U20170 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17274), .A(n17003), .ZN(
        n16996) );
  XNOR2_X1 U20171 ( .A(n16995), .B(n16999), .ZN(n17331) );
  OAI22_X1 U20172 ( .A1(n16997), .A2(n16996), .B1(n17274), .B2(n17331), .ZN(
        P3_U2679) );
  NOR3_X1 U20173 ( .A1(n16998), .A2(n17038), .A3(n17004), .ZN(n17018) );
  AOI21_X1 U20174 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17274), .A(n17018), .ZN(
        n17002) );
  OAI21_X1 U20175 ( .B1(n17001), .B2(n17000), .A(n16999), .ZN(n17336) );
  OAI22_X1 U20176 ( .A1(n17003), .A2(n17002), .B1(n17274), .B2(n17336), .ZN(
        P3_U2680) );
  INV_X1 U20177 ( .A(n17004), .ZN(n17036) );
  AOI22_X1 U20178 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17274), .B1(
        P3_EBX_REG_21__SCAN_IN), .B2(n17036), .ZN(n17017) );
  INV_X1 U20179 ( .A(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17006) );
  AOI22_X1 U20180 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17005) );
  OAI21_X1 U20181 ( .B1(n12100), .B2(n17006), .A(n17005), .ZN(n17016) );
  AOI22_X1 U20182 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17014) );
  OAI22_X1 U20183 ( .A1(n17163), .A2(n17007), .B1(n17167), .B2(n17131), .ZN(
        n17012) );
  AOI22_X1 U20184 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17010) );
  AOI22_X1 U20185 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17009) );
  AOI22_X1 U20186 ( .A1(n12616), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17209), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17008) );
  NAND3_X1 U20187 ( .A1(n17010), .A2(n17009), .A3(n17008), .ZN(n17011) );
  AOI211_X1 U20188 ( .C1(n17230), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n17012), .B(n17011), .ZN(n17013) );
  OAI211_X1 U20189 ( .C1(n17227), .C2(n17256), .A(n17014), .B(n17013), .ZN(
        n17015) );
  AOI211_X1 U20190 ( .C1(n17231), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n17016), .B(n17015), .ZN(n17339) );
  OAI22_X1 U20191 ( .A1(n17018), .A2(n17017), .B1(n17339), .B2(n17274), .ZN(
        P3_U2681) );
  OAI21_X1 U20192 ( .B1(n17019), .B2(n17065), .A(n17274), .ZN(n17052) );
  AOI22_X1 U20193 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U20194 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17021) );
  OAI21_X1 U20195 ( .B1(n9699), .B2(n17022), .A(n17021), .ZN(n17031) );
  AOI22_X1 U20196 ( .A1(n9631), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9633), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20197 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17024) );
  AOI22_X1 U20198 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17101), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17023) );
  OAI211_X1 U20199 ( .C1(n17235), .C2(n17025), .A(n17024), .B(n17023), .ZN(
        n17026) );
  AOI21_X1 U20200 ( .B1(n9630), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n17026), .ZN(n17027) );
  OAI211_X1 U20201 ( .C1(n17205), .C2(n17029), .A(n17028), .B(n17027), .ZN(
        n17030) );
  AOI211_X1 U20202 ( .C1(n17230), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n17031), .B(n17030), .ZN(n17032) );
  OAI211_X1 U20203 ( .C1(n17035), .C2(n17034), .A(n17033), .B(n17032), .ZN(
        n17344) );
  AOI22_X1 U20204 ( .A1(n17282), .A2(n17344), .B1(n17036), .B2(n17038), .ZN(
        n17037) );
  OAI21_X1 U20205 ( .B1(n17038), .B2(n17052), .A(n17037), .ZN(P3_U2682) );
  AOI22_X1 U20206 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17039) );
  OAI21_X1 U20207 ( .B1(n12562), .B2(n17040), .A(n17039), .ZN(n17050) );
  AOI22_X1 U20208 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17225), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17048) );
  OAI22_X1 U20209 ( .A1(n17163), .A2(n17041), .B1(n17099), .B2(n18525), .ZN(
        n17046) );
  AOI22_X1 U20210 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U20211 ( .A1(n17202), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U20212 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17209), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17042) );
  NAND3_X1 U20213 ( .A1(n17044), .A2(n17043), .A3(n17042), .ZN(n17045) );
  AOI211_X1 U20214 ( .C1(n12616), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n17046), .B(n17045), .ZN(n17047) );
  OAI211_X1 U20215 ( .C1(n17227), .C2(n17266), .A(n17048), .B(n17047), .ZN(
        n17049) );
  AOI211_X1 U20216 ( .C1(n17230), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n17050), .B(n17049), .ZN(n17352) );
  NOR2_X1 U20217 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17051), .ZN(n17053) );
  OAI22_X1 U20218 ( .A1(n17352), .A2(n17274), .B1(n17053), .B2(n17052), .ZN(
        P3_U2683) );
  AOI22_X1 U20219 ( .A1(n17204), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9630), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17064) );
  AOI22_X1 U20220 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17055) );
  AOI22_X1 U20221 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17161), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17054) );
  OAI211_X1 U20222 ( .C1(n17235), .C2(n17056), .A(n17055), .B(n17054), .ZN(
        n17062) );
  AOI22_X1 U20223 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17060) );
  AOI22_X1 U20224 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17059) );
  AOI22_X1 U20225 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17058) );
  NAND2_X1 U20226 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n17057) );
  NAND4_X1 U20227 ( .A1(n17060), .A2(n17059), .A3(n17058), .A4(n17057), .ZN(
        n17061) );
  AOI211_X1 U20228 ( .C1(n12616), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n17062), .B(n17061), .ZN(n17063) );
  OAI211_X1 U20229 ( .C1(n17217), .C2(n17171), .A(n17064), .B(n17063), .ZN(
        n17353) );
  INV_X1 U20230 ( .A(n17353), .ZN(n17067) );
  OAI21_X1 U20231 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17082), .A(n17065), .ZN(
        n17066) );
  AOI22_X1 U20232 ( .A1(n17282), .A2(n17067), .B1(n17066), .B2(n17274), .ZN(
        P3_U2684) );
  OAI21_X1 U20233 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17068), .A(n17274), .ZN(
        n17081) );
  AOI22_X1 U20234 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17079) );
  AOI22_X1 U20235 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17070) );
  AOI22_X1 U20236 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17069) );
  OAI211_X1 U20237 ( .C1(n17235), .C2(n17071), .A(n17070), .B(n17069), .ZN(
        n17077) );
  AOI22_X1 U20238 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17075) );
  AOI22_X1 U20239 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17074) );
  AOI22_X1 U20240 ( .A1(n17228), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17073) );
  NAND2_X1 U20241 ( .A1(n12616), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n17072) );
  NAND4_X1 U20242 ( .A1(n17075), .A2(n17074), .A3(n17073), .A4(n17072), .ZN(
        n17076) );
  AOI211_X1 U20243 ( .C1(n9630), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n17077), .B(n17076), .ZN(n17078) );
  OAI211_X1 U20244 ( .C1(n17227), .C2(n17276), .A(n17079), .B(n17078), .ZN(
        n17358) );
  INV_X1 U20245 ( .A(n17358), .ZN(n17080) );
  OAI22_X1 U20246 ( .A1(n17082), .A2(n17081), .B1(n17080), .B2(n17274), .ZN(
        P3_U2685) );
  AOI22_X1 U20247 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17101), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17092) );
  AOI22_X1 U20248 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17161), .ZN(n17084) );
  AOI22_X1 U20249 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17229), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17083) );
  OAI211_X1 U20250 ( .C1(n17207), .C2(n17235), .A(n17084), .B(n17083), .ZN(
        n17090) );
  AOI22_X1 U20251 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17088) );
  AOI22_X1 U20252 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17185), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17223), .ZN(n17087) );
  AOI22_X1 U20253 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12616), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17086) );
  NAND2_X1 U20254 ( .A1(n17204), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n17085) );
  NAND4_X1 U20255 ( .A1(n17088), .A2(n17087), .A3(n17086), .A4(n17085), .ZN(
        n17089) );
  AOI211_X1 U20256 ( .C1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .C2(n9630), .A(
        n17090), .B(n17089), .ZN(n17091) );
  OAI211_X1 U20257 ( .C1(n17093), .C2(n12608), .A(n17092), .B(n17091), .ZN(
        n17364) );
  INV_X1 U20258 ( .A(n17364), .ZN(n17097) );
  OAI21_X1 U20259 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17095), .A(n17094), .ZN(
        n17096) );
  AOI22_X1 U20260 ( .A1(n17282), .A2(n17097), .B1(n17096), .B2(n17274), .ZN(
        P3_U2686) );
  NAND4_X1 U20261 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(P3_EBX_REG_13__SCAN_IN), .A4(n17160), .ZN(n17128) );
  AOI22_X1 U20262 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17098) );
  OAI21_X1 U20263 ( .B1(n17099), .B2(n18513), .A(n17098), .ZN(n17110) );
  AOI22_X1 U20264 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17108) );
  AOI22_X1 U20265 ( .A1(n17204), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17209), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17100) );
  INV_X1 U20266 ( .A(n17100), .ZN(n17106) );
  AOI22_X1 U20267 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17104) );
  AOI22_X1 U20268 ( .A1(n17202), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17103) );
  AOI22_X1 U20269 ( .A1(n12616), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9630), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17102) );
  NAND3_X1 U20270 ( .A1(n17104), .A2(n17103), .A3(n17102), .ZN(n17105) );
  AOI211_X1 U20271 ( .C1(n17230), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n17106), .B(n17105), .ZN(n17107) );
  OAI211_X1 U20272 ( .C1(n17217), .C2(n17240), .A(n17108), .B(n17107), .ZN(
        n17109) );
  AOI211_X1 U20273 ( .C1(n17161), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n17110), .B(n17109), .ZN(n17375) );
  NAND3_X1 U20274 ( .A1(n17128), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n17274), 
        .ZN(n17111) );
  OAI221_X1 U20275 ( .B1(n17128), .B2(P3_EBX_REG_16__SCAN_IN), .C1(n17274), 
        .C2(n17375), .A(n17111), .ZN(P3_U2687) );
  AOI22_X1 U20276 ( .A1(n17202), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17112) );
  OAI21_X1 U20277 ( .B1(n17114), .B2(n17113), .A(n17112), .ZN(n17126) );
  INV_X1 U20278 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17124) );
  AOI22_X1 U20279 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17123) );
  OAI22_X1 U20280 ( .A1(n17205), .A2(n17116), .B1(n12562), .B2(n17115), .ZN(
        n17121) );
  AOI22_X1 U20281 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17231), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17119) );
  AOI22_X1 U20282 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17118) );
  AOI22_X1 U20283 ( .A1(n9630), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17209), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17117) );
  NAND3_X1 U20284 ( .A1(n17119), .A2(n17118), .A3(n17117), .ZN(n17120) );
  AOI211_X1 U20285 ( .C1(n17204), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n17121), .B(n17120), .ZN(n17122) );
  OAI211_X1 U20286 ( .C1(n17241), .C2(n17124), .A(n17123), .B(n17122), .ZN(
        n17125) );
  AOI211_X1 U20287 ( .C1(n17225), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n17126), .B(n17125), .ZN(n17379) );
  INV_X1 U20288 ( .A(n17127), .ZN(n17144) );
  OAI211_X1 U20289 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n17144), .A(n17128), .B(
        n17274), .ZN(n17129) );
  OAI21_X1 U20290 ( .B1(n17379), .B2(n17274), .A(n17129), .ZN(P3_U2688) );
  AOI22_X1 U20291 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17274), .B1(
        P3_EBX_REG_13__SCAN_IN), .B2(n17160), .ZN(n17143) );
  AOI22_X1 U20292 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17225), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17130) );
  OAI21_X1 U20293 ( .B1(n17184), .B2(n17131), .A(n17130), .ZN(n17141) );
  INV_X1 U20294 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17139) );
  AOI22_X1 U20295 ( .A1(n9631), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17138) );
  AOI22_X1 U20296 ( .A1(n12616), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17132) );
  OAI21_X1 U20297 ( .B1(n12100), .B2(n18532), .A(n17132), .ZN(n17136) );
  AOI22_X1 U20298 ( .A1(n17202), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17134) );
  AOI22_X1 U20299 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17133) );
  OAI211_X1 U20300 ( .C1(n17235), .C2(n17256), .A(n17134), .B(n17133), .ZN(
        n17135) );
  AOI211_X1 U20301 ( .C1(n9630), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n17136), .B(n17135), .ZN(n17137) );
  OAI211_X1 U20302 ( .C1(n17241), .C2(n17139), .A(n17138), .B(n17137), .ZN(
        n17140) );
  AOI211_X1 U20303 ( .C1(n17142), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n17141), .B(n17140), .ZN(n17385) );
  OAI22_X1 U20304 ( .A1(n17144), .A2(n17143), .B1(n17385), .B2(n17274), .ZN(
        P3_U2689) );
  OAI22_X1 U20305 ( .A1(n17227), .A2(n17145), .B1(n12100), .B2(n18525), .ZN(
        n17157) );
  AOI22_X1 U20306 ( .A1(n17229), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U20307 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17154) );
  INV_X1 U20308 ( .A(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17147) );
  AOI22_X1 U20309 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17146) );
  OAI21_X1 U20310 ( .B1(n17167), .B2(n17147), .A(n17146), .ZN(n17152) );
  AOI22_X1 U20311 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17150) );
  AOI22_X1 U20312 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17161), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17149) );
  OAI211_X1 U20313 ( .C1(n17235), .C2(n17266), .A(n17150), .B(n17149), .ZN(
        n17151) );
  AOI211_X1 U20314 ( .C1(n12616), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n17152), .B(n17151), .ZN(n17153) );
  NAND3_X1 U20315 ( .A1(n17155), .A2(n17154), .A3(n17153), .ZN(n17156) );
  AOI211_X1 U20316 ( .C1(n17225), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n17157), .B(n17156), .ZN(n17393) );
  AOI22_X1 U20317 ( .A1(n17291), .A2(n17158), .B1(P3_EBX_REG_12__SCAN_IN), 
        .B2(n17274), .ZN(n17159) );
  OAI22_X1 U20318 ( .A1(n17393), .A2(n17274), .B1(n17160), .B2(n17159), .ZN(
        P3_U2691) );
  AOI22_X1 U20319 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17176) );
  AOI22_X1 U20320 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17175) );
  OAI22_X1 U20321 ( .A1(n17163), .A2(n17162), .B1(n12100), .B2(n18522), .ZN(
        n17173) );
  AOI22_X1 U20322 ( .A1(n17204), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17209), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17170) );
  AOI22_X1 U20323 ( .A1(n17202), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17165) );
  AOI22_X1 U20324 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17225), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17164) );
  OAI211_X1 U20325 ( .C1(n17167), .C2(n17166), .A(n17165), .B(n17164), .ZN(
        n17168) );
  AOI21_X1 U20326 ( .B1(n12616), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n17168), .ZN(n17169) );
  OAI211_X1 U20327 ( .C1(n17241), .C2(n17171), .A(n17170), .B(n17169), .ZN(
        n17172) );
  AOI211_X1 U20328 ( .C1(n17230), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n17173), .B(n17172), .ZN(n17174) );
  NAND3_X1 U20329 ( .A1(n17176), .A2(n17175), .A3(n17174), .ZN(n17397) );
  INV_X1 U20330 ( .A(n17397), .ZN(n17180) );
  INV_X1 U20331 ( .A(n17177), .ZN(n17222) );
  NAND2_X1 U20332 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17249), .ZN(n17220) );
  INV_X1 U20333 ( .A(n17220), .ZN(n17198) );
  AND2_X1 U20334 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17198), .ZN(n17200) );
  OAI21_X1 U20335 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17200), .A(n17178), .ZN(
        n17179) );
  AOI22_X1 U20336 ( .A1(n17282), .A2(n17180), .B1(n17179), .B2(n17274), .ZN(
        P3_U2692) );
  AOI22_X1 U20337 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17196) );
  AOI22_X1 U20338 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17182) );
  OAI21_X1 U20339 ( .B1(n17184), .B2(n17183), .A(n17182), .ZN(n17194) );
  AOI22_X1 U20340 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17192) );
  INV_X1 U20341 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17189) );
  AOI22_X1 U20342 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17188) );
  AOI22_X1 U20343 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17187) );
  OAI211_X1 U20344 ( .C1(n17205), .C2(n17189), .A(n17188), .B(n17187), .ZN(
        n17190) );
  AOI21_X1 U20345 ( .B1(n9630), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n17190), .ZN(n17191) );
  OAI211_X1 U20346 ( .C1(n17235), .C2(n17276), .A(n17192), .B(n17191), .ZN(
        n17193) );
  AOI211_X1 U20347 ( .C1(n17202), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n17194), .B(n17193), .ZN(n17195) );
  OAI211_X1 U20348 ( .C1(n17227), .C2(n17197), .A(n17196), .B(n17195), .ZN(
        n17400) );
  INV_X1 U20349 ( .A(n17400), .ZN(n17201) );
  OAI21_X1 U20350 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17198), .A(n17274), .ZN(
        n17199) );
  OAI22_X1 U20351 ( .A1(n17201), .A2(n17274), .B1(n17200), .B2(n17199), .ZN(
        P3_U2693) );
  AOI22_X1 U20352 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9633), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17203) );
  OAI21_X1 U20353 ( .B1(n18516), .B2(n12100), .A(n17203), .ZN(n17219) );
  AOI22_X1 U20354 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17204), .B1(
        n17225), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17216) );
  OAI22_X1 U20355 ( .A1(n17208), .A2(n17207), .B1(n17206), .B2(n17205), .ZN(
        n17214) );
  AOI22_X1 U20356 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17223), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17229), .ZN(n17212) );
  AOI22_X1 U20357 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17161), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17211) );
  AOI22_X1 U20358 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n9630), .B1(
        n17209), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17210) );
  NAND3_X1 U20359 ( .A1(n17212), .A2(n17211), .A3(n17210), .ZN(n17213) );
  AOI211_X1 U20360 ( .C1(n17228), .C2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n17214), .B(n17213), .ZN(n17215) );
  OAI211_X1 U20361 ( .C1(n17217), .C2(n18601), .A(n17216), .B(n17215), .ZN(
        n17218) );
  AOI211_X1 U20362 ( .C1(n17101), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n17219), .B(n17218), .ZN(n17404) );
  OAI21_X1 U20363 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17249), .A(n17220), .ZN(
        n17221) );
  AOI22_X1 U20364 ( .A1(n17282), .A2(n17404), .B1(n17221), .B2(n17274), .ZN(
        P3_U2694) );
  OAI21_X1 U20365 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17222), .A(n17274), .ZN(
        n17248) );
  AOI22_X1 U20366 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17246) );
  AOI22_X1 U20367 ( .A1(n17225), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17161), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17245) );
  OAI22_X1 U20368 ( .A1(n17227), .A2(n17226), .B1(n12100), .B2(n18513), .ZN(
        n17243) );
  AOI22_X1 U20369 ( .A1(n12616), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17228), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17239) );
  AOI22_X1 U20370 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17233) );
  AOI22_X1 U20371 ( .A1(n17231), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17232) );
  OAI211_X1 U20372 ( .C1(n17235), .C2(n17234), .A(n17233), .B(n17232), .ZN(
        n17236) );
  AOI21_X1 U20373 ( .B1(n9630), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n17236), .ZN(n17238) );
  OAI211_X1 U20374 ( .C1(n17241), .C2(n17240), .A(n17239), .B(n17238), .ZN(
        n17242) );
  AOI211_X1 U20375 ( .C1(n9635), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n17243), .B(n17242), .ZN(n17244) );
  NAND3_X1 U20376 ( .A1(n17246), .A2(n17245), .A3(n17244), .ZN(n17408) );
  INV_X1 U20377 ( .A(n17408), .ZN(n17247) );
  OAI22_X1 U20378 ( .A1(n17249), .A2(n17248), .B1(n17247), .B2(n17274), .ZN(
        P3_U2695) );
  NAND2_X1 U20379 ( .A1(n17291), .A2(n17250), .ZN(n17252) );
  NOR2_X1 U20380 ( .A1(n17282), .A2(n17250), .ZN(n17253) );
  AOI22_X1 U20381 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17282), .B1(
        P3_EBX_REG_7__SCAN_IN), .B2(n17253), .ZN(n17251) );
  OAI21_X1 U20382 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17252), .A(n17251), .ZN(
        P3_U2696) );
  INV_X1 U20383 ( .A(n17257), .ZN(n17254) );
  OAI21_X1 U20384 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17254), .A(n17253), .ZN(
        n17255) );
  OAI21_X1 U20385 ( .B1(n17274), .B2(n17256), .A(n17255), .ZN(P3_U2697) );
  OAI21_X1 U20386 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17258), .A(n17257), .ZN(
        n17259) );
  AOI22_X1 U20387 ( .A1(n17282), .A2(n17260), .B1(n17259), .B2(n17274), .ZN(
        P3_U2698) );
  NAND2_X1 U20388 ( .A1(n17261), .A2(n17281), .ZN(n17272) );
  NOR2_X1 U20389 ( .A1(n17267), .A2(n17272), .ZN(n17271) );
  NOR2_X1 U20390 ( .A1(n17282), .A2(n17262), .ZN(n17264) );
  OAI22_X1 U20391 ( .A1(n17271), .A2(n17264), .B1(n17263), .B2(n17279), .ZN(
        n17265) );
  OAI21_X1 U20392 ( .B1(n17274), .B2(n17266), .A(n17265), .ZN(P3_U2699) );
  OAI21_X1 U20393 ( .B1(n17267), .B2(n17282), .A(n17272), .ZN(n17268) );
  INV_X1 U20394 ( .A(n17268), .ZN(n17270) );
  OAI22_X1 U20395 ( .A1(n17271), .A2(n17270), .B1(n17269), .B2(n17274), .ZN(
        P3_U2700) );
  OAI221_X1 U20396 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n17285), .C1(
        P3_EBX_REG_2__SCAN_IN), .C2(n17273), .A(n17272), .ZN(n17275) );
  AOI22_X1 U20397 ( .A1(n17282), .A2(n17276), .B1(n17275), .B2(n17274), .ZN(
        P3_U2701) );
  INV_X1 U20398 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17277) );
  AOI22_X1 U20399 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17282), .B1(
        n17281), .B2(n17284), .ZN(n17283) );
  OAI21_X1 U20400 ( .B1(n17285), .B2(n17284), .A(n17283), .ZN(P3_U2703) );
  INV_X1 U20401 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17511) );
  INV_X1 U20402 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17507) );
  INV_X1 U20403 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17552) );
  NAND2_X1 U20404 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n17440) );
  INV_X1 U20405 ( .A(n17440), .ZN(n17433) );
  NAND4_X1 U20406 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17286) );
  NOR2_X1 U20407 ( .A1(n17438), .A2(n17286), .ZN(n17287) );
  NAND4_X1 U20408 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(n17433), .A4(n17287), .ZN(n17410) );
  NAND4_X1 U20409 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .A4(P3_EAX_REG_10__SCAN_IN), .ZN(n17380)
         );
  NAND3_X1 U20410 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(P3_EAX_REG_14__SCAN_IN), .ZN(n17288) );
  NOR2_X2 U20411 ( .A1(n17552), .A2(n17382), .ZN(n17376) );
  INV_X1 U20412 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17493) );
  INV_X1 U20413 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17491) );
  NOR2_X1 U20414 ( .A1(n17493), .A2(n17491), .ZN(n17338) );
  NAND4_X1 U20415 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .A4(n17338), .ZN(n17337) );
  INV_X1 U20416 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17499) );
  NOR3_X2 U20417 ( .A1(n17372), .A2(n17337), .A3(n17499), .ZN(n17333) );
  NAND2_X1 U20418 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17333), .ZN(n17332) );
  NAND2_X1 U20419 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17328), .ZN(n17327) );
  NAND2_X1 U20420 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17305), .ZN(n17300) );
  NAND2_X1 U20421 ( .A1(n17296), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17295) );
  NAND2_X1 U20422 ( .A1(n17292), .A2(n17389), .ZN(n17369) );
  OAI22_X1 U20423 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17414), .B1(n17389), 
        .B2(n17296), .ZN(n17293) );
  AOI22_X1 U20424 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17370), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17293), .ZN(n17294) );
  OAI21_X1 U20425 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17295), .A(n17294), .ZN(
        P3_U2704) );
  NAND2_X1 U20426 ( .A1(n18286), .A2(n17389), .ZN(n17363) );
  AOI22_X1 U20427 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17371), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17370), .ZN(n17298) );
  OAI211_X1 U20428 ( .C1(n17296), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17432), .B(
        n17295), .ZN(n17297) );
  OAI211_X1 U20429 ( .C1(n17299), .C2(n17444), .A(n17298), .B(n17297), .ZN(
        P3_U2705) );
  AOI22_X1 U20430 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17371), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17370), .ZN(n17302) );
  OAI211_X1 U20431 ( .C1(n17305), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17432), .B(
        n17300), .ZN(n17301) );
  OAI211_X1 U20432 ( .C1(n17303), .C2(n17444), .A(n17302), .B(n17301), .ZN(
        P3_U2706) );
  INV_X1 U20433 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n17309) );
  AOI22_X1 U20434 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17371), .B1(n17409), .B2(
        n17304), .ZN(n17308) );
  AOI211_X1 U20435 ( .C1(n17511), .C2(n17313), .A(n17305), .B(n17389), .ZN(
        n17306) );
  INV_X1 U20436 ( .A(n17306), .ZN(n17307) );
  OAI211_X1 U20437 ( .C1(n17369), .C2(n17309), .A(n17308), .B(n17307), .ZN(
        P3_U2707) );
  OAI21_X1 U20438 ( .B1(n17312), .B2(n17311), .A(n17310), .ZN(n17316) );
  AOI22_X1 U20439 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17371), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17370), .ZN(n17315) );
  OAI211_X1 U20440 ( .C1(n17318), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17432), .B(
        n17313), .ZN(n17314) );
  OAI211_X1 U20441 ( .C1(n17316), .C2(n17444), .A(n17315), .B(n17314), .ZN(
        P3_U2708) );
  INV_X1 U20442 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n19260) );
  AOI22_X1 U20443 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17371), .B1(n17409), .B2(
        n17317), .ZN(n17321) );
  AOI211_X1 U20444 ( .C1(n17507), .C2(n17322), .A(n17318), .B(n17389), .ZN(
        n17319) );
  INV_X1 U20445 ( .A(n17319), .ZN(n17320) );
  OAI211_X1 U20446 ( .C1(n17369), .C2(n19260), .A(n17321), .B(n17320), .ZN(
        P3_U2709) );
  AOI22_X1 U20447 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17371), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17370), .ZN(n17325) );
  OAI211_X1 U20448 ( .C1(n17323), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17432), .B(
        n17322), .ZN(n17324) );
  OAI211_X1 U20449 ( .C1(n17326), .C2(n17444), .A(n17325), .B(n17324), .ZN(
        P3_U2710) );
  AOI22_X1 U20450 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17371), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17370), .ZN(n17330) );
  OAI211_X1 U20451 ( .C1(n17328), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17432), .B(
        n17327), .ZN(n17329) );
  OAI211_X1 U20452 ( .C1(n17331), .C2(n17444), .A(n17330), .B(n17329), .ZN(
        P3_U2711) );
  AOI22_X1 U20453 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17371), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17370), .ZN(n17335) );
  OAI211_X1 U20454 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17333), .A(n17432), .B(
        n17332), .ZN(n17334) );
  OAI211_X1 U20455 ( .C1(n17336), .C2(n17444), .A(n17335), .B(n17334), .ZN(
        P3_U2712) );
  INV_X1 U20456 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18289) );
  NOR3_X1 U20457 ( .A1(n18294), .A2(n17372), .A3(n17337), .ZN(n17342) );
  NAND2_X1 U20458 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17366), .ZN(n17365) );
  NAND2_X1 U20459 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17354), .ZN(n17349) );
  NAND2_X1 U20460 ( .A1(n17432), .A2(n17349), .ZN(n17345) );
  OAI21_X1 U20461 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17414), .A(n17345), .ZN(
        n17341) );
  INV_X1 U20462 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n19282) );
  OAI22_X1 U20463 ( .A1(n17339), .A2(n17444), .B1(n19282), .B2(n17369), .ZN(
        n17340) );
  AOI221_X1 U20464 ( .B1(n17342), .B2(n17499), .C1(n17341), .C2(
        P3_EAX_REG_22__SCAN_IN), .A(n17340), .ZN(n17343) );
  OAI21_X1 U20465 ( .B1(n18289), .B2(n17363), .A(n17343), .ZN(P3_U2713) );
  AOI22_X1 U20466 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17370), .B1(n17409), .B2(
        n17344), .ZN(n17348) );
  INV_X1 U20467 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18285) );
  INV_X1 U20468 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17497) );
  OAI22_X1 U20469 ( .A1(n18285), .A2(n17363), .B1(n17497), .B2(n17345), .ZN(
        n17346) );
  INV_X1 U20470 ( .A(n17346), .ZN(n17347) );
  OAI211_X1 U20471 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n17349), .A(n17348), .B(
        n17347), .ZN(P3_U2714) );
  AOI22_X1 U20472 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17371), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17370), .ZN(n17351) );
  OAI211_X1 U20473 ( .C1(n17354), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17432), .B(
        n17349), .ZN(n17350) );
  OAI211_X1 U20474 ( .C1(n17352), .C2(n17444), .A(n17351), .B(n17350), .ZN(
        P3_U2715) );
  AOI22_X1 U20475 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17371), .B1(n17409), .B2(
        n17353), .ZN(n17357) );
  NAND2_X1 U20476 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17360), .ZN(n17359) );
  AOI211_X1 U20477 ( .C1(n17493), .C2(n17359), .A(n17354), .B(n17389), .ZN(
        n17355) );
  INV_X1 U20478 ( .A(n17355), .ZN(n17356) );
  OAI211_X1 U20479 ( .C1(n17369), .C2(n13996), .A(n17357), .B(n17356), .ZN(
        P3_U2716) );
  INV_X1 U20480 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18272) );
  AOI22_X1 U20481 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17370), .B1(n17409), .B2(
        n17358), .ZN(n17362) );
  OAI211_X1 U20482 ( .C1(n17360), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17432), .B(
        n17359), .ZN(n17361) );
  OAI211_X1 U20483 ( .C1(n17363), .C2(n18272), .A(n17362), .B(n17361), .ZN(
        P3_U2717) );
  AOI22_X1 U20484 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17371), .B1(n17409), .B2(
        n17364), .ZN(n17368) );
  OAI211_X1 U20485 ( .C1(n17366), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17432), .B(
        n17365), .ZN(n17367) );
  OAI211_X1 U20486 ( .C1(n17369), .C2(n13902), .A(n17368), .B(n17367), .ZN(
        P3_U2718) );
  AOI22_X1 U20487 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17371), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17370), .ZN(n17374) );
  OAI211_X1 U20488 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17376), .A(n17432), .B(
        n17372), .ZN(n17373) );
  OAI211_X1 U20489 ( .C1(n17375), .C2(n17444), .A(n17374), .B(n17373), .ZN(
        P3_U2719) );
  AOI211_X1 U20490 ( .C1(n17552), .C2(n17382), .A(n17389), .B(n17376), .ZN(
        n17377) );
  AOI21_X1 U20491 ( .B1(n17439), .B2(BUF2_REG_15__SCAN_IN), .A(n17377), .ZN(
        n17378) );
  OAI21_X1 U20492 ( .B1(n17379), .B2(n17444), .A(n17378), .ZN(P3_U2720) );
  NOR2_X1 U20493 ( .A1(n18294), .A2(n17410), .ZN(n17417) );
  NAND3_X1 U20494 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(n17417), .ZN(n17402) );
  NOR3_X1 U20495 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17380), .A3(n17402), .ZN(
        n17381) );
  AOI21_X1 U20496 ( .B1(n17439), .B2(BUF2_REG_14__SCAN_IN), .A(n17381), .ZN(
        n17384) );
  NAND3_X1 U20497 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17432), .A3(n17382), 
        .ZN(n17383) );
  OAI211_X1 U20498 ( .C1(n17385), .C2(n17444), .A(n17384), .B(n17383), .ZN(
        P3_U2721) );
  NAND2_X1 U20499 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .ZN(n17386) );
  NOR2_X1 U20500 ( .A1(n17386), .A2(n17402), .ZN(n17392) );
  NAND2_X1 U20501 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17392), .ZN(n17391) );
  NAND2_X1 U20502 ( .A1(n17391), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n17390) );
  AOI22_X1 U20503 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17439), .B1(n17409), .B2(
        n17387), .ZN(n17388) );
  OAI221_X1 U20504 ( .B1(n17391), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n17390), 
        .C2(n17389), .A(n17388), .ZN(P3_U2722) );
  INV_X1 U20505 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17396) );
  INV_X1 U20506 ( .A(n17391), .ZN(n17395) );
  AOI21_X1 U20507 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17432), .A(n17392), .ZN(
        n17394) );
  OAI222_X1 U20508 ( .A1(n17437), .A2(n17396), .B1(n17395), .B2(n17394), .C1(
        n17444), .C2(n17393), .ZN(P3_U2723) );
  INV_X1 U20509 ( .A(n17402), .ZN(n17406) );
  NAND2_X1 U20510 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17406), .ZN(n17399) );
  INV_X1 U20511 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17539) );
  INV_X1 U20512 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17537) );
  OAI21_X1 U20513 ( .B1(n17537), .B2(n17402), .A(n17432), .ZN(n17403) );
  AOI22_X1 U20514 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17439), .B1(n17409), .B2(
        n17397), .ZN(n17398) );
  OAI221_X1 U20515 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17399), .C1(n17539), 
        .C2(n17403), .A(n17398), .ZN(P3_U2724) );
  AOI22_X1 U20516 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17439), .B1(n17409), .B2(
        n17400), .ZN(n17401) );
  OAI221_X1 U20517 ( .B1(n17403), .B2(n17537), .C1(n17403), .C2(n17402), .A(
        n17401), .ZN(P3_U2725) );
  INV_X1 U20518 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17407) );
  AOI22_X1 U20519 ( .A1(n17417), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17432), .ZN(n17405) );
  OAI222_X1 U20520 ( .A1(n17437), .A2(n17407), .B1(n17406), .B2(n17405), .C1(
        n17444), .C2(n17404), .ZN(P3_U2726) );
  INV_X1 U20521 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17413) );
  INV_X1 U20522 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17533) );
  AOI22_X1 U20523 ( .A1(n17409), .A2(n17408), .B1(n17417), .B2(n17533), .ZN(
        n17412) );
  NAND3_X1 U20524 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17432), .A3(n17410), .ZN(
        n17411) );
  OAI211_X1 U20525 ( .C1(n17437), .C2(n17413), .A(n17412), .B(n17411), .ZN(
        P3_U2727) );
  INV_X1 U20526 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18296) );
  INV_X1 U20527 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17529) );
  INV_X1 U20528 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17525) );
  INV_X1 U20529 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17521) );
  NAND2_X1 U20530 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17436), .ZN(n17425) );
  NOR2_X1 U20531 ( .A1(n17525), .A2(n17425), .ZN(n17428) );
  NAND2_X1 U20532 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17428), .ZN(n17418) );
  NOR2_X1 U20533 ( .A1(n17529), .A2(n17418), .ZN(n17421) );
  AOI21_X1 U20534 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17432), .A(n17421), .ZN(
        n17416) );
  OAI222_X1 U20535 ( .A1(n17437), .A2(n18296), .B1(n17417), .B2(n17416), .C1(
        n17444), .C2(n17415), .ZN(P3_U2728) );
  INV_X1 U20536 ( .A(n17418), .ZN(n17424) );
  AOI21_X1 U20537 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17432), .A(n17424), .ZN(
        n17420) );
  OAI222_X1 U20538 ( .A1(n18289), .A2(n17437), .B1(n17421), .B2(n17420), .C1(
        n17444), .C2(n17419), .ZN(P3_U2729) );
  AOI21_X1 U20539 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17432), .A(n17428), .ZN(
        n17423) );
  OAI222_X1 U20540 ( .A1(n18285), .A2(n17437), .B1(n17424), .B2(n17423), .C1(
        n17444), .C2(n17422), .ZN(P3_U2730) );
  INV_X1 U20541 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18280) );
  INV_X1 U20542 ( .A(n17425), .ZN(n17431) );
  AOI21_X1 U20543 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17432), .A(n17431), .ZN(
        n17427) );
  OAI222_X1 U20544 ( .A1(n18280), .A2(n17437), .B1(n17428), .B2(n17427), .C1(
        n17444), .C2(n17426), .ZN(P3_U2731) );
  INV_X1 U20545 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18276) );
  AOI21_X1 U20546 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17432), .A(n17436), .ZN(
        n17430) );
  OAI222_X1 U20547 ( .A1(n18276), .A2(n17437), .B1(n17431), .B2(n17430), .C1(
        n17444), .C2(n17429), .ZN(P3_U2732) );
  AOI22_X1 U20548 ( .A1(n17441), .A2(n17433), .B1(P3_EAX_REG_2__SCAN_IN), .B2(
        n17432), .ZN(n17435) );
  OAI222_X1 U20549 ( .A1(n18272), .A2(n17437), .B1(n17436), .B2(n17435), .C1(
        n17444), .C2(n17434), .ZN(P3_U2733) );
  AOI22_X1 U20550 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17439), .B1(
        P3_EAX_REG_1__SCAN_IN), .B2(n17438), .ZN(n17443) );
  OAI211_X1 U20551 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(P3_EAX_REG_0__SCAN_IN), 
        .A(n17441), .B(n17440), .ZN(n17442) );
  OAI211_X1 U20552 ( .C1(n17445), .C2(n17444), .A(n17443), .B(n17442), .ZN(
        P3_U2734) );
  NOR2_X2 U20553 ( .A1(n18905), .A2(n18791), .ZN(n18929) );
  NOR2_X4 U20554 ( .A1(n18929), .A2(n17464), .ZN(n17461) );
  AND2_X1 U20555 ( .A1(n17461), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20556 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17515) );
  NAND2_X1 U20557 ( .A1(n17464), .A2(n18267), .ZN(n17463) );
  AOI22_X1 U20558 ( .A1(n18929), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17461), .ZN(n17447) );
  OAI21_X1 U20559 ( .B1(n17515), .B2(n17463), .A(n17447), .ZN(P3_U2737) );
  INV_X1 U20560 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17513) );
  AOI22_X1 U20561 ( .A1(n18929), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17448) );
  OAI21_X1 U20562 ( .B1(n17513), .B2(n17463), .A(n17448), .ZN(P3_U2738) );
  AOI22_X1 U20563 ( .A1(n18929), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17449) );
  OAI21_X1 U20564 ( .B1(n17511), .B2(n17463), .A(n17449), .ZN(P3_U2739) );
  INV_X1 U20565 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17509) );
  AOI22_X1 U20566 ( .A1(n18929), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17450) );
  OAI21_X1 U20567 ( .B1(n17509), .B2(n17463), .A(n17450), .ZN(P3_U2740) );
  AOI22_X1 U20568 ( .A1(n18929), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17451) );
  OAI21_X1 U20569 ( .B1(n17507), .B2(n17463), .A(n17451), .ZN(P3_U2741) );
  INV_X1 U20570 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17505) );
  AOI22_X1 U20571 ( .A1(n18929), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17452) );
  OAI21_X1 U20572 ( .B1(n17505), .B2(n17463), .A(n17452), .ZN(P3_U2742) );
  INV_X1 U20573 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17503) );
  AOI22_X1 U20574 ( .A1(n18929), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17453) );
  OAI21_X1 U20575 ( .B1(n17503), .B2(n17463), .A(n17453), .ZN(P3_U2743) );
  INV_X1 U20576 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17501) );
  CLKBUF_X1 U20577 ( .A(n18929), .Z(n17480) );
  AOI22_X1 U20578 ( .A1(n17480), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17454) );
  OAI21_X1 U20579 ( .B1(n17501), .B2(n17463), .A(n17454), .ZN(P3_U2744) );
  AOI22_X1 U20580 ( .A1(n17480), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17455) );
  OAI21_X1 U20581 ( .B1(n17499), .B2(n17463), .A(n17455), .ZN(P3_U2745) );
  AOI22_X1 U20582 ( .A1(n17480), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17456) );
  OAI21_X1 U20583 ( .B1(n17497), .B2(n17463), .A(n17456), .ZN(P3_U2746) );
  INV_X1 U20584 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17495) );
  AOI22_X1 U20585 ( .A1(n17480), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17457) );
  OAI21_X1 U20586 ( .B1(n17495), .B2(n17463), .A(n17457), .ZN(P3_U2747) );
  AOI22_X1 U20587 ( .A1(n17480), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17458) );
  OAI21_X1 U20588 ( .B1(n17493), .B2(n17463), .A(n17458), .ZN(P3_U2748) );
  AOI22_X1 U20589 ( .A1(n17480), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17459) );
  OAI21_X1 U20590 ( .B1(n17491), .B2(n17463), .A(n17459), .ZN(P3_U2749) );
  INV_X1 U20591 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17489) );
  AOI22_X1 U20592 ( .A1(n17480), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17460) );
  OAI21_X1 U20593 ( .B1(n17489), .B2(n17463), .A(n17460), .ZN(P3_U2750) );
  INV_X1 U20594 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17487) );
  AOI22_X1 U20595 ( .A1(n17480), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17462) );
  OAI21_X1 U20596 ( .B1(n17487), .B2(n17463), .A(n17462), .ZN(P3_U2751) );
  AOI22_X1 U20597 ( .A1(n17480), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17465) );
  OAI21_X1 U20598 ( .B1(n17552), .B2(n17482), .A(n17465), .ZN(P3_U2752) );
  INV_X1 U20599 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17547) );
  AOI22_X1 U20600 ( .A1(n17480), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17466) );
  OAI21_X1 U20601 ( .B1(n17547), .B2(n17482), .A(n17466), .ZN(P3_U2753) );
  INV_X1 U20602 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17544) );
  AOI22_X1 U20603 ( .A1(n17480), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17467) );
  OAI21_X1 U20604 ( .B1(n17544), .B2(n17482), .A(n17467), .ZN(P3_U2754) );
  INV_X1 U20605 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17542) );
  AOI22_X1 U20606 ( .A1(n17480), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17468) );
  OAI21_X1 U20607 ( .B1(n17542), .B2(n17482), .A(n17468), .ZN(P3_U2755) );
  AOI22_X1 U20608 ( .A1(n17480), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17469) );
  OAI21_X1 U20609 ( .B1(n17539), .B2(n17482), .A(n17469), .ZN(P3_U2756) );
  AOI22_X1 U20610 ( .A1(n17480), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17470) );
  OAI21_X1 U20611 ( .B1(n17537), .B2(n17482), .A(n17470), .ZN(P3_U2757) );
  INV_X1 U20612 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17535) );
  AOI22_X1 U20613 ( .A1(n17480), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17471) );
  OAI21_X1 U20614 ( .B1(n17535), .B2(n17482), .A(n17471), .ZN(P3_U2758) );
  AOI22_X1 U20615 ( .A1(n17480), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17472) );
  OAI21_X1 U20616 ( .B1(n17533), .B2(n17482), .A(n17472), .ZN(P3_U2759) );
  INV_X1 U20617 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17531) );
  AOI22_X1 U20618 ( .A1(n17480), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17473) );
  OAI21_X1 U20619 ( .B1(n17531), .B2(n17482), .A(n17473), .ZN(P3_U2760) );
  AOI22_X1 U20620 ( .A1(n17480), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17474) );
  OAI21_X1 U20621 ( .B1(n17529), .B2(n17482), .A(n17474), .ZN(P3_U2761) );
  INV_X1 U20622 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17527) );
  AOI22_X1 U20623 ( .A1(n17480), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17475) );
  OAI21_X1 U20624 ( .B1(n17527), .B2(n17482), .A(n17475), .ZN(P3_U2762) );
  AOI22_X1 U20625 ( .A1(n17480), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17476) );
  OAI21_X1 U20626 ( .B1(n17525), .B2(n17482), .A(n17476), .ZN(P3_U2763) );
  INV_X1 U20627 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17523) );
  AOI22_X1 U20628 ( .A1(n17480), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17477) );
  OAI21_X1 U20629 ( .B1(n17523), .B2(n17482), .A(n17477), .ZN(P3_U2764) );
  AOI22_X1 U20630 ( .A1(n17480), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17478) );
  OAI21_X1 U20631 ( .B1(n17521), .B2(n17482), .A(n17478), .ZN(P3_U2765) );
  INV_X1 U20632 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17519) );
  AOI22_X1 U20633 ( .A1(n17480), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17479) );
  OAI21_X1 U20634 ( .B1(n17519), .B2(n17482), .A(n17479), .ZN(P3_U2766) );
  AOI22_X1 U20635 ( .A1(n17480), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17461), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17481) );
  OAI21_X1 U20636 ( .B1(n17517), .B2(n17482), .A(n17481), .ZN(P3_U2767) );
  NAND2_X1 U20637 ( .A1(n18932), .A2(n17485), .ZN(n18775) );
  AOI22_X1 U20638 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17549), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17548), .ZN(n17486) );
  OAI21_X1 U20639 ( .B1(n17487), .B2(n17551), .A(n17486), .ZN(P3_U2768) );
  AOI22_X1 U20640 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17549), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17548), .ZN(n17488) );
  OAI21_X1 U20641 ( .B1(n17489), .B2(n17551), .A(n17488), .ZN(P3_U2769) );
  AOI22_X1 U20642 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17549), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17548), .ZN(n17490) );
  OAI21_X1 U20643 ( .B1(n17491), .B2(n17551), .A(n17490), .ZN(P3_U2770) );
  AOI22_X1 U20644 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17540), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17548), .ZN(n17492) );
  OAI21_X1 U20645 ( .B1(n17493), .B2(n17551), .A(n17492), .ZN(P3_U2771) );
  AOI22_X1 U20646 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17540), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17548), .ZN(n17494) );
  OAI21_X1 U20647 ( .B1(n17495), .B2(n17551), .A(n17494), .ZN(P3_U2772) );
  AOI22_X1 U20648 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17540), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17548), .ZN(n17496) );
  OAI21_X1 U20649 ( .B1(n17497), .B2(n17551), .A(n17496), .ZN(P3_U2773) );
  AOI22_X1 U20650 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17540), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17548), .ZN(n17498) );
  OAI21_X1 U20651 ( .B1(n17499), .B2(n17551), .A(n17498), .ZN(P3_U2774) );
  AOI22_X1 U20652 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17540), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17548), .ZN(n17500) );
  OAI21_X1 U20653 ( .B1(n17501), .B2(n17551), .A(n17500), .ZN(P3_U2775) );
  AOI22_X1 U20654 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17540), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17548), .ZN(n17502) );
  OAI21_X1 U20655 ( .B1(n17503), .B2(n17551), .A(n17502), .ZN(P3_U2776) );
  AOI22_X1 U20656 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17540), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17548), .ZN(n17504) );
  OAI21_X1 U20657 ( .B1(n17505), .B2(n17551), .A(n17504), .ZN(P3_U2777) );
  AOI22_X1 U20658 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17540), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17548), .ZN(n17506) );
  OAI21_X1 U20659 ( .B1(n17507), .B2(n17551), .A(n17506), .ZN(P3_U2778) );
  AOI22_X1 U20660 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17540), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17548), .ZN(n17508) );
  OAI21_X1 U20661 ( .B1(n17509), .B2(n17551), .A(n17508), .ZN(P3_U2779) );
  AOI22_X1 U20662 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17549), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17548), .ZN(n17510) );
  OAI21_X1 U20663 ( .B1(n17511), .B2(n17551), .A(n17510), .ZN(P3_U2780) );
  AOI22_X1 U20664 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17549), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17548), .ZN(n17512) );
  OAI21_X1 U20665 ( .B1(n17513), .B2(n17551), .A(n17512), .ZN(P3_U2781) );
  AOI22_X1 U20666 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17549), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17548), .ZN(n17514) );
  OAI21_X1 U20667 ( .B1(n17515), .B2(n17551), .A(n17514), .ZN(P3_U2782) );
  AOI22_X1 U20668 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17549), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17548), .ZN(n17516) );
  OAI21_X1 U20669 ( .B1(n17517), .B2(n17551), .A(n17516), .ZN(P3_U2783) );
  AOI22_X1 U20670 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17549), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17548), .ZN(n17518) );
  OAI21_X1 U20671 ( .B1(n17519), .B2(n17551), .A(n17518), .ZN(P3_U2784) );
  AOI22_X1 U20672 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17549), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17548), .ZN(n17520) );
  OAI21_X1 U20673 ( .B1(n17521), .B2(n17551), .A(n17520), .ZN(P3_U2785) );
  AOI22_X1 U20674 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17549), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17545), .ZN(n17522) );
  OAI21_X1 U20675 ( .B1(n17523), .B2(n17551), .A(n17522), .ZN(P3_U2786) );
  AOI22_X1 U20676 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17549), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17545), .ZN(n17524) );
  OAI21_X1 U20677 ( .B1(n17525), .B2(n17551), .A(n17524), .ZN(P3_U2787) );
  AOI22_X1 U20678 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17549), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17545), .ZN(n17526) );
  OAI21_X1 U20679 ( .B1(n17527), .B2(n17551), .A(n17526), .ZN(P3_U2788) );
  AOI22_X1 U20680 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17549), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17545), .ZN(n17528) );
  OAI21_X1 U20681 ( .B1(n17529), .B2(n17551), .A(n17528), .ZN(P3_U2789) );
  AOI22_X1 U20682 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17549), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17545), .ZN(n17530) );
  OAI21_X1 U20683 ( .B1(n17531), .B2(n17551), .A(n17530), .ZN(P3_U2790) );
  AOI22_X1 U20684 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17549), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17545), .ZN(n17532) );
  OAI21_X1 U20685 ( .B1(n17533), .B2(n17551), .A(n17532), .ZN(P3_U2791) );
  AOI22_X1 U20686 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17549), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17545), .ZN(n17534) );
  OAI21_X1 U20687 ( .B1(n17535), .B2(n17551), .A(n17534), .ZN(P3_U2792) );
  AOI22_X1 U20688 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17540), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17548), .ZN(n17536) );
  OAI21_X1 U20689 ( .B1(n17537), .B2(n17551), .A(n17536), .ZN(P3_U2793) );
  AOI22_X1 U20690 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17549), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17545), .ZN(n17538) );
  OAI21_X1 U20691 ( .B1(n17539), .B2(n17551), .A(n17538), .ZN(P3_U2794) );
  AOI22_X1 U20692 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17540), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17548), .ZN(n17541) );
  OAI21_X1 U20693 ( .B1(n17542), .B2(n17551), .A(n17541), .ZN(P3_U2795) );
  AOI22_X1 U20694 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17549), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17545), .ZN(n17543) );
  OAI21_X1 U20695 ( .B1(n17544), .B2(n17551), .A(n17543), .ZN(P3_U2796) );
  AOI22_X1 U20696 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17549), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17545), .ZN(n17546) );
  OAI21_X1 U20697 ( .B1(n17547), .B2(n17551), .A(n17546), .ZN(P3_U2797) );
  AOI22_X1 U20698 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17549), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17548), .ZN(n17550) );
  OAI21_X1 U20699 ( .B1(n17552), .B2(n17551), .A(n17550), .ZN(P3_U2798) );
  AOI21_X1 U20700 ( .B1(n17770), .B2(n17554), .A(n17553), .ZN(n17570) );
  NOR2_X1 U20701 ( .A1(n17902), .A2(n17828), .ZN(n17671) );
  OAI22_X1 U20702 ( .A1(n17920), .A2(n17916), .B1(n17919), .B2(n17758), .ZN(
        n17589) );
  NOR2_X1 U20703 ( .A1(n17918), .A2(n17589), .ZN(n17577) );
  NOR3_X1 U20704 ( .A1(n17671), .A2(n17577), .A3(n17555), .ZN(n17560) );
  AOI211_X1 U20705 ( .C1(n17558), .C2(n17557), .A(n17556), .B(n17831), .ZN(
        n17559) );
  AOI211_X1 U20706 ( .C1(n17561), .C2(n17718), .A(n17560), .B(n17559), .ZN(
        n17569) );
  NOR3_X1 U20707 ( .A1(n17722), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        n17564), .ZN(n17579) );
  OAI21_X1 U20708 ( .B1(n17562), .B2(n18791), .A(n17912), .ZN(n17563) );
  AOI21_X1 U20709 ( .B1(n17820), .B2(n17564), .A(n17563), .ZN(n17593) );
  OAI21_X1 U20710 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17665), .A(
        n17593), .ZN(n17580) );
  OAI21_X1 U20711 ( .B1(n17579), .B2(n17580), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17568) );
  NAND3_X1 U20712 ( .A1(n17566), .A2(n17748), .A3(n17565), .ZN(n17567) );
  NAND4_X1 U20713 ( .A1(n17570), .A2(n17569), .A3(n17568), .A4(n17567), .ZN(
        P3_U2802) );
  NOR2_X1 U20714 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17571), .ZN(
        n17576) );
  INV_X1 U20715 ( .A(n17572), .ZN(n17573) );
  NAND2_X1 U20716 ( .A1(n17574), .A2(n17573), .ZN(n17575) );
  XOR2_X1 U20717 ( .A(n17815), .B(n17575), .Z(n17932) );
  OAI22_X1 U20718 ( .A1(n17577), .A2(n17576), .B1(n17932), .B2(n17831), .ZN(
        n17578) );
  AOI211_X1 U20719 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17580), .A(
        n17579), .B(n17578), .ZN(n17581) );
  NAND2_X1 U20720 ( .A1(n18071), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17930) );
  OAI211_X1 U20721 ( .C1(n17754), .C2(n17582), .A(n17581), .B(n17930), .ZN(
        P3_U2803) );
  AOI21_X1 U20722 ( .B1(n18304), .B2(n17583), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17592) );
  NAND2_X1 U20723 ( .A1(n17754), .A2(n17665), .ZN(n17696) );
  AOI22_X1 U20724 ( .A1(n18071), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n17584), 
        .B2(n17696), .ZN(n17591) );
  AOI21_X1 U20725 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17586), .A(
        n17585), .ZN(n17938) );
  NAND3_X1 U20726 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17598), .A3(
        n10019), .ZN(n17934) );
  OAI22_X1 U20727 ( .A1(n17938), .A2(n17831), .B1(n17587), .B2(n17934), .ZN(
        n17588) );
  AOI21_X1 U20728 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17589), .A(
        n17588), .ZN(n17590) );
  OAI211_X1 U20729 ( .C1(n17593), .C2(n17592), .A(n17591), .B(n17590), .ZN(
        P3_U2804) );
  INV_X1 U20730 ( .A(n18791), .ZN(n17636) );
  OAI21_X1 U20731 ( .B1(n17594), .B2(n18592), .A(n17912), .ZN(n17595) );
  AOI21_X1 U20732 ( .B1(n17636), .B2(n17596), .A(n17595), .ZN(n17621) );
  OAI21_X1 U20733 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17665), .A(
        n17621), .ZN(n17615) );
  AOI22_X1 U20734 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17615), .B1(
        n17770), .B2(n17597), .ZN(n17609) );
  NAND2_X1 U20735 ( .A1(n17598), .A2(n17974), .ZN(n17599) );
  XOR2_X1 U20736 ( .A(n17599), .B(n17939), .Z(n17951) );
  XOR2_X1 U20737 ( .A(n17600), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17953) );
  OAI21_X1 U20738 ( .B1(n17815), .B2(n17602), .A(n17601), .ZN(n17603) );
  XOR2_X1 U20739 ( .A(n17603), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17949) );
  OAI22_X1 U20740 ( .A1(n17916), .A2(n17953), .B1(n17831), .B2(n17949), .ZN(
        n17604) );
  AOI21_X1 U20741 ( .B1(n17828), .B2(n17951), .A(n17604), .ZN(n17608) );
  NAND2_X1 U20742 ( .A1(n18071), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17947) );
  NOR2_X1 U20743 ( .A1(n17722), .A2(n17605), .ZN(n17617) );
  OAI211_X1 U20744 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17617), .B(n17606), .ZN(n17607) );
  NAND4_X1 U20745 ( .A1(n17609), .A2(n17608), .A3(n17947), .A4(n17607), .ZN(
        P3_U2805) );
  AOI21_X1 U20746 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17611), .A(
        n17610), .ZN(n17966) );
  INV_X1 U20747 ( .A(n17612), .ZN(n17613) );
  OAI22_X1 U20748 ( .A1(n18140), .A2(n18856), .B1(n17754), .B2(n17613), .ZN(
        n17614) );
  AOI221_X1 U20749 ( .B1(n17617), .B2(n17616), .C1(n17615), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17614), .ZN(n17620) );
  NOR2_X1 U20750 ( .A1(n17618), .A2(n18062), .ZN(n17954) );
  OAI22_X1 U20751 ( .A1(n17955), .A2(n17916), .B1(n17954), .B2(n17758), .ZN(
        n17630) );
  NOR2_X1 U20752 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17618), .ZN(
        n17963) );
  AOI22_X1 U20753 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17630), .B1(
        n17718), .B2(n17963), .ZN(n17619) );
  OAI211_X1 U20754 ( .C1(n17966), .C2(n17831), .A(n17620), .B(n17619), .ZN(
        P3_U2806) );
  AOI221_X1 U20755 ( .B1(n17623), .B2(n17622), .C1(n18592), .C2(n17622), .A(
        n17621), .ZN(n17624) );
  AOI221_X1 U20756 ( .B1(n17770), .B2(n17625), .C1(n17664), .C2(n17625), .A(
        n17624), .ZN(n17634) );
  AOI22_X1 U20757 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17815), .B1(
        n17627), .B2(n17644), .ZN(n17628) );
  NAND2_X1 U20758 ( .A1(n17626), .A2(n17628), .ZN(n17629) );
  XOR2_X1 U20759 ( .A(n17629), .B(n17631), .Z(n17967) );
  AOI22_X1 U20760 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17630), .B1(
        n17810), .B2(n17967), .ZN(n17633) );
  NAND4_X1 U20761 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17984), .A3(
        n17718), .A4(n17631), .ZN(n17632) );
  NAND2_X1 U20762 ( .A1(n18071), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17972) );
  NAND4_X1 U20763 ( .A1(n17634), .A2(n17633), .A3(n17632), .A4(n17972), .ZN(
        P3_U2807) );
  NAND2_X1 U20764 ( .A1(n17984), .A2(n17718), .ZN(n17649) );
  NAND2_X1 U20765 ( .A1(n17638), .A2(n17748), .ZN(n17652) );
  AOI221_X1 U20766 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n17651), .C2(n17639), .A(
        n17652), .ZN(n17641) );
  NAND2_X1 U20767 ( .A1(n17636), .A2(n17635), .ZN(n17637) );
  OAI211_X1 U20768 ( .C1(n17638), .C2(n17750), .A(n17912), .B(n17637), .ZN(
        n17669) );
  AOI21_X1 U20769 ( .B1(n17664), .B2(n17662), .A(n17669), .ZN(n17650) );
  OAI22_X1 U20770 ( .A1(n17650), .A2(n17639), .B1(n18140), .B2(n18852), .ZN(
        n17640) );
  AOI211_X1 U20771 ( .C1(n17642), .C2(n17770), .A(n17641), .B(n17640), .ZN(
        n17648) );
  INV_X1 U20772 ( .A(n17720), .ZN(n18067) );
  OAI22_X1 U20773 ( .A1(n17916), .A2(n18067), .B1(n17758), .B2(n17974), .ZN(
        n17717) );
  INV_X1 U20774 ( .A(n17717), .ZN(n17670) );
  OAI21_X1 U20775 ( .B1(n17984), .B2(n17671), .A(n17670), .ZN(n17659) );
  INV_X1 U20776 ( .A(n17626), .ZN(n17643) );
  AOI221_X1 U20777 ( .B1(n17645), .B2(n17644), .C1(n17655), .C2(n17644), .A(
        n17643), .ZN(n17646) );
  XOR2_X1 U20778 ( .A(n17646), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(
        n17989) );
  AOI22_X1 U20779 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17659), .B1(
        n17810), .B2(n17989), .ZN(n17647) );
  OAI211_X1 U20780 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17649), .A(
        n17648), .B(n17647), .ZN(P3_U2808) );
  NAND2_X1 U20781 ( .A1(n17980), .A2(n18000), .ZN(n18006) );
  NAND2_X1 U20782 ( .A1(n18028), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17996) );
  INV_X1 U20783 ( .A(n17996), .ZN(n17993) );
  NAND2_X1 U20784 ( .A1(n17718), .A2(n17993), .ZN(n17684) );
  NAND2_X1 U20785 ( .A1(n18071), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18004) );
  OAI221_X1 U20786 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17652), .C1(
        n17651), .C2(n17650), .A(n18004), .ZN(n17653) );
  AOI21_X1 U20787 ( .B1(n17770), .B2(n17654), .A(n17653), .ZN(n17661) );
  INV_X1 U20788 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17977) );
  NOR3_X1 U20789 ( .A1(n17977), .A2(n17815), .A3(n17655), .ZN(n17679) );
  INV_X1 U20790 ( .A(n17656), .ZN(n17691) );
  AOI22_X1 U20791 ( .A1(n17980), .A2(n17679), .B1(n17691), .B2(n17657), .ZN(
        n17658) );
  XOR2_X1 U20792 ( .A(n18000), .B(n17658), .Z(n18003) );
  AOI22_X1 U20793 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17659), .B1(
        n17810), .B2(n18003), .ZN(n17660) );
  OAI211_X1 U20794 ( .C1(n18006), .C2(n17684), .A(n17661), .B(n17660), .ZN(
        P3_U2809) );
  INV_X1 U20795 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17978) );
  NAND2_X1 U20796 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17978), .ZN(
        n18016) );
  OAI21_X1 U20797 ( .B1(n18592), .B2(n17663), .A(n17662), .ZN(n17668) );
  INV_X1 U20798 ( .A(n17664), .ZN(n17665) );
  NAND2_X1 U20799 ( .A1(n18071), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18014) );
  OAI221_X1 U20800 ( .B1(n17666), .B2(n17754), .C1(n17666), .C2(n17665), .A(
        n18014), .ZN(n17667) );
  AOI21_X1 U20801 ( .B1(n17669), .B2(n17668), .A(n17667), .ZN(n17674) );
  NOR2_X1 U20802 ( .A1(n18021), .A2(n17996), .ZN(n18008) );
  OAI21_X1 U20803 ( .B1(n17671), .B2(n18008), .A(n17670), .ZN(n17681) );
  OAI221_X1 U20804 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17690), 
        .C1(n18021), .C2(n17679), .A(n17626), .ZN(n17672) );
  XOR2_X1 U20805 ( .A(n17978), .B(n17672), .Z(n18012) );
  AOI22_X1 U20806 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17681), .B1(
        n17810), .B2(n18012), .ZN(n17673) );
  OAI211_X1 U20807 ( .C1(n17684), .C2(n18016), .A(n17674), .B(n17673), .ZN(
        P3_U2810) );
  AOI21_X1 U20808 ( .B1(n17820), .B2(n9887), .A(n17818), .ZN(n17697) );
  OAI21_X1 U20809 ( .B1(n17675), .B2(n18791), .A(n17697), .ZN(n17687) );
  INV_X1 U20810 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18846) );
  NOR2_X1 U20811 ( .A1(n18140), .A2(n18846), .ZN(n18017) );
  OAI211_X1 U20812 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n16710), .B(n17748), .ZN(n17677) );
  OAI22_X1 U20813 ( .A1(n10169), .A2(n17677), .B1(n17676), .B2(n17754), .ZN(
        n17678) );
  AOI211_X1 U20814 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n17687), .A(
        n18017), .B(n17678), .ZN(n17683) );
  AOI21_X1 U20815 ( .B1(n17690), .B2(n17691), .A(n17679), .ZN(n17680) );
  XOR2_X1 U20816 ( .A(n18021), .B(n17680), .Z(n18018) );
  AOI22_X1 U20817 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17681), .B1(
        n17810), .B2(n18018), .ZN(n17682) );
  OAI211_X1 U20818 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17684), .A(
        n17683), .B(n17682), .ZN(P3_U2811) );
  AOI21_X1 U20819 ( .B1(n17718), .B2(n17693), .A(n17717), .ZN(n17707) );
  NOR2_X1 U20820 ( .A1(n17722), .A2(n9887), .ZN(n17689) );
  INV_X1 U20821 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17688) );
  OAI22_X1 U20822 ( .A1(n18140), .A2(n18844), .B1(n17754), .B2(n17685), .ZN(
        n17686) );
  AOI221_X1 U20823 ( .B1(n17689), .B2(n17688), .C1(n17687), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17686), .ZN(n17695) );
  AOI21_X1 U20824 ( .B1(n10022), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17690), .ZN(n17692) );
  XOR2_X1 U20825 ( .A(n17692), .B(n17691), .Z(n18037) );
  NOR2_X1 U20826 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17693), .ZN(
        n18036) );
  AOI22_X1 U20827 ( .A1(n17810), .A2(n18037), .B1(n17718), .B2(n18036), .ZN(
        n17694) );
  OAI211_X1 U20828 ( .C1(n17707), .C2(n17977), .A(n17695), .B(n17694), .ZN(
        P3_U2812) );
  NOR2_X1 U20829 ( .A1(n18140), .A2(n18843), .ZN(n17701) );
  AOI221_X1 U20830 ( .B1(n18592), .B2(n17699), .C1(n17698), .C2(n17699), .A(
        n17697), .ZN(n17700) );
  AOI211_X1 U20831 ( .C1(n17702), .C2(n17696), .A(n17701), .B(n17700), .ZN(
        n17706) );
  OAI21_X1 U20832 ( .B1(n17704), .B2(n18029), .A(n17703), .ZN(n18042) );
  NOR2_X1 U20833 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18053), .ZN(
        n18041) );
  AOI22_X1 U20834 ( .A1(n17810), .A2(n18042), .B1(n17718), .B2(n18041), .ZN(
        n17705) );
  OAI211_X1 U20835 ( .C1(n17707), .C2(n18029), .A(n17706), .B(n17705), .ZN(
        P3_U2813) );
  NOR2_X1 U20836 ( .A1(n17815), .A2(n17708), .ZN(n17795) );
  OAI22_X1 U20837 ( .A1(n10022), .A2(n17709), .B1(n17803), .B2(n18035), .ZN(
        n17710) );
  XOR2_X1 U20838 ( .A(n18053), .B(n17710), .Z(n18058) );
  OAI211_X1 U20839 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17711), .B(n17748), .ZN(n17715) );
  INV_X1 U20840 ( .A(n17711), .ZN(n17721) );
  AOI21_X1 U20841 ( .B1(n17820), .B2(n17721), .A(n17818), .ZN(n17738) );
  OAI21_X1 U20842 ( .B1(n17712), .B2(n18791), .A(n17738), .ZN(n17725) );
  AOI22_X1 U20843 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17725), .B1(
        n17770), .B2(n17713), .ZN(n17714) );
  NAND2_X1 U20844 ( .A1(n18071), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n18056) );
  OAI211_X1 U20845 ( .C1(n10170), .C2(n17715), .A(n17714), .B(n18056), .ZN(
        n17716) );
  AOI221_X1 U20846 ( .B1(n17718), .B2(n18053), .C1(n17717), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n17716), .ZN(n17719) );
  OAI21_X1 U20847 ( .B1(n18058), .B2(n17831), .A(n17719), .ZN(P3_U2814) );
  NOR2_X1 U20848 ( .A1(n17743), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18066) );
  NAND2_X1 U20849 ( .A1(n17902), .A2(n17720), .ZN(n17735) );
  NOR2_X1 U20850 ( .A1(n17722), .A2(n17721), .ZN(n17727) );
  INV_X1 U20851 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17726) );
  OAI22_X1 U20852 ( .A1(n18140), .A2(n18838), .B1(n17754), .B2(n17723), .ZN(
        n17724) );
  AOI221_X1 U20853 ( .B1(n17727), .B2(n17726), .C1(n17725), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17724), .ZN(n17734) );
  NAND3_X1 U20854 ( .A1(n17771), .A2(n18076), .A3(n17815), .ZN(n17736) );
  NAND4_X1 U20855 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18114), .A3(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(n17728), .ZN(n17729) );
  NAND2_X1 U20856 ( .A1(n17736), .A2(n17729), .ZN(n17730) );
  OAI221_X1 U20857 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18083), 
        .C1(n18092), .C2(n10022), .A(n17730), .ZN(n17731) );
  XOR2_X1 U20858 ( .A(n18074), .B(n17731), .Z(n18070) );
  NOR2_X1 U20859 ( .A1(n17974), .A2(n17758), .ZN(n17732) );
  OAI21_X1 U20860 ( .B1(n18049), .B2(n17782), .A(n18074), .ZN(n18061) );
  AOI22_X1 U20861 ( .A1(n17810), .A2(n18070), .B1(n17732), .B2(n18061), .ZN(
        n17733) );
  OAI211_X1 U20862 ( .C1(n18066), .C2(n17735), .A(n17734), .B(n17733), .ZN(
        P3_U2815) );
  OAI22_X1 U20863 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17736), .B1(
        n17803), .B2(n18060), .ZN(n17737) );
  XOR2_X1 U20864 ( .A(n18083), .B(n17737), .Z(n18090) );
  AOI221_X1 U20865 ( .B1(n18592), .B2(n17740), .C1(n17739), .C2(n17740), .A(
        n17738), .ZN(n17741) );
  NOR2_X1 U20866 ( .A1(n18140), .A2(n18837), .ZN(n18085) );
  AOI211_X1 U20867 ( .C1(n17742), .C2(n17696), .A(n17741), .B(n18085), .ZN(
        n17747) );
  NOR2_X1 U20868 ( .A1(n18123), .A2(n18108), .ZN(n18098) );
  INV_X1 U20869 ( .A(n18098), .ZN(n17744) );
  AOI221_X1 U20870 ( .B1(n18076), .B2(n18083), .C1(n17744), .C2(n18083), .A(
        n17743), .ZN(n18086) );
  NAND2_X1 U20871 ( .A1(n18075), .A2(n18121), .ZN(n18100) );
  NOR2_X1 U20872 ( .A1(n18049), .A2(n17782), .ZN(n17745) );
  AOI221_X1 U20873 ( .B1(n18076), .B2(n18083), .C1(n18100), .C2(n18083), .A(
        n17745), .ZN(n18087) );
  AOI22_X1 U20874 ( .A1(n17902), .A2(n18086), .B1(n17828), .B2(n18087), .ZN(
        n17746) );
  OAI211_X1 U20875 ( .C1(n18090), .C2(n17831), .A(n17747), .B(n17746), .ZN(
        P3_U2816) );
  NAND2_X1 U20876 ( .A1(n18075), .A2(n18076), .ZN(n18106) );
  NAND2_X1 U20877 ( .A1(n16695), .A2(n17748), .ZN(n17767) );
  AOI211_X1 U20878 ( .C1(n17766), .C2(n17755), .A(n17749), .B(n17767), .ZN(
        n17757) );
  OAI21_X1 U20879 ( .B1(n16695), .B2(n17750), .A(n18791), .ZN(n17751) );
  AOI21_X1 U20880 ( .B1(n17752), .B2(n17751), .A(n17818), .ZN(n17765) );
  OAI22_X1 U20881 ( .A1(n17765), .A2(n17755), .B1(n17754), .B2(n17753), .ZN(
        n17756) );
  AOI211_X1 U20882 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n18071), .A(n17757), 
        .B(n17756), .ZN(n17764) );
  INV_X1 U20883 ( .A(n18100), .ZN(n17759) );
  OAI22_X1 U20884 ( .A1(n18098), .A2(n17916), .B1(n17759), .B2(n17758), .ZN(
        n17773) );
  AOI22_X1 U20885 ( .A1(n17728), .A2(n18075), .B1(n18092), .B2(n17815), .ZN(
        n17760) );
  NOR2_X1 U20886 ( .A1(n17761), .A2(n17760), .ZN(n17762) );
  XOR2_X1 U20887 ( .A(n17762), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n18091) );
  AOI22_X1 U20888 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17773), .B1(
        n17810), .B2(n18091), .ZN(n17763) );
  OAI211_X1 U20889 ( .C1(n17813), .C2(n18106), .A(n17764), .B(n17763), .ZN(
        P3_U2817) );
  NAND2_X1 U20890 ( .A1(n18071), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18116) );
  OAI221_X1 U20891 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17767), .C1(
        n17766), .C2(n17765), .A(n18116), .ZN(n17768) );
  AOI21_X1 U20892 ( .B1(n17770), .B2(n17769), .A(n17768), .ZN(n17777) );
  AOI22_X1 U20893 ( .A1(n18114), .A2(n17795), .B1(n17771), .B2(n17815), .ZN(
        n17772) );
  XOR2_X1 U20894 ( .A(n18092), .B(n17772), .Z(n18115) );
  AOI22_X1 U20895 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17773), .B1(
        n17810), .B2(n18115), .ZN(n17776) );
  NAND3_X1 U20896 ( .A1(n18114), .A2(n18092), .A3(n17774), .ZN(n17775) );
  NAND3_X1 U20897 ( .A1(n17777), .A2(n17776), .A3(n17775), .ZN(P3_U2818) );
  NAND2_X1 U20898 ( .A1(n18126), .A2(n18093), .ZN(n18133) );
  NAND3_X1 U20899 ( .A1(n18304), .A2(n17788), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17793) );
  INV_X1 U20900 ( .A(n17909), .ZN(n17869) );
  NAND2_X1 U20901 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n17869), .ZN(
        n17778) );
  AOI22_X1 U20902 ( .A1(n18304), .A2(n16695), .B1(n17793), .B2(n17778), .ZN(
        n17780) );
  INV_X1 U20903 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18830) );
  NOR2_X1 U20904 ( .A1(n18140), .A2(n18830), .ZN(n17779) );
  AOI211_X1 U20905 ( .C1(n17781), .C2(n17696), .A(n17780), .B(n17779), .ZN(
        n17787) );
  AOI22_X1 U20906 ( .A1(n17902), .A2(n18123), .B1(n17828), .B2(n17782), .ZN(
        n17812) );
  OAI21_X1 U20907 ( .B1(n18126), .B2(n17813), .A(n17812), .ZN(n17785) );
  NAND2_X1 U20908 ( .A1(n17783), .A2(n10018), .ZN(n17804) );
  OAI22_X1 U20909 ( .A1(n18095), .A2(n17803), .B1(n17799), .B2(n17804), .ZN(
        n17784) );
  XOR2_X1 U20910 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17784), .Z(
        n18119) );
  AOI22_X1 U20911 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17785), .B1(
        n17810), .B2(n18119), .ZN(n17786) );
  OAI211_X1 U20912 ( .C1(n17813), .C2(n18133), .A(n17787), .B(n17786), .ZN(
        P3_U2819) );
  AND2_X1 U20913 ( .A1(n17788), .A2(n18304), .ZN(n17808) );
  AOI21_X1 U20914 ( .B1(n17869), .B2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n17808), .ZN(n17789) );
  INV_X1 U20915 ( .A(n17789), .ZN(n17792) );
  OAI22_X1 U20916 ( .A1(n17897), .A2(n17790), .B1(n18140), .B2(n18828), .ZN(
        n17791) );
  AOI21_X1 U20917 ( .B1(n17793), .B2(n17792), .A(n17791), .ZN(n17802) );
  NOR4_X1 U20918 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n10022), .A3(
        n18134), .A4(n17794), .ZN(n17797) );
  AOI221_X1 U20919 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n17803), 
        .C1(n18134), .C2(n17795), .A(n18146), .ZN(n17796) );
  AOI211_X1 U20920 ( .C1(n17798), .C2(n17804), .A(n17797), .B(n17796), .ZN(
        n18135) );
  NOR2_X1 U20921 ( .A1(n18126), .A2(n17813), .ZN(n17800) );
  AOI22_X1 U20922 ( .A1(n17810), .A2(n18135), .B1(n17800), .B2(n17799), .ZN(
        n17801) );
  OAI211_X1 U20923 ( .C1(n17812), .C2(n18134), .A(n17802), .B(n17801), .ZN(
        P3_U2820) );
  NAND2_X1 U20924 ( .A1(n17804), .A2(n17803), .ZN(n17805) );
  XOR2_X1 U20925 ( .A(n17805), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18150) );
  NOR2_X1 U20926 ( .A1(n18140), .A2(n18826), .ZN(n18152) );
  NOR2_X1 U20927 ( .A1(n18592), .A2(n17819), .ZN(n17832) );
  AOI22_X1 U20928 ( .A1(n17816), .A2(n17832), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17869), .ZN(n17807) );
  OAI22_X1 U20929 ( .A1(n17808), .A2(n17807), .B1(n17897), .B2(n17806), .ZN(
        n17809) );
  AOI211_X1 U20930 ( .C1(n17810), .C2(n18150), .A(n18152), .B(n17809), .ZN(
        n17811) );
  OAI221_X1 U20931 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17813), .C1(
        n18146), .C2(n17812), .A(n17811), .ZN(P3_U2821) );
  AOI21_X1 U20932 ( .B1(n17815), .B2(n17827), .A(n17814), .ZN(n18171) );
  AOI211_X1 U20933 ( .C1(n17821), .C2(n17817), .A(n17816), .B(n18592), .ZN(
        n17823) );
  AOI21_X1 U20934 ( .B1(n17820), .B2(n17819), .A(n17818), .ZN(n17835) );
  OAI22_X1 U20935 ( .A1(n18140), .A2(n18824), .B1(n17821), .B2(n17835), .ZN(
        n17822) );
  AOI211_X1 U20936 ( .C1(n17824), .C2(n17696), .A(n17823), .B(n17822), .ZN(
        n17830) );
  AOI21_X1 U20937 ( .B1(n17826), .B2(n10018), .A(n17825), .ZN(n18165) );
  INV_X1 U20938 ( .A(n17827), .ZN(n18167) );
  AOI22_X1 U20939 ( .A1(n17902), .A2(n18165), .B1(n17828), .B2(n18167), .ZN(
        n17829) );
  OAI211_X1 U20940 ( .C1(n18171), .C2(n17831), .A(n17830), .B(n17829), .ZN(
        P3_U2822) );
  INV_X1 U20941 ( .A(n17832), .ZN(n17833) );
  NAND2_X1 U20942 ( .A1(n18071), .A2(P3_REIP_REG_7__SCAN_IN), .ZN(n18179) );
  OAI221_X1 U20943 ( .B1(n17835), .B2(n17834), .C1(n17833), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18179), .ZN(n17836) );
  INV_X1 U20944 ( .A(n17836), .ZN(n17844) );
  NAND2_X1 U20945 ( .A1(n17838), .A2(n17837), .ZN(n17839) );
  XOR2_X1 U20946 ( .A(n17839), .B(n18175), .Z(n18173) );
  INV_X1 U20947 ( .A(n17840), .ZN(n17841) );
  AOI21_X1 U20948 ( .B1(n18175), .B2(n17842), .A(n17841), .ZN(n18172) );
  AOI22_X1 U20949 ( .A1(n17902), .A2(n18173), .B1(n9659), .B2(n18172), .ZN(
        n17843) );
  OAI211_X1 U20950 ( .C1(n17897), .C2(n17845), .A(n17844), .B(n17843), .ZN(
        P3_U2823) );
  AOI21_X1 U20951 ( .B1(n17847), .B2(n17846), .A(n9754), .ZN(n18182) );
  NOR2_X1 U20952 ( .A1(n18140), .A2(n18820), .ZN(n18181) );
  INV_X1 U20953 ( .A(n17853), .ZN(n17848) );
  NOR3_X1 U20954 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17848), .A3(
        n18592), .ZN(n17849) );
  AOI211_X1 U20955 ( .C1(n9659), .C2(n18182), .A(n18181), .B(n17849), .ZN(
        n17855) );
  AOI21_X1 U20956 ( .B1(n17852), .B2(n17851), .A(n17850), .ZN(n18183) );
  AOI21_X1 U20957 ( .B1(n17853), .B2(n18304), .A(n17909), .ZN(n17864) );
  AOI22_X1 U20958 ( .A1(n17902), .A2(n18183), .B1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17864), .ZN(n17854) );
  OAI211_X1 U20959 ( .C1(n17897), .C2(n17856), .A(n17855), .B(n17854), .ZN(
        P3_U2824) );
  AOI21_X1 U20960 ( .B1(n17859), .B2(n17858), .A(n17857), .ZN(n18188) );
  AOI22_X1 U20961 ( .A1(n17902), .A2(n18188), .B1(n18071), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17866) );
  AOI21_X1 U20962 ( .B1(n18189), .B2(n17861), .A(n17860), .ZN(n18187) );
  NAND3_X1 U20963 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(n17912), .ZN(n17868) );
  OAI21_X1 U20964 ( .B1(n17880), .B2(n17868), .A(n17862), .ZN(n17863) );
  AOI22_X1 U20965 ( .A1(n9659), .A2(n18187), .B1(n17864), .B2(n17863), .ZN(
        n17865) );
  OAI211_X1 U20966 ( .C1(n17897), .C2(n17867), .A(n17866), .B(n17865), .ZN(
        P3_U2825) );
  NAND2_X1 U20967 ( .A1(n17869), .A2(n17868), .ZN(n17889) );
  AOI21_X1 U20968 ( .B1(n17872), .B2(n17871), .A(n17870), .ZN(n18204) );
  NOR2_X1 U20969 ( .A1(n18140), .A2(n18816), .ZN(n18201) );
  NOR3_X1 U20970 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17873), .A3(
        n18592), .ZN(n17874) );
  AOI211_X1 U20971 ( .C1(n17902), .C2(n18204), .A(n18201), .B(n17874), .ZN(
        n17879) );
  AOI21_X1 U20972 ( .B1(n9765), .B2(n17876), .A(n17875), .ZN(n18202) );
  AOI22_X1 U20973 ( .A1(n9659), .A2(n18202), .B1(n17877), .B2(n17696), .ZN(
        n17878) );
  OAI211_X1 U20974 ( .C1(n17880), .C2(n17889), .A(n17879), .B(n17878), .ZN(
        P3_U2826) );
  AOI21_X1 U20975 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17912), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17890) );
  AOI21_X1 U20976 ( .B1(n17883), .B2(n17882), .A(n17881), .ZN(n18213) );
  AOI22_X1 U20977 ( .A1(n17902), .A2(n18213), .B1(n18071), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17888) );
  AOI21_X1 U20978 ( .B1(n18216), .B2(n17885), .A(n17884), .ZN(n18209) );
  AOI22_X1 U20979 ( .A1(n9659), .A2(n18209), .B1(n17886), .B2(n17696), .ZN(
        n17887) );
  OAI211_X1 U20980 ( .C1(n17890), .C2(n17889), .A(n17888), .B(n17887), .ZN(
        P3_U2827) );
  AOI21_X1 U20981 ( .B1(n17893), .B2(n17892), .A(n17891), .ZN(n18225) );
  NOR2_X1 U20982 ( .A1(n18140), .A2(n18812), .ZN(n18217) );
  XNOR2_X1 U20983 ( .A(n17895), .B(n17894), .ZN(n18229) );
  OAI22_X1 U20984 ( .A1(n17897), .A2(n17896), .B1(n17916), .B2(n18229), .ZN(
        n17898) );
  AOI211_X1 U20985 ( .C1(n9659), .C2(n18225), .A(n18217), .B(n17898), .ZN(
        n17899) );
  OAI221_X1 U20986 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18592), .C1(
        n17900), .C2(n17912), .A(n17899), .ZN(P3_U2828) );
  NOR2_X1 U20987 ( .A1(n17911), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17901) );
  XNOR2_X1 U20988 ( .A(n17901), .B(n17904), .ZN(n18237) );
  AOI22_X1 U20989 ( .A1(n17902), .A2(n18237), .B1(n18071), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17907) );
  AOI21_X1 U20990 ( .B1(n17904), .B2(n17910), .A(n17903), .ZN(n18231) );
  AOI22_X1 U20991 ( .A1(n9659), .A2(n18231), .B1(n17908), .B2(n17696), .ZN(
        n17906) );
  OAI211_X1 U20992 ( .C1(n17909), .C2(n17908), .A(n17907), .B(n17906), .ZN(
        P3_U2829) );
  OAI21_X1 U20993 ( .B1(n17911), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17910), .ZN(n18245) );
  INV_X1 U20994 ( .A(n18245), .ZN(n18247) );
  NAND3_X1 U20995 ( .A1(n18905), .A2(n18791), .A3(n17912), .ZN(n17913) );
  AOI22_X1 U20996 ( .A1(n18071), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17913), .ZN(n17914) );
  OAI221_X1 U20997 ( .B1(n18247), .B2(n17916), .C1(n18245), .C2(n17915), .A(
        n17914), .ZN(P3_U2830) );
  AOI221_X1 U20998 ( .B1(n17982), .B2(n17918), .C1(n17917), .C2(n17918), .A(
        n18161), .ZN(n17929) );
  OAI22_X1 U20999 ( .A1(n17920), .A2(n18097), .B1(n17919), .B2(n18120), .ZN(
        n17927) );
  NOR2_X1 U21000 ( .A1(n18717), .A2(n18738), .ZN(n18196) );
  INV_X1 U21001 ( .A(n18196), .ZN(n18221) );
  OAI21_X1 U21002 ( .B1(n18251), .B2(n17921), .A(n18738), .ZN(n17987) );
  OAI21_X1 U21003 ( .B1(n17922), .B2(n18196), .A(n17987), .ZN(n17957) );
  AOI21_X1 U21004 ( .B1(n17923), .B2(n18221), .A(n17957), .ZN(n17945) );
  NAND2_X1 U21005 ( .A1(n18128), .A2(n18721), .ZN(n18232) );
  OAI21_X1 U21006 ( .B1(n17940), .B2(n17924), .A(n18232), .ZN(n17925) );
  OAI211_X1 U21007 ( .C1(n18740), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17945), .B(n17925), .ZN(n17926) );
  NOR2_X1 U21008 ( .A1(n17927), .A2(n17926), .ZN(n17933) );
  OAI211_X1 U21009 ( .C1(n18740), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17933), .ZN(n17928) );
  AOI22_X1 U21010 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18242), .B1(
        n17929), .B2(n17928), .ZN(n17931) );
  OAI211_X1 U21011 ( .C1(n17932), .C2(n18170), .A(n17931), .B(n17930), .ZN(
        P3_U2835) );
  OAI22_X1 U21012 ( .A1(n17982), .A2(n17934), .B1(n17933), .B2(n10019), .ZN(
        n17935) );
  AOI22_X1 U21013 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18242), .B1(
        n18243), .B2(n17935), .ZN(n17937) );
  NAND2_X1 U21014 ( .A1(n18071), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17936) );
  OAI211_X1 U21015 ( .C1(n17938), .C2(n18170), .A(n17937), .B(n17936), .ZN(
        P3_U2836) );
  NOR2_X1 U21016 ( .A1(n17940), .A2(n17939), .ZN(n17944) );
  AOI21_X1 U21017 ( .B1(n17942), .B2(n17941), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17943) );
  AOI211_X1 U21018 ( .C1(n17945), .C2(n17944), .A(n17943), .B(n18161), .ZN(
        n17946) );
  AOI21_X1 U21019 ( .B1(n18242), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17946), .ZN(n17948) );
  OAI211_X1 U21020 ( .C1(n17949), .C2(n18170), .A(n17948), .B(n17947), .ZN(
        n17950) );
  AOI21_X1 U21021 ( .B1(n18166), .B2(n17951), .A(n17950), .ZN(n17952) );
  OAI21_X1 U21022 ( .B1(n18230), .B2(n17953), .A(n17952), .ZN(P3_U2837) );
  OAI22_X1 U21023 ( .A1(n17955), .A2(n18097), .B1(n17954), .B2(n18120), .ZN(
        n17956) );
  NOR3_X1 U21024 ( .A1(n18242), .A2(n17957), .A3(n17956), .ZN(n17961) );
  OAI211_X1 U21025 ( .C1(n17958), .C2(n18721), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n17961), .ZN(n17959) );
  AND2_X1 U21026 ( .A1(n18140), .A2(n17959), .ZN(n17969) );
  AOI21_X1 U21027 ( .B1(n18052), .B2(n17961), .A(n17960), .ZN(n17962) );
  AOI22_X1 U21028 ( .A1(n17994), .A2(n17963), .B1(n17969), .B2(n17962), .ZN(
        n17965) );
  NAND2_X1 U21029 ( .A1(n18071), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17964) );
  OAI211_X1 U21030 ( .C1(n17966), .C2(n18170), .A(n17965), .B(n17964), .ZN(
        P3_U2838) );
  INV_X1 U21031 ( .A(n17967), .ZN(n17973) );
  NOR3_X1 U21032 ( .A1(n18242), .A2(n17982), .A3(n17968), .ZN(n17970) );
  OAI21_X1 U21033 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17970), .A(
        n17969), .ZN(n17971) );
  OAI211_X1 U21034 ( .C1(n17973), .C2(n18170), .A(n17972), .B(n17971), .ZN(
        P3_U2839) );
  OAI22_X1 U21035 ( .A1(n18067), .A2(n18097), .B1(n17974), .B2(n18120), .ZN(
        n17995) );
  NOR2_X1 U21036 ( .A1(n18750), .A2(n18101), .ZN(n18125) );
  AOI21_X1 U21037 ( .B1(n18028), .B2(n17975), .A(n18721), .ZN(n18025) );
  AOI21_X1 U21038 ( .B1(n18024), .B2(n18008), .A(n18740), .ZN(n17976) );
  AOI211_X1 U21039 ( .C1(n18751), .C2(n17977), .A(n18025), .B(n17976), .ZN(
        n18007) );
  NAND2_X1 U21040 ( .A1(n18717), .A2(n17978), .ZN(n17979) );
  OAI211_X1 U21041 ( .C1(n17984), .C2(n18125), .A(n18007), .B(n17979), .ZN(
        n17998) );
  OAI22_X1 U21042 ( .A1(n18138), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n17980), .B2(n18721), .ZN(n17981) );
  NOR4_X1 U21043 ( .A1(n17992), .A2(n17995), .A3(n17998), .A4(n17981), .ZN(
        n17986) );
  INV_X1 U21044 ( .A(n17982), .ZN(n17983) );
  AOI21_X1 U21045 ( .B1(n17984), .B2(n17983), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17985) );
  AOI211_X1 U21046 ( .C1(n17987), .C2(n17986), .A(n17985), .B(n18161), .ZN(
        n17988) );
  AOI21_X1 U21047 ( .B1(n17989), .B2(n18151), .A(n17988), .ZN(n17991) );
  NAND2_X1 U21048 ( .A1(n18071), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17990) );
  OAI211_X1 U21049 ( .C1(n18233), .C2(n17992), .A(n17991), .B(n17990), .ZN(
        P3_U2840) );
  NAND2_X1 U21050 ( .A1(n17994), .A2(n17993), .ZN(n18022) );
  NOR2_X1 U21051 ( .A1(n18161), .A2(n17995), .ZN(n18051) );
  OAI21_X1 U21052 ( .B1(n18045), .B2(n17996), .A(n18738), .ZN(n17997) );
  NAND2_X1 U21053 ( .A1(n18051), .A2(n17997), .ZN(n18010) );
  AOI211_X1 U21054 ( .C1(n17999), .C2(n18232), .A(n17998), .B(n18010), .ZN(
        n18001) );
  NOR3_X1 U21055 ( .A1(n18071), .A2(n18001), .A3(n18000), .ZN(n18002) );
  AOI21_X1 U21056 ( .B1(n18151), .B2(n18003), .A(n18002), .ZN(n18005) );
  OAI211_X1 U21057 ( .C1(n18006), .C2(n18022), .A(n18005), .B(n18004), .ZN(
        P3_U2841) );
  NAND3_X1 U21058 ( .A1(n18021), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(n18232), 
        .ZN(n18011) );
  OAI21_X1 U21059 ( .B1(n18008), .B2(n18125), .A(n18007), .ZN(n18009) );
  OAI21_X1 U21060 ( .B1(n18010), .B2(n18009), .A(n18140), .ZN(n18020) );
  NAND2_X1 U21061 ( .A1(n18011), .A2(n18020), .ZN(n18013) );
  AOI22_X1 U21062 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18013), .B1(
        n18151), .B2(n18012), .ZN(n18015) );
  OAI211_X1 U21063 ( .C1(n18022), .C2(n18016), .A(n18015), .B(n18014), .ZN(
        P3_U2842) );
  AOI21_X1 U21064 ( .B1(n18151), .B2(n18018), .A(n18017), .ZN(n18019) );
  OAI221_X1 U21065 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18022), 
        .C1(n18021), .C2(n18020), .A(n18019), .ZN(P3_U2843) );
  NOR2_X1 U21066 ( .A1(n18128), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18219) );
  INV_X1 U21067 ( .A(n18219), .ZN(n18023) );
  NAND3_X1 U21068 ( .A1(n18024), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18023), .ZN(n18026) );
  AOI21_X1 U21069 ( .B1(n18221), .B2(n18026), .A(n18025), .ZN(n18027) );
  OAI211_X1 U21070 ( .C1(n18028), .C2(n18125), .A(n18051), .B(n18027), .ZN(
        n18040) );
  OAI221_X1 U21071 ( .B1(n18040), .B2(n18029), .C1(n18040), .C2(n18221), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18039) );
  INV_X1 U21072 ( .A(n18030), .ZN(n18034) );
  AOI22_X1 U21073 ( .A1(n18751), .A2(n18031), .B1(n18197), .B2(n18218), .ZN(
        n18210) );
  NOR2_X1 U21074 ( .A1(n18210), .A2(n18032), .ZN(n18177) );
  NAND2_X1 U21075 ( .A1(n18033), .A2(n18177), .ZN(n18059) );
  NAND2_X1 U21076 ( .A1(n18034), .A2(n18059), .ZN(n18113) );
  NAND2_X1 U21077 ( .A1(n18243), .A2(n18113), .ZN(n18155) );
  NOR2_X1 U21078 ( .A1(n18035), .A2(n18155), .ZN(n18054) );
  AOI22_X1 U21079 ( .A1(n18151), .A2(n18037), .B1(n18054), .B2(n18036), .ZN(
        n18038) );
  OAI221_X1 U21080 ( .B1(n18071), .B2(n18039), .C1(n18140), .C2(n18844), .A(
        n18038), .ZN(P3_U2844) );
  NAND2_X1 U21081 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18040), .ZN(
        n18044) );
  AOI22_X1 U21082 ( .A1(n18151), .A2(n18042), .B1(n18054), .B2(n18041), .ZN(
        n18043) );
  OAI221_X1 U21083 ( .B1(n18071), .B2(n18044), .C1(n18140), .C2(n18843), .A(
        n18043), .ZN(P3_U2845) );
  INV_X1 U21084 ( .A(n18045), .ZN(n18046) );
  AOI21_X1 U21085 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18128), .A(
        n18046), .ZN(n18048) );
  NAND2_X1 U21086 ( .A1(n18751), .A2(n18047), .ZN(n18124) );
  NAND2_X1 U21087 ( .A1(n18717), .A2(n18094), .ZN(n18136) );
  NAND2_X1 U21088 ( .A1(n18124), .A2(n18136), .ZN(n18145) );
  AOI211_X1 U21089 ( .C1(n18050), .C2(n18049), .A(n18048), .B(n18145), .ZN(
        n18063) );
  AOI221_X1 U21090 ( .B1(n18052), .B2(n18051), .C1(n18063), .C2(n18051), .A(
        n18071), .ZN(n18055) );
  AOI22_X1 U21091 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18055), .B1(
        n18054), .B2(n18053), .ZN(n18057) );
  OAI211_X1 U21092 ( .C1(n18058), .C2(n18170), .A(n18057), .B(n18056), .ZN(
        P3_U2846) );
  NOR2_X1 U21093 ( .A1(n18060), .A2(n18059), .ZN(n18080) );
  AOI21_X1 U21094 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18080), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18065) );
  NAND3_X1 U21095 ( .A1(n18101), .A2(n18062), .A3(n18061), .ZN(n18064) );
  AOI221_X1 U21096 ( .B1(n18065), .B2(n18064), .C1(n18063), .C2(n18064), .A(
        n18161), .ZN(n18069) );
  NOR3_X1 U21097 ( .A1(n18067), .A2(n18066), .A3(n18230), .ZN(n18068) );
  AOI211_X1 U21098 ( .C1(n18070), .C2(n18151), .A(n18069), .B(n18068), .ZN(
        n18073) );
  NAND2_X1 U21099 ( .A1(n18071), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18072) );
  OAI211_X1 U21100 ( .C1(n18233), .C2(n18074), .A(n18073), .B(n18072), .ZN(
        P3_U2847) );
  AOI21_X1 U21101 ( .B1(n18075), .B2(n18107), .A(n18128), .ZN(n18103) );
  AOI211_X1 U21102 ( .C1(n18076), .C2(n18232), .A(n18103), .B(n18145), .ZN(
        n18077) );
  OAI211_X1 U21103 ( .C1(n18138), .C2(n18078), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18077), .ZN(n18079) );
  NAND2_X1 U21104 ( .A1(n18243), .A2(n18079), .ZN(n18082) );
  INV_X1 U21105 ( .A(n18080), .ZN(n18081) );
  AOI222_X1 U21106 ( .A1(n18083), .A2(n18082), .B1(n18083), .B2(n18081), .C1(
        n18082), .C2(n18233), .ZN(n18084) );
  AOI211_X1 U21107 ( .C1(n18086), .C2(n18246), .A(n18085), .B(n18084), .ZN(
        n18089) );
  NAND2_X1 U21108 ( .A1(n18166), .A2(n18087), .ZN(n18088) );
  OAI211_X1 U21109 ( .C1(n18090), .C2(n18170), .A(n18089), .B(n18088), .ZN(
        P3_U2848) );
  AOI22_X1 U21110 ( .A1(n18071), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18151), 
        .B2(n18091), .ZN(n18105) );
  AOI21_X1 U21111 ( .B1(n18717), .B2(n18093), .A(n18092), .ZN(n18110) );
  OAI21_X1 U21112 ( .B1(n18095), .B2(n18094), .A(n18717), .ZN(n18096) );
  OAI21_X1 U21113 ( .B1(n18114), .B2(n18721), .A(n18096), .ZN(n18130) );
  OAI21_X1 U21114 ( .B1(n18098), .B2(n18097), .A(n18124), .ZN(n18099) );
  AOI211_X1 U21115 ( .C1(n18101), .C2(n18100), .A(n18130), .B(n18099), .ZN(
        n18109) );
  OAI211_X1 U21116 ( .C1(n18138), .C2(n18110), .A(n18243), .B(n18109), .ZN(
        n18102) );
  OAI211_X1 U21117 ( .C1(n18103), .C2(n18102), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18140), .ZN(n18104) );
  OAI211_X1 U21118 ( .C1(n18106), .C2(n18155), .A(n18105), .B(n18104), .ZN(
        P3_U2849) );
  INV_X1 U21119 ( .A(n18107), .ZN(n18144) );
  NOR2_X1 U21120 ( .A1(n18108), .A2(n18144), .ZN(n18111) );
  OAI211_X1 U21121 ( .C1(n18111), .C2(n18128), .A(n18110), .B(n18109), .ZN(
        n18112) );
  OAI221_X1 U21122 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18114), 
        .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18113), .A(n18112), .ZN(
        n18118) );
  AOI22_X1 U21123 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18242), .B1(
        n18151), .B2(n18115), .ZN(n18117) );
  OAI211_X1 U21124 ( .C1(n18161), .C2(n18118), .A(n18117), .B(n18116), .ZN(
        P3_U2850) );
  AOI22_X1 U21125 ( .A1(n18071), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18151), 
        .B2(n18119), .ZN(n18132) );
  OAI21_X1 U21126 ( .B1(n18121), .B2(n18120), .A(n18243), .ZN(n18122) );
  AOI21_X1 U21127 ( .B1(n18750), .B2(n18123), .A(n18122), .ZN(n18148) );
  OAI211_X1 U21128 ( .C1(n18126), .C2(n18125), .A(n18148), .B(n18124), .ZN(
        n18127) );
  AOI221_X1 U21129 ( .B1(n18146), .B2(n18738), .C1(n18144), .C2(n18738), .A(
        n18127), .ZN(n18137) );
  OAI21_X1 U21130 ( .B1(n18128), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18137), .ZN(n18129) );
  OAI211_X1 U21131 ( .C1(n18130), .C2(n18129), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18140), .ZN(n18131) );
  OAI211_X1 U21132 ( .C1(n18133), .C2(n18155), .A(n18132), .B(n18131), .ZN(
        P3_U2851) );
  NAND2_X1 U21133 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18134), .ZN(
        n18143) );
  AOI22_X1 U21134 ( .A1(n18071), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18151), 
        .B2(n18135), .ZN(n18142) );
  OAI211_X1 U21135 ( .C1(n18138), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18137), .B(n18136), .ZN(n18139) );
  NAND3_X1 U21136 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18140), .A3(
        n18139), .ZN(n18141) );
  OAI211_X1 U21137 ( .C1(n18143), .C2(n18155), .A(n18142), .B(n18141), .ZN(
        P3_U2852) );
  OAI21_X1 U21138 ( .B1(n18738), .B2(n18145), .A(n18144), .ZN(n18147) );
  AOI211_X1 U21139 ( .C1(n18148), .C2(n18147), .A(n18071), .B(n18146), .ZN(
        n18149) );
  AOI21_X1 U21140 ( .B1(n18151), .B2(n18150), .A(n18149), .ZN(n18154) );
  INV_X1 U21141 ( .A(n18152), .ZN(n18153) );
  OAI211_X1 U21142 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18155), .A(
        n18154), .B(n18153), .ZN(P3_U2853) );
  OAI22_X1 U21143 ( .A1(n18157), .A2(n18196), .B1(n18156), .B2(n18721), .ZN(
        n18158) );
  OAI21_X1 U21144 ( .B1(n18158), .B2(n18219), .A(n18243), .ZN(n18159) );
  INV_X1 U21145 ( .A(n18159), .ZN(n18190) );
  AOI21_X1 U21146 ( .B1(n18160), .B2(n18162), .A(n18190), .ZN(n18174) );
  AOI21_X1 U21147 ( .B1(n18174), .B2(n18233), .A(n10018), .ZN(n18164) );
  NOR3_X1 U21148 ( .A1(n18210), .A2(n18161), .A3(n18216), .ZN(n18203) );
  NAND3_X1 U21149 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n18203), .ZN(n18186) );
  NOR3_X1 U21150 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18162), .A3(
        n18186), .ZN(n18163) );
  AOI211_X1 U21151 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n18071), .A(n18164), .B(
        n18163), .ZN(n18169) );
  AOI22_X1 U21152 ( .A1(n18167), .A2(n18166), .B1(n18246), .B2(n18165), .ZN(
        n18168) );
  OAI211_X1 U21153 ( .C1(n18171), .C2(n18170), .A(n18169), .B(n18168), .ZN(
        P3_U2854) );
  AOI22_X1 U21154 ( .A1(n18246), .A2(n18173), .B1(n18248), .B2(n18172), .ZN(
        n18180) );
  OAI21_X1 U21155 ( .B1(n18175), .B2(n18233), .A(n18174), .ZN(n18176) );
  OAI221_X1 U21156 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18177), .A(n18176), .ZN(
        n18178) );
  NAND3_X1 U21157 ( .A1(n18180), .A2(n18179), .A3(n18178), .ZN(P3_U2855) );
  AOI221_X1 U21158 ( .B1(n18242), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        n18190), .C2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n18181), .ZN(
        n18185) );
  AOI22_X1 U21159 ( .A1(n18246), .A2(n18183), .B1(n18248), .B2(n18182), .ZN(
        n18184) );
  OAI211_X1 U21160 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n18186), .A(
        n18185), .B(n18184), .ZN(P3_U2856) );
  AOI22_X1 U21161 ( .A1(n18246), .A2(n18188), .B1(n18248), .B2(n18187), .ZN(
        n18194) );
  NAND2_X1 U21162 ( .A1(n18071), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18193) );
  NAND3_X1 U21163 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18203), .A3(
        n18189), .ZN(n18192) );
  OAI21_X1 U21164 ( .B1(n18242), .B2(n18190), .A(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18191) );
  NAND4_X1 U21165 ( .A1(n18194), .A2(n18193), .A3(n18192), .A4(n18191), .ZN(
        P3_U2857) );
  NAND2_X1 U21166 ( .A1(n18751), .A2(n18195), .ZN(n18222) );
  OAI211_X1 U21167 ( .C1(n18197), .C2(n18196), .A(n18222), .B(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18198) );
  OAI21_X1 U21168 ( .B1(n18198), .B2(n18219), .A(n18243), .ZN(n18199) );
  INV_X1 U21169 ( .A(n18199), .ZN(n18212) );
  AOI21_X1 U21170 ( .B1(n18212), .B2(n18200), .A(n18242), .ZN(n18208) );
  AOI21_X1 U21171 ( .B1(n18202), .B2(n18248), .A(n18201), .ZN(n18206) );
  AOI22_X1 U21172 ( .A1(n18204), .A2(n18246), .B1(n18203), .B2(n18207), .ZN(
        n18205) );
  OAI211_X1 U21173 ( .C1(n18208), .C2(n18207), .A(n18206), .B(n18205), .ZN(
        P3_U2858) );
  AOI22_X1 U21174 ( .A1(n18071), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18248), 
        .B2(n18209), .ZN(n18215) );
  NAND2_X1 U21175 ( .A1(n18210), .A2(n18216), .ZN(n18211) );
  AOI22_X1 U21176 ( .A1(n18246), .A2(n18213), .B1(n18212), .B2(n18211), .ZN(
        n18214) );
  OAI211_X1 U21177 ( .C1(n18216), .C2(n18233), .A(n18215), .B(n18214), .ZN(
        P3_U2859) );
  AOI21_X1 U21178 ( .B1(n18242), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n18217), .ZN(n18228) );
  NAND2_X1 U21179 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18218), .ZN(
        n18224) );
  NOR3_X1 U21180 ( .A1(n18721), .A2(n18251), .A3(n18890), .ZN(n18220) );
  AOI211_X1 U21181 ( .C1(n18890), .C2(n18221), .A(n18220), .B(n18219), .ZN(
        n18223) );
  OAI221_X1 U21182 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n18224), .C1(
        n12642), .C2(n18223), .A(n18222), .ZN(n18226) );
  AOI22_X1 U21183 ( .A1(n18243), .A2(n18226), .B1(n18248), .B2(n18225), .ZN(
        n18227) );
  OAI211_X1 U21184 ( .C1(n18230), .C2(n18229), .A(n18228), .B(n18227), .ZN(
        P3_U2860) );
  INV_X1 U21185 ( .A(n18231), .ZN(n18241) );
  NAND3_X1 U21186 ( .A1(n18243), .A2(n18251), .A3(n18232), .ZN(n18249) );
  AOI21_X1 U21187 ( .B1(n18233), .B2(n18249), .A(n18890), .ZN(n18236) );
  AOI211_X1 U21188 ( .C1(n18740), .C2(n18251), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18234), .ZN(n18235) );
  AOI211_X1 U21189 ( .C1(n18246), .C2(n18237), .A(n18236), .B(n18235), .ZN(
        n18239) );
  NAND2_X1 U21190 ( .A1(n18071), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18238) );
  OAI211_X1 U21191 ( .C1(n18241), .C2(n18240), .A(n18239), .B(n18238), .ZN(
        P3_U2861) );
  AOI21_X1 U21192 ( .B1(n18243), .B2(n18717), .A(n18242), .ZN(n18252) );
  AND2_X1 U21193 ( .A1(n18071), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18244) );
  AOI221_X1 U21194 ( .B1(n18248), .B2(n18247), .C1(n18246), .C2(n18245), .A(
        n18244), .ZN(n18250) );
  OAI211_X1 U21195 ( .C1(n18252), .C2(n18251), .A(n18250), .B(n18249), .ZN(
        P3_U2862) );
  AOI211_X1 U21196 ( .C1(n18255), .C2(n18254), .A(n18253), .B(n18905), .ZN(
        n18778) );
  OAI21_X1 U21197 ( .B1(n18778), .B2(n18256), .A(n18261), .ZN(n18257) );
  OAI221_X1 U21198 ( .B1(n18539), .B2(n18926), .C1(n18539), .C2(n18261), .A(
        n18257), .ZN(P3_U2863) );
  INV_X1 U21199 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18762) );
  NAND2_X1 U21200 ( .A1(n18761), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18482) );
  INV_X1 U21201 ( .A(n18482), .ZN(n18563) );
  NAND2_X1 U21202 ( .A1(n18762), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18411) );
  INV_X1 U21203 ( .A(n18411), .ZN(n18435) );
  NOR2_X1 U21204 ( .A1(n18563), .A2(n18435), .ZN(n18258) );
  OAI22_X1 U21205 ( .A1(n18260), .A2(n18762), .B1(n18259), .B2(n18258), .ZN(
        P3_U2866) );
  NOR2_X1 U21206 ( .A1(n18763), .A2(n18261), .ZN(P3_U2867) );
  INV_X1 U21207 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18262) );
  NOR2_X1 U21208 ( .A1(n18592), .A2(n18262), .ZN(n18594) );
  INV_X1 U21209 ( .A(n18594), .ZN(n18661) );
  NAND2_X1 U21210 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18263) );
  NAND2_X1 U21211 ( .A1(n18539), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18410) );
  NOR2_X2 U21212 ( .A1(n18263), .A2(n18410), .ZN(n18642) );
  INV_X1 U21213 ( .A(n18642), .ZN(n18651) );
  INV_X1 U21214 ( .A(n18263), .ZN(n18657) );
  NAND2_X1 U21215 ( .A1(n18657), .A2(n18743), .ZN(n18593) );
  NOR2_X2 U21216 ( .A1(n18539), .A2(n18593), .ZN(n18704) );
  AND2_X1 U21217 ( .A1(n18568), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18654) );
  NAND3_X1 U21218 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n18434), .ZN(n18711) );
  NAND2_X1 U21219 ( .A1(n18743), .A2(n18539), .ZN(n18744) );
  NAND2_X1 U21220 ( .A1(n18761), .A2(n18762), .ZN(n18343) );
  NOR2_X2 U21221 ( .A1(n18744), .A2(n18343), .ZN(n18363) );
  INV_X1 U21222 ( .A(n18363), .ZN(n18361) );
  AOI21_X1 U21223 ( .B1(n18711), .B2(n18361), .A(n18653), .ZN(n18297) );
  AOI22_X1 U21224 ( .A1(n18704), .A2(n18655), .B1(n18654), .B2(n18297), .ZN(
        n18269) );
  INV_X1 U21225 ( .A(n18410), .ZN(n18506) );
  NOR2_X1 U21226 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18539), .ZN(
        n18480) );
  NOR2_X1 U21227 ( .A1(n18506), .A2(n18480), .ZN(n18566) );
  NOR2_X1 U21228 ( .A1(n18566), .A2(n18263), .ZN(n18627) );
  NAND2_X1 U21229 ( .A1(n18568), .A2(n18264), .ZN(n18507) );
  AOI21_X1 U21230 ( .B1(n18711), .B2(n18361), .A(n18507), .ZN(n18324) );
  AOI21_X1 U21231 ( .B1(n18304), .B2(n18627), .A(n18324), .ZN(n18299) );
  NOR2_X1 U21232 ( .A1(n18266), .A2(n18265), .ZN(n18295) );
  NAND2_X1 U21233 ( .A1(n18267), .A2(n18295), .ZN(n18542) );
  INV_X1 U21234 ( .A(n18542), .ZN(n18658) );
  AOI22_X1 U21235 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18299), .B1(
        n18363), .B2(n18658), .ZN(n18268) );
  OAI211_X1 U21236 ( .C1(n18661), .C2(n18651), .A(n18269), .B(n18268), .ZN(
        P3_U2868) );
  NOR2_X1 U21237 ( .A1(n18592), .A2(n13902), .ZN(n18663) );
  INV_X1 U21238 ( .A(n18663), .ZN(n18573) );
  NAND2_X1 U21239 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18304), .ZN(n18667) );
  INV_X1 U21240 ( .A(n18667), .ZN(n18598) );
  AND2_X1 U21241 ( .A1(n18568), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18662) );
  AOI22_X1 U21242 ( .A1(n18704), .A2(n18598), .B1(n18297), .B2(n18662), .ZN(
        n18271) );
  INV_X1 U21243 ( .A(n18295), .ZN(n18290) );
  NOR2_X2 U21244 ( .A1(n18932), .A2(n18290), .ZN(n18664) );
  AOI22_X1 U21245 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18299), .B1(
        n18363), .B2(n18664), .ZN(n18270) );
  OAI211_X1 U21246 ( .C1(n18651), .C2(n18573), .A(n18271), .B(n18270), .ZN(
        P3_U2869) );
  NAND2_X1 U21247 ( .A1(n18304), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18464) );
  NAND2_X1 U21248 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18304), .ZN(n18673) );
  INV_X1 U21249 ( .A(n18673), .ZN(n18602) );
  NOR2_X2 U21250 ( .A1(n18345), .A2(n18272), .ZN(n18668) );
  AOI22_X1 U21251 ( .A1(n18704), .A2(n18602), .B1(n18297), .B2(n18668), .ZN(
        n18275) );
  NOR2_X2 U21252 ( .A1(n18273), .A2(n18290), .ZN(n18670) );
  AOI22_X1 U21253 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18299), .B1(
        n18363), .B2(n18670), .ZN(n18274) );
  OAI211_X1 U21254 ( .C1(n18651), .C2(n18464), .A(n18275), .B(n18274), .ZN(
        P3_U2870) );
  NOR2_X1 U21255 ( .A1(n18592), .A2(n13996), .ZN(n18675) );
  INV_X1 U21256 ( .A(n18675), .ZN(n18610) );
  NAND2_X1 U21257 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18304), .ZN(n18679) );
  INV_X1 U21258 ( .A(n18679), .ZN(n18606) );
  NOR2_X2 U21259 ( .A1(n18345), .A2(n18276), .ZN(n18674) );
  AOI22_X1 U21260 ( .A1(n18704), .A2(n18606), .B1(n18297), .B2(n18674), .ZN(
        n18279) );
  NOR2_X2 U21261 ( .A1(n18277), .A2(n18290), .ZN(n18676) );
  AOI22_X1 U21262 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18299), .B1(
        n18363), .B2(n18676), .ZN(n18278) );
  OAI211_X1 U21263 ( .C1(n18651), .C2(n18610), .A(n18279), .B(n18278), .ZN(
        P3_U2871) );
  NAND2_X1 U21264 ( .A1(n18304), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18685) );
  NAND2_X1 U21265 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18304), .ZN(n18552) );
  INV_X1 U21266 ( .A(n18552), .ZN(n18681) );
  NOR2_X2 U21267 ( .A1(n18345), .A2(n18280), .ZN(n18680) );
  AOI22_X1 U21268 ( .A1(n18704), .A2(n18681), .B1(n18297), .B2(n18680), .ZN(
        n18283) );
  NOR2_X2 U21269 ( .A1(n18281), .A2(n18290), .ZN(n18682) );
  AOI22_X1 U21270 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18299), .B1(
        n18363), .B2(n18682), .ZN(n18282) );
  OAI211_X1 U21271 ( .C1(n18651), .C2(n18685), .A(n18283), .B(n18282), .ZN(
        P3_U2872) );
  INV_X1 U21272 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18284) );
  NOR2_X1 U21273 ( .A1(n18592), .A2(n18284), .ZN(n18688) );
  INV_X1 U21274 ( .A(n18688), .ZN(n18471) );
  NAND2_X1 U21275 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18304), .ZN(n18692) );
  INV_X1 U21276 ( .A(n18692), .ZN(n18526) );
  NOR2_X2 U21277 ( .A1(n18345), .A2(n18285), .ZN(n18687) );
  AOI22_X1 U21278 ( .A1(n18704), .A2(n18526), .B1(n18297), .B2(n18687), .ZN(
        n18288) );
  NOR2_X2 U21279 ( .A1(n18286), .A2(n18290), .ZN(n18689) );
  AOI22_X1 U21280 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18299), .B1(
        n18363), .B2(n18689), .ZN(n18287) );
  OAI211_X1 U21281 ( .C1(n18651), .C2(n18471), .A(n18288), .B(n18287), .ZN(
        P3_U2873) );
  NOR2_X1 U21282 ( .A1(n18592), .A2(n19282), .ZN(n18694) );
  INV_X1 U21283 ( .A(n18694), .ZN(n18645) );
  NAND2_X1 U21284 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18304), .ZN(n18700) );
  INV_X1 U21285 ( .A(n18700), .ZN(n18641) );
  NOR2_X2 U21286 ( .A1(n18345), .A2(n18289), .ZN(n18693) );
  AOI22_X1 U21287 ( .A1(n18704), .A2(n18641), .B1(n18297), .B2(n18693), .ZN(
        n18293) );
  NOR2_X2 U21288 ( .A1(n9649), .A2(n18290), .ZN(n18695) );
  AOI22_X1 U21289 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18299), .B1(
        n18363), .B2(n18695), .ZN(n18292) );
  OAI211_X1 U21290 ( .C1(n18651), .C2(n18645), .A(n18293), .B(n18292), .ZN(
        P3_U2874) );
  NAND2_X1 U21291 ( .A1(n18295), .A2(n18294), .ZN(n18710) );
  AND2_X1 U21292 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18304), .ZN(n18703) );
  NOR2_X2 U21293 ( .A1(n18296), .A2(n18345), .ZN(n18702) );
  AOI22_X1 U21294 ( .A1(n18642), .A2(n18703), .B1(n18297), .B2(n18702), .ZN(
        n18301) );
  NOR2_X2 U21295 ( .A1(n18592), .A2(n18298), .ZN(n18706) );
  AOI22_X1 U21296 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18299), .B1(
        n18704), .B2(n18706), .ZN(n18300) );
  OAI211_X1 U21297 ( .C1(n18361), .C2(n18710), .A(n18301), .B(n18300), .ZN(
        P3_U2875) );
  INV_X1 U21298 ( .A(n18653), .ZN(n18623) );
  NAND2_X1 U21299 ( .A1(n18743), .A2(n18623), .ZN(n18481) );
  NOR2_X1 U21300 ( .A1(n18343), .A2(n18481), .ZN(n18319) );
  AOI22_X1 U21301 ( .A1(n18642), .A2(n18655), .B1(n18654), .B2(n18319), .ZN(
        n18306) );
  NAND2_X1 U21302 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18434), .ZN(
        n18652) );
  INV_X1 U21303 ( .A(n18652), .ZN(n18303) );
  INV_X1 U21304 ( .A(n18343), .ZN(n18346) );
  NAND2_X1 U21305 ( .A1(n18568), .A2(n18302), .ZN(n18590) );
  NOR2_X1 U21306 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18590), .ZN(
        n18484) );
  AOI22_X1 U21307 ( .A1(n18304), .A2(n18303), .B1(n18346), .B2(n18484), .ZN(
        n18320) );
  NAND2_X1 U21308 ( .A1(n18346), .A2(n18480), .ZN(n18381) );
  INV_X1 U21309 ( .A(n18381), .ZN(n18385) );
  AOI22_X1 U21310 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18320), .B1(
        n18658), .B2(n18385), .ZN(n18305) );
  OAI211_X1 U21311 ( .C1(n18711), .C2(n18661), .A(n18306), .B(n18305), .ZN(
        P3_U2876) );
  AOI22_X1 U21312 ( .A1(n18642), .A2(n18598), .B1(n18662), .B2(n18319), .ZN(
        n18308) );
  AOI22_X1 U21313 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18320), .B1(
        n18664), .B2(n18385), .ZN(n18307) );
  OAI211_X1 U21314 ( .C1(n18711), .C2(n18573), .A(n18308), .B(n18307), .ZN(
        P3_U2877) );
  AOI22_X1 U21315 ( .A1(n18642), .A2(n18602), .B1(n18668), .B2(n18319), .ZN(
        n18310) );
  AOI22_X1 U21316 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18320), .B1(
        n18670), .B2(n18385), .ZN(n18309) );
  OAI211_X1 U21317 ( .C1(n18711), .C2(n18464), .A(n18310), .B(n18309), .ZN(
        P3_U2878) );
  AOI22_X1 U21318 ( .A1(n18642), .A2(n18606), .B1(n18674), .B2(n18319), .ZN(
        n18312) );
  AOI22_X1 U21319 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18320), .B1(
        n18676), .B2(n18385), .ZN(n18311) );
  OAI211_X1 U21320 ( .C1(n18711), .C2(n18610), .A(n18312), .B(n18311), .ZN(
        P3_U2879) );
  AOI22_X1 U21321 ( .A1(n18642), .A2(n18681), .B1(n18680), .B2(n18319), .ZN(
        n18314) );
  AOI22_X1 U21322 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18320), .B1(
        n18682), .B2(n18385), .ZN(n18313) );
  OAI211_X1 U21323 ( .C1(n18711), .C2(n18685), .A(n18314), .B(n18313), .ZN(
        P3_U2880) );
  INV_X1 U21324 ( .A(n18711), .ZN(n18696) );
  AOI22_X1 U21325 ( .A1(n18696), .A2(n18688), .B1(n18687), .B2(n18319), .ZN(
        n18316) );
  AOI22_X1 U21326 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18320), .B1(
        n18689), .B2(n18385), .ZN(n18315) );
  OAI211_X1 U21327 ( .C1(n18651), .C2(n18692), .A(n18316), .B(n18315), .ZN(
        P3_U2881) );
  AOI22_X1 U21328 ( .A1(n18642), .A2(n18641), .B1(n18693), .B2(n18319), .ZN(
        n18318) );
  AOI22_X1 U21329 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18320), .B1(
        n18695), .B2(n18385), .ZN(n18317) );
  OAI211_X1 U21330 ( .C1(n18711), .C2(n18645), .A(n18318), .B(n18317), .ZN(
        P3_U2882) );
  AOI22_X1 U21331 ( .A1(n18696), .A2(n18703), .B1(n18702), .B2(n18319), .ZN(
        n18322) );
  AOI22_X1 U21332 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18320), .B1(
        n18642), .B2(n18706), .ZN(n18321) );
  OAI211_X1 U21333 ( .C1(n18710), .C2(n18381), .A(n18322), .B(n18321), .ZN(
        P3_U2883) );
  NOR2_X2 U21334 ( .A1(n18343), .A2(n18410), .ZN(n18406) );
  INV_X1 U21335 ( .A(n18406), .ZN(n18404) );
  NAND2_X1 U21336 ( .A1(n18381), .A2(n18404), .ZN(n18323) );
  INV_X1 U21337 ( .A(n18323), .ZN(n18367) );
  NOR2_X1 U21338 ( .A1(n18653), .A2(n18367), .ZN(n18339) );
  AOI22_X1 U21339 ( .A1(n18363), .A2(n18594), .B1(n18654), .B2(n18339), .ZN(
        n18326) );
  INV_X1 U21340 ( .A(n18507), .ZN(n18624) );
  AOI22_X1 U21341 ( .A1(n18626), .A2(n18324), .B1(n18624), .B2(n18323), .ZN(
        n18340) );
  AOI22_X1 U21342 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18340), .B1(
        n18696), .B2(n18655), .ZN(n18325) );
  OAI211_X1 U21343 ( .C1(n18542), .C2(n18404), .A(n18326), .B(n18325), .ZN(
        P3_U2884) );
  AOI22_X1 U21344 ( .A1(n18696), .A2(n18598), .B1(n18662), .B2(n18339), .ZN(
        n18328) );
  AOI22_X1 U21345 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18340), .B1(
        n18664), .B2(n18406), .ZN(n18327) );
  OAI211_X1 U21346 ( .C1(n18361), .C2(n18573), .A(n18328), .B(n18327), .ZN(
        P3_U2885) );
  INV_X1 U21347 ( .A(n18464), .ZN(n18669) );
  AOI22_X1 U21348 ( .A1(n18363), .A2(n18669), .B1(n18668), .B2(n18339), .ZN(
        n18330) );
  AOI22_X1 U21349 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18340), .B1(
        n18670), .B2(n18406), .ZN(n18329) );
  OAI211_X1 U21350 ( .C1(n18711), .C2(n18673), .A(n18330), .B(n18329), .ZN(
        P3_U2886) );
  AOI22_X1 U21351 ( .A1(n18696), .A2(n18606), .B1(n18674), .B2(n18339), .ZN(
        n18332) );
  AOI22_X1 U21352 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18340), .B1(
        n18676), .B2(n18406), .ZN(n18331) );
  OAI211_X1 U21353 ( .C1(n18361), .C2(n18610), .A(n18332), .B(n18331), .ZN(
        P3_U2887) );
  AOI22_X1 U21354 ( .A1(n18696), .A2(n18681), .B1(n18680), .B2(n18339), .ZN(
        n18334) );
  AOI22_X1 U21355 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18340), .B1(
        n18682), .B2(n18406), .ZN(n18333) );
  OAI211_X1 U21356 ( .C1(n18361), .C2(n18685), .A(n18334), .B(n18333), .ZN(
        P3_U2888) );
  AOI22_X1 U21357 ( .A1(n18696), .A2(n18526), .B1(n18687), .B2(n18339), .ZN(
        n18336) );
  AOI22_X1 U21358 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18340), .B1(
        n18689), .B2(n18406), .ZN(n18335) );
  OAI211_X1 U21359 ( .C1(n18361), .C2(n18471), .A(n18336), .B(n18335), .ZN(
        P3_U2889) );
  AOI22_X1 U21360 ( .A1(n18363), .A2(n18694), .B1(n18693), .B2(n18339), .ZN(
        n18338) );
  AOI22_X1 U21361 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18340), .B1(
        n18695), .B2(n18406), .ZN(n18337) );
  OAI211_X1 U21362 ( .C1(n18711), .C2(n18700), .A(n18338), .B(n18337), .ZN(
        P3_U2890) );
  AOI22_X1 U21363 ( .A1(n18696), .A2(n18706), .B1(n18702), .B2(n18339), .ZN(
        n18342) );
  AOI22_X1 U21364 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18340), .B1(
        n18363), .B2(n18703), .ZN(n18341) );
  OAI211_X1 U21365 ( .C1(n18710), .C2(n18404), .A(n18342), .B(n18341), .ZN(
        P3_U2891) );
  NOR2_X1 U21366 ( .A1(n18743), .A2(n18343), .ZN(n18389) );
  AND2_X1 U21367 ( .A1(n18623), .A2(n18389), .ZN(n18362) );
  AOI22_X1 U21368 ( .A1(n18363), .A2(n18655), .B1(n18654), .B2(n18362), .ZN(
        n18348) );
  OAI21_X1 U21369 ( .B1(n18345), .B2(n18344), .A(n18592), .ZN(n18656) );
  NAND2_X1 U21370 ( .A1(n18346), .A2(n18656), .ZN(n18364) );
  NAND2_X1 U21371 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18389), .ZN(
        n18428) );
  INV_X1 U21372 ( .A(n18428), .ZN(n18430) );
  AOI22_X1 U21373 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18364), .B1(
        n18658), .B2(n18430), .ZN(n18347) );
  OAI211_X1 U21374 ( .C1(n18661), .C2(n18381), .A(n18348), .B(n18347), .ZN(
        P3_U2892) );
  AOI22_X1 U21375 ( .A1(n18663), .A2(n18385), .B1(n18662), .B2(n18362), .ZN(
        n18350) );
  AOI22_X1 U21376 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18364), .B1(
        n18664), .B2(n18430), .ZN(n18349) );
  OAI211_X1 U21377 ( .C1(n18361), .C2(n18667), .A(n18350), .B(n18349), .ZN(
        P3_U2893) );
  AOI22_X1 U21378 ( .A1(n18669), .A2(n18385), .B1(n18668), .B2(n18362), .ZN(
        n18352) );
  AOI22_X1 U21379 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18364), .B1(
        n18670), .B2(n18430), .ZN(n18351) );
  OAI211_X1 U21380 ( .C1(n18361), .C2(n18673), .A(n18352), .B(n18351), .ZN(
        P3_U2894) );
  AOI22_X1 U21381 ( .A1(n18675), .A2(n18385), .B1(n18674), .B2(n18362), .ZN(
        n18354) );
  AOI22_X1 U21382 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18364), .B1(
        n18676), .B2(n18430), .ZN(n18353) );
  OAI211_X1 U21383 ( .C1(n18361), .C2(n18679), .A(n18354), .B(n18353), .ZN(
        P3_U2895) );
  INV_X1 U21384 ( .A(n18685), .ZN(n18549) );
  AOI22_X1 U21385 ( .A1(n18549), .A2(n18385), .B1(n18680), .B2(n18362), .ZN(
        n18356) );
  AOI22_X1 U21386 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18364), .B1(
        n18682), .B2(n18430), .ZN(n18355) );
  OAI211_X1 U21387 ( .C1(n18361), .C2(n18552), .A(n18356), .B(n18355), .ZN(
        P3_U2896) );
  AOI22_X1 U21388 ( .A1(n18363), .A2(n18526), .B1(n18687), .B2(n18362), .ZN(
        n18358) );
  AOI22_X1 U21389 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18364), .B1(
        n18689), .B2(n18430), .ZN(n18357) );
  OAI211_X1 U21390 ( .C1(n18471), .C2(n18381), .A(n18358), .B(n18357), .ZN(
        P3_U2897) );
  AOI22_X1 U21391 ( .A1(n18694), .A2(n18385), .B1(n18693), .B2(n18362), .ZN(
        n18360) );
  AOI22_X1 U21392 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18364), .B1(
        n18695), .B2(n18430), .ZN(n18359) );
  OAI211_X1 U21393 ( .C1(n18361), .C2(n18700), .A(n18360), .B(n18359), .ZN(
        P3_U2898) );
  AOI22_X1 U21394 ( .A1(n18703), .A2(n18385), .B1(n18702), .B2(n18362), .ZN(
        n18366) );
  AOI22_X1 U21395 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18364), .B1(
        n18363), .B2(n18706), .ZN(n18365) );
  OAI211_X1 U21396 ( .C1(n18710), .C2(n18428), .A(n18366), .B(n18365), .ZN(
        P3_U2899) );
  NOR2_X2 U21397 ( .A1(n18744), .A2(n18411), .ZN(n18452) );
  INV_X1 U21398 ( .A(n18452), .ZN(n18450) );
  AOI21_X1 U21399 ( .B1(n18428), .B2(n18450), .A(n18653), .ZN(n18384) );
  AOI22_X1 U21400 ( .A1(n18655), .A2(n18385), .B1(n18654), .B2(n18384), .ZN(
        n18370) );
  AOI221_X1 U21401 ( .B1(n18367), .B2(n18428), .C1(n18508), .C2(n18428), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18368) );
  OAI21_X1 U21402 ( .B1(n18452), .B2(n18368), .A(n18568), .ZN(n18386) );
  AOI22_X1 U21403 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18386), .B1(
        n18594), .B2(n18406), .ZN(n18369) );
  OAI211_X1 U21404 ( .C1(n18542), .C2(n18450), .A(n18370), .B(n18369), .ZN(
        P3_U2900) );
  AOI22_X1 U21405 ( .A1(n18663), .A2(n18406), .B1(n18662), .B2(n18384), .ZN(
        n18372) );
  AOI22_X1 U21406 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18386), .B1(
        n18664), .B2(n18452), .ZN(n18371) );
  OAI211_X1 U21407 ( .C1(n18667), .C2(n18381), .A(n18372), .B(n18371), .ZN(
        P3_U2901) );
  AOI22_X1 U21408 ( .A1(n18669), .A2(n18406), .B1(n18668), .B2(n18384), .ZN(
        n18374) );
  AOI22_X1 U21409 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18386), .B1(
        n18670), .B2(n18452), .ZN(n18373) );
  OAI211_X1 U21410 ( .C1(n18673), .C2(n18381), .A(n18374), .B(n18373), .ZN(
        P3_U2902) );
  AOI22_X1 U21411 ( .A1(n18675), .A2(n18406), .B1(n18674), .B2(n18384), .ZN(
        n18376) );
  AOI22_X1 U21412 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18386), .B1(
        n18676), .B2(n18452), .ZN(n18375) );
  OAI211_X1 U21413 ( .C1(n18679), .C2(n18381), .A(n18376), .B(n18375), .ZN(
        P3_U2903) );
  AOI22_X1 U21414 ( .A1(n18549), .A2(n18406), .B1(n18680), .B2(n18384), .ZN(
        n18378) );
  AOI22_X1 U21415 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18386), .B1(
        n18682), .B2(n18452), .ZN(n18377) );
  OAI211_X1 U21416 ( .C1(n18552), .C2(n18381), .A(n18378), .B(n18377), .ZN(
        P3_U2904) );
  AOI22_X1 U21417 ( .A1(n18688), .A2(n18406), .B1(n18687), .B2(n18384), .ZN(
        n18380) );
  AOI22_X1 U21418 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18386), .B1(
        n18689), .B2(n18452), .ZN(n18379) );
  OAI211_X1 U21419 ( .C1(n18692), .C2(n18381), .A(n18380), .B(n18379), .ZN(
        P3_U2905) );
  AOI22_X1 U21420 ( .A1(n18641), .A2(n18385), .B1(n18693), .B2(n18384), .ZN(
        n18383) );
  AOI22_X1 U21421 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18386), .B1(
        n18695), .B2(n18452), .ZN(n18382) );
  OAI211_X1 U21422 ( .C1(n18645), .C2(n18404), .A(n18383), .B(n18382), .ZN(
        P3_U2906) );
  AOI22_X1 U21423 ( .A1(n18703), .A2(n18406), .B1(n18702), .B2(n18384), .ZN(
        n18388) );
  AOI22_X1 U21424 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18386), .B1(
        n18706), .B2(n18385), .ZN(n18387) );
  OAI211_X1 U21425 ( .C1(n18710), .C2(n18450), .A(n18388), .B(n18387), .ZN(
        P3_U2907) );
  NAND2_X1 U21426 ( .A1(n18435), .A2(n18480), .ZN(n18474) );
  NOR2_X1 U21427 ( .A1(n18411), .A2(n18481), .ZN(n18405) );
  AOI22_X1 U21428 ( .A1(n18594), .A2(n18430), .B1(n18654), .B2(n18405), .ZN(
        n18391) );
  AOI22_X1 U21429 ( .A1(n18304), .A2(n18389), .B1(n18435), .B2(n18484), .ZN(
        n18407) );
  AOI22_X1 U21430 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18407), .B1(
        n18655), .B2(n18406), .ZN(n18390) );
  OAI211_X1 U21431 ( .C1(n18542), .C2(n18474), .A(n18391), .B(n18390), .ZN(
        P3_U2908) );
  AOI22_X1 U21432 ( .A1(n18598), .A2(n18406), .B1(n18662), .B2(n18405), .ZN(
        n18393) );
  INV_X1 U21433 ( .A(n18474), .ZN(n18476) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18407), .B1(
        n18664), .B2(n18476), .ZN(n18392) );
  OAI211_X1 U21435 ( .C1(n18573), .C2(n18428), .A(n18393), .B(n18392), .ZN(
        P3_U2909) );
  AOI22_X1 U21436 ( .A1(n18669), .A2(n18430), .B1(n18668), .B2(n18405), .ZN(
        n18395) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18407), .B1(
        n18670), .B2(n18476), .ZN(n18394) );
  OAI211_X1 U21438 ( .C1(n18673), .C2(n18404), .A(n18395), .B(n18394), .ZN(
        P3_U2910) );
  AOI22_X1 U21439 ( .A1(n18675), .A2(n18430), .B1(n18674), .B2(n18405), .ZN(
        n18397) );
  AOI22_X1 U21440 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18407), .B1(
        n18676), .B2(n18476), .ZN(n18396) );
  OAI211_X1 U21441 ( .C1(n18679), .C2(n18404), .A(n18397), .B(n18396), .ZN(
        P3_U2911) );
  AOI22_X1 U21442 ( .A1(n18681), .A2(n18406), .B1(n18680), .B2(n18405), .ZN(
        n18399) );
  AOI22_X1 U21443 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18407), .B1(
        n18682), .B2(n18476), .ZN(n18398) );
  OAI211_X1 U21444 ( .C1(n18685), .C2(n18428), .A(n18399), .B(n18398), .ZN(
        P3_U2912) );
  AOI22_X1 U21445 ( .A1(n18526), .A2(n18406), .B1(n18687), .B2(n18405), .ZN(
        n18401) );
  AOI22_X1 U21446 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18407), .B1(
        n18689), .B2(n18476), .ZN(n18400) );
  OAI211_X1 U21447 ( .C1(n18471), .C2(n18428), .A(n18401), .B(n18400), .ZN(
        P3_U2913) );
  AOI22_X1 U21448 ( .A1(n18694), .A2(n18430), .B1(n18693), .B2(n18405), .ZN(
        n18403) );
  AOI22_X1 U21449 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18407), .B1(
        n18695), .B2(n18476), .ZN(n18402) );
  OAI211_X1 U21450 ( .C1(n18700), .C2(n18404), .A(n18403), .B(n18402), .ZN(
        P3_U2914) );
  AOI22_X1 U21451 ( .A1(n18703), .A2(n18430), .B1(n18702), .B2(n18405), .ZN(
        n18409) );
  AOI22_X1 U21452 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18407), .B1(
        n18706), .B2(n18406), .ZN(n18408) );
  OAI211_X1 U21453 ( .C1(n18710), .C2(n18474), .A(n18409), .B(n18408), .ZN(
        P3_U2915) );
  NOR2_X2 U21454 ( .A1(n18411), .A2(n18410), .ZN(n18502) );
  INV_X1 U21455 ( .A(n18502), .ZN(n18500) );
  NOR2_X1 U21456 ( .A1(n18476), .A2(n18502), .ZN(n18456) );
  NOR2_X1 U21457 ( .A1(n18653), .A2(n18456), .ZN(n18429) );
  AOI22_X1 U21458 ( .A1(n18655), .A2(n18430), .B1(n18654), .B2(n18429), .ZN(
        n18415) );
  NOR2_X1 U21459 ( .A1(n18430), .A2(n18452), .ZN(n18412) );
  OAI21_X1 U21460 ( .B1(n18412), .B2(n18508), .A(n18456), .ZN(n18413) );
  OAI211_X1 U21461 ( .C1(n18502), .C2(n18883), .A(n18568), .B(n18413), .ZN(
        n18431) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18431), .B1(
        n18594), .B2(n18452), .ZN(n18414) );
  OAI211_X1 U21463 ( .C1(n18542), .C2(n18500), .A(n18415), .B(n18414), .ZN(
        P3_U2916) );
  AOI22_X1 U21464 ( .A1(n18598), .A2(n18430), .B1(n18662), .B2(n18429), .ZN(
        n18417) );
  AOI22_X1 U21465 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18431), .B1(
        n18664), .B2(n18502), .ZN(n18416) );
  OAI211_X1 U21466 ( .C1(n18573), .C2(n18450), .A(n18417), .B(n18416), .ZN(
        P3_U2917) );
  AOI22_X1 U21467 ( .A1(n18669), .A2(n18452), .B1(n18668), .B2(n18429), .ZN(
        n18419) );
  AOI22_X1 U21468 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18431), .B1(
        n18670), .B2(n18502), .ZN(n18418) );
  OAI211_X1 U21469 ( .C1(n18673), .C2(n18428), .A(n18419), .B(n18418), .ZN(
        P3_U2918) );
  AOI22_X1 U21470 ( .A1(n18606), .A2(n18430), .B1(n18674), .B2(n18429), .ZN(
        n18421) );
  AOI22_X1 U21471 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18431), .B1(
        n18676), .B2(n18502), .ZN(n18420) );
  OAI211_X1 U21472 ( .C1(n18610), .C2(n18450), .A(n18421), .B(n18420), .ZN(
        P3_U2919) );
  AOI22_X1 U21473 ( .A1(n18681), .A2(n18430), .B1(n18680), .B2(n18429), .ZN(
        n18423) );
  AOI22_X1 U21474 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18431), .B1(
        n18682), .B2(n18502), .ZN(n18422) );
  OAI211_X1 U21475 ( .C1(n18685), .C2(n18450), .A(n18423), .B(n18422), .ZN(
        P3_U2920) );
  AOI22_X1 U21476 ( .A1(n18688), .A2(n18452), .B1(n18687), .B2(n18429), .ZN(
        n18425) );
  AOI22_X1 U21477 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18431), .B1(
        n18689), .B2(n18502), .ZN(n18424) );
  OAI211_X1 U21478 ( .C1(n18692), .C2(n18428), .A(n18425), .B(n18424), .ZN(
        P3_U2921) );
  AOI22_X1 U21479 ( .A1(n18694), .A2(n18452), .B1(n18693), .B2(n18429), .ZN(
        n18427) );
  AOI22_X1 U21480 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18431), .B1(
        n18695), .B2(n18502), .ZN(n18426) );
  OAI211_X1 U21481 ( .C1(n18700), .C2(n18428), .A(n18427), .B(n18426), .ZN(
        P3_U2922) );
  AOI22_X1 U21482 ( .A1(n18703), .A2(n18452), .B1(n18702), .B2(n18429), .ZN(
        n18433) );
  AOI22_X1 U21483 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18431), .B1(
        n18706), .B2(n18430), .ZN(n18432) );
  OAI211_X1 U21484 ( .C1(n18710), .C2(n18500), .A(n18433), .B(n18432), .ZN(
        P3_U2923) );
  NAND2_X1 U21485 ( .A1(n18762), .A2(n18434), .ZN(n18483) );
  NOR2_X2 U21486 ( .A1(n18539), .A2(n18483), .ZN(n18535) );
  INV_X1 U21487 ( .A(n18535), .ZN(n18519) );
  NOR2_X1 U21488 ( .A1(n18653), .A2(n18483), .ZN(n18451) );
  AOI22_X1 U21489 ( .A1(n18594), .A2(n18476), .B1(n18654), .B2(n18451), .ZN(
        n18437) );
  NAND2_X1 U21490 ( .A1(n18435), .A2(n18656), .ZN(n18453) );
  AOI22_X1 U21491 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18453), .B1(
        n18655), .B2(n18452), .ZN(n18436) );
  OAI211_X1 U21492 ( .C1(n18542), .C2(n18519), .A(n18437), .B(n18436), .ZN(
        P3_U2924) );
  AOI22_X1 U21493 ( .A1(n18663), .A2(n18476), .B1(n18662), .B2(n18451), .ZN(
        n18439) );
  AOI22_X1 U21494 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18453), .B1(
        n18664), .B2(n18535), .ZN(n18438) );
  OAI211_X1 U21495 ( .C1(n18667), .C2(n18450), .A(n18439), .B(n18438), .ZN(
        P3_U2925) );
  AOI22_X1 U21496 ( .A1(n18602), .A2(n18452), .B1(n18668), .B2(n18451), .ZN(
        n18441) );
  AOI22_X1 U21497 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18453), .B1(
        n18670), .B2(n18535), .ZN(n18440) );
  OAI211_X1 U21498 ( .C1(n18464), .C2(n18474), .A(n18441), .B(n18440), .ZN(
        P3_U2926) );
  AOI22_X1 U21499 ( .A1(n18675), .A2(n18476), .B1(n18674), .B2(n18451), .ZN(
        n18443) );
  AOI22_X1 U21500 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18453), .B1(
        n18676), .B2(n18535), .ZN(n18442) );
  OAI211_X1 U21501 ( .C1(n18679), .C2(n18450), .A(n18443), .B(n18442), .ZN(
        P3_U2927) );
  AOI22_X1 U21502 ( .A1(n18549), .A2(n18476), .B1(n18680), .B2(n18451), .ZN(
        n18445) );
  AOI22_X1 U21503 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18453), .B1(
        n18682), .B2(n18535), .ZN(n18444) );
  OAI211_X1 U21504 ( .C1(n18552), .C2(n18450), .A(n18445), .B(n18444), .ZN(
        P3_U2928) );
  AOI22_X1 U21505 ( .A1(n18688), .A2(n18476), .B1(n18687), .B2(n18451), .ZN(
        n18447) );
  AOI22_X1 U21506 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18453), .B1(
        n18689), .B2(n18535), .ZN(n18446) );
  OAI211_X1 U21507 ( .C1(n18692), .C2(n18450), .A(n18447), .B(n18446), .ZN(
        P3_U2929) );
  AOI22_X1 U21508 ( .A1(n18694), .A2(n18476), .B1(n18693), .B2(n18451), .ZN(
        n18449) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18453), .B1(
        n18695), .B2(n18535), .ZN(n18448) );
  OAI211_X1 U21510 ( .C1(n18700), .C2(n18450), .A(n18449), .B(n18448), .ZN(
        P3_U2930) );
  AOI22_X1 U21511 ( .A1(n18703), .A2(n18476), .B1(n18702), .B2(n18451), .ZN(
        n18455) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18453), .B1(
        n18706), .B2(n18452), .ZN(n18454) );
  OAI211_X1 U21513 ( .C1(n18710), .C2(n18519), .A(n18455), .B(n18454), .ZN(
        P3_U2931) );
  NOR2_X2 U21514 ( .A1(n18744), .A2(n18482), .ZN(n18559) );
  INV_X1 U21515 ( .A(n18559), .ZN(n18557) );
  NOR2_X1 U21516 ( .A1(n18535), .A2(n18559), .ZN(n18510) );
  NOR2_X1 U21517 ( .A1(n18653), .A2(n18510), .ZN(n18475) );
  AOI22_X1 U21518 ( .A1(n18594), .A2(n18502), .B1(n18654), .B2(n18475), .ZN(
        n18459) );
  OAI21_X1 U21519 ( .B1(n18456), .B2(n18508), .A(n18510), .ZN(n18457) );
  OAI211_X1 U21520 ( .C1(n18559), .C2(n18883), .A(n18568), .B(n18457), .ZN(
        n18477) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18477), .B1(
        n18655), .B2(n18476), .ZN(n18458) );
  OAI211_X1 U21522 ( .C1(n18542), .C2(n18557), .A(n18459), .B(n18458), .ZN(
        P3_U2932) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18477), .B1(
        n18662), .B2(n18475), .ZN(n18461) );
  AOI22_X1 U21524 ( .A1(n18664), .A2(n18559), .B1(n18598), .B2(n18476), .ZN(
        n18460) );
  OAI211_X1 U21525 ( .C1(n18573), .C2(n18500), .A(n18461), .B(n18460), .ZN(
        P3_U2933) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18477), .B1(
        n18668), .B2(n18475), .ZN(n18463) );
  AOI22_X1 U21527 ( .A1(n18670), .A2(n18559), .B1(n18602), .B2(n18476), .ZN(
        n18462) );
  OAI211_X1 U21528 ( .C1(n18464), .C2(n18500), .A(n18463), .B(n18462), .ZN(
        P3_U2934) );
  AOI22_X1 U21529 ( .A1(n18675), .A2(n18502), .B1(n18674), .B2(n18475), .ZN(
        n18466) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18477), .B1(
        n18676), .B2(n18559), .ZN(n18465) );
  OAI211_X1 U21531 ( .C1(n18679), .C2(n18474), .A(n18466), .B(n18465), .ZN(
        P3_U2935) );
  AOI22_X1 U21532 ( .A1(n18549), .A2(n18502), .B1(n18680), .B2(n18475), .ZN(
        n18468) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18477), .B1(
        n18682), .B2(n18559), .ZN(n18467) );
  OAI211_X1 U21534 ( .C1(n18552), .C2(n18474), .A(n18468), .B(n18467), .ZN(
        P3_U2936) );
  AOI22_X1 U21535 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18477), .B1(
        n18687), .B2(n18475), .ZN(n18470) );
  AOI22_X1 U21536 ( .A1(n18689), .A2(n18559), .B1(n18526), .B2(n18476), .ZN(
        n18469) );
  OAI211_X1 U21537 ( .C1(n18471), .C2(n18500), .A(n18470), .B(n18469), .ZN(
        P3_U2937) );
  AOI22_X1 U21538 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18477), .B1(
        n18693), .B2(n18475), .ZN(n18473) );
  AOI22_X1 U21539 ( .A1(n18694), .A2(n18502), .B1(n18695), .B2(n18559), .ZN(
        n18472) );
  OAI211_X1 U21540 ( .C1(n18700), .C2(n18474), .A(n18473), .B(n18472), .ZN(
        P3_U2938) );
  AOI22_X1 U21541 ( .A1(n18703), .A2(n18502), .B1(n18702), .B2(n18475), .ZN(
        n18479) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18477), .B1(
        n18706), .B2(n18476), .ZN(n18478) );
  OAI211_X1 U21543 ( .C1(n18710), .C2(n18557), .A(n18479), .B(n18478), .ZN(
        P3_U2939) );
  NAND2_X1 U21544 ( .A1(n18563), .A2(n18480), .ZN(n18582) );
  NOR2_X1 U21545 ( .A1(n18482), .A2(n18481), .ZN(n18501) );
  AOI22_X1 U21546 ( .A1(n18655), .A2(n18502), .B1(n18654), .B2(n18501), .ZN(
        n18487) );
  INV_X1 U21547 ( .A(n18483), .ZN(n18485) );
  AOI22_X1 U21548 ( .A1(n18304), .A2(n18485), .B1(n18563), .B2(n18484), .ZN(
        n18503) );
  AOI22_X1 U21549 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18503), .B1(
        n18594), .B2(n18535), .ZN(n18486) );
  OAI211_X1 U21550 ( .C1(n18542), .C2(n18582), .A(n18487), .B(n18486), .ZN(
        P3_U2940) );
  AOI22_X1 U21551 ( .A1(n18598), .A2(n18502), .B1(n18662), .B2(n18501), .ZN(
        n18489) );
  INV_X1 U21552 ( .A(n18582), .ZN(n18586) );
  AOI22_X1 U21553 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18503), .B1(
        n18664), .B2(n18586), .ZN(n18488) );
  OAI211_X1 U21554 ( .C1(n18573), .C2(n18519), .A(n18489), .B(n18488), .ZN(
        P3_U2941) );
  AOI22_X1 U21555 ( .A1(n18669), .A2(n18535), .B1(n18668), .B2(n18501), .ZN(
        n18491) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18503), .B1(
        n18670), .B2(n18586), .ZN(n18490) );
  OAI211_X1 U21557 ( .C1(n18673), .C2(n18500), .A(n18491), .B(n18490), .ZN(
        P3_U2942) );
  AOI22_X1 U21558 ( .A1(n18606), .A2(n18502), .B1(n18674), .B2(n18501), .ZN(
        n18493) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18503), .B1(
        n18676), .B2(n18586), .ZN(n18492) );
  OAI211_X1 U21560 ( .C1(n18610), .C2(n18519), .A(n18493), .B(n18492), .ZN(
        P3_U2943) );
  AOI22_X1 U21561 ( .A1(n18549), .A2(n18535), .B1(n18680), .B2(n18501), .ZN(
        n18495) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18503), .B1(
        n18682), .B2(n18586), .ZN(n18494) );
  OAI211_X1 U21563 ( .C1(n18552), .C2(n18500), .A(n18495), .B(n18494), .ZN(
        P3_U2944) );
  AOI22_X1 U21564 ( .A1(n18688), .A2(n18535), .B1(n18687), .B2(n18501), .ZN(
        n18497) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18503), .B1(
        n18689), .B2(n18586), .ZN(n18496) );
  OAI211_X1 U21566 ( .C1(n18692), .C2(n18500), .A(n18497), .B(n18496), .ZN(
        P3_U2945) );
  AOI22_X1 U21567 ( .A1(n18694), .A2(n18535), .B1(n18693), .B2(n18501), .ZN(
        n18499) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18503), .B1(
        n18695), .B2(n18586), .ZN(n18498) );
  OAI211_X1 U21569 ( .C1(n18700), .C2(n18500), .A(n18499), .B(n18498), .ZN(
        P3_U2946) );
  AOI22_X1 U21570 ( .A1(n18703), .A2(n18535), .B1(n18702), .B2(n18501), .ZN(
        n18505) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18503), .B1(
        n18706), .B2(n18502), .ZN(n18504) );
  OAI211_X1 U21572 ( .C1(n18710), .C2(n18582), .A(n18505), .B(n18504), .ZN(
        P3_U2947) );
  NAND2_X1 U21573 ( .A1(n18563), .A2(n18506), .ZN(n18617) );
  INV_X1 U21574 ( .A(n18617), .ZN(n18619) );
  NOR2_X1 U21575 ( .A1(n18586), .A2(n18619), .ZN(n18509) );
  AOI21_X1 U21576 ( .B1(n18582), .B2(n18617), .A(n18653), .ZN(n18534) );
  AOI22_X1 U21577 ( .A1(n18655), .A2(n18535), .B1(n18654), .B2(n18534), .ZN(
        n18512) );
  AOI22_X1 U21578 ( .A1(n18594), .A2(n18559), .B1(n18658), .B2(n18619), .ZN(
        n18511) );
  OAI211_X1 U21579 ( .C1(n18533), .C2(n18513), .A(n18512), .B(n18511), .ZN(
        P3_U2948) );
  AOI22_X1 U21580 ( .A1(n18598), .A2(n18535), .B1(n18662), .B2(n18534), .ZN(
        n18515) );
  AOI22_X1 U21581 ( .A1(n18663), .A2(n18559), .B1(n18664), .B2(n18619), .ZN(
        n18514) );
  OAI211_X1 U21582 ( .C1(n18533), .C2(n18516), .A(n18515), .B(n18514), .ZN(
        P3_U2949) );
  AOI22_X1 U21583 ( .A1(n18669), .A2(n18559), .B1(n18668), .B2(n18534), .ZN(
        n18518) );
  INV_X1 U21584 ( .A(n18533), .ZN(n18536) );
  AOI22_X1 U21585 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18536), .B1(
        n18670), .B2(n18619), .ZN(n18517) );
  OAI211_X1 U21586 ( .C1(n18673), .C2(n18519), .A(n18518), .B(n18517), .ZN(
        P3_U2950) );
  AOI22_X1 U21587 ( .A1(n18675), .A2(n18559), .B1(n18674), .B2(n18534), .ZN(
        n18521) );
  AOI22_X1 U21588 ( .A1(n18676), .A2(n18619), .B1(n18606), .B2(n18535), .ZN(
        n18520) );
  OAI211_X1 U21589 ( .C1(n18533), .C2(n18522), .A(n18521), .B(n18520), .ZN(
        P3_U2951) );
  AOI22_X1 U21590 ( .A1(n18549), .A2(n18559), .B1(n18680), .B2(n18534), .ZN(
        n18524) );
  AOI22_X1 U21591 ( .A1(n18682), .A2(n18619), .B1(n18681), .B2(n18535), .ZN(
        n18523) );
  OAI211_X1 U21592 ( .C1(n18533), .C2(n18525), .A(n18524), .B(n18523), .ZN(
        P3_U2952) );
  AOI22_X1 U21593 ( .A1(n18688), .A2(n18559), .B1(n18687), .B2(n18534), .ZN(
        n18528) );
  AOI22_X1 U21594 ( .A1(n18689), .A2(n18619), .B1(n18526), .B2(n18535), .ZN(
        n18527) );
  OAI211_X1 U21595 ( .C1(n18533), .C2(n18529), .A(n18528), .B(n18527), .ZN(
        P3_U2953) );
  AOI22_X1 U21596 ( .A1(n18641), .A2(n18535), .B1(n18693), .B2(n18534), .ZN(
        n18531) );
  AOI22_X1 U21597 ( .A1(n18694), .A2(n18559), .B1(n18695), .B2(n18619), .ZN(
        n18530) );
  OAI211_X1 U21598 ( .C1(n18533), .C2(n18532), .A(n18531), .B(n18530), .ZN(
        P3_U2954) );
  AOI22_X1 U21599 ( .A1(n18703), .A2(n18559), .B1(n18702), .B2(n18534), .ZN(
        n18538) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18536), .B1(
        n18706), .B2(n18535), .ZN(n18537) );
  OAI211_X1 U21601 ( .C1(n18710), .C2(n18617), .A(n18538), .B(n18537), .ZN(
        P3_U2955) );
  NAND2_X1 U21602 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18563), .ZN(
        n18591) );
  NOR2_X2 U21603 ( .A1(n18539), .A2(n18591), .ZN(n18647) );
  INV_X1 U21604 ( .A(n18647), .ZN(n18640) );
  NOR2_X1 U21605 ( .A1(n18653), .A2(n18591), .ZN(n18558) );
  AOI22_X1 U21606 ( .A1(n18594), .A2(n18586), .B1(n18654), .B2(n18558), .ZN(
        n18541) );
  NAND2_X1 U21607 ( .A1(n18563), .A2(n18656), .ZN(n18560) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18560), .B1(
        n18655), .B2(n18559), .ZN(n18540) );
  OAI211_X1 U21609 ( .C1(n18542), .C2(n18640), .A(n18541), .B(n18540), .ZN(
        P3_U2956) );
  AOI22_X1 U21610 ( .A1(n18663), .A2(n18586), .B1(n18662), .B2(n18558), .ZN(
        n18544) );
  AOI22_X1 U21611 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18560), .B1(
        n18664), .B2(n18647), .ZN(n18543) );
  OAI211_X1 U21612 ( .C1(n18667), .C2(n18557), .A(n18544), .B(n18543), .ZN(
        P3_U2957) );
  AOI22_X1 U21613 ( .A1(n18669), .A2(n18586), .B1(n18668), .B2(n18558), .ZN(
        n18546) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18560), .B1(
        n18670), .B2(n18647), .ZN(n18545) );
  OAI211_X1 U21615 ( .C1(n18673), .C2(n18557), .A(n18546), .B(n18545), .ZN(
        P3_U2958) );
  AOI22_X1 U21616 ( .A1(n18606), .A2(n18559), .B1(n18674), .B2(n18558), .ZN(
        n18548) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18560), .B1(
        n18676), .B2(n18647), .ZN(n18547) );
  OAI211_X1 U21618 ( .C1(n18610), .C2(n18582), .A(n18548), .B(n18547), .ZN(
        P3_U2959) );
  AOI22_X1 U21619 ( .A1(n18549), .A2(n18586), .B1(n18680), .B2(n18558), .ZN(
        n18551) );
  AOI22_X1 U21620 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18560), .B1(
        n18682), .B2(n18647), .ZN(n18550) );
  OAI211_X1 U21621 ( .C1(n18552), .C2(n18557), .A(n18551), .B(n18550), .ZN(
        P3_U2960) );
  AOI22_X1 U21622 ( .A1(n18688), .A2(n18586), .B1(n18687), .B2(n18558), .ZN(
        n18554) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18560), .B1(
        n18689), .B2(n18647), .ZN(n18553) );
  OAI211_X1 U21624 ( .C1(n18692), .C2(n18557), .A(n18554), .B(n18553), .ZN(
        P3_U2961) );
  AOI22_X1 U21625 ( .A1(n18694), .A2(n18586), .B1(n18693), .B2(n18558), .ZN(
        n18556) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18560), .B1(
        n18695), .B2(n18647), .ZN(n18555) );
  OAI211_X1 U21627 ( .C1(n18700), .C2(n18557), .A(n18556), .B(n18555), .ZN(
        P3_U2962) );
  AOI22_X1 U21628 ( .A1(n18706), .A2(n18559), .B1(n18702), .B2(n18558), .ZN(
        n18562) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18560), .B1(
        n18703), .B2(n18586), .ZN(n18561) );
  OAI211_X1 U21630 ( .C1(n18710), .C2(n18640), .A(n18562), .B(n18561), .ZN(
        P3_U2963) );
  NOR2_X2 U21631 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18593), .ZN(
        n18705) );
  INV_X1 U21632 ( .A(n18705), .ZN(n18699) );
  NAND2_X1 U21633 ( .A1(n18640), .A2(n18699), .ZN(n18625) );
  INV_X1 U21634 ( .A(n18625), .ZN(n18564) );
  NOR2_X1 U21635 ( .A1(n18653), .A2(n18564), .ZN(n18585) );
  AOI22_X1 U21636 ( .A1(n18655), .A2(n18586), .B1(n18654), .B2(n18585), .ZN(
        n18570) );
  NAND2_X1 U21637 ( .A1(n18626), .A2(n18563), .ZN(n18565) );
  OAI21_X1 U21638 ( .B1(n18566), .B2(n18565), .A(n18564), .ZN(n18567) );
  OAI211_X1 U21639 ( .C1(n18705), .C2(n18883), .A(n18568), .B(n18567), .ZN(
        n18587) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18587), .B1(
        n18658), .B2(n18705), .ZN(n18569) );
  OAI211_X1 U21641 ( .C1(n18661), .C2(n18617), .A(n18570), .B(n18569), .ZN(
        P3_U2964) );
  AOI22_X1 U21642 ( .A1(n18598), .A2(n18586), .B1(n18662), .B2(n18585), .ZN(
        n18572) );
  AOI22_X1 U21643 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18587), .B1(
        n18664), .B2(n18705), .ZN(n18571) );
  OAI211_X1 U21644 ( .C1(n18573), .C2(n18617), .A(n18572), .B(n18571), .ZN(
        P3_U2965) );
  AOI22_X1 U21645 ( .A1(n18669), .A2(n18619), .B1(n18668), .B2(n18585), .ZN(
        n18575) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18587), .B1(
        n18670), .B2(n18705), .ZN(n18574) );
  OAI211_X1 U21647 ( .C1(n18673), .C2(n18582), .A(n18575), .B(n18574), .ZN(
        P3_U2966) );
  AOI22_X1 U21648 ( .A1(n18675), .A2(n18619), .B1(n18674), .B2(n18585), .ZN(
        n18577) );
  AOI22_X1 U21649 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18587), .B1(
        n18676), .B2(n18705), .ZN(n18576) );
  OAI211_X1 U21650 ( .C1(n18679), .C2(n18582), .A(n18577), .B(n18576), .ZN(
        P3_U2967) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18587), .B1(
        n18680), .B2(n18585), .ZN(n18579) );
  AOI22_X1 U21652 ( .A1(n18682), .A2(n18705), .B1(n18681), .B2(n18586), .ZN(
        n18578) );
  OAI211_X1 U21653 ( .C1(n18685), .C2(n18617), .A(n18579), .B(n18578), .ZN(
        P3_U2968) );
  AOI22_X1 U21654 ( .A1(n18688), .A2(n18619), .B1(n18687), .B2(n18585), .ZN(
        n18581) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18587), .B1(
        n18689), .B2(n18705), .ZN(n18580) );
  OAI211_X1 U21656 ( .C1(n18692), .C2(n18582), .A(n18581), .B(n18580), .ZN(
        P3_U2969) );
  AOI22_X1 U21657 ( .A1(n18641), .A2(n18586), .B1(n18693), .B2(n18585), .ZN(
        n18584) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18587), .B1(
        n18695), .B2(n18705), .ZN(n18583) );
  OAI211_X1 U21659 ( .C1(n18645), .C2(n18617), .A(n18584), .B(n18583), .ZN(
        P3_U2970) );
  AOI22_X1 U21660 ( .A1(n18706), .A2(n18586), .B1(n18702), .B2(n18585), .ZN(
        n18589) );
  AOI22_X1 U21661 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18587), .B1(
        n18703), .B2(n18619), .ZN(n18588) );
  OAI211_X1 U21662 ( .C1(n18710), .C2(n18699), .A(n18589), .B(n18588), .ZN(
        P3_U2971) );
  OAI22_X1 U21663 ( .A1(n18592), .A2(n18591), .B1(n18593), .B2(n18590), .ZN(
        n18607) );
  NOR2_X1 U21664 ( .A1(n18653), .A2(n18593), .ZN(n18618) );
  AOI22_X1 U21665 ( .A1(n18655), .A2(n18619), .B1(n18654), .B2(n18618), .ZN(
        n18596) );
  AOI22_X1 U21666 ( .A1(n18594), .A2(n18647), .B1(n18658), .B2(n18704), .ZN(
        n18595) );
  OAI211_X1 U21667 ( .C1(n18597), .C2(n18607), .A(n18596), .B(n18595), .ZN(
        P3_U2972) );
  AOI22_X1 U21668 ( .A1(n18663), .A2(n18647), .B1(n18662), .B2(n18618), .ZN(
        n18600) );
  AOI22_X1 U21669 ( .A1(n18704), .A2(n18664), .B1(n18598), .B2(n18619), .ZN(
        n18599) );
  OAI211_X1 U21670 ( .C1(n18601), .C2(n18607), .A(n18600), .B(n18599), .ZN(
        P3_U2973) );
  AOI22_X1 U21671 ( .A1(n18602), .A2(n18619), .B1(n18668), .B2(n18618), .ZN(
        n18604) );
  AOI22_X1 U21672 ( .A1(n18704), .A2(n18670), .B1(n18669), .B2(n18647), .ZN(
        n18603) );
  OAI211_X1 U21673 ( .C1(n18605), .C2(n18607), .A(n18604), .B(n18603), .ZN(
        P3_U2974) );
  AOI22_X1 U21674 ( .A1(n18606), .A2(n18619), .B1(n18674), .B2(n18618), .ZN(
        n18609) );
  INV_X1 U21675 ( .A(n18607), .ZN(n18620) );
  AOI22_X1 U21676 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18620), .B1(
        n18704), .B2(n18676), .ZN(n18608) );
  OAI211_X1 U21677 ( .C1(n18610), .C2(n18640), .A(n18609), .B(n18608), .ZN(
        P3_U2975) );
  AOI22_X1 U21678 ( .A1(n18681), .A2(n18619), .B1(n18680), .B2(n18618), .ZN(
        n18612) );
  AOI22_X1 U21679 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18620), .B1(
        n18704), .B2(n18682), .ZN(n18611) );
  OAI211_X1 U21680 ( .C1(n18685), .C2(n18640), .A(n18612), .B(n18611), .ZN(
        P3_U2976) );
  AOI22_X1 U21681 ( .A1(n18688), .A2(n18647), .B1(n18687), .B2(n18618), .ZN(
        n18614) );
  AOI22_X1 U21682 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18620), .B1(
        n18704), .B2(n18689), .ZN(n18613) );
  OAI211_X1 U21683 ( .C1(n18692), .C2(n18617), .A(n18614), .B(n18613), .ZN(
        P3_U2977) );
  AOI22_X1 U21684 ( .A1(n18694), .A2(n18647), .B1(n18693), .B2(n18618), .ZN(
        n18616) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18620), .B1(
        n18704), .B2(n18695), .ZN(n18615) );
  OAI211_X1 U21686 ( .C1(n18700), .C2(n18617), .A(n18616), .B(n18615), .ZN(
        P3_U2978) );
  INV_X1 U21687 ( .A(n18704), .ZN(n18686) );
  AOI22_X1 U21688 ( .A1(n18706), .A2(n18619), .B1(n18702), .B2(n18618), .ZN(
        n18622) );
  AOI22_X1 U21689 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18620), .B1(
        n18703), .B2(n18647), .ZN(n18621) );
  OAI211_X1 U21690 ( .C1(n18686), .C2(n18710), .A(n18622), .B(n18621), .ZN(
        P3_U2979) );
  AND2_X1 U21691 ( .A1(n18623), .A2(n18627), .ZN(n18646) );
  AOI22_X1 U21692 ( .A1(n18655), .A2(n18647), .B1(n18654), .B2(n18646), .ZN(
        n18629) );
  OAI221_X1 U21693 ( .B1(n18627), .B2(n18626), .C1(n18627), .C2(n18625), .A(
        n18624), .ZN(n18648) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18648), .B1(
        n18642), .B2(n18658), .ZN(n18628) );
  OAI211_X1 U21695 ( .C1(n18661), .C2(n18699), .A(n18629), .B(n18628), .ZN(
        P3_U2980) );
  AOI22_X1 U21696 ( .A1(n18663), .A2(n18705), .B1(n18662), .B2(n18646), .ZN(
        n18631) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18648), .B1(
        n18642), .B2(n18664), .ZN(n18630) );
  OAI211_X1 U21698 ( .C1(n18667), .C2(n18640), .A(n18631), .B(n18630), .ZN(
        P3_U2981) );
  AOI22_X1 U21699 ( .A1(n18669), .A2(n18705), .B1(n18668), .B2(n18646), .ZN(
        n18633) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18648), .B1(
        n18642), .B2(n18670), .ZN(n18632) );
  OAI211_X1 U21701 ( .C1(n18673), .C2(n18640), .A(n18633), .B(n18632), .ZN(
        P3_U2982) );
  AOI22_X1 U21702 ( .A1(n18675), .A2(n18705), .B1(n18674), .B2(n18646), .ZN(
        n18635) );
  AOI22_X1 U21703 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18648), .B1(
        n18642), .B2(n18676), .ZN(n18634) );
  OAI211_X1 U21704 ( .C1(n18679), .C2(n18640), .A(n18635), .B(n18634), .ZN(
        P3_U2983) );
  AOI22_X1 U21705 ( .A1(n18681), .A2(n18647), .B1(n18680), .B2(n18646), .ZN(
        n18637) );
  AOI22_X1 U21706 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18648), .B1(
        n18642), .B2(n18682), .ZN(n18636) );
  OAI211_X1 U21707 ( .C1(n18685), .C2(n18699), .A(n18637), .B(n18636), .ZN(
        P3_U2984) );
  AOI22_X1 U21708 ( .A1(n18688), .A2(n18705), .B1(n18687), .B2(n18646), .ZN(
        n18639) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18648), .B1(
        n18642), .B2(n18689), .ZN(n18638) );
  OAI211_X1 U21710 ( .C1(n18692), .C2(n18640), .A(n18639), .B(n18638), .ZN(
        P3_U2985) );
  AOI22_X1 U21711 ( .A1(n18641), .A2(n18647), .B1(n18693), .B2(n18646), .ZN(
        n18644) );
  AOI22_X1 U21712 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18648), .B1(
        n18642), .B2(n18695), .ZN(n18643) );
  OAI211_X1 U21713 ( .C1(n18645), .C2(n18699), .A(n18644), .B(n18643), .ZN(
        P3_U2986) );
  AOI22_X1 U21714 ( .A1(n18706), .A2(n18647), .B1(n18702), .B2(n18646), .ZN(
        n18650) );
  AOI22_X1 U21715 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18648), .B1(
        n18703), .B2(n18705), .ZN(n18649) );
  OAI211_X1 U21716 ( .C1(n18651), .C2(n18710), .A(n18650), .B(n18649), .ZN(
        P3_U2987) );
  NOR2_X1 U21717 ( .A1(n18653), .A2(n18652), .ZN(n18701) );
  AOI22_X1 U21718 ( .A1(n18655), .A2(n18705), .B1(n18654), .B2(n18701), .ZN(
        n18660) );
  NAND2_X1 U21719 ( .A1(n18657), .A2(n18656), .ZN(n18707) );
  AOI22_X1 U21720 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18707), .B1(
        n18696), .B2(n18658), .ZN(n18659) );
  OAI211_X1 U21721 ( .C1(n18661), .C2(n18686), .A(n18660), .B(n18659), .ZN(
        P3_U2988) );
  AOI22_X1 U21722 ( .A1(n18704), .A2(n18663), .B1(n18662), .B2(n18701), .ZN(
        n18666) );
  AOI22_X1 U21723 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18707), .B1(
        n18696), .B2(n18664), .ZN(n18665) );
  OAI211_X1 U21724 ( .C1(n18667), .C2(n18699), .A(n18666), .B(n18665), .ZN(
        P3_U2989) );
  AOI22_X1 U21725 ( .A1(n18704), .A2(n18669), .B1(n18668), .B2(n18701), .ZN(
        n18672) );
  AOI22_X1 U21726 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18707), .B1(
        n18696), .B2(n18670), .ZN(n18671) );
  OAI211_X1 U21727 ( .C1(n18673), .C2(n18699), .A(n18672), .B(n18671), .ZN(
        P3_U2990) );
  AOI22_X1 U21728 ( .A1(n18704), .A2(n18675), .B1(n18674), .B2(n18701), .ZN(
        n18678) );
  AOI22_X1 U21729 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18707), .B1(
        n18696), .B2(n18676), .ZN(n18677) );
  OAI211_X1 U21730 ( .C1(n18679), .C2(n18699), .A(n18678), .B(n18677), .ZN(
        P3_U2991) );
  AOI22_X1 U21731 ( .A1(n18681), .A2(n18705), .B1(n18680), .B2(n18701), .ZN(
        n18684) );
  AOI22_X1 U21732 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18707), .B1(
        n18696), .B2(n18682), .ZN(n18683) );
  OAI211_X1 U21733 ( .C1(n18686), .C2(n18685), .A(n18684), .B(n18683), .ZN(
        P3_U2992) );
  AOI22_X1 U21734 ( .A1(n18688), .A2(n18704), .B1(n18687), .B2(n18701), .ZN(
        n18691) );
  AOI22_X1 U21735 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18707), .B1(
        n18696), .B2(n18689), .ZN(n18690) );
  OAI211_X1 U21736 ( .C1(n18692), .C2(n18699), .A(n18691), .B(n18690), .ZN(
        P3_U2993) );
  AOI22_X1 U21737 ( .A1(n18694), .A2(n18704), .B1(n18693), .B2(n18701), .ZN(
        n18698) );
  AOI22_X1 U21738 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18707), .B1(
        n18696), .B2(n18695), .ZN(n18697) );
  OAI211_X1 U21739 ( .C1(n18700), .C2(n18699), .A(n18698), .B(n18697), .ZN(
        P3_U2994) );
  AOI22_X1 U21740 ( .A1(n18704), .A2(n18703), .B1(n18702), .B2(n18701), .ZN(
        n18709) );
  AOI22_X1 U21741 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18707), .B1(
        n18706), .B2(n18705), .ZN(n18708) );
  OAI211_X1 U21742 ( .C1(n18711), .C2(n18710), .A(n18709), .B(n18708), .ZN(
        P3_U2995) );
  INV_X1 U21743 ( .A(n18712), .ZN(n18729) );
  OAI21_X1 U21744 ( .B1(n18715), .B2(n18714), .A(n18713), .ZN(n18726) );
  AOI22_X1 U21745 ( .A1(n18729), .A2(n18717), .B1(n18716), .B2(n18726), .ZN(
        n18719) );
  NAND2_X1 U21746 ( .A1(n18719), .A2(n18718), .ZN(n18887) );
  NOR2_X1 U21747 ( .A1(n18766), .A2(n18887), .ZN(n18724) );
  NOR3_X1 U21748 ( .A1(n18727), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        n18720), .ZN(n18741) );
  OAI22_X1 U21749 ( .A1(n18741), .A2(n18729), .B1(n18722), .B2(n18721), .ZN(
        n18884) );
  NAND2_X1 U21750 ( .A1(n12014), .A2(n18884), .ZN(n18723) );
  OAI22_X1 U21751 ( .A1(n18724), .A2(n12014), .B1(n18766), .B2(n18723), .ZN(
        n18774) );
  AOI21_X1 U21752 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18738), .A(
        n18727), .ZN(n18725) );
  NOR3_X1 U21753 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18725), .A3(
        n12023), .ZN(n18735) );
  AOI21_X1 U21754 ( .B1(n12023), .B2(n18727), .A(n18726), .ZN(n18733) );
  NAND2_X1 U21755 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18728), .ZN(
        n18732) );
  OAI211_X1 U21756 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n18730), .B(n18729), .ZN(
        n18731) );
  OAI21_X1 U21757 ( .B1(n18733), .B2(n18732), .A(n18731), .ZN(n18734) );
  AOI211_X1 U21758 ( .C1(n18751), .C2(n18736), .A(n18735), .B(n18734), .ZN(
        n18893) );
  INV_X1 U21759 ( .A(n18766), .ZN(n18737) );
  AOI22_X1 U21760 ( .A1(n18766), .A2(n18897), .B1(n18893), .B2(n18737), .ZN(
        n18760) );
  NOR2_X1 U21761 ( .A1(n18739), .A2(n18738), .ZN(n18742) );
  AOI22_X1 U21762 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18740), .B1(
        n18742), .B2(n18912), .ZN(n18746) );
  OAI22_X1 U21763 ( .A1(n18742), .A2(n18898), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18741), .ZN(n18903) );
  AOI21_X1 U21764 ( .B1(n18746), .B2(n18743), .A(n18903), .ZN(n18745) );
  OAI21_X1 U21765 ( .B1(n18766), .B2(n18745), .A(n18744), .ZN(n18748) );
  INV_X1 U21766 ( .A(n18746), .ZN(n18906) );
  NAND3_X1 U21767 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n18906), .ZN(n18747) );
  OAI211_X1 U21768 ( .C1(n18761), .C2(n18760), .A(n18748), .B(n18747), .ZN(
        n18758) );
  INV_X1 U21769 ( .A(n18760), .ZN(n18749) );
  OAI221_X1 U21770 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n18758), .A(n18749), .ZN(
        n18773) );
  NOR2_X1 U21771 ( .A1(n18751), .A2(n18750), .ZN(n18753) );
  OAI222_X1 U21772 ( .A1(n18757), .A2(n18756), .B1(n18755), .B2(n18754), .C1(
        n18753), .C2(n18752), .ZN(n18925) );
  INV_X1 U21773 ( .A(n18758), .ZN(n18759) );
  AOI21_X1 U21774 ( .B1(n18761), .B2(n18760), .A(n18759), .ZN(n18771) );
  NAND2_X1 U21775 ( .A1(n18763), .A2(n18762), .ZN(n18770) );
  AOI211_X1 U21776 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18766), .A(
        n18765), .B(n18764), .ZN(n18769) );
  OAI21_X1 U21777 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18767), .ZN(n18768) );
  OAI211_X1 U21778 ( .C1(n18771), .C2(n18770), .A(n18769), .B(n18768), .ZN(
        n18772) );
  AOI211_X1 U21779 ( .C1(n18774), .C2(n18773), .A(n18925), .B(n18772), .ZN(
        n18782) );
  AOI22_X1 U21780 ( .A1(n18909), .A2(n18935), .B1(n18785), .B2(n18929), .ZN(
        n18779) );
  OAI211_X1 U21781 ( .C1(n18776), .C2(n18775), .A(n18927), .B(n18782), .ZN(
        n18882) );
  OAI211_X1 U21782 ( .C1(P3_STATE2_REG_2__SCAN_IN), .C2(n18933), .A(n18777), 
        .B(n18882), .ZN(n18787) );
  OAI22_X1 U21783 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18779), .B1(n18778), 
        .B2(n18787), .ZN(n18780) );
  OAI21_X1 U21784 ( .B1(n18782), .B2(n18781), .A(n18780), .ZN(P3_U2996) );
  NOR4_X1 U21785 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18783), .A3(n18905), 
        .A4(n18933), .ZN(n18789) );
  AOI211_X1 U21786 ( .C1(n18785), .C2(n18929), .A(n18784), .B(n18789), .ZN(
        n18786) );
  OAI21_X1 U21787 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n18787), .A(n18786), 
        .ZN(P3_U2997) );
  OAI21_X1 U21788 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18788), .ZN(n18790) );
  AOI21_X1 U21789 ( .B1(n18791), .B2(n18790), .A(n18789), .ZN(P3_U2998) );
  AND2_X1 U21790 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18879), .ZN(
        P3_U2999) );
  AND2_X1 U21791 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18792), .ZN(
        P3_U3000) );
  AND2_X1 U21792 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18879), .ZN(
        P3_U3001) );
  AND2_X1 U21793 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18879), .ZN(
        P3_U3002) );
  AND2_X1 U21794 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18879), .ZN(
        P3_U3003) );
  AND2_X1 U21795 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18879), .ZN(
        P3_U3004) );
  AND2_X1 U21796 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18879), .ZN(
        P3_U3005) );
  AND2_X1 U21797 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18879), .ZN(
        P3_U3006) );
  AND2_X1 U21798 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18879), .ZN(
        P3_U3007) );
  AND2_X1 U21799 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18879), .ZN(
        P3_U3008) );
  AND2_X1 U21800 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18879), .ZN(
        P3_U3009) );
  AND2_X1 U21801 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18792), .ZN(
        P3_U3010) );
  AND2_X1 U21802 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18792), .ZN(
        P3_U3011) );
  AND2_X1 U21803 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18792), .ZN(
        P3_U3012) );
  AND2_X1 U21804 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18792), .ZN(
        P3_U3013) );
  AND2_X1 U21805 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18792), .ZN(
        P3_U3014) );
  AND2_X1 U21806 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18792), .ZN(
        P3_U3015) );
  AND2_X1 U21807 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18792), .ZN(
        P3_U3016) );
  AND2_X1 U21808 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18792), .ZN(
        P3_U3017) );
  AND2_X1 U21809 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18792), .ZN(
        P3_U3018) );
  AND2_X1 U21810 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18792), .ZN(
        P3_U3019) );
  AND2_X1 U21811 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18879), .ZN(
        P3_U3020) );
  AND2_X1 U21812 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18879), .ZN(P3_U3021) );
  AND2_X1 U21813 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18792), .ZN(P3_U3022) );
  AND2_X1 U21814 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18879), .ZN(P3_U3023) );
  AND2_X1 U21815 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18879), .ZN(P3_U3024) );
  AND2_X1 U21816 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18879), .ZN(P3_U3025) );
  AND2_X1 U21817 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18879), .ZN(P3_U3026) );
  AND2_X1 U21818 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18879), .ZN(P3_U3027) );
  AND2_X1 U21819 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18879), .ZN(P3_U3028) );
  INV_X1 U21820 ( .A(n18798), .ZN(n18797) );
  OAI21_X1 U21821 ( .B1(n18793), .B2(n21063), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18794) );
  AOI22_X1 U21822 ( .A1(n18807), .A2(n18809), .B1(n18941), .B2(n18794), .ZN(
        n18796) );
  NAND3_X1 U21823 ( .A1(NA), .A2(n18807), .A3(n18799), .ZN(n18795) );
  OAI211_X1 U21824 ( .C1(n18933), .C2(n18797), .A(n18796), .B(n18795), .ZN(
        P3_U3029) );
  NAND2_X1 U21825 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n18802) );
  AOI22_X1 U21826 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n18802), .B1(HOLD), 
        .B2(n18798), .ZN(n18800) );
  NOR2_X1 U21827 ( .A1(n18933), .A2(n18799), .ZN(n18801) );
  INV_X1 U21828 ( .A(n18801), .ZN(n18803) );
  OAI211_X1 U21829 ( .C1(n18800), .C2(n18807), .A(n18803), .B(n18930), .ZN(
        P3_U3030) );
  INV_X1 U21830 ( .A(NA), .ZN(n21031) );
  AOI221_X1 U21831 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n18807), .C1(n21031), 
        .C2(n18807), .A(n18801), .ZN(n18808) );
  INV_X1 U21832 ( .A(n18802), .ZN(n18805) );
  OAI22_X1 U21833 ( .A1(NA), .A2(n18803), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18804) );
  OAI22_X1 U21834 ( .A1(n18805), .A2(n18804), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18806) );
  OAI22_X1 U21835 ( .A1(n18808), .A2(n18809), .B1(n18807), .B2(n18806), .ZN(
        P3_U3031) );
  INV_X1 U21836 ( .A(n18941), .ZN(n18940) );
  OAI222_X1 U21837 ( .A1(n18811), .A2(n18873), .B1(n18810), .B2(n18940), .C1(
        n18812), .C2(n18862), .ZN(P3_U3032) );
  INV_X1 U21838 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18814) );
  OAI222_X1 U21839 ( .A1(n18862), .A2(n18814), .B1(n18813), .B2(n18870), .C1(
        n18812), .C2(n18873), .ZN(P3_U3033) );
  OAI222_X1 U21840 ( .A1(n18862), .A2(n18816), .B1(n18815), .B2(n18940), .C1(
        n18814), .C2(n18873), .ZN(P3_U3034) );
  OAI222_X1 U21841 ( .A1(n18862), .A2(n18818), .B1(n18817), .B2(n18870), .C1(
        n18816), .C2(n18873), .ZN(P3_U3035) );
  OAI222_X1 U21842 ( .A1(n18862), .A2(n18820), .B1(n18819), .B2(n18940), .C1(
        n18818), .C2(n18873), .ZN(P3_U3036) );
  OAI222_X1 U21843 ( .A1(n18862), .A2(n18822), .B1(n18821), .B2(n18940), .C1(
        n18820), .C2(n18873), .ZN(P3_U3037) );
  OAI222_X1 U21844 ( .A1(n18862), .A2(n18824), .B1(n18823), .B2(n18870), .C1(
        n18822), .C2(n18873), .ZN(P3_U3038) );
  OAI222_X1 U21845 ( .A1(n18862), .A2(n18826), .B1(n18825), .B2(n18940), .C1(
        n18824), .C2(n18873), .ZN(P3_U3039) );
  OAI222_X1 U21846 ( .A1(n18862), .A2(n18828), .B1(n18827), .B2(n18940), .C1(
        n18826), .C2(n18873), .ZN(P3_U3040) );
  OAI222_X1 U21847 ( .A1(n18862), .A2(n18830), .B1(n18829), .B2(n18940), .C1(
        n18828), .C2(n18873), .ZN(P3_U3041) );
  OAI222_X1 U21848 ( .A1(n18862), .A2(n18832), .B1(n18831), .B2(n18940), .C1(
        n18830), .C2(n18873), .ZN(P3_U3042) );
  OAI222_X1 U21849 ( .A1(n18862), .A2(n18834), .B1(n18833), .B2(n18940), .C1(
        n18832), .C2(n18873), .ZN(P3_U3043) );
  OAI222_X1 U21850 ( .A1(n18862), .A2(n18837), .B1(n18835), .B2(n18940), .C1(
        n18834), .C2(n18873), .ZN(P3_U3044) );
  OAI222_X1 U21851 ( .A1(n18837), .A2(n18873), .B1(n18836), .B2(n18940), .C1(
        n18838), .C2(n18862), .ZN(P3_U3045) );
  OAI222_X1 U21852 ( .A1(n18862), .A2(n18840), .B1(n18839), .B2(n18940), .C1(
        n18838), .C2(n18873), .ZN(P3_U3046) );
  OAI222_X1 U21853 ( .A1(n18862), .A2(n18843), .B1(n18841), .B2(n18940), .C1(
        n18840), .C2(n18873), .ZN(P3_U3047) );
  OAI222_X1 U21854 ( .A1(n18843), .A2(n18873), .B1(n18842), .B2(n18940), .C1(
        n18844), .C2(n18862), .ZN(P3_U3048) );
  OAI222_X1 U21855 ( .A1(n18862), .A2(n18846), .B1(n18845), .B2(n18940), .C1(
        n18844), .C2(n18873), .ZN(P3_U3049) );
  OAI222_X1 U21856 ( .A1(n18862), .A2(n18849), .B1(n18847), .B2(n18940), .C1(
        n18846), .C2(n18873), .ZN(P3_U3050) );
  OAI222_X1 U21857 ( .A1(n18849), .A2(n18873), .B1(n18848), .B2(n18940), .C1(
        n18850), .C2(n18862), .ZN(P3_U3051) );
  OAI222_X1 U21858 ( .A1(n18862), .A2(n18852), .B1(n18851), .B2(n18940), .C1(
        n18850), .C2(n18873), .ZN(P3_U3052) );
  OAI222_X1 U21859 ( .A1(n18862), .A2(n18854), .B1(n18853), .B2(n18940), .C1(
        n18852), .C2(n18873), .ZN(P3_U3053) );
  OAI222_X1 U21860 ( .A1(n18862), .A2(n18856), .B1(n18855), .B2(n18870), .C1(
        n18854), .C2(n18873), .ZN(P3_U3054) );
  INV_X1 U21861 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18858) );
  OAI222_X1 U21862 ( .A1(n18862), .A2(n18858), .B1(n18857), .B2(n18870), .C1(
        n18856), .C2(n18873), .ZN(P3_U3055) );
  OAI222_X1 U21863 ( .A1(n18862), .A2(n18860), .B1(n18859), .B2(n18870), .C1(
        n18858), .C2(n18873), .ZN(P3_U3056) );
  OAI222_X1 U21864 ( .A1(n18862), .A2(n18863), .B1(n18861), .B2(n18870), .C1(
        n18860), .C2(n18873), .ZN(P3_U3057) );
  OAI222_X1 U21865 ( .A1(n18862), .A2(n18866), .B1(n18864), .B2(n18870), .C1(
        n18863), .C2(n18873), .ZN(P3_U3058) );
  OAI222_X1 U21866 ( .A1(n18866), .A2(n18873), .B1(n18865), .B2(n18870), .C1(
        n18867), .C2(n18862), .ZN(P3_U3059) );
  OAI222_X1 U21867 ( .A1(n18862), .A2(n18872), .B1(n18868), .B2(n18870), .C1(
        n18867), .C2(n18873), .ZN(P3_U3060) );
  INV_X1 U21868 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18871) );
  OAI222_X1 U21869 ( .A1(n18873), .A2(n18872), .B1(n18871), .B2(n18870), .C1(
        n18869), .C2(n18862), .ZN(P3_U3061) );
  OAI22_X1 U21870 ( .A1(n18941), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18940), .ZN(n18874) );
  INV_X1 U21871 ( .A(n18874), .ZN(P3_U3274) );
  OAI22_X1 U21872 ( .A1(n18941), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18940), .ZN(n18875) );
  INV_X1 U21873 ( .A(n18875), .ZN(P3_U3275) );
  OAI22_X1 U21874 ( .A1(n18941), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18940), .ZN(n18876) );
  INV_X1 U21875 ( .A(n18876), .ZN(P3_U3276) );
  OAI22_X1 U21876 ( .A1(n18941), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18870), .ZN(n18877) );
  INV_X1 U21877 ( .A(n18877), .ZN(P3_U3277) );
  INV_X1 U21878 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18915) );
  AOI21_X1 U21879 ( .B1(n18879), .B2(n18915), .A(n18878), .ZN(P3_U3280) );
  AOI21_X1 U21880 ( .B1(n18879), .B2(P3_DATAWIDTH_REG_1__SCAN_IN), .A(n18878), 
        .ZN(n18880) );
  INV_X1 U21881 ( .A(n18880), .ZN(P3_U3281) );
  OAI221_X1 U21882 ( .B1(n18883), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18883), 
        .C2(n18882), .A(n18881), .ZN(P3_U3282) );
  NOR2_X1 U21883 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18892), .ZN(
        n18885) );
  AOI22_X1 U21884 ( .A1(n18909), .A2(n18886), .B1(n18885), .B2(n18884), .ZN(
        n18889) );
  AOI21_X1 U21885 ( .B1(n18902), .B2(n18887), .A(n18913), .ZN(n18888) );
  OAI22_X1 U21886 ( .A1(n18913), .A2(n18889), .B1(n18888), .B2(n12014), .ZN(
        P3_U3285) );
  NAND2_X1 U21887 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18908) );
  AOI22_X1 U21888 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18891), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n18890), .ZN(n18900) );
  OAI22_X1 U21889 ( .A1(n18893), .A2(n18892), .B1(n18908), .B2(n18900), .ZN(
        n18894) );
  AOI21_X1 U21890 ( .B1(n18909), .B2(n18895), .A(n18894), .ZN(n18896) );
  AOI22_X1 U21891 ( .A1(n18913), .A2(n18897), .B1(n18896), .B2(n18910), .ZN(
        P3_U3288) );
  INV_X1 U21892 ( .A(n18898), .ZN(n18901) );
  INV_X1 U21893 ( .A(n18908), .ZN(n18899) );
  AOI222_X1 U21894 ( .A1(n18903), .A2(n18902), .B1(n18909), .B2(n18901), .C1(
        n18900), .C2(n18899), .ZN(n18904) );
  AOI22_X1 U21895 ( .A1(n18913), .A2(n12023), .B1(n18904), .B2(n18910), .ZN(
        P3_U3289) );
  OAI21_X1 U21896 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18906), .A(n18905), 
        .ZN(n18907) );
  AOI22_X1 U21897 ( .A1(n18909), .A2(n18912), .B1(n18908), .B2(n18907), .ZN(
        n18911) );
  AOI22_X1 U21898 ( .A1(n18913), .A2(n18912), .B1(n18911), .B2(n18910), .ZN(
        P3_U3290) );
  NOR3_X1 U21899 ( .A1(n18915), .A2(P3_REIP_REG_0__SCAN_IN), .A3(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18914) );
  AOI221_X1 U21900 ( .B1(n18916), .B2(n18915), .C1(P3_REIP_REG_1__SCAN_IN), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n18914), .ZN(n18918) );
  INV_X1 U21901 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18917) );
  INV_X1 U21902 ( .A(n18922), .ZN(n18919) );
  AOI22_X1 U21903 ( .A1(n18922), .A2(n18918), .B1(n18917), .B2(n18919), .ZN(
        P3_U3292) );
  NOR2_X1 U21904 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n18921) );
  INV_X1 U21905 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18920) );
  AOI22_X1 U21906 ( .A1(n18922), .A2(n18921), .B1(n18920), .B2(n18919), .ZN(
        P3_U3293) );
  INV_X1 U21907 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18923) );
  AOI22_X1 U21908 ( .A1(n18940), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18923), 
        .B2(n18941), .ZN(P3_U3294) );
  MUX2_X1 U21909 ( .A(P3_MORE_REG_SCAN_IN), .B(n18925), .S(n18924), .Z(
        P3_U3295) );
  OAI21_X1 U21910 ( .B1(n18927), .B2(n18926), .A(n18946), .ZN(n18928) );
  AOI21_X1 U21911 ( .B1(n18929), .B2(n18933), .A(n18928), .ZN(n18939) );
  AOI21_X1 U21912 ( .B1(n18932), .B2(n18931), .A(n18930), .ZN(n18934) );
  OAI211_X1 U21913 ( .C1(n18945), .C2(n18934), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18933), .ZN(n18936) );
  AOI21_X1 U21914 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18936), .A(n18935), 
        .ZN(n18938) );
  NAND2_X1 U21915 ( .A1(n18939), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18937) );
  OAI21_X1 U21916 ( .B1(n18939), .B2(n18938), .A(n18937), .ZN(P3_U3296) );
  OAI22_X1 U21917 ( .A1(n18941), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18940), .ZN(n18942) );
  INV_X1 U21918 ( .A(n18942), .ZN(P3_U3297) );
  OR2_X1 U21919 ( .A1(n18944), .A2(n18943), .ZN(n18949) );
  OAI22_X1 U21920 ( .A1(n18949), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18946), 
        .B2(n18945), .ZN(n18947) );
  INV_X1 U21921 ( .A(n18947), .ZN(P3_U3298) );
  OAI21_X1 U21922 ( .B1(n18949), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n18948), 
        .ZN(n18950) );
  INV_X1 U21923 ( .A(n18950), .ZN(P3_U3299) );
  INV_X1 U21924 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19872) );
  NAND2_X1 U21925 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19872), .ZN(n19861) );
  INV_X1 U21926 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19854) );
  AOI22_X1 U21927 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19861), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n19854), .ZN(n19928) );
  AOI21_X1 U21928 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19928), .ZN(n18951) );
  INV_X1 U21929 ( .A(n18951), .ZN(P2_U2815) );
  INV_X1 U21930 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18953) );
  NAND2_X1 U21931 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18952), .ZN(n19846) );
  OAI22_X1 U21932 ( .A1(n19980), .A2(n18953), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19846), .ZN(P2_U2816) );
  INV_X1 U21933 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19864) );
  OR2_X1 U21934 ( .A1(n19864), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n19997) );
  AOI22_X1 U21935 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(n19997), .B1(n19863), .B2(
        n19854), .ZN(n18954) );
  OAI21_X1 U21936 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n19997), .A(n18954), 
        .ZN(P2_U2817) );
  OAI21_X1 U21937 ( .B1(n19863), .B2(BS16), .A(n19928), .ZN(n19926) );
  OAI21_X1 U21938 ( .B1(n19928), .B2(n19643), .A(n19926), .ZN(P2_U2818) );
  NOR4_X1 U21939 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18958) );
  NOR4_X1 U21940 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18957) );
  NOR4_X1 U21941 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18956) );
  NOR4_X1 U21942 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18955) );
  NAND4_X1 U21943 ( .A1(n18958), .A2(n18957), .A3(n18956), .A4(n18955), .ZN(
        n18964) );
  NOR4_X1 U21944 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18962) );
  AOI211_X1 U21945 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n18961) );
  NOR4_X1 U21946 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18960) );
  NOR4_X1 U21947 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18959) );
  NAND4_X1 U21948 ( .A1(n18962), .A2(n18961), .A3(n18960), .A4(n18959), .ZN(
        n18963) );
  NOR2_X1 U21949 ( .A1(n18964), .A2(n18963), .ZN(n18974) );
  INV_X1 U21950 ( .A(n18974), .ZN(n18972) );
  NOR2_X1 U21951 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18972), .ZN(n18967) );
  INV_X1 U21952 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18965) );
  AOI22_X1 U21953 ( .A1(n18967), .A2(n11457), .B1(n18972), .B2(n18965), .ZN(
        P2_U2820) );
  OR3_X1 U21954 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18971) );
  INV_X1 U21955 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18966) );
  AOI22_X1 U21956 ( .A1(n18967), .A2(n18971), .B1(n18972), .B2(n18966), .ZN(
        P2_U2821) );
  INV_X1 U21957 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19927) );
  NAND2_X1 U21958 ( .A1(n18967), .A2(n19927), .ZN(n18970) );
  OAI21_X1 U21959 ( .B1(n11445), .B2(n11457), .A(n18974), .ZN(n18968) );
  OAI21_X1 U21960 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18974), .A(n18968), 
        .ZN(n18969) );
  OAI221_X1 U21961 ( .B1(n18970), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18970), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18969), .ZN(P2_U2822) );
  INV_X1 U21962 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18973) );
  OAI221_X1 U21963 ( .B1(n18974), .B2(n18973), .C1(n18972), .C2(n18971), .A(
        n18970), .ZN(P2_U2823) );
  AOI22_X1 U21964 ( .A1(n19135), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n19076), .ZN(n18975) );
  OAI21_X1 U21965 ( .B1(n11846), .B2(n19073), .A(n18975), .ZN(n18978) );
  NOR2_X1 U21966 ( .A1(n18976), .A2(n19101), .ZN(n18977) );
  AOI211_X1 U21967 ( .C1(n19122), .C2(n18979), .A(n18978), .B(n18977), .ZN(
        n18986) );
  AOI211_X1 U21968 ( .C1(n18982), .C2(n18980), .A(n18981), .B(n19851), .ZN(
        n18983) );
  AOI21_X1 U21969 ( .B1(n19129), .B2(n18984), .A(n18983), .ZN(n18985) );
  NAND2_X1 U21970 ( .A1(n18986), .A2(n18985), .ZN(P2_U2834) );
  AOI22_X1 U21971 ( .A1(n18987), .A2(n19131), .B1(P2_REIP_REG_20__SCAN_IN), 
        .B2(n19076), .ZN(n18998) );
  AOI22_X1 U21972 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n19135), .B1(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19142), .ZN(n18997) );
  NOR2_X1 U21973 ( .A1(n18988), .A2(n19137), .ZN(n18989) );
  AOI21_X1 U21974 ( .B1(n18990), .B2(n19129), .A(n18989), .ZN(n18996) );
  AOI21_X1 U21975 ( .B1(n18993), .B2(n18991), .A(n18992), .ZN(n18994) );
  NAND2_X1 U21976 ( .A1(n19123), .A2(n18994), .ZN(n18995) );
  NAND4_X1 U21977 ( .A1(n18998), .A2(n18997), .A3(n18996), .A4(n18995), .ZN(
        P2_U2835) );
  AOI211_X1 U21978 ( .C1(n18999), .C2(n19001), .A(n19851), .B(n19000), .ZN(
        n19008) );
  AOI22_X1 U21979 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(n19135), .B1(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19142), .ZN(n19002) );
  OAI211_X1 U21980 ( .C1(n19133), .C2(n19895), .A(n19002), .B(n19113), .ZN(
        n19003) );
  AOI21_X1 U21981 ( .B1(n19004), .B2(n19122), .A(n19003), .ZN(n19005) );
  OAI21_X1 U21982 ( .B1(n19006), .B2(n19101), .A(n19005), .ZN(n19007) );
  NOR2_X1 U21983 ( .A1(n19008), .A2(n19007), .ZN(n19009) );
  OAI21_X1 U21984 ( .B1(n19010), .B2(n19127), .A(n19009), .ZN(P2_U2836) );
  INV_X1 U21985 ( .A(n19011), .ZN(n19023) );
  AOI22_X1 U21986 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(n19135), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n19142), .ZN(n19012) );
  OAI211_X1 U21987 ( .C1(n19133), .C2(n19892), .A(n19012), .B(n19113), .ZN(
        n19013) );
  INV_X1 U21988 ( .A(n19013), .ZN(n19014) );
  OAI21_X1 U21989 ( .B1(n19015), .B2(n19137), .A(n19014), .ZN(n19020) );
  AOI211_X1 U21990 ( .C1(n19018), .C2(n19017), .A(n19851), .B(n19016), .ZN(
        n19019) );
  AOI211_X1 U21991 ( .C1(n19131), .C2(n19021), .A(n19020), .B(n19019), .ZN(
        n19022) );
  OAI21_X1 U21992 ( .B1(n19023), .B2(n19127), .A(n19022), .ZN(P2_U2838) );
  INV_X1 U21993 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n19036) );
  OAI22_X1 U21994 ( .A1(n19025), .A2(n19101), .B1(n19073), .B2(n19024), .ZN(
        n19026) );
  AOI211_X1 U21995 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n19076), .A(n15544), 
        .B(n19026), .ZN(n19035) );
  NOR2_X1 U21996 ( .A1(n19105), .A2(n19027), .ZN(n19028) );
  XNOR2_X1 U21997 ( .A(n19029), .B(n19028), .ZN(n19033) );
  OAI22_X1 U21998 ( .A1(n19031), .A2(n19127), .B1(n19137), .B2(n19030), .ZN(
        n19032) );
  AOI21_X1 U21999 ( .B1(n19033), .B2(n19123), .A(n19032), .ZN(n19034) );
  OAI211_X1 U22000 ( .C1(n19100), .C2(n19036), .A(n19035), .B(n19034), .ZN(
        P2_U2839) );
  NOR2_X1 U22001 ( .A1(n19105), .A2(n19037), .ZN(n19039) );
  XOR2_X1 U22002 ( .A(n19039), .B(n19038), .Z(n19049) );
  AOI22_X1 U22003 ( .A1(n19040), .A2(n19131), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19142), .ZN(n19041) );
  OAI21_X1 U22004 ( .B1(n19100), .B2(n19042), .A(n19041), .ZN(n19043) );
  AOI211_X1 U22005 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19076), .A(n15544), 
        .B(n19043), .ZN(n19048) );
  INV_X1 U22006 ( .A(n19044), .ZN(n19045) );
  OAI22_X1 U22007 ( .A1(n19154), .A2(n19127), .B1(n19137), .B2(n19045), .ZN(
        n19046) );
  INV_X1 U22008 ( .A(n19046), .ZN(n19047) );
  OAI211_X1 U22009 ( .C1(n19851), .C2(n19049), .A(n19048), .B(n19047), .ZN(
        P2_U2841) );
  NAND2_X1 U22010 ( .A1(n12794), .A2(n19050), .ZN(n19052) );
  XOR2_X1 U22011 ( .A(n19052), .B(n19051), .Z(n19060) );
  AOI22_X1 U22012 ( .A1(n19053), .A2(n19131), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19142), .ZN(n19054) );
  OAI211_X1 U22013 ( .C1(n11895), .C2(n19133), .A(n19054), .B(n19113), .ZN(
        n19058) );
  OAI22_X1 U22014 ( .A1(n19056), .A2(n19127), .B1(n19137), .B2(n19055), .ZN(
        n19057) );
  AOI211_X1 U22015 ( .C1(P2_EBX_REG_13__SCAN_IN), .C2(n19135), .A(n19058), .B(
        n19057), .ZN(n19059) );
  OAI21_X1 U22016 ( .B1(n19060), .B2(n19851), .A(n19059), .ZN(P2_U2842) );
  NOR2_X1 U22017 ( .A1(n19105), .A2(n19071), .ZN(n19062) );
  XOR2_X1 U22018 ( .A(n19062), .B(n19061), .Z(n19070) );
  AOI22_X1 U22019 ( .A1(P2_EBX_REG_12__SCAN_IN), .A2(n19135), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19142), .ZN(n19063) );
  OAI21_X1 U22020 ( .B1(n19064), .B2(n19101), .A(n19063), .ZN(n19065) );
  AOI211_X1 U22021 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19076), .A(n15544), 
        .B(n19065), .ZN(n19069) );
  AOI22_X1 U22022 ( .A1(n19067), .A2(n19122), .B1(n19129), .B2(n19066), .ZN(
        n19068) );
  OAI211_X1 U22023 ( .C1(n19851), .C2(n19070), .A(n19069), .B(n19068), .ZN(
        P2_U2843) );
  AOI211_X1 U22024 ( .C1(n19084), .C2(n19072), .A(n19071), .B(n19145), .ZN(
        n19083) );
  OAI22_X1 U22025 ( .A1(n19100), .A2(n11705), .B1(n19074), .B2(n19073), .ZN(
        n19075) );
  AOI211_X1 U22026 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n19076), .A(n15544), 
        .B(n19075), .ZN(n19077) );
  OAI21_X1 U22027 ( .B1(n19078), .B2(n19127), .A(n19077), .ZN(n19081) );
  NOR2_X1 U22028 ( .A1(n19079), .A2(n19101), .ZN(n19080) );
  OR2_X1 U22029 ( .A1(n19081), .A2(n19080), .ZN(n19082) );
  NOR2_X1 U22030 ( .A1(n19083), .A2(n19082), .ZN(n19086) );
  AOI22_X1 U22031 ( .A1(n10163), .A2(n19122), .B1(n19141), .B2(n19084), .ZN(
        n19085) );
  NAND2_X1 U22032 ( .A1(n19086), .A2(n19085), .ZN(P2_U2844) );
  NAND2_X1 U22033 ( .A1(n12794), .A2(n19087), .ZN(n19089) );
  XOR2_X1 U22034 ( .A(n19089), .B(n19088), .Z(n19097) );
  AOI22_X1 U22035 ( .A1(n19090), .A2(n19131), .B1(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19142), .ZN(n19091) );
  OAI211_X1 U22036 ( .C1(n11879), .C2(n19133), .A(n19091), .B(n19113), .ZN(
        n19095) );
  OAI22_X1 U22037 ( .A1(n19093), .A2(n19127), .B1(n19137), .B2(n19092), .ZN(
        n19094) );
  AOI211_X1 U22038 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n19135), .A(n19095), .B(
        n19094), .ZN(n19096) );
  OAI21_X1 U22039 ( .B1(n19097), .B2(n19851), .A(n19096), .ZN(P2_U2846) );
  OAI21_X1 U22040 ( .B1(n11869), .B2(n19133), .A(n19113), .ZN(n19103) );
  OAI22_X1 U22041 ( .A1(n9809), .A2(n19101), .B1(n19100), .B2(n19099), .ZN(
        n19102) );
  AOI211_X1 U22042 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19142), .A(
        n19103), .B(n19102), .ZN(n19111) );
  NOR2_X1 U22043 ( .A1(n19105), .A2(n19104), .ZN(n19107) );
  XNOR2_X1 U22044 ( .A(n19107), .B(n19106), .ZN(n19109) );
  AOI22_X1 U22045 ( .A1(n19109), .A2(n19123), .B1(n19122), .B2(n19108), .ZN(
        n19110) );
  OAI211_X1 U22046 ( .C1(n19127), .C2(n19112), .A(n19111), .B(n19110), .ZN(
        P2_U2849) );
  OAI21_X1 U22047 ( .B1(n11864), .B2(n19133), .A(n19113), .ZN(n19117) );
  AOI22_X1 U22048 ( .A1(n19114), .A2(n19131), .B1(P2_EBX_REG_5__SCAN_IN), .B2(
        n19135), .ZN(n19115) );
  INV_X1 U22049 ( .A(n19115), .ZN(n19116) );
  AOI211_X1 U22050 ( .C1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n19142), .A(
        n19117), .B(n19116), .ZN(n19126) );
  NAND2_X1 U22051 ( .A1(n12794), .A2(n19118), .ZN(n19119) );
  XNOR2_X1 U22052 ( .A(n19120), .B(n19119), .ZN(n19124) );
  AOI22_X1 U22053 ( .A1(n19124), .A2(n19123), .B1(n19122), .B2(n19121), .ZN(
        n19125) );
  OAI211_X1 U22054 ( .C1(n19127), .C2(n19173), .A(n19126), .B(n19125), .ZN(
        P2_U2850) );
  INV_X1 U22055 ( .A(n19128), .ZN(n19193) );
  AOI22_X1 U22056 ( .A1(n19131), .A2(n19130), .B1(n19129), .B2(n19193), .ZN(
        n19132) );
  OAI21_X1 U22057 ( .B1(n11457), .B2(n19133), .A(n19132), .ZN(n19134) );
  AOI21_X1 U22058 ( .B1(n19135), .B2(P2_EBX_REG_0__SCAN_IN), .A(n19134), .ZN(
        n19136) );
  OAI21_X1 U22059 ( .B1(n19138), .B2(n19137), .A(n19136), .ZN(n19139) );
  AOI21_X1 U22060 ( .B1(n19297), .B2(n19140), .A(n19139), .ZN(n19144) );
  OAI21_X1 U22061 ( .B1(n19142), .B2(n19141), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19143) );
  OAI211_X1 U22062 ( .C1(n19146), .C2(n19145), .A(n19144), .B(n19143), .ZN(
        P2_U2855) );
  AOI22_X1 U22063 ( .A1(n19148), .A2(n19189), .B1(n19147), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19151) );
  AOI22_X1 U22064 ( .A1(n19149), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19188), .ZN(n19150) );
  NAND2_X1 U22065 ( .A1(n19151), .A2(n19150), .ZN(P2_U2888) );
  AOI22_X1 U22066 ( .A1(n19167), .A2(n19152), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19188), .ZN(n19153) );
  OAI21_X1 U22067 ( .B1(n19174), .B2(n19154), .A(n19153), .ZN(P2_U2905) );
  AOI22_X1 U22068 ( .A1(n19167), .A2(n19155), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n19188), .ZN(n19156) );
  OAI21_X1 U22069 ( .B1(n19174), .B2(n19157), .A(n19156), .ZN(P2_U2907) );
  INV_X1 U22070 ( .A(n19158), .ZN(n19161) );
  AOI22_X1 U22071 ( .A1(n19167), .A2(n19159), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n19188), .ZN(n19160) );
  OAI21_X1 U22072 ( .B1(n19174), .B2(n19161), .A(n19160), .ZN(P2_U2909) );
  INV_X1 U22073 ( .A(n19162), .ZN(n19165) );
  AOI22_X1 U22074 ( .A1(n19167), .A2(n19163), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n19188), .ZN(n19164) );
  OAI21_X1 U22075 ( .B1(n19174), .B2(n19165), .A(n19164), .ZN(P2_U2911) );
  INV_X1 U22076 ( .A(n19276), .ZN(n19166) );
  AOI22_X1 U22077 ( .A1(n19167), .A2(n19166), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19188), .ZN(n19172) );
  INV_X1 U22078 ( .A(n19168), .ZN(n19169) );
  NAND3_X1 U22079 ( .A1(n19170), .A2(n19169), .A3(n19191), .ZN(n19171) );
  OAI211_X1 U22080 ( .C1(n19174), .C2(n19173), .A(n19172), .B(n19171), .ZN(
        P2_U2914) );
  AOI22_X1 U22081 ( .A1(n19936), .A2(n19189), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19188), .ZN(n19180) );
  AOI21_X1 U22082 ( .B1(n19177), .B2(n19176), .A(n19175), .ZN(n19178) );
  OR2_X1 U22083 ( .A1(n19178), .A2(n19183), .ZN(n19179) );
  OAI211_X1 U22084 ( .C1(n19266), .C2(n19196), .A(n19180), .B(n19179), .ZN(
        P2_U2916) );
  AOI22_X1 U22085 ( .A1(n19189), .A2(n19954), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19188), .ZN(n19186) );
  AOI21_X1 U22086 ( .B1(n19190), .B2(n19182), .A(n19181), .ZN(n19184) );
  OR2_X1 U22087 ( .A1(n19184), .A2(n19183), .ZN(n19185) );
  OAI211_X1 U22088 ( .C1(n19187), .C2(n19196), .A(n19186), .B(n19185), .ZN(
        P2_U2918) );
  AOI22_X1 U22089 ( .A1(n19189), .A2(n19193), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19188), .ZN(n19195) );
  INV_X1 U22090 ( .A(n19190), .ZN(n19192) );
  OAI211_X1 U22091 ( .C1(n19297), .C2(n19193), .A(n19192), .B(n19191), .ZN(
        n19194) );
  OAI211_X1 U22092 ( .C1(n19248), .C2(n19196), .A(n19195), .B(n19194), .ZN(
        P2_U2919) );
  AND2_X1 U22093 ( .A1(n19211), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22094 ( .A1(n19982), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19198) );
  OAI21_X1 U22095 ( .B1(n12966), .B2(n19230), .A(n19198), .ZN(P2_U2936) );
  AOI22_X1 U22096 ( .A1(n19982), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19199) );
  OAI21_X1 U22097 ( .B1(n19200), .B2(n19230), .A(n19199), .ZN(P2_U2937) );
  AOI22_X1 U22098 ( .A1(n19982), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19201) );
  OAI21_X1 U22099 ( .B1(n19202), .B2(n19230), .A(n19201), .ZN(P2_U2938) );
  AOI22_X1 U22100 ( .A1(n19982), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19203) );
  OAI21_X1 U22101 ( .B1(n19204), .B2(n19230), .A(n19203), .ZN(P2_U2939) );
  AOI22_X1 U22102 ( .A1(n19982), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19205) );
  OAI21_X1 U22103 ( .B1(n19206), .B2(n19230), .A(n19205), .ZN(P2_U2940) );
  AOI22_X1 U22104 ( .A1(n19982), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19207) );
  OAI21_X1 U22105 ( .B1(n19208), .B2(n19230), .A(n19207), .ZN(P2_U2941) );
  AOI22_X1 U22106 ( .A1(n19982), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19209) );
  OAI21_X1 U22107 ( .B1(n19210), .B2(n19230), .A(n19209), .ZN(P2_U2942) );
  AOI22_X1 U22108 ( .A1(n19982), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19211), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19212) );
  OAI21_X1 U22109 ( .B1(n19213), .B2(n19230), .A(n19212), .ZN(P2_U2943) );
  AOI22_X1 U22110 ( .A1(n19982), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19214) );
  OAI21_X1 U22111 ( .B1(n19215), .B2(n19230), .A(n19214), .ZN(P2_U2944) );
  AOI22_X1 U22112 ( .A1(n19982), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19216) );
  OAI21_X1 U22113 ( .B1(n19217), .B2(n19230), .A(n19216), .ZN(P2_U2945) );
  INV_X1 U22114 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19219) );
  AOI22_X1 U22115 ( .A1(n19982), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19218) );
  OAI21_X1 U22116 ( .B1(n19219), .B2(n19230), .A(n19218), .ZN(P2_U2946) );
  INV_X1 U22117 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19221) );
  AOI22_X1 U22118 ( .A1(n19982), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19220) );
  OAI21_X1 U22119 ( .B1(n19221), .B2(n19230), .A(n19220), .ZN(P2_U2947) );
  INV_X1 U22120 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19223) );
  AOI22_X1 U22121 ( .A1(n19982), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19222) );
  OAI21_X1 U22122 ( .B1(n19223), .B2(n19230), .A(n19222), .ZN(P2_U2948) );
  INV_X1 U22123 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19225) );
  AOI22_X1 U22124 ( .A1(n19982), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19224) );
  OAI21_X1 U22125 ( .B1(n19225), .B2(n19230), .A(n19224), .ZN(P2_U2949) );
  INV_X1 U22126 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19227) );
  AOI22_X1 U22127 ( .A1(n19982), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19226) );
  OAI21_X1 U22128 ( .B1(n19227), .B2(n19230), .A(n19226), .ZN(P2_U2950) );
  AOI22_X1 U22129 ( .A1(n19982), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19228), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19229) );
  OAI21_X1 U22130 ( .B1(n13020), .B2(n19230), .A(n19229), .ZN(P2_U2951) );
  AOI22_X1 U22131 ( .A1(n19231), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n11988), .ZN(n19238) );
  OAI22_X1 U22132 ( .A1(n19233), .A2(n11993), .B1(n13736), .B2(n19232), .ZN(
        n19234) );
  AOI21_X1 U22133 ( .B1(n19236), .B2(n19235), .A(n19234), .ZN(n19237) );
  OAI211_X1 U22134 ( .C1(n19240), .C2(n19239), .A(n19238), .B(n19237), .ZN(
        P2_U3010) );
  INV_X1 U22135 ( .A(n19330), .ZN(n19241) );
  AOI21_X1 U22136 ( .B1(n19842), .B2(n19241), .A(n19643), .ZN(n19242) );
  NOR2_X1 U22137 ( .A1(n19242), .A2(n19719), .ZN(n19249) );
  INV_X1 U22138 ( .A(n19243), .ZN(n19244) );
  AND2_X1 U22139 ( .A1(n19244), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19783) );
  NAND2_X1 U22140 ( .A1(n19938), .A2(n19946), .ZN(n19365) );
  INV_X1 U22141 ( .A(n19365), .ZN(n19363) );
  NAND2_X1 U22142 ( .A1(n19363), .A2(n19956), .ZN(n19303) );
  NOR2_X1 U22143 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19303), .ZN(
        n19289) );
  NOR2_X1 U22144 ( .A1(n19783), .A2(n19289), .ZN(n19252) );
  AOI21_X1 U22145 ( .B1(n19245), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19246) );
  OAI21_X1 U22146 ( .B1(n19246), .B2(n19289), .A(n19781), .ZN(n19247) );
  AOI22_X1 U22147 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19292), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19291), .ZN(n19787) );
  INV_X1 U22148 ( .A(n19274), .ZN(n19287) );
  AND2_X1 U22149 ( .A1(n11388), .A2(n19287), .ZN(n19716) );
  AOI22_X1 U22150 ( .A1(n19682), .A2(n19820), .B1(n19716), .B2(n19289), .ZN(
        n19255) );
  NOR2_X2 U22151 ( .A1(n19248), .A2(n19466), .ZN(n19727) );
  INV_X1 U22152 ( .A(n19249), .ZN(n19253) );
  OAI21_X1 U22153 ( .B1(n19250), .B2(n19289), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19251) );
  AOI22_X1 U22154 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19292), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19291), .ZN(n19623) );
  AOI22_X1 U22155 ( .A1(n19727), .A2(n19293), .B1(n19330), .B2(n19784), .ZN(
        n19254) );
  OAI211_X1 U22156 ( .C1(n19296), .C2(n19256), .A(n19255), .B(n19254), .ZN(
        P2_U3048) );
  AOI22_X1 U22157 ( .A1(n19731), .A2(n19820), .B1(n19730), .B2(n19289), .ZN(
        n19258) );
  AOI22_X1 U22158 ( .A1(n19732), .A2(n19293), .B1(n19330), .B2(n19791), .ZN(
        n19257) );
  OAI211_X1 U22159 ( .C1(n19296), .C2(n19259), .A(n19258), .B(n19257), .ZN(
        P2_U3049) );
  INV_X1 U22160 ( .A(n19291), .ZN(n19281) );
  INV_X1 U22161 ( .A(n19292), .ZN(n19283) );
  OAI22_X2 U22162 ( .A1(n19260), .A2(n19281), .B1(n20262), .B2(n19283), .ZN(
        n19798) );
  NOR2_X2 U22163 ( .A1(n11413), .A2(n19274), .ZN(n19736) );
  AOI22_X1 U22164 ( .A1(n19798), .A2(n19820), .B1(n19736), .B2(n19289), .ZN(
        n19263) );
  NOR2_X2 U22165 ( .A1(n19261), .A2(n19466), .ZN(n19737) );
  AOI22_X2 U22166 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19292), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19291), .ZN(n19801) );
  INV_X1 U22167 ( .A(n19801), .ZN(n19381) );
  AOI22_X1 U22168 ( .A1(n19737), .A2(n19293), .B1(n19330), .B2(n19381), .ZN(
        n19262) );
  OAI211_X1 U22169 ( .C1(n19296), .C2(n19264), .A(n19263), .B(n19262), .ZN(
        P2_U3050) );
  AOI22_X1 U22170 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19292), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19291), .ZN(n19694) );
  AND2_X1 U22171 ( .A1(n19265), .A2(n19287), .ZN(n19740) );
  AOI22_X1 U22172 ( .A1(n19805), .A2(n19820), .B1(n19740), .B2(n19289), .ZN(
        n19268) );
  NOR2_X2 U22173 ( .A1(n19266), .A2(n19466), .ZN(n19741) );
  AOI22_X1 U22174 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19292), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19291), .ZN(n19808) );
  INV_X1 U22175 ( .A(n19808), .ZN(n19691) );
  AOI22_X1 U22176 ( .A1(n19741), .A2(n19293), .B1(n19330), .B2(n19691), .ZN(
        n19267) );
  OAI211_X1 U22177 ( .C1(n19296), .C2(n19269), .A(n19268), .B(n19267), .ZN(
        P2_U3051) );
  AOI22_X1 U22178 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19292), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19291), .ZN(n19699) );
  NOR2_X2 U22179 ( .A1(n11390), .A2(n19274), .ZN(n19744) );
  AOI22_X1 U22180 ( .A1(n19812), .A2(n19820), .B1(n19744), .B2(n19289), .ZN(
        n19272) );
  NOR2_X2 U22181 ( .A1(n19270), .A2(n19466), .ZN(n19746) );
  AOI22_X1 U22182 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19292), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19291), .ZN(n19815) );
  INV_X1 U22183 ( .A(n19815), .ZN(n19696) );
  AOI22_X1 U22184 ( .A1(n19746), .A2(n19293), .B1(n19330), .B2(n19696), .ZN(
        n19271) );
  OAI211_X1 U22185 ( .C1(n19296), .C2(n19273), .A(n19272), .B(n19271), .ZN(
        P2_U3052) );
  AOI22_X2 U22186 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19291), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19292), .ZN(n19824) );
  INV_X1 U22187 ( .A(n19824), .ZN(n19669) );
  NOR2_X2 U22188 ( .A1(n19275), .A2(n19274), .ZN(n19749) );
  AOI22_X1 U22189 ( .A1(n19669), .A2(n19820), .B1(n19749), .B2(n19289), .ZN(
        n19278) );
  NOR2_X2 U22190 ( .A1(n19276), .A2(n19466), .ZN(n19750) );
  AOI22_X1 U22191 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19292), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19291), .ZN(n19672) );
  AOI22_X1 U22192 ( .A1(n19750), .A2(n19293), .B1(n19330), .B2(n19819), .ZN(
        n19277) );
  OAI211_X1 U22193 ( .C1(n19296), .C2(n13216), .A(n19278), .B(n19277), .ZN(
        P2_U3053) );
  AOI22_X1 U22194 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19291), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19292), .ZN(n19758) );
  INV_X1 U22195 ( .A(n19758), .ZN(n19828) );
  AND2_X1 U22196 ( .A1(n19279), .A2(n19287), .ZN(n19753) );
  AOI22_X1 U22197 ( .A1(n19828), .A2(n19820), .B1(n19753), .B2(n19289), .ZN(
        n19285) );
  NOR2_X2 U22198 ( .A1(n19280), .A2(n19466), .ZN(n19755) );
  AOI22_X1 U22199 ( .A1(n19755), .A2(n19293), .B1(n19330), .B2(n19754), .ZN(
        n19284) );
  OAI211_X1 U22200 ( .C1(n19296), .C2(n19286), .A(n19285), .B(n19284), .ZN(
        P2_U3054) );
  AOI22_X1 U22201 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19292), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19291), .ZN(n19768) );
  AND2_X1 U22202 ( .A1(n19288), .A2(n19287), .ZN(n19760) );
  AOI22_X1 U22203 ( .A1(n19837), .A2(n19820), .B1(n19760), .B2(n19289), .ZN(
        n19295) );
  NOR2_X2 U22204 ( .A1(n19290), .A2(n19466), .ZN(n19763) );
  INV_X1 U22205 ( .A(n19843), .ZN(n19761) );
  AOI22_X1 U22206 ( .A1(n19763), .A2(n19293), .B1(n19330), .B2(n19761), .ZN(
        n19294) );
  OAI211_X1 U22207 ( .C1(n19296), .C2(n14302), .A(n19295), .B(n19294), .ZN(
        P2_U3055) );
  NAND2_X1 U22208 ( .A1(n19956), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19549) );
  NOR2_X1 U22209 ( .A1(n19549), .A2(n19365), .ZN(n19306) );
  OR2_X1 U22210 ( .A1(n19306), .A2(n19769), .ZN(n19298) );
  NOR2_X1 U22211 ( .A1(n11568), .A2(n19298), .ZN(n19302) );
  OAI21_X1 U22212 ( .B1(n19303), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19769), 
        .ZN(n19299) );
  INV_X1 U22213 ( .A(n19299), .ZN(n19300) );
  INV_X1 U22214 ( .A(n19727), .ZN(n19775) );
  INV_X1 U22215 ( .A(n19716), .ZN(n19774) );
  INV_X1 U22216 ( .A(n19306), .ZN(n19327) );
  OAI22_X1 U22217 ( .A1(n19328), .A2(n19775), .B1(n19774), .B2(n19327), .ZN(
        n19301) );
  INV_X1 U22218 ( .A(n19301), .ZN(n19308) );
  NAND2_X1 U22219 ( .A1(n19932), .A2(n19941), .ZN(n19304) );
  AOI21_X1 U22220 ( .B1(n19304), .B2(n19303), .A(n19302), .ZN(n19305) );
  OAI211_X1 U22221 ( .C1(n19306), .C2(n19645), .A(n19305), .B(n19781), .ZN(
        n19331) );
  AOI22_X1 U22222 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19331), .B1(
        n19330), .B2(n19682), .ZN(n19307) );
  OAI211_X1 U22223 ( .C1(n19623), .C2(n19356), .A(n19308), .B(n19307), .ZN(
        P2_U3056) );
  INV_X1 U22224 ( .A(n19732), .ZN(n19789) );
  OAI22_X1 U22225 ( .A1(n19328), .A2(n19789), .B1(n19788), .B2(n19327), .ZN(
        n19309) );
  INV_X1 U22226 ( .A(n19309), .ZN(n19311) );
  AOI22_X1 U22227 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19331), .B1(
        n19330), .B2(n19731), .ZN(n19310) );
  OAI211_X1 U22228 ( .C1(n19735), .C2(n19356), .A(n19311), .B(n19310), .ZN(
        P2_U3057) );
  INV_X1 U22229 ( .A(n19737), .ZN(n19796) );
  INV_X1 U22230 ( .A(n19736), .ZN(n19795) );
  OAI22_X1 U22231 ( .A1(n19328), .A2(n19796), .B1(n19795), .B2(n19327), .ZN(
        n19312) );
  INV_X1 U22232 ( .A(n19312), .ZN(n19314) );
  AOI22_X1 U22233 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19331), .B1(
        n19330), .B2(n19798), .ZN(n19313) );
  OAI211_X1 U22234 ( .C1(n19801), .C2(n19356), .A(n19314), .B(n19313), .ZN(
        P2_U3058) );
  INV_X1 U22235 ( .A(n19741), .ZN(n19803) );
  INV_X1 U22236 ( .A(n19740), .ZN(n19802) );
  OAI22_X1 U22237 ( .A1(n19328), .A2(n19803), .B1(n19802), .B2(n19327), .ZN(
        n19315) );
  INV_X1 U22238 ( .A(n19315), .ZN(n19317) );
  AOI22_X1 U22239 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19331), .B1(
        n19330), .B2(n19805), .ZN(n19316) );
  OAI211_X1 U22240 ( .C1(n19808), .C2(n19356), .A(n19317), .B(n19316), .ZN(
        P2_U3059) );
  INV_X1 U22241 ( .A(n19746), .ZN(n19810) );
  INV_X1 U22242 ( .A(n19744), .ZN(n19809) );
  OAI22_X1 U22243 ( .A1(n19328), .A2(n19810), .B1(n19809), .B2(n19327), .ZN(
        n19318) );
  INV_X1 U22244 ( .A(n19318), .ZN(n19320) );
  AOI22_X1 U22245 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19331), .B1(
        n19330), .B2(n19812), .ZN(n19319) );
  OAI211_X1 U22246 ( .C1(n19815), .C2(n19356), .A(n19320), .B(n19319), .ZN(
        P2_U3060) );
  INV_X1 U22247 ( .A(n19750), .ZN(n19817) );
  INV_X1 U22248 ( .A(n19749), .ZN(n19816) );
  OAI22_X1 U22249 ( .A1(n19328), .A2(n19817), .B1(n19816), .B2(n19327), .ZN(
        n19321) );
  INV_X1 U22250 ( .A(n19321), .ZN(n19323) );
  AOI22_X1 U22251 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19331), .B1(
        n19330), .B2(n19669), .ZN(n19322) );
  OAI211_X1 U22252 ( .C1(n19672), .C2(n19356), .A(n19323), .B(n19322), .ZN(
        P2_U3061) );
  INV_X1 U22253 ( .A(n19754), .ZN(n19831) );
  INV_X1 U22254 ( .A(n19755), .ZN(n19826) );
  INV_X1 U22255 ( .A(n19753), .ZN(n19825) );
  OAI22_X1 U22256 ( .A1(n19328), .A2(n19826), .B1(n19825), .B2(n19327), .ZN(
        n19324) );
  INV_X1 U22257 ( .A(n19324), .ZN(n19326) );
  AOI22_X1 U22258 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19331), .B1(
        n19330), .B2(n19828), .ZN(n19325) );
  OAI211_X1 U22259 ( .C1(n19831), .C2(n19356), .A(n19326), .B(n19325), .ZN(
        P2_U3062) );
  INV_X1 U22260 ( .A(n19763), .ZN(n19834) );
  INV_X1 U22261 ( .A(n19760), .ZN(n19833) );
  OAI22_X1 U22262 ( .A1(n19328), .A2(n19834), .B1(n19833), .B2(n19327), .ZN(
        n19329) );
  INV_X1 U22263 ( .A(n19329), .ZN(n19333) );
  AOI22_X1 U22264 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19331), .B1(
        n19330), .B2(n19837), .ZN(n19332) );
  OAI211_X1 U22265 ( .C1(n19843), .C2(n19356), .A(n19333), .B(n19332), .ZN(
        P2_U3063) );
  NOR2_X1 U22266 ( .A1(n19956), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19578) );
  AND2_X1 U22267 ( .A1(n19578), .A2(n19363), .ZN(n19357) );
  OAI21_X1 U22268 ( .B1(n19338), .B2(n19357), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19335) );
  NOR2_X1 U22269 ( .A1(n19580), .A2(n19365), .ZN(n19336) );
  INV_X1 U22270 ( .A(n19336), .ZN(n19334) );
  NAND2_X1 U22271 ( .A1(n19335), .A2(n19334), .ZN(n19358) );
  AOI22_X1 U22272 ( .A1(n19358), .A2(n19727), .B1(n19716), .B2(n19357), .ZN(
        n19343) );
  NAND2_X1 U22273 ( .A1(n19400), .A2(n19356), .ZN(n19337) );
  AOI21_X1 U22274 ( .B1(n19337), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19336), 
        .ZN(n19340) );
  AOI21_X1 U22275 ( .B1(n19338), .B2(n19645), .A(n19357), .ZN(n19339) );
  MUX2_X1 U22276 ( .A(n19340), .B(n19339), .S(n19719), .Z(n19341) );
  AOI22_X1 U22277 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19360), .B1(
        n19388), .B2(n19784), .ZN(n19342) );
  OAI211_X1 U22278 ( .C1(n19787), .C2(n19356), .A(n19343), .B(n19342), .ZN(
        P2_U3064) );
  AOI22_X1 U22279 ( .A1(n19358), .A2(n19732), .B1(n19730), .B2(n19357), .ZN(
        n19345) );
  AOI22_X1 U22280 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19360), .B1(
        n19388), .B2(n19791), .ZN(n19344) );
  OAI211_X1 U22281 ( .C1(n19794), .C2(n19356), .A(n19345), .B(n19344), .ZN(
        P2_U3065) );
  AOI22_X1 U22282 ( .A1(n19358), .A2(n19737), .B1(n19736), .B2(n19357), .ZN(
        n19347) );
  INV_X1 U22283 ( .A(n19356), .ZN(n19359) );
  AOI22_X1 U22284 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19360), .B1(
        n19359), .B2(n19798), .ZN(n19346) );
  OAI211_X1 U22285 ( .C1(n19801), .C2(n19400), .A(n19347), .B(n19346), .ZN(
        P2_U3066) );
  AOI22_X1 U22286 ( .A1(n19358), .A2(n19741), .B1(n19740), .B2(n19357), .ZN(
        n19349) );
  AOI22_X1 U22287 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19360), .B1(
        n19359), .B2(n19805), .ZN(n19348) );
  OAI211_X1 U22288 ( .C1(n19808), .C2(n19400), .A(n19349), .B(n19348), .ZN(
        P2_U3067) );
  AOI22_X1 U22289 ( .A1(n19358), .A2(n19746), .B1(n19744), .B2(n19357), .ZN(
        n19351) );
  AOI22_X1 U22290 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19360), .B1(
        n19359), .B2(n19812), .ZN(n19350) );
  OAI211_X1 U22291 ( .C1(n19815), .C2(n19400), .A(n19351), .B(n19350), .ZN(
        P2_U3068) );
  AOI22_X1 U22292 ( .A1(n19358), .A2(n19750), .B1(n19749), .B2(n19357), .ZN(
        n19353) );
  AOI22_X1 U22293 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19360), .B1(
        n19388), .B2(n19819), .ZN(n19352) );
  OAI211_X1 U22294 ( .C1(n19824), .C2(n19356), .A(n19353), .B(n19352), .ZN(
        P2_U3069) );
  AOI22_X1 U22295 ( .A1(n19358), .A2(n19755), .B1(n19753), .B2(n19357), .ZN(
        n19355) );
  AOI22_X1 U22296 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19360), .B1(
        n19388), .B2(n19754), .ZN(n19354) );
  OAI211_X1 U22297 ( .C1(n19758), .C2(n19356), .A(n19355), .B(n19354), .ZN(
        P2_U3070) );
  AOI22_X1 U22298 ( .A1(n19358), .A2(n19763), .B1(n19760), .B2(n19357), .ZN(
        n19362) );
  AOI22_X1 U22299 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19360), .B1(
        n19359), .B2(n19837), .ZN(n19361) );
  OAI211_X1 U22300 ( .C1(n19843), .C2(n19400), .A(n19362), .B(n19361), .ZN(
        P2_U3071) );
  NAND2_X1 U22301 ( .A1(n19932), .A2(n19619), .ZN(n19364) );
  NAND2_X1 U22302 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19363), .ZN(
        n19371) );
  NAND2_X1 U22303 ( .A1(n19364), .A2(n19371), .ZN(n19369) );
  NAND2_X1 U22304 ( .A1(n11566), .A2(n19645), .ZN(n19367) );
  NOR2_X1 U22305 ( .A1(n19609), .A2(n19365), .ZN(n19395) );
  INV_X1 U22306 ( .A(n19395), .ZN(n19366) );
  NAND2_X1 U22307 ( .A1(n19367), .A2(n19366), .ZN(n19368) );
  MUX2_X1 U22308 ( .A(n19369), .B(n19368), .S(n19719), .Z(n19370) );
  NAND2_X1 U22309 ( .A1(n19370), .A2(n19781), .ZN(n19397) );
  INV_X1 U22310 ( .A(n19397), .ZN(n19385) );
  INV_X1 U22311 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n19377) );
  AOI22_X1 U22312 ( .A1(n19784), .A2(n19431), .B1(n19395), .B2(n19716), .ZN(
        n19376) );
  INV_X1 U22313 ( .A(n19371), .ZN(n19372) );
  NAND2_X1 U22314 ( .A1(n19372), .A2(n19939), .ZN(n19374) );
  OAI21_X1 U22315 ( .B1(n11566), .B2(n19395), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19373) );
  NAND2_X1 U22316 ( .A1(n19374), .A2(n19373), .ZN(n19396) );
  AOI22_X1 U22317 ( .A1(n19727), .A2(n19396), .B1(n19388), .B2(n19682), .ZN(
        n19375) );
  OAI211_X1 U22318 ( .C1(n19385), .C2(n19377), .A(n19376), .B(n19375), .ZN(
        P2_U3072) );
  INV_X1 U22319 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n19380) );
  AOI22_X1 U22320 ( .A1(n19791), .A2(n19431), .B1(n19395), .B2(n19730), .ZN(
        n19379) );
  AOI22_X1 U22321 ( .A1(n19732), .A2(n19396), .B1(n19388), .B2(n19731), .ZN(
        n19378) );
  OAI211_X1 U22322 ( .C1(n19385), .C2(n19380), .A(n19379), .B(n19378), .ZN(
        P2_U3073) );
  INV_X1 U22323 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n19384) );
  AOI22_X1 U22324 ( .A1(n19381), .A2(n19431), .B1(n19395), .B2(n19736), .ZN(
        n19383) );
  AOI22_X1 U22325 ( .A1(n19737), .A2(n19396), .B1(n19388), .B2(n19798), .ZN(
        n19382) );
  OAI211_X1 U22326 ( .C1(n19385), .C2(n19384), .A(n19383), .B(n19382), .ZN(
        P2_U3074) );
  AOI22_X1 U22327 ( .A1(n19691), .A2(n19431), .B1(n19395), .B2(n19740), .ZN(
        n19387) );
  AOI22_X1 U22328 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19397), .B1(
        n19741), .B2(n19396), .ZN(n19386) );
  OAI211_X1 U22329 ( .C1(n19694), .C2(n19400), .A(n19387), .B(n19386), .ZN(
        P2_U3075) );
  AOI22_X1 U22330 ( .A1(n19812), .A2(n19388), .B1(n19395), .B2(n19744), .ZN(
        n19390) );
  AOI22_X1 U22331 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19397), .B1(
        n19746), .B2(n19396), .ZN(n19389) );
  OAI211_X1 U22332 ( .C1(n19815), .C2(n19428), .A(n19390), .B(n19389), .ZN(
        P2_U3076) );
  AOI22_X1 U22333 ( .A1(n19819), .A2(n19431), .B1(n19395), .B2(n19749), .ZN(
        n19392) );
  AOI22_X1 U22334 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19397), .B1(
        n19750), .B2(n19396), .ZN(n19391) );
  OAI211_X1 U22335 ( .C1(n19824), .C2(n19400), .A(n19392), .B(n19391), .ZN(
        P2_U3077) );
  AOI22_X1 U22336 ( .A1(n19754), .A2(n19431), .B1(n19395), .B2(n19753), .ZN(
        n19394) );
  AOI22_X1 U22337 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19397), .B1(
        n19755), .B2(n19396), .ZN(n19393) );
  OAI211_X1 U22338 ( .C1(n19758), .C2(n19400), .A(n19394), .B(n19393), .ZN(
        P2_U3078) );
  AOI22_X1 U22339 ( .A1(n19761), .A2(n19431), .B1(n19395), .B2(n19760), .ZN(
        n19399) );
  AOI22_X1 U22340 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19397), .B1(
        n19763), .B2(n19396), .ZN(n19398) );
  OAI211_X1 U22341 ( .C1(n19768), .C2(n19400), .A(n19399), .B(n19398), .ZN(
        P2_U3079) );
  NAND2_X1 U22342 ( .A1(n11572), .A2(n19645), .ZN(n19402) );
  NAND3_X1 U22343 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19938), .A3(
        n19956), .ZN(n19438) );
  NOR2_X1 U22344 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19438), .ZN(
        n19429) );
  NOR2_X1 U22345 ( .A1(n19939), .A2(n19429), .ZN(n19401) );
  NAND2_X1 U22346 ( .A1(n19402), .A2(n19401), .ZN(n19409) );
  INV_X1 U22347 ( .A(n19403), .ZN(n19405) );
  NOR2_X1 U22348 ( .A1(n19405), .A2(n19404), .ZN(n19652) );
  NAND2_X1 U22349 ( .A1(n19652), .A2(n19938), .ZN(n19411) );
  OAI21_X1 U22350 ( .B1(n19431), .B2(n19455), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19406) );
  NAND2_X1 U22351 ( .A1(n19411), .A2(n19406), .ZN(n19407) );
  AND2_X1 U22352 ( .A1(n19781), .A2(n19407), .ZN(n19408) );
  INV_X1 U22353 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n19414) );
  OAI21_X1 U22354 ( .B1(n11572), .B2(n19429), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19410) );
  OAI21_X1 U22355 ( .B1(n19411), .B2(n19719), .A(n19410), .ZN(n19430) );
  AOI22_X1 U22356 ( .A1(n19430), .A2(n19727), .B1(n19716), .B2(n19429), .ZN(
        n19413) );
  AOI22_X1 U22357 ( .A1(n19455), .A2(n19784), .B1(n19431), .B2(n19682), .ZN(
        n19412) );
  OAI211_X1 U22358 ( .C1(n19415), .C2(n19414), .A(n19413), .B(n19412), .ZN(
        P2_U3080) );
  AOI22_X1 U22359 ( .A1(n19430), .A2(n19732), .B1(n19730), .B2(n19429), .ZN(
        n19417) );
  AOI22_X1 U22360 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19432), .B1(
        n19455), .B2(n19791), .ZN(n19416) );
  OAI211_X1 U22361 ( .C1(n19794), .C2(n19428), .A(n19417), .B(n19416), .ZN(
        P2_U3081) );
  AOI22_X1 U22362 ( .A1(n19430), .A2(n19737), .B1(n19736), .B2(n19429), .ZN(
        n19419) );
  AOI22_X1 U22363 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19432), .B1(
        n19431), .B2(n19798), .ZN(n19418) );
  OAI211_X1 U22364 ( .C1(n19801), .C2(n19454), .A(n19419), .B(n19418), .ZN(
        P2_U3082) );
  AOI22_X1 U22365 ( .A1(n19430), .A2(n19741), .B1(n19740), .B2(n19429), .ZN(
        n19421) );
  AOI22_X1 U22366 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19432), .B1(
        n19431), .B2(n19805), .ZN(n19420) );
  OAI211_X1 U22367 ( .C1(n19808), .C2(n19454), .A(n19421), .B(n19420), .ZN(
        P2_U3083) );
  AOI22_X1 U22368 ( .A1(n19430), .A2(n19746), .B1(n19744), .B2(n19429), .ZN(
        n19423) );
  AOI22_X1 U22369 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19432), .B1(
        n19431), .B2(n19812), .ZN(n19422) );
  OAI211_X1 U22370 ( .C1(n19815), .C2(n19454), .A(n19423), .B(n19422), .ZN(
        P2_U3084) );
  AOI22_X1 U22371 ( .A1(n19430), .A2(n19750), .B1(n19749), .B2(n19429), .ZN(
        n19425) );
  AOI22_X1 U22372 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19432), .B1(
        n19455), .B2(n19819), .ZN(n19424) );
  OAI211_X1 U22373 ( .C1(n19824), .C2(n19428), .A(n19425), .B(n19424), .ZN(
        P2_U3085) );
  AOI22_X1 U22374 ( .A1(n19430), .A2(n19755), .B1(n19753), .B2(n19429), .ZN(
        n19427) );
  AOI22_X1 U22375 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19432), .B1(
        n19455), .B2(n19754), .ZN(n19426) );
  OAI211_X1 U22376 ( .C1(n19758), .C2(n19428), .A(n19427), .B(n19426), .ZN(
        P2_U3086) );
  AOI22_X1 U22377 ( .A1(n19430), .A2(n19763), .B1(n19760), .B2(n19429), .ZN(
        n19434) );
  AOI22_X1 U22378 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19432), .B1(
        n19431), .B2(n19837), .ZN(n19433) );
  OAI211_X1 U22379 ( .C1(n19843), .C2(n19454), .A(n19434), .B(n19433), .ZN(
        P2_U3087) );
  NOR2_X1 U22380 ( .A1(n19966), .A2(n19438), .ZN(n19464) );
  AOI22_X1 U22381 ( .A1(n19682), .A2(n19455), .B1(n19716), .B2(n19464), .ZN(
        n19441) );
  AOI21_X1 U22382 ( .B1(n19932), .B2(n10178), .A(n19719), .ZN(n19436) );
  NOR2_X1 U22383 ( .A1(n11565), .A2(n19464), .ZN(n19437) );
  AOI22_X1 U22384 ( .A1(n19436), .A2(n19438), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19437), .ZN(n19435) );
  OAI211_X1 U22385 ( .C1(n19464), .C2(n19645), .A(n19435), .B(n19781), .ZN(
        n19457) );
  INV_X1 U22386 ( .A(n19436), .ZN(n19439) );
  OAI22_X1 U22387 ( .A1(n19439), .A2(n19438), .B1(n19437), .B2(n19769), .ZN(
        n19456) );
  AOI22_X1 U22388 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19457), .B1(
        n19727), .B2(n19456), .ZN(n19440) );
  OAI211_X1 U22389 ( .C1(n19623), .C2(n19482), .A(n19441), .B(n19440), .ZN(
        P2_U3088) );
  AOI22_X1 U22390 ( .A1(n19731), .A2(n19455), .B1(n19730), .B2(n19464), .ZN(
        n19443) );
  AOI22_X1 U22391 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19457), .B1(
        n19732), .B2(n19456), .ZN(n19442) );
  OAI211_X1 U22392 ( .C1(n19735), .C2(n19482), .A(n19443), .B(n19442), .ZN(
        P2_U3089) );
  AOI22_X1 U22393 ( .A1(n19798), .A2(n19455), .B1(n19736), .B2(n19464), .ZN(
        n19445) );
  AOI22_X1 U22394 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19457), .B1(
        n19737), .B2(n19456), .ZN(n19444) );
  OAI211_X1 U22395 ( .C1(n19801), .C2(n19482), .A(n19445), .B(n19444), .ZN(
        P2_U3090) );
  AOI22_X1 U22396 ( .A1(n19805), .A2(n19455), .B1(n19464), .B2(n19740), .ZN(
        n19447) );
  AOI22_X1 U22397 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19457), .B1(
        n19741), .B2(n19456), .ZN(n19446) );
  OAI211_X1 U22398 ( .C1(n19808), .C2(n19482), .A(n19447), .B(n19446), .ZN(
        P2_U3091) );
  AOI22_X1 U22399 ( .A1(n19696), .A2(n19485), .B1(n19744), .B2(n19464), .ZN(
        n19449) );
  AOI22_X1 U22400 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19457), .B1(
        n19746), .B2(n19456), .ZN(n19448) );
  OAI211_X1 U22401 ( .C1(n19699), .C2(n19454), .A(n19449), .B(n19448), .ZN(
        P2_U3092) );
  AOI22_X1 U22402 ( .A1(n19819), .A2(n19485), .B1(n19464), .B2(n19749), .ZN(
        n19451) );
  AOI22_X1 U22403 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19457), .B1(
        n19750), .B2(n19456), .ZN(n19450) );
  OAI211_X1 U22404 ( .C1(n19824), .C2(n19454), .A(n19451), .B(n19450), .ZN(
        P2_U3093) );
  AOI22_X1 U22405 ( .A1(n19754), .A2(n19485), .B1(n19753), .B2(n19464), .ZN(
        n19453) );
  AOI22_X1 U22406 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19457), .B1(
        n19755), .B2(n19456), .ZN(n19452) );
  OAI211_X1 U22407 ( .C1(n19758), .C2(n19454), .A(n19453), .B(n19452), .ZN(
        P2_U3094) );
  AOI22_X1 U22408 ( .A1(n19837), .A2(n19455), .B1(n19760), .B2(n19464), .ZN(
        n19459) );
  AOI22_X1 U22409 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19457), .B1(
        n19763), .B2(n19456), .ZN(n19458) );
  OAI211_X1 U22410 ( .C1(n19843), .C2(n19482), .A(n19459), .B(n19458), .ZN(
        P2_U3095) );
  NOR2_X1 U22411 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19493), .ZN(
        n19483) );
  NOR2_X1 U22412 ( .A1(n19464), .A2(n19483), .ZN(n19460) );
  OR2_X1 U22413 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19460), .ZN(n19461) );
  NOR3_X1 U22414 ( .A1(n11562), .A2(n19483), .A3(n19769), .ZN(n19465) );
  AOI21_X1 U22415 ( .B1(n19769), .B2(n19461), .A(n19465), .ZN(n19484) );
  AOI22_X1 U22416 ( .A1(n19484), .A2(n19727), .B1(n19716), .B2(n19483), .ZN(
        n19469) );
  AOI21_X1 U22417 ( .B1(n19482), .B2(n19513), .A(n19643), .ZN(n19463) );
  AOI221_X1 U22418 ( .B1(n19645), .B2(n19464), .C1(n19645), .C2(n19463), .A(
        n19483), .ZN(n19467) );
  AOI22_X1 U22419 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19486), .B1(
        n19516), .B2(n19784), .ZN(n19468) );
  OAI211_X1 U22420 ( .C1(n19787), .C2(n19482), .A(n19469), .B(n19468), .ZN(
        P2_U3096) );
  AOI22_X1 U22421 ( .A1(n19484), .A2(n19732), .B1(n19730), .B2(n19483), .ZN(
        n19471) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19486), .B1(
        n19516), .B2(n19791), .ZN(n19470) );
  OAI211_X1 U22423 ( .C1(n19794), .C2(n19482), .A(n19471), .B(n19470), .ZN(
        P2_U3097) );
  AOI22_X1 U22424 ( .A1(n19484), .A2(n19737), .B1(n19736), .B2(n19483), .ZN(
        n19473) );
  AOI22_X1 U22425 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19486), .B1(
        n19485), .B2(n19798), .ZN(n19472) );
  OAI211_X1 U22426 ( .C1(n19801), .C2(n19513), .A(n19473), .B(n19472), .ZN(
        P2_U3098) );
  AOI22_X1 U22427 ( .A1(n19484), .A2(n19741), .B1(n19740), .B2(n19483), .ZN(
        n19475) );
  AOI22_X1 U22428 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19486), .B1(
        n19485), .B2(n19805), .ZN(n19474) );
  OAI211_X1 U22429 ( .C1(n19808), .C2(n19513), .A(n19475), .B(n19474), .ZN(
        P2_U3099) );
  AOI22_X1 U22430 ( .A1(n19484), .A2(n19746), .B1(n19744), .B2(n19483), .ZN(
        n19477) );
  AOI22_X1 U22431 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19486), .B1(
        n19516), .B2(n19696), .ZN(n19476) );
  OAI211_X1 U22432 ( .C1(n19699), .C2(n19482), .A(n19477), .B(n19476), .ZN(
        P2_U3100) );
  AOI22_X1 U22433 ( .A1(n19484), .A2(n19750), .B1(n19749), .B2(n19483), .ZN(
        n19479) );
  AOI22_X1 U22434 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19486), .B1(
        n19516), .B2(n19819), .ZN(n19478) );
  OAI211_X1 U22435 ( .C1(n19824), .C2(n19482), .A(n19479), .B(n19478), .ZN(
        P2_U3101) );
  AOI22_X1 U22436 ( .A1(n19484), .A2(n19755), .B1(n19753), .B2(n19483), .ZN(
        n19481) );
  AOI22_X1 U22437 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19486), .B1(
        n19516), .B2(n19754), .ZN(n19480) );
  OAI211_X1 U22438 ( .C1(n19758), .C2(n19482), .A(n19481), .B(n19480), .ZN(
        P2_U3102) );
  AOI22_X1 U22439 ( .A1(n19484), .A2(n19763), .B1(n19760), .B2(n19483), .ZN(
        n19488) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19486), .B1(
        n19485), .B2(n19837), .ZN(n19487) );
  OAI211_X1 U22441 ( .C1(n19843), .C2(n19513), .A(n19488), .B(n19487), .ZN(
        P2_U3103) );
  INV_X1 U22442 ( .A(n11567), .ZN(n19491) );
  AND2_X1 U22443 ( .A1(n19524), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19490) );
  NAND2_X1 U22444 ( .A1(n19491), .A2(n19490), .ZN(n19497) );
  OAI21_X1 U22445 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19493), .A(n19769), 
        .ZN(n19492) );
  AND2_X1 U22446 ( .A1(n19497), .A2(n19492), .ZN(n19515) );
  INV_X1 U22447 ( .A(n19524), .ZN(n19514) );
  AOI22_X1 U22448 ( .A1(n19515), .A2(n19727), .B1(n19514), .B2(n19716), .ZN(
        n19500) );
  INV_X1 U22449 ( .A(n19932), .ZN(n19495) );
  OAI21_X1 U22450 ( .B1(n19495), .B2(n19494), .A(n19493), .ZN(n19498) );
  NAND2_X1 U22451 ( .A1(n19524), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19496) );
  NAND4_X1 U22452 ( .A1(n19498), .A2(n19781), .A3(n19497), .A4(n19496), .ZN(
        n19517) );
  AOI22_X1 U22453 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19517), .B1(
        n19516), .B2(n19682), .ZN(n19499) );
  OAI211_X1 U22454 ( .C1(n19623), .C2(n19540), .A(n19500), .B(n19499), .ZN(
        P2_U3104) );
  AOI22_X1 U22455 ( .A1(n19515), .A2(n19732), .B1(n19514), .B2(n19730), .ZN(
        n19502) );
  AOI22_X1 U22456 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19517), .B1(
        n19516), .B2(n19731), .ZN(n19501) );
  OAI211_X1 U22457 ( .C1(n19735), .C2(n19540), .A(n19502), .B(n19501), .ZN(
        P2_U3105) );
  AOI22_X1 U22458 ( .A1(n19515), .A2(n19737), .B1(n19514), .B2(n19736), .ZN(
        n19504) );
  AOI22_X1 U22459 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19517), .B1(
        n19516), .B2(n19798), .ZN(n19503) );
  OAI211_X1 U22460 ( .C1(n19801), .C2(n19540), .A(n19504), .B(n19503), .ZN(
        P2_U3106) );
  AOI22_X1 U22461 ( .A1(n19515), .A2(n19741), .B1(n19514), .B2(n19740), .ZN(
        n19506) );
  AOI22_X1 U22462 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19517), .B1(
        n19516), .B2(n19805), .ZN(n19505) );
  OAI211_X1 U22463 ( .C1(n19808), .C2(n19540), .A(n19506), .B(n19505), .ZN(
        P2_U3107) );
  AOI22_X1 U22464 ( .A1(n19515), .A2(n19746), .B1(n19514), .B2(n19744), .ZN(
        n19508) );
  AOI22_X1 U22465 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19517), .B1(
        n19516), .B2(n19812), .ZN(n19507) );
  OAI211_X1 U22466 ( .C1(n19815), .C2(n19540), .A(n19508), .B(n19507), .ZN(
        P2_U3108) );
  AOI22_X1 U22467 ( .A1(n19515), .A2(n19750), .B1(n19514), .B2(n19749), .ZN(
        n19510) );
  AOI22_X1 U22468 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19517), .B1(
        n19544), .B2(n19819), .ZN(n19509) );
  OAI211_X1 U22469 ( .C1(n19824), .C2(n19513), .A(n19510), .B(n19509), .ZN(
        P2_U3109) );
  AOI22_X1 U22470 ( .A1(n19515), .A2(n19755), .B1(n19514), .B2(n19753), .ZN(
        n19512) );
  AOI22_X1 U22471 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19517), .B1(
        n19544), .B2(n19754), .ZN(n19511) );
  OAI211_X1 U22472 ( .C1(n19758), .C2(n19513), .A(n19512), .B(n19511), .ZN(
        P2_U3110) );
  AOI22_X1 U22473 ( .A1(n19515), .A2(n19763), .B1(n19514), .B2(n19760), .ZN(
        n19519) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19517), .B1(
        n19516), .B2(n19837), .ZN(n19518) );
  OAI211_X1 U22475 ( .C1(n19843), .C2(n19540), .A(n19519), .B(n19518), .ZN(
        P2_U3111) );
  NAND2_X1 U22476 ( .A1(n19946), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19607) );
  INV_X1 U22477 ( .A(n19607), .ZN(n19610) );
  NAND2_X1 U22478 ( .A1(n19610), .A2(n19956), .ZN(n19555) );
  NOR2_X1 U22479 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19555), .ZN(
        n19543) );
  AOI22_X1 U22480 ( .A1(n19784), .A2(n19569), .B1(n19543), .B2(n19716), .ZN(
        n19529) );
  NAND2_X1 U22481 ( .A1(n19540), .A2(n19577), .ZN(n19520) );
  AOI21_X1 U22482 ( .B1(n19520), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19719), 
        .ZN(n19523) );
  AOI21_X1 U22483 ( .B1(n11554), .B2(n19645), .A(n19939), .ZN(n19521) );
  AOI21_X1 U22484 ( .B1(n19523), .B2(n19524), .A(n19521), .ZN(n19522) );
  OAI21_X1 U22485 ( .B1(n19543), .B2(n19522), .A(n19781), .ZN(n19546) );
  INV_X1 U22486 ( .A(n19523), .ZN(n19527) );
  OAI21_X1 U22487 ( .B1(n11554), .B2(n19543), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19526) );
  NOR2_X1 U22488 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19543), .ZN(n19525) );
  AOI22_X1 U22489 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19546), .B1(
        n19727), .B2(n19545), .ZN(n19528) );
  OAI211_X1 U22490 ( .C1(n19787), .C2(n19540), .A(n19529), .B(n19528), .ZN(
        P2_U3112) );
  AOI22_X1 U22491 ( .A1(n19791), .A2(n19569), .B1(n19730), .B2(n19543), .ZN(
        n19531) );
  AOI22_X1 U22492 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19546), .B1(
        n19545), .B2(n19732), .ZN(n19530) );
  OAI211_X1 U22493 ( .C1(n19794), .C2(n19540), .A(n19531), .B(n19530), .ZN(
        P2_U3113) );
  AOI22_X1 U22494 ( .A1(n19798), .A2(n19544), .B1(n19736), .B2(n19543), .ZN(
        n19533) );
  AOI22_X1 U22495 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19546), .B1(
        n19545), .B2(n19737), .ZN(n19532) );
  OAI211_X1 U22496 ( .C1(n19801), .C2(n19577), .A(n19533), .B(n19532), .ZN(
        P2_U3114) );
  AOI22_X1 U22497 ( .A1(n19691), .A2(n19569), .B1(n19543), .B2(n19740), .ZN(
        n19535) );
  AOI22_X1 U22498 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19546), .B1(
        n19545), .B2(n19741), .ZN(n19534) );
  OAI211_X1 U22499 ( .C1(n19694), .C2(n19540), .A(n19535), .B(n19534), .ZN(
        P2_U3115) );
  AOI22_X1 U22500 ( .A1(n19812), .A2(n19544), .B1(n19543), .B2(n19744), .ZN(
        n19537) );
  AOI22_X1 U22501 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19546), .B1(
        n19545), .B2(n19746), .ZN(n19536) );
  OAI211_X1 U22502 ( .C1(n19815), .C2(n19577), .A(n19537), .B(n19536), .ZN(
        P2_U3116) );
  AOI22_X1 U22503 ( .A1(n19819), .A2(n19569), .B1(n19543), .B2(n19749), .ZN(
        n19539) );
  AOI22_X1 U22504 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19546), .B1(
        n19545), .B2(n19750), .ZN(n19538) );
  OAI211_X1 U22505 ( .C1(n19824), .C2(n19540), .A(n19539), .B(n19538), .ZN(
        P2_U3117) );
  AOI22_X1 U22506 ( .A1(n19828), .A2(n19544), .B1(n19543), .B2(n19753), .ZN(
        n19542) );
  AOI22_X1 U22507 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19546), .B1(
        n19545), .B2(n19755), .ZN(n19541) );
  OAI211_X1 U22508 ( .C1(n19831), .C2(n19577), .A(n19542), .B(n19541), .ZN(
        P2_U3118) );
  AOI22_X1 U22509 ( .A1(n19837), .A2(n19544), .B1(n19543), .B2(n19760), .ZN(
        n19548) );
  AOI22_X1 U22510 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19546), .B1(
        n19545), .B2(n19763), .ZN(n19547) );
  OAI211_X1 U22511 ( .C1(n19843), .C2(n19577), .A(n19548), .B(n19547), .ZN(
        P2_U3119) );
  NOR2_X1 U22512 ( .A1(n19549), .A2(n19607), .ZN(n19572) );
  AOI22_X1 U22513 ( .A1(n19682), .A2(n19569), .B1(n19716), .B2(n19572), .ZN(
        n19558) );
  INV_X1 U22514 ( .A(n19572), .ZN(n19582) );
  NAND3_X1 U22515 ( .A1(n19550), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19582), 
        .ZN(n19552) );
  AOI21_X1 U22516 ( .B1(n19777), .B2(n19941), .A(n19719), .ZN(n19553) );
  AOI22_X1 U22517 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19582), .B1(n19553), 
        .B2(n19555), .ZN(n19551) );
  NAND3_X1 U22518 ( .A1(n19552), .A2(n19551), .A3(n19781), .ZN(n19574) );
  INV_X1 U22519 ( .A(n19553), .ZN(n19556) );
  OAI21_X1 U22520 ( .B1(n11556), .B2(n19572), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19554) );
  AOI22_X1 U22521 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19574), .B1(
        n19727), .B2(n19573), .ZN(n19557) );
  OAI211_X1 U22522 ( .C1(n19623), .C2(n19597), .A(n19558), .B(n19557), .ZN(
        P2_U3120) );
  AOI22_X1 U22523 ( .A1(n19791), .A2(n19602), .B1(n19730), .B2(n19572), .ZN(
        n19560) );
  AOI22_X1 U22524 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19574), .B1(
        n19732), .B2(n19573), .ZN(n19559) );
  OAI211_X1 U22525 ( .C1(n19794), .C2(n19577), .A(n19560), .B(n19559), .ZN(
        P2_U3121) );
  AOI22_X1 U22526 ( .A1(n19798), .A2(n19569), .B1(n19736), .B2(n19572), .ZN(
        n19562) );
  AOI22_X1 U22527 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19574), .B1(
        n19737), .B2(n19573), .ZN(n19561) );
  OAI211_X1 U22528 ( .C1(n19801), .C2(n19597), .A(n19562), .B(n19561), .ZN(
        P2_U3122) );
  AOI22_X1 U22529 ( .A1(n19805), .A2(n19569), .B1(n19740), .B2(n19572), .ZN(
        n19564) );
  AOI22_X1 U22530 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19574), .B1(
        n19741), .B2(n19573), .ZN(n19563) );
  OAI211_X1 U22531 ( .C1(n19808), .C2(n19597), .A(n19564), .B(n19563), .ZN(
        P2_U3123) );
  AOI22_X1 U22532 ( .A1(n19696), .A2(n19602), .B1(n19744), .B2(n19572), .ZN(
        n19566) );
  AOI22_X1 U22533 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19574), .B1(
        n19746), .B2(n19573), .ZN(n19565) );
  OAI211_X1 U22534 ( .C1(n19699), .C2(n19577), .A(n19566), .B(n19565), .ZN(
        P2_U3124) );
  AOI22_X1 U22535 ( .A1(n19669), .A2(n19569), .B1(n19749), .B2(n19572), .ZN(
        n19568) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19574), .B1(
        n19750), .B2(n19573), .ZN(n19567) );
  OAI211_X1 U22537 ( .C1(n19672), .C2(n19597), .A(n19568), .B(n19567), .ZN(
        P2_U3125) );
  AOI22_X1 U22538 ( .A1(n19828), .A2(n19569), .B1(n19753), .B2(n19572), .ZN(
        n19571) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19574), .B1(
        n19755), .B2(n19573), .ZN(n19570) );
  OAI211_X1 U22540 ( .C1(n19831), .C2(n19597), .A(n19571), .B(n19570), .ZN(
        P2_U3126) );
  AOI22_X1 U22541 ( .A1(n19761), .A2(n19602), .B1(n19760), .B2(n19572), .ZN(
        n19576) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19574), .B1(
        n19763), .B2(n19573), .ZN(n19575) );
  OAI211_X1 U22543 ( .C1(n19768), .C2(n19577), .A(n19576), .B(n19575), .ZN(
        P2_U3127) );
  AND2_X1 U22544 ( .A1(n19578), .A2(n19610), .ZN(n19600) );
  OAI21_X1 U22545 ( .B1(n11553), .B2(n19600), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19579) );
  OAI21_X1 U22546 ( .B1(n19607), .B2(n19580), .A(n19579), .ZN(n19601) );
  AOI22_X1 U22547 ( .A1(n19601), .A2(n19727), .B1(n19716), .B2(n19600), .ZN(
        n19586) );
  OAI21_X1 U22548 ( .B1(n19626), .B2(n19602), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19583) );
  NOR2_X1 U22549 ( .A1(n11553), .A2(n19769), .ZN(n19581) );
  AOI211_X1 U22550 ( .C1(n19583), .C2(n19582), .A(P2_STATE2_REG_3__SCAN_IN), 
        .B(n19581), .ZN(n19584) );
  OAI21_X1 U22551 ( .B1(n19584), .B2(n19600), .A(n19781), .ZN(n19603) );
  AOI22_X1 U22552 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19603), .B1(
        n19626), .B2(n19784), .ZN(n19585) );
  OAI211_X1 U22553 ( .C1(n19787), .C2(n19597), .A(n19586), .B(n19585), .ZN(
        P2_U3128) );
  AOI22_X1 U22554 ( .A1(n19601), .A2(n19732), .B1(n19730), .B2(n19600), .ZN(
        n19588) );
  AOI22_X1 U22555 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19603), .B1(
        n19626), .B2(n19791), .ZN(n19587) );
  OAI211_X1 U22556 ( .C1(n19794), .C2(n19597), .A(n19588), .B(n19587), .ZN(
        P2_U3129) );
  AOI22_X1 U22557 ( .A1(n19601), .A2(n19737), .B1(n19736), .B2(n19600), .ZN(
        n19590) );
  AOI22_X1 U22558 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19603), .B1(
        n19602), .B2(n19798), .ZN(n19589) );
  OAI211_X1 U22559 ( .C1(n19801), .C2(n19642), .A(n19590), .B(n19589), .ZN(
        P2_U3130) );
  AOI22_X1 U22560 ( .A1(n19601), .A2(n19741), .B1(n19740), .B2(n19600), .ZN(
        n19592) );
  AOI22_X1 U22561 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19603), .B1(
        n19626), .B2(n19691), .ZN(n19591) );
  OAI211_X1 U22562 ( .C1(n19694), .C2(n19597), .A(n19592), .B(n19591), .ZN(
        P2_U3131) );
  AOI22_X1 U22563 ( .A1(n19601), .A2(n19746), .B1(n19744), .B2(n19600), .ZN(
        n19594) );
  AOI22_X1 U22564 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19603), .B1(
        n19602), .B2(n19812), .ZN(n19593) );
  OAI211_X1 U22565 ( .C1(n19815), .C2(n19642), .A(n19594), .B(n19593), .ZN(
        P2_U3132) );
  AOI22_X1 U22566 ( .A1(n19601), .A2(n19750), .B1(n19749), .B2(n19600), .ZN(
        n19596) );
  AOI22_X1 U22567 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19603), .B1(
        n19626), .B2(n19819), .ZN(n19595) );
  OAI211_X1 U22568 ( .C1(n19824), .C2(n19597), .A(n19596), .B(n19595), .ZN(
        P2_U3133) );
  AOI22_X1 U22569 ( .A1(n19601), .A2(n19755), .B1(n19753), .B2(n19600), .ZN(
        n19599) );
  AOI22_X1 U22570 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19603), .B1(
        n19602), .B2(n19828), .ZN(n19598) );
  OAI211_X1 U22571 ( .C1(n19831), .C2(n19642), .A(n19599), .B(n19598), .ZN(
        P2_U3134) );
  AOI22_X1 U22572 ( .A1(n19601), .A2(n19763), .B1(n19760), .B2(n19600), .ZN(
        n19605) );
  AOI22_X1 U22573 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19603), .B1(
        n19602), .B2(n19837), .ZN(n19604) );
  OAI211_X1 U22574 ( .C1(n19843), .C2(n19642), .A(n19605), .B(n19604), .ZN(
        P2_U3135) );
  NAND2_X1 U22575 ( .A1(n19606), .A2(n19619), .ZN(n19668) );
  NOR2_X1 U22576 ( .A1(n19956), .A2(n19607), .ZN(n19620) );
  INV_X1 U22577 ( .A(n19620), .ZN(n19608) );
  OR2_X1 U22578 ( .A1(n19608), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19614) );
  INV_X1 U22579 ( .A(n19609), .ZN(n19611) );
  NAND2_X1 U22580 ( .A1(n19611), .A2(n19610), .ZN(n19615) );
  NAND2_X1 U22581 ( .A1(n19615), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19612) );
  NOR2_X1 U22582 ( .A1(n19613), .A2(n19612), .ZN(n19617) );
  AOI21_X1 U22583 ( .B1(n19769), .B2(n19614), .A(n19617), .ZN(n19638) );
  INV_X1 U22584 ( .A(n19615), .ZN(n19637) );
  AOI22_X1 U22585 ( .A1(n19638), .A2(n19727), .B1(n19716), .B2(n19637), .ZN(
        n19622) );
  OAI21_X1 U22586 ( .B1(n19637), .B2(n19645), .A(n19781), .ZN(n19616) );
  NOR2_X1 U22587 ( .A1(n19617), .A2(n19616), .ZN(n19618) );
  OAI221_X1 U22588 ( .B1(n19620), .B2(n19619), .C1(n19620), .C2(n19777), .A(
        n19618), .ZN(n19639) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19639), .B1(
        n19626), .B2(n19682), .ZN(n19621) );
  OAI211_X1 U22590 ( .C1(n19623), .C2(n19668), .A(n19622), .B(n19621), .ZN(
        P2_U3136) );
  AOI22_X1 U22591 ( .A1(n19638), .A2(n19732), .B1(n19730), .B2(n19637), .ZN(
        n19625) );
  AOI22_X1 U22592 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19639), .B1(
        n19626), .B2(n19731), .ZN(n19624) );
  OAI211_X1 U22593 ( .C1(n19735), .C2(n19668), .A(n19625), .B(n19624), .ZN(
        P2_U3137) );
  AOI22_X1 U22594 ( .A1(n19638), .A2(n19737), .B1(n19736), .B2(n19637), .ZN(
        n19628) );
  AOI22_X1 U22595 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19639), .B1(
        n19626), .B2(n19798), .ZN(n19627) );
  OAI211_X1 U22596 ( .C1(n19801), .C2(n19668), .A(n19628), .B(n19627), .ZN(
        P2_U3138) );
  AOI22_X1 U22597 ( .A1(n19638), .A2(n19741), .B1(n19740), .B2(n19637), .ZN(
        n19630) );
  AOI22_X1 U22598 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19639), .B1(
        n19677), .B2(n19691), .ZN(n19629) );
  OAI211_X1 U22599 ( .C1(n19694), .C2(n19642), .A(n19630), .B(n19629), .ZN(
        P2_U3139) );
  AOI22_X1 U22600 ( .A1(n19638), .A2(n19746), .B1(n19744), .B2(n19637), .ZN(
        n19632) );
  AOI22_X1 U22601 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19639), .B1(
        n19677), .B2(n19696), .ZN(n19631) );
  OAI211_X1 U22602 ( .C1(n19699), .C2(n19642), .A(n19632), .B(n19631), .ZN(
        P2_U3140) );
  AOI22_X1 U22603 ( .A1(n19638), .A2(n19750), .B1(n19749), .B2(n19637), .ZN(
        n19634) );
  AOI22_X1 U22604 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19639), .B1(
        n19677), .B2(n19819), .ZN(n19633) );
  OAI211_X1 U22605 ( .C1(n19824), .C2(n19642), .A(n19634), .B(n19633), .ZN(
        P2_U3141) );
  AOI22_X1 U22606 ( .A1(n19638), .A2(n19755), .B1(n19753), .B2(n19637), .ZN(
        n19636) );
  AOI22_X1 U22607 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19639), .B1(
        n19677), .B2(n19754), .ZN(n19635) );
  OAI211_X1 U22608 ( .C1(n19758), .C2(n19642), .A(n19636), .B(n19635), .ZN(
        P2_U3142) );
  AOI22_X1 U22609 ( .A1(n19638), .A2(n19763), .B1(n19760), .B2(n19637), .ZN(
        n19641) );
  AOI22_X1 U22610 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19639), .B1(
        n19677), .B2(n19761), .ZN(n19640) );
  OAI211_X1 U22611 ( .C1(n19768), .C2(n19642), .A(n19641), .B(n19640), .ZN(
        P2_U3143) );
  AOI21_X1 U22612 ( .B1(n19668), .B2(n19703), .A(n19643), .ZN(n19644) );
  AOI21_X1 U22613 ( .B1(n19652), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n19644), .ZN(n19651) );
  NAND2_X1 U22614 ( .A1(n11557), .A2(n19645), .ZN(n19648) );
  NOR2_X1 U22615 ( .A1(n19646), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19675) );
  INV_X1 U22616 ( .A(n19675), .ZN(n19647) );
  NAND3_X1 U22617 ( .A1(n19648), .A2(n19647), .A3(n19719), .ZN(n19649) );
  NAND2_X1 U22618 ( .A1(n19649), .A2(n19781), .ZN(n19650) );
  INV_X1 U22619 ( .A(n19678), .ZN(n19659) );
  INV_X1 U22620 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n19658) );
  INV_X1 U22621 ( .A(n19652), .ZN(n19654) );
  OAI21_X1 U22622 ( .B1(n11557), .B2(n19675), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19653) );
  OAI21_X1 U22623 ( .B1(n19655), .B2(n19654), .A(n19653), .ZN(n19676) );
  AOI22_X1 U22624 ( .A1(n19676), .A2(n19727), .B1(n19716), .B2(n19675), .ZN(
        n19657) );
  AOI22_X1 U22625 ( .A1(n19710), .A2(n19784), .B1(n19677), .B2(n19682), .ZN(
        n19656) );
  OAI211_X1 U22626 ( .C1(n19659), .C2(n19658), .A(n19657), .B(n19656), .ZN(
        P2_U3144) );
  AOI22_X1 U22627 ( .A1(n19676), .A2(n19732), .B1(n19730), .B2(n19675), .ZN(
        n19661) );
  AOI22_X1 U22628 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19678), .B1(
        n19677), .B2(n19731), .ZN(n19660) );
  OAI211_X1 U22629 ( .C1(n19735), .C2(n19703), .A(n19661), .B(n19660), .ZN(
        P2_U3145) );
  AOI22_X1 U22630 ( .A1(n19676), .A2(n19737), .B1(n19736), .B2(n19675), .ZN(
        n19663) );
  AOI22_X1 U22631 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19678), .B1(
        n19677), .B2(n19798), .ZN(n19662) );
  OAI211_X1 U22632 ( .C1(n19801), .C2(n19703), .A(n19663), .B(n19662), .ZN(
        P2_U3146) );
  AOI22_X1 U22633 ( .A1(n19676), .A2(n19741), .B1(n19740), .B2(n19675), .ZN(
        n19665) );
  AOI22_X1 U22634 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19678), .B1(
        n19677), .B2(n19805), .ZN(n19664) );
  OAI211_X1 U22635 ( .C1(n19808), .C2(n19703), .A(n19665), .B(n19664), .ZN(
        P2_U3147) );
  AOI22_X1 U22636 ( .A1(n19676), .A2(n19746), .B1(n19744), .B2(n19675), .ZN(
        n19667) );
  AOI22_X1 U22637 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19678), .B1(
        n19710), .B2(n19696), .ZN(n19666) );
  OAI211_X1 U22638 ( .C1(n19699), .C2(n19668), .A(n19667), .B(n19666), .ZN(
        P2_U3148) );
  AOI22_X1 U22639 ( .A1(n19676), .A2(n19750), .B1(n19749), .B2(n19675), .ZN(
        n19671) );
  AOI22_X1 U22640 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19678), .B1(
        n19677), .B2(n19669), .ZN(n19670) );
  OAI211_X1 U22641 ( .C1(n19672), .C2(n19703), .A(n19671), .B(n19670), .ZN(
        P2_U3149) );
  AOI22_X1 U22642 ( .A1(n19676), .A2(n19755), .B1(n19753), .B2(n19675), .ZN(
        n19674) );
  AOI22_X1 U22643 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19678), .B1(
        n19677), .B2(n19828), .ZN(n19673) );
  OAI211_X1 U22644 ( .C1(n19831), .C2(n19703), .A(n19674), .B(n19673), .ZN(
        P2_U3150) );
  AOI22_X1 U22645 ( .A1(n19676), .A2(n19763), .B1(n19760), .B2(n19675), .ZN(
        n19680) );
  AOI22_X1 U22646 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19678), .B1(
        n19677), .B2(n19837), .ZN(n19679) );
  OAI211_X1 U22647 ( .C1(n19843), .C2(n19703), .A(n19680), .B(n19679), .ZN(
        P2_U3151) );
  INV_X1 U22648 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n19685) );
  OAI22_X1 U22649 ( .A1(n19708), .A2(n19775), .B1(n19707), .B2(n19774), .ZN(
        n19681) );
  INV_X1 U22650 ( .A(n19681), .ZN(n19684) );
  AOI22_X1 U22651 ( .A1(n19745), .A2(n19784), .B1(n19710), .B2(n19682), .ZN(
        n19683) );
  OAI211_X1 U22652 ( .C1(n19686), .C2(n19685), .A(n19684), .B(n19683), .ZN(
        P2_U3152) );
  OAI22_X1 U22653 ( .A1(n19708), .A2(n19796), .B1(n19707), .B2(n19795), .ZN(
        n19687) );
  INV_X1 U22654 ( .A(n19687), .ZN(n19689) );
  AOI22_X1 U22655 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19711), .B1(
        n19710), .B2(n19798), .ZN(n19688) );
  OAI211_X1 U22656 ( .C1(n19801), .C2(n19767), .A(n19689), .B(n19688), .ZN(
        P2_U3154) );
  OAI22_X1 U22657 ( .A1(n19708), .A2(n19803), .B1(n19707), .B2(n19802), .ZN(
        n19690) );
  INV_X1 U22658 ( .A(n19690), .ZN(n19693) );
  AOI22_X1 U22659 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19711), .B1(
        n19745), .B2(n19691), .ZN(n19692) );
  OAI211_X1 U22660 ( .C1(n19694), .C2(n19703), .A(n19693), .B(n19692), .ZN(
        P2_U3155) );
  OAI22_X1 U22661 ( .A1(n19708), .A2(n19810), .B1(n19707), .B2(n19809), .ZN(
        n19695) );
  INV_X1 U22662 ( .A(n19695), .ZN(n19698) );
  AOI22_X1 U22663 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19711), .B1(
        n19745), .B2(n19696), .ZN(n19697) );
  OAI211_X1 U22664 ( .C1(n19699), .C2(n19703), .A(n19698), .B(n19697), .ZN(
        P2_U3156) );
  OAI22_X1 U22665 ( .A1(n19708), .A2(n19817), .B1(n19707), .B2(n19816), .ZN(
        n19700) );
  INV_X1 U22666 ( .A(n19700), .ZN(n19702) );
  AOI22_X1 U22667 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19711), .B1(
        n19745), .B2(n19819), .ZN(n19701) );
  OAI211_X1 U22668 ( .C1(n19824), .C2(n19703), .A(n19702), .B(n19701), .ZN(
        P2_U3157) );
  OAI22_X1 U22669 ( .A1(n19708), .A2(n19826), .B1(n19707), .B2(n19825), .ZN(
        n19704) );
  INV_X1 U22670 ( .A(n19704), .ZN(n19706) );
  AOI22_X1 U22671 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19711), .B1(
        n19710), .B2(n19828), .ZN(n19705) );
  OAI211_X1 U22672 ( .C1(n19831), .C2(n19767), .A(n19706), .B(n19705), .ZN(
        P2_U3158) );
  OAI22_X1 U22673 ( .A1(n19708), .A2(n19834), .B1(n19707), .B2(n19833), .ZN(
        n19709) );
  INV_X1 U22674 ( .A(n19709), .ZN(n19713) );
  AOI22_X1 U22675 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19711), .B1(
        n19710), .B2(n19837), .ZN(n19712) );
  OAI211_X1 U22676 ( .C1(n19843), .C2(n19767), .A(n19713), .B(n19712), .ZN(
        P2_U3159) );
  NAND2_X1 U22677 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19715), .ZN(
        n19779) );
  NOR2_X1 U22678 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19779), .ZN(
        n19759) );
  AOI22_X1 U22679 ( .A1(n19784), .A2(n19838), .B1(n19716), .B2(n19759), .ZN(
        n19729) );
  OAI21_X1 U22680 ( .B1(n19838), .B2(n19745), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19717) );
  NAND2_X1 U22681 ( .A1(n19717), .A2(n19939), .ZN(n19726) );
  NOR2_X1 U22682 ( .A1(n19759), .A2(n19718), .ZN(n19725) );
  INV_X1 U22683 ( .A(n19725), .ZN(n19723) );
  INV_X1 U22684 ( .A(n11564), .ZN(n19721) );
  INV_X1 U22685 ( .A(n19759), .ZN(n19720) );
  OAI211_X1 U22686 ( .C1(n19721), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19720), 
        .B(n19719), .ZN(n19722) );
  OAI211_X1 U22687 ( .C1(n19726), .C2(n19723), .A(n19781), .B(n19722), .ZN(
        n19764) );
  OAI21_X1 U22688 ( .B1(n11564), .B2(n19759), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19724) );
  AOI22_X1 U22689 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19764), .B1(
        n19727), .B2(n19762), .ZN(n19728) );
  OAI211_X1 U22690 ( .C1(n19787), .C2(n19767), .A(n19729), .B(n19728), .ZN(
        P2_U3160) );
  AOI22_X1 U22691 ( .A1(n19731), .A2(n19745), .B1(n19730), .B2(n19759), .ZN(
        n19734) );
  AOI22_X1 U22692 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19764), .B1(
        n19732), .B2(n19762), .ZN(n19733) );
  OAI211_X1 U22693 ( .C1(n19735), .C2(n19823), .A(n19734), .B(n19733), .ZN(
        P2_U3161) );
  AOI22_X1 U22694 ( .A1(n19798), .A2(n19745), .B1(n19736), .B2(n19759), .ZN(
        n19739) );
  AOI22_X1 U22695 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19764), .B1(
        n19737), .B2(n19762), .ZN(n19738) );
  OAI211_X1 U22696 ( .C1(n19801), .C2(n19823), .A(n19739), .B(n19738), .ZN(
        P2_U3162) );
  AOI22_X1 U22697 ( .A1(n19805), .A2(n19745), .B1(n19740), .B2(n19759), .ZN(
        n19743) );
  AOI22_X1 U22698 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19764), .B1(
        n19741), .B2(n19762), .ZN(n19742) );
  OAI211_X1 U22699 ( .C1(n19808), .C2(n19823), .A(n19743), .B(n19742), .ZN(
        P2_U3163) );
  AOI22_X1 U22700 ( .A1(n19812), .A2(n19745), .B1(n19744), .B2(n19759), .ZN(
        n19748) );
  AOI22_X1 U22701 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19764), .B1(
        n19746), .B2(n19762), .ZN(n19747) );
  OAI211_X1 U22702 ( .C1(n19815), .C2(n19823), .A(n19748), .B(n19747), .ZN(
        P2_U3164) );
  AOI22_X1 U22703 ( .A1(n19819), .A2(n19838), .B1(n19749), .B2(n19759), .ZN(
        n19752) );
  AOI22_X1 U22704 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19764), .B1(
        n19750), .B2(n19762), .ZN(n19751) );
  OAI211_X1 U22705 ( .C1(n19824), .C2(n19767), .A(n19752), .B(n19751), .ZN(
        P2_U3165) );
  AOI22_X1 U22706 ( .A1(n19754), .A2(n19838), .B1(n19753), .B2(n19759), .ZN(
        n19757) );
  AOI22_X1 U22707 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19764), .B1(
        n19755), .B2(n19762), .ZN(n19756) );
  OAI211_X1 U22708 ( .C1(n19758), .C2(n19767), .A(n19757), .B(n19756), .ZN(
        P2_U3166) );
  AOI22_X1 U22709 ( .A1(n19761), .A2(n19838), .B1(n19760), .B2(n19759), .ZN(
        n19766) );
  AOI22_X1 U22710 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19764), .B1(
        n19763), .B2(n19762), .ZN(n19765) );
  OAI211_X1 U22711 ( .C1(n19768), .C2(n19767), .A(n19766), .B(n19765), .ZN(
        P2_U3167) );
  OR2_X1 U22712 ( .A1(n19783), .A2(n19769), .ZN(n19770) );
  NOR2_X1 U22713 ( .A1(n19771), .A2(n19770), .ZN(n19778) );
  INV_X1 U22714 ( .A(n19779), .ZN(n19772) );
  AOI21_X1 U22715 ( .B1(n19645), .B2(n19772), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19773) );
  OR2_X1 U22716 ( .A1(n19778), .A2(n19773), .ZN(n19835) );
  INV_X1 U22717 ( .A(n19783), .ZN(n19832) );
  OAI22_X1 U22718 ( .A1(n19835), .A2(n19775), .B1(n19774), .B2(n19832), .ZN(
        n19776) );
  INV_X1 U22719 ( .A(n19776), .ZN(n19786) );
  NAND2_X1 U22720 ( .A1(n19777), .A2(n19931), .ZN(n19780) );
  AOI21_X1 U22721 ( .B1(n19780), .B2(n19779), .A(n19778), .ZN(n19782) );
  OAI211_X1 U22722 ( .C1(n19783), .C2(n19645), .A(n19782), .B(n19781), .ZN(
        n19839) );
  AOI22_X1 U22723 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19839), .B1(
        n19820), .B2(n19784), .ZN(n19785) );
  OAI211_X1 U22724 ( .C1(n19787), .C2(n19823), .A(n19786), .B(n19785), .ZN(
        P2_U3168) );
  OAI22_X1 U22725 ( .A1(n19835), .A2(n19789), .B1(n19788), .B2(n19832), .ZN(
        n19790) );
  INV_X1 U22726 ( .A(n19790), .ZN(n19793) );
  AOI22_X1 U22727 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19839), .B1(
        n19820), .B2(n19791), .ZN(n19792) );
  OAI211_X1 U22728 ( .C1(n19794), .C2(n19823), .A(n19793), .B(n19792), .ZN(
        P2_U3169) );
  OAI22_X1 U22729 ( .A1(n19835), .A2(n19796), .B1(n19795), .B2(n19832), .ZN(
        n19797) );
  INV_X1 U22730 ( .A(n19797), .ZN(n19800) );
  AOI22_X1 U22731 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19839), .B1(
        n19838), .B2(n19798), .ZN(n19799) );
  OAI211_X1 U22732 ( .C1(n19801), .C2(n19842), .A(n19800), .B(n19799), .ZN(
        P2_U3170) );
  OAI22_X1 U22733 ( .A1(n19835), .A2(n19803), .B1(n19802), .B2(n19832), .ZN(
        n19804) );
  INV_X1 U22734 ( .A(n19804), .ZN(n19807) );
  AOI22_X1 U22735 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19839), .B1(
        n19838), .B2(n19805), .ZN(n19806) );
  OAI211_X1 U22736 ( .C1(n19808), .C2(n19842), .A(n19807), .B(n19806), .ZN(
        P2_U3171) );
  OAI22_X1 U22737 ( .A1(n19835), .A2(n19810), .B1(n19809), .B2(n19832), .ZN(
        n19811) );
  INV_X1 U22738 ( .A(n19811), .ZN(n19814) );
  AOI22_X1 U22739 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19839), .B1(
        n19838), .B2(n19812), .ZN(n19813) );
  OAI211_X1 U22740 ( .C1(n19815), .C2(n19842), .A(n19814), .B(n19813), .ZN(
        P2_U3172) );
  OAI22_X1 U22741 ( .A1(n19835), .A2(n19817), .B1(n19816), .B2(n19832), .ZN(
        n19818) );
  INV_X1 U22742 ( .A(n19818), .ZN(n19822) );
  AOI22_X1 U22743 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19839), .B1(
        n19820), .B2(n19819), .ZN(n19821) );
  OAI211_X1 U22744 ( .C1(n19824), .C2(n19823), .A(n19822), .B(n19821), .ZN(
        P2_U3173) );
  OAI22_X1 U22745 ( .A1(n19835), .A2(n19826), .B1(n19825), .B2(n19832), .ZN(
        n19827) );
  INV_X1 U22746 ( .A(n19827), .ZN(n19830) );
  AOI22_X1 U22747 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19839), .B1(
        n19838), .B2(n19828), .ZN(n19829) );
  OAI211_X1 U22748 ( .C1(n19831), .C2(n19842), .A(n19830), .B(n19829), .ZN(
        P2_U3174) );
  OAI22_X1 U22749 ( .A1(n19835), .A2(n19834), .B1(n19833), .B2(n19832), .ZN(
        n19836) );
  INV_X1 U22750 ( .A(n19836), .ZN(n19841) );
  AOI22_X1 U22751 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19839), .B1(
        n19838), .B2(n19837), .ZN(n19840) );
  OAI211_X1 U22752 ( .C1(n19843), .C2(n19842), .A(n19841), .B(n19840), .ZN(
        P2_U3175) );
  NOR2_X1 U22753 ( .A1(n11444), .A2(n19985), .ZN(n19850) );
  NAND2_X1 U22754 ( .A1(n19848), .A2(n19844), .ZN(n19849) );
  OAI21_X1 U22755 ( .B1(n19867), .B2(n19846), .A(n19845), .ZN(n19847) );
  AOI22_X1 U22756 ( .A1(n19850), .A2(n19849), .B1(n19848), .B2(n19847), .ZN(
        n19852) );
  NAND2_X1 U22757 ( .A1(n19852), .A2(n19851), .ZN(P2_U3177) );
  INV_X1 U22758 ( .A(n19928), .ZN(n19853) );
  AND2_X1 U22759 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19853), .ZN(
        P2_U3179) );
  AND2_X1 U22760 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19853), .ZN(
        P2_U3180) );
  AND2_X1 U22761 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19853), .ZN(
        P2_U3181) );
  AND2_X1 U22762 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19853), .ZN(
        P2_U3182) );
  AND2_X1 U22763 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19853), .ZN(
        P2_U3183) );
  AND2_X1 U22764 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19853), .ZN(
        P2_U3184) );
  AND2_X1 U22765 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19853), .ZN(
        P2_U3185) );
  AND2_X1 U22766 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19853), .ZN(
        P2_U3186) );
  AND2_X1 U22767 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19853), .ZN(
        P2_U3187) );
  AND2_X1 U22768 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19853), .ZN(
        P2_U3188) );
  AND2_X1 U22769 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19853), .ZN(
        P2_U3189) );
  AND2_X1 U22770 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19853), .ZN(
        P2_U3190) );
  AND2_X1 U22771 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19853), .ZN(
        P2_U3191) );
  AND2_X1 U22772 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19853), .ZN(
        P2_U3192) );
  AND2_X1 U22773 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19853), .ZN(
        P2_U3193) );
  AND2_X1 U22774 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19853), .ZN(
        P2_U3194) );
  AND2_X1 U22775 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19853), .ZN(
        P2_U3195) );
  AND2_X1 U22776 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19853), .ZN(
        P2_U3196) );
  AND2_X1 U22777 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19853), .ZN(
        P2_U3197) );
  AND2_X1 U22778 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19853), .ZN(
        P2_U3198) );
  AND2_X1 U22779 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19853), .ZN(
        P2_U3199) );
  AND2_X1 U22780 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19853), .ZN(
        P2_U3200) );
  AND2_X1 U22781 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19853), .ZN(P2_U3201) );
  AND2_X1 U22782 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19853), .ZN(P2_U3202) );
  AND2_X1 U22783 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19853), .ZN(P2_U3203) );
  AND2_X1 U22784 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19853), .ZN(P2_U3204) );
  AND2_X1 U22785 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19853), .ZN(P2_U3205) );
  AND2_X1 U22786 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19853), .ZN(P2_U3206) );
  AND2_X1 U22787 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19853), .ZN(P2_U3207) );
  AND2_X1 U22788 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19853), .ZN(P2_U3208) );
  NOR2_X1 U22789 ( .A1(n19864), .A2(n19985), .ZN(n19862) );
  INV_X1 U22790 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19995) );
  OR3_X1 U22791 ( .A1(n19862), .A2(n19995), .A3(n19854), .ZN(n19856) );
  INV_X2 U22792 ( .A(n19997), .ZN(n19918) );
  AOI211_X1 U22793 ( .C1(n21063), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n19863), .B(n19918), .ZN(n19855) );
  NOR3_X1 U22794 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n21031), .ZN(n19869) );
  AOI211_X1 U22795 ( .C1(n19872), .C2(n19856), .A(n19855), .B(n19869), .ZN(
        n19857) );
  INV_X1 U22796 ( .A(n19857), .ZN(P2_U3209) );
  AOI21_X1 U22797 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21063), .A(n19872), 
        .ZN(n19865) );
  NOR3_X1 U22798 ( .A1(n19865), .A2(n19995), .A3(n19854), .ZN(n19858) );
  NOR2_X1 U22799 ( .A1(n19858), .A2(n19862), .ZN(n19860) );
  OAI211_X1 U22800 ( .C1(n21063), .C2(n19861), .A(n19860), .B(n19859), .ZN(
        P2_U3210) );
  AOI22_X1 U22801 ( .A1(n19863), .A2(n19995), .B1(n19862), .B2(n21031), .ZN(
        n19871) );
  OAI21_X1 U22802 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n19870) );
  NOR2_X1 U22803 ( .A1(n19864), .A2(n19872), .ZN(n19866) );
  AOI21_X1 U22804 ( .B1(n19867), .B2(n19866), .A(n19865), .ZN(n19868) );
  OAI22_X1 U22805 ( .A1(n19871), .A2(n19870), .B1(n19869), .B2(n19868), .ZN(
        P2_U3211) );
  NAND2_X1 U22806 ( .A1(n19918), .A2(n19872), .ZN(n19921) );
  CLKBUF_X1 U22807 ( .A(n19921), .Z(n19915) );
  OAI222_X1 U22808 ( .A1(n19915), .A2(n11440), .B1(n19873), .B2(n19918), .C1(
        n11445), .C2(n19916), .ZN(P2_U3212) );
  OAI222_X1 U22809 ( .A1(n19921), .A2(n11430), .B1(n19874), .B2(n19918), .C1(
        n11440), .C2(n19916), .ZN(P2_U3213) );
  OAI222_X1 U22810 ( .A1(n19921), .A2(n11860), .B1(n19875), .B2(n19918), .C1(
        n11430), .C2(n19916), .ZN(P2_U3214) );
  OAI222_X1 U22811 ( .A1(n19921), .A2(n11864), .B1(n19876), .B2(n19918), .C1(
        n11860), .C2(n19916), .ZN(P2_U3215) );
  OAI222_X1 U22812 ( .A1(n19921), .A2(n11869), .B1(n19877), .B2(n19918), .C1(
        n11864), .C2(n19916), .ZN(P2_U3216) );
  OAI222_X1 U22813 ( .A1(n19921), .A2(n19879), .B1(n19878), .B2(n19918), .C1(
        n11869), .C2(n19916), .ZN(P2_U3217) );
  OAI222_X1 U22814 ( .A1(n19921), .A2(n13590), .B1(n19880), .B2(n19918), .C1(
        n19879), .C2(n19916), .ZN(P2_U3218) );
  OAI222_X1 U22815 ( .A1(n19915), .A2(n11879), .B1(n19881), .B2(n19918), .C1(
        n13590), .C2(n19916), .ZN(P2_U3219) );
  OAI222_X1 U22816 ( .A1(n19915), .A2(n13578), .B1(n19882), .B2(n19918), .C1(
        n11879), .C2(n19916), .ZN(P2_U3220) );
  OAI222_X1 U22817 ( .A1(n19915), .A2(n11888), .B1(n19883), .B2(n19918), .C1(
        n13578), .C2(n19916), .ZN(P2_U3221) );
  OAI222_X1 U22818 ( .A1(n19915), .A2(n12425), .B1(n19884), .B2(n19918), .C1(
        n11888), .C2(n19916), .ZN(P2_U3222) );
  OAI222_X1 U22819 ( .A1(n19915), .A2(n11895), .B1(n19885), .B2(n19918), .C1(
        n12425), .C2(n19916), .ZN(P2_U3223) );
  OAI222_X1 U22820 ( .A1(n19915), .A2(n11902), .B1(n19886), .B2(n19918), .C1(
        n11895), .C2(n19916), .ZN(P2_U3224) );
  OAI222_X1 U22821 ( .A1(n19915), .A2(n19888), .B1(n19887), .B2(n19918), .C1(
        n11902), .C2(n19916), .ZN(P2_U3225) );
  OAI222_X1 U22822 ( .A1(n19921), .A2(n19890), .B1(n19889), .B2(n19918), .C1(
        n19888), .C2(n19916), .ZN(P2_U3226) );
  OAI222_X1 U22823 ( .A1(n19921), .A2(n19892), .B1(n19891), .B2(n19918), .C1(
        n19890), .C2(n19916), .ZN(P2_U3227) );
  OAI222_X1 U22824 ( .A1(n19921), .A2(n15223), .B1(n19893), .B2(n19918), .C1(
        n19892), .C2(n19916), .ZN(P2_U3228) );
  OAI222_X1 U22825 ( .A1(n19921), .A2(n19895), .B1(n19894), .B2(n19918), .C1(
        n15223), .C2(n19916), .ZN(P2_U3229) );
  OAI222_X1 U22826 ( .A1(n19915), .A2(n15485), .B1(n19896), .B2(n19918), .C1(
        n19895), .C2(n19916), .ZN(P2_U3230) );
  OAI222_X1 U22827 ( .A1(n19915), .A2(n19898), .B1(n19897), .B2(n19918), .C1(
        n15485), .C2(n19916), .ZN(P2_U3231) );
  OAI222_X1 U22828 ( .A1(n19915), .A2(n19900), .B1(n19899), .B2(n19918), .C1(
        n19898), .C2(n19916), .ZN(P2_U3232) );
  OAI222_X1 U22829 ( .A1(n19915), .A2(n19902), .B1(n19901), .B2(n19918), .C1(
        n19900), .C2(n19916), .ZN(P2_U3233) );
  OAI222_X1 U22830 ( .A1(n19915), .A2(n11935), .B1(n19903), .B2(n19918), .C1(
        n19902), .C2(n19916), .ZN(P2_U3234) );
  OAI222_X1 U22831 ( .A1(n19915), .A2(n19905), .B1(n19904), .B2(n19918), .C1(
        n11935), .C2(n19916), .ZN(P2_U3235) );
  OAI222_X1 U22832 ( .A1(n19915), .A2(n19907), .B1(n19906), .B2(n19918), .C1(
        n19905), .C2(n19916), .ZN(P2_U3236) );
  OAI222_X1 U22833 ( .A1(n19915), .A2(n19910), .B1(n19908), .B2(n19918), .C1(
        n19907), .C2(n19916), .ZN(P2_U3237) );
  OAI222_X1 U22834 ( .A1(n19916), .A2(n19910), .B1(n19909), .B2(n19918), .C1(
        n19911), .C2(n19915), .ZN(P2_U3238) );
  OAI222_X1 U22835 ( .A1(n19915), .A2(n19913), .B1(n19912), .B2(n19918), .C1(
        n19911), .C2(n19916), .ZN(P2_U3239) );
  OAI222_X1 U22836 ( .A1(n19915), .A2(n19917), .B1(n19914), .B2(n19918), .C1(
        n19913), .C2(n19916), .ZN(P2_U3240) );
  INV_X1 U22837 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19919) );
  OAI222_X1 U22838 ( .A1(n19921), .A2(n19920), .B1(n19919), .B2(n19918), .C1(
        n19917), .C2(n19916), .ZN(P2_U3241) );
  OAI22_X1 U22839 ( .A1(n19997), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19918), .ZN(n19922) );
  INV_X1 U22840 ( .A(n19922), .ZN(P2_U3585) );
  MUX2_X1 U22841 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19997), .Z(P2_U3586) );
  OAI22_X1 U22842 ( .A1(n19997), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19918), .ZN(n19923) );
  INV_X1 U22843 ( .A(n19923), .ZN(P2_U3587) );
  OAI22_X1 U22844 ( .A1(n19997), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19918), .ZN(n19924) );
  INV_X1 U22845 ( .A(n19924), .ZN(P2_U3588) );
  OAI21_X1 U22846 ( .B1(n19928), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19926), 
        .ZN(n19925) );
  INV_X1 U22847 ( .A(n19925), .ZN(P2_U3591) );
  OAI21_X1 U22848 ( .B1(n19928), .B2(n19927), .A(n19926), .ZN(P2_U3592) );
  INV_X1 U22849 ( .A(n19965), .ZN(n19964) );
  NAND3_X1 U22850 ( .A1(n19931), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19929), 
        .ZN(n19930) );
  NAND2_X1 U22851 ( .A1(n19930), .A2(n19947), .ZN(n19940) );
  NAND3_X1 U22852 ( .A1(n19932), .A2(n19939), .A3(n19931), .ZN(n19933) );
  OAI21_X1 U22853 ( .B1(n19940), .B2(n19934), .A(n19933), .ZN(n19935) );
  AOI21_X1 U22854 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19936), .A(n19935), 
        .ZN(n19937) );
  AOI22_X1 U22855 ( .A1(n19964), .A2(n19938), .B1(n19937), .B2(n19965), .ZN(
        P2_U3602) );
  NAND2_X1 U22856 ( .A1(n19939), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19951) );
  AOI211_X1 U22857 ( .C1(n19942), .C2(n19951), .A(n19941), .B(n19940), .ZN(
        n19943) );
  AOI21_X1 U22858 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19944), .A(n19943), 
        .ZN(n19945) );
  AOI22_X1 U22859 ( .A1(n19964), .A2(n19946), .B1(n19945), .B2(n19965), .ZN(
        P2_U3603) );
  INV_X1 U22860 ( .A(n19947), .ZN(n19960) );
  AND2_X1 U22861 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19948) );
  OR3_X1 U22862 ( .A1(n19949), .A2(n19960), .A3(n19948), .ZN(n19950) );
  OAI21_X1 U22863 ( .B1(n19952), .B2(n19951), .A(n19950), .ZN(n19953) );
  AOI21_X1 U22864 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19954), .A(n19953), 
        .ZN(n19955) );
  AOI22_X1 U22865 ( .A1(n19964), .A2(n19956), .B1(n19955), .B2(n19965), .ZN(
        P2_U3604) );
  INV_X1 U22866 ( .A(n19957), .ZN(n19959) );
  OAI22_X1 U22867 ( .A1(n19961), .A2(n19960), .B1(n19959), .B2(n19958), .ZN(
        n19962) );
  AOI21_X1 U22868 ( .B1(n19966), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19962), 
        .ZN(n19963) );
  OAI22_X1 U22869 ( .A1(n19966), .A2(n19965), .B1(n19964), .B2(n19963), .ZN(
        P2_U3605) );
  INV_X1 U22870 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19967) );
  AOI22_X1 U22871 ( .A1(n19918), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19967), 
        .B2(n19997), .ZN(P2_U3608) );
  INV_X1 U22872 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n19977) );
  INV_X1 U22873 ( .A(n19968), .ZN(n19972) );
  AOI22_X1 U22874 ( .A1(n19972), .A2(n19971), .B1(n19970), .B2(n19969), .ZN(
        n19973) );
  NOR2_X1 U22875 ( .A1(n19973), .A2(n11397), .ZN(n19974) );
  OAI21_X1 U22876 ( .B1(n19975), .B2(n19974), .A(n19978), .ZN(n19976) );
  OAI21_X1 U22877 ( .B1(n19978), .B2(n19977), .A(n19976), .ZN(P2_U3609) );
  AOI21_X1 U22878 ( .B1(n19979), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19981) );
  AOI211_X1 U22879 ( .C1(n19985), .C2(n19982), .A(n19981), .B(n19980), .ZN(
        n19983) );
  INV_X1 U22880 ( .A(n19983), .ZN(n19996) );
  AOI21_X1 U22881 ( .B1(n19985), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n19984), 
        .ZN(n19993) );
  AOI21_X1 U22882 ( .B1(n19988), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19986), 
        .ZN(n19991) );
  NOR3_X1 U22883 ( .A1(n19988), .A2(n19987), .A3(n11388), .ZN(n19990) );
  MUX2_X1 U22884 ( .A(n19991), .B(n19990), .S(n19989), .Z(n19992) );
  OAI21_X1 U22885 ( .B1(n19993), .B2(n19992), .A(n19996), .ZN(n19994) );
  OAI21_X1 U22886 ( .B1(n19996), .B2(n19995), .A(n19994), .ZN(P2_U3610) );
  OAI22_X1 U22887 ( .A1(n19997), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19918), .ZN(n19998) );
  INV_X1 U22888 ( .A(n19998), .ZN(P2_U3611) );
  AOI21_X1 U22889 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20853), .A(n20847), 
        .ZN(n20849) );
  INV_X1 U22890 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19999) );
  NAND2_X1 U22891 ( .A1(n20847), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20899) );
  AOI21_X1 U22892 ( .B1(n20849), .B2(n19999), .A(n20923), .ZN(P1_U2802) );
  INV_X1 U22893 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n21044) );
  AOI21_X1 U22894 ( .B1(n20001), .B2(n20000), .A(n21044), .ZN(n20002) );
  AOI21_X1 U22895 ( .B1(n20003), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20002), 
        .ZN(n20004) );
  INV_X1 U22896 ( .A(n20004), .ZN(P1_U2803) );
  NOR2_X1 U22897 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20006) );
  OAI21_X1 U22898 ( .B1(n20006), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20899), .ZN(
        n20005) );
  OAI21_X1 U22899 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20899), .A(n20005), 
        .ZN(P1_U2804) );
  NOR2_X1 U22900 ( .A1(n20923), .A2(n20849), .ZN(n20904) );
  OAI21_X1 U22901 ( .B1(BS16), .B2(n20006), .A(n20904), .ZN(n20902) );
  OAI21_X1 U22902 ( .B1(n20904), .B2(n21034), .A(n20902), .ZN(P1_U2805) );
  OAI21_X1 U22903 ( .B1(n20009), .B2(n20008), .A(n20007), .ZN(P1_U2806) );
  NOR4_X1 U22904 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20013) );
  NOR4_X1 U22905 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20012) );
  NOR4_X1 U22906 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20011) );
  NOR4_X1 U22907 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20010) );
  NAND4_X1 U22908 ( .A1(n20013), .A2(n20012), .A3(n20011), .A4(n20010), .ZN(
        n20019) );
  NOR4_X1 U22909 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20017) );
  AOI211_X1 U22910 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20016) );
  NOR4_X1 U22911 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20015) );
  NOR4_X1 U22912 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20014) );
  NAND4_X1 U22913 ( .A1(n20017), .A2(n20016), .A3(n20015), .A4(n20014), .ZN(
        n20018) );
  NOR2_X1 U22914 ( .A1(n20019), .A2(n20018), .ZN(n20909) );
  INV_X1 U22915 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21068) );
  NOR3_X1 U22916 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20021) );
  OAI21_X1 U22917 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20021), .A(n20909), .ZN(
        n20020) );
  OAI21_X1 U22918 ( .B1(n20909), .B2(n21068), .A(n20020), .ZN(P1_U2807) );
  INV_X1 U22919 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20903) );
  AOI21_X1 U22920 ( .B1(n20855), .B2(n20903), .A(n20021), .ZN(n20022) );
  INV_X1 U22921 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21015) );
  INV_X1 U22922 ( .A(n20909), .ZN(n20907) );
  AOI22_X1 U22923 ( .A1(n20909), .A2(n20022), .B1(n21015), .B2(n20907), .ZN(
        P1_U2808) );
  AOI22_X1 U22924 ( .A1(n20089), .A2(n20024), .B1(n20023), .B2(n13869), .ZN(
        n20034) );
  OAI22_X1 U22925 ( .A1(n20026), .A2(n13869), .B1(n20025), .B2(n14519), .ZN(
        n20027) );
  AOI211_X1 U22926 ( .C1(n20091), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n20167), .B(n20027), .ZN(n20033) );
  OAI22_X1 U22927 ( .A1(n20030), .A2(n20029), .B1(n20078), .B2(n20028), .ZN(
        n20031) );
  INV_X1 U22928 ( .A(n20031), .ZN(n20032) );
  NAND3_X1 U22929 ( .A1(n20034), .A2(n20033), .A3(n20032), .ZN(P1_U2831) );
  NOR2_X1 U22930 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20044), .ZN(n20040) );
  AOI22_X1 U22931 ( .A1(n20089), .A2(n20035), .B1(n20088), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n20036) );
  OAI211_X1 U22932 ( .C1(n20067), .C2(n20037), .A(n20036), .B(n20064), .ZN(
        n20038) );
  AOI21_X1 U22933 ( .B1(n20040), .B2(n20039), .A(n20038), .ZN(n20048) );
  INV_X1 U22934 ( .A(n20041), .ZN(n20045) );
  OAI21_X1 U22935 ( .B1(n20043), .B2(n20052), .A(n20042), .ZN(n20082) );
  OAI21_X1 U22936 ( .B1(n20045), .B2(n20044), .A(n20082), .ZN(n20057) );
  AOI22_X1 U22937 ( .A1(n20046), .A2(n20058), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n20057), .ZN(n20047) );
  OAI211_X1 U22938 ( .C1(n20049), .C2(n20078), .A(n20048), .B(n20047), .ZN(
        P1_U2833) );
  NAND2_X1 U22939 ( .A1(n20051), .A2(n20050), .ZN(n20097) );
  NOR2_X1 U22940 ( .A1(n20052), .A2(n20097), .ZN(n20069) );
  NAND2_X1 U22941 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n20069), .ZN(n20055) );
  AOI22_X1 U22942 ( .A1(n20089), .A2(n20053), .B1(n20088), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n20054) );
  OAI21_X1 U22943 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n20055), .A(n20054), .ZN(
        n20056) );
  AOI211_X1 U22944 ( .C1(n20091), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20167), .B(n20056), .ZN(n20061) );
  AOI22_X1 U22945 ( .A1(n20059), .A2(n20058), .B1(P1_REIP_REG_6__SCAN_IN), 
        .B2(n20057), .ZN(n20060) );
  OAI211_X1 U22946 ( .C1(n20062), .C2(n20078), .A(n20061), .B(n20060), .ZN(
        P1_U2834) );
  INV_X1 U22947 ( .A(n20082), .ZN(n20070) );
  INV_X1 U22948 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20862) );
  AOI22_X1 U22949 ( .A1(n20089), .A2(n20063), .B1(n20088), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n20065) );
  OAI211_X1 U22950 ( .C1(n20067), .C2(n20066), .A(n20065), .B(n20064), .ZN(
        n20068) );
  AOI221_X1 U22951 ( .B1(n20070), .B2(P1_REIP_REG_5__SCAN_IN), .C1(n20069), 
        .C2(n20862), .A(n20068), .ZN(n20073) );
  NAND2_X1 U22952 ( .A1(n20071), .A2(n20099), .ZN(n20072) );
  OAI211_X1 U22953 ( .C1(n20078), .C2(n20074), .A(n20073), .B(n20072), .ZN(
        P1_U2835) );
  INV_X1 U22954 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20859) );
  NOR3_X1 U22955 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20859), .A3(n20097), .ZN(
        n20075) );
  AOI211_X1 U22956 ( .C1(n20091), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20167), .B(n20075), .ZN(n20085) );
  INV_X1 U22957 ( .A(n20076), .ZN(n20173) );
  INV_X1 U22958 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20857) );
  NAND2_X1 U22959 ( .A1(n20077), .A2(n20094), .ZN(n20081) );
  NOR2_X1 U22960 ( .A1(n20078), .A2(n20177), .ZN(n20079) );
  AOI21_X1 U22961 ( .B1(n20088), .B2(P1_EBX_REG_4__SCAN_IN), .A(n20079), .ZN(
        n20080) );
  OAI211_X1 U22962 ( .C1(n20857), .C2(n20082), .A(n20081), .B(n20080), .ZN(
        n20083) );
  AOI21_X1 U22963 ( .B1(n20173), .B2(n20099), .A(n20083), .ZN(n20084) );
  OAI211_X1 U22964 ( .C1(n20086), .C2(n20181), .A(n20085), .B(n20084), .ZN(
        P1_U2836) );
  INV_X1 U22965 ( .A(n20087), .ZN(n20191) );
  AOI22_X1 U22966 ( .A1(n20089), .A2(n20191), .B1(n20088), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n20102) );
  INV_X1 U22967 ( .A(n20090), .ZN(n20092) );
  AOI22_X1 U22968 ( .A1(n20093), .A2(n20092), .B1(n20091), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20096) );
  NAND2_X1 U22969 ( .A1(n13423), .A2(n20094), .ZN(n20095) );
  OAI211_X1 U22970 ( .C1(n20097), .C2(P1_REIP_REG_3__SCAN_IN), .A(n20096), .B(
        n20095), .ZN(n20098) );
  AOI21_X1 U22971 ( .B1(n20100), .B2(n20099), .A(n20098), .ZN(n20101) );
  OAI211_X1 U22972 ( .C1(n20859), .C2(n20103), .A(n20102), .B(n20101), .ZN(
        P1_U2837) );
  AOI22_X1 U22973 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20104) );
  OAI21_X1 U22974 ( .B1(n13252), .B2(n20127), .A(n20104), .ZN(P1_U2921) );
  INV_X1 U22975 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20106) );
  AOI22_X1 U22976 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20105) );
  OAI21_X1 U22977 ( .B1(n20106), .B2(n20127), .A(n20105), .ZN(P1_U2922) );
  AOI22_X1 U22978 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20107) );
  OAI21_X1 U22979 ( .B1(n14854), .B2(n20127), .A(n20107), .ZN(P1_U2923) );
  AOI22_X1 U22980 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20108) );
  OAI21_X1 U22981 ( .B1(n14029), .B2(n20127), .A(n20108), .ZN(P1_U2924) );
  AOI22_X1 U22982 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20109) );
  OAI21_X1 U22983 ( .B1(n13968), .B2(n20127), .A(n20109), .ZN(P1_U2925) );
  AOI22_X1 U22984 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20110) );
  OAI21_X1 U22985 ( .B1(n13866), .B2(n20127), .A(n20110), .ZN(P1_U2926) );
  AOI22_X1 U22986 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20111) );
  OAI21_X1 U22987 ( .B1(n13806), .B2(n20127), .A(n20111), .ZN(P1_U2927) );
  AOI22_X1 U22988 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20919), .B1(n15983), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20112) );
  OAI21_X1 U22989 ( .B1(n13705), .B2(n20127), .A(n20112), .ZN(P1_U2928) );
  AOI22_X1 U22990 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20125), .B1(n15983), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20113) );
  OAI21_X1 U22991 ( .B1(n10564), .B2(n20127), .A(n20113), .ZN(P1_U2929) );
  AOI22_X1 U22992 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20125), .B1(n15983), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20114) );
  OAI21_X1 U22993 ( .B1(n10546), .B2(n20127), .A(n20114), .ZN(P1_U2930) );
  AOI22_X1 U22994 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20125), .B1(n15983), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20115) );
  OAI21_X1 U22995 ( .B1(n20116), .B2(n20127), .A(n20115), .ZN(P1_U2931) );
  AOI22_X1 U22996 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20125), .B1(n15983), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20117) );
  OAI21_X1 U22997 ( .B1(n20118), .B2(n20127), .A(n20117), .ZN(P1_U2932) );
  AOI22_X1 U22998 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20125), .B1(n15983), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20119) );
  OAI21_X1 U22999 ( .B1(n20120), .B2(n20127), .A(n20119), .ZN(P1_U2933) );
  AOI22_X1 U23000 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20125), .B1(n15983), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20121) );
  OAI21_X1 U23001 ( .B1(n20122), .B2(n20127), .A(n20121), .ZN(P1_U2934) );
  AOI22_X1 U23002 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20125), .B1(n15983), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20123) );
  OAI21_X1 U23003 ( .B1(n20124), .B2(n20127), .A(n20123), .ZN(P1_U2935) );
  AOI22_X1 U23004 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20125), .B1(n15983), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20126) );
  OAI21_X1 U23005 ( .B1(n20128), .B2(n20127), .A(n20126), .ZN(P1_U2936) );
  AOI22_X1 U23006 ( .A1(n20164), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20135), .ZN(n20131) );
  INV_X1 U23007 ( .A(n20129), .ZN(n20130) );
  NAND2_X1 U23008 ( .A1(n20149), .A2(n20130), .ZN(n20151) );
  NAND2_X1 U23009 ( .A1(n20131), .A2(n20151), .ZN(P1_U2945) );
  AOI22_X1 U23010 ( .A1(n20164), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20135), .ZN(n20134) );
  INV_X1 U23011 ( .A(n20132), .ZN(n20133) );
  NAND2_X1 U23012 ( .A1(n20149), .A2(n20133), .ZN(n20153) );
  NAND2_X1 U23013 ( .A1(n20134), .A2(n20153), .ZN(P1_U2946) );
  AOI22_X1 U23014 ( .A1(n20164), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20135), .ZN(n20138) );
  INV_X1 U23015 ( .A(n20136), .ZN(n20137) );
  NAND2_X1 U23016 ( .A1(n20149), .A2(n20137), .ZN(n20155) );
  NAND2_X1 U23017 ( .A1(n20138), .A2(n20155), .ZN(P1_U2947) );
  AOI22_X1 U23018 ( .A1(n20164), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20159), .ZN(n20141) );
  INV_X1 U23019 ( .A(n20139), .ZN(n20140) );
  NAND2_X1 U23020 ( .A1(n20149), .A2(n20140), .ZN(n20157) );
  NAND2_X1 U23021 ( .A1(n20141), .A2(n20157), .ZN(P1_U2948) );
  AOI22_X1 U23022 ( .A1(n20164), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20159), .ZN(n20144) );
  INV_X1 U23023 ( .A(n20142), .ZN(n20143) );
  NAND2_X1 U23024 ( .A1(n20149), .A2(n20143), .ZN(n20160) );
  NAND2_X1 U23025 ( .A1(n20144), .A2(n20160), .ZN(P1_U2949) );
  AOI22_X1 U23026 ( .A1(n20164), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20159), .ZN(n20147) );
  INV_X1 U23027 ( .A(n20145), .ZN(n20146) );
  NAND2_X1 U23028 ( .A1(n20149), .A2(n20146), .ZN(n20162) );
  NAND2_X1 U23029 ( .A1(n20147), .A2(n20162), .ZN(P1_U2950) );
  AOI22_X1 U23030 ( .A1(n20164), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20159), .ZN(n20150) );
  NAND2_X1 U23031 ( .A1(n20149), .A2(n20148), .ZN(n20165) );
  NAND2_X1 U23032 ( .A1(n20150), .A2(n20165), .ZN(P1_U2951) );
  AOI22_X1 U23033 ( .A1(n20164), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20159), .ZN(n20152) );
  NAND2_X1 U23034 ( .A1(n20152), .A2(n20151), .ZN(P1_U2960) );
  AOI22_X1 U23035 ( .A1(n20164), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20159), .ZN(n20154) );
  NAND2_X1 U23036 ( .A1(n20154), .A2(n20153), .ZN(P1_U2961) );
  AOI22_X1 U23037 ( .A1(n20164), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20159), .ZN(n20156) );
  NAND2_X1 U23038 ( .A1(n20156), .A2(n20155), .ZN(P1_U2962) );
  AOI22_X1 U23039 ( .A1(n20164), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20159), .ZN(n20158) );
  NAND2_X1 U23040 ( .A1(n20158), .A2(n20157), .ZN(P1_U2963) );
  AOI22_X1 U23041 ( .A1(n20164), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20159), .ZN(n20161) );
  NAND2_X1 U23042 ( .A1(n20161), .A2(n20160), .ZN(P1_U2964) );
  AOI22_X1 U23043 ( .A1(n20164), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20159), .ZN(n20163) );
  NAND2_X1 U23044 ( .A1(n20163), .A2(n20162), .ZN(P1_U2965) );
  AOI22_X1 U23045 ( .A1(n20164), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20135), .ZN(n20166) );
  NAND2_X1 U23046 ( .A1(n20166), .A2(n20165), .ZN(P1_U2966) );
  AOI22_X1 U23047 ( .A1(n20168), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20167), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20176) );
  OAI21_X1 U23048 ( .B1(n20171), .B2(n20170), .A(n20169), .ZN(n20172) );
  INV_X1 U23049 ( .A(n20172), .ZN(n20184) );
  AOI22_X1 U23050 ( .A1(n20184), .A2(n20174), .B1(n20239), .B2(n20173), .ZN(
        n20175) );
  OAI211_X1 U23051 ( .C1(n20178), .C2(n20177), .A(n20176), .B(n20175), .ZN(
        P1_U2995) );
  INV_X1 U23052 ( .A(n20179), .ZN(n20180) );
  AOI21_X1 U23053 ( .B1(n20209), .B2(n20208), .A(n20180), .ZN(n20198) );
  OAI22_X1 U23054 ( .A1(n20182), .A2(n20181), .B1(n20857), .B2(n20225), .ZN(
        n20183) );
  AOI21_X1 U23055 ( .B1(n20184), .B2(n20206), .A(n20183), .ZN(n20187) );
  OAI211_X1 U23056 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20193), .B(n20185), .ZN(n20186) );
  OAI211_X1 U23057 ( .C1(n20198), .C2(n20188), .A(n20187), .B(n20186), .ZN(
        P1_U3027) );
  INV_X1 U23058 ( .A(n20189), .ZN(n20190) );
  AOI21_X1 U23059 ( .B1(n20228), .B2(n20191), .A(n20190), .ZN(n20196) );
  INV_X1 U23060 ( .A(n20192), .ZN(n20194) );
  AOI22_X1 U23061 ( .A1(n20194), .A2(n20206), .B1(n20197), .B2(n20193), .ZN(
        n20195) );
  OAI211_X1 U23062 ( .C1(n20198), .C2(n20197), .A(n20196), .B(n20195), .ZN(
        P1_U3028) );
  INV_X1 U23063 ( .A(n20199), .ZN(n20202) );
  INV_X1 U23064 ( .A(n20200), .ZN(n20201) );
  AOI21_X1 U23065 ( .B1(n20228), .B2(n20202), .A(n20201), .ZN(n20218) );
  INV_X1 U23066 ( .A(n20203), .ZN(n20207) );
  AOI22_X1 U23067 ( .A1(n20207), .A2(n20206), .B1(n20205), .B2(n20204), .ZN(
        n20217) );
  NAND2_X1 U23068 ( .A1(n20209), .A2(n20208), .ZN(n20216) );
  NAND2_X1 U23069 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20211) );
  OAI22_X1 U23070 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20212), .B1(
        n20211), .B2(n20210), .ZN(n20213) );
  OAI21_X1 U23071 ( .B1(n20214), .B2(n20213), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20215) );
  NAND4_X1 U23072 ( .A1(n20218), .A2(n20217), .A3(n20216), .A4(n20215), .ZN(
        P1_U3029) );
  NAND2_X1 U23073 ( .A1(n20220), .A2(n20219), .ZN(n20234) );
  INV_X1 U23074 ( .A(n20221), .ZN(n20224) );
  OR3_X1 U23075 ( .A1(n20224), .A2(n20223), .A3(n20222), .ZN(n20230) );
  NOR2_X1 U23076 ( .A1(n20225), .A2(n20855), .ZN(n20226) );
  AOI21_X1 U23077 ( .B1(n20228), .B2(n20227), .A(n20226), .ZN(n20229) );
  AND2_X1 U23078 ( .A1(n20230), .A2(n20229), .ZN(n20231) );
  OAI221_X1 U23079 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20234), .C1(
        n20233), .C2(n20232), .A(n20231), .ZN(P1_U3030) );
  NOR2_X1 U23080 ( .A1(n20236), .A2(n20235), .ZN(P1_U3032) );
  NAND2_X1 U23081 ( .A1(n20237), .A2(n20239), .ZN(n20288) );
  INV_X1 U23082 ( .A(n20288), .ZN(n20285) );
  NAND2_X1 U23083 ( .A1(n20239), .A2(n20238), .ZN(n20286) );
  INV_X1 U23084 ( .A(n20286), .ZN(n20284) );
  INV_X1 U23085 ( .A(n20326), .ZN(n20241) );
  INV_X1 U23086 ( .A(n20621), .ZN(n20242) );
  AOI22_X1 U23087 ( .A1(DATAI_24_), .A2(n20285), .B1(BUF1_REG_24__SCAN_IN), 
        .B2(n20284), .ZN(n20787) );
  INV_X1 U23088 ( .A(n20787), .ZN(n20731) );
  NAND3_X1 U23089 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20914), .A3(n20243), 
        .ZN(n20275) );
  NAND2_X1 U23090 ( .A1(n20290), .A2(n20244), .ZN(n20647) );
  NOR3_X1 U23091 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20303) );
  INV_X1 U23092 ( .A(n20303), .ZN(n20298) );
  NOR2_X1 U23093 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20298), .ZN(
        n20291) );
  AOI22_X1 U23094 ( .A1(n20829), .A2(n20731), .B1(n20774), .B2(n20291), .ZN(
        n20256) );
  INV_X1 U23095 ( .A(n20252), .ZN(n20245) );
  NOR2_X1 U23096 ( .A1(n20245), .A2(n20837), .ZN(n20400) );
  NOR3_X1 U23097 ( .A1(n20314), .A2(n20829), .A3(n20781), .ZN(n20246) );
  NOR2_X1 U23098 ( .A1(n20246), .A2(n20328), .ZN(n20254) );
  INV_X1 U23099 ( .A(n20254), .ZN(n20249) );
  OR2_X1 U23100 ( .A1(n13423), .A2(n20247), .ZN(n20331) );
  OR2_X1 U23101 ( .A1(n20331), .A2(n9665), .ZN(n20253) );
  INV_X1 U23102 ( .A(n20520), .ZN(n20248) );
  NAND2_X1 U23103 ( .A1(n20248), .A2(n20575), .ZN(n20403) );
  AOI22_X1 U23104 ( .A1(n20249), .A2(n20253), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20403), .ZN(n20250) );
  NOR2_X2 U23105 ( .A1(n20251), .A2(n20299), .ZN(n20773) );
  OR2_X1 U23106 ( .A1(n20252), .A2(n20837), .ZN(n20579) );
  OAI22_X1 U23107 ( .A1(n20254), .A2(n20253), .B1(n20579), .B2(n20403), .ZN(
        n20293) );
  AOI22_X1 U23108 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20294), .B1(
        n20773), .B2(n20293), .ZN(n20255) );
  OAI211_X1 U23109 ( .C1(n20734), .C2(n20325), .A(n20256), .B(n20255), .ZN(
        P1_U3033) );
  INV_X1 U23110 ( .A(DATAI_17_), .ZN(n20932) );
  OAI22_X1 U23111 ( .A1(n20257), .A2(n20286), .B1(n20932), .B2(n20288), .ZN(
        n20790) );
  INV_X1 U23112 ( .A(n20790), .ZN(n20738) );
  AOI22_X1 U23113 ( .A1(DATAI_25_), .A2(n20285), .B1(BUF1_REG_25__SCAN_IN), 
        .B2(n20284), .ZN(n20793) );
  INV_X1 U23114 ( .A(n20793), .ZN(n20735) );
  NAND2_X1 U23115 ( .A1(n20290), .A2(n20258), .ZN(n20660) );
  AOI22_X1 U23116 ( .A1(n20829), .A2(n20735), .B1(n20789), .B2(n20291), .ZN(
        n20261) );
  NOR2_X2 U23117 ( .A1(n20259), .A2(n20299), .ZN(n20788) );
  AOI22_X1 U23118 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20294), .B1(
        n20788), .B2(n20293), .ZN(n20260) );
  OAI211_X1 U23119 ( .C1(n20738), .C2(n20325), .A(n20261), .B(n20260), .ZN(
        P1_U3034) );
  AOI22_X1 U23120 ( .A1(DATAI_18_), .A2(n20285), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20284), .ZN(n20742) );
  INV_X1 U23121 ( .A(DATAI_26_), .ZN(n20936) );
  OAI22_X1 U23122 ( .A1(n20262), .A2(n20286), .B1(n20936), .B2(n20288), .ZN(
        n20739) );
  NAND2_X1 U23123 ( .A1(n20290), .A2(n20263), .ZN(n20664) );
  AOI22_X1 U23124 ( .A1(n20829), .A2(n20739), .B1(n20795), .B2(n20291), .ZN(
        n20266) );
  NOR2_X2 U23125 ( .A1(n20264), .A2(n20299), .ZN(n20794) );
  AOI22_X1 U23126 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20294), .B1(
        n20794), .B2(n20293), .ZN(n20265) );
  OAI211_X1 U23127 ( .C1(n20742), .C2(n20325), .A(n20266), .B(n20265), .ZN(
        P1_U3035) );
  INV_X1 U23128 ( .A(DATAI_27_), .ZN(n21014) );
  OAI22_X1 U23129 ( .A1(n15329), .A2(n20286), .B1(n21014), .B2(n20288), .ZN(
        n20743) );
  NAND2_X1 U23130 ( .A1(n20290), .A2(n20267), .ZN(n20668) );
  AOI22_X1 U23131 ( .A1(n20829), .A2(n20743), .B1(n20801), .B2(n20291), .ZN(
        n20270) );
  NOR2_X2 U23132 ( .A1(n20268), .A2(n20299), .ZN(n20800) );
  AOI22_X1 U23133 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20294), .B1(
        n20800), .B2(n20293), .ZN(n20269) );
  OAI211_X1 U23134 ( .C1(n20746), .C2(n20325), .A(n20270), .B(n20269), .ZN(
        P1_U3036) );
  AOI22_X1 U23135 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20284), .B1(DATAI_20_), 
        .B2(n20285), .ZN(n20750) );
  INV_X1 U23136 ( .A(DATAI_28_), .ZN(n21037) );
  OAI22_X1 U23137 ( .A1(n15322), .A2(n20286), .B1(n21037), .B2(n20288), .ZN(
        n20747) );
  NAND2_X1 U23138 ( .A1(n20290), .A2(n20271), .ZN(n20672) );
  AOI22_X1 U23139 ( .A1(n20829), .A2(n20747), .B1(n20807), .B2(n20291), .ZN(
        n20274) );
  NOR2_X2 U23140 ( .A1(n20299), .A2(n20272), .ZN(n20806) );
  AOI22_X1 U23141 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20294), .B1(
        n20806), .B2(n20293), .ZN(n20273) );
  OAI211_X1 U23142 ( .C1(n20750), .C2(n20325), .A(n20274), .B(n20273), .ZN(
        P1_U3037) );
  AOI22_X1 U23143 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20284), .B1(DATAI_21_), 
        .B2(n20285), .ZN(n20754) );
  INV_X1 U23144 ( .A(DATAI_29_), .ZN(n20928) );
  OAI22_X1 U23145 ( .A1(n15317), .A2(n20286), .B1(n20928), .B2(n20288), .ZN(
        n20751) );
  NOR2_X2 U23146 ( .A1(n20275), .A2(n10304), .ZN(n20812) );
  AOI22_X1 U23147 ( .A1(n20829), .A2(n20751), .B1(n20812), .B2(n20291), .ZN(
        n20278) );
  NOR2_X2 U23148 ( .A1(n20299), .A2(n20276), .ZN(n20813) );
  AOI22_X1 U23149 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20294), .B1(
        n20813), .B2(n20293), .ZN(n20277) );
  OAI211_X1 U23150 ( .C1(n20754), .C2(n20325), .A(n20278), .B(n20277), .ZN(
        P1_U3038) );
  INV_X1 U23151 ( .A(DATAI_22_), .ZN(n20930) );
  OAI22_X1 U23152 ( .A1(n20279), .A2(n20286), .B1(n20930), .B2(n20288), .ZN(
        n20820) );
  INV_X1 U23153 ( .A(n20820), .ZN(n20758) );
  INV_X1 U23154 ( .A(n20823), .ZN(n20755) );
  NAND2_X1 U23155 ( .A1(n20290), .A2(n20280), .ZN(n20680) );
  AOI22_X1 U23156 ( .A1(n20829), .A2(n20755), .B1(n20819), .B2(n20291), .ZN(
        n20283) );
  NOR2_X2 U23157 ( .A1(n20299), .A2(n20281), .ZN(n20818) );
  AOI22_X1 U23158 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20294), .B1(
        n20818), .B2(n20293), .ZN(n20282) );
  OAI211_X1 U23159 ( .C1(n20758), .C2(n20325), .A(n20283), .B(n20282), .ZN(
        P1_U3039) );
  AOI22_X1 U23160 ( .A1(DATAI_23_), .A2(n20285), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n20284), .ZN(n20766) );
  INV_X1 U23161 ( .A(DATAI_31_), .ZN(n21038) );
  OAI22_X1 U23162 ( .A1(n21038), .A2(n20288), .B1(n20287), .B2(n20286), .ZN(
        n20761) );
  NAND2_X1 U23163 ( .A1(n20290), .A2(n20289), .ZN(n20685) );
  AOI22_X1 U23164 ( .A1(n20829), .A2(n20761), .B1(n20827), .B2(n20291), .ZN(
        n20296) );
  NOR2_X2 U23165 ( .A1(n20299), .A2(n20292), .ZN(n20825) );
  AOI22_X1 U23166 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20294), .B1(
        n20825), .B2(n20293), .ZN(n20295) );
  OAI211_X1 U23167 ( .C1(n20766), .C2(n20325), .A(n20296), .B(n20295), .ZN(
        P1_U3040) );
  NOR2_X1 U23168 ( .A1(n20692), .A2(n20298), .ZN(n20320) );
  INV_X1 U23169 ( .A(n20331), .ZN(n20367) );
  INV_X1 U23170 ( .A(n20297), .ZN(n20693) );
  AOI21_X1 U23171 ( .B1(n20367), .B2(n20693), .A(n20320), .ZN(n20300) );
  OAI22_X1 U23172 ( .A1(n20300), .A2(n20781), .B1(n20298), .B2(n20837), .ZN(
        n20319) );
  AOI22_X1 U23173 ( .A1(n20774), .A2(n20320), .B1(n20773), .B2(n20319), .ZN(
        n20305) );
  INV_X1 U23174 ( .A(n20369), .ZN(n20301) );
  OAI211_X1 U23175 ( .C1(n20301), .C2(n20548), .A(n20783), .B(n20300), .ZN(
        n20302) );
  OAI211_X1 U23176 ( .C1(n20783), .C2(n20303), .A(n20779), .B(n20302), .ZN(
        n20322) );
  INV_X1 U23177 ( .A(n20364), .ZN(n20321) );
  INV_X1 U23178 ( .A(n20734), .ZN(n20784) );
  AOI22_X1 U23179 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20322), .B1(
        n20321), .B2(n20784), .ZN(n20304) );
  OAI211_X1 U23180 ( .C1(n20787), .C2(n20325), .A(n20305), .B(n20304), .ZN(
        P1_U3041) );
  AOI22_X1 U23181 ( .A1(n20789), .A2(n20320), .B1(n20788), .B2(n20319), .ZN(
        n20307) );
  AOI22_X1 U23182 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20322), .B1(
        n20321), .B2(n20790), .ZN(n20306) );
  OAI211_X1 U23183 ( .C1(n20793), .C2(n20325), .A(n20307), .B(n20306), .ZN(
        P1_U3042) );
  AOI22_X1 U23184 ( .A1(n20795), .A2(n20320), .B1(n20794), .B2(n20319), .ZN(
        n20309) );
  AOI22_X1 U23185 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20322), .B1(
        n20314), .B2(n20739), .ZN(n20308) );
  OAI211_X1 U23186 ( .C1(n20742), .C2(n20364), .A(n20309), .B(n20308), .ZN(
        P1_U3043) );
  AOI22_X1 U23187 ( .A1(n20801), .A2(n20320), .B1(n20800), .B2(n20319), .ZN(
        n20311) );
  AOI22_X1 U23188 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20322), .B1(
        n20314), .B2(n20743), .ZN(n20310) );
  OAI211_X1 U23189 ( .C1(n20746), .C2(n20364), .A(n20311), .B(n20310), .ZN(
        P1_U3044) );
  INV_X1 U23190 ( .A(n20747), .ZN(n20811) );
  AOI22_X1 U23191 ( .A1(n20807), .A2(n20320), .B1(n20806), .B2(n20319), .ZN(
        n20313) );
  INV_X1 U23192 ( .A(n20750), .ZN(n20808) );
  AOI22_X1 U23193 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20322), .B1(
        n20321), .B2(n20808), .ZN(n20312) );
  OAI211_X1 U23194 ( .C1(n20811), .C2(n20325), .A(n20313), .B(n20312), .ZN(
        P1_U3045) );
  AOI22_X1 U23195 ( .A1(n20813), .A2(n20319), .B1(n20812), .B2(n20320), .ZN(
        n20316) );
  AOI22_X1 U23196 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20322), .B1(
        n20314), .B2(n20751), .ZN(n20315) );
  OAI211_X1 U23197 ( .C1(n20754), .C2(n20364), .A(n20316), .B(n20315), .ZN(
        P1_U3046) );
  AOI22_X1 U23198 ( .A1(n20819), .A2(n20320), .B1(n20818), .B2(n20319), .ZN(
        n20318) );
  AOI22_X1 U23199 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20322), .B1(
        n20321), .B2(n20820), .ZN(n20317) );
  OAI211_X1 U23200 ( .C1(n20823), .C2(n20325), .A(n20318), .B(n20317), .ZN(
        P1_U3047) );
  INV_X1 U23201 ( .A(n20761), .ZN(n20834) );
  AOI22_X1 U23202 ( .A1(n20827), .A2(n20320), .B1(n20825), .B2(n20319), .ZN(
        n20324) );
  INV_X1 U23203 ( .A(n20766), .ZN(n20828) );
  AOI22_X1 U23204 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20322), .B1(
        n20321), .B2(n20828), .ZN(n20323) );
  OAI211_X1 U23205 ( .C1(n20834), .C2(n20325), .A(n20324), .B(n20323), .ZN(
        P1_U3048) );
  NAND3_X1 U23206 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20645), .A3(
        n20646), .ZN(n20372) );
  NOR2_X1 U23207 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20372), .ZN(
        n20351) );
  INV_X1 U23208 ( .A(n20351), .ZN(n20358) );
  OAI22_X1 U23209 ( .A1(n20364), .A2(n20787), .B1(n20358), .B2(n20647), .ZN(
        n20327) );
  INV_X1 U23210 ( .A(n20327), .ZN(n20338) );
  NAND3_X1 U23211 ( .A1(n20394), .A2(n20364), .A3(n20783), .ZN(n20330) );
  INV_X1 U23212 ( .A(n20328), .ZN(n20329) );
  NAND2_X1 U23213 ( .A1(n20330), .A2(n20329), .ZN(n20333) );
  OR2_X1 U23214 ( .A1(n20331), .A2(n20651), .ZN(n20335) );
  AOI22_X1 U23215 ( .A1(n20333), .A2(n20335), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20358), .ZN(n20332) );
  OAI21_X1 U23216 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20575), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20457) );
  NAND3_X1 U23217 ( .A1(n20577), .A2(n20332), .A3(n20457), .ZN(n20361) );
  INV_X1 U23218 ( .A(n20333), .ZN(n20336) );
  INV_X1 U23219 ( .A(n20575), .ZN(n20334) );
  NAND2_X1 U23220 ( .A1(n20334), .A2(n20645), .ZN(n20460) );
  OAI22_X1 U23221 ( .A1(n20336), .A2(n20335), .B1(n20579), .B2(n20460), .ZN(
        n20360) );
  AOI22_X1 U23222 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20361), .B1(
        n20773), .B2(n20360), .ZN(n20337) );
  OAI211_X1 U23223 ( .C1(n20734), .C2(n20394), .A(n20338), .B(n20337), .ZN(
        P1_U3049) );
  OAI22_X1 U23224 ( .A1(n20364), .A2(n20793), .B1(n20358), .B2(n20660), .ZN(
        n20339) );
  INV_X1 U23225 ( .A(n20339), .ZN(n20341) );
  AOI22_X1 U23226 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20361), .B1(
        n20788), .B2(n20360), .ZN(n20340) );
  OAI211_X1 U23227 ( .C1(n20738), .C2(n20394), .A(n20341), .B(n20340), .ZN(
        P1_U3050) );
  INV_X1 U23228 ( .A(n20739), .ZN(n20799) );
  OAI22_X1 U23229 ( .A1(n20394), .A2(n20742), .B1(n20664), .B2(n20358), .ZN(
        n20342) );
  INV_X1 U23230 ( .A(n20342), .ZN(n20344) );
  AOI22_X1 U23231 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20361), .B1(
        n20794), .B2(n20360), .ZN(n20343) );
  OAI211_X1 U23232 ( .C1(n20799), .C2(n20364), .A(n20344), .B(n20343), .ZN(
        P1_U3051) );
  INV_X1 U23233 ( .A(n20743), .ZN(n20805) );
  OAI22_X1 U23234 ( .A1(n20394), .A2(n20746), .B1(n20358), .B2(n20668), .ZN(
        n20345) );
  INV_X1 U23235 ( .A(n20345), .ZN(n20347) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20361), .B1(
        n20800), .B2(n20360), .ZN(n20346) );
  OAI211_X1 U23237 ( .C1(n20805), .C2(n20364), .A(n20347), .B(n20346), .ZN(
        P1_U3052) );
  OAI22_X1 U23238 ( .A1(n20394), .A2(n20750), .B1(n20672), .B2(n20358), .ZN(
        n20348) );
  INV_X1 U23239 ( .A(n20348), .ZN(n20350) );
  AOI22_X1 U23240 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20361), .B1(
        n20806), .B2(n20360), .ZN(n20349) );
  OAI211_X1 U23241 ( .C1(n20811), .C2(n20364), .A(n20350), .B(n20349), .ZN(
        P1_U3053) );
  INV_X1 U23242 ( .A(n20751), .ZN(n20817) );
  INV_X1 U23243 ( .A(n20394), .ZN(n20352) );
  INV_X1 U23244 ( .A(n20754), .ZN(n20814) );
  AOI22_X1 U23245 ( .A1(n20352), .A2(n20814), .B1(n20812), .B2(n20351), .ZN(
        n20354) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20361), .B1(
        n20813), .B2(n20360), .ZN(n20353) );
  OAI211_X1 U23247 ( .C1(n20817), .C2(n20364), .A(n20354), .B(n20353), .ZN(
        P1_U3054) );
  OAI22_X1 U23248 ( .A1(n20364), .A2(n20823), .B1(n20358), .B2(n20680), .ZN(
        n20355) );
  INV_X1 U23249 ( .A(n20355), .ZN(n20357) );
  AOI22_X1 U23250 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20361), .B1(
        n20818), .B2(n20360), .ZN(n20356) );
  OAI211_X1 U23251 ( .C1(n20758), .C2(n20394), .A(n20357), .B(n20356), .ZN(
        P1_U3055) );
  OAI22_X1 U23252 ( .A1(n20394), .A2(n20766), .B1(n20358), .B2(n20685), .ZN(
        n20359) );
  INV_X1 U23253 ( .A(n20359), .ZN(n20363) );
  AOI22_X1 U23254 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20361), .B1(
        n20825), .B2(n20360), .ZN(n20362) );
  OAI211_X1 U23255 ( .C1(n20834), .C2(n20364), .A(n20363), .B(n20362), .ZN(
        P1_U3056) );
  OR2_X1 U23256 ( .A1(n20610), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20393) );
  OAI22_X1 U23257 ( .A1(n20394), .A2(n20787), .B1(n20393), .B2(n20647), .ZN(
        n20365) );
  INV_X1 U23258 ( .A(n20365), .ZN(n20376) );
  AND2_X1 U23259 ( .A1(n9645), .A2(n10445), .ZN(n20767) );
  INV_X1 U23260 ( .A(n20393), .ZN(n20387) );
  AOI21_X1 U23261 ( .B1(n20367), .B2(n20767), .A(n20387), .ZN(n20374) );
  AOI21_X1 U23262 ( .B1(n20369), .B2(n20368), .A(n20781), .ZN(n20371) );
  AOI22_X1 U23263 ( .A1(n20374), .A2(n20371), .B1(n20781), .B2(n20372), .ZN(
        n20370) );
  NAND2_X1 U23264 ( .A1(n20779), .A2(n20370), .ZN(n20397) );
  INV_X1 U23265 ( .A(n20371), .ZN(n20373) );
  OAI22_X1 U23266 ( .A1(n20374), .A2(n20373), .B1(n20837), .B2(n20372), .ZN(
        n20396) );
  AOI22_X1 U23267 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20397), .B1(
        n20773), .B2(n20396), .ZN(n20375) );
  OAI211_X1 U23268 ( .C1(n20734), .C2(n20428), .A(n20376), .B(n20375), .ZN(
        P1_U3057) );
  OAI22_X1 U23269 ( .A1(n20394), .A2(n20793), .B1(n20393), .B2(n20660), .ZN(
        n20377) );
  INV_X1 U23270 ( .A(n20377), .ZN(n20379) );
  AOI22_X1 U23271 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20397), .B1(
        n20788), .B2(n20396), .ZN(n20378) );
  OAI211_X1 U23272 ( .C1(n20738), .C2(n20428), .A(n20379), .B(n20378), .ZN(
        P1_U3058) );
  INV_X1 U23273 ( .A(n20742), .ZN(n20796) );
  AOI22_X1 U23274 ( .A1(n20420), .A2(n20796), .B1(n20795), .B2(n20387), .ZN(
        n20381) );
  AOI22_X1 U23275 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20397), .B1(
        n20794), .B2(n20396), .ZN(n20380) );
  OAI211_X1 U23276 ( .C1(n20799), .C2(n20394), .A(n20381), .B(n20380), .ZN(
        P1_U3059) );
  OAI22_X1 U23277 ( .A1(n20394), .A2(n20805), .B1(n20393), .B2(n20668), .ZN(
        n20382) );
  INV_X1 U23278 ( .A(n20382), .ZN(n20384) );
  AOI22_X1 U23279 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20397), .B1(
        n20800), .B2(n20396), .ZN(n20383) );
  OAI211_X1 U23280 ( .C1(n20746), .C2(n20428), .A(n20384), .B(n20383), .ZN(
        P1_U3060) );
  AOI22_X1 U23281 ( .A1(n20420), .A2(n20808), .B1(n20807), .B2(n20387), .ZN(
        n20386) );
  AOI22_X1 U23282 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20397), .B1(
        n20806), .B2(n20396), .ZN(n20385) );
  OAI211_X1 U23283 ( .C1(n20811), .C2(n20394), .A(n20386), .B(n20385), .ZN(
        P1_U3061) );
  AOI22_X1 U23284 ( .A1(n20420), .A2(n20814), .B1(n20387), .B2(n20812), .ZN(
        n20389) );
  AOI22_X1 U23285 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20397), .B1(
        n20813), .B2(n20396), .ZN(n20388) );
  OAI211_X1 U23286 ( .C1(n20817), .C2(n20394), .A(n20389), .B(n20388), .ZN(
        P1_U3062) );
  OAI22_X1 U23287 ( .A1(n20394), .A2(n20823), .B1(n20393), .B2(n20680), .ZN(
        n20390) );
  INV_X1 U23288 ( .A(n20390), .ZN(n20392) );
  AOI22_X1 U23289 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20397), .B1(
        n20818), .B2(n20396), .ZN(n20391) );
  OAI211_X1 U23290 ( .C1(n20758), .C2(n20428), .A(n20392), .B(n20391), .ZN(
        P1_U3063) );
  OAI22_X1 U23291 ( .A1(n20394), .A2(n20834), .B1(n20393), .B2(n20685), .ZN(
        n20395) );
  INV_X1 U23292 ( .A(n20395), .ZN(n20399) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20397), .B1(
        n20825), .B2(n20396), .ZN(n20398) );
  OAI211_X1 U23294 ( .C1(n20766), .C2(n20428), .A(n20399), .B(n20398), .ZN(
        P1_U3064) );
  NOR3_X1 U23295 ( .A1(n20646), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20433) );
  INV_X1 U23296 ( .A(n20433), .ZN(n20429) );
  NOR2_X1 U23297 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20429), .ZN(
        n20424) );
  INV_X1 U23298 ( .A(n20400), .ZN(n20723) );
  NOR2_X1 U23299 ( .A1(n13416), .A2(n20401), .ZN(n20491) );
  NAND3_X1 U23300 ( .A1(n20491), .A2(n20783), .A3(n20651), .ZN(n20402) );
  OAI21_X1 U23301 ( .B1(n20403), .B2(n20723), .A(n20402), .ZN(n20423) );
  AOI22_X1 U23302 ( .A1(n20774), .A2(n20424), .B1(n20773), .B2(n20423), .ZN(
        n20409) );
  INV_X1 U23303 ( .A(n20491), .ZN(n20405) );
  OAI21_X1 U23304 ( .B1(n20420), .B2(n20451), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20404) );
  OAI21_X1 U23305 ( .B1(n9665), .B2(n20405), .A(n20404), .ZN(n20407) );
  OAI221_X1 U23306 ( .B1(n20424), .B2(n20525), .C1(n20424), .C2(n20407), .A(
        n20729), .ZN(n20425) );
  AOI22_X1 U23307 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20425), .B1(
        n20420), .B2(n20731), .ZN(n20408) );
  OAI211_X1 U23308 ( .C1(n20734), .C2(n20448), .A(n20409), .B(n20408), .ZN(
        P1_U3065) );
  AOI22_X1 U23309 ( .A1(n20789), .A2(n20424), .B1(n20788), .B2(n20423), .ZN(
        n20411) );
  AOI22_X1 U23310 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20425), .B1(
        n20420), .B2(n20735), .ZN(n20410) );
  OAI211_X1 U23311 ( .C1(n20738), .C2(n20448), .A(n20411), .B(n20410), .ZN(
        P1_U3066) );
  AOI22_X1 U23312 ( .A1(n20795), .A2(n20424), .B1(n20794), .B2(n20423), .ZN(
        n20413) );
  AOI22_X1 U23313 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20425), .B1(
        n20451), .B2(n20796), .ZN(n20412) );
  OAI211_X1 U23314 ( .C1(n20799), .C2(n20428), .A(n20413), .B(n20412), .ZN(
        P1_U3067) );
  AOI22_X1 U23315 ( .A1(n20801), .A2(n20424), .B1(n20800), .B2(n20423), .ZN(
        n20415) );
  INV_X1 U23316 ( .A(n20746), .ZN(n20802) );
  AOI22_X1 U23317 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20425), .B1(
        n20451), .B2(n20802), .ZN(n20414) );
  OAI211_X1 U23318 ( .C1(n20805), .C2(n20428), .A(n20415), .B(n20414), .ZN(
        P1_U3068) );
  AOI22_X1 U23319 ( .A1(n20807), .A2(n20424), .B1(n20806), .B2(n20423), .ZN(
        n20417) );
  AOI22_X1 U23320 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20425), .B1(
        n20451), .B2(n20808), .ZN(n20416) );
  OAI211_X1 U23321 ( .C1(n20811), .C2(n20428), .A(n20417), .B(n20416), .ZN(
        P1_U3069) );
  AOI22_X1 U23322 ( .A1(n20813), .A2(n20423), .B1(n20812), .B2(n20424), .ZN(
        n20419) );
  AOI22_X1 U23323 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20425), .B1(
        n20451), .B2(n20814), .ZN(n20418) );
  OAI211_X1 U23324 ( .C1(n20817), .C2(n20428), .A(n20419), .B(n20418), .ZN(
        P1_U3070) );
  AOI22_X1 U23325 ( .A1(n20819), .A2(n20424), .B1(n20818), .B2(n20423), .ZN(
        n20422) );
  AOI22_X1 U23326 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20425), .B1(
        n20420), .B2(n20755), .ZN(n20421) );
  OAI211_X1 U23327 ( .C1(n20758), .C2(n20448), .A(n20422), .B(n20421), .ZN(
        P1_U3071) );
  AOI22_X1 U23328 ( .A1(n20827), .A2(n20424), .B1(n20825), .B2(n20423), .ZN(
        n20427) );
  AOI22_X1 U23329 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20425), .B1(
        n20451), .B2(n20828), .ZN(n20426) );
  OAI211_X1 U23330 ( .C1(n20834), .C2(n20428), .A(n20427), .B(n20426), .ZN(
        P1_U3072) );
  NOR2_X1 U23331 ( .A1(n20692), .A2(n20429), .ZN(n20450) );
  AOI21_X1 U23332 ( .B1(n20491), .B2(n20693), .A(n20450), .ZN(n20430) );
  OAI22_X1 U23333 ( .A1(n20430), .A2(n20781), .B1(n20429), .B2(n20837), .ZN(
        n20449) );
  AOI22_X1 U23334 ( .A1(n20774), .A2(n20450), .B1(n20773), .B2(n20449), .ZN(
        n20435) );
  OAI21_X1 U23335 ( .B1(n20431), .B2(n20548), .A(n20430), .ZN(n20432) );
  OAI221_X1 U23336 ( .B1(n20783), .B2(n20433), .C1(n20781), .C2(n20432), .A(
        n20779), .ZN(n20452) );
  AOI22_X1 U23337 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20452), .B1(
        n20451), .B2(n20731), .ZN(n20434) );
  OAI211_X1 U23338 ( .C1(n20734), .C2(n20489), .A(n20435), .B(n20434), .ZN(
        P1_U3073) );
  AOI22_X1 U23339 ( .A1(n20789), .A2(n20450), .B1(n20788), .B2(n20449), .ZN(
        n20437) );
  AOI22_X1 U23340 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20452), .B1(
        n20451), .B2(n20735), .ZN(n20436) );
  OAI211_X1 U23341 ( .C1(n20738), .C2(n20489), .A(n20437), .B(n20436), .ZN(
        P1_U3074) );
  AOI22_X1 U23342 ( .A1(n20795), .A2(n20450), .B1(n20794), .B2(n20449), .ZN(
        n20439) );
  INV_X1 U23343 ( .A(n20489), .ZN(n20468) );
  AOI22_X1 U23344 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20452), .B1(
        n20468), .B2(n20796), .ZN(n20438) );
  OAI211_X1 U23345 ( .C1(n20799), .C2(n20448), .A(n20439), .B(n20438), .ZN(
        P1_U3075) );
  AOI22_X1 U23346 ( .A1(n20801), .A2(n20450), .B1(n20800), .B2(n20449), .ZN(
        n20441) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20452), .B1(
        n20451), .B2(n20743), .ZN(n20440) );
  OAI211_X1 U23348 ( .C1(n20746), .C2(n20489), .A(n20441), .B(n20440), .ZN(
        P1_U3076) );
  AOI22_X1 U23349 ( .A1(n20807), .A2(n20450), .B1(n20806), .B2(n20449), .ZN(
        n20443) );
  AOI22_X1 U23350 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20452), .B1(
        n20468), .B2(n20808), .ZN(n20442) );
  OAI211_X1 U23351 ( .C1(n20811), .C2(n20448), .A(n20443), .B(n20442), .ZN(
        P1_U3077) );
  AOI22_X1 U23352 ( .A1(n20813), .A2(n20449), .B1(n20812), .B2(n20450), .ZN(
        n20445) );
  AOI22_X1 U23353 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20452), .B1(
        n20468), .B2(n20814), .ZN(n20444) );
  OAI211_X1 U23354 ( .C1(n20817), .C2(n20448), .A(n20445), .B(n20444), .ZN(
        P1_U3078) );
  AOI22_X1 U23355 ( .A1(n20819), .A2(n20450), .B1(n20818), .B2(n20449), .ZN(
        n20447) );
  AOI22_X1 U23356 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20452), .B1(
        n20468), .B2(n20820), .ZN(n20446) );
  OAI211_X1 U23357 ( .C1(n20823), .C2(n20448), .A(n20447), .B(n20446), .ZN(
        P1_U3079) );
  AOI22_X1 U23358 ( .A1(n20827), .A2(n20450), .B1(n20825), .B2(n20449), .ZN(
        n20454) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20452), .B1(
        n20451), .B2(n20761), .ZN(n20453) );
  OAI211_X1 U23360 ( .C1(n20766), .C2(n20489), .A(n20454), .B(n20453), .ZN(
        P1_U3080) );
  NAND2_X1 U23361 ( .A1(n20692), .A2(n10147), .ZN(n20483) );
  OAI22_X1 U23362 ( .A1(n20512), .A2(n20734), .B1(n20647), .B2(n20483), .ZN(
        n20455) );
  INV_X1 U23363 ( .A(n20455), .ZN(n20464) );
  NAND2_X1 U23364 ( .A1(n20512), .A2(n20489), .ZN(n20456) );
  AOI21_X1 U23365 ( .B1(n20456), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20781), 
        .ZN(n20459) );
  NAND2_X1 U23366 ( .A1(n20491), .A2(n9665), .ZN(n20461) );
  AOI22_X1 U23367 ( .A1(n20459), .A2(n20461), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20483), .ZN(n20458) );
  NAND3_X1 U23368 ( .A1(n20729), .A2(n20458), .A3(n20457), .ZN(n20486) );
  INV_X1 U23369 ( .A(n20459), .ZN(n20462) );
  OAI22_X1 U23370 ( .A1(n20462), .A2(n20461), .B1(n20460), .B2(n20723), .ZN(
        n20485) );
  AOI22_X1 U23371 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20486), .B1(
        n20773), .B2(n20485), .ZN(n20463) );
  OAI211_X1 U23372 ( .C1(n20787), .C2(n20489), .A(n20464), .B(n20463), .ZN(
        P1_U3081) );
  OAI22_X1 U23373 ( .A1(n20489), .A2(n20793), .B1(n20660), .B2(n20483), .ZN(
        n20465) );
  INV_X1 U23374 ( .A(n20465), .ZN(n20467) );
  AOI22_X1 U23375 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20486), .B1(
        n20788), .B2(n20485), .ZN(n20466) );
  OAI211_X1 U23376 ( .C1(n20738), .C2(n20512), .A(n20467), .B(n20466), .ZN(
        P1_U3082) );
  INV_X1 U23377 ( .A(n20483), .ZN(n20477) );
  AOI22_X1 U23378 ( .A1(n20468), .A2(n20739), .B1(n20795), .B2(n20477), .ZN(
        n20470) );
  AOI22_X1 U23379 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20486), .B1(
        n20794), .B2(n20485), .ZN(n20469) );
  OAI211_X1 U23380 ( .C1(n20742), .C2(n20512), .A(n20470), .B(n20469), .ZN(
        P1_U3083) );
  OAI22_X1 U23381 ( .A1(n20489), .A2(n20805), .B1(n20668), .B2(n20483), .ZN(
        n20471) );
  INV_X1 U23382 ( .A(n20471), .ZN(n20473) );
  AOI22_X1 U23383 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20486), .B1(
        n20800), .B2(n20485), .ZN(n20472) );
  OAI211_X1 U23384 ( .C1(n20746), .C2(n20512), .A(n20473), .B(n20472), .ZN(
        P1_U3084) );
  OAI22_X1 U23385 ( .A1(n20489), .A2(n20811), .B1(n20672), .B2(n20483), .ZN(
        n20474) );
  INV_X1 U23386 ( .A(n20474), .ZN(n20476) );
  AOI22_X1 U23387 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20486), .B1(
        n20806), .B2(n20485), .ZN(n20475) );
  OAI211_X1 U23388 ( .C1(n20750), .C2(n20512), .A(n20476), .B(n20475), .ZN(
        P1_U3085) );
  AOI22_X1 U23389 ( .A1(n20515), .A2(n20814), .B1(n20812), .B2(n20477), .ZN(
        n20479) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20486), .B1(
        n20813), .B2(n20485), .ZN(n20478) );
  OAI211_X1 U23391 ( .C1(n20817), .C2(n20489), .A(n20479), .B(n20478), .ZN(
        P1_U3086) );
  OAI22_X1 U23392 ( .A1(n20512), .A2(n20758), .B1(n20680), .B2(n20483), .ZN(
        n20480) );
  INV_X1 U23393 ( .A(n20480), .ZN(n20482) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20486), .B1(
        n20818), .B2(n20485), .ZN(n20481) );
  OAI211_X1 U23395 ( .C1(n20823), .C2(n20489), .A(n20482), .B(n20481), .ZN(
        P1_U3087) );
  OAI22_X1 U23396 ( .A1(n20512), .A2(n20766), .B1(n20685), .B2(n20483), .ZN(
        n20484) );
  INV_X1 U23397 ( .A(n20484), .ZN(n20488) );
  AOI22_X1 U23398 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20486), .B1(
        n20825), .B2(n20485), .ZN(n20487) );
  OAI211_X1 U23399 ( .C1(n20834), .C2(n20489), .A(n20488), .B(n20487), .ZN(
        P1_U3088) );
  NAND2_X1 U23400 ( .A1(n20490), .A2(n20621), .ZN(n20519) );
  INV_X1 U23401 ( .A(n20492), .ZN(n20514) );
  NAND2_X1 U23402 ( .A1(n20491), .A2(n20767), .ZN(n20493) );
  NAND2_X1 U23403 ( .A1(n20493), .A2(n20492), .ZN(n20494) );
  NAND2_X1 U23404 ( .A1(n20494), .A2(n20783), .ZN(n20496) );
  NAND2_X1 U23405 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n10147), .ZN(n20495) );
  NAND2_X1 U23406 ( .A1(n20496), .A2(n20495), .ZN(n20513) );
  AOI22_X1 U23407 ( .A1(n20774), .A2(n20514), .B1(n20773), .B2(n20513), .ZN(
        n20499) );
  OAI21_X1 U23408 ( .B1(n10147), .B2(n20497), .A(n20779), .ZN(n20516) );
  AOI22_X1 U23409 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20731), .ZN(n20498) );
  OAI211_X1 U23410 ( .C1(n20734), .C2(n20519), .A(n20499), .B(n20498), .ZN(
        P1_U3089) );
  AOI22_X1 U23411 ( .A1(n20789), .A2(n20514), .B1(n20788), .B2(n20513), .ZN(
        n20501) );
  AOI22_X1 U23412 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20516), .B1(
        n20542), .B2(n20790), .ZN(n20500) );
  OAI211_X1 U23413 ( .C1(n20793), .C2(n20512), .A(n20501), .B(n20500), .ZN(
        P1_U3090) );
  AOI22_X1 U23414 ( .A1(n20795), .A2(n20514), .B1(n20794), .B2(n20513), .ZN(
        n20503) );
  AOI22_X1 U23415 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20739), .ZN(n20502) );
  OAI211_X1 U23416 ( .C1(n20742), .C2(n20519), .A(n20503), .B(n20502), .ZN(
        P1_U3091) );
  AOI22_X1 U23417 ( .A1(n20801), .A2(n20514), .B1(n20800), .B2(n20513), .ZN(
        n20505) );
  AOI22_X1 U23418 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20743), .ZN(n20504) );
  OAI211_X1 U23419 ( .C1(n20746), .C2(n20519), .A(n20505), .B(n20504), .ZN(
        P1_U3092) );
  AOI22_X1 U23420 ( .A1(n20807), .A2(n20514), .B1(n20806), .B2(n20513), .ZN(
        n20507) );
  AOI22_X1 U23421 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20747), .ZN(n20506) );
  OAI211_X1 U23422 ( .C1(n20750), .C2(n20519), .A(n20507), .B(n20506), .ZN(
        P1_U3093) );
  AOI22_X1 U23423 ( .A1(n20813), .A2(n20513), .B1(n20812), .B2(n20514), .ZN(
        n20509) );
  AOI22_X1 U23424 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20751), .ZN(n20508) );
  OAI211_X1 U23425 ( .C1(n20754), .C2(n20519), .A(n20509), .B(n20508), .ZN(
        P1_U3094) );
  AOI22_X1 U23426 ( .A1(n20819), .A2(n20514), .B1(n20818), .B2(n20513), .ZN(
        n20511) );
  AOI22_X1 U23427 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20516), .B1(
        n20542), .B2(n20820), .ZN(n20510) );
  OAI211_X1 U23428 ( .C1(n20823), .C2(n20512), .A(n20511), .B(n20510), .ZN(
        P1_U3095) );
  AOI22_X1 U23429 ( .A1(n20827), .A2(n20514), .B1(n20825), .B2(n20513), .ZN(
        n20518) );
  AOI22_X1 U23430 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20761), .ZN(n20517) );
  OAI211_X1 U23431 ( .C1(n20766), .C2(n20519), .A(n20518), .B(n20517), .ZN(
        P1_U3096) );
  NOR3_X1 U23432 ( .A1(n20645), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20550) );
  INV_X1 U23433 ( .A(n20550), .ZN(n20546) );
  NOR2_X1 U23434 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20546), .ZN(
        n20541) );
  AND2_X1 U23435 ( .A1(n13423), .A2(n13416), .ZN(n20611) );
  AOI21_X1 U23436 ( .B1(n20611), .B2(n20651), .A(n20541), .ZN(n20522) );
  AND2_X1 U23437 ( .A1(n20520), .A2(n20575), .ZN(n20653) );
  INV_X1 U23438 ( .A(n20653), .ZN(n20655) );
  OAI22_X1 U23439 ( .A1(n20522), .A2(n20781), .B1(n20579), .B2(n20655), .ZN(
        n20540) );
  AOI22_X1 U23440 ( .A1(n20774), .A2(n20541), .B1(n20773), .B2(n20540), .ZN(
        n20527) );
  INV_X1 U23441 ( .A(n20571), .ZN(n20521) );
  OAI21_X1 U23442 ( .B1(n20521), .B2(n20542), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20523) );
  NAND2_X1 U23443 ( .A1(n20523), .A2(n20522), .ZN(n20524) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20543), .B1(
        n20542), .B2(n20731), .ZN(n20526) );
  OAI211_X1 U23445 ( .C1(n20734), .C2(n20571), .A(n20527), .B(n20526), .ZN(
        P1_U3097) );
  AOI22_X1 U23446 ( .A1(n20789), .A2(n20541), .B1(n20788), .B2(n20540), .ZN(
        n20529) );
  AOI22_X1 U23447 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20543), .B1(
        n20542), .B2(n20735), .ZN(n20528) );
  OAI211_X1 U23448 ( .C1(n20738), .C2(n20571), .A(n20529), .B(n20528), .ZN(
        P1_U3098) );
  AOI22_X1 U23449 ( .A1(n20795), .A2(n20541), .B1(n20794), .B2(n20540), .ZN(
        n20531) );
  AOI22_X1 U23450 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20543), .B1(
        n20542), .B2(n20739), .ZN(n20530) );
  OAI211_X1 U23451 ( .C1(n20742), .C2(n20571), .A(n20531), .B(n20530), .ZN(
        P1_U3099) );
  AOI22_X1 U23452 ( .A1(n20801), .A2(n20541), .B1(n20800), .B2(n20540), .ZN(
        n20533) );
  AOI22_X1 U23453 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20543), .B1(
        n20542), .B2(n20743), .ZN(n20532) );
  OAI211_X1 U23454 ( .C1(n20746), .C2(n20571), .A(n20533), .B(n20532), .ZN(
        P1_U3100) );
  AOI22_X1 U23455 ( .A1(n20807), .A2(n20541), .B1(n20806), .B2(n20540), .ZN(
        n20535) );
  AOI22_X1 U23456 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20543), .B1(
        n20542), .B2(n20747), .ZN(n20534) );
  OAI211_X1 U23457 ( .C1(n20750), .C2(n20571), .A(n20535), .B(n20534), .ZN(
        P1_U3101) );
  AOI22_X1 U23458 ( .A1(n20813), .A2(n20540), .B1(n20812), .B2(n20541), .ZN(
        n20537) );
  AOI22_X1 U23459 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20543), .B1(
        n20542), .B2(n20751), .ZN(n20536) );
  OAI211_X1 U23460 ( .C1(n20754), .C2(n20571), .A(n20537), .B(n20536), .ZN(
        P1_U3102) );
  AOI22_X1 U23461 ( .A1(n20819), .A2(n20541), .B1(n20818), .B2(n20540), .ZN(
        n20539) );
  AOI22_X1 U23462 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20543), .B1(
        n20542), .B2(n20755), .ZN(n20538) );
  OAI211_X1 U23463 ( .C1(n20758), .C2(n20571), .A(n20539), .B(n20538), .ZN(
        P1_U3103) );
  AOI22_X1 U23464 ( .A1(n20827), .A2(n20541), .B1(n20825), .B2(n20540), .ZN(
        n20545) );
  AOI22_X1 U23465 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20543), .B1(
        n20542), .B2(n20761), .ZN(n20544) );
  OAI211_X1 U23466 ( .C1(n20766), .C2(n20571), .A(n20545), .B(n20544), .ZN(
        P1_U3104) );
  NOR2_X1 U23467 ( .A1(n20692), .A2(n20546), .ZN(n20567) );
  AOI21_X1 U23468 ( .B1(n20611), .B2(n20693), .A(n20567), .ZN(n20547) );
  OAI22_X1 U23469 ( .A1(n20547), .A2(n20781), .B1(n20546), .B2(n20837), .ZN(
        n20566) );
  AOI22_X1 U23470 ( .A1(n20774), .A2(n20567), .B1(n20773), .B2(n20566), .ZN(
        n20553) );
  OAI211_X1 U23471 ( .C1(n20618), .C2(n20548), .A(n20783), .B(n20547), .ZN(
        n20549) );
  OAI211_X1 U23472 ( .C1(n20783), .C2(n20550), .A(n20779), .B(n20549), .ZN(
        n20568) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20568), .B1(
        n20597), .B2(n20784), .ZN(n20552) );
  OAI211_X1 U23474 ( .C1(n20787), .C2(n20571), .A(n20553), .B(n20552), .ZN(
        P1_U3105) );
  AOI22_X1 U23475 ( .A1(n20789), .A2(n20567), .B1(n20788), .B2(n20566), .ZN(
        n20555) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20568), .B1(
        n20597), .B2(n20790), .ZN(n20554) );
  OAI211_X1 U23477 ( .C1(n20793), .C2(n20571), .A(n20555), .B(n20554), .ZN(
        P1_U3106) );
  AOI22_X1 U23478 ( .A1(n20795), .A2(n20567), .B1(n20794), .B2(n20566), .ZN(
        n20557) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20568), .B1(
        n20597), .B2(n20796), .ZN(n20556) );
  OAI211_X1 U23480 ( .C1(n20799), .C2(n20571), .A(n20557), .B(n20556), .ZN(
        P1_U3107) );
  AOI22_X1 U23481 ( .A1(n20801), .A2(n20567), .B1(n20800), .B2(n20566), .ZN(
        n20559) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20568), .B1(
        n20597), .B2(n20802), .ZN(n20558) );
  OAI211_X1 U23483 ( .C1(n20805), .C2(n20571), .A(n20559), .B(n20558), .ZN(
        P1_U3108) );
  AOI22_X1 U23484 ( .A1(n20807), .A2(n20567), .B1(n20806), .B2(n20566), .ZN(
        n20561) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20568), .B1(
        n20597), .B2(n20808), .ZN(n20560) );
  OAI211_X1 U23486 ( .C1(n20811), .C2(n20571), .A(n20561), .B(n20560), .ZN(
        P1_U3109) );
  AOI22_X1 U23487 ( .A1(n20813), .A2(n20566), .B1(n20812), .B2(n20567), .ZN(
        n20563) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20568), .B1(
        n20597), .B2(n20814), .ZN(n20562) );
  OAI211_X1 U23489 ( .C1(n20817), .C2(n20571), .A(n20563), .B(n20562), .ZN(
        P1_U3110) );
  AOI22_X1 U23490 ( .A1(n20819), .A2(n20567), .B1(n20818), .B2(n20566), .ZN(
        n20565) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20568), .B1(
        n20597), .B2(n20820), .ZN(n20564) );
  OAI211_X1 U23492 ( .C1(n20823), .C2(n20571), .A(n20565), .B(n20564), .ZN(
        P1_U3111) );
  AOI22_X1 U23493 ( .A1(n20827), .A2(n20567), .B1(n20825), .B2(n20566), .ZN(
        n20570) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20568), .B1(
        n20597), .B2(n20828), .ZN(n20569) );
  OAI211_X1 U23495 ( .C1(n20834), .C2(n20571), .A(n20570), .B(n20569), .ZN(
        P1_U3112) );
  NOR3_X1 U23496 ( .A1(n20645), .A2(n20572), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20620) );
  NAND2_X1 U23497 ( .A1(n20692), .A2(n20620), .ZN(n20603) );
  OAI22_X1 U23498 ( .A1(n20609), .A2(n20787), .B1(n20647), .B2(n20603), .ZN(
        n20573) );
  INV_X1 U23499 ( .A(n20573), .ZN(n20583) );
  NAND2_X1 U23500 ( .A1(n20644), .A2(n20609), .ZN(n20574) );
  AOI21_X1 U23501 ( .B1(n20574), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20781), 
        .ZN(n20578) );
  NAND2_X1 U23502 ( .A1(n20611), .A2(n9665), .ZN(n20580) );
  AOI22_X1 U23503 ( .A1(n20578), .A2(n20580), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20603), .ZN(n20576) );
  OR2_X1 U23504 ( .A1(n20575), .A2(n20645), .ZN(n20724) );
  NAND2_X1 U23505 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20724), .ZN(n20728) );
  NAND3_X1 U23506 ( .A1(n20577), .A2(n20576), .A3(n20728), .ZN(n20606) );
  INV_X1 U23507 ( .A(n20578), .ZN(n20581) );
  AOI22_X1 U23508 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20606), .B1(
        n20773), .B2(n20605), .ZN(n20582) );
  OAI211_X1 U23509 ( .C1(n20734), .C2(n20644), .A(n20583), .B(n20582), .ZN(
        P1_U3113) );
  OAI22_X1 U23510 ( .A1(n20609), .A2(n20793), .B1(n20660), .B2(n20603), .ZN(
        n20584) );
  INV_X1 U23511 ( .A(n20584), .ZN(n20586) );
  AOI22_X1 U23512 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20606), .B1(
        n20788), .B2(n20605), .ZN(n20585) );
  OAI211_X1 U23513 ( .C1(n20738), .C2(n20644), .A(n20586), .B(n20585), .ZN(
        P1_U3114) );
  OAI22_X1 U23514 ( .A1(n20644), .A2(n20742), .B1(n20664), .B2(n20603), .ZN(
        n20587) );
  INV_X1 U23515 ( .A(n20587), .ZN(n20589) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20606), .B1(
        n20794), .B2(n20605), .ZN(n20588) );
  OAI211_X1 U23517 ( .C1(n20799), .C2(n20609), .A(n20589), .B(n20588), .ZN(
        P1_U3115) );
  OAI22_X1 U23518 ( .A1(n20644), .A2(n20746), .B1(n20668), .B2(n20603), .ZN(
        n20590) );
  INV_X1 U23519 ( .A(n20590), .ZN(n20592) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20606), .B1(
        n20800), .B2(n20605), .ZN(n20591) );
  OAI211_X1 U23521 ( .C1(n20805), .C2(n20609), .A(n20592), .B(n20591), .ZN(
        P1_U3116) );
  OAI22_X1 U23522 ( .A1(n20609), .A2(n20811), .B1(n20672), .B2(n20603), .ZN(
        n20593) );
  INV_X1 U23523 ( .A(n20593), .ZN(n20595) );
  AOI22_X1 U23524 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20606), .B1(
        n20806), .B2(n20605), .ZN(n20594) );
  OAI211_X1 U23525 ( .C1(n20750), .C2(n20644), .A(n20595), .B(n20594), .ZN(
        P1_U3117) );
  INV_X1 U23526 ( .A(n20603), .ZN(n20596) );
  AOI22_X1 U23527 ( .A1(n20597), .A2(n20751), .B1(n20812), .B2(n20596), .ZN(
        n20599) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20606), .B1(
        n20813), .B2(n20605), .ZN(n20598) );
  OAI211_X1 U23529 ( .C1(n20754), .C2(n20644), .A(n20599), .B(n20598), .ZN(
        P1_U3118) );
  OAI22_X1 U23530 ( .A1(n20644), .A2(n20758), .B1(n20680), .B2(n20603), .ZN(
        n20600) );
  INV_X1 U23531 ( .A(n20600), .ZN(n20602) );
  AOI22_X1 U23532 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20606), .B1(
        n20818), .B2(n20605), .ZN(n20601) );
  OAI211_X1 U23533 ( .C1(n20823), .C2(n20609), .A(n20602), .B(n20601), .ZN(
        P1_U3119) );
  OAI22_X1 U23534 ( .A1(n20644), .A2(n20766), .B1(n20685), .B2(n20603), .ZN(
        n20604) );
  INV_X1 U23535 ( .A(n20604), .ZN(n20608) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20606), .B1(
        n20825), .B2(n20605), .ZN(n20607) );
  OAI211_X1 U23537 ( .C1(n20834), .C2(n20609), .A(n20608), .B(n20607), .ZN(
        P1_U3120) );
  OR2_X1 U23538 ( .A1(n20610), .A2(n20645), .ZN(n20612) );
  INV_X1 U23539 ( .A(n20612), .ZN(n20639) );
  NAND2_X1 U23540 ( .A1(n20611), .A2(n20767), .ZN(n20613) );
  NAND2_X1 U23541 ( .A1(n20613), .A2(n20612), .ZN(n20616) );
  NAND2_X1 U23542 ( .A1(n20616), .A2(n20783), .ZN(n20615) );
  NAND2_X1 U23543 ( .A1(n20620), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20614) );
  NAND2_X1 U23544 ( .A1(n20615), .A2(n20614), .ZN(n20638) );
  AOI22_X1 U23545 ( .A1(n20774), .A2(n20639), .B1(n20773), .B2(n20638), .ZN(
        n20624) );
  INV_X1 U23546 ( .A(n20616), .ZN(n20617) );
  OAI211_X1 U23547 ( .C1(n20618), .C2(n20777), .A(n20783), .B(n20617), .ZN(
        n20619) );
  OAI211_X1 U23548 ( .C1(n20783), .C2(n20620), .A(n20779), .B(n20619), .ZN(
        n20641) );
  AOI22_X1 U23549 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20784), .ZN(n20623) );
  OAI211_X1 U23550 ( .C1(n20787), .C2(n20644), .A(n20624), .B(n20623), .ZN(
        P1_U3121) );
  AOI22_X1 U23551 ( .A1(n20789), .A2(n20639), .B1(n20788), .B2(n20638), .ZN(
        n20626) );
  INV_X1 U23552 ( .A(n20644), .ZN(n20633) );
  AOI22_X1 U23553 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20641), .B1(
        n20633), .B2(n20735), .ZN(n20625) );
  OAI211_X1 U23554 ( .C1(n20738), .C2(n20691), .A(n20626), .B(n20625), .ZN(
        P1_U3122) );
  AOI22_X1 U23555 ( .A1(n20795), .A2(n20639), .B1(n20794), .B2(n20638), .ZN(
        n20628) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20796), .ZN(n20627) );
  OAI211_X1 U23557 ( .C1(n20799), .C2(n20644), .A(n20628), .B(n20627), .ZN(
        P1_U3123) );
  AOI22_X1 U23558 ( .A1(n20801), .A2(n20639), .B1(n20800), .B2(n20638), .ZN(
        n20630) );
  AOI22_X1 U23559 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20802), .ZN(n20629) );
  OAI211_X1 U23560 ( .C1(n20805), .C2(n20644), .A(n20630), .B(n20629), .ZN(
        P1_U3124) );
  AOI22_X1 U23561 ( .A1(n20807), .A2(n20639), .B1(n20806), .B2(n20638), .ZN(
        n20632) );
  AOI22_X1 U23562 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20808), .ZN(n20631) );
  OAI211_X1 U23563 ( .C1(n20811), .C2(n20644), .A(n20632), .B(n20631), .ZN(
        P1_U3125) );
  AOI22_X1 U23564 ( .A1(n20813), .A2(n20638), .B1(n20812), .B2(n20639), .ZN(
        n20635) );
  AOI22_X1 U23565 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20641), .B1(
        n20633), .B2(n20751), .ZN(n20634) );
  OAI211_X1 U23566 ( .C1(n20754), .C2(n20691), .A(n20635), .B(n20634), .ZN(
        P1_U3126) );
  AOI22_X1 U23567 ( .A1(n20819), .A2(n20639), .B1(n20818), .B2(n20638), .ZN(
        n20637) );
  AOI22_X1 U23568 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20820), .ZN(n20636) );
  OAI211_X1 U23569 ( .C1(n20823), .C2(n20644), .A(n20637), .B(n20636), .ZN(
        P1_U3127) );
  AOI22_X1 U23570 ( .A1(n20827), .A2(n20639), .B1(n20825), .B2(n20638), .ZN(
        n20643) );
  AOI22_X1 U23571 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20828), .ZN(n20642) );
  OAI211_X1 U23572 ( .C1(n20834), .C2(n20644), .A(n20643), .B(n20642), .ZN(
        P1_U3128) );
  NOR3_X1 U23573 ( .A1(n20646), .A2(n20645), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20697) );
  NAND2_X1 U23574 ( .A1(n20692), .A2(n20697), .ZN(n20684) );
  OAI22_X1 U23575 ( .A1(n20718), .A2(n20734), .B1(n20647), .B2(n20684), .ZN(
        n20648) );
  INV_X1 U23576 ( .A(n20648), .ZN(n20659) );
  NAND2_X1 U23577 ( .A1(n20691), .A2(n20718), .ZN(n20649) );
  AOI21_X1 U23578 ( .B1(n20649), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20781), 
        .ZN(n20654) );
  NOR2_X1 U23579 ( .A1(n13416), .A2(n20650), .ZN(n20768) );
  NAND2_X1 U23580 ( .A1(n20768), .A2(n20651), .ZN(n20656) );
  AOI22_X1 U23581 ( .A1(n20654), .A2(n20656), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20684), .ZN(n20652) );
  OAI211_X1 U23582 ( .C1(n20653), .C2(n20837), .A(n20729), .B(n20652), .ZN(
        n20688) );
  INV_X1 U23583 ( .A(n20654), .ZN(n20657) );
  OAI22_X1 U23584 ( .A1(n20657), .A2(n20656), .B1(n20723), .B2(n20655), .ZN(
        n20687) );
  AOI22_X1 U23585 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20688), .B1(
        n20773), .B2(n20687), .ZN(n20658) );
  OAI211_X1 U23586 ( .C1(n20787), .C2(n20691), .A(n20659), .B(n20658), .ZN(
        P1_U3129) );
  OAI22_X1 U23587 ( .A1(n20718), .A2(n20738), .B1(n20660), .B2(n20684), .ZN(
        n20661) );
  INV_X1 U23588 ( .A(n20661), .ZN(n20663) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20688), .B1(
        n20788), .B2(n20687), .ZN(n20662) );
  OAI211_X1 U23590 ( .C1(n20793), .C2(n20691), .A(n20663), .B(n20662), .ZN(
        P1_U3130) );
  OAI22_X1 U23591 ( .A1(n20718), .A2(n20742), .B1(n20664), .B2(n20684), .ZN(
        n20665) );
  INV_X1 U23592 ( .A(n20665), .ZN(n20667) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20688), .B1(
        n20794), .B2(n20687), .ZN(n20666) );
  OAI211_X1 U23594 ( .C1(n20799), .C2(n20691), .A(n20667), .B(n20666), .ZN(
        P1_U3131) );
  OAI22_X1 U23595 ( .A1(n20718), .A2(n20746), .B1(n20668), .B2(n20684), .ZN(
        n20669) );
  INV_X1 U23596 ( .A(n20669), .ZN(n20671) );
  AOI22_X1 U23597 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20688), .B1(
        n20800), .B2(n20687), .ZN(n20670) );
  OAI211_X1 U23598 ( .C1(n20805), .C2(n20691), .A(n20671), .B(n20670), .ZN(
        P1_U3132) );
  OAI22_X1 U23599 ( .A1(n20718), .A2(n20750), .B1(n20672), .B2(n20684), .ZN(
        n20673) );
  INV_X1 U23600 ( .A(n20673), .ZN(n20675) );
  AOI22_X1 U23601 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20688), .B1(
        n20806), .B2(n20687), .ZN(n20674) );
  OAI211_X1 U23602 ( .C1(n20811), .C2(n20691), .A(n20675), .B(n20674), .ZN(
        P1_U3133) );
  INV_X1 U23603 ( .A(n20718), .ZN(n20677) );
  INV_X1 U23604 ( .A(n20684), .ZN(n20676) );
  AOI22_X1 U23605 ( .A1(n20677), .A2(n20814), .B1(n20812), .B2(n20676), .ZN(
        n20679) );
  AOI22_X1 U23606 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20688), .B1(
        n20813), .B2(n20687), .ZN(n20678) );
  OAI211_X1 U23607 ( .C1(n20817), .C2(n20691), .A(n20679), .B(n20678), .ZN(
        P1_U3134) );
  OAI22_X1 U23608 ( .A1(n20718), .A2(n20758), .B1(n20680), .B2(n20684), .ZN(
        n20681) );
  INV_X1 U23609 ( .A(n20681), .ZN(n20683) );
  AOI22_X1 U23610 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20688), .B1(
        n20818), .B2(n20687), .ZN(n20682) );
  OAI211_X1 U23611 ( .C1(n20823), .C2(n20691), .A(n20683), .B(n20682), .ZN(
        P1_U3135) );
  OAI22_X1 U23612 ( .A1(n20718), .A2(n20766), .B1(n20685), .B2(n20684), .ZN(
        n20686) );
  INV_X1 U23613 ( .A(n20686), .ZN(n20690) );
  AOI22_X1 U23614 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20688), .B1(
        n20825), .B2(n20687), .ZN(n20689) );
  OAI211_X1 U23615 ( .C1(n20834), .C2(n20691), .A(n20690), .B(n20689), .ZN(
        P1_U3136) );
  INV_X1 U23616 ( .A(n20697), .ZN(n20694) );
  NOR2_X1 U23617 ( .A1(n20692), .A2(n20694), .ZN(n20714) );
  AOI21_X1 U23618 ( .B1(n20768), .B2(n20693), .A(n20714), .ZN(n20695) );
  OAI22_X1 U23619 ( .A1(n20695), .A2(n20781), .B1(n20694), .B2(n20837), .ZN(
        n20713) );
  AOI22_X1 U23620 ( .A1(n20774), .A2(n20714), .B1(n20773), .B2(n20713), .ZN(
        n20700) );
  OAI21_X1 U23621 ( .B1(n20697), .B2(n20696), .A(n20779), .ZN(n20715) );
  NOR2_X2 U23622 ( .A1(n20778), .A2(n20698), .ZN(n20762) );
  AOI22_X1 U23623 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20715), .B1(
        n20762), .B2(n20784), .ZN(n20699) );
  OAI211_X1 U23624 ( .C1(n20787), .C2(n20718), .A(n20700), .B(n20699), .ZN(
        P1_U3137) );
  AOI22_X1 U23625 ( .A1(n20789), .A2(n20714), .B1(n20788), .B2(n20713), .ZN(
        n20702) );
  AOI22_X1 U23626 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20715), .B1(
        n20762), .B2(n20790), .ZN(n20701) );
  OAI211_X1 U23627 ( .C1(n20793), .C2(n20718), .A(n20702), .B(n20701), .ZN(
        P1_U3138) );
  AOI22_X1 U23628 ( .A1(n20795), .A2(n20714), .B1(n20794), .B2(n20713), .ZN(
        n20704) );
  AOI22_X1 U23629 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20715), .B1(
        n20762), .B2(n20796), .ZN(n20703) );
  OAI211_X1 U23630 ( .C1(n20799), .C2(n20718), .A(n20704), .B(n20703), .ZN(
        P1_U3139) );
  AOI22_X1 U23631 ( .A1(n20801), .A2(n20714), .B1(n20800), .B2(n20713), .ZN(
        n20706) );
  AOI22_X1 U23632 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20715), .B1(
        n20762), .B2(n20802), .ZN(n20705) );
  OAI211_X1 U23633 ( .C1(n20805), .C2(n20718), .A(n20706), .B(n20705), .ZN(
        P1_U3140) );
  AOI22_X1 U23634 ( .A1(n20807), .A2(n20714), .B1(n20806), .B2(n20713), .ZN(
        n20708) );
  AOI22_X1 U23635 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20715), .B1(
        n20762), .B2(n20808), .ZN(n20707) );
  OAI211_X1 U23636 ( .C1(n20811), .C2(n20718), .A(n20708), .B(n20707), .ZN(
        P1_U3141) );
  AOI22_X1 U23637 ( .A1(n20813), .A2(n20713), .B1(n20812), .B2(n20714), .ZN(
        n20710) );
  AOI22_X1 U23638 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20715), .B1(
        n20762), .B2(n20814), .ZN(n20709) );
  OAI211_X1 U23639 ( .C1(n20817), .C2(n20718), .A(n20710), .B(n20709), .ZN(
        P1_U3142) );
  AOI22_X1 U23640 ( .A1(n20819), .A2(n20714), .B1(n20818), .B2(n20713), .ZN(
        n20712) );
  AOI22_X1 U23641 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20715), .B1(
        n20762), .B2(n20820), .ZN(n20711) );
  OAI211_X1 U23642 ( .C1(n20823), .C2(n20718), .A(n20712), .B(n20711), .ZN(
        P1_U3143) );
  AOI22_X1 U23643 ( .A1(n20827), .A2(n20714), .B1(n20825), .B2(n20713), .ZN(
        n20717) );
  AOI22_X1 U23644 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20715), .B1(
        n20762), .B2(n20828), .ZN(n20716) );
  OAI211_X1 U23645 ( .C1(n20834), .C2(n20718), .A(n20717), .B(n20716), .ZN(
        P1_U3144) );
  INV_X1 U23646 ( .A(n20782), .ZN(n20721) );
  NOR2_X1 U23647 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20721), .ZN(
        n20760) );
  NAND3_X1 U23648 ( .A1(n20768), .A2(n9665), .A3(n20783), .ZN(n20722) );
  OAI21_X1 U23649 ( .B1(n20724), .B2(n20723), .A(n20722), .ZN(n20759) );
  AOI22_X1 U23650 ( .A1(n20774), .A2(n20760), .B1(n20773), .B2(n20759), .ZN(
        n20733) );
  INV_X1 U23651 ( .A(n20762), .ZN(n20725) );
  AOI21_X1 U23652 ( .B1(n20725), .B2(n20833), .A(n21034), .ZN(n20726) );
  AOI21_X1 U23653 ( .B1(n20768), .B2(n9665), .A(n20726), .ZN(n20727) );
  NOR2_X1 U23654 ( .A1(n20727), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20730) );
  AOI22_X1 U23655 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20763), .B1(
        n20762), .B2(n20731), .ZN(n20732) );
  OAI211_X1 U23656 ( .C1(n20734), .C2(n20833), .A(n20733), .B(n20732), .ZN(
        P1_U3145) );
  AOI22_X1 U23657 ( .A1(n20789), .A2(n20760), .B1(n20788), .B2(n20759), .ZN(
        n20737) );
  AOI22_X1 U23658 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20763), .B1(
        n20762), .B2(n20735), .ZN(n20736) );
  OAI211_X1 U23659 ( .C1(n20738), .C2(n20833), .A(n20737), .B(n20736), .ZN(
        P1_U3146) );
  AOI22_X1 U23660 ( .A1(n20795), .A2(n20760), .B1(n20794), .B2(n20759), .ZN(
        n20741) );
  AOI22_X1 U23661 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20763), .B1(
        n20762), .B2(n20739), .ZN(n20740) );
  OAI211_X1 U23662 ( .C1(n20742), .C2(n20833), .A(n20741), .B(n20740), .ZN(
        P1_U3147) );
  AOI22_X1 U23663 ( .A1(n20801), .A2(n20760), .B1(n20800), .B2(n20759), .ZN(
        n20745) );
  AOI22_X1 U23664 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20763), .B1(
        n20762), .B2(n20743), .ZN(n20744) );
  OAI211_X1 U23665 ( .C1(n20746), .C2(n20833), .A(n20745), .B(n20744), .ZN(
        P1_U3148) );
  AOI22_X1 U23666 ( .A1(n20807), .A2(n20760), .B1(n20806), .B2(n20759), .ZN(
        n20749) );
  AOI22_X1 U23667 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20763), .B1(
        n20762), .B2(n20747), .ZN(n20748) );
  OAI211_X1 U23668 ( .C1(n20750), .C2(n20833), .A(n20749), .B(n20748), .ZN(
        P1_U3149) );
  AOI22_X1 U23669 ( .A1(n20813), .A2(n20759), .B1(n20812), .B2(n20760), .ZN(
        n20753) );
  AOI22_X1 U23670 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20763), .B1(
        n20762), .B2(n20751), .ZN(n20752) );
  OAI211_X1 U23671 ( .C1(n20754), .C2(n20833), .A(n20753), .B(n20752), .ZN(
        P1_U3150) );
  AOI22_X1 U23672 ( .A1(n20819), .A2(n20760), .B1(n20818), .B2(n20759), .ZN(
        n20757) );
  AOI22_X1 U23673 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20763), .B1(
        n20762), .B2(n20755), .ZN(n20756) );
  OAI211_X1 U23674 ( .C1(n20758), .C2(n20833), .A(n20757), .B(n20756), .ZN(
        P1_U3151) );
  AOI22_X1 U23675 ( .A1(n20827), .A2(n20760), .B1(n20825), .B2(n20759), .ZN(
        n20765) );
  AOI22_X1 U23676 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20763), .B1(
        n20762), .B2(n20761), .ZN(n20764) );
  OAI211_X1 U23677 ( .C1(n20766), .C2(n20833), .A(n20765), .B(n20764), .ZN(
        P1_U3152) );
  INV_X1 U23678 ( .A(n20769), .ZN(n20826) );
  NAND2_X1 U23679 ( .A1(n20768), .A2(n20767), .ZN(n20770) );
  NAND2_X1 U23680 ( .A1(n20770), .A2(n20769), .ZN(n20775) );
  NAND2_X1 U23681 ( .A1(n20775), .A2(n20783), .ZN(n20772) );
  NAND2_X1 U23682 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20782), .ZN(n20771) );
  NAND2_X1 U23683 ( .A1(n20772), .A2(n20771), .ZN(n20824) );
  AOI22_X1 U23684 ( .A1(n20774), .A2(n20826), .B1(n20773), .B2(n20824), .ZN(
        n20786) );
  INV_X1 U23685 ( .A(n20775), .ZN(n20776) );
  OAI21_X1 U23686 ( .B1(n20778), .B2(n20777), .A(n20776), .ZN(n20780) );
  OAI221_X1 U23687 ( .B1(n20783), .B2(n20782), .C1(n20781), .C2(n20780), .A(
        n20779), .ZN(n20830) );
  AOI22_X1 U23688 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20830), .B1(
        n20829), .B2(n20784), .ZN(n20785) );
  OAI211_X1 U23689 ( .C1(n20787), .C2(n20833), .A(n20786), .B(n20785), .ZN(
        P1_U3153) );
  AOI22_X1 U23690 ( .A1(n20789), .A2(n20826), .B1(n20788), .B2(n20824), .ZN(
        n20792) );
  AOI22_X1 U23691 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20830), .B1(
        n20829), .B2(n20790), .ZN(n20791) );
  OAI211_X1 U23692 ( .C1(n20793), .C2(n20833), .A(n20792), .B(n20791), .ZN(
        P1_U3154) );
  AOI22_X1 U23693 ( .A1(n20795), .A2(n20826), .B1(n20794), .B2(n20824), .ZN(
        n20798) );
  AOI22_X1 U23694 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20830), .B1(
        n20829), .B2(n20796), .ZN(n20797) );
  OAI211_X1 U23695 ( .C1(n20799), .C2(n20833), .A(n20798), .B(n20797), .ZN(
        P1_U3155) );
  AOI22_X1 U23696 ( .A1(n20801), .A2(n20826), .B1(n20800), .B2(n20824), .ZN(
        n20804) );
  AOI22_X1 U23697 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20830), .B1(
        n20829), .B2(n20802), .ZN(n20803) );
  OAI211_X1 U23698 ( .C1(n20805), .C2(n20833), .A(n20804), .B(n20803), .ZN(
        P1_U3156) );
  AOI22_X1 U23699 ( .A1(n20807), .A2(n20826), .B1(n20806), .B2(n20824), .ZN(
        n20810) );
  AOI22_X1 U23700 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20830), .B1(
        n20829), .B2(n20808), .ZN(n20809) );
  OAI211_X1 U23701 ( .C1(n20811), .C2(n20833), .A(n20810), .B(n20809), .ZN(
        P1_U3157) );
  AOI22_X1 U23702 ( .A1(n20813), .A2(n20824), .B1(n20812), .B2(n20826), .ZN(
        n20816) );
  AOI22_X1 U23703 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20830), .B1(
        n20829), .B2(n20814), .ZN(n20815) );
  OAI211_X1 U23704 ( .C1(n20817), .C2(n20833), .A(n20816), .B(n20815), .ZN(
        P1_U3158) );
  AOI22_X1 U23705 ( .A1(n20819), .A2(n20826), .B1(n20818), .B2(n20824), .ZN(
        n20822) );
  AOI22_X1 U23706 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20830), .B1(
        n20829), .B2(n20820), .ZN(n20821) );
  OAI211_X1 U23707 ( .C1(n20823), .C2(n20833), .A(n20822), .B(n20821), .ZN(
        P1_U3159) );
  AOI22_X1 U23708 ( .A1(n20827), .A2(n20826), .B1(n20825), .B2(n20824), .ZN(
        n20832) );
  AOI22_X1 U23709 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20830), .B1(
        n20829), .B2(n20828), .ZN(n20831) );
  OAI211_X1 U23710 ( .C1(n20834), .C2(n20833), .A(n20832), .B(n20831), .ZN(
        P1_U3160) );
  OAI221_X1 U23711 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20838), .C1(n20837), 
        .C2(n20836), .A(n20835), .ZN(P1_U3163) );
  AND2_X1 U23712 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20839), .ZN(
        P1_U3164) );
  AND2_X1 U23713 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20839), .ZN(
        P1_U3165) );
  AND2_X1 U23714 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20839), .ZN(
        P1_U3166) );
  AND2_X1 U23715 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20839), .ZN(
        P1_U3167) );
  AND2_X1 U23716 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20839), .ZN(
        P1_U3168) );
  AND2_X1 U23717 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20839), .ZN(
        P1_U3169) );
  AND2_X1 U23718 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20839), .ZN(
        P1_U3170) );
  AND2_X1 U23719 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20839), .ZN(
        P1_U3171) );
  AND2_X1 U23720 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20839), .ZN(
        P1_U3172) );
  AND2_X1 U23721 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20839), .ZN(
        P1_U3173) );
  AND2_X1 U23722 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20839), .ZN(
        P1_U3174) );
  AND2_X1 U23723 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20839), .ZN(
        P1_U3175) );
  AND2_X1 U23724 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20839), .ZN(
        P1_U3176) );
  AND2_X1 U23725 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20839), .ZN(
        P1_U3177) );
  AND2_X1 U23726 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20839), .ZN(
        P1_U3178) );
  AND2_X1 U23727 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20839), .ZN(
        P1_U3179) );
  AND2_X1 U23728 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20839), .ZN(
        P1_U3180) );
  AND2_X1 U23729 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20839), .ZN(
        P1_U3181) );
  AND2_X1 U23730 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20839), .ZN(
        P1_U3182) );
  AND2_X1 U23731 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20839), .ZN(
        P1_U3183) );
  AND2_X1 U23732 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20839), .ZN(
        P1_U3184) );
  AND2_X1 U23733 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20839), .ZN(
        P1_U3185) );
  AND2_X1 U23734 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20839), .ZN(P1_U3186) );
  AND2_X1 U23735 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20839), .ZN(P1_U3187) );
  AND2_X1 U23736 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20839), .ZN(P1_U3188) );
  AND2_X1 U23737 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20839), .ZN(P1_U3189) );
  AND2_X1 U23738 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20839), .ZN(P1_U3190) );
  AND2_X1 U23739 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20839), .ZN(P1_U3191) );
  AND2_X1 U23740 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20839), .ZN(P1_U3192) );
  AND2_X1 U23741 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20839), .ZN(P1_U3193) );
  AND2_X1 U23742 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20840), .ZN(n20852) );
  INV_X1 U23743 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21035) );
  INV_X1 U23744 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20844) );
  OAI22_X1 U23745 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21031), .B1(n20844), 
        .B2(n21063), .ZN(n20841) );
  NOR3_X1 U23746 ( .A1(n20842), .A2(n21035), .A3(n20841), .ZN(n20843) );
  OAI22_X1 U23747 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20852), .B1(n20923), 
        .B2(n20843), .ZN(P1_U3194) );
  NOR2_X1 U23748 ( .A1(n20844), .A2(n20853), .ZN(n20846) );
  NOR2_X1 U23749 ( .A1(n20847), .A2(n21035), .ZN(n20845) );
  OAI22_X1 U23750 ( .A1(n20846), .A2(n21031), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20845), .ZN(n20851) );
  NOR3_X1 U23751 ( .A1(NA), .A2(n20847), .A3(n20918), .ZN(n20848) );
  OAI22_X1 U23752 ( .A1(n20849), .A2(n20848), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n21035), .ZN(n20850) );
  OAI22_X1 U23753 ( .A1(n20852), .A2(n20851), .B1(n21063), .B2(n20850), .ZN(
        P1_U3196) );
  OR2_X1 U23754 ( .A1(n20853), .A2(n20899), .ZN(n20892) );
  NAND2_X1 U23755 ( .A1(n20853), .A2(n20923), .ZN(n20895) );
  INV_X1 U23756 ( .A(n20895), .ZN(n20890) );
  AOI22_X1 U23757 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n20899), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20890), .ZN(n20854) );
  OAI21_X1 U23758 ( .B1(n20855), .B2(n20892), .A(n20854), .ZN(P1_U3197) );
  INV_X1 U23759 ( .A(n20892), .ZN(n20893) );
  AOI22_X1 U23760 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20899), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20893), .ZN(n20856) );
  OAI21_X1 U23761 ( .B1(n20859), .B2(n20895), .A(n20856), .ZN(P1_U3198) );
  OAI222_X1 U23762 ( .A1(n20892), .A2(n20859), .B1(n20858), .B2(n20923), .C1(
        n20857), .C2(n20895), .ZN(P1_U3199) );
  INV_X1 U23763 ( .A(n20923), .ZN(n20922) );
  AOI222_X1 U23764 ( .A1(n20890), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20893), .ZN(n20860) );
  INV_X1 U23765 ( .A(n20860), .ZN(P1_U3200) );
  AOI22_X1 U23766 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n20899), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n20890), .ZN(n20861) );
  OAI21_X1 U23767 ( .B1(n20862), .B2(n20892), .A(n20861), .ZN(P1_U3201) );
  INV_X1 U23768 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20864) );
  AOI22_X1 U23769 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20899), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20890), .ZN(n20863) );
  OAI21_X1 U23770 ( .B1(n20864), .B2(n20892), .A(n20863), .ZN(P1_U3202) );
  AOI22_X1 U23771 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20899), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20893), .ZN(n20865) );
  OAI21_X1 U23772 ( .B1(n20866), .B2(n20895), .A(n20865), .ZN(P1_U3203) );
  AOI222_X1 U23773 ( .A1(n20890), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20893), .ZN(n20867) );
  INV_X1 U23774 ( .A(n20867), .ZN(P1_U3204) );
  AOI222_X1 U23775 ( .A1(n20893), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20890), .ZN(n20868) );
  INV_X1 U23776 ( .A(n20868), .ZN(P1_U3205) );
  AOI222_X1 U23777 ( .A1(n20893), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20890), .ZN(n20869) );
  INV_X1 U23778 ( .A(n20869), .ZN(P1_U3206) );
  AOI222_X1 U23779 ( .A1(n20893), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20890), .ZN(n20870) );
  INV_X1 U23780 ( .A(n20870), .ZN(P1_U3207) );
  AOI222_X1 U23781 ( .A1(n20893), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20890), .ZN(n20871) );
  INV_X1 U23782 ( .A(n20871), .ZN(P1_U3208) );
  AOI22_X1 U23783 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20899), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20890), .ZN(n20872) );
  OAI21_X1 U23784 ( .B1(n20873), .B2(n20892), .A(n20872), .ZN(P1_U3209) );
  AOI22_X1 U23785 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20899), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20893), .ZN(n20874) );
  OAI21_X1 U23786 ( .B1(n20875), .B2(n20895), .A(n20874), .ZN(P1_U3210) );
  AOI222_X1 U23787 ( .A1(n20893), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20890), .ZN(n20876) );
  INV_X1 U23788 ( .A(n20876), .ZN(P1_U3211) );
  AOI222_X1 U23789 ( .A1(n20893), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20890), .ZN(n20877) );
  INV_X1 U23790 ( .A(n20877), .ZN(P1_U3212) );
  AOI222_X1 U23791 ( .A1(n20893), .A2(P1_REIP_REG_17__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n20890), .ZN(n20878) );
  INV_X1 U23792 ( .A(n20878), .ZN(P1_U3213) );
  AOI222_X1 U23793 ( .A1(n20893), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20890), .ZN(n20879) );
  INV_X1 U23794 ( .A(n20879), .ZN(P1_U3214) );
  AOI222_X1 U23795 ( .A1(n20893), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n20890), .ZN(n20880) );
  INV_X1 U23796 ( .A(n20880), .ZN(P1_U3215) );
  AOI222_X1 U23797 ( .A1(n20890), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n20893), .ZN(n20881) );
  INV_X1 U23798 ( .A(n20881), .ZN(P1_U3216) );
  AOI222_X1 U23799 ( .A1(n20893), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20890), .ZN(n20882) );
  INV_X1 U23800 ( .A(n20882), .ZN(P1_U3217) );
  AOI222_X1 U23801 ( .A1(n20893), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20890), .ZN(n20883) );
  INV_X1 U23802 ( .A(n20883), .ZN(P1_U3218) );
  AOI222_X1 U23803 ( .A1(n20890), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20893), .ZN(n20884) );
  INV_X1 U23804 ( .A(n20884), .ZN(P1_U3219) );
  AOI222_X1 U23805 ( .A1(n20890), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20893), .ZN(n20885) );
  INV_X1 U23806 ( .A(n20885), .ZN(P1_U3220) );
  AOI222_X1 U23807 ( .A1(n20893), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20890), .ZN(n20886) );
  INV_X1 U23808 ( .A(n20886), .ZN(P1_U3221) );
  AOI222_X1 U23809 ( .A1(n20890), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20893), .ZN(n20887) );
  INV_X1 U23810 ( .A(n20887), .ZN(P1_U3222) );
  AOI222_X1 U23811 ( .A1(n20890), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20893), .ZN(n20888) );
  INV_X1 U23812 ( .A(n20888), .ZN(P1_U3223) );
  AOI222_X1 U23813 ( .A1(n20893), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20922), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20890), .ZN(n20889) );
  INV_X1 U23814 ( .A(n20889), .ZN(P1_U3224) );
  AOI22_X1 U23815 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(n20899), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(n20890), .ZN(n20891) );
  OAI21_X1 U23816 ( .B1(n21052), .B2(n20892), .A(n20891), .ZN(P1_U3225) );
  AOI22_X1 U23817 ( .A1(P1_ADDRESS_REG_29__SCAN_IN), .A2(n20899), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(n20893), .ZN(n20894) );
  OAI21_X1 U23818 ( .B1(n21032), .B2(n20895), .A(n20894), .ZN(P1_U3226) );
  OAI22_X1 U23819 ( .A1(n20922), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20923), .ZN(n20896) );
  INV_X1 U23820 ( .A(n20896), .ZN(P1_U3458) );
  OAI22_X1 U23821 ( .A1(n20922), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20923), .ZN(n20897) );
  INV_X1 U23822 ( .A(n20897), .ZN(P1_U3459) );
  OAI22_X1 U23823 ( .A1(n20922), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20923), .ZN(n20898) );
  INV_X1 U23824 ( .A(n20898), .ZN(P1_U3460) );
  OAI22_X1 U23825 ( .A1(n20899), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20923), .ZN(n20900) );
  INV_X1 U23826 ( .A(n20900), .ZN(P1_U3461) );
  OAI21_X1 U23827 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20904), .A(n20902), 
        .ZN(n20901) );
  INV_X1 U23828 ( .A(n20901), .ZN(P1_U3464) );
  OAI21_X1 U23829 ( .B1(n20904), .B2(n20903), .A(n20902), .ZN(P1_U3465) );
  AOI211_X1 U23830 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_REIP_REG_1__SCAN_IN), .B(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20905) );
  AOI21_X1 U23831 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20905), .ZN(n20906) );
  INV_X1 U23832 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21053) );
  AOI22_X1 U23833 ( .A1(n20909), .A2(n20906), .B1(n21053), .B2(n20907), .ZN(
        P1_U3481) );
  NOR2_X1 U23834 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20908) );
  INV_X1 U23835 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20941) );
  AOI22_X1 U23836 ( .A1(n20909), .A2(n20908), .B1(n20941), .B2(n20907), .ZN(
        P1_U3482) );
  AOI22_X1 U23837 ( .A1(n20923), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21028), 
        .B2(n20922), .ZN(P1_U3483) );
  NAND2_X1 U23838 ( .A1(n20910), .A2(n21034), .ZN(n20911) );
  AND4_X1 U23839 ( .A1(n20912), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n20918), 
        .A4(n20911), .ZN(n20915) );
  OAI21_X1 U23840 ( .B1(n20915), .B2(n20914), .A(n20913), .ZN(n20921) );
  AOI211_X1 U23841 ( .C1(n20919), .C2(n20918), .A(n20917), .B(n20916), .ZN(
        n20920) );
  MUX2_X1 U23842 ( .A(n20921), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20920), 
        .Z(P1_U3485) );
  INV_X1 U23843 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n20957) );
  AOI22_X1 U23844 ( .A1(n20923), .A2(n20957), .B1(n20979), .B2(n20922), .ZN(
        P1_U3486) );
  INV_X1 U23845 ( .A(keyinput_f24), .ZN(n21012) );
  AOI22_X1 U23846 ( .A1(n13250), .A2(keyinput_f17), .B1(keyinput_f47), .B2(
        n21028), .ZN(n20924) );
  OAI221_X1 U23847 ( .B1(n13250), .B2(keyinput_f17), .C1(n21028), .C2(
        keyinput_f47), .A(n20924), .ZN(n21010) );
  AOI22_X1 U23848 ( .A1(n21059), .A2(keyinput_f61), .B1(keyinput_f22), .B2(
        n21087), .ZN(n20925) );
  OAI221_X1 U23849 ( .B1(n21059), .B2(keyinput_f61), .C1(n21087), .C2(
        keyinput_f22), .A(n20925), .ZN(n21009) );
  INV_X1 U23850 ( .A(DATAI_23_), .ZN(n20927) );
  OAI22_X1 U23851 ( .A1(n20928), .A2(keyinput_f3), .B1(n20927), .B2(
        keyinput_f9), .ZN(n20926) );
  AOI221_X1 U23852 ( .B1(n20928), .B2(keyinput_f3), .C1(keyinput_f9), .C2(
        n20927), .A(n20926), .ZN(n20945) );
  AOI22_X1 U23853 ( .A1(n13405), .A2(keyinput_f28), .B1(n20930), .B2(
        keyinput_f10), .ZN(n20929) );
  OAI221_X1 U23854 ( .B1(n13405), .B2(keyinput_f28), .C1(n20930), .C2(
        keyinput_f10), .A(n20929), .ZN(n20940) );
  AOI22_X1 U23855 ( .A1(n13401), .A2(keyinput_f27), .B1(keyinput_f15), .B2(
        n20932), .ZN(n20931) );
  OAI221_X1 U23856 ( .B1(n13401), .B2(keyinput_f27), .C1(n20932), .C2(
        keyinput_f15), .A(n20931), .ZN(n20939) );
  INV_X1 U23857 ( .A(READY1), .ZN(n20934) );
  AOI22_X1 U23858 ( .A1(n20934), .A2(keyinput_f36), .B1(keyinput_f54), .B2(
        n21052), .ZN(n20933) );
  OAI221_X1 U23859 ( .B1(n20934), .B2(keyinput_f36), .C1(n21052), .C2(
        keyinput_f54), .A(n20933), .ZN(n20938) );
  AOI22_X1 U23860 ( .A1(n21037), .A2(keyinput_f4), .B1(keyinput_f6), .B2(
        n20936), .ZN(n20935) );
  OAI221_X1 U23861 ( .B1(n21037), .B2(keyinput_f4), .C1(n20936), .C2(
        keyinput_f6), .A(n20935), .ZN(n20937) );
  NOR4_X1 U23862 ( .A1(n20940), .A2(n20939), .A3(n20938), .A4(n20937), .ZN(
        n20944) );
  XOR2_X1 U23863 ( .A(keyinput_f48), .B(n20941), .Z(n20943) );
  XOR2_X1 U23864 ( .A(keyinput_f50), .B(n21053), .Z(n20942) );
  NAND4_X1 U23865 ( .A1(n20945), .A2(n20944), .A3(n20943), .A4(n20942), .ZN(
        n21008) );
  OAI22_X1 U23866 ( .A1(DATAI_11_), .A2(keyinput_f21), .B1(
        P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_f40), .ZN(n20946) );
  AOI221_X1 U23867 ( .B1(DATAI_11_), .B2(keyinput_f21), .C1(keyinput_f40), 
        .C2(P1_CODEFETCH_REG_SCAN_IN), .A(n20946), .ZN(n21006) );
  OAI22_X1 U23868 ( .A1(DATAI_9_), .A2(keyinput_f23), .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_f42), .ZN(n20947) );
  AOI221_X1 U23869 ( .B1(DATAI_9_), .B2(keyinput_f23), .C1(keyinput_f42), .C2(
        P1_D_C_N_REG_SCAN_IN), .A(n20947), .ZN(n21005) );
  AOI22_X1 U23870 ( .A1(DATAI_16_), .A2(keyinput_f16), .B1(DATAI_6_), .B2(
        keyinput_f26), .ZN(n20948) );
  OAI221_X1 U23871 ( .B1(DATAI_16_), .B2(keyinput_f16), .C1(DATAI_6_), .C2(
        keyinput_f26), .A(n20948), .ZN(n20955) );
  AOI22_X1 U23872 ( .A1(DATAI_30_), .A2(keyinput_f2), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(keyinput_f53), .ZN(n20949) );
  OAI221_X1 U23873 ( .B1(DATAI_30_), .B2(keyinput_f2), .C1(
        P1_REIP_REG_30__SCAN_IN), .C2(keyinput_f53), .A(n20949), .ZN(n20954)
         );
  AOI22_X1 U23874 ( .A1(DATAI_14_), .A2(keyinput_f18), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(keyinput_f60), .ZN(n20950) );
  OAI221_X1 U23875 ( .B1(DATAI_14_), .B2(keyinput_f18), .C1(
        P1_REIP_REG_23__SCAN_IN), .C2(keyinput_f60), .A(n20950), .ZN(n20953)
         );
  AOI22_X1 U23876 ( .A1(keyinput_f34), .A2(NA), .B1(DATAI_24_), .B2(
        keyinput_f8), .ZN(n20951) );
  OAI221_X1 U23877 ( .B1(keyinput_f34), .B2(NA), .C1(DATAI_24_), .C2(
        keyinput_f8), .A(n20951), .ZN(n20952) );
  NOR4_X1 U23878 ( .A1(n20955), .A2(n20954), .A3(n20953), .A4(n20952), .ZN(
        n20959) );
  OAI22_X1 U23879 ( .A1(n20957), .A2(keyinput_f0), .B1(keyinput_f11), .B2(
        DATAI_21_), .ZN(n20956) );
  AOI221_X1 U23880 ( .B1(n20957), .B2(keyinput_f0), .C1(DATAI_21_), .C2(
        keyinput_f11), .A(n20956), .ZN(n20958) );
  OAI211_X1 U23881 ( .C1(DATAI_12_), .C2(keyinput_f20), .A(n20959), .B(n20958), 
        .ZN(n20960) );
  AOI21_X1 U23882 ( .B1(DATAI_12_), .B2(keyinput_f20), .A(n20960), .ZN(n21004)
         );
  OAI22_X1 U23883 ( .A1(DATAI_31_), .A2(keyinput_f1), .B1(keyinput_f32), .B2(
        DATAI_0_), .ZN(n20961) );
  AOI221_X1 U23884 ( .B1(DATAI_31_), .B2(keyinput_f1), .C1(DATAI_0_), .C2(
        keyinput_f32), .A(n20961), .ZN(n20969) );
  OAI22_X1 U23885 ( .A1(DATAI_2_), .A2(keyinput_f30), .B1(READY2), .B2(
        keyinput_f37), .ZN(n20962) );
  AOI221_X1 U23886 ( .B1(DATAI_2_), .B2(keyinput_f30), .C1(keyinput_f37), .C2(
        READY2), .A(n20962), .ZN(n20968) );
  INV_X1 U23887 ( .A(DATAI_3_), .ZN(n20964) );
  OAI22_X1 U23888 ( .A1(n20964), .A2(keyinput_f29), .B1(n21015), .B2(
        keyinput_f51), .ZN(n20963) );
  AOI221_X1 U23889 ( .B1(n20964), .B2(keyinput_f29), .C1(keyinput_f51), .C2(
        n21015), .A(n20963), .ZN(n20967) );
  OAI22_X1 U23890 ( .A1(n21035), .A2(keyinput_f43), .B1(keyinput_f12), .B2(
        DATAI_20_), .ZN(n20965) );
  AOI221_X1 U23891 ( .B1(n21035), .B2(keyinput_f43), .C1(DATAI_20_), .C2(
        keyinput_f12), .A(n20965), .ZN(n20966) );
  NAND4_X1 U23892 ( .A1(n20969), .A2(n20968), .A3(n20967), .A4(n20966), .ZN(
        n21002) );
  OAI22_X1 U23893 ( .A1(DATAI_7_), .A2(keyinput_f25), .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_f46), .ZN(n20970) );
  AOI221_X1 U23894 ( .B1(DATAI_7_), .B2(keyinput_f25), .C1(keyinput_f46), .C2(
        P1_FLUSH_REG_SCAN_IN), .A(n20970), .ZN(n20977) );
  OAI22_X1 U23895 ( .A1(P1_REIP_REG_31__SCAN_IN), .A2(keyinput_f52), .B1(
        keyinput_f5), .B2(DATAI_27_), .ZN(n20971) );
  AOI221_X1 U23896 ( .B1(P1_REIP_REG_31__SCAN_IN), .B2(keyinput_f52), .C1(
        DATAI_27_), .C2(keyinput_f5), .A(n20971), .ZN(n20976) );
  OAI22_X1 U23897 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(keyinput_f59), .B1(
        P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_f38), .ZN(n20972) );
  AOI221_X1 U23898 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(keyinput_f59), .C1(
        keyinput_f38), .C2(P1_READREQUEST_REG_SCAN_IN), .A(n20972), .ZN(n20975) );
  OAI22_X1 U23899 ( .A1(DATAI_25_), .A2(keyinput_f7), .B1(keyinput_f45), .B2(
        P1_MORE_REG_SCAN_IN), .ZN(n20973) );
  AOI221_X1 U23900 ( .B1(DATAI_25_), .B2(keyinput_f7), .C1(P1_MORE_REG_SCAN_IN), .C2(keyinput_f45), .A(n20973), .ZN(n20974) );
  NAND4_X1 U23901 ( .A1(n20977), .A2(n20976), .A3(n20975), .A4(n20974), .ZN(
        n21001) );
  OAI22_X1 U23902 ( .A1(n21019), .A2(keyinput_f57), .B1(n20979), .B2(
        keyinput_f41), .ZN(n20978) );
  AOI221_X1 U23903 ( .B1(n21019), .B2(keyinput_f57), .C1(keyinput_f41), .C2(
        n20979), .A(n20978), .ZN(n20989) );
  INV_X1 U23904 ( .A(DATAI_18_), .ZN(n21021) );
  INV_X1 U23905 ( .A(keyinput_f39), .ZN(n20981) );
  OAI22_X1 U23906 ( .A1(n21021), .A2(keyinput_f14), .B1(n20981), .B2(
        P1_ADS_N_REG_SCAN_IN), .ZN(n20980) );
  AOI221_X1 U23907 ( .B1(n21021), .B2(keyinput_f14), .C1(P1_ADS_N_REG_SCAN_IN), 
        .C2(n20981), .A(n20980), .ZN(n20988) );
  INV_X1 U23908 ( .A(DATAI_19_), .ZN(n20983) );
  OAI22_X1 U23909 ( .A1(n14897), .A2(keyinput_f58), .B1(n20983), .B2(
        keyinput_f13), .ZN(n20982) );
  AOI221_X1 U23910 ( .B1(n14897), .B2(keyinput_f58), .C1(keyinput_f13), .C2(
        n20983), .A(n20982), .ZN(n20987) );
  OAI22_X1 U23911 ( .A1(n20985), .A2(keyinput_f63), .B1(n21029), .B2(
        keyinput_f35), .ZN(n20984) );
  AOI221_X1 U23912 ( .B1(n20985), .B2(keyinput_f63), .C1(keyinput_f35), .C2(
        n21029), .A(n20984), .ZN(n20986) );
  NAND4_X1 U23913 ( .A1(n20989), .A2(n20988), .A3(n20987), .A4(n20986), .ZN(
        n21000) );
  OAI22_X1 U23914 ( .A1(n21034), .A2(keyinput_f44), .B1(n21065), .B2(
        keyinput_f55), .ZN(n20990) );
  AOI221_X1 U23915 ( .B1(n21034), .B2(keyinput_f44), .C1(keyinput_f55), .C2(
        n21065), .A(n20990), .ZN(n20998) );
  INV_X1 U23916 ( .A(DATAI_1_), .ZN(n21022) );
  OAI22_X1 U23917 ( .A1(n21060), .A2(keyinput_f56), .B1(n21022), .B2(
        keyinput_f31), .ZN(n20991) );
  AOI221_X1 U23918 ( .B1(n21060), .B2(keyinput_f56), .C1(keyinput_f31), .C2(
        n21022), .A(n20991), .ZN(n20997) );
  OAI22_X1 U23919 ( .A1(n21050), .A2(keyinput_f19), .B1(n21068), .B2(
        keyinput_f49), .ZN(n20992) );
  AOI221_X1 U23920 ( .B1(n21050), .B2(keyinput_f19), .C1(keyinput_f49), .C2(
        n21068), .A(n20992), .ZN(n20996) );
  OAI22_X1 U23921 ( .A1(n20994), .A2(keyinput_f62), .B1(n21063), .B2(
        keyinput_f33), .ZN(n20993) );
  AOI221_X1 U23922 ( .B1(n20994), .B2(keyinput_f62), .C1(keyinput_f33), .C2(
        n21063), .A(n20993), .ZN(n20995) );
  NAND4_X1 U23923 ( .A1(n20998), .A2(n20997), .A3(n20996), .A4(n20995), .ZN(
        n20999) );
  NOR4_X1 U23924 ( .A1(n21002), .A2(n21001), .A3(n21000), .A4(n20999), .ZN(
        n21003) );
  NAND4_X1 U23925 ( .A1(n21006), .A2(n21005), .A3(n21004), .A4(n21003), .ZN(
        n21007) );
  NOR4_X1 U23926 ( .A1(n21010), .A2(n21009), .A3(n21008), .A4(n21007), .ZN(
        n21011) );
  AOI221_X1 U23927 ( .B1(DATAI_8_), .B2(n21012), .C1(n21119), .C2(keyinput_f24), .A(n21011), .ZN(n21118) );
  AOI22_X1 U23928 ( .A1(n21015), .A2(keyinput_g51), .B1(n21014), .B2(
        keyinput_g5), .ZN(n21013) );
  OAI221_X1 U23929 ( .B1(n21015), .B2(keyinput_g51), .C1(n21014), .C2(
        keyinput_g5), .A(n21013), .ZN(n21026) );
  AOI22_X1 U23930 ( .A1(n21017), .A2(keyinput_g23), .B1(n14897), .B2(
        keyinput_g58), .ZN(n21016) );
  OAI221_X1 U23931 ( .B1(n21017), .B2(keyinput_g23), .C1(n14897), .C2(
        keyinput_g58), .A(n21016), .ZN(n21025) );
  AOI22_X1 U23932 ( .A1(n13401), .A2(keyinput_g27), .B1(n21019), .B2(
        keyinput_g57), .ZN(n21018) );
  OAI221_X1 U23933 ( .B1(n13401), .B2(keyinput_g27), .C1(n21019), .C2(
        keyinput_g57), .A(n21018), .ZN(n21024) );
  AOI22_X1 U23934 ( .A1(n21022), .A2(keyinput_g31), .B1(n21021), .B2(
        keyinput_g14), .ZN(n21020) );
  OAI221_X1 U23935 ( .B1(n21022), .B2(keyinput_g31), .C1(n21021), .C2(
        keyinput_g14), .A(n21020), .ZN(n21023) );
  NOR4_X1 U23936 ( .A1(n21026), .A2(n21025), .A3(n21024), .A4(n21023), .ZN(
        n21077) );
  AOI22_X1 U23937 ( .A1(n21029), .A2(keyinput_g35), .B1(n21028), .B2(
        keyinput_g47), .ZN(n21027) );
  OAI221_X1 U23938 ( .B1(n21029), .B2(keyinput_g35), .C1(n21028), .C2(
        keyinput_g47), .A(n21027), .ZN(n21042) );
  AOI22_X1 U23939 ( .A1(n21032), .A2(keyinput_g52), .B1(keyinput_g34), .B2(
        n21031), .ZN(n21030) );
  OAI221_X1 U23940 ( .B1(n21032), .B2(keyinput_g52), .C1(n21031), .C2(
        keyinput_g34), .A(n21030), .ZN(n21041) );
  AOI22_X1 U23941 ( .A1(n21035), .A2(keyinput_g43), .B1(n21034), .B2(
        keyinput_g44), .ZN(n21033) );
  OAI221_X1 U23942 ( .B1(n21035), .B2(keyinput_g43), .C1(n21034), .C2(
        keyinput_g44), .A(n21033), .ZN(n21040) );
  AOI22_X1 U23943 ( .A1(n21038), .A2(keyinput_g1), .B1(keyinput_g4), .B2(
        n21037), .ZN(n21036) );
  OAI221_X1 U23944 ( .B1(n21038), .B2(keyinput_g1), .C1(n21037), .C2(
        keyinput_g4), .A(n21036), .ZN(n21039) );
  NOR4_X1 U23945 ( .A1(n21042), .A2(n21041), .A3(n21040), .A4(n21039), .ZN(
        n21076) );
  INV_X1 U23946 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n21045) );
  AOI22_X1 U23947 ( .A1(n21045), .A2(keyinput_g38), .B1(keyinput_g40), .B2(
        n21044), .ZN(n21043) );
  OAI221_X1 U23948 ( .B1(n21045), .B2(keyinput_g38), .C1(n21044), .C2(
        keyinput_g40), .A(n21043), .ZN(n21057) );
  INV_X1 U23949 ( .A(DATAI_21_), .ZN(n21048) );
  AOI22_X1 U23950 ( .A1(n21048), .A2(keyinput_g11), .B1(n21047), .B2(
        keyinput_g21), .ZN(n21046) );
  OAI221_X1 U23951 ( .B1(n21048), .B2(keyinput_g11), .C1(n21047), .C2(
        keyinput_g21), .A(n21046), .ZN(n21056) );
  AOI22_X1 U23952 ( .A1(n13405), .A2(keyinput_g28), .B1(n21050), .B2(
        keyinput_g19), .ZN(n21049) );
  OAI221_X1 U23953 ( .B1(n13405), .B2(keyinput_g28), .C1(n21050), .C2(
        keyinput_g19), .A(n21049), .ZN(n21055) );
  AOI22_X1 U23954 ( .A1(n21053), .A2(keyinput_g50), .B1(n21052), .B2(
        keyinput_g54), .ZN(n21051) );
  OAI221_X1 U23955 ( .B1(n21053), .B2(keyinput_g50), .C1(n21052), .C2(
        keyinput_g54), .A(n21051), .ZN(n21054) );
  NOR4_X1 U23956 ( .A1(n21057), .A2(n21056), .A3(n21055), .A4(n21054), .ZN(
        n21075) );
  AOI22_X1 U23957 ( .A1(n21060), .A2(keyinput_g56), .B1(n21059), .B2(
        keyinput_g61), .ZN(n21058) );
  OAI221_X1 U23958 ( .B1(n21060), .B2(keyinput_g56), .C1(n21059), .C2(
        keyinput_g61), .A(n21058), .ZN(n21073) );
  AOI22_X1 U23959 ( .A1(n21063), .A2(keyinput_g33), .B1(n21062), .B2(
        keyinput_g20), .ZN(n21061) );
  OAI221_X1 U23960 ( .B1(n21063), .B2(keyinput_g33), .C1(n21062), .C2(
        keyinput_g20), .A(n21061), .ZN(n21072) );
  INV_X1 U23961 ( .A(DATAI_20_), .ZN(n21066) );
  AOI22_X1 U23962 ( .A1(n21066), .A2(keyinput_g12), .B1(n21065), .B2(
        keyinput_g55), .ZN(n21064) );
  OAI221_X1 U23963 ( .B1(n21066), .B2(keyinput_g12), .C1(n21065), .C2(
        keyinput_g55), .A(n21064), .ZN(n21071) );
  AOI22_X1 U23964 ( .A1(n21069), .A2(keyinput_g45), .B1(keyinput_g49), .B2(
        n21068), .ZN(n21067) );
  OAI221_X1 U23965 ( .B1(n21069), .B2(keyinput_g45), .C1(n21068), .C2(
        keyinput_g49), .A(n21067), .ZN(n21070) );
  NOR4_X1 U23966 ( .A1(n21073), .A2(n21072), .A3(n21071), .A4(n21070), .ZN(
        n21074) );
  NAND4_X1 U23967 ( .A1(n21077), .A2(n21076), .A3(n21075), .A4(n21074), .ZN(
        n21116) );
  AOI22_X1 U23968 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(keyinput_g46), .B1(
        DATAI_17_), .B2(keyinput_g15), .ZN(n21078) );
  OAI221_X1 U23969 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_g46), .C1(
        DATAI_17_), .C2(keyinput_g15), .A(n21078), .ZN(n21085) );
  AOI22_X1 U23970 ( .A1(DATAI_0_), .A2(keyinput_g32), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(keyinput_g53), .ZN(n21079) );
  OAI221_X1 U23971 ( .B1(DATAI_0_), .B2(keyinput_g32), .C1(
        P1_REIP_REG_30__SCAN_IN), .C2(keyinput_g53), .A(n21079), .ZN(n21084)
         );
  AOI22_X1 U23972 ( .A1(DATAI_26_), .A2(keyinput_g6), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(keyinput_g60), .ZN(n21080) );
  OAI221_X1 U23973 ( .B1(DATAI_26_), .B2(keyinput_g6), .C1(
        P1_REIP_REG_23__SCAN_IN), .C2(keyinput_g60), .A(n21080), .ZN(n21083)
         );
  AOI22_X1 U23974 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(keyinput_g39), .B1(DATAI_7_), .B2(keyinput_g25), .ZN(n21081) );
  OAI221_X1 U23975 ( .B1(P1_ADS_N_REG_SCAN_IN), .B2(keyinput_g39), .C1(
        DATAI_7_), .C2(keyinput_g25), .A(n21081), .ZN(n21082) );
  NOR4_X1 U23976 ( .A1(n21085), .A2(n21084), .A3(n21083), .A4(n21082), .ZN(
        n21114) );
  XNOR2_X1 U23977 ( .A(DATAI_2_), .B(keyinput_g30), .ZN(n21093) );
  AOI22_X1 U23978 ( .A1(DATAI_3_), .A2(keyinput_g29), .B1(n21087), .B2(
        keyinput_g22), .ZN(n21086) );
  OAI221_X1 U23979 ( .B1(DATAI_3_), .B2(keyinput_g29), .C1(n21087), .C2(
        keyinput_g22), .A(n21086), .ZN(n21092) );
  AOI22_X1 U23980 ( .A1(P1_BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_g48), .B1(
        DATAI_23_), .B2(keyinput_g9), .ZN(n21088) );
  OAI221_X1 U23981 ( .B1(P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_g48), 
        .C1(DATAI_23_), .C2(keyinput_g9), .A(n21088), .ZN(n21091) );
  AOI22_X1 U23982 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(keyinput_g59), .ZN(n21089) );
  OAI221_X1 U23983 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        P1_REIP_REG_24__SCAN_IN), .C2(keyinput_g59), .A(n21089), .ZN(n21090)
         );
  NOR4_X1 U23984 ( .A1(n21093), .A2(n21092), .A3(n21091), .A4(n21090), .ZN(
        n21113) );
  AOI22_X1 U23985 ( .A1(DATAI_14_), .A2(keyinput_g18), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(keyinput_g63), .ZN(n21094) );
  OAI221_X1 U23986 ( .B1(DATAI_14_), .B2(keyinput_g18), .C1(
        P1_REIP_REG_20__SCAN_IN), .C2(keyinput_g63), .A(n21094), .ZN(n21102)
         );
  AOI22_X1 U23987 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(keyinput_g42), .B1(
        DATAI_30_), .B2(keyinput_g2), .ZN(n21095) );
  OAI221_X1 U23988 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_g42), .C1(
        DATAI_30_), .C2(keyinput_g2), .A(n21095), .ZN(n21101) );
  INV_X1 U23989 ( .A(DATAI_25_), .ZN(n21097) );
  AOI22_X1 U23990 ( .A1(DATAI_29_), .A2(keyinput_g3), .B1(n21097), .B2(
        keyinput_g7), .ZN(n21096) );
  OAI221_X1 U23991 ( .B1(DATAI_29_), .B2(keyinput_g3), .C1(n21097), .C2(
        keyinput_g7), .A(n21096), .ZN(n21100) );
  AOI22_X1 U23992 ( .A1(DATAI_16_), .A2(keyinput_g16), .B1(DATAI_6_), .B2(
        keyinput_g26), .ZN(n21098) );
  OAI221_X1 U23993 ( .B1(DATAI_16_), .B2(keyinput_g16), .C1(DATAI_6_), .C2(
        keyinput_g26), .A(n21098), .ZN(n21099) );
  NOR4_X1 U23994 ( .A1(n21102), .A2(n21101), .A3(n21100), .A4(n21099), .ZN(
        n21112) );
  AOI22_X1 U23995 ( .A1(DATAI_22_), .A2(keyinput_g10), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(keyinput_g62), .ZN(n21103) );
  OAI221_X1 U23996 ( .B1(DATAI_22_), .B2(keyinput_g10), .C1(
        P1_REIP_REG_21__SCAN_IN), .C2(keyinput_g62), .A(n21103), .ZN(n21110)
         );
  AOI22_X1 U23997 ( .A1(DATAI_24_), .A2(keyinput_g8), .B1(READY1), .B2(
        keyinput_g36), .ZN(n21104) );
  OAI221_X1 U23998 ( .B1(DATAI_24_), .B2(keyinput_g8), .C1(READY1), .C2(
        keyinput_g36), .A(n21104), .ZN(n21109) );
  AOI22_X1 U23999 ( .A1(P1_M_IO_N_REG_SCAN_IN), .A2(keyinput_g41), .B1(
        DATAI_19_), .B2(keyinput_g13), .ZN(n21105) );
  OAI221_X1 U24000 ( .B1(P1_M_IO_N_REG_SCAN_IN), .B2(keyinput_g41), .C1(
        DATAI_19_), .C2(keyinput_g13), .A(n21105), .ZN(n21108) );
  AOI22_X1 U24001 ( .A1(DATAI_15_), .A2(keyinput_g17), .B1(READY2), .B2(
        keyinput_g37), .ZN(n21106) );
  OAI221_X1 U24002 ( .B1(DATAI_15_), .B2(keyinput_g17), .C1(READY2), .C2(
        keyinput_g37), .A(n21106), .ZN(n21107) );
  NOR4_X1 U24003 ( .A1(n21110), .A2(n21109), .A3(n21108), .A4(n21107), .ZN(
        n21111) );
  NAND4_X1 U24004 ( .A1(n21114), .A2(n21113), .A3(n21112), .A4(n21111), .ZN(
        n21115) );
  OAI22_X1 U24005 ( .A1(keyinput_g24), .A2(n21119), .B1(n21116), .B2(n21115), 
        .ZN(n21117) );
  AOI211_X1 U24006 ( .C1(keyinput_g24), .C2(n21119), .A(n21118), .B(n21117), 
        .ZN(n21121) );
  AOI22_X1 U24007 ( .A1(n16543), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16545), .ZN(n21120) );
  XNOR2_X1 U24008 ( .A(n21121), .B(n21120), .ZN(U355) );
  AND2_X1 U11487 ( .A1(n10193), .A2(n15163), .ZN(n10836) );
  NAND2_X1 U14171 ( .A1(n11312), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14290) );
  NAND4_X1 U11160 ( .A1(n11452), .A2(n11461), .A3(n11460), .A4(n11459), .ZN(
        n11471) );
  INV_X1 U11472 ( .A(n11496), .ZN(n11502) );
  NOR2_X1 U12742 ( .A1(n12833), .A2(n12834), .ZN(n14153) );
  INV_X1 U11480 ( .A(n11330), .ZN(n9648) );
  NAND2_X1 U14325 ( .A1(n11399), .A2(n11381), .ZN(n11397) );
  AND2_X2 U12499 ( .A1(n11367), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11625) );
  INV_X2 U11099 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16338) );
  AND2_X2 U11125 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11221) );
  CLKBUF_X1 U11129 ( .A(n11428), .Z(n16386) );
  CLKBUF_X1 U11130 ( .A(n20064), .Z(n20225) );
  CLKBUF_X1 U11191 ( .A(n15780), .Z(n9646) );
  CLKBUF_X1 U11242 ( .A(n11426), .Z(n12811) );
  CLKBUF_X1 U11247 ( .A(n11683), .Z(n11790) );
  CLKBUF_X1 U11410 ( .A(n13089), .Z(n19982) );
  CLKBUF_X1 U11470 ( .A(n17905), .Z(n9659) );
  CLKBUF_X1 U11502 ( .A(n10427), .Z(n20837) );
  CLKBUF_X1 U11503 ( .A(n17540), .Z(n17549) );
endmodule

